
module global_region (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
