
module dual_region (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
