`ifndef GENCORES_SIM_DEFS_SV
 `define GENCORES_SIM_DEFS_SV 1

typedef byte unsigned uint8_t;
typedef longint unsigned uint64_t;
typedef int unsigned uint32_t;
typedef shortint unsigned uint16_t;

typedef uint64_t u64_vector_t[$];
typedef uint32_t u32_vector_t[$];
typedef uint16_t u16_vector_t[$];
typedef byte u8_vector_t[$];

`endif
