`ifndef SIMDRV_DEFS_SV
 `define SIMDRV_DEFS_SV 1

`include "gencores_sim_defs.svh"

import gencores_sim_pkg::*;

`endif