// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gotGNDsNDrzpLsTY6uFyGlU3sOCQyNUzFCF+D1jsW3QNZSe30hCgXY6XQWkC93rU
lHihKGcGmXz3izmBFo2fNMMzyzqnGerA/IGJkuQxODaMDfO+GR9K/sQMTQBQWBNT
DDvd6IhQM9zWfXMz9QAg4Q13nvjAoYXHKb1kF8i8u6A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70016)
wp7+5sRWYoBUuWQuZ8cIfVdzP/Aei9pctafTd6jsQ1g/NLCnowuFTqaPTOQNdabQ
7z+z82yqnqpEv6ccV2L4aUhABnR0pyL18ttnc2uhboxGRiPkYnGKMjoG2T93BIkR
t2K4eNntsoSYon8fI8dKd+6FTJfXEUHsG+F/WsBGRCtoIyFVL1rwkyN6oxRiEGJ/
160TmnQ6gles6PrONRt9sOukkBbcGk19Cphf4uD0AephS2vQIrgb6pbuRhsVmCDx
Voo+xXp2wyfS571YRqPHIJirx3hzEUiP6+B1g4bWljf/0NAdpUYcErjAZArVtPoj
awfVly0fGcCWIBmru/CkYTZMCwIzmjjWR1iI1h0BUiOKSbP1OUnqQ9sHV+HK0Zc7
VqGi7zMTFO9A9rPVXRpv3uXSOJSyyjKLoFAWnzoMuWw8wbqjCW59cqRnALxLJMpO
Ddgbm0MlO5tCplfpfZpI0Y81wVq/URJZIffBWnVuEklxdWMd87ch1krkSfnF65jn
HvQckaa13Tq49f0CyXLpTFmVbj9i1Bvuh1C41+Z9MCs4q6TJRBdLAID+a9XcZcT+
JRtdudflHtnl1EtH9KmEa7sZ3L8GqvKOJKFNmfkIF+CCLUv+erS6uVP0O0Y/XSCP
JJeVWyPIjeEhz7z19wpcxxE2cyT35rSjiMCWxVTdJJ3fvds199R+OHZIkxtlQde4
TEsJG2FRDqD/N5m85Ez1e1/tciZsveK4dER7TsWFTEQwg2kElGQ/OSe9kmoFbJmG
WSd25MCcP5UfXeFZDCFHo77dlp7WrCm92r8RUX8jcqE/aPbv9En1rB+7SUiJtVGH
Y66N3YO1tLrzhkn0aDrSpAEVMboxww4fRkqZUpOPkZnkxBQXSh4tLJvB5Lmz0Zc6
Ugoszvt5XRuTZmwdMLKLeOBzVNnkt2vX7lQOh/rwovou4I/6Ne9rG6+S2Z6uFMza
fk04UU0lWYJKU/YP5EpJOvjwse9QyMH/AYEPs0KeHiyrWoQjiyM7QtR/KndnCmZ0
6vSh94xbzkrAJikidypXbg5tIKJTR/w+gtEv96gg9gkHP3CJCisj0xMMgVIxBTXD
Ptoa1NnrfB8XW9VanOys6jHiMaAytv+P4mLuMEZPjHB50OytVIAM52MGq5vUNBy5
5lvdGO0SfXLaelGfEMFqlUm8woWwH9TMHpZdsvvDy2Nq3VfJd+F8T/a1H+V4JzpT
4i5XFQ6h9dsGr2DFcbC2PQZPLjx3do+HXN/VMMRQA9gs510p+xn7CqmTWFyugTfu
TOahZig3qlkcmGzUiswtIE4en/75JLGmKKkE16RaDZLiS1xcTGWHgxlZYwf7ZwVa
8rfRE4DhrwSSeICjFRa6VklO+V0wac8RfbxhCqOCkcPAzIFM8HH4vltVhGbUs3DC
K15Nm4nwfGVzWZ9qMdMxVXCONtSwN5W9yT/Wo8r6iKvaBseKaz47KfrJvlGkID9o
PYlwD6Zc6/Po/vcCFLvYyjiesWPDHMo5pD8V2kjBXFXVw8WCRzkd1DpOekgnYM3k
S5ThVoAwJUNLS4uxUEdV3yzr3v84pJEJpaBcvp8T2HEBGMisqqclMePkpnSUGl1G
He2MtanyxtPXWZs99SMmgV0yilriq2DwnupH3Sqki4QT2a4RIiaTbqDJMYI/EqzR
cQbhZoGkJafUp/52Q4TbJgnoF2gmkVBR+/EDx8oHBydy3jIetiiph6ogEHA7uom4
SA92XgzOY1bhyV+xn6vbsrceXgHDkJZSsaTZgW9Z+KvSvflZQ6IkbPVNr8fZ/bp8
oYKORdMWC6Cc6/LpV1wK/5phwP+7u2jms9LSFhm8AtCSA26Dp0LEslFYHU4YHoRt
Q57PceeA5/4TEVWpJ6+EjDtiVezx1cBxisti+Z6WFeaXzqsvXed8jz8MV9teCyPp
8jqSyQ5zToEyXwxYtPDLVh6w4UvNkRXr39hzWu8AoTP24DXUjHSQeH7Oqn4i9MUn
UrCmhpG6jQx77JUoDwNriJ1RWHxacodIbPTlswyfF9iqVsgaWdOYGRM9eH2tGl89
ELwsIsin5i9FUP8zb+BMq5uecH7oGgO7WT06Ykvu9/e3ENEEzljA38RaqmRFZU0K
ug+k4luY5pzUGC9KNo7/Q2goHu4PHAkeK7oeM311QQMfM7QMRdNmlVu0CTbZ6fdK
ZlMmMBB77oFgFL2+kudLw4KodOXZ6ynctp9If6Cqz//cMmUR9t/agiy7pgxIw/dt
F9MNLkvJ6zPU+wa2p1LGzwhPm6RZCeEEqrdJQgtqGMlmdje2dy4S2w/IfxoKcunF
zF86b4IwH+lOGAki2sL75ZU17aua7fxG+vhrmk1UWzLaqbdRMa7snB80ZQmHPhX7
bbamzI1J9Owa7OTzQpHEq2EXPdKH4D7ctR/W/Ity5rUkLeVjSP2DOmfgyspCaiaT
sBiKJlxKcoaL3wCmSDI8cG3xCtsa56mHK2hx7gFNRDBD1/4eY3qcKZEMi3tL8M12
mkzTpdpsceiaECV1ZP8AT8mm68MpghpThz4QH/CtstZkeH1IOFjTMRN+VicR5Pa1
WwmoQbbSHsOORayHyQDiyoa8CnWHwJE92rKlVOWtaDv4ov19/5/CiFgppjAOAXly
PloEpC1oT36l1RApXOGjBvIjEVaRFLAse5lo+yzK4+MgPzcBqq9cF+eNVKpSET6m
47YUr+euKZv6Ft3pf1R44Rny8ME8xUBRz80FnzPyJbtAcO3lLOoIoQTZ4Hhnek1O
p2s7pfeWdg4OLx76HpDFOZN3Bf7LZtPrWguIOK0tc7VjPny3/fUudAJ9JiVVRGa9
Bap30G0QWLYwfN0pllHYs+Loc8HTs4JqtiAgApJLLxy5RcVuzP2mSTL/6kM9QNYF
TgYBJLM15jeFmd01VzKn8sXD/sfNMOSolzDcXJsRgRPuYh2zxn54eol/TcJcBoNn
1cJRL3rfQX3kn0hSk5Vx8SRRKVwkxX+OTX7NTCJTao3gD3DgWZ5Ok2eKG3C5L8S+
lO1U6ywDRWS96N/JHyvn95dLqxIhaOI0Obhh0851O1XXAQPCkIDp3A7k0Z6T+Tte
fwUUQqcMalEsYxVlIMTB4NXbQMPTpdVuZaXadRKTOtxGF6TGS8/njQ/ZCPGaLBtm
3Lk0Yb3P0YlA9RQcnksgO1ah3Ph4qVCjh4PKll8Q0eMZuAezrG9Lg3yyUMvVkosf
ciaUXOyzvXE7bK3hIZz51ODlsDlhM/vyyjgjh4BsrNgxJxpu+q8DQ1SMCrV3lWLo
K8iY7HR3h+gOayHmn/QekrC57uSAoIEoiOmJaD3+25i0JYiCLFtJ3/sQTRD9xfFp
fTSe3BJFOmCGHUcFlNq1vp2d1V7zIjzpLQyoC/w42O1tsVXKNIamZc+NI/9ZL8R4
09YbuOn4V7yVmrhMgVj3XCs22NyDaZUudhBLAAqDhzyAO/CPQMnsDVh9M1WZ5Mz4
eNnAfFAcQegQ1uFr45TSTKiAb28USf5eBDIWnGjvEMmi1om1ueM18CZoQwTaEQSc
Y4KRdCMU16IkkNkR7GnHRMyPasoqPLyEdCfCgslwxhpYvwRWUJC7EOtOlaReWa6S
LQ+kBLEWlK/WvdrsUqlVpTO++DsKCZNnd1a/F59KV8WsKXWeWPOb+6r/G9yEHuic
pb/ByPxQXz56zlSD+GIjyvuS/1E76cvuu4OM7+Fue0dVfmgHchAj3uqTMaClKTRK
2t6nIDUUNuK2t5FCZHSjYHbcNx9Aihn22l2NEoDm1JGFqIg+TW7AOae/LN3nIpVa
Gpzxd1InCKTPu6mqLRCjGNY/ETPdXIfUc+GC95jwnOGmu5fAHcO/ceoRdZOX+J8F
rISgjhLaXiosgu0ONAeFfYcEEFHGSYn+n0Y5wlTzg69iw3CzN1hUi1Rz5hAE14Zy
g6K8WKwlUDOVfFu3OJleBio+kHuS95vE1rSvxRUr/ZZN0eCnvoUywdg+PocFe+Jh
o1qyI1yRwSRh7qn684uJSk2TlZWNFWU+xwgoTvQ3OSMhSkWL4ZXwXHDkijnszd+h
h0LW0JWnaU/Q8pqt72LYo6ECqGAywb+z/Aw041JVD4g1yz/rOE5NR0AfxhuI7gtx
OTi9tlnbLEZjWsC9giQyu/VZ3Xwrh/QZQ+9nACiLOzb5EK3h1WQPNxML3mCbzuxm
Kapgv75GeJtVGpidZ79MXpgTOg5Untz+VdhCrnOhg5sBPFZNLEuPDH9Qh+Mqw0k9
L0CcK3vtmeeU1wTIUwCiErfK62LPAXxIJRl3nAMY53WCIDwkmA6Au1F2l7JUHfHF
/u6BPKdkqJVpfCpaSauTpEqJCizu7COsGTptuVh3ifQJLxDZzn9Jc3SPPy1G1gf/
VilWf0/V7GVJfglWFNl7VWRYjXcac2G6k4GWEdm8mewvFTO1IlegpjVqprzk2Sf5
g+wFP2JdN5VxsnUe2SxRPEMBKtNUOMKChaD3JO6bzGbjBugcSF8svEU42QdEw73D
H2eldPuU7iqtEfVjkJ+VYujlE+MYqLYdbjy1tyWR9sPgUkojBr/5AYDmdohhxglz
azV2ujuguhE8n2VRHLcRuZxDzFtIFVp/5WCouKEf2/tnmx4ZNoG0Orbt1LmuoTxp
oYPX0GHEkA7ih3/8qAjSBAsh1P/2Df4RuioqbhO7dD1Et8wzn5lPfhElGUFkZuYO
JLMs6gsK/ICvftsYJ0FSC9pzIYzZJiVcXDFpYYjnIZ5HFx5Oa1CLmiY2IJWZlZf5
g8IXvyplOH59KGFVRxposO/d7N75tAv4sUeBz5/7ygtVHIu/JIxKFGMPemrTeh+V
xN1p7UDaJzX1rtG7Qd9QDw3wNLUcEACCXLNpx4R3rNbE3OYZAkA9ACs9AX8Ga1zL
/LUvF978jbk9bTqjJo/Ng4HZ+H77JxeVjms5WxH9yNnB3adYTd6m21OOkYWlW8sM
fUs34/HQHyB0Is7OeGcsUBMriORgzfK7ZU+MLT1h51xRjph6zSZWo9a7egNsp4ew
h3o/tNQxBx2BDSr4OI8v0GQQKbfDbwBVXJme/JSur+tDda9KrxN2WEh1ENCi85Qb
M1tbx2TXL6aIqmjybPImjI9MZPSdNA56hd3Eu7xpuoA6n3/roM1T1lqbjsfzOJDf
WO2V2w8FitRLFN635MKObnFm4ByzPPH7FkTgNaZyyj7ejr1casJQjgh8WhI/ZB3V
bziHSarUurzHFyuiL/DbkknLFQttl0HYSXwBKqlDdzrB8jPndcGE9yZ52qrQavZq
W8vwWoVxJRRsoMWa96gitm7k9L1CnfNhFshFn1QX953Dw79BaVg4DA1lU3MmQBX2
9xmmNeZW5NB8EA6KIZ6sNxIs82aKhkBNxhQU+KNK235sUqXV9KNdZYWOL70GNCYt
1Sdhooe4wiXfNYWN6l7W3b7OaICffbyJReOkEMdqjbcjS6tsbMVK56gvAc6QS73d
Gc+Qju0cXzSuuqolUS/CuQs5bBRgMu7/xJBtC/Ju4Wy/RYhFdf8/XMSODV4tMuVV
G1n3/7U4cYZgm6XcsxmHZGwBFcXsMvrc0pwkqtpb8dqdo8nYrySwjWinvr1zNVqN
RO4cwcL7mvtR+5ASpM4dxcQwjnwJ/ARt/XAituKICRi12wNHqcAKMoXkflInVn64
D3JII1/mqm3Wjrk+0at2IWEs8yByXJEySZQF1XDTwKWdtAkMc8B2gOoiNkzlvfzk
Tq8P8B36YW6w6ytE/9iUTmwWlp5SezN+PjpYET23B2vXY4jXOLM9GDcmx8UFOOrz
yTKsVudfAxh+qS9+4GWgA7O/9y27VYYuE7xu6DB5Funt+i502R5rjR4myOSRow+T
9oRnq3Ky+zUk+AMN2tfr/HYe1Uj/I6hX1wTYTHTz9ivLjIKF4Usb+8drJ2/ZR43t
/5mjq39xzFZasAJ0ELTHCM2rjmkieR9UE6k8CuiRF2ojQPzmZvw5cytPFPyNki+A
TblG7uGEgTg1JgPZUhLFSB88HA4KibPQY39NVGuvZlST779gCOwLoeUFTW8EMkTH
eJqT7C1wFnlSmiI6p3aBZVmeuja7kgBULwAfU6iC+RwwVZdDyFqNANvDkQc1rh3w
lcSksfPndzEm4DicK4EHC/oASlTEXpMEmdUeafG0Uic7ViksvBejiTiwmTKA6l1E
jJfxu3tdBqS2YbvmkVW5b3zdfhmTb5xB/2NVRMHiVjK1AQ1TbAYM5BRAldfPp4xI
xHd3UCOD/JYBJW2/G18oxZ0QQ6QzZhzmpPkfAkHJ4awcw6BIokOobtvNAbc7WVvj
CY/8aqa7oOGZZaSI+0XefxTjwjoOfM/4cJfBltiJ114HENeTxIQIBhXV38OQcgkY
cJF0K3xYgyffKZfzLvdmzmzVoF2OrkZfxxvd4qo0BkJpFkHgO7MVzXJ6MeEKQ0rl
nQCAvsJJ+vRNmlSr0tgDe7xv/LZuDo0Q3RjGx2+Llu4i8WBuCqEk2FDiS+R7TDWu
nZhhBaHiQDdTVXd34kmXozq2egAw6ri6QHMTGN/tQ5q34AAWceiXHTMWg05LnBTv
Zu1V1edniCrJD/NHv7cIlj5Lvkq7KMIby9FScTDhzuSG4eti/Ir0v4ViGuSH97mB
Cwt0pb3m7wekYBgMqKNNMHLqubkRNZV+J4G0MymiTsQFhWyNUkyP6lXRLdUgpjK2
M0gotSknmZX68G6nzxZ6G6kUuDmSBf+wVxtzWJy7YSGYk9aHnGpB5tiOU4onY3FP
BxQ1ZTj2TdjY1NAHFc4DOVYg5CFIeSHti8Mqb6F/8yTLpqnq3LtXLjbAYEdVxINZ
DwR5uAcri0AElLqprNxmLqOSNtD3KJtdwKFvDBc5eyieFAIeF2C4a/ZSjYueS0XA
IE6u5NRmaYy13yrbFWIDs1XYhlulu9PKaNPM9ddoIERhUEtE2hzDtB5JL8r9VgzY
52z16D7/EvKPNyuhiYLkoVLXz8nCWZrBirpNzZIGT8RWo1bCv/00Wx6dQsvfah2K
HdqdhPU+VZEVqhcknGDtM/diXxXkXFZBlkJWWmmK2u/gftFdlYWm5uEW04xQEUXt
PlBUFp55rhLrHnttuXOihmLLiuydgxHVUzBrK+g33Ws2+9V8lkSEsCN8thFsMFGY
PHvonNyfhOYIPbq8wrCq0PQXjIKnyV1bpdWY//fR3U8QYgBnQUMg5DiPctG91D/J
b3OH/u56NjejOajgiVLNtR2IpeMPOjQ92BOcRM7PX8omJiVZYDQrI8Zfcroux+5X
R5LKOb8jZsWvepzZ5Bk/zvAjvQIHJrJiFVF2dRrj8u2bTz6ZhPkTQn2dvL4mU6sG
ZnWzlzD7o+ji8uqxHzGa5zY2kbkt429L4YLCd8ntB8jJjf5mYhJX+P9TR7DKOSpj
wPDvRo59lwAyc77ibFqT/UEm6uxVs1MCzeo3GTLwdAC9sefhOtpSLAwpCP28dgEK
LttTLFk4jf3whxbW5TnTuCVZ86qi+gc1u8fmTmSG0uXQkLTY6Lp0/ei8mnhOubIN
YSiw1s7cOw3eUxukwIK4Kcbwl/eYAsW3jrxtvhb7Cv2/x+jL2zGj5Gd+6x0STyl8
8VqXuZYDbVMydBtIBlkJp7JM0Z4wSdhrYVVreOOzlSls8s4J4q/C/RweLJwoHEcN
ODFeb506IxfZehXOYFd73/SBZTjhNUatBuN4Z6c0nQKbiTpambFFXpRBR8nOxdh9
WBNOxWWgI2pyyoaduXTUf4yQrZJJnNWU1e/t0oiDeYFi/hIop9/f0pn28//ntOo4
xc5TWi2/f1VllX6ggPXcDygLk+BknzZOgjrQFh3Qf3ywf8Sf2n8Fv9x/ByYLoQwO
ayOFRvTxIvZElf6THvIjLy65oNwMAeG6zEbkknrx3s99/NJpc/WiBnCvQMG/g+/a
CVAoS1iDukD7sRXsDeAWIHrDlO7yvmO4UCkZELMB4dAOepVJ8ckAes6PRYfpbNUA
wLgwRbIPjBCcmViE7qgBM3qHO8HU4cw3amCd+eRuSuXCh/Hpk+mntfJh/zOtGE29
/5oMVHXbIgzNvH9+37u/4haIKd+Mrvl/xDAPCHcENYyvMXFMj7TFXqc1P5OYqlGa
2lzvD/z3Qj8u5c/+C58tnf/xtQ3NS6duqC3XPXH0vPR+ybMbTTHoE6Y/lbpyEMrK
45LF+mZE9PJ6t5z27FNQgFJCKPBnvM5WAKJropiBfIIMIMdS3YvV2K3uPmFMxMRv
UxL0GQtwKrJ1J1SqdM55ZmkJupd08suaKNTxZH1gn0mI0zbnigSRn1/AQj3bAZUx
uYyIXx/Yw/YtPDvSxOMXrx66wYw5QPL8C0M7MTtgjPjw5OqymC+3P2E+b8GVwBA2
SIArVXVoKKSHws3ESfesFrKioswwCPxTQ4GJ8bSl5asDDUoeTj+mZZTbymGXapwh
HSYgU6NXFKwI7MKNakePh8XNJSFSk1sf2pN5PH917hoJfZAPAyvTBKtC4/D6pSBF
pJAYvwCnsddqzNHma35HRM5c7T8ollSTMbOU0rZYJ18qGg1FdVDy7/Ml2hSeuKvW
cOLo6B9KF4roB/m0Mdc8w2WDxQKzLUSCyI5LXVjI9/hWfKn/i0yNgWgFMa1JJr9r
V3v6PXj3Gu0dV/SvYJOaIgKCJ8C5T/lGwTxG/MRXyWARsnFcJLubNHwJWxC2YXnw
UuSXvfT8RoSNMCiwuAHzwzpRBs3OkrTbunF2vPQv1Bzy/DwLS3ccy92IDG3J57dB
SEpuIlh+IwvZVKTUSN0SkcmQnrtro81q+2WrzKQ9gQNl4XfykweVcRi5Rai4xo5K
F841KECEqMoW2WCpk3byXJpf+AZ+ePsZlRYMDKMar5LHtIQjhLJV0ZUr1VXeRoYU
AZYmQ556oMGCNhEDFHHY2NvuDOYHj5hClQkeTK4OsDOxGeYo8x/S86rxp/Nv7gYI
a4H0xtBo5rTglCWzh9prdpYj1BETQzrIEhyz1L01ZxMiT/iMtfeXYlhxJyZUtWuj
azPdvD/VfvxaxDh6siABt6uyMFkm+zenMoAVljEYpaXEjnu14sb56NnTelFJrwNx
iqsLF8RcU6yYDQtcRm9KFcNf2yXRPiig1TlALoW6r/tlZU+rPfxH7mBKlCwB56iR
qGWTSLYcLeY7U249ivsiU9dzlfZNpyGaYC4eqsH1fDX/WaDqA67jVVUHdpgM2A8Y
wN2jdWOARvMxypGsr9OYTqEGFDSF+lQxzLO/vCHZQfWoUJsmCEPWwvWvlSZetpC7
RrNOgbtE1hlh8HEAw+HxfEziBC/uKHvS+68e0EsiBElB17NX+S2NejKisH4eg6mo
RLg02nH2//6ECaBedRkMlzblX2nERWCZMNFSwYWe+KOaZME1sYnpl7c17rezgt0T
viZ5rFV16fOaFXjeGhGNX1vvg39lSCHcsVCylK4wQFNEbL5uWkSC/g7BbHauONkL
dsDAk+MH1jw/vJmZ6OXAiSS0ab+4KyMv1W99aJLk14oFUq2DhvtbbkFKxKePz/xW
lu8PG0wb6CXPguhOfGRhauNuehUTnZEO3oLMWnJ2IZUrKZ6hlCYDy6E51D4TD/fT
L2csHP6UAJAC/M8PoYRZPrp+Rg8PwiXIfKCTb2+qwrJ0nMwl67S+vMhEXOK1ls7U
Hx8xGcqXyI9RUZXE/hEiP/Nri7eX5Ns09esP+rWfpMMs/8lMRSMiAJsX6U+Lov80
96VhxDT3csLLdZ0IS0cg5TwEkNrmOkgybjP/fQ+JEsA516a+Z287zuwSFNbBHw6t
cq3gUYioUPrANxFsWseZ2ErGQDJpbIwn5Xdlm0a/XSgPKI+zQ+0uqo2onaHk5Qef
78eB/qmbFWCEIgPPvMc7QYUMrydDlnBUoJFjCqftYiS4u7d6/+SJtU+WPKw6tN6L
JAfDCT2w+OUpXIG8lA0KhTrmdeBd4eADfnCj6kOle0jHXgrZQDLnW/B+nvXjeugn
opAaIxMlJCui8SXO8K2Dri18V/RZcJ8i99tCXWx5rJy4m7vot2x05TXMm8/kkWnv
E2OoZSkfOokd7jlgQHuwyrZuVlRCPFD9RiQoR7uy95ru3MlPsleoW8pjwyIUx9yx
r+Y+SHq6fSgNhWi8a9BXa1iBQYwkQafTauroPfzX1mXMc4M9Isw7b9yslfKALzkV
URV0gza0Os9SEDrsmSgCLnIM/jzeHENMbzaeTw3NMMiq2Ae9BpeAhC2h0Dt1mnKP
+QDShYvzZttlr5tTf2h6O7Or/1Px8VYK9ULDaW5J1SCc/RthtMKkUA5tg55TDjCU
YzeXTyVMQIfpi0CuRZKRYRod7MPaodlVY6JhZ0aBgdM27drQ6TLMWS403/AKLNWW
LnuboSES+NIEQxrx24BFbcV+dUQJQ+ooViwWljbRFKCpSYT0gIlgJeguEP4lubv0
TQ2zDN56t9RQ4LqrjXQlRFHa8O3vO29U1Bm2ZFfbuQ6szmXfYNjvlY7iKWnFsiHx
LJoA0t1HOLCIQSEPMYfks/2b+JgzbDf7+BPo5SRWxP+j7e1yis/SMWk1FzMDQmPa
zrBaj9tlRqOVe29Wm+7O1D4nD/ZnsxBHgb1pKTzaRN6ItyysSxQXSZDNzfbVnGCX
OzoNU8P7BGxL44o6iMHHox0Xu86e0JdSsp1sIc9XnPbCJUXdD9TV/X+n/HCJavvL
h1oKD0O4C2RHf0fQ5x+jZC4rkIirON+ryKK6CZT/CfnNZ9xPrB+CtPrTP1JKcL+c
L45KlaTy3vQdRKSTGkL+RerNQaJbJK8gGX5MKN+LwkM/fdZkWOnimQ4q2/9gRl2y
xhSEerr+LLDA45ARM7SxbE13edWS+H9d3T8qCZRUwOLt299WFbr3AK46GZXEv9wg
8YqSALH627RJjIEPIv6bwslM648nz6O2ZcOpiOzHFd/8VmksvH7iw7KoB27Ah6n7
Bt3UAxEVT1Th7REbkvZwGiDq6yaoWoar4xMTPVbHLvAv23j97cFQuB38lNLd44q3
db85SRZHUsXpcjZt/NHwO8WoRvn4z7G/O18oF7rwHPfmdWw9nEis9cFozUil9o2M
ppGzVQM51beUKp4+4Lv854KjQg6lnd3+RRgu5N7AA0x1IAZVoSUFWFuWuKc4ILYz
pvW2f4H1tCxsiuoYLXIPkckb4GS4JzaY+ov/UnZSJduJi8U0At6D+ffVo9MT0+tu
GHY3FqfT1huBPoue+LLBESUFDJbQXxQe8iaGjfeks3zBdEIIBxFHauajjQnPRONX
I/1itxRHn8qLmX5e+s+hvrJKeYRfHv3L1PFNkr0TurcF7Lf49RCmqysWvZ85iXCY
83sUa1BhT2kpRH9Aiz2nKoDNIzusi9SlRsmjiGwXyi5RE0jzbmxD5hEzPJE6nH7P
grwx4YuhLkhm4NtpiRQ/ZxKq9UW7tTNlf7xfth9kcRzJfPE2G4zNhyYAVUdJzbNI
DHjGiCCRLEr4VoMrw718wYwgpaUPJuP0+VG3gT86+U3wgMMb77fnblBZQfa0QGZ0
0ycHTWdBrNEK+B5P3aeQbzTCxd/RMxwP4By5/aE/deEDDFG9cTDjh/XXdz2tU3Os
zkEMTgvfetQOk0raLFAd4TSmHqXap0RcY/0Zpe4ltqmryFn864B6IzMrUon8WEmz
Sy+0Vr97skDbsfeikz+l1kRhAxNnotOfaLJIga7KnssRmQJIFh+fUl0mzHKMqePN
itFlQWUcTJAdbu+K3ZnIbDwGdyPn1iENTqqgn9SPscWiGXt1yf0ji0J5TGmMuXAf
+NyWkUGi6ayEvI2OdGw0ueO1M09JfdNAHyGI8HJGNkxpOJhW9s+hse0od8LbmQBA
JXJPDi4JQLAg9xSpdihQ1xN37Q19MRfKlkzrEb9qwXCSYAI5c8xgZ0Usub7InuF1
QMNJI8o5KOKrf4BCqx1QJIJ/uy6yJ6N8iMAkiGVoDr/YuPZUKZy5DS8HDKzUh2eM
GvcLIqLmZ5UCCdiqSQST3De2Mnxqx3PXEjj5lGVjlPmKWDA8WBR36Gk2ZSe0Afsb
Z5gUo5/dujVv+RAfYSsjZEhxsVxBhER9YP+eKXZ+oO9xfEDAcKz1LkFzvh5sKtEn
OG91LOE7bEHkwwD6Dit+Z4xawjZ2b8cnoTzE1Wyhl7k6HHRhcEZOo5pt2YZMQkCz
qZMY53s0LUFcs54gQGenRn2g6CIwQfxCq28yjmuvuYh3jVeJcG6ZiQ5+p2L9je7i
QM8KN8T23BMkzAd0LTa2i+3EJaUS/wcgOb6MbLXn5HbmZEt/JUsy+BhRYZL2+YnY
ZsNjZaIJS/+TECVxdwxOB5e+waHBMyevlxLrEEiQN0qe00E0sQ6cPL5GZRNlAy7K
WYZmZ/8VzuNOcQ/TDozCLDIapCFW2RyOP3gs5nAYLUTLvkXYSITpFuTUFMbAsFKu
lb+eq1ns20ejBuM8VytWebjm7z6QmErHhQlPpC79hYlQfEkDUUjbwnWxtJtJ6whj
Uk4kJuGWinSkLXROXxWheZtdcT8c0mMQSor4EndWpUcgQr+dTdB44l/6BHTJD77Y
sgzqtcwHenq9zcacBF2rI14gcFlrhe3zwd+bqxMN7STr6thOsuKA3i4itnYR7IhP
9b+WvzSMoSgR255zNcI1caVWMVT36d2Bae5oD7aOwj/Me5TC6dZAEhcH+KdH0O4z
MiguMQKdKtmcMI9DFFDu9n6veRs211hL5f9g/CY8jEBj5dHt4rjw/5RGvHauhuFV
4ICEkU6VvZ8sGIgvE+tehtNciJZgJmXWWfL0cl00Wj/D79zW6QqCSye8w9QlWXYZ
mrHoSlrHW1565Hyq7NfPzjcnmwS0Tn1WcMkS7xbXLpkLtk39Jt12KWW6hW1MXXph
pIwu1VXD3/EdB76w2vYfk4nIosj42BVUh27ZVk9Oy/I9a2vW8XpRG880Io/QZmDi
IByN+W5WatvawXeWqQ9Dm9zEdRz1p//yWlKJwxOXE//7NCjybdcMsVSxWfNdCFaX
KyJfhmahzvjKC0LIYOoXAH/lpmEWd+W82hQL7XuJ7tS+cByCCEVnMdPl9PSMOsSX
cdnLKosUtcSURu2rebF5LSJENAY0mqIlaeClVX/s7wKiQ5k36T67cPYUmzRcWZXX
J1hIHgT+yX1cmQyHag1fHTa3Uco0R0bNl60p/cFCSLcf1G0Y2D0CKihg7E0hM3D6
dQr7MtIPs+6pRlvVNbUv804XzUKErbFPTo78CfQnO80k//ZklJgRPa2XqZ5z0hD9
ilUFkpMQKLadn8vxBxcdaDKTi9v9wkAcWp9yI5MsUsxbIog0i4I90jrHResFrW6i
l5dq7qonACjOF4xBA9Nlg8hxuRicIIJPiCXklw91Avvn+YVV4VKWxtU5xZqKiixh
rJa4rjrNeVG10UUWHG0x9x+1z2eHItQEd/W0PfBho1NMhzcFwsmE2vs/OQfzV8Ur
Q0ZPnj1mm17VV+Am4YDC5W6UfASggIF5IEuFFw23bNgLFJduk84NqtElEPhBkyJ7
OAWaYj8KLGINMtjqZnqGx59WCoSap9KZodAUF1dy+v+ow0eG8/d+OusEmS8uzK6C
GwN4abbEMS5uDyUs1YPJ72zvpM8sF3EroAcMmu406Nya+EU0LTrYXSQTh8ga0+cd
mfScBHKBHlOyINgvOv8Z5LjqgK4QRSfafuEclrBqBWwAEvjgvCBvwiywEVcUheRk
t7E4pO/hcvXWQBYULLwqb67Z2kj6jvhLPmli1yifH6achc3TUKNGoztVNe56oDQJ
ccRTtfdUp8GX4fUrzflxcy276AhKwF6uBG/ljWSeRnIKX0HtuJsqo9XywzqMtIec
1OexKsyaiG6HBvIgiIP5zW3/N16vy8hx5tL6d8KJ7GISNLeBh3C8pYam3dMzW8/m
wn+iqEIbsNkC5J8JeBlTFyaZ/iMGmg8vfBDL5y2bVD4VRPkxBjoO1C53dBX+hXgM
YVW+HWW2fPGv7JJybZM71tZTrD3wvHmWpzL4P1pwptfhKtV27YSpdJrWqlqkVxDb
E2kPmJ7EokNQxVqSHor6Ky0CnezrQoYLwUsjQVnIbt/EHDZ8B1nnBKqERJINfXPd
sm2DvlzvHCgFK9yheJiRaUcl2NQYbJs3Tz094guHB55TcvfhgAwOpoYg5yXKRpea
lXJLER7BRtzaMOq9zrvo7XukWv4Qd82I/jb+AgnSQtOinGSu2NjY/q8cc2uBRJ+H
OW4XRc03ZPnaH6XJglJnoGd8UZcdGDfFKq6A9/s+748E4y5gqXul+KbV/aEXc6Hw
LTlE7FNzyZ9T16L0qKIU2p0rF/FwzEObKRuTcUkpHi3nExd5Qd25vSbCUlrX7Lyu
qCVDxKEXmuPtFyAtS95ROHTDFQDwzy51r92izrhMLSe02seqpz+BqZ3nofRv1ZbR
9R08cNkU0Vm/fSQudXMfAI4kKWbXLYGgF+/ZTj867Uc4si5KCOZvwuTXoTq/7qjd
xWRjOXYiX/3pxetKVMgVR42QDRExb6XrdXsINONWB8nIoU+szOIsqp+Tu2vyxCNS
tS3lnFhur7OH6wCA9AonY+QjDVXkqFhI3ABK8jwj0q0cVwyK0aSPKKvAgEQp/Qky
FOs/uTOsJo5nosNtaQkyxpFjLgAehi5ULqLHqpwYwORafu6Jxns/Hrlunz0zXL2V
GnuVoy9kknsGpoKH6EoSFnOXm15Tkr64suxd6IekTaVD6YNQNq5I5e9a5M5jVvGR
parZtEeQILv0L74tyqmarL/mk5IyBoke8wUVGTKh/zGo6ry4vHTJ+QlqsBzxQCIz
0dqXtGAXm7UiVvFWSTJj1ucF9LBflnhA2iCBPPjEVikf8NHaTX8ME+jkP07zMrTc
RubhZXxwGETK/cbML4ajYr4Rkv+U5RXz36ZnRPXm9fROip8h8zXU3oSsLt0BfnIA
zf+Vcp2hohupSdcjp76DWOQMErNzERBBsZibbyrUS+T7Ls5xTemHWRFqDGCZH+Xp
CvczLIQbvY+/YO909GmWAKHVDOezRKHLlgyVIDeojNLX14NvK07GICJ6nu0OENFH
yNnuwFj9BSaqt+PiJccjjBj5MjR+tpoC7NY+lZfzZqAs6P6XHJMH0ZhHIywyYV/p
Nzq4pT4BGFpoBRis4ea4t25qSauCa0GINrctMBZmUqulCWEEQHQKA4duzBszhgBM
+APamQqJmcMgBVldPBYKNcQJhWA30uMUBMyonUI3pSaP9E2fgLOSoetIR1merMQz
qq8mbtVvU4NsGHzOmBd6K0x6xmmJx436LLw8Sfy+0iJMJWr5SQKx1kHK9XvHumYS
s/HlOpYglQZTq/4EpbL+mkhUJK2yU/0QkeAPQWvGeo6x9hQjYiiJBz8SlFfofb/5
TKYpuTDtMESTqgzZrHgLS/9OAO42AYX3nj/vYhISYuBy5kEVlJfVAhiC2Qiirnhu
1i3E3HjaZ1jj+yEJHobb09x9PaQjQQmsC3snx4EGHRLUmIZ5MXX9pG38Jw3FE1ju
EI6H5XXWByP/UPNM23JH8/2x9xVzRoaUNPK89TrFpDY/gRmf1SFmuH8xm+yqtOAC
gqq8qQ0hzGlc57vD7NPHGtpk8QxwY5a2ZrQJYsFUgrLwENOabdGIJv5/+ZOxuEip
PRm/ATRTCJA2BnuLa/aGMGhGf4TgeOzhvroxTdI9pRp9f9ryMeusY2hTeyr6U9OM
qFnl9WPVFipzdqGYXA0Xlz7LP0KD7dKdTcyCtjofufTszsISAdovyJZx5mjlelSn
+Bv0vjhQFj/AgYU6PhUwtPXXxUWhYSWvX1+C4WhGBWlWb5z2yp0orqn83MgFDksM
CeMSacEYOup6JMUk2xGsyx8MJTD7mKJylrRTGv6HWml8eh64o6YG1vhyXPN+CIuW
xmCqhU5YPN13iFWYZDvScFf7E3M4ef8P+bhnI7fvUEG4gJ2MXoEvOzMSCJXhnLTx
XHjTSpWcBC61nFXQne6b8coTzl+/SwLZ5OcZANF9MLGoTruxrQLIJjb3im3jl6Uy
zQlnAXty0zRTT3CuhObDW0HDoUSM1RcxxEDLgmmb4wZoKzcPItvewmWS+k45tf/m
Ruk9UYiOvq60LjPbVNPXTkV6zgEqTtjvadB6pNxIATqEeP4VoGTWSwNw3CgheU5i
jDI38Mhf4R7A+zwSiit0simg4TiK/9K515pnGYs72hdVE9T/2TqTSGK0KibXVY3z
4FEWlXDuUynR27ol3JNRmgtgQ7HSWL2iN9WuCBdInYakLLsJziYqkSUwjVMueMgI
MCZdJktSeguN61QttZph/2QxWDz/P7s16+oCLn65pVfMr5Di+CcmykIU07xsY+qu
3gOB5uu7NjdhF8/w55h+XQ+1ehJ5QXYML8tjY2nSlBuPxQKPYNCCWhYSZVpwdF37
zkheKReT9pVsjgCDBanQHI/Xxw7zGZFYNN8ZizVowyACQKxLwrtAv3bOkn/rDmy2
4YBuFYML4vuGgKvTSz4yhgCInTIJMIHa0QJFIJJv1RfUaBDBDFcwI1zykqSRG8Vi
ehE/bwNf9AA70YYXHV1T5iVo+F07vliKoP8pcDC/p6rRbi3NgCLw7+ZNNz18viJy
aPFkGy0lNPPpW853FugK54Tmtm6mVcQwrUsG42lH/LoHnyMfiL4OthOEJMQqw6Ls
Cuf+Pq8BFhIgffRq7gZdzbU9Ueu2dbm21pAVvy94JCoAqR+RMrhyvOGyfHxhCpFn
D+7xv58AoH9spQ/hX49UCtrqtMZvTv5eubr1Ppk0YHjpxQiloS0hSISuVqQLSSn7
Q9xMtbl3hbVsuHQOkJomkcckJpZvEYHiZa7TycJODAWVOdcdfqixqQQWyPK+Nemu
dYbnjBrGojoPwfmYZRUNbbSD+onhbXVDi2h65Dek0Kc6EjxBYnzclIqiuyO1mKgK
1OebLJ59R9VWvq469PzbW7LRsJiU4IFea1BwyIvT6sFqG2kKxLwlZdJEjp+6C43y
iSyA8Htqk3xPmd3H7qobFJwLi53rAweykFLEN7IzNwCcDqadiIDhCrCB6Apm5w1O
RYAbNugspb0ywJ+4lorAZBnVmOcPnfsfCiYzoUV7i1zwBUN+Uh8AvCTLEpKT1sRD
k9qBH9Rc+SIZCJ5StZvjl7EzQyUf5mVc8qETNur/fmjgsu9QoGW5DkJv1bqBwKu8
iaW3IOsC8R0/8DPdQpmWjCGbm0yLcdMYcav1/hARAOiazCXeCYYrUNtuiJUGHPcH
BhyLXPpG1KDQYAeilVrAjbv4k8U4mBsLxdufUBQCxvq8yOfgvWm14Pu5pScpVUH7
SZBHfHNM2l4eq2S9LUH6am29tQDFTm5xfT0bVUy8wsei9AXXRZ8PhjNucAIWTHcQ
sIx6Dhx7fblbsl1DDGhHRHQOX8WfDz+nOYTwgOEtPclHsjDDwUCX08ibTn8i36Kz
KU9CcPL8xBRY1Wc4OwWom/gkop/xzICZVv4qdshGrz76dshuJEG0khrt+3+gEyFG
H67UP8MgXCUjV+o3+dOCaDi+rQZS+sU1AmNiKN8AWGnz1SU/NTGznvDSNQMpr8mA
2+OgNA3vmasndGeGUweoACEZdavpKY9JwIKWJ5WJMqMz6gCze6v+01TyJXl7DEa8
M8D5e2cpRByMUHV+9RIOX+hl6o4Rn1/pe6kyhDNaEQKvrB5dRSeKH2ahpS42pOGC
OeGJtyJ8JggsavzXy0xJJ93p9em+OPOr7Kn6V+xZENAyBOYnpp0PQIEf/ECVBG7a
/z6f8G6zCPooL9hUGOd9sOIKjjg9HbnD9WLD7tNhLtJp6w8CIN9YNiojzUyIbp+V
xL1PZwVb8dGeBy6y1yFL5XN0LeE8290LZxcuAh2W5wKDMsRxUBZKAnVYjmoRhenb
9D2ZzQX7Pxo0k/9PI8e2cKLeAYE+rdaPcBuXcpLKXLR5CTWetWgNUIrkzBgE1lPc
muYrX+QFQLw/HUmTEv/VgfWSYk3YCCwNosJ5g3lb/RsdUd87VVMT5XX8oktURKbW
liW4IAmJfac+wPWNvnNCP0qnGcRaxEl71fGIUZ8nW4aNg/T26SGLbWMnr6qwFWAU
VIG6NI1YDTJb3EHUsRJwPcWXYxSNr0MxBg8ScUUfntQhaNi2yytlntya0ppVJ5qE
UyAEybAXpGtHMV/5o1et0d8/dDSyXwCKPWFCbCkEYDuaTLHl/O9NwlnpdR7KlsjO
NZDzv7ZoijxSJMCkGub/IoXnvsqb7bQJuweE67V/n04ZgO7dm2Tv81Lod8/qFXF2
1ciiHfFFNkZ9P0/k6GGBvfgEpYTHBuVVl2mmZHF+19Hr8TZHLtY0uL4Y9JRKcyu1
nru+ILUjzgxbFRoQj5gmmD0cpGsfFvNBK05YMGrLYa/cpQsNgw6INMlJLy6E5kKm
DLdMlx6yHFF210L9/B31mIWbYYc4tO2NOvcpintmajFpVp6YMQv/iIu71O2gW5oy
ouijy/aLTwEkdt0HUqEHYk2UjbMZFmiJSaJjRDsCaGVwJH61VscUdUO1P5bvE17A
JJf4q7c5H2HSilWZrN5SX3ATFLV/QCEy5GoAUamC0QkwaVwLyLwaDk/voM1nIm8T
vbqsHxqmluNlCSTGRPSjKhjKnUqhRCnfPwiHUtljP5m2G0I6IKHh4Jlh6PEk+8hZ
SPcK+xZ+NxsPJdLQr+tUYEMrwWbIeLrE/tLC09MTtnQzakTWRUAHHdZseC5W9fx3
i7sPUc+oXpxktm6us2j6uD8E91kvbMRU21KOMl81meFhRopE0LqjQSe+VAeZlxl7
/TFjw44PA3wdY4JtWYbXxtJmQk06Hu8Cq4q6MbzeSMrLczM7H6vFGbCVcvbUSY/W
7VCErz1CE4JkEy+NSu21yqRJ5jR2pOkaFYkZNSSu1b/rolDFjuiJE+sBaz9SHcCn
c4AqQt+rtYsv/d9hOmyA6yF4fJCn5mc57vqkXYEg37A+Bop2KtMn7WRjvLvYX8a7
lVHZ5u0vIgaFKefZOpr19/3fAZzRpF6Xo1D5ITqnX7re4TB4jdrjGNCbg3WHcq3J
3YCa/ZyypbPmg+yBj3tZJa2QDaw4PirfIjeSWPjwlNwx04RVWOAOfJmSzuNQVq/X
VAmC+87Kc3+UsscDwoqCVafgWaTtF4YSlOZPt5G9AZ6LBSXb+xSoKLcMcanrhmd0
8WdlYq1KNYf6vM4NX6nph0yoULMS0hNtjbh8Mr5fXw7A72AcgDEmTxJP3fXI/MRy
g0Yxv3Hm2im0UYJwTfUxY9Ddg2ZCI6UzBBDhFNia3+LHxJPl3LcRio5YqNUDuzTo
uzdhOkw1I6jmz36RPJ8+6azlZ/UihQO9ZGxXK9YrbQAVILy1tfb/ZopKyRtXm2Io
kb2PXGykbiVBRtRkRBft3E1ySpeytyPy7bVNHSrc8BnPP5lIXI83727Rp97ybsV6
DCc9j2dAjjK94CNmdBsGvgLHuDDYaloPlR0Dr6rPWPxANqins8ne6Yfn14vR06d5
ATw96Wa1ykkqXUBReIog04ciJqxeymXN+PZu9So/vqZ/0P7niX/8AUtu7nY+mMnN
goRzwWz5gVr6hwu52Uy2Dz0AGZK80TIUciS/m6ZViVVg02QP+ERk0k0ZdJ4LndI+
eT/WB5f4BFhdIqjskTYUTVy6Exm5Axx+BBhBqxTH/j2UW3PuJmUiwdsQ9R7nKZUm
717amw3RivVAi5ELeokfu4KaDTf+QsIEvelosI7Hu+VR/K+2OfQCelvkYYJxORh/
KmBDas+SvTSynMvoE2mZbqcK+Rqshyr9RbXOQj4WKe4Kz+j2jOM5ianSYn10P8v4
SJ+Pk8AN+9NhAnnqZB+5TNZ0h/YcBeG2RvKkzUiCUtbPujdlvcfRhjBnNyWNpBLw
AoN8xaezD3e5QtC4icPwrQjtN9GwjoGhV3bToLo3V4LytYA40Q7ETF4w8EhWOXEM
GWD4nChJv9upiQcRuTbGbiFDi8V25B3PypDiPpRfsaX6ATvCzqjpEbzRhokqMWS+
qjFCr0Qjce00AZLCaB+t2F/oqCJTpBwsfJbk9wAsJY10fJZUeFe1Q3mBpMSUPMND
xvaA6mWXej7XkHKh9QRFo/J7/1BI4KhnfWlfDaU4Ro4obRQ5y4R3/bvSmtn0tz+H
qXBVkOToobtv+jY31S95oy4Gi1rlLTqYBZaVfPMn6LqVf/J0ReAH8NYpy2my6jrh
8JKTPue+/6mLOWegLJTVmvegMF+xH/xPQ11brDYbDfMb+PjRiBKEiVJuvuhrwZZW
LhhS0VPuCUePm3sl5hAIwvRnrM2B/yAAIKzCdjqE20KNf92T/JXwxhzcNFs3jSSk
7PZkLXt+X5+RhVt/dbFMJcUv9G513KGrjMdiSKLHygrI5zYWfA63Y8K+jLcaGYmL
zo58lXNjRh3vYoTbSwUxo0Kxdfvn5Tr0aGiUkmcIir/eqCGQwlxfGtHRKdwPLYTS
rDoQphbH46OIbaTi7G1npunbDfaf5wgXhDp8kF/5bnplQDvbNAjwouRnbUNXiHCE
+l6ENGdczgbsXtrfcAPHx2OVtIWD6uzuLi1FWiN2N3wxgpg8XxQpQVp8dL7VLw3B
t+TrVjwG1RIl3IUVp9U3ZBERtIjV+D1mWTPFYULzW95bIXcK6U9FuFGB6IUUVUUK
YbaSpp1SquJ8ZUMLKX/c7c/zoItGkQqrm4y3bXccYd2Q7kDKGqltboBTSOCajCqH
rnUMsDDrmVJ9NNuQfI7xmJZ9wgiWxYn0icSXjyR3/inmjk4/tY2EExFuxDzhW9of
aD4fM7vJMAfXIw7hIv0sgB/KpGGHe5XePuZFOdcT24igpUw1D1YOdbz5NBuVM45e
PKDPwMEJ2vVyuUDONikiiOsOsfC6anjCat41zijFXFBqbDdAPSJ5N8hB4VToEHaP
DgLwNmd86GbO8M1zHjBCioAX+6DYtRTzQ2qyHTzJVQgez+w4EmUj0raP23NN+WjT
tk+RFGQnkubzpS2qvbJvxtGJPUrDX2wRkgroK4nLFHdEQNp8Ir4NNinkRWSK9FMW
QRoxmVkt4kYN7cEnLoXRLKeJkieu35FkGKY6zD28glVpHP4JSNdl70XCSNDpCR2t
k7gUliyZBCS/S10kLWcP2t9z2zN28ULdemwvBYitS6r/nRD/nNSzUZEWHBBr3bWH
tG65X+BHLyiN/RGhSc2owjQ8uwPVMWjppN85OJIdLNEiplLDU3h3g7K545ibCIZc
zDNc+NlwA5BBiGdc6xerhe3aAJvvP9OzmR5DEn6R6hfU5O0pN8JC2pZvY1N+uDmp
fvjAZUKt4/+qt2CaQLnFD49XWVjG0xLbFF6Gbahn/jJH3jIcOzsflDZySr+6wSwF
XzCZGyGSXShNPri11+QljW/I35jdJTMv1QpXlOpRJOdz8+FtwJjxriH2ZqhpZhh1
WksBvnGj7ply6tam551pIc1gCWv11J3iQqdwI2YSI4wMsXIgGe9mahe4H7+mdciH
1Mu6tQ5BZzAKoAwqkcCq31v7nCehR8sF980V9rpFsaC+4l/Vul4k5TO8NZX7lItR
NY0/Gb+h23+IGwjyQzKkfkrwYcjDZtxDfH9SrRFIGv/7gDkqNGWFW0sAzQkqrzE2
c4USTwHXR648QqPO/el8UbYTdGX1LNkwlM5GbZSRk8MrHuIcA00G2AFs0yt/uLM1
IE1Ma87XUCqdtPe+52L8cW0TdgaUiwN7t4ck3GvY/wxw8JDcOPS4qifYKSqIXsPr
uPkhnyOmZSpJJgM6yrmivALmzgH6CQJQa4/+G3q/Wq8Sx+JRqg1gO4iINmZbinPA
UnPo05MgKPWDslPyOj3l/lNxV9REn+H6zE1tnV05ARVxK3y2tSCm+iMGTJpV2meo
HV6RD4JGZfq8zd4GpU//CNE1sNISnmJ7h9rAF/hU0k80MNPjFmwDHZzv6CEnysJR
0F51ooD40lbfulB5eWFil4nZj1kzTkpGZEB1HvnlFFv+g25K+YDkoOR7s5+Z36uT
KxVoqZb/02zP0O2BkxrfGDDyxLWja/9TXaKi3HyMY0jnQj1Bo+UZUr1ecjsc6OK1
eT3n47OO2QYe7GVH/kQDVBnICvtpZwPJqNCx97fhoTdUI2ESbemu5wSyUiBaaNS3
ih+nj9gyE3ms6oDYpQyuukqwO+caKQg+dl7wXwQopIdNoZEQAwRIW0SqX+SmIJYW
CfexJ4F/iPP72oYR5xNv1cWANCXOtG4jhj43z5N2W0085A6GkaxQqOIFxdvXHSCz
HPC+QazwfeqTPG1N5Ed2QX6Ut79i1BT1w3UzCcYrJ/PWZ70UfclIsZ88+fXLCwSA
vbMUUWmwegTZJtO8d53NpcvWUA4M2Oy9gKZH9VSgTiT7Pqk74cXjAgVeVB+FG5Oh
8ICvjIdI/Do50svyNNjfv7PK5HYLehnedzK5kKnERSeJL/Ue77dXnOHanvbdLSRC
2ebD3N8JpYhcVg7uZK9AJHe+AOXeuyOrz1GOrnzi5GBCR6lBvVcCPgOHPl+D95OW
eBi8bipk7rBbQS3X4bjjMirVbmdLSInuGFqxMAjdtJXKBDX3IRYLVdOe5RYqYz7w
ISIlC5kMzAsCs0q2gMpNMUgvQmG2ioLltzSlHyLV+oPWiwSRlfXJzn8/v4QySL+K
JQjAWSe5Q1BrvR8O9/84HZUjfV9+fJFbCxwKRmR35l0T4PB/bH41t++2zqiqGxVB
siwRQCx+cWFg/HV7F1O17+BmM+fiENGKnMCyzwjsk1jLzRBdfKdOSsLU90jkSw17
l0dbljpUPBC8fhgDfO2BnRhRNvdqqnsRgVxL9oUcx+mo+rPqRsvwpKeL4hfq8IWV
tVeMxp3chOYGNZ/fznRUoddFJKBXfhm5L6/1GSWR+gy+wRXPg1Eag/Xf/jw+r3qq
AtLXAsKrJubdY8EnmPQDdKvSOGdIMFHTh7kk267E61F03TNeBaoOvVFxkir+5SQP
Uru4qDOwCcYGPIGR7JupW2yphnsDxlb+Ar8hVeEZzNA7QdwwE06RN7uFvdqzlJR0
ompqFVKP92zpP4nkFBNfPAi57LfW3kFy5CRz/AV/SaJppmc44Tz6Lihu+i38l6wU
KREk3zpMJnBPkQJ6bYPn4H1yizuS5lJIEtogQRMIQSuz5KWQE8EfkCMvLyyZyLeq
gL+nW4SvObLMM6paxmiZjx6TDfQk5S53R23hhRy+iIjYhri/FhfVSVAJjw6zK6ia
+X1qOnVFegfoLMix+Tnm0kxPc94gAC3GxFLe6Oyq3IyfXMl3aYWNDxYY/yNZG4JD
judmwKW+FXxD+OZ/dPLs6F8lYFZiAvhtAEfPuoZNMvCyHmmvE0rboWCpF+6EjdnF
6nAdJ2qdoYlBgjfDULSOVq80m1awzdoFEG+vTDoUArfZInripEholo7s0kT/E8hO
U350cVhDhJZjtaqOOYxPV0AiLDmdHvY3j7dZtf1ugtx3ZbYrM8w5vx1nyJvsxHqO
pzpnyklfoIG3JwGKn24k+M3P00huFfT80lx/HUkyLY9MNY1VYu5G4yy+b5DCVNHj
NIjH095f0r6pkae0gdGegKP8hfAhdsitMMIyNQ15GyJpyyoZwnBxyzx1Y9PWyltp
DJKy1LEIcmPA/YVifjPPPJ6v/xR/+CxYAgSi8/SVyWJK3fy+Bzy+J7I4VhlBIwFv
4+tbLC7/cpws+qAjdEUdUtr++syROcwoebH2rXi/NPCL25Zw2Hw3tsDdOdeXLGqh
/W4+Z7bEdMEITBJ7dsC2qpNqOFK7wlWMbBBylMEtxwmf2Uo76BuA2KriaM9vmPRz
OGQ0+K2MLDZBZ7/NUGjfN7mCaMqoli0ytGtmtmycdkhcWmcTxnn+WmJKWXLJQgEV
8pOcJaT497jNOujL+Jblq14AsSovgZyGBM4d4U1vMZn47Ycq+f2lNeDaenjpeX1v
ht5oSMjkBrIa9tnPMwIq7k7LNiOWnyfLdXPJ1TYutumh+tyJTUarweLqEDJ1orAM
G/DR5AAdSaMZci0jf6lrQtvcuE5EOnzzl6fBwZR9O2CjgXrQqhuH2iX6w5eVrD4X
dkWrhSS8pPlklpWwLbEGhw+3t3aUWxl2t3Yar77XB/EgZJ+BUXjZnMXH4p/WGmFU
S0DeslyUtNMwwxr8eJepm4JURc/6ffGmYOlAfoRHSpSmNSGYpl9ER0wj5pq1TMht
YhZkudqCnAE4lTsbdx3Rb5AshfCWsjTaiNhzCyJ3gD2p8aViI4+/I7NZzZX5JEl+
3rTH1gdUANo1X8Mo9p6LK/Dh10YWm3XzHeM8m0/+HiroUzleN8MepSi8CBgPMtNA
lFo7EXeAjtiurXoTx3mzomkz/bu8VHicgcYmQ9CfqMCk/uHQIyd88uc1uCBxjC9+
11MvvvwoDXEBTmLEZrz+PSKqXH3BopXA+ZUJMtwi1BdLS58V9BsBlVQRNQiqwzYz
bLpBj1YRkbAOcB29sYGUmi76DRWmBGKOSgIev+dufehr/MJpWaWRUqo4PgzdhLgq
2lF18m1l1PhXOvqCT3j87dL8Zag3z4Re9jxrHXMG5Px1G+xINb96V7vIZGQNaMP5
mcsBKfXDPoTlequgHOIy/qEKgarwZnhPu3kM2LYh96TIoUwjL6zD/uX/9p5qvIVT
hpOMVknzRrVTjFLa2SvxFbzA74FiWqUSAgtITgMw8VvLl4zydBxnjeM9XKDNFDYh
91//U5w4GRFhB5O7HCPrRZqYUnHRphI8PUj9Vvg9JkB3V+sr8XJTucStTdO/HMFG
rDFulnCRvfJjKWyX859864zcO39rjH/7HxLF3uotNIDuPceEjdHS457Vyi0CJGHk
p7DFsG1Q2WIRoyiCTrlxtLajO6TaYgctETl9blcUp2Cwo3btNfxAP4umKnRnwiL1
PKgCYWMhVnqc9IaeFCsxVvMhd1Gt7nAuo5LgNa4CK1VuUhXm2ictrH9DK9zQX7V1
+zthL/1/iNZUY3D+0FIuEL/hl5Abku2YtnwADvD7qTqb2DB9iUJz4Xtg5ologX/t
h62S0yCfQXWFC2R4fBc2cRrLIZtscRoNg3ZErTCE5fJwUfDYuq8IVOHPOsBAhraF
KcUPjJN/DAYCCDPrVXPqNeFA6M0hRhK+CaVoBHOC6HRy9g8qVaxj/OVMGgkOO6XG
0cVUwMozKEtM3gILgcBt9tkKTSJV07kWdNyk9Sm3/g6Lp10cx8QY+HhUZyvFV+/a
Pron9WMW/dMskT/zESkJo37LH0ul7mW4B0RsuN/jU3g8H4f4275Jb5AiEETSWFlj
xs1rJ7cb07trU2gfOYRnBzpfhdv7qsJLlYaFkrnLPKV3Lr0Bjurn/KWIWcAP3ZCo
cBH7Klbis3mlg2vegj6YVj5g8XYgtGDT30nO3Q3ScmsNK30x4F8EOk/4PKbjLclI
yxMyNOlg+zfsjoQiIqafUhRDvONNId3FRH4qGx+iW4hKa28X/6c5JQkGct4p26I9
NjsvlM7ZyS05JhTLvKMW+IcYZowZJaV3ki0LTG/9D4y0Mf5BR8iwhkrOduGqh11o
4Ro8WptDdaD/jK8F09ehjT5PZ7ahQT46PMX+bJVy9bbENUL0Equl43e4jfgWgAGd
JwGAK3tmdIw+UTjsL5EYeEYwqyNCTJ8zgd0xj+UA96xsrtI1fLh8JlBmAadep5Ri
ls2OcPZEMIOC9pbtN09ZVcys0mhqrVXLe2AJgbMNjIROPA+gpQAkUQRdSaV1qZ3a
AiaF9bqSRcF9ZMPOGiCL+FGivY6PSkNb/znyAVTLvjg1IczLk3VPOVkc9oxsnbJk
mUxb72CUioz2IIUb3SqViqP6qFSQA1J8OaUXw81oDBvre2kbY+sWQDIEJiYvEpsb
6a9B6x0jI/AyvbgzFSYsHk+uKKav4Dw1/8/Th4Xje8R4fRxUVjiFHqFGRG9lSgFt
owor9JYq8zvuWZNNha4nA6wDpGPGKKdohbDS2c0ObqQ8DCP/b2VQ2GFB6tIKsutI
L5cqZoK3eFCo/w9kK9yIgjr4lnD71cuGJutrooDoskNMEJDQhFzAa30psg8jO0sW
r+YqcLud4a7+ItBdt1XyhUXc7IvGaIgrMV+i3f7AZQFkSGeQUXCLw2DY6dbQpcys
sjr7JSK10cOhs22ly3fEaMi5wd2Sg16It6dcWOh/LlbCAqGyY0X6QdVgHG2G3XyF
8PQu6XmJB0mTYKGX74t5NgOb+pVlqzjsNtMTauwcYG8ts2onbBKnZ4RMMJsTa1Ys
O3zWWhPYgX71LnxknBQosKV/DPD5MVvGY0Vceb4UsloEiI5p7hGK45bJtCNPtiwR
j8XrrtIVWDAK6CCTmdutFxa+G324hWDzh0kmEj87zrm93JvPh7I15rDdAFr3qgcp
lxbzAc98oXwsw/jN+ZNUa40C+rfEoexFVZJUMGxQnWGhuiv8zeypG1Hhz7NpzaNa
QOQPqHtL+HbgaMGfV9Ka6FSJlfyB6zLVp7q7VOgTutmL+ZkW/PYLfVJoCeFo/Ldq
OV+P0FpybGQJv8ayQD7zmKEKV8lMyipTH5SON10dJB17+iRiQdQ26UaSFcxjbEOy
dAwXOALp6r2VyQTqXhmZf+60YSKYwdEaJBY89HGfIkQcXtj/OKuvEMvfmmQZ9vWy
MaXmjoqhtsoB0vYf0xvozZGviWOoFBKQK1jsz+eqHjyo4491/wCGc7T85PHFontm
a26pKWDdMOyFeeaTGOx7Uf4NXpMAMPTkif9AfUW2w3qDxfjvaejiUZu+ejwiv+UC
kp5KpTKohCPQ3VVd2qm04CoSCH74+wFw83QB9IzN6QDkVh41j6myt2naxu+VwZ/g
P8iGTCxxQMuOCZzMq57usFpXdpzR9rmn3RD0yCTiXi6M/PJsJz8X339snp5ufCRw
ZR+62JoOYmfsYG4TXMtKpwQeE7y/Nl1bPgXajtS38EYTYP509bO41Wp1GM+iJlcj
URYEoZxE9qV+zwLbU52n40wVPnNJD8K2MWelNlb7sGuRCAfH13laxL19Wqxc97uf
SwBtNEMhlV4cPXe/mR0Nsn0prSPU7yPF4WwRfJZjXn1t9TXEM+j29RLoM0k4Bn14
x8nEtmf1y6UDeAU2XBOYPP2jnVE0utxsaxL49kXmtMYN8fl4AYx/wkPD/seFlSA1
pJZC1jSxcGqFB0glqKMRP+WEqKPiwB12oObdTYHYlobjpMBEt5gAQml9rUJCybM+
tfoFrhBdNnvVffkOlnODF/mj2ez5Mz5GDwYhD+8lMtvLOb0iNid1qgGLUevdam7P
o+acHuZ0+avk7R8hyJs5IEtiGdkTsvcU+5XakQ2dW9fZTo0hiGnbi0uSPM7rR4z2
eHtg7yQsN2xMfl9d3GuXVE/3DNoQvWnZQeOriKkHOEH+qI9gx8s3BA4FwKbIHGQi
2ByxVk1XoNn5pkratXLYRCw8bbaLZViH+j5s3BxPWoPnvasD7vka+nX9PN/5dn7x
M0/z9S/jvVea0dEuGMlglbWggjZ2pRrViZ766NQPoLIyqe+298aLN1KI0UQr5dHz
tx3cfwZ189BNFzrVCrtYIaCbEfKd3arz504DnQqnnjmNVilYxz9aLAYTepwPsMy4
IfICn+ZkogOFMqItPaY/Fd3xe6yBDz+AegwO4zexKIuAIyrBOQtv4Cvvdr7m601x
5RwXoDAjqnZpG0EHcr0litwvf4Ppt37PDEh62KQzfIYGeUgOAGzhbhljPC+TO7bc
V3IPZOMkMLe1zXC4SurpfzhdsMZtJ954X5s+L0b5GgqzZq2lm48hLvLFpGmw7On/
sIxHKksiiO8rmSXB4Qe1+ezi3kehIVPmuJIXeLRzIWghAJ4WwcxQQAEEJBYFgaSN
9hrQu+5K07DD55+VI6z5bNgy/+Vjfiyw7sN3Ty8+QEJ6+vvfebK4xUL6FodTRPab
zUC7H7/p19EgwvFnYmzgTukeUHo1c5xoRPXU8ms9fpEGmY34PjwSkaix9b8I4o4v
QwVzxvHHYovOjTN2wtg9B8cM9lXFbOyed8s3bFv1sBgJ24XZ++kgvgTBmsAlTQrC
Jebz0yBxrHfB/gCAECOE3Jd8a8OQom5MkIthTFhBMErsYY6JDGpHAeDo8Y2iKY5Z
qfpyqg0m9zbM/BSVJJlUb0wKYv7tgqeR9oBJO9hGAb3H9el3zeQf67lOVZIJCMzP
12G+kVg5OeFZWG+74bWmoYwwWwHqEeLtEUFLidI6cUpzNRu0sRe1+YrNDu8zwfpo
CQrheLuzyR95OB1Zo3bgw7Nr6R3cR6KOO0E8C5bg7s3ynYvgv7YXOvrEvhrn1JJG
GDNkP+bPoKX4NpGp+HABEvtKUONRElEWaXjmc+Uy44wlGtIgH2MaZ6fj1KddaPNV
DBUUhpkXsKEDfZqXEuj2BUMgkUtrPUVw/1boNUaRX9YWG3f2jdpncghu8tXlUM6F
rw+DUC1p5huYY909ws9GK/5nprLERVZSpXRWzimci/N66Xf6YtAs4hgPFt74zKLY
tKTDHc5CQudZMRP2oOH8G8HoKaUaE6+mT/xEbskoeNZtdpz1dlsKuf5eVmMngWGv
gqRvc9jH3/inAxxQGMNgHrI1DUfKlydcxDaNmvHRzejzQAysl2gtLqwWnAP2TOFi
qCdYuN+GUYkA9k/d8bfaasmBcd3Fh0J79wPKz1c2nN1FQKrsI0tZMF5Cc8TurBOq
cV+0lqUzVxU5/Llfbb7iwbYhBHGBzvU+/blOrLJ2WJUZvZqclonKcAO8UhgsmW+F
l59SxpZv22pFk9ddA8KP01n5F0O7uYx8uenKVK/F9FKNaTsGQd+vEFi0dW3heqOR
EgrA5zTJz3LUdE4asrrhehg3KhUH+JP+TMXUQNacGez2k1Bl0apS0BRyxospD7Sk
1pyi9Y8SU+VmNS0r3EsgedsPOsT8NGICC/ymBDeQgLlSz/627tralmiT7gE7GAk3
HZd4QFCY+ngpjtfL3Sku7enMC0DVbPtrljTdESjsK1lLWEMelPuHQs+kQOd2lutZ
yn18AYUdJfPuGsJ65RIgtlxNoGY7+3hmK8FgzkPsBvcrifaLGm4FvY6By7lYPa7t
JmpVpbdVDzrStsiw/rrS45O0jDWSWh0PcQ7qsD8r1qSnvebyy60x1aGvln+AMJDu
OPOf2T3M75188eZDnHIs4kIAgXRUC60bVk8FKy9guoP1rmOM4MIKrhlUG6kyJdkY
vVpyUReY+PuZmFEakmUrhKTOGDlUVpgl406Ep1gZQLCCO9BPR1cGi6PYuRMfaalG
9zfHZ/ThT5osYgP+FXhnhTQ0oPg0ExnXWxVn8UdDJAz3XavrcIoAPXtTtbXdFaDR
zkvlaktxzBk8hzvZTp3zJps1q0zTkaohkgv9ALpz1lrlBWGVIPWxXvV/4IlidWFg
C8h0L8MDDRgZn6N8o982HmU7khVBN5nflxzbhKEY0hR6UGfi1aZpszhDLwvClGKa
csGfUu9xIh/mA99D4TlO9M5qy2tFVWAHXY8x+XFj0sx4XfHgQH3/H54becuP30/6
V8zM2Scgo6/nujOqycYPntET/mW5+jI1m+BrVji62ABfLzZD5UrWB1zNO1VFXemX
MHzzC5HLGsvVySbfi1fSioSe+CX2MAe3Hn+nFmUF3+D0xFdr7/JdgXbZvLWZ1jF5
TZNxeOVrJAApY9zE+RNWc8abicypEKkp3MToqjzUpmzqljndo3Qjob5e5FamxgC1
30e6KKfAn+niJKw87sbCV6/cREsZq6PJ5GC5BCU0oTiybX4r1ccgbK3OrHitBB5k
nIbxj3B+fzNR6fbpusTY3xgGVKs5oRihmm9N7uRuNLcyEOEhKW/+BJ9rDIvgKe24
VgAaTriW7OvwlzH+eqIMXQtHngG3rNTFOCJsdq2Dzsu9gLm57GyhagWX8EhUehy0
qB86tCVcXiPzibDzPYME1UaJe6DuQa+EUfUxAqVe3lU0M1J3Ba+Iis4WgM3PvFHE
KCpWuRJR9uNn1m2dKNiy/9+n5UrbF12gFmc468RtT263uYUqrivugERjRV3B7MD7
x/DmHXtjQxbAusar4LKLQKcLwMcKtcbd1L1KTOKFihwqlSt23/gKHdhPS5xBwJZC
Mj4/xf/zgtr5+GqpSMfHpbrGQuxEf8ekQlK0oNnqzjHgv8wdbSFUYV16bJgd7GrR
oYtljDZpQTURwYcYL9Wgcun/PJcJKljhXydhYOyZNE1bHckmvkYI9bN2K+jTU7XW
TWbA32mIiruBM48fPvmXdpW4hJfKTxWk10TsAeN1/1hSt1Ax8cw68d8eJLDFVWAt
bivK+sljp8dPF0VwbDpg/31xR2Ij7fU1XS/Te9VRp0n2Sv8oLJALfuIJNUBVLdCz
9PmAFW77LyMO1zrSgru9UvVJ1Ly0IGsd+ioehfcfhhlO/LlDjOTNQSvm49/ISqyA
5fTBIVE+0Va5VDfX/snEAU31GrU9RS1/+TvPDslNOGRQvLeOm9zbGPXXZIQStrZW
9i6lsBw4IVMeMqFTDVhpOhr1tM5zeCQzWG/tvxiPDGjyaA5DHce1gwCt2usM+pMv
t8izpO6fwLZ+VzhAgmrz+l1R9NiV/Cn4fTS+zNtVxA4giqIn5+ywNd02Mh+NFQB2
Bgols7dPI8zAnYrdI6kt9fORbD7wcUfYKIeljGEGcqFiBlCaVHhSBS1jwhybTebi
yV4Y9sjLeG+8jziGCYV8q5v2YvHeNm5I4090jCSR9SIEkwaUhmM0cIXYVPRREwqD
w0VEk1lUnP9LTM+Ey+vnJURTY3v+exQifXFsTGvzgT/2uWY3rqkQ+lRm4r9ocL6E
O0PIgmP+AxilmpfG22b4/oKBJgjq2zMv3UGxYHfoGirwrnZwqGy9euo18YXmh3n+
FufWsXP33PBolesYowoGLKoOQNo9B2ZKOBZllMl/3wHdNh0MlKARi1NhqrxcUW0L
m3wsFS6Kzyh0dV2vFr01DxdqXYhLoYpRLqyK1qp6eUv0sAk354JOmBtLUKduy/qE
H4dS5mjUXSray0HPrUE85eZvn5yq3uOG6QgAvIJNLX/v4NaU89amwO5NZSprj4kJ
/oGVB2sBZGUQ/SHkfXA/j3RTY2nSUsF3mnVy6Oz0vCTZzqU5PeBZxjP0sE1VruJx
GDjdL5pVfb6FinyYnfMcaqZndNNB1toCB1kZ2vGceCUlVl8NhdOw3nPkCyX8hal3
g0HtwCyrYvUR5BLriSPl4+384OZKrRJxKOP0TZdgCcY0hRLbRgtRRy0fMFVMnnbH
IkmX2xLGye+RA6BXaPsFGbm1CgnGjLReZH3sfmJGpUpTNSyRyStJZ00Im0pvJcmA
ljDoYs7FBmzY5h1WptTF0rKMyaiK5DKSabwTILdNQAlGke32OOPsOSdxMZnSfQRo
k678PLp3r4HU4l1LSQY3OJRx541XJEhX6eQ/6xZ/yn3DKKrzhC47qUYmgborvg/O
8g59kOPZzn9Ou0LupAomZk/n+XD7D7Wn9qQUt4eUWFgGj2AfM086Rc7dQfTUtys5
e/x6SOPmtcSGvhvgw/y08fo4Gogf54LNV/HUKGlmsUUZgSwsggjNnHHtbnGtvBvz
T2GmgkzE32Kc29EWSrLUVyI/rGrQHPMQXQr94f3hr/HwE63vV334YCTQgyC6h59M
z3kmkkX9FUS8H8XCya+CxkqLQbIzXcQE91+m/BX7bzcIesuxBTL3L6tqoRGsUUH6
yO6gmkHsPKdvEbGa/psysG+aMR6/Qb3ppl5FOjr6sJInOLjvYvAI7FaWvY67sVaM
WjLAj4C72wK0yRrpbLxohN6mdYQjduOvzEnt5GljZnXhGt+pmXQScZN5oDyFxAa2
QeOISuMnLZ2VIufGfvohdymFiUcnVnqkbzuUCAdvnn6cgF/gXSBA51hHPKqSxa18
KoSAEi2OP9CxJ4+svtFnIAa/UxW2Wo8CBApoDon4WhlYX2xqu0b/6B3dt9kLmCjU
KEORIUAtaIh2BnauhPsHJwYWVJ9w0Vl57ffQEdFNpqbeom/lpq6VIG3begdjJOWo
Ya192hX4LDcIBUYoNMSrg4qDbBKR0izzvomGloi0VyuLB7MqY4iC7L86C5LQ8QSg
bvj31345i+YZUQLEAOhcg1KOhDyM8CKw0i4/if1zuq4mbRBzETrqIcH2Ve/Uyj5S
5bx5bnVle8b6NGq+7/MgKdWBC9J1x9FyORAlAgtW9ZJnAStmo6JqiGD5jDEhhHrs
EF/aEXfpYq8+V2JqC/afGy8mlDI0y1qujQ2SYmK3kfOcKirDamJ2RhImHj/+vxCV
HA/DDNEpK9jkesDeLxTlC4f/pgZu3DjjUhDW3G3kj1mG6ka496UHvJs3JqgEu/sU
oEeP6bwk/mnZlQWM3el5vwgL2hc6lJqboAJFp+WiFyKca/zFp3fsZ2XpsocsCeFS
V+gYsjuoc2/O+D3r7yGtzeF4TMMJtnUGLtoSZ7lOs9OzTikEtWUkn89SJVFrF6gk
RZ+daGIbc9KOtDINgB7op/q20xkop/7fyLJy02tMXUEmHKpUbww/BwzIvNp9HHCn
aM2z4vxzhnF2rblecfWOnYfo1puE4ypQ9wmifwX5dAb9xHB7OiEz7uXX9zKk7TkE
yALoToGYGEMRGWeCXX1huziNeSGxfXuE3bn7e7QXsM/DpmiQ9M5e+GxJhr/PhYD4
qj/4TxM37ayoC+butJRQoqAzk8vTp3gBz/IkrWSL9Njk8wxeHgh52V94mnooghsM
6S9g+MGvvTOnaFdo6/YEBMv54mB5BTOnVJz7gT5ANrQz+2pVTig1wxpfmqu4qpKb
RDiSRKKyfYFhRkwxfxJa0Z3eHxmfAIXrxnJFrBWJrg42HZDsf9jrHSY3fiFJzpgM
dzivz8jFYlvFyTsYW2m+QN0xCKYurv70f/i0k2RkbAmXTZleBQmVLdfAhGqaNyCW
2g5N+cMVY4C4+AtwaUvlww+pc8pZh7a8LTpmJ94u3QSSy6c4JlklmP0lMjipHOBn
okk3TXS39tNl6diXI6+ont+giRpKeY4jgqYf7xCbiC9QoVh+y7dUhtCxxNqMSKlj
V1JEt0txG3TSlwpSlX46lcogHomYkQ8jo8wgJZoifRgWge4ea6qnnbbN3DtQHNdJ
pUjXI/v4OqBp8b0dWhS3B1VPCS7cuUT2U2wZLEtaHTG/Gz1JW7KmSsmjaAqeUocq
g5V3A1KSYB5XgryEsuSqdmtfhJnemj4V9IFOP7ElrgUyPuVfpiWPAPag07irgoFW
9lVDaEU4oRJkRBiPUHbePWQwgboxE7Eat+2pVIYenugulAqk+I/kxEvlhK1xnjAF
AxW1PC5KHtwPR4cQRagOH9Xr7wgs71Y7jDpStA2V4f5ecf6/kKLIyr8hUaFHxzbB
lvRqOlCy4e6nBCJOQa2UERfbnkceIPzzkH4uDowjCY6DNMnNPxx9ASy+Fk09LIAS
mZEa4FM9zpB3PXLbR/uxWZDqPtpXxctUnut+gpI6Sip9aSLtmIuLF+SPfJ8Zavh/
Kw+QskL2locFtSbyg4IE4itIuR8NIpckU/w/noWoX4YBCpyPXJFZHIhAG+KtUvUL
BrGLsNtmpTKHPXU8ZF+qDq8uaKB+8zzFzbv4s12+DXBA/F96IyR2FQe1Cohlj3AK
jL6caEFjlQW2KfgUEOvjENiiky20HPiG9CZy+zKay1EIqaRFnL+sxHONcF++smZn
tt3KerggpztxrxgmUvOvqeoLf+8yFf9IROah5PFu+F+m0F2qB0HZp8tnT/nJacDo
lsUXU0aGH5Jl9NKbSl/1MjfGhckZNMXsnpfuvISwGYewBcb7691WKyOsLoiyqsgt
yU2lBuhBEXNER5JjGGBm53FMqTy8QfKE/ITZx4OHGtuvm2njDBZCnUvNJnHUcRKr
Pgp5gU9dr3MdClW+3shzuwi0FNzFXAjC7PqU5XK6zFrO5UK4kYRge+IYwtDyzziW
fTk3bw2mgjni0mA4wVYHWpUFJlHgs5aQKEma//nwHji+lS+KKiIRNPqTlKnxwwiG
CynQPyaw/Nwl9BKBljVmZ/Mwy5kkixqwd8YhywTfgvr0aOYs0/PZ8Qsf7Lu2nb0t
zf/rjNNVuoWQfVdmMg+4INrUXZ9G4E1561SDSgypK9Dnkavsjz+pYtyMMmftKaEs
PlbekrAxHUJ89EPK+mfWHkSYmTpNMSH+dodsP4oRltbYxMsQy3GDdi8gt6H6qCC1
KJU8nT43Dn4YP1AJqnL4F7ufw6CkP+FNdxwKbyWtyYwDhdzBAELrPf/cIGdZaUKh
4as79U0CgOMI+b3CLDkmVZ6jbv5E0ITTyvLo0wvrjUwtwpKsJVDv1IjGlQvcxCYQ
0D3+zRvAhKx1I0KsKm4I9TmClFPHQp9UaQ7fdNtjCWLhOjPd+EL144uokww6i/6K
JtpaoZlkhvQxt5eR+JTU8nnZSShhIDG8vJXUd2/kN7gX2o9SG0WOIQqOosvuItD+
LJ9YI04rPJ1dC/xMlJ+p5JfpTRndGIcARzBf12npVKfE0WkWO1Ddkts4wuJTfAV4
yhah4wiQf/uqYSYYDXMVIpszVq/my0l2GFsDFgf+g9SiJHvBfKIRvNOl1K79P2zV
xP4kUSLDCHKNdvSZcV48CbxbfcJjvtLWHudFMBimTcvHmY6zbExf4hHWdgPfsSts
eSoV0Wewekw1+zqE89NdHdxORHt5iQqhsbwXmEwG9vRzLzKpfs6ydQ8zxBYBW2tM
aUGAlGogqnu/gQT/IJzyrFxOFDxk0kEX7V9N/F5W8OrgKPOQtrzPBdiQAcrB41ja
Y2n2a5fnG/1FcIW7fGAaOV2sIcSH2RyL8Z25L/aHlNDTFsqMPwEYuTmwpN0B1Sd8
6WIaZcd19YOJQ+wnV9KvQCBG4xBC+r3FH8vh/MthmwcJgBXEEVV9lOIw/yBWwW/e
9yEHaEZDQ9lxQhEMLK7R/G5iP0me9BupQWDXmnfLGDMRnvlls+UtJPqsfYksA8f2
u35AN3xWhyaoogQ7ry2f6lenK99w8RCPjfteWC2pFithOgZCi61UNV6RlblnK0QO
Q5jMIrpx7SXSqlFoFdGndB2BwsF7eCpO33Cvroc6M/laE41FTjWTpiExnxtuAYDG
5FWjYyhbjHoF8LceD4zyVqSjzEEobe0Iv0BiFJ0OJgQSGqJeyXEvoW8vWnbZvnAn
bqTLVC7vxbuYvR/JetNwVz7bnOtU5tj0P5xYFNlHNK+keCULTiq9r+mXihNDEoTs
OTlIqypmwJgupIKAZXw53O0PKhcD8MTLakrmyEzlH0JEIaEfP3DUOrBufthgRB4R
3c9TDqaXiywhT0dCIjuaFQishtLrC+zh2NTBd5+eaOOI74bxNdS7qWBijzZUo7pS
aexUqt+aDwh0yZWCTcACGGXBr8ifL2eSjH7vrrr9qY73iHN81z4Z6WCvZNNQ6zRU
tywtU4sYVHHknIlE9uBZKA+jb2pLLa+yQWUoKczMh25eJn4xeydwHsGg/YndFwn2
B1OVBUHmve+AOHws5WzCyjntnsSELNCdbB52j5b6EK6tOvPYgxRqJhZzZui35MIO
IYgBRf70kRXOl0Y4n19NoIF/B44lHjxID9Z+7gTOrMC1DNm82U8zyXTy6eF8fPYs
AQ8pCSai7E16xEO16N75oxyUXpGe1usx1CGLFtgphpHqEQwNKz3MsaSw0MM9yNNc
tzxbR1gcdOBgh8pq2H9T3tYabzBc+E4Y5WiNhiM20Sqht3HItXV1lMhHz+v/UTr6
u0E4G8O/tu9HJho8SCHNiTKACOMOVr+rvca1geiKt+0YC/HgPKTPQDYY9lb/gneT
c6OrxN9PBO7s+Th7lPRE3P32Mouenq91hs+B1Uv3h2ZRmB74cfhhYX/hbaudL4b+
sq5dYKqICOi6KVNe3xJ1f89QjCuFaNrk+B5XFiEWNielStgwWyHdPkQrTBUO3QM8
96BcfLSTwtbOw6x78I0THs0x6Oa9X4XvYSZXGOXLt/iDEe4nfd9iYiVGRDaZDTSw
nW+dluDrYSqLdCBDINaQKykyNIjDR46Tg9lWTOr3fh3FZspbIuuKLb2ogTWEvnoQ
w28+MelbDEL6lDHmvvxoVJ8kyJ4Q6m21s63oN3Lizfwguz9Gh9z0gEqz5qiDCYyR
4OdqyDoMW3RzBN2Ac9YrVwXvOn3WRRISK7t/vIMblRyHEvO235H3LZIqkb2aoIt9
A/jQy/MnG04Kv3r7JMGkSeDrJEDdix5rLyJt8EwOp8xZypXsOlsCvR7M7mamBcgF
2Meq/dQLKtQ7I4TRTo07HPTzriSJP0zE824FVQy4GuV9KknwV3Y6g4i0IM5VyIt3
pxdzq3t6LZD+9qUWNGtsKS3e/DKxXsK+Ik+OnCOrZry9JBswjnT7tVSREEgk4Xdt
xpolHuRSXooXaiUCkb+jCqe/wIYQUkFSiE9T8omZtprGvADdDGeEbv/caOnBI16k
Tc+0LlnpHgbCCwiDM6Fk8auQLcA+lxR7q42uM/9uNvHvFiwcSL/CWytwW8fVP0/m
9bKi1b5bCpRkm/q6uODiRHtH78w3KGaTPBtEHL4Z0+EBAXw0+Epz+KZl+6IJb94f
TDmdf0l7pnBidvitK/H4eTuF2qJdsTjVIDhPeQqNYsZHvuAbcZsbdDAHPCUL3U8w
Epyi7Ae4ElTaSBmOf0W6OykH6KjQjv/Vys49Wk2pJlkjFKU+OGl5f3LPgkMlAkx6
4lcIelUJpmNB5pCGr7XV8sy12j/i5Q0MkFhHIz3GGii3AMIRwXZ8b/ssQ61YG2+2
RmAqO43Z2RsnIjKihuk9RDrcMUWd7J6gacCrhGVi55kXzrf0Bym4j1Fj8mambfL5
2SDQN6f7UpA0DjN1tUPOU94D01NHi6AzHP59j+KNiYgR1P+4lfna/g2O0LiXTmII
yJ78vTuHyxCbw2r9YDbtWAP0ocHFIvC54YKxAKBKsRPqngRrlnCpNL2dEvD/Fsgy
CGSxhwMNnP/n8wolMUsFUkDmsJ1z55FEME9wVB74jlJAUUUzslopmj4t+f7U/RSW
KVpzJ/5TdYTU0vgq60YnXVWTXSUl+r5rJz75cZd08j4uL8T8z8VnkbpRdAodSna3
NzLrM1LLv4L/OkWwPvVS2oenFwBzhUNqgfWMFMON2A2y/piWnAyTwqUFvW4N+KnM
zY31jkIUZv5b+UNYZIxWxMefYuAaUWVfnVQEgu5zbS8rGE16VqRoK3kzFGNk1s+i
gHJVWYrOXaKTOMHqU410OkVodbs6QDh/EpPme/ZqplesPsr3sG9nouZo473Ckjnd
ngmeunxpGCZ/q+xwzQdsE2F5DocpVbCXHtfSia5nhVR19wTPYFTAu2mYTdnJodMp
XwBpuXBs8KNK6x/amhicH2Yow/4/a3XnvMBCr71GirKS9uNOeLTeTQfN5WafroIg
ca70sXmgHsUUrgpkynhX8vxyqVe1bPL+nNTd/h7hAnU6TvWynyUVm7Wrzboz8RhU
0ycx01Yhsrjyd5syFFMrQ2gVfSym/mDbCIx4Wjsi32QNsLWSDkQ3H/0icuknks4Y
YRXwCwQPMWrkZzOVfD2CivUiK9Nwz4d/DETaDbXXPNe2ppxWdzmTgx03WZvtF3qg
7iJfPjktJ4mLqFEYUAeLxBVD5MgWOCxED/mm5hoQuaLr+Fa+ZywsLHhavZqP/e1M
D+M+u3ZbUNgS4QqzlaKm4bAE2Mu0el3CAbVqhMGN8R8wzJvZX8yZCPN/tYkV+ajH
E58rmwmIeE+83xD/48UQ68wrZvMZyCkX7R76ANLdPwDeoFQjJsKJIhDNiBJkihlU
WNPCytBxUxsVNA015DaFVMN4rvleLvsfY0cp4FcB61KYHnRjEQLEFNsihbOENOQ7
jmyZXkxbM8sc2zU+2Tby0ovTGmmIj68IYVGLqSMvBzg1y34DBO6PL+aNTyrlfkVE
2SmHBV1y6ixKswuAKwreei04k85KG2iG8FEf4AhqBYJAmijE4dWUHoO8cO6TY7SS
MnnEwPzvmFJ0pKC2gO+vWLuDay5nqPboqCxoyJS2A6PwWL247ecp6HcNKKlU6Kji
3z3+Ufb5Lc5XQxlnhWfsrkVHTa/XpgqQl58laflBlb53XCss5L74jbSSSMrgUskH
qnuydfi9+Nb6DNbfXqyHuwKUVsG/GXCBrhn1IyAMcAl52NxAkw5pHGAUbG+tjWOS
3/KY6gFU31AXf6fUE6L5cMY9bBzFobSTYNzY3hjROYNU25Gt8TA3Skfb3UWGbvT/
bFDWhVpf8pyAJw0l2zB5lh+21NJVHS3ILrJv/8zg19P4I53Ps+4XLSNFEjvzPMYU
3sX3ko/YGlIdcKQbiWMaRdMtIP+4RcQiQCXYoNLJOafDhQ/kOk1yVfhS/qEh2rFD
4716T55FiTUoBVNTxyLtQC12q7nAMPv16pUCEDCzWnC1b7XWC0ul/ezbcBVs+P5E
Gr/8q93NXZxLaoiGgSkGX3wBaqQH5+fsa6uBPaYqjBySl5bMHK5inUMqTl41DsxB
nE+4KTXXzrO1+dQnN7L5s68WnTK4l86i6kOd9W49vQSVLHpS8wft33ZsHiY7qvQC
DQwbpV8ZmdM4Ic7RX/WRzdSHn9b+X+Ta4X3X5WV3rwmKVKJQ4rOYhk1oIR5R/jjq
ZSN+kloBOkW2p7EniMhYgjNXNM/KkE55N5YC9cW2PJJJu7bcfxypiMHAo5gkqRSR
Jeo7cVixoRJqzpUKbTiLbOdpl/4/KduO39zQi7xUK6DABeCyhWpuNkibpdKZ7Grn
EN0ZioHQTjwmLXJ0PvNxtzKQK7yDn/m+OhK8RHJiEoKxk1VlHFTAiHNiKjwjDQiz
3TWM8lwfqOhiy+O8zvgUTygtNv1Z8MUa2MPcKwbu6B6JqXiKlXDhmF5RHZ7DBDDY
+9yDlhHgThqhCVjQe9Ug3JOj6ExbapFNr/+ePLQBiMAkFX2I2RdPuLswGBaGnWDm
0FZGL8W2+JsYG/HIeNSJgNO3JzC0ebEPQVHCH7gB2125aPlylduh+WYKJYqNhKiR
o8cCY39A31bWBsYZ1WxkNOJ/qqD+Gr0JXbP/ioUiP9zLGIw50fGXFppuhReOMGHG
RsLdPgl2dwpI7kqyCWt1xizfyqBEXvwXFJdSlVVgGkJ9Y3G4jbNZFS8ht+xUX1kz
YUNx9IaBceF0EpPRT09j53UWrzEX3N/Oy8mA4i8F59Y4NHUlyqERb0l044UsxuUA
Go7gpwHExl8JyMpU+yMtNtl9JQdeJYlLddwwGSi0yjpTrQrhZ+ciP3Xj0WFQOhnP
SNTb0bRQY7QiQzcnF6y2cQKHFSCnv6fAC4QlTj0EJB5zAfA35/0K3ETRN46KTeql
SEuPzlK2BGgDZkkQZaapyk9M8ccZhcnAp+cewtUvoJnZNXYw4XWNBPriBlEuuceS
be0Acm15hsZPLGUT0pXlIM+ZAxB/KJdEloXqG4Kdo0cZGiW3qObRY63jbrCuWcAn
+vo/qHCKNjv0BdZfod7ai3/vrNNvP2BV43gUArijdZc61O1A8b/1DVyEaeVx14yl
rBEgw5PM4ISs9lzh301opCQn3HRG7EIZlSRZSCHZSVnZju9DdDnKJRbEjArpvNNP
NsMYRWNghIJpzB+kH9PXZdYFLg2NcLaB1b7BecAxEUDKHBDtPrO8y5HzG/rRM3u1
mUonVDhZF9zTsZSe8JqbOSt8cxpgVr8xVI0fLvEeinjEGiRzRyg7vSqeG2Dl8LZh
YgcXQ4VGcodB0AwfQicRN/8EhTvxaw/9ZaCpzfuBpRoinDfYqnO5PMiaL5anrqNY
lsgIcVypjs0dXhmCzRnos/VeQ13P8sKzHby0wIIgyGCiIA4X4ocWa0btg+CDtm3F
tVaLx/MJBZIt5u4hqcYVDdw8CDCfNKlUZUyQgjLMZuZROZcH6SazLxJPkujKMjLp
bHMkhwfUJksTfscVfRjx9ooY79DzwX/z1A7/AtTcaUq+OukdB0/8FaIMZt19Q85n
IQESgx2qzJFLNKZRUrMp8njB/92ITFuY+kuKohAiR8f1TSx6/6kFabb+SZNPS5Wg
JQyxXctzJ83cQ2cMHpRBe1L+7ovsDEEdS6/KVGHSZac1f2/rxCi1VNj1l7MIHFYH
jCUlJYl+y4oj/OqHeGPnc/x+HNN5aMcLn418h7tT14jI1DONNN3v71Ks7qjBtYf+
B6mCTuZAqAQK8UPNnKS8EbJj8FIPLGgqdH+T4+Y1qTZi++0j/VcEYrmkrLzgh/W+
52tWxqAhz47DeFkRZ34Bvt99dJghJROI8aAfdLgV6ArDzp7YpcFG6lwl4sLg3T53
vLYRcQuYABYhnUMXWGyT0f1UjKGIVcmIyXj9mTrgh3JmCxA9XPY6exPx0xeSWn+X
90uFKIDvWdJNdpoPBtnpvxW/eqf5KIUWGRlxj1SaqBbJCE+s/3S0bwIlzNzaENv2
XVl7O7MLXD/AsLmu7iuIiD1eJ4HK48eZUaE6Tlu+S8vLr15sGRGEWVI67eCwe6Zq
MZkpsHwwlV4W2dvyIGd3UklLAfMUxV1zHvB3wPwrXaRU4he6tATDdlBrlt4VS6lp
d0Sx3ScCUgxQWf6yAMFUY2g8D3NLAiAZ4NDgxLV9hXLxoF6MXkhOiukYIVy3y6uP
1P2tZnmo0Wh7Ji467wErwYNHjQO6QzTn93+T+DQ3qtceQLWZ6CZ0FEjoIOQyBvBS
EGE9Wqbw6h58zqAUk/Q71iCj7Bwj0mNWEDshLlIiUtzexCnIJCXdn33Mp7bbhTgM
8yEXIXVWVNceiBRjhDx9C9BBIUCUgvnt2zunvWrPvawIg9SgkX9+9jZgM6yTjGj5
mav1ukC7cv/KxmZGVF1F5SnTOWHrvaO5JD1cxCQyxEk9a4wcvrTbF6TkhxZnxzRF
8IQTaC51FbAnDh1Qkn3eJ0t8TvQ0wv+nMXJzQRscnFNMHOr6ssyc33ZHDc+is5JW
gAEj1V8jfL/guJ/QapmV8BRetbl5A1JpHq2R5gKkMHtYzofk/lPEzRlm8DKro/HO
qoqusvHnylA1PNsS6gdpHR2BNQlJ0j5PRK5o+bBKTeDV8pplDBWkv08mwPKtCAhX
aELU+lWga8bTR8aYvCfUYD9LspBBDX9TbW0NlgNA0mO02iC32cSKCLcrILrl0MRL
6dipBE5yiZJahWFqAiU2pMsPxjRKNJ0Xt4WZIqecpE2xj8zUWQSVzGLatDn8BXgg
wAIZRAECknvfwnYDZ1KMorpXwFgdhWGH3ONIVYfUafQqFfUHSx3y0WMibYkUaY6N
9ToYGumFEd/yAew6olGkVr5ENBhIUquHAW7Jz7N4fd3iiKefxNGDw9y3oQHhUHsK
FUMOi9ng+BXhSHA0BeeDCn8K9tj8eVBwqeZyIxTu6Z8AkNHCo/jewCpo/3UNCb5p
8doFRmCDLNBzR5si5WpPbYsFy9M1gUi7UKfmf1tc/8A9nlbaD6wTU3cvHbtSbAfj
eXW0NLR7izeeJ594g7oDDY6QoyajpULg++SxbSyKSN2lVLhAJIwGJsjjO+itSMU9
L+67pS/nt+tDcM+qtkuvb/LtQX//cFWUJgBw0eVVEhMECo75qk43HW9hBPICrXwp
97YYWhdbyZtxx/4u9kGRpRh5p5vnq8C5hew25unI45iMVhQyT8gQ16VhDkIno+ZE
3dYi7vnvAHbRnMWkc56RIy+vn+yeXhsnfs3en1auCNermW4xeuX0NIjwe1edqbrf
KOb3lEcejbcb9W1YkNQszFlU7sRO2KgXhK9ie2SCKyim5sh3jfBnz742zcE7pBOO
FinICpthiT667khcohs6nv0e0Pd3CoOsAefPNo2K5E4tKGtpPYfl5s7ZG5aTM3S5
W0D9YphkR2uasStuVvZUJlraE4z8vQrfbL+iuWHeKImqcPj/FNmqklyIJhfGRjMu
4jOEG4jlY8ulf+jupclY7zF8miyqafrh9IZ8Ei+GXobHROzsTYZOEQHrICMtENta
feBHjH6FraxP3aTAxYrGh6dBm+rMC2MtrcAPLW6djMakYYGQ6wTsQtXAs9ut+2TR
KigX0q6lak82sbdbjalJjOnwcTLUBxcgHR7j2R3PdLrbcunqimtZMT18oLSi2hSQ
7v7xlJsgxAIM86bqoyMf1v+HAL69NjpxtR6xHXFO7GMcv20EjXBQrfOb7lBEMtZ4
y8c+68zvuhbYgQAlpAs4IpH6q33i735OF1ByaHlD0HYaKJCMSIzZB/fyUWr0k+sZ
TxIrrL2+IAQqEzBY9F2Nk3AxFEhFAvRActMuoOJFoP4FYpVkNBPMaIeVpmSS4FTx
36hTtiIYoxOH5fI16Ho1wrUWf1K/sJuvkRNnP/nGr3CpVAEdHZiBsXEyASP558hR
egF3QCrTjN5rHTjgs0ZWyZ2qQn0snIw3tYy+l1inghueIkPpap3TZ5AUPmczs5Ww
d5oebQgG/V73Q05ItxnVxh3YC6Ta9IYjkMThzXkbV6i+3h69nnqcsBr9m+VT4eH8
XEHb6V5ov4+CjTgbeGprRPB+iZ7QCdNGmq0gET73rErF9ocn033F05oG/WObQ+B2
qf8oiWl0Sp/8MnTKJksXHF1MEf1+04/FgUSTRaYciMFnHoEuYw1a5Skz2Vk7ianA
qJv0U3nvEtIi6AJ+X6NI/E6CCqtKS3af1CCGiYDCClXfBRKVQ/Xpbcm+4WDTwAOJ
d34+HEmGrguJ4oGxiz/+d73gIO7Bq+Ph13D4OB3mSBcvSsGsA7cgJL3HPlWuRxxv
zuYIJFLh9CNMm6C0NADVNzqJfPIAY+LEL+hxMGwmts0gR5YK3NDi3Sllyo50jFcr
N1SQ7NDDfMFHAtQa/kCKpJM7T7kigFmveSBoSsgpY+hYqGblKbRx4TjWpn4A8BH4
NXhsD0o8WlMC4lF+5LMW1lD4Eo/C1I4uBGg+4L8VHRi2KmMAhTSs6w/mc+b4/dee
oXHof+6t32Yxujri1Wofq9aNCaeb0YCMuqnFGMWipStfxp9jEaKoyR00Qhmbjy0b
qJmTGZUXyxqKIWfUtGBnmRzZ9h2uLKJk/Sh/2ZoTSSTnfIb/gpLXPOCadiA58D0P
53WJyfzFqak8feVKpMibNZbrKX45AxTZtfClscL2sNqeOFJ+vNKEIeT8sqjPd1Yx
pQ62Q7PUMzV3X1vd5/GD58Nwr9ebIcQgjQ8fH46irRPrRl4DaMAFrpKd+M/6FRw/
tqLZQHj/+UPyuiQW5xZ1wfTFYDQAcYLxpysdGoQVr3GO3n4gm5mcus9YE8rsdfB3
9DAl76tzRZHCw3jH+7Bp0OPgh0K9czQhwhFKf1+xFjevbp1NJOarHvRvjPYkuNKE
6uTgvWmKwjaaTAEJHrm+eVImxs/soL2w5yDOSw/YOzhGe1Kdr/MmJnLu+K887y6w
yUQiej4K3nsBBj4FNjqQf5Wk+/5fMKVVFJMsenTmRE5hhccZ1+6DO0qDQxfzMd0F
kMieO7OYE8dqIKFsLcmHMvbpGoJPxomNsmIplHPIEJmiP9NPnyto3CrWy6Zck4uX
QlPU8rF8jGmgwVVX8XLmF81ATEvRki0aMP//aRam3cVOiC6KQzODOdUmEemkNj/C
wCv7p/zfvBQdu1R/69fyR4CHekpdhn2wF1niv7DlDXO8pzTb8gGsYs50w/14eDgi
R1aX8cZ7zznhB//UyR6V/jt4niAHnG/nyqW9tqZdNJHE4zngECBPG2K6EMm5Yn6t
D5KN7OOYcDbgFc6UOzKd+9jyvAshB1+v5TOi2yamRFG3NXUQvN1Mu5HIzgxgi+pe
/mO/sAEjDyyy/j4kkEfg66JSwRd0Qbm4hpu0A+lTKKfWa+y2hqeOrG/5vEc3KQJO
Ix4ofw5AlTEDq4FLGBh6fUN4Z5qBcODFvQWgqxCLIlriiIOmvF6dP7TdpeJzfcQk
JTGA4ksku3ASqMsPNAJ0AHSeL5WKz8okHJFJLZSz87M6lOkKnkDmY53xJVRuMjUR
vBgXMCNG97IvDPWEAKAS4wTSGdV9yw0zv8uaLBKvO+XN9zgcpgZ/pUs2r0X4e2qS
On/2bHKPDhYG65Rw81H6cJokulhN5GPGeb5YBZK8d2EDZ5IlwwnW2QtUwgUp+2B+
HWikBDamG144XbCnVIIsAIIJ1z6IW/cHYlG4ksOaVNxb3UDB/VYl6h6PXrdRMFFi
NnOnajOuiVqqRx9tfRBwe55tNAGlhR3Ue9tM7960I2nMneCSa5DoFVIf6UX3Aqcf
lgdxLl0iUka2e4HbysiDXmE/2B3ooO/1CwKjy/mQi/wAHIBrdENbg6htSKfMFJKL
siO18UMSEmMjG2PmI2Nj+UrGG8yF834y2MOgRQLz6b9DZEiJtO+Anz1lWMz15qiI
R9tR8Cj3oZfBAYJ5q9CjJmdOYybQPp6FVH5uEvggFyS6Ln4RcIkMe0W33IgH4enr
r2Up1o4X3srZ9xObrgE4zOlYLAbrcXLGDD/p62mkvQjX+qpLUpPdA83jWWR4JW5y
B2sUL5MqZz90+nQfXaJATcyWmuyTro4IitGAUHo+WrW+fzwMzeAgRfmtzh+JnxMG
d6xDoJnzF3jtwblNzHki+H5Rgnko0F10TtyQiq5mrLl0ybbrDu+MI+M5X97j0yGh
KKNZ4DaProWU4KJeUpZuXWauVfgg32Sh0xsAdIyzniYESIZMsjgAqUA5ZUSSGFoX
3U4j0OpKFaa6sOo6QYSmU1bsS98LDC/LaVFn+tER/Rbz+wgMuxou4iIaPGJWmflF
d5OdZiPk9O49fvz5OsIx9+xi+L1oxqWZUyZaK/zBqcpGYuV4QjjjkwbfwJEOwdSH
4J5U1JebeFmzlOd6JZST2aOq/Ve4suaqF6wpRS8mcKPsZ6np0LjvxZ2+MiDUx5sA
+N60CXJy9oY3a4xkfQzX8fBKf3brSHqYoERbZjnwbeyS2gcY3eA8CuXXnwSSVEjY
nGmYXtyrr9Ob1vMBkycnHuZfy8hY3OnioC+OaA0Nd0NTeSK+JBX+g9rbSHEWOFDP
Xhr+zQhbruk+wYyFAafhTxSwSBKnkPPS6qKJXde2t5tV0ZxacP++wsOvV7o7ewXm
+PPYJLlRCgQnMSbpAD6Kt+A53Zra4KAhNDVmWQ5Qw7EK1+SOeFryTqdkZ0dm+cVm
zdkPsKil8+E2Kl3xhH8KUCRekd69rL7hLWctF/RGl0mikNYIRJALuuC6SAe1GYQX
z9Fq8rgSgbmE2Vtm0TFPANjGgN9IcgPtMsGXb7cB7QXA2ltzfNAPIOwff8vWSEDc
La+AM7PQNZPfr1cbRK/fXIF8Tobqix14qQrzJmTYk5brksIzhiZofYtVoElWM+Od
JKXHu5UzmpIX7Xp02d3nFd8JzInvuyTSFJM2rmKdiYSHj7M9+Cfd36hXw3CKT6SF
m/0NWOMka5UahrElEn1RtCmxXmbHuV5HFgvn99XZUGX1872E61aWRZ6Wbb1Kxl2w
rVMXR6HcyegMbXtyzawb2yBw2bJKweBqqW0yydIcr3kgaPGU1bCI/HQpFzer23Lz
eTGv0lf+wUgwekLyjfiOfWOM3J787d2BzN+FlD17ZPVt5Jb0V+bf6ozfuPnOE9Vw
6ewQzyaQmWmswVmJUb4YjysGJYESgeQkYL6fO1IL4qqFVTmDjrbT0Limxe7kfKVk
BWUEXL2x3V9ofSX3jRnW3wZuxNO4JKDHIYDrORVM3H/ihCbaoZDykIUh/E09DHLP
fHsgSnQQht5zhvxq+youS8WhaE37thOaKVxOquBTIs/p8d0MwJv9VmmksJbwTkY6
3f7q5pNRuJJbkgr2x2qzrGQKQ6vm6tNvIkhy0967UqQEwe/sX9K3erEUuqYxgNZY
r4lIWXCXEWn4v65Y+PsoH0UopANEd6KWi5hXEzCdl84wL0/AQ4qO3PCRTNEx56Fu
PS9AIv86KKhzP9zTwOrcj6wmcrB5EtB0j6nz0XRhe8ZH8T0q3BnCpQZ0C1xfgvFz
ubCL9EsCGs9D3YEYdVucI47JscB6ViG+TRhN2YgxBCZHQUubmvI2/WlDEUDry2+G
pye2oiHXofaRheKKQWgeOXOff4W1I/vMknXsjIPZqu5mxNhp6Y2zjSbn/5DdmDtl
eiXtQsdOCquWu31dy7LF0ii2dOXISCiV789JE7jNQmI58m+UA6WRYAa+OetL0aUS
v0kggnl+lfTJq9rFvEgzNXN+3SKKLrx30eZqjmwhcEJbFU9jaQ9Gke9Z3hDo+HtK
zVtSQw0O9cF6oIIJ8vuERxH3TRb5d0Tynmoprf5hWl3auyk6MjuZV0kTzIji/LbG
CuQXhAPHhxW3pciFKwWbbPdQ6vMN3vNSjtTqHKUU9dlVxc+1MJfZLNpN6AGXIxh8
FyLUcjm/nlpzKYMbHKB7nCwODEuWDlulcTCnQPXFK5MdOblLrgtyAsLFdkEBY5ps
zdhDvirn5WbSIl/9ks+of5GFVLyJu0LTNFJzCBeEunsTrGdMbIu8k3kLF8T1GZhr
B/o5eAspanXh5fR05B/Vsoui2tDw2wJMBunTBMWXu366Qum64G8s0kwb3G9anebz
Cvj9yS/Kwo6pKyFXkLnP2JpzGOo+pwVrLapHiD4QYIDJZ9XhHW51wbcglx/FMb2F
aJQUKvoRFVmciyKWYhf1Obu5TLU2MWyeScWMQCc5ZLmBB6v/VS6wHEnmpsAzxa+C
nZBEO68d+UXWu0u4RjiPoeA+QzZxiEMAUpHYe+Uh8H9nPAqtfdIIzK6pHeT458lu
VEg4ESkUTgEb3JuSpOJYzLNUQBdHOrk6sWj+wDMNSeIMQRv4V9NxmkkepiX/EBzb
tfH75/oWxZLLzsBLZ7LtpzRMECAjirHPF4LIDZezDiRJ1Y/KtNrxVZdFf1Wp5G0l
ibQT4z8VAZNg+5R3nD7fkcDIFs/i+GZZH/3TcpuzN+TTqdQNVVcGt256juTZ0MED
2HWsKb6ncY/lH0OLJ5sxRlAgZ1VNnM1ETQ/9M9CD6J88GJbEiU8v7Nq84xCi7i2D
7w3RM+VVNRRNNi5bSdJkC9eZb3JMWRLqm1KEpNOmLH7Hp5kk1pwzWyozvLPTkdOb
HGvdDCFE/w+iJAYa9JIPo549QtfHvDBN3q82daMcY8TSwerxsp7XtKZ4qGYIlkN7
mnwvZOb3RLngJJiAeuiYbpugeWWtcnuTyBYY/dtuNu0LsiQeAEToDGBzWjx9RyKs
NG1bF4ffrnML7mROV0pKFhrcSlV4HLqK6CMTfsb66qNq4oqUrdqE4n9OnOo5Lk0I
/Xleo9WxcmRJOHzmkV/aX3u/RSwEtG+hh1iZhZqHDkNpCDnj/0Vm2+56vmqWI/Gq
TCS7IXsI1nL0hmxODp6de20bw5VXXbQKhz4OB5W38XaqkTeQ0KNRDmMz4WzW9Oko
WM+2LMacW5mC0jTZoXMSsg2S1e/8xfXleFi/61cunEjTQ/dFBobpKCP54YBg2eNA
+wb8ZfmECth+qoxC3b3cvGclb41MXTuz0gt41xtz0CeO69vNbBP47Nb6eX6Dy9uX
s8cWkoQqLo+iTAdOn6inFKWnr5XmBVt7KCF1+UHYZ+YqAeeUQnNpebe/fIxjUMek
tD9y27PVYJB/E7lR36ZDo4EyzZfegQMffvpBR2sBmd2n88tROH7BeNHQ92LXJMiZ
BPYfDg5F407TfSIUY204maa9Q2JIO7B6WRQ8kZ09fJdAqW2BpsudUyCtSDJe++Xa
Kn/dgKL5D3OqjEkk+XOBjYQy1yMk56MDYzd3vr6ehwN+Mnd2J6OKFNlZHwA74yu8
g1kgH6lH5xL71eLf2H1rQFh1vDpX9jpMbmSyOj5GPs8MGagDa0xE9Dj8aNQXI6J/
W3QpktoBwctsHyaJdQ06BYfhSA1Sy/p3Z249vA1ixhMvk6fdJ96k670brHGwODpb
aqhDjL6Be+HFeQvBth4BGkUaF9GqNUncbd5Z9LqAaL95xjVM1OHvs+AYsv9Minte
tVJM33kt4t/XVWI0wrG+LdDGJEFzwLJE50CQ2GGQI4gvWYIvV2nXhSeXDr/IU4Hp
Lk0gRqLAQbNGzGQg1QkQTwqEPw9KqGrnoEmmoIvu5JwV7IlibhEh5/5BS6LQxD2j
yZ0MxsNaVHCNlhVDnLVcwBEWFb1dQB1Co1xdlMP9u/8wcppnAVrMZQJiG/XwshTO
JMNe0NUbx1pDIhE7FHU9A/iKxdfMaeYgFZUTlMfFk6rjrplZcVDb2IAkeaGaLgad
TnoO2xL4XNXOMzwjZVLvm0jpuD0lXJ/gSKLvq8LoDRXUiYKnreDMVV0DT29srPQI
gr4BwdtLloNBn/rxOlZyasf8NDBXyRD3UGxFghY2eBP427qut9I0QCo46WAU+5RS
063o9Ae/sqiI9LSWGvFrvfW1ox8L7HHWZUCPzt+PmAmwdBglOj96su03Z1ejuyoL
94teq39INRz76Efo2MB8i02tkd/J4+DlSEXKV89IAEQ21zXIeHJp3ww6xKmImdDt
eEDFCBD5KyeCrTqIFsJYOvezjOrsXSMnR4I3P8y8mY7TaET2Z8UmvxHmPpntTuPf
4JuAxmWVk0v6QQD+xguo9mdk6+/DF+0K0ojbrG3lb/HdueAy8IZRKBdUq46U6s2B
LtyjBunPqO+FMgQGG0gTlvzLrxreAVBtUkb6HXIz6FxtxQ4QWBIY6KMCi0QVSPDj
UN2tBLUSUOZYJtcmYgZIlzYKCLaA1Pfq/BpWJ/ubJCeJXMkzmSnAxrXXsEDnMNZ9
huz3IdIb2dIuhLg8AgZUgndtfmVrwcQdSCvOc/FSvnZFF8DrlDzW0Kb7ZHc3AYV7
8V/fvHFE7OntwyGwzhcqg0wLuYGtr4BCRI2MX1x70LKLS8yICeLHsYFcrxkTSAzM
sRLQ2llEllR/WYN/8tvFdnz0hZHRWKN0MUvvi2QKvqOwcKzaCNp2gaDGYHNavImr
VwYC/4gQP7/W3UHNw68LclApbXIpLYpk/PqaaXVVv8kPBFxaAN0pLRdWSfbvAQVj
iPjyTJsFm9Ro9L5c3YU9txhmg4aVGZuMe+DnPMcd1Rq1jd+Lz2rFD/bSqNmmXsgX
zh3bFEKnsjNtwSgglZ1wsxnM6x5v8QwtrXVyO6LYFmBsGas6KeNsz7x2Qrt2h/X4
JjHwgmzb9C8pzB8Rv86bUtYbTyABYdfuC8KJIludhFA9ygqlCz+wfRS8eJQX6iKP
/OJzo/NaLJUXYlBj/Gzq0J+CjZ1iDe4hmktYC1khgFKdfDv/Es8dNXXO1nggRMUi
lroGRUkdXBNulUjNF0sXytP2xYdMcJXJaXbGfp+2LfMDYjs6ZhRJt/dT6f7JpCre
eKU5L1Dm1I3LAoul4EXA60i9YBnQNXuQRKWBnajLN7CaP2wayPfFdkPYQvUmBCAE
HEaytLDw6OVeirTG1qYKVYuaXGrCz1hNLDezAJ0766XDSigU97/8Znlr8rZbNDFY
EYVdLkMB4MtwlqTrNSsBR/LGyHXvmTch9uIgDagteLj7Xyp1N3JfYz5s5U8g2NxS
XAyQSGnHc/Ec6a2wKmm5beuHyjXNO3oZDHox5Ae9PAflKoJYygbTWT6uKVQQZiiH
93L1RTNFvhU4G+GlMc/jGIEDRv6MtRbRJ1ePsn5y/0ovkIPr4ClvukLL6bYFHW+9
2Riml+jEy0rPs6VPwp0y1nyb71VgpoONSry1ybcaNACNDXJtgldCMKL5kosXwICU
zrUYjL9I2tZQqC9ETe095StQ9DCIWDB9BW3/nF3sW4jwaAbCQ8ULayaUGOTqRIWB
lphTqpyEZL58PN6SedKr/JLtKH/1+t5QluRAiet+xC7IZCo/asB9pOOVh3VT8ayl
s1NpLs22jir+BoaYn1P6Nqf9EEivzWYcQBu9Af4DKzOT80LASBHZ9NaLgJEE3cFa
pnpxs3tThuMqcPPB7JkZ2DtAaYCV0kl0ZYfnhgbNKjKvQvzmGjlA91typSPWtP4J
8hsgVvgEqZrzLTIiFCKfzHYFNhGujJhJuVfRbFQxgBRIonZbCst5efTTkbYB4Dp6
OAucvCyJ8Y2XArWmuS6eYPvG+7fglAD7VrVKp35dVe/ZlpOPe5f/seskwEKW40mr
POqtpJ39grc3tVCVSafkYG1JIvgcg/lUPmRopp5z9WKsr2TERoyWxQ6vYWQkA92O
GjYsq3MJtwR1/oMswmWOxzYtDIhjRM/0/l66BOSGB60zgBiwtDaoDVrd83ktHPhJ
LAffkULWgoKNERfSuJIEy0RGgC5Op6znw6ADjp26B9WI4d/f93URrcG+YKMlNLQU
L1kdj4fA8YMI/USm2AhabXK7KJ2CvaEOQqTkDwlyRC7q5YCRDMdIVr7g0HZSMOCS
TZX8Fdgj+8mkQOq+gWulPG13B7n+U5z0xvirde9QI2LKmUI4StoxI0C8dXW8BTOd
+5GwNwE4pNTWocvlJmcRSaEjgGZIWDQsmsPL5Q55uBdDCRvE8FXCFBeH0pnZBNdn
JmdaJAKDLGEh50VrMFb36d6eIcXrQ9J+3lw/LvZCAlr5ca08rwk2j7SAxD81Tw9r
cKbEl3ygrLVXZF8Zt88hGlC6eRYNdXEfL1pfwFfQ5sE8tyMVun8Y2oY399SwrnSp
vO9+R1SCcDg7+T0CV1HmSLUvQYqoV/3a0lIbRiVu6qJ6Bg2Re74+CvDh70pAMvra
iUy9nDgCv72Q2fe4vHmfLDFgwj6aH/b88jVDg+JijiVhL2G1x0I3mtQiZheyegnu
dzdVJG9PX9IUYbm04hsZ3Hrlmv37rjJEUiQel96OXe3ndp2SA1G1fS8ONd7mhY+B
lqwdw6fOCw5yB7+g7aJX3VEDD5x8yG7ej0ooXULvD3ha9f8MS/1d+dMbqerhkIAP
PIrZryxN7IHakf1t14/LPTMOZjTFnmkL8QgP3H/Kvqx2368ufHJdgVhA4ohBHWLJ
35wyibtArP1xutalNEzugrArO5w4ljiqKmaflMx/1THw4oR9EQDCz5BiL8dQRud5
a3oVw6jSu/iJlvx6eKvOh9sNaIX7UmW+FMlLJQg6ELALVqVfGmwVbZEjWuKc5mel
Ne4O8WSvv2qYHRnaAm96ca1owWzpyqD0cV6DPZKuksaH6rZdHbrS4gcccgw4+HzJ
3/kJR1o9ldnn6n2vFI7O3z+cDp0KUB0XtLQEP8nqhNNzouOinrE3y4Suy9hLQh0x
NJhmOZDYvMQNRmU15Z3F8zal2TR1n+EVqPUkgxC8KsFtKULmdkIyKZ29x4Dxm4S0
3et//Sc25VOOpLFrLYYwOu3oouobBlj7f7J3Tp0xqttccip5wa3sg/qQSmx4ix/n
/7otFDFKcqaB3GsvI6KV0MaboSDUFXwFrLmaTpWcSHZdV7H/9c7aZDdsx71xMIr1
/bbN0oRz4MTAHLxp9xh+4MEPhtdclaHLO29iSZQbolX9OwS0L2bweTqxwA+KKJKD
gigwIgasBZKP6wU8Bre437wAOp+sES1a7ga2bJ60uOZmVXGajMbeRnrCIN8fKwAW
kovj4AUhgy8h+NtkrIzsJGDDv8XrHsMtUYwsINctrljOWw769Wc0t56/x3KSqWIJ
cAgWvpR9MNwr8skXqOD7Ohml+aRQSFMruMpcf2KVNnBBWCiOu6AFD5s4ZX/jEf2g
AGsVOTj9IzxzsvPFN6ko8OUdC2TFWUOlf5Lx9IlH/MHCEYncWT2Lm4wMSpAQ5wip
/OHX2TCEMMIZeLvfw1a3EIPDIjny/MHv3hkVpHsAov1K0T2BeVmxuUUZkgorMabD
2KXNicorkHv1pmJCM0HdNsYvHHCwiWYCyeST3ExZFH5sPMVCJ9kOZn5b8/FXqyyc
8hYHzhDrU+7Lxe2ojc+m/brfNJk7jjSWK2j4SVyTkMNj0x6oTMu/wUlaoqYU50pc
+ARuwbwlLWgj+SUmdsSl1CYd+EsjysqAX0hfr6TZn/V9/gG0jUpgvZctZnMC6zMb
/qXqZMqFC1fOLwI7ZyGIa0BkMWZ4lVav69FL+tfWscEYB+XUczyTs0o0Lb0Vcy6d
lwInnu6M2GlDxYqAV0C5eZ4VIMiIN0uOWP0lX2w9ehbrCm6zAw2VLTZIZB2YF++B
opqvLFFXy2LECtL634HiLJuHbsquGG3ZK51BL/qCPrfLv0MWoj6cx2PcuMZdS565
tHXn3KRPqcJLWOaUnR2Q5BjIUGL7Wc/LwvIwiKsio5GnXvh1p6OmBtLuwnIid+X0
vhgHq+1rWLRBcIubQ/Ac793HpTsxj3S4pXemwaBuoysv+ESnsgrvBGWPe3e/YZ1O
QE/IJ9vKJpD5REaU9vnUn0X9od2wAkpJ7zs024lqdNTOPLENaN43bMnSNervbDaR
/y07xuuB09u25sSflPw+1Wjx9YhAIKq6ap851AWLk6kon6TBjRwd2WkEFotkUIpB
vCCzZMtiKo5I1V3UKy10B8dk3yAz1LSytXtc326vMojE/+SkzR/3cLw1yngNGY7s
C/+y1qAyR58UJ5LO3NywPe3M/YVDJX4wnzThIZhfAVCoxnyXG02HssUqsDvpsaFS
6EJyrGOyFB1LWgLsbkNep0p9Py8o245ckM0i86yHlohlRwlEa8sDkjw/qiP2qWzy
BaqHQXcEyKI+nile27jH4kctc8xVa8i/yGbPSolgK3Kbm8gSUXKa65WkuxxaVpvk
uGtHVWfkTfEnryIoC/6xhvLXCItdWHG93iIDDvdVXvUyrExnMGK/+zvuTdQUhjWZ
9+CoEfPPQUV4eiRWRpB7QjHgiGjkW9xdyFNlG2Smhm2NbBBk4VR3ppY0NWTyJvA0
h60vG2BNgQ1IefV05v7uahKTsyLjADN9/LnCsfQGvpZjdKGGCjvrxyS1Ls1QA5PO
XDv/tTSaRRjGeBzYsffD9bVIF67+BCU0IsDqyWZnkgZeJeR+SIsg3e1uOnlM5nbd
wPz/W6UxO8Utm8kxmc00XrkOeIiUht7uw31OaxC4g/08XOz/u6rGGy6ZRwrOmXr7
c8amxxKZoyobnB/84gnE3lVMADIriEo5SSg1ajlE6m7rL0xLRTke1IJEiqBlWCc4
9itr4xp70zOmS9MAWv7T7NnMv8U65BGNWm4ZH6igWlXeA4+h4x04/oqChKvIJ7qN
A1x2dtI0fiUrY7cPk15ajYMsAy0nkcFdos/YxxuzXmSo2FAQS/nVxaCT+2bMTDvZ
8HifU7p+Y6jv5m7PtjebFOMRmj42ct3IyT8h4xO84Kqo5GzZHgMS72Iq2l1TRALh
L0SUuftsoRL8nN4M/fYTZpwIZeoWQqE8GF+A3OFZho5GeDgIiD+M5lAE92KFBLWO
+IL24eWrCFXsH4ZILRSOXTxjCFpLndFw/vWlHigatf+xeyN3ccAGRln6ayadBkuY
+TUe3s+q4OXP1pTYLfKX5XeyWPEW6I0BLrA3gt32sgjrRMWT91kHgmv/42++pgJr
LhxUM0JLfBIFmUeDmMJGVHTbN3a2A7zmjhCE//veI8OVz8kmk/MITd//ACFPFXAH
a+39JxuxGDvWCOtkpW4LPZHu6icquESFr/qjPOiNu9Z1y69LlcO1aDpkMwUoQ/3j
XIbB0O1bvdtog8mzsaR21JTEFA/gCuOhoOwe+Q8dPxF1UokW0LbsnAdUul0nnbi0
5fNmwtlQ3SWxJDMtIxmkoGlmQ0GLrOVFo/3sExNzmTc+ilG/TKnxu6nwP7EoAUNu
5xP6yD3WaitpMLcbS5N/pFZ2LPY4ceO2GC4rSyTOZAhKJCCWQZmzipOOe+fIQ6mV
k8u183H89Mx9tkQE2ZJo+tfh086fntckVZnJrIrdnvUIi/aQSW/135/lkAYbSFXf
7mDstLF61rDhaEYnhmBkls42GvWHiueE4EH3X/BzFlfujjNIoiQJAFY+FXU/eqaD
tGcxou7tjzq3g0CghIYc9NQPZNc5+7LecX9Pv+XDz1JpXVVGpbO3tlB2mTb3ulI7
M1eA4CXUUOln1qMcIg75+M+i5NntzqsCNcNmx1uI/BDd/eXWoPOzfFi5NmO9wtv1
H8XlKhImb4147tOWDVFCE5vSAtj7cVFBS4bCHzsCEvFr0rZZhux0wqcg0jz0mNv3
pGMEea1iscJ3SXh4xY+RbINUg5GWQ28jpE0+29Q/nNEVxSXmI9vMQ9JC/lFcaYiu
clQiw/8P6lKB00YuhBd8fVD0B+Y3OR9IC56L1JUYD3o/Io1GLMzt9C/KUT8lr/+x
7GXDMnDcY0Pyv4dtU/oVF1dTMelPpcqzr5n5YoCkfR2ctk/wYuH4bpInygfRT4Fo
O97nfKEZzAdbwYgyFkn565WPqG9HPCw7+HoRHm807Z6ERmdNJJqUxQ7YiYsR29Ft
BAiJqlP1AagUyGITiX7WLbBYxSam51jEPvAMERx/XybhxO6zDTfmssTgLFT79wmm
BRHSwI0UkShc++XeOW9CjE7uYBf5gA4tLqupYm8xCjHXqfulP6h+ZJtyB+jhynmM
r+liOdfEFqQJNOP+19+SSd3k0OsNFKgY5x7TAyoggHO6Xka90t0sbjG/7Y5yL84A
/07/MV5Z1JCvpwhcZs9qyC2nSRcAOG91mAkYDvYg4gb9uAD24bROO3nQP/mwQUUE
xIBPIcSSU3O+UN4Ii46oJqlPnrDNoRJThkCRu42Rtmx/8CVHC7ZnQbXltlpWnKwg
N4St/b1SoFQm+0qFGM+/VQimNOueG7IEBVAwE1u3kVtAJGxoxUkrPc0uHfZfZ5rJ
vnI2tAGV4xW3cnnkBrMIeMzLnbxYMsdSBY1UKVG+0kJuG6b9y5xwKnf5fzqqgOLN
5I8cdUW9uibMWMSH1UR7m6zeiwOh2KnIVZsTxhDXGQvm06NlR3LaW21JJknbdAIM
KiaMNRG08Hp0QUUJMFBlBRSUkSCRjIB8HLQhcF9LDAuzy/fOft9WPRPsQx8nceik
1W0qb3/HKaAKgHZ3fzhRq8xY2EVwJJrjIC5pykjoc+Kdnvbg2ojN6em4vpbkDSJG
XyWtQr3z1PTzpm0eLC6eDxR/OhwJ1W/cSEf7+KbqkNcH2NneZPwg98maBori+Qvf
o+olaKhx2sl72rU595M4s2wKdsOzKsZjBfE/fYf6AFCdZBrFl+q/L0MI0YkXjRUu
SeHfSyLJIOXS1lRZTHXvvD+CEQfDJuJ6fuR/RkB+pO+PZ/M2RWjytkSlac8cImei
KQkAt6NqIM9MZ+rXLLsRjg5Z+3yMsItH7ngmyE6lzJ7n4x8zImh19VSySx539q+u
IK3OahRtmUrQaLvYf6JR7hMjZ/58Ow35O0E0lBFbrQhEorjLudOenEMfFRT3+gHS
I+N9QnSuIjsXiFejj2QH/1nb/l8KmLr1C70ZsE2gjGl+8rj00k+B83biCD1+J2tC
R+lUtz3XLDybQPMGZKkt0b/lomGMtIqh4fvHfpgv0GhOj+zMmCk1YwpIF4YUt4B9
eDgZxxU517Fb8AaKxkrwkwzkhKN7jmT3/7JKyAgvOGIPEwJ1eEuWAE3jyHgovxsM
7WlGdgWTNcZgZ3lfO9jLaShiHXd06b7VfGxqiBc9gWXCGTJVxdvMDnHwn9y2bNXB
ZjoXw+i/aqLnN7OjXyL1ltqz3t6z5imp32yABjbt4P/5xcrWcukjG3/7MQ5U8S3y
ZivTetNMpS4Q2BWpAor3pR+iAyco2si1c1Y8x2ikn2uHxgh2tilXxltXq4vKYItE
0XC3qN/dQXUmvD7ZzVOhz2HWAvPF2wPASz2Ms77NodDfmnCCA5gz+40rvf2Ei3/V
Snkr9yTSoMr0s3S4M6G3PdpDT6K1KCeIV2wqFoQ+pKiqxYCua3c2VvAAIUKCVceW
DFAsqEg43siVNUcGb1vxhjCN1Q2ByLmyiDy7avrV2XfEIPdiqc8dKq1zVskg8wQ8
wzKG9aDyO+HyCKbCKRMC35wxLFj1zHVEjQEis76ul8b1GtD55Hijil0B9KiM4yoF
xYoheyBj7dwGLsdr5bzpLMStbqFZW8Fh3ea9F/JQpoa8QV1jOW/tZ1hO7/RVF1iI
5aoMBH8dGtX2LDXJq7VJKvDcHudao9OMF7422SYYDczAhJDHXaHvt8aTR3Z8aE9M
UDK334yKdCf9oBM+PHoJC2xDfx4PuSTcWZgw0rDGWlWgiUD4RaLb3+mmGw/nmN28
+dDVamI4taXzgIv09FkJTuW09/zrCICYpzn6HmxYEhw8Ze8ma4kfAlrBzqD1JMXv
O4ixvML4JG8Fa/gIgDGWT4gjOGX0AeRg6K8XHEbNAegILWq8GltyKrmTQtxUspS4
0VE3eqii73EmMwspABB6Nmq83DRBLHDVNN8FFfQwrE8vm87MDmbi7IsiIRmlDnxa
y+h1VnYM+lWcj0itGe1gHTunF5bwGsx/F+pUuNhBGa476HTNy+AI6NSOXRvRppZI
+NP+9E0u7uVVe6pecMORJOA2OWhwi0IOUBfGgaGK+GLh1ptfm5NyrkWz/J3oF4Ms
gGHnaslxOVxlpx5Zjy7iqPunNhxhbRwgtPZYJBfmnEWYkJyD8EE+2rFfsyF+S0TQ
5VaktNZtKYfupLLWzk3P+DVSX27mCTycnj2A58ZNPzkt7pFMbXLeO2lNqewG8Lia
zzMggs41ZCVM6/KmN6WWFG/1iEYeV8nJpZHvQVa9Tn6rpboV+CwFiZOp0yuFsyHK
XEiwHtBtNjaHWLtySms8QcPOGTz7dC/Eon7RpCAFbOXKXZfGLmOdvEEIpigGyMbf
dIkWcdIeFIJsEaTwDPH26cvciMdeJkNjRp14yBIuJizlds8oElDeDL9QT8HS6eqs
NHvpRBdTh1qT42KjUlg1tLwQ2ZE5mbeB657rTywrlKRF67Pd8giEED1LdSnjwGcL
ag8lxR2a3+n6lJV8notRxn0JcltFHhRqnG95FIXh0ExXM1Stf6AH9iT3ZqnF3dCj
BqdjJFpG/anRO8Uqh+GljBpo0FLVIo9KwBd31+TFTnG1LdxN0osK8m1/CWCkPSVr
ezsJ6sJfxL42r8/ZlcEZZlzYtc3l7figOF4Nrx1XJe7/SfH+sRtLwR+xHesLqgtd
sHDnIsfciANnSbCXjTbmzC3HVkXBOK5iXC+oi9Zy4yRRVUtvpL2zYhaUxjW9Js6T
GSmegYl52A8TYVOuwgtMxPDvLaugVQc4qfjxhj7eEMikvZbDMePEkW5gLVNvjQWY
oXSGdrkVNL3mgUG+yuBwAe9mY25SkGL+nE6qnUMHBuhjY6OAa+8cPdWaggBbNs6w
mVwVxziB5ePZI644rmHRqNA5AGI70gkbZDe5L3mleOYIiipHaoi7i6e4qRGyymbu
8T8TQcOKVkMFdsJ4bux3/pvxMJgZ4LyXESmALFxG5uheKR1FB5dvv022dGgOob7E
q1ds8RUQX61Zc4iMIZBSZb+osVy0LEjbeX8hdtzmxR6HtThjwtgtu0JnBLZ5DyqU
0hzWyhhQXHR7nqCqZguSc9GrgP/1AZmY6PCqI58Toyx84AV4GNWFOeHqCsqyFUSV
o0E9h6+SW1BIY7om3ziLBZD7IsiZ+5yzedzjBLgz+PnKJgxyRmxEI2ITD7R5ZCs8
5MCEzQxjq42GtI/UP929y/L4KAKv53Tk7QnRkPqAlrlKnxyQF1p1kyAZAfnlxWBx
no5o33pCIdZD8Kss2lsAGDxSVw97B7Q13Etdfr7ac8WjxBNOLfEvBbjBUvYazxrW
E7bsouTIZRtVaHCjUgNMzjHzfahxxAVM14JaY2ibgIBS07jqMaep4gUsO60MddOB
DU7KufAda2Nm0CiYre3Tdt7WPvAcZtwb39Kye9R7TT2j4pSfqyvZJLJP9Ad+d3ts
KTWUsZPcTeER9ClhUewYU+uKzjRT+MBjjgjXbDlgE2cyRhYGGjIEWxuBrqAwkhuI
+EabJb9LKA2U/8J0s36LNzvB7m410RyPhAWiRHLnVrKeqCRn97OCRopG3RQWtaIs
8Z3+jhxrwq9s+dPSMnXwub9+Cb+HWFuW1WKEShBpxVuN7HadYNDpbDGydIKGDVyk
SBu7yuq+S/w45iD4BmKnSSR70wVjWsiUs9BjiMbtoGBafc/gNaLd+wOvIodXNcEU
tkD9RFcRPYpuiXghrnbTKZPSb1dStLxpXCKjvcs6orezXhtpV2mp2PJeyA2/Otlo
jwWM+kEr5bI0zhxGt1JvYvG7Q90ZE1GcLA61X0Q4+LESRhyjyb9HjOokG9u6IcY2
IFA77mk1tCzTaJFlhpT2MztIYNc8LaIbkRktk41sPtZDu7gcdq536+BFQMN86ow4
foArCJGHNmh1Yqut/GuBdMZAMNU6Bsa0J6Ni3/h8ovxs4mZxgBPaHtt2kqaN3R8g
Gp+DpcAf6sWQOkQxE6dwC4ntIifLlo+gsgkIs7oQnlU+/Mr81bCcB2G6NjzMnUAK
liLR412QJJZPnoQjlU6f5AMFfAr8enqeLZl/VriKChztQyssPYCF8IckI2ncoD3y
cLjSXkBcMS/x8bH+bQHk3cz89RDWQI38SrtQovzY1HSW3m4snjQk7xmG/MWWuw+I
GTKk3RYZ8Yi6UFOmt44DEooWBYCxmDBGudK0Q+9ShKwLXKWsvu8DjmCdVmln9m7s
L1HWYXPoIQWo8SjIzYeY3JG2iSjF+EpyCH+5yeVSu0tYN1COGio1JfXs/hchNzYS
H455fqDzTbMRwhS3vd0oda3hXUL1hXhJ6mXZV9fxjIZRfHZknVw+lWcaWyECVB2+
r3ZkMdtqG9RASehuWFcIWN/eqJSl+q0E+TkI/D64vSbMAHA2hPz98O0OrpAvCIwj
clYbsntm06yKbwtULOIhvRK8dJ6Dg650H9OnkS3EIiXGDAcwZZfeLF0Aj5PYlFWn
Ez+AaQsSfDwPMmDZfQ4l2r1RVusMHyTV+BEqH2HdaaM8fRAKQ3cTVakSgSQcIjHI
qs31S+m0g4gvjRwiBHdDrFhNyWY+FrH1qpxWeHioycSyakPot3JYXrCgcAwIx7Sh
gMi4BKG8A/QKl0QzweWjMTNG6cwhVzFiK4fuCHobvpZADpE5rbXIqe/xPDxBuWXP
iNdg5ru2poUP9jS7Bz6P31c+/3ZaYS8G5h2FnajYFhpRSVoZo3Vy7fdbmJWua9oy
yHkiQmgZYNDCe6u7+WGMH5XdgoQ7m8x53QbxGKCMfEjhqc6+YCuUct3Jn8MtZEIf
jaK1416yZfYtbPCTPqpmkOgSUtYNOz6uZeZneE46hXOIXi4Yffne/IqC8gLEimwq
FOBLKVsxVhzXXcIY1iNVGVQQiplcSp53aLm45gPntvPmFQRmJWCcZs+/1lG4Zvz5
/zmWpLGBNdRbnllpIUuoEMsjLuACKHxrlNaruGZSVM3qDM9ct33gn4dmuNxDeCTf
xDdbLsdCwIQ1Ojmqo65B6S/fOlQe7zfvu5VMgsLsfj1pAapclLnezKs+vWrh4snZ
ywg5G9EDunjD6DaYzJBWDMwtHopcSfkSZFagJ2U/DRgX7k0KhDgIlAZdzB3OqWhK
qUg9nS8ZGDCGVutisvi5nqo6GdgwBusgaFz5v4N6pyuXpwlj43omSvpTfxnthxP7
cvGsCVTrPLe59HCL8FGmjIIs2mTB/dw7sEzw7oS/npUTJfzqdjUTTJ73KNpm/jMJ
/RNdi4iX2TxYxAESiR+H7+iLT1GscAUJ9RQRUehZzksmEXW1fiTREMRGGztld5xN
V6kLZrthxfnNaBtyDMt95rFTlbue+3qSiTqf8BYkjZ1dbRlztkBBlUuw286CNusl
L9rCf/ilNExvV13zNxn2WgpoAm+uM9HYLaM67+d0WIFxEkO700Dg29JcIxM3l5j5
rJizbX7y9IaapG7IaQ1EfFxFCPF3xkLOVdIqbW8cyCpHSUmSGwNnA9F73T+kw+HY
uEwVjNxAwMNN9mGkM36ObQjtDuRv5o8/gvjPSNIt/wrgcuI3SHsa10C2Z8rDBwcY
zPOuGv0iiHSV2vrMOQP/rYtWsQp6rfwfzoPO+KI/m8QfKWnWbLDwtCysGvEchjRm
YcGTnU0C2P+esTUSh441gWnabHrro4uBXNkAPhC9/npJF4hH7QHgPmURPlbqiAHP
G6yFyx9IGjT0LqesL1JZjOlWcu0DoWqpSj7OPcq0JNBI8ipVb7FbXZXuXR8uXY77
01oxFhqhiDRBWgYBGwYWwjFwWcSxSHzp1kdh5XYcQADTToSJ3DoWn2ZP8DzKhInt
fjuUB9dbrSw1YunV3z0PQtSH0PQFOAJ7ZfDCT4L1enQlRQSR97fOjdOyhqLqmpM+
ExqTwywqxFbSmmVdb8k33S63sHWVsZQeQ8wyWmvkDg4m9lCj/F6e9Wx3x1no0gNJ
fje56nDTFiv0+CXM+VJAS6uZfTYVL4zxn6DUmOqsunD3Hh+Eefn/dsEHbqkWWAn0
TTe4suHE3riVZ0MDymZlxaYNKTqRlIjx1NPEvU5Tnz//ImMk7Et5YLC8uZDufpX1
Cwwv1PaRh4spNIx7E6ZuT/mBWVBnZbcn+fnb/A52HMORPy+7NgcDtFovoKUbUvd5
K6ItvszAsCezommxV/D18pLfUBT5tMUwDFwDS5jZU2L2VBajai6s/LQcKIDdgQVY
oZEGodygHzUz65HEY0z6r0zLGw7ICNRCThk50lc5+T+agkLg2Ut4ltN7G+FpQNg+
/uhG2dRo9N/xPD9oMcGAb18LDMpRyIGSMEI/A8e/lvNRrLxslkTogLqbKh8pGBOq
iB72h7AMOXlVdwTCYctXuEW3e2MP06Pq94gZC3XH1Pxyzn/7rDB3Y9X8y5NOFX4i
6SbNLz/uUMpQTgTEXJ+HI5OCUP6vYNRrUikbYYEqdE6N7I/Vlc3ku9ujGGyC2VM9
oJqkld18pJWv19+puz/9EnqxWkX+ttWyVskFtACu2BCdTP3s1W6vgwZVNQbG1oRm
SKpWITe8jB2H6ZxucXwFqOTppEYohwnwXB4LN12PfW24Z6wFNv2t3/LxNov+WrIN
D9lTRIMc031ItsRAm5m05o0I8C1ba0+3lYir1lrW/LU/pY3TMefCIsXYL84cBCIb
R/TBnZSsdUTrRktBDX+PDAPmPWVjSvvfdwZnUP+t59CQtC+0gZkrGsSHJ30y4fm3
iFjCm0jZM5dfztxKRCBs9rQqeFZqc6CLxow8oJLbnvxRec4KLi+stvcV99JQ3095
eXR2meHICn7LV8HVcClxU6fLAGUs1OjPvmyp0qszI4BS1eSqk5rjN41onpRkpD+z
JXj7qCTUSF+5Eu0FxMXbBPjQp/dYcM+cICTE6RVuPbxwv1FEJmYTI+xV0TDtG7ka
isZDkDWZC7rQB7g8Trb3ygCtRSYsmTwQ7BawG7+LTDAT50lVNa4MuhH7t/RlRLaK
/QjnjKfmukkOJDq20sm3cSxZudOJn9Y9mgAcwtPKebl1t4ZRxJtc3dMxG/smUceJ
C6lytbCz1OmwPANfsONc3CkJM067ScidOSUGERuXl/UbAuRoL+N40xKYAMiYMrLl
e5AqhN7ANiI6UZ6MnGRaO/Pmf92TFgTAri8KFCr/JyTBRwEwutUitKk3aJvlfeBO
/XiZ73fmRo0Ty4cHtoqGebNw7mnqILOVTju3Ds+WxSWHLZh9gsT7KnqRNgYJceYe
040hj0oi76k72IKQv3+tTCFOfDDg3k9r3YtB2yqXflbV68OmktKLdGQP96LGsmLK
GmIKUTtiasZ5aNQ5nRpFc3fRMkRxhGQV1MUvkBkFbRBHfF3q/o8UbMB9SqA6Q/cV
ktQTLpElt8sDQCCGwONK1hP0x+3LtBQpaFnB8piVcZAuQOZNzaADQDuAycpacr8K
KjpJj0vSNgqucHBZaq7psSFTGYeV2FhxlvP5sFAH6NF7K3005qbvE6m75kDxXh8y
AO8bX3RaIwPh44PUGi4QVwtUlsvEfJnMAP84JpkXuVvQY6G0cFXvdHLtS1CuTU23
cv96I4S8Lv4OTVwQiN1CH8ZmXOVrAczy5b7yTpNTOj1EkSTytLl8iMrczQ9DEc8V
6q9C9Wb5ndK5gilCCwUtW5ZcPOvFMMi2d7EH6sFEieDmPGf3Up8erV1ACXXrxA+4
IsXB5jeJ48UW8KZVtlCTqvWoshWWnknsGa7T1xlwcBqS50Xgv9VgaE0JcHp8lIb0
SfkbOo0d8ZnmR05OzWq7GoflXAAVvttmTLtSF/nDJnEE/HU/c1PGH9n7FKDSwimr
oBJSnHaWD95k4azzroG7Ppc5+7lqOwdr6fWih5w1ODsUeUx0S2uk+KVJsdwRwv0r
66O4fxBPuoPIEGpMsKuA6dyQ2aEZIM0TvQTPOLCa+DmBvfQLm4vMdMfu8ukkFEYV
u4g5s8w8h6K//68Ooo4SA+uRjjtxQUMfyzmkeQabhamuEBI9BeQjuqWONtzOo8he
sChKZmvrPkNM/GWBcbDC6rZMvoz2NFCjeU1Q4++M+S1i+K4wq+aA4txgQ/ZHEDVg
8JurWtmNT1J9QQ3vVAvk4tfGmc9qzJkFecBgbsQp617eVPp2GlRYzqCXK6rK6V9m
Ss+VrAU8nPpc6RpVPQsyBeu3rFPIwWOW2FbtZ1llRFRMBN2TDuSNizAJo6xe2RDE
+RwOf5PK0R1BFCEp88EjBl4U0Cw35bIa8jj/wyRRBdPkFVzui09q7y57X687xdY/
wLAxwM6AH44OUfETARS8BOS18FWuN7qog7cyFb/dQqPLK9PCrgWf4PpgQHelAEDE
pZqtwz4OJQ1+ZtQpSdCj+L/YhPD+oMWUOHwTJuuZ3mUPW/bM/lkZAydwxURK3HRo
8KOz49rJaUivsamOssA8JIcV6K+9poSZyZunTqrE3UdK7eigxBRkD+c5ddl0/W79
UqVJgNHIGpkrnoI7LwE8Re86Bkl/WHFMDMnDOFOUfHwQIy8C7gwNVtC8iy/w0B/x
Rb2LDUPC1itBRzma8Su6IAFggl50Z2vXisPQ0F4rO56ZZ0I4jSrJKl4+xzCx/4d3
IB6XncGtBQ3fIlkh72Y46VIYgzq4BvVhvixGaL+gtGvEw7JXF/6t7wSWDLCrNFow
FO6AXHvxWfWz/GFb22UH+6/Z59+98TUxDP7Yb6WpFk4WEzkytZEdJr7FdDw/IFNs
OvfzFpb3dKZS7QUzU8h6oWnVLCDVB1XJSZohKOy5NlMS5VCvOlfmzaOT9owVxIPF
J1Z2nUgV3pzL7uvnqRLz2PzaIdrttWy2O5Sk5QVS9kepQkoPNeZblhR0lqRLfitU
xqvGvXnKwnvk5f6DwHALB0MnVX9dPxxnX/PPpGqZMd09tvZTtpZ7CTUr7pqIfgY+
NjgkhVWO3VysQ9XbqE4FBhfE6hjnQRhRI47ExiR6TXp+VWBjYVVkD4upjI2kzCDd
+B/iJl1ZBwJ68ZlLTwL5EIWJnSGmwSwP+j0JBmreUa9FsvWR6V+/godZfMHlgjlf
dqgPGLBeJSQ8T1lRkMN9Xege4LGosrRtZ0LOPlzSmvbphd7X9oCPiVwo1vuv6L8a
UuqegTBOGl1omKrSPkaMf0fWCXPkYhSJpC+ttPB4qfveK2nkMECudHxS31xMD8Z3
vy4NQo5casmG9wni2jNFU0XQhQ85CTcE3gsZr1qDLoO5cgwbXp/DIwOoWbaSDmhX
I+/Wfnoe/8dFiU+2xGWD8P+XDtJOVKfAf4QTYwXvp1k1Z4bx+nuTPkMFtB2b35bB
Qc121wwhJt2+bstJI4zjw0U9ahxNBxf29bIQ8j2p4LbIlZx89HZ2pG8Nvyhrb43B
Shd/l2kPdPYVdqEyWoOLClo6wm+qskEtIYbsodTIfSjVC6jncJlKStLsYd+BRft7
9vjovy22Yh5ehTvC0qtNj+yjgvUuuFnttqfsy2f6agTF7KmHkmMYmYIj2Lvp3yAt
nuO/aOn8Xj+aKunSu+u3vWjQGc/kNJOMcZ7TrUdECV77P2fbbAso9LMqyX0MUUno
PZaZedJLpf9HC6gZM+n6Fi50udT7gskR26BLPljP9hLscoZ9oh3sokDiuMmbfrQB
M95lJaxWHtU9jgCTNajy2yIk2R0eoNUfeJ4W2ztmv8GipdT7mJyhRgy4LLrbcwYq
kKmKd5RuEkUUdhaH6XU7o62049bgGQnPaz2BNN9IyYKCEVVHIRXKz6QCLA8cu1WC
XKLrnZgFYKHYJd6742dxRYoPdyTi1lFgMmjtcuGQPAIobsTM+rwRkj8959UKmAeI
Ueew9uG1w5fmfp2szEFOoznYjEQxm9GcYTKSg884MxxTXnd2/Pa8Cuu0Rsz75DDD
Ov2Omb/19c02kWjSkcHGuUlVlNGb8W1XBK2LFueyDkiTiLtK7ontSDRjwm8fNyIL
gVtN90K1TBzCo43A6u+CwVMInGlXGNxwLlgKt6l7lG5VlwBr2eWwjd92zcWYgsCy
huJOuNedS6px6KmpsWV27B4x/JzYAsREnbXDGtYqUoGFcro8GAo4soPB70m3gD0S
pLfLoS+DT5+Jnp1ha2kTJZqMgvynRYRMVDQD5Vb1GXEkLtCxnie3Ohf12nzwjMmv
WrTcnBV3I+whc2JqMY+LNP71M1woleCRWUQ7bwJVG/wPK3dP31I9qPY3VJhu9pO9
Xxoj3vhp5VrLofFQlxKZgOTZvjShYwPXbXz8oKYTmDlBJifgb52TFlH0oz9fKovU
ZwDRo7lYOXXGkC7EqVe1Q4k/03AXVQq4B4PTSDKotU7/ClqJ2Ju5ggs0jWDVxTS1
+dGhGIAmZm80kjdw5o8/a/5y18+PL9OGihZZnNpazeuHWs0cEg06NTBnE8s/JgP7
8SON2MknBMvyNVTMkCqzramQtKObViWZUVIXk6e9GPFh7JlVAfNDCg/J5NFcu0IR
GvOtwTTnlNiacFFpczTrCPYySDWW/NdofL7fW/jArWJ/Vy2B0ql91ZxGQuy5biyl
8e7tqftFH52CWjxVBmTwlsIuB6ga3ejSLLbhxfX+DMhiBp9pKeICQInWqMWv1XEH
yNCVzKEfrU7zrIwwn/yHa+KVGK6REFuti9jlgi2EFc/mRQYRaRzvt+r6L67aS1Dp
m8rtJ83FPg/qmiQlmIUp4SSL6rKNt5gbU5x7jLjibhaYGNW3JzkgOwgaY4Gl62xw
O7t5bHbNP83zQnExd58jtYZS35Z681fMPgYy3dsv/pEgc0y5p2vhGmmb5q71eSlf
T6UdwY/nMs6dr1+4YQuhYBHpDzlGDbKy0asgHWHuDwBboUaNuz1vtDp7G2JL1fpf
Sl7OREUbEzh2uQYrW5z/e1XQg2YZX88cn8XmLWgITqp3nP47rCwXvDchPIFmBEhH
ErIX8fn77S3WOpfZgT8nhMUNzE/mdlm7EbjzSZ7wY/0CEa5M71aUqYDNN2bT4bTg
wf+w0YMH7qUwUEZdtntnmK6MjsctDVppXfHTQvv8cnAD1d61dr/RL6X1X7w+0cHN
24+zuPMaBzJ5vW4CFY1NS6rU1F5i01W+Zy//Or3bI1bE1VTvp9/wSsJFy7JiYA/f
+xjOHPyU03pmY/RoKDYIRwXDivdjh8iy7bVyFcTFzzvmWk8kTphiEQ9Tt2RP6rs4
VimVAhzvl/EkmboY6zwPjLNtqSE3/X7G1hjAQORJ4mFjnOjTeSvz1FnHct8qfoHI
IHGdUv8v3GgOES8LRaRYlAWVjFm1Sy+dYWTQ92CiukW2ZBRh/FSwcl2ljL6m0qpW
8RtYg23tX1oW+FdJbz2anATaSG3owM/7m8bxxKFese6Oc+k+7Peucu9lf/fG244H
5f68P6gs5DTnPt3uq9cMpIda/zPEABXUEJQVffEcYnVPoqA1jUq33keP5jNQuW5C
KJRcaFJsj/OyMZFC9Ulh1t/wa83GAnE8qMqDmckbafdvOf0NnUb0nafJG/Md5GoB
UgivVuyu0QsEl9eC1OBruodIWIOX2nA14cWi4DD0wCp9XvuCrCD6W5UFP1M36sOK
vYUpcGvUeJ6HwzQTGE/BdJoEnudp9aImQc0rLsx6qBjpTXIhO5pGBxe8/LxgZUBK
57KyAcPrutZIHRuPjhC5qhYMvQeRII1V1O+N4vt+rZL6lUdeXmtyAkzHY6zTUZKc
C+aA2IetQ8txCBT7Z9dTms/DKt0B2v4rk0o6Fmc3j6lkX2Ocg8xNcYGBTKndqEQ1
PsPaATrfPB+Qp/yG4l46oOtEVFjP1ayP5aO7IpOCHy6HBNHp1porR9yjoWVP0x0q
nAcodEC5OD/ZGdb+mGLnMLtyFdcoxRPvYY1iFm6+yvIE8s2iDVhX3inOsbOqoTQp
bRLIybqUXymacQDTdZe6rsLMy9Mwl171U0cLOQBGOyDbaz/vJkE5CH2rOfR0LxLT
VnManEah9NhBx3pYcIdeKRYn9+Q0dYrJ3WpQwMsWlTPZYJFcz5hYhS6SFuGsiWKb
FTW04ZJYJbH3hC11gs9pGZEUZ38Fa3+RgKqJcFJwFv4oLG6jm8EKP4mxwD6aSXa4
n2hWu/r8/hRWS4QuWMgpJIoezsQd02/W/Jd30sJ4uu8H+5/g7z0omNZhFcNSqL/7
FPhI72AzDAww3/Nn08ooDNTGQfHs8ac0QvnOeoDtFBT8duD+rM13jb8oXuSh719l
u/UphmZlR3vnnWbQWRlbFcozdMrnShNWQOa+u1OpFlVy32W3LZZhZr8NErY2E2mg
XBYkSgCbc94YUO6/BnLyKw5ycQnwPpzmLIhcrJdfZauGr3uDMHxjtQHbShKtAL0D
i2BaX2zvyVC6L/7ucBYnBTQM/5d375k9m7hEBp9p1skrRTaE54Ibf9HUrBBHsF3C
sI4mcJbCgzMq+kGO0qjEObBqG7AS+BORKKhhMnyAWnRa2s4HffVwTSvhrGuGrR41
eyHwiOddtAGAZLqvFbFj0aPkJk1T9Tm1oH5UV5FNZx9Y+PVU6OzGyIMpq5LaLA9i
sPbheeAp6UacQ/sRjlD13rqtMg8nkFH1qT6yGbQtjdjoT1cMms9XvOUkW8ZqZJKP
gLbpgOwrAHvKxvJ0gTGEOILj/bdgOULEBokwSZMD0esV5m0oCpUMKQvoHMUB4rSc
cgWwYvZLK9VEdt3+NxImdPNNL+wBW3s7Hyk8HzJxuvw3F4QVOaFlBrNQLf+1qZtW
26onaYrPGVWpwLGTEKR8k4wnZkFTvTrRS4UdTa1OGP6TuU0cYWOSIluTMrfq7SM7
sDaM6HzURiZtEPio12p/eCnQB8b+oACu0GFuvfmvydFCmezZjeml8Pq0K/GdhFFA
kZzFjhrTL+AmYdrGz0QTeMlaR+waxYElYIKtP/frIGH06lDJ/+bt+vhB1WIevJEe
AKW7nRCahi3/ry/B0NpwY8h6NHLyoaVik9xKI11Z6mhJSo9cOXBTZbxF1KGrV8Ts
bq/OtHeUHMEBvqoKmJ7/TKDEXHKGs95r13ayqKdyEZbjhjDjRHoE0QAdV/+PoKvH
jCigQv7I0+FPAz2gCk8geLZ47hGtLTajXf61OKh9B6QdXq5PX4sP40T3QXMh6qi5
kgNTW2cNqB5ReWGz9i6v0H9w+h0c5iRLnXipTOaxJP3GWrWL0eRHo4+c6GsUP1Kk
XeN5dK+dF1sWGKI10uVDiZyLakJFWH+U9J82yidxU4tQjJV2NijkAidihizbIURV
QaHw4NF0/96sXrrvViuxJb1HkvpnWH3Z02y+VZ2Mm5Pfz4G0pQlSQT2SIIbvL/Sf
ZOrgIL9q4tKoTm9zGThDJJeYVl3zJLT9z9O2Fp/l3NTWSuQ3NfSlkocgrq69wiQM
lhH85WwHs/7sEyeFzRpLJskJdcI6cVEzwstK7RVGNwSCTrzQBFVkX6TSmH1gMnpw
FL+gq/aLlbRIfUnDFMUN9H8C7Tu+kZIawVB0SDTvQfW1SVT8j4+UDO88Q3AfnsWG
gKjOPgQk2/C4PR6i60effnNARjuYaCV57lFgjnK52q+lYU0OnZkqldBqnNV9tLw7
1FR8VP0tOEYLJZPQqSkqJIV3gRr+VL+exaGZuJQsJqnP7vwIJrtvgln3+6knC2II
G7O+r95bJicL7CocKjAeImpfimiWZvnk6Ywk4Hin7tkKJYtbY+SNqA8DFTl8G+OR
GHLTYfvFLiDZgM+V5b91Ocker7lHz9AXYdvZEaIg4oWPVqr8gIXpo/099UE1tgI5
mcAE+YszrMfeMW4SsTy7XGuER2UO6DAyaeeNRIAvppUbBbE0rDyvfEkSdP0mIesI
IyBffSwzeCy8Ekxf7+3XJ16srJhDiFx7MLHBlfH+5RxFZ3EpOBnsQTHebxM2Wxeq
eQa9bJAJ4KX2fXwZ+Pk2lYoFQtRh7DUae8VlTCi6AZLedH/Q8k4sATv6wg0Ou+yB
pGYaInHV3PZBeF1/0jIK1BWuKLRWquzh1ze2Fx/qpm2rQolSArQJQwxy2gITELfW
O+B05rlMuVFen3rLB7XLPMPIX7NqFLSsA6uL7VozSjDVFp9S//hvbTf3AYSEcXKW
bIoEudV/s6a7+9klqxKrO1tUwDZR3QVp8m5UNVmx39Plgt0/WYo166yCUmphEreF
U4uGOZOzsuaCkYZ9KiJaDYulYwVGHh16u7oVwP1KMGTakhjVYq6OfE9YFQPNBx45
p7iJPkw/vCFYYjfHQtAIDgm5HEjAwvgqQ8yd2EcZs2lm7f5hkCu4ObDf9iFydgKc
gOYhKIHvYnBW2GE0Qx3IPXbZ5x/sEvtrAGPYDJFnm7nnAvMbB2ek0YTOQXpGr3Fw
Cd6HOgHjh1uhkvny3ogaw+HPAyNzShKKmxL2BiOHiTqmEZKRwm6CV9AYdhq1DJu6
0KlzZELW+DhLLHt+H3maLl4JYTjsCEHbyYbCO7vygLQJfD/yBsSkfjTdFBwBHZ26
7bRIbNzwiNnZBiySwag5mH06/q+kmtqNUiHdMy17fU4yW+ys1BcRPfEdyJt330gb
zfXoUgimMOYFBENmGcJW4fIlth184Mtbz8amAOyPgkOSvIM/biftf2XgNUJtu7SL
ILMTdIdBp0VuN42LrjUBcpcwKUm5TFZLi9o3RdEWHbQJbarWi9dmllyHNlmPUtkT
lTN5nkanZwceWjVSZ7Wmv4m1s8cN7mD0rAWQ0UA8kn5Ch9znWP3MeTagdF4AAs2H
1okYIMeXxhdBIpP0jmgTxoBDUNY1UhJnQgQ5H6UGC2/5/2U72eQ4ucMlzQkUQj2M
qNHTbcBBcvgZsMFDsawcQB3xcGh8CKEfSdTPXr3DSydYVCQzS7hOdPsfeM4T6JeM
j1vSDXqi/J/PSSI4htE7YShmbD6X+61De7pGh+Ifymh+phJqspl5MMTWePkqZ+KV
K0eRcCNl3VUhqYceJzinEOoEjNVAgH4h/mgDTm4EE5VMl88I5OcT5L9Uuglo+db6
Bq9Yv8VMkzEuT1ctWWRWV+YZgPF4JzeHmw9NQjOsa++7b72FG6C/MuiDqu/sItNH
nsgEdVa5rui9g1aLKEKd0CUgMAEcT339gOBP3c+Wi0wBYlV/nsm+9M7Qap4bGlMf
B7DyYjeAnDIPQlAWLNY02mJF97yBtE5dOwpKHgLzcasKJ5GU2SCtFTgMNdChWiYv
nECv4T81I1o4E9Ni2q8siEPs2c+sT3nlzO7VSxtu9BOXmIhRM8fkfg4Nulik4Cl0
jJ6cYapRzftr7Lcn/lL0xn+qTkqd8zikrSTIT7eZqh/rTGJnCxtfp257sWteUy0I
F6WPv/MnnWQrQpTI77V4opcCVbpBbADa3j+kR3mkr3yIrMQM1FG6ghSu6Vr1qacx
uToS2qiZntvUMKEIvYmpukX3Pxp3s3S15XYCrdJWB0zM/D54kPCaf6A6MKIRpb99
vVHzJlm/9UV5jLn7ej2+uf2H2gw6Py5HoWmAHq9XjoTkvSYb5Z6G333vBwxJpY3a
VSfKuFEf3P/GlszgJCgKrS7TdyxxLcQC5cKstmSeCa1yL4S6UfRJiFOrDI1WzNLa
PIl1OIVykNmJj2Ub1ee/WAi4NWv47HezQ0TAXhiGGdH6ZLi5utu4GfVw3M3aGXq3
HRLARbdvk+DK7D+GNmbZoQkN3ncW/ECF7cDAzKQzlFkIkIoISwJ7uTGPWIbmw+RQ
KkAOH5zU/vXJ+ZuzVzQ2sfalavj0CRYhOmAjiLc7Ivu4E+CJHHVo/BTvBRStcDFw
L4s5YqKGi5D/fAumR3QFwFkmxRDAQNry0g7TOfIVSJ4DDd59FBKbVKLZeuqI4tal
4aWfi416i58aQvpebi1qsmYELggwkaQMC0k7yE8ek8hKfiWLpx/6PFYB0wG+EVTn
WDXxDf7waznkWX1/4niNc9B0ucGLI/LP9BN/zxzmCAj61c1+5q9LprRzOH0taboH
j5iGem1oXCksKUXg1Itb6AG7KdxsGy+Pkb9KAKVsHokSGMNZYMZG1999jClZEOCw
ut0fCXu+Du4yt3Uq+fMuD4/rl3H9V40FWl8XrvXQN1MvUns+s2zn4+Rh10fkr5ez
O7nlE1bEXPkfZ4PBconl/n76QdR8Nxmt93+mavV/kpKOF0iY9k6NP+VTTSREplsn
NyOwEpedWw3pqSEhFo6uzW/Ykns63+IF4jDZd7g9MkwD/86iUG4ANA2l6A/T4Ioi
AYCzfddJYwuIIynTaOAK8mEzPsuR3PEJwTnk07d+YfIHiL4u5uTXmLd2bBthRMFs
WcVPMfZcMtkNJx8N1hMJBc32scTjR2thaWriOC8k8a3o9fiV94oKvJ73LYUkN2SS
WU90aamSnd5pK3Ktc72t6P1UAIefQ0JzYVG7PuNohqvCuCZPvpI8839u/Rwx0w3V
sFXbGcDLxeQ1f4dhEPhZ5MoLaAldRRE0shzrEkuodu4/xoPm3f+qq7Nu6r2E3czx
it8RSa+XTs6vs40JriyTh0KbbmTVCnB+jVTBSgZHT1aGyO4ujjFhAwfyFZ3wfmCy
uXzaA+QjAUPUg5BSPXtdvYOsPfzd7r7vher9/ODX9xuMlbQxM/nmaVhtZHozfQQ5
zveJJYCUgvgWuDffmTGoTwaHjkRB4tueummMdYnqyA5kra41S2PYJQbGHNWBRxpJ
2FJ7I72cdvnfJLSFJ46M86fEVGXHXPsfMr7bzsY3wDRPCzpZIdu8lxgyp+liHIOm
Jt4LI/19sr/I1lMZ31Lm8KJGECvOF3W/UY9ksqs6qbdVSXNHRxiMFTEYVyCw9gB2
34f5vrDHU+ZSNr0fAiME8ynWRCNUBVbIUNlSSPTeDF5YedytqSAzbJRXS2yY53wM
hPZeOgV9Zcg/ZIUtaIZCbdgNCdgB0czH1TaGmQg3K19HVfQ3MBLN1A/sNA6dlwkB
VqA+nixOhy/aOEwV8418EUZ4CrOHGpGkNbWg9CEB0k6afR1RGYkZKxzR15uc+m4Z
Hk5h3TS9S+6ldMG4vtEgUK4Dx6GWaLIpUasX7j4KkTrS68zY+Ls9thWwKB0B6OAV
b3BNVe5gJHHGgFD7PR37m9j7DSfJGbAT5FOifzqkPOaEWFW2zBnm6kZUVU1IrzkR
/0P2XG/ol9AwOaQkkuXOzgZwpF9+Yef609FH4OJKnQhpDYP5iIAEZF582B8xn8qO
VVxIJ3IkIWgfU2NEc2J8LakdkuExKEze7Kpqgv5+asNl/GrU6Mi/TCh1XRaUQytW
T+LTSoTgWtA6hLYsp7AyXV4yq5yas88hsf+wczqU9TNjWEFTyhJjZBiEi2hrPic8
olKdthWPZqrVpuySkyilf3LKlyJscu6e4uUNdYp0287D3an6TxlG48tYxM0x6tjX
Mmmh21PLduByVWjzDYrLio5l2GY9t0GS6nbpsnsbZ90n38IbStEuB6+14KsGPMKn
sprVdrr2wYusXlELeJhl2y1iGenZdG9NSQbT54I/K6Jp7Ks9PqIza9lsBqYTIyRw
V8KFExIzPLGXMrwESnHj+zoXCHu8ZJCDivA7ix6Uxx7U7vE1P+eDkgqTwND90Pfj
w8BiAuZh5Yr4+Vj8jSLum1pCiwPEQFSWSzAU3+105RKRJTwoze2rIJpsfaRo9w47
Cqj5+X/O4hhyRiSFgt5NDgTRA4FLVGU9TjNvPrWz7sug2GY5XzHVXDOmP1MM3ZJl
4U2KMhap/QubolEn2qe4gCoeq0ZHAxzVkByPJcfnUWaSS2bneWcxqaSOX+RFMuTS
7/P02OHplKcKDUI0gk+/cCQFaCUI5h370TFo5rNgqkbHAWCt6wWfiCy1lS6pGOqf
86rB2ALOsnvKEmrmq0muTF/7RZT2HsdSn8NOwEeTZMJExpZ24JWI8hql/75VFG06
vAqGRza33zWmaIdvpq+uMmMBrRsrH/719msAaF6av+4g1qsr5AhPJJV7i3bcbD1V
O9aYNm+kTsbEpywZlE8HRkVCuexSk7xPsue37XWIGh7djZvkurMklNssAkuk+tF9
Sk9qkdqM1Z57KCDm8hMKXEfK/S7teecpAT8zIuMlHADOrWjpQXvIgGB2vYIgPlVA
ezlXqaBhnIQrNSQd5JwoQoHMCBW7NuTwHJBtdmoqy1/rg0diDfwMUiLvSe4HYTKM
6UydAbg0rmiYxaX9FZY8VygO1Kb0Nu/WK7+sm0+F7h/r94eyBfPWyXPGnRYaX1xh
bkkrOuxZcCV23Lzf5Kx8IgVw7CrZGzAXZs4fmyVLvid2GY28hfvbIa/DRzxhGvcb
O9hopqBspQ3xg0kQBm421bQvntZkOQnll2ILpitVcf1PNDq7A7ib3FA4JsystYBW
y0qb23WrS+j0mzzVDqwgkHmQ6U5u13rSbFv61+8iqNNkWfqF/2NAMY+0tnNnyXXf
KGSk2NK/EDbqJrU4uTDWyJW1W/+JVgMZupiKUoMRKUctdiFZGqrEiHVaMncoxSZo
Ip1nbJ1sfoSrcAUootRb6c8EGSQ4ar+Xmh7QXO7ANjydRxxifKKFFZr0urM1Cmey
iSKxobVAxyhrOHZa9v8REygPexwOkH7I9k3Q568R/yGvfOcI9vbdQaV3QfoJpOcJ
ta+nH8tHL3A2iaUsg37w8/ryNM+CSDYoNxgFr8zLM68cp3bLXlUJLwIUHgVB3uD2
h+leoVII17YFXDrq8VhOaJ78tTfXw7ICyGhakHInvEiT2mDtPQv7tWeS6fYUwKRi
1F1D3WjVH0lUKMBoikBEPkO8nKLc+FyYx3x5jjYp1uhsrQu3aa4+DUfpar5VDC94
Z7iDfj0bsh5ufY3IjafKs3wdP1EaZix4KyIdeTl+z9zLnqKbuSg4IUrM1h0YqG+c
fsvnCAneIb7xjbEdzLdBiJjpJAGY6wVo8hrAwoIs40P7GA4aau27MjWezuObZH+h
xyEOjLHpaY2ZkYwkXjy7lZ1hTSn/k02oA5s38V5MuCBweIsCGcW/L/7t1AUDwgno
VA1LZBqGeKSF2/0SbY44SE2JY1VbLwTCPtF1GyA99Su7EVg87u7FbZXMrZFrPTlm
IiHYtmJWW4QzpckaBVya1Pv5Ew7QrrEGn5KcPlumzmMCEhFQQTgM88PG/7EeJXev
WOrXN0HJGl78tCeIYaY40BV3syHGaRqJYT2khEWXDD2HAWRNgSNRotDvkDzmT5vu
t4HGACr1M79Q6D+9nhObbjcO+uXZJVkmUXbasmKIrVZ7X75ikORoNCANriwjpAeK
gJedo812KlghHLs3g65Cfqz1uqT4YuA6g41/yWiRRE0vFtsmCev5R2ZG8RzCmC1H
bcGp7vS+2w81KgwZ57dtqJZRdWMY/6E+W1tsWSseHQQJg0LA47p7FEirnH4s5I5c
CSvI+pOZ7T46j5AxXBtspcLHR3FBrO+rlpfxlv5+bIjA8J92LAUpyveDF9veMRl+
ALagHhpRMtdT5dEwSVjAElLKKyvwDbtgjHht+GqheWjiPVYSwrCzoI2NZotaoWNE
J7UOUWZ7AcvnZuBQZgjixIE/FxOTIS5dLy1zv/avwVLbiLq5BlVVlnWXYPcJA+5b
hMnJk055JVmZDhqUJHcLH9SqGDMwGpeO5o6N6JcDY3cQA37u8koqtd19ru3r4gUn
It0Sv6MX8Mtdv6S2yhyjY8vydNgiX5v7Wssy0cqWs/1k2nhAkKYQ/J0VTs3PXXpd
Jtmq88eVQlklELCz30QSCX43GCHKDX4Q18AlbSLz07iJpJQyDsdMYkNky7cH3Ojv
jUMeVx4qwoEgZkRbL2nR2sUzjU0dE5NHAP9YPBpWC5F+xQA7yBgL+WdqOmNVefgj
d+BPBJjLZ4cBSv4j9woFQv6IH5MXlzLi2Pwn+BSvSbbLaB3HL+Nx5OYrqFva68eo
9E8EHUYfLGr9B33kcMYHIzadJi2uobzvL4DHkGSPZX37SYhmArPU1YBqwjfsA4rt
la5W/rFu5xyWfqQ9WoEW+mT2w9/0WOv788FvX3jojRdTxLQbJ/VJ10cKsm/XWiaI
zhCD2RfbRRiTeKfrgYcRsZ/eXRdczo8yI396WM5NYAx5NmkfluPydJpWia6ReykS
6Bp3eV0hJmOWe+NdS3vMhcUXXi/MvZbQXhpoWQMOe7BYZg3ThX5KGlaFFpI/Hqp+
ZPrGB3HUIkRDGJ92l2I3zn2vfmytNvqnpjwqtysCu7zhoDYGRUqB8w7Cqch+10dn
2KmSK8yapN0Ei0M7P1djJe03+1iG/+zVsyiE7ql4Hsjkc74h8oT2CH9BMs5yCkFT
uVTuBWfZtgGoD4erBU5pf7Ftv/SUPskjRZ/8n2ss4+4HHmorDOIbPUMzsDIxtsor
f+lgXMOhKEK9s/AL2q1ZtpZ6I8C1iq28ANNB9Uwo7RWx+9WUHXeRpyrQ5IjFLss3
sLq8eTF1T5YijfUY9lzFzbVXSrlZCqEoLGCNNfGLi2cIs26qx07H3KuvfGa+IQ2y
7SuWXT4QKIaoqCMvuVUcGNiyw1AAgY1LVON/ZvUJAl8EaRAjyttmbgAnkkSnZkEO
otAyYpA7LZtoRrxGLoylaOhYaeJNv7vLiFu/cYw8NKWf5oVLD1Y2R6Un3IHRGUsi
skUGaf2XhaB9V2IhP8hbQLrXRdoAIzPMNbAdvvJi20l12ARdYfbt2MJG1Od59/21
5uHeYAFqofF1B7JxTyH+SCmw+0VqmQcSU04xCtrrQD/32qj3nylTuK+R3ruWZ3Hl
chv/hvpe2avuvKHbrnKDA32wFKKOxZq6IL1LWN9KykDvdbrj2fD4cQgL2UK9uYjQ
TytUZKEI8/0XEY5euksLJW6pIyssrEJoNF2KP2H01vpZDuBX+uGewsaIJrNfW14Z
pI0RNZhp7GMnlXYskhSt+Cdzq7WZJZxC/LZT4DV/kZ5k1PkTOLY1s+tjqagzpr4j
kH4DdnTwW0Op7PHOlsLd8f+iqMbkh4+Ng52Ip+WwMvYyKZOhLcZcgAsbKMnYuyYH
xlTPAjJUvhqY6WBcCG2v6r4RNVxPX0uma5E17H4Bzm+JZwJXWMKuKjsTu5LtMwiw
v7JjUwTY13/NSLgmqsBNa2+GxBGWgzdCByCy6YvXj9l8MKiBaqS8ORNJbbMrgFKl
oEwr6TKigm4BJibffJGDUnZlKZZyUHN0sG3lF8SK15dJgPBK5+RDTekvRtDAhzXs
bCiXbJ4hbhX0l0o4BOcFg+mDetHDjZ0isAs62lrzgbUANX/cVztGRllKxYxUpHOh
NbKkEqiAY8JHI0esXZ/Kq1ePIhN+TQ3eKlEOyYFdV9Cgslt2R0N/CbxVz7Liv+7P
3QEAUcjpOFlBgHPmtJigtNoFQt9e0SyfYl4J4qbMtidsvIy8ms8PUZDdoCsEoW9h
niQethbwYPA9Le26vikxMx8uMHSx4pfRUMLFiwGaS9dSeD/rlMcMhOqAwF8pFxso
W1q+knUqaF56vB0041go/RcraNkGUzsJV4mbwbpeJUd1jlAHQ2D5+3mElrNVHNfW
iXPSL9h8H8osyLdVB8iuxejCWfPSaRkffmIsfSCLOOTiJSirQbx7S8mAvsdX0TjH
mEv4D9r99CNBsY/8ETSEIShvY41MuaHEpHblk6DbbXHJncPN44HxPi3fyXi60Zm0
Pp+3bkJ9sPbttBtxw31hJR5UzpDiODFNVkRokF9ODmGtM8BJ6Sxn/RKOBJ2VPg3/
r+bJDeAE+V6A5xIH7YsjPh9RBOkBpA9puhufa0JoUuAPDEOk0OUpnttzyOr7qgNf
OEdeRvvpwFh2Kog+r7i1OKDABKJdAyAeqrP6ngDG+CcNiDk8CLm7g+PwzDddQUch
61fV7Olf1n1Z3BrOvwzC9vjF0g2OZjuLMrpSUmGIbqMSMp0yGhHsQmWPjWitQydz
9DRXYGweYk6GSTpwOxD65LvRqe3Z61BsDc5hhYEMBDmhvITlXIVozPbm06hlG4Hy
5Gfa3KzSOMTvq92u0viTsYWCxipLEdotstlpGgzhhyPHlRR1MEGu2NBLQVnbYGDy
wrL6fVAp6iuHRwMEjFmtSPA0zsq+g7NyHPt3hkiaKWDRKfvEr25mvBL8Sah9FJ+4
xs96jOprT/CJ2riaWCtTxBA7hvww1Yu+yfiJKYwJlqK1CAbv48LdRuD5aEJxzpe+
BV7zGc31jaaOOFbxEMueZ5RjdhAPQFJQxb/jPfzqvWK0jqKshqn19A+Sitmqx7X4
XGAyb+CC9TCIYXv9Pny7nUl3H0vTT+rNMRJi83Zc/jdTYPU8CMNYkPhrFyh0Cttl
bxzhgFvrNGdxHF1QSqkGJZaudkyYWbbBos76ri8xQb5Ah8drMU84bCFVx4kTPGt9
S1bEmYg6PTTjq2EhoC0yaEJ4p9nZcgjQxl3J1sbCFhyMLe9mgZ2Iv0f2znlLCtuw
sgGRjb+jzjnqsde+XmxO/nvcjkuOyCV1vCuPiRFXvk/3ARUI4i2aLcpjas8PvgmW
tOuQIJexq68EHGj0Y/UwzTupj33ngzOeZJSGy6HWYB9u2wauoxLpO5fhgeF7hICs
kwi00BSKaUohqOg6h1RKS/qKZDT9a8nr/UUepcMwfJALc30+AVxKbceRLyUkOZ0P
pCHQae9uJE3bk5Q+6htDV+YVHO4FVZwNGhKzafTVLV/aNSW8MYXOcs2azvzs4v2Y
kq0B72BwoGk7bcJ8caELcrnDbYeuQhk2sA+iBsEtmtQVTDhmUOcnsF0MRF8uh6SR
4KjD4XPLxO0vYJSAe48TwKeg6ag8/4E6EfHNAt2/HqiGEDn/I5mhH13JQ6K6uApI
NC6bTaN2+yWSy1PjP4kE5JDNqivcKu/4cjn5NsdL7ZHFYOLbPVsXpa/ynH4lVBdZ
kND/KEhQFShZNlhhMXZNQJV2WpXorqX+4YO6lkFLMFBJcS3O5KKPQvufcSWRTMta
WY7oYsKC2DVECMhZ+swhDaw74CX1YMZNAW71T0QyuGwnjFjII2cq1u6AE+SAuMVu
IgFevIdY5jQZoocyZNklPyQXrBpeRleWTeWSHOBXLsk2uz0USAj6nVl9IdR6YuIu
YUKoJpam1+VUACAbjYyCapTaUDK31/uZnble5dDzjTMIwNg33ZLLECerRVktHjk9
jw/fS5BYI43wWnrOky/MXazYN5RYQtYO7bhLoNIYgWK7C8vGo8jZtLE+5TYaAVGa
rYtybfo2BZTKlm56x8qEWaHrHNHVfst+mb2KimZCeFP97JDM5k43yqyit0B4ULr4
K2UIt6g8Q7N5R4VpMwHF0qTV0dVg6xra058sNJ51DbUj2P9MaWnHAgs/EtnlNXa8
DEszohx3VjwnLi7hkcTQZgbMilZ6ouORhXD86sh+myuCeC4hZRNJk7uVmc7rvkcG
PXb8YqHQfXe9gtgq/xF/c/OEPvu8EkvWTyEVMO2UPpsSjVbdKwH1q9tfxJP5revA
Yai5Vpc5NpH1J1DtLzVeuBHHR87L262VASupO7uG0DpGi5C59nOnh1+Yl4KFK+tn
IRviYmezweY+fJLiWylR0eoeTqczmo62HqNq/sdBPQC9zwWfsBNi05MqssqME2sF
QEzeFk9yQ9Ew4mUBJyzrSRDWCnhDGXNq9hUr8d5SMsZzvQcbIujzw6OJvzvCaYmm
TYh8zOTEuZfmSLOaXen0q0Au7ayRkN6GTEBKakJfjQ6XKCD//xdJ+jzo8wnfbM1R
xy69q2hwxjO2YbC4L5RfApXSAcYkeH6V+4ekgdGRBDcpQHXnAgJGTHzGUmYLI0Tn
KXGMIcYLQalzISrWhgB77LY55KslRsa1+jnlrRiq40hq6h4RB4RJ7mZfspRHjP2s
/B261W4f3BZRjnyWRb+i1OIe/9VZiQb/ON+tOt2Kq9lnAEoCnUEMoTEjLM4fE9UU
0B3j4my3ijIfdfU7mPFa9dXMNfnVC0tNis20uNFAGQv+rm+CVLEmLGfhHOYS3P4V
vfk1AwOro5iyY17hTPhSX2XfnpCAu9BrdLa6SEGcnnsICQbRvZkPGJIJDXFIQxXM
3+TVgD18nXvU9TzzRvmbllOyMlRJS51KnakcTS99amXZed7gO6gEvswj8GnMXFWt
hjUsuWT4mGgYBlxK26me6sq5o/E1geqX+sRKnNpPjHpiI+MsCOAqR8A0SYF3jsU0
48qRoJqenvBiaqxpX/kwQa8owYFboup9vCS1Nc9iJrV6UsTuRuX/pWSiOVPTXO3n
X5fNijpRlyMecdOF5p7WeCOwpDb4Tmi/vSIFn27wdBPq5O8cWAewQg4eQ8YJZ8lH
KrlJUALBeRxFdkTXCWhE+B3Jx2M4cp79rvNZbrA2l7Hjx/MxDXm5Bq+Z/NeyOl3L
mG9F6gM1UgeLImFKM9W7lhpOPNZxcAtybytErO5zYK+/UkCRUvVhDh+arInq/Y60
nmwo+g+RChgys5EVrZK5MWwY7+QzIq6yPUfhoUxI9UnG1UTpPM3TjS10Q20WmIGV
tb1hzuNPbB0ouoEA4RS7R6S7IdA3m2NYLRfP87TIZuTj+yFS+ikH+BziIQO+LlOw
8SEutnoSPIBO97DWc+MUZHkiOvNh2l1BzejZG9TsFsXsi7cD5we6V/YOqft5GyP9
ZgT8aQn4e+JzD0g5J/LhhnkwTyZOCkiM7OZGAii1Pty71WA20RnjiKvxggb/AeWS
3Jo9PeMl8iwqlxRmdSxSOeF7axFbwaPVRarA+kAFkCfvDdWu4E3/WryqUydXLeYl
yX4au+1KWFoEkhH4AYbis1ZAT7gOU3ZwJVgPKIW6zCIOcHY8S+LgZ2RCpe5xX4t4
jIDFgpUrHQQv8EAcAMLSmYHr5A+uCINB7hvU0n0GaM8E710L/KoZGZZpLcYINVLQ
AIc4w9ivpuiPO6P3MYIvyQDuzSMBv0M2aV5qAJ9/uiE4lk7iTUjKPjAHmgc7zwGB
CTsujZOwKse3FKHQKhFw0BzeJdtG1DKOitLX7tB5uATuSlGJyLs6PTG10GkBd9Ml
JkXT5lucKNSuzXfW2u+EtXfMdKx1r9NldZOa4qF4/gioJCH+TH/eaFJz3xLA4vSN
tb1Hz/EN7HXHgNi1QmQu/Oh7+25sPKd5slnIhFhC64D7ZFFzbOH/YHx7JD4EQp1n
emqu+S1vnhBhPyaR+vBCfovpDv9QBzMiabTFzIRx8rDmokhHeSktp2gUzM40f/Dz
hOq8RFmItBEaGroGZaLbcK7i2TZBqBM+7ZNktRnmXDvuW9/XqVHk1x37vXXSrjMO
keNoZoqPEFZKctVvt9TKCBZJFMmY5cYkqGh7bvCLI93A0QIE9NTj7bxnkcUiatm4
F8go+Xz5KemUeEUsYLHz1DN3wxmBKP6iNtfbwEgmnFDTxPiAThA4JXyMeQESxdkY
GaZcxs4TFhvok5N2S5Z4PwKxNf2/vQrR+VPEUO8kZ+tC47zlTg1CW/zS7LO3ALl6
bayXEnV3JouUoMl9ZWMtU616lNEGBSAxcVkfnO55UZSPvBR8ukuHspkjk+ugHHns
BZnbe7iWjL9TcfSj24t5tNJ3VThfPHtsm9oqvnnWX353R0txE0a+Puc6lSKoj/IS
2Ev1+xNHrQW1n8Qe5PszBjnsYIgLWX92CDsHUBb1AS5oABDefjeYkm9oSG4/j0LK
kVlcZ4IsYSQVYBjjnrWnDbZv0AjDAbpf36gzM2W7ygSgMAoU74RsLpoYNIEV7hog
QLwTNa6fRIYyUXUptbgxUICSXeDTdndBMj/gzT5dTYSoH/Nz5vkAAQNwbSqfGASS
ibF9yG0PHI0R0gMEXDd78T0TUJ2Qu81oNnSD4MoaLEWOMwOq7IumRzUDrfNDK8h+
ruM6EI5nPYsoJ9Toz9UyyDW1uJJu+zEU3bb9e/crM4BhczxGJXI7Q33jToG7epV6
eYnuAZQceIo03fLIhVw7mofWJlH6T55gtIpZaviJUCTYwr+l/BcCcrNNOR0NNM7l
eb5IF6kx7449y1LtkYkh1WThSQOoTuSrQtE8SGgLERPo6EpMOEa9bBCNrLNxvbEs
E4NseabEGhtEyNU9dHk5H+o6k7Hfx1O3crQg8zRpHIYAKTrMNv8ve59Bx/ap2IvM
jsegXbvuToLeQf+wTq94NdEXMnupXtGvXRHStKj0XQDYaccSrhfXmSk3eR878PpK
Wp/f8E9b21+Dh1XtHsYoBdr/ZvcmsF9fe5ecikPKPuVBFVyD/mG9eFvacVl3frE1
lIor+OBhyOD2MobBvpDsQHDaw6TbgDjX7zWMMy6rgbrKptWFkPx7bHBz0g6/hZda
nVbxr+czbflAhSXM7RrR/E0HqY10pWWNvAyZgpUvJxq4CauD/t3WEFsOV06ZOY0+
ehRGKy/Ks/JhPjrN54P2Hi6lfA0kjkSVkgx6h0dM8SGP+KrwcsOD5qAjfXAsH4PQ
wEs3pUU2U0zoP8jnXTCbIWtuT4n4T8NcT8+L3KtK/59/qa/rwPghdxP8xKi70G3m
DrfuS2c44PfG0jjuDqVP7SlMr1JMOWJ+rdR/AE+aBvZrlkfWeRhj4opmgF5ABhZg
2L5gd+ewevcO5Ut2YrZ33NWIUqRAnH8OM3ExuE6EBWjOKsfmKHXbded9I5k+Dtoh
DTr4SGpfquxCp6LA52nwQD71c0XZfftP4Dtj6RrABpmHUVKMn2B/UaELxUntb9Tu
mX8Ybv8zhGK9WMssQNMhPG2UflLEampmqHTx30H9Hb6As+eQ9sh3dqqhBfGw/lCK
CHzK3ytDILE9/4cAD/B9RgW2ZkSRWEn7OqS1m/RCBmIiYPOB7fA0SKh42mDhpQUc
fjh/lpl8Y2JWovcD+X8VNEd2pD3NT7IDuTaaiEVbYntGhtujv92a5Ykupef//dCs
N7rjvGql/wXcaMt8AHWyn5Gq1Gr+F1JgLLHwB+UiYCHAK/OIDC/fNWP4hwKQDPGP
WUOTPGedUsh8Nj6zski++dCIeIqxLLO/PYtxyQnomqSLs2ANPacDUlecBgCIkTbX
kyRWb1EIBiehrC5TK7aYSl8GAPSSsjCMgAOZoy43Pcc46zAifyG6vCEzdJxkPriT
i/bAp+r/e0oY6Q93K1cmzGww6m1V4+ZA6BZKgxqHsCwM9h5BNvw+8ok69CvzkiGT
0RJn99xVtIobsqVvaXMpAC+uBqQVPzbahFW8TRo2G/wezOcw1/YB6XZ6xdXfaYn+
GyGJn620KaqN5QadC9LMHj0npLqAdqvdHaZv5Z+2qmlBiTfKpTn7YMZupPSX+asi
GNOK0KlxK9I2ydu5vi+mT0Zwg/5gTN7YmfonT0d3vsAdFy1y+VCYdK+BaTHTKN8e
q2h2itNaXNslg1VNjoH4VRo4BK3MH4gzaC2xV6cWdt8KwkNfvU9Rb9H/aofbmQrs
hy+J5hK5/HoGlndjaqBbfeFQwHLAKtjo551afX40RXKhvXWUc5oKyrHvCuC5tpAu
AWITmf9x7hgf33Kr2MyRgRXOiFjvMPbXR8Ng2MDIiDZu/n2EwQXHsXfkSHuWHM+/
9SIbYHQLtvpLWGxGkYazV5q7F2RXF2fFNoH0Snj9obvWkl+SoYim38CyRpYJwHBt
YhRLidalV4BYsofcLeInLx/RoQWZfTuA+xHkj6eT9P4AHUYCtQecw4iUDBwB8Z7i
i5SAz+qhGXSUJ8egztwL7RwHeovxtChb9n8M0bRG3INOJhngI49Ul5Ptxd3sVyj3
ZKzqbftG4BB/THhZCP9WwHVT3aFKSorhPg8fP90wkXiUGkLfHMP18+LRjLfk/Aqu
+dA9RQBKcG4BSdXUDMsV96LPmrBFzXKX469aOzCVyV4wzK4SERdCD0N+YHL6P0OJ
AkcDYNMzJBKMo3p01BUgS1s6XMp9oSnE/ki4JblMOtFWW/tV/bhcAWZWb8LPKK34
X83KPtg8YQrOpvDMuM8qEeaPUg6SsJuzfZEq2fvJyWz7cR21ZRzVfZBIhcvMOB10
WaV0pGEEbwWCOF1J+gOIQFcitVIhRVHGrE+eFiwbXKYSXn18Zp31oGRaEVV9zVVC
hbCzehlEt60ML+dar+bSfkmznCeZf2ZPJj8QMA3e5TEb064M1urCTa2SxOAN3mVc
gUqLCD0lJSrNOGUg2bjMUCb2aX0chekbBO5v7b+FuwaZQWiRK+AywNYjV5X2ow1M
OOqXxwOru4lZRwI8rU1yQ3WJhLlFmtTHveJP1dVl12qvuBMRE19CiOxnAA5k6ACA
lpQyIpnE4F8/XN23+vsBHJwTqiGlkXSLg7Eqs8/XGXUknd0WSDbMqrJD7i7CMTHi
8m9sVw/mrTsR5Z5cWc89rZtQ0NX7UyXSHg2ekkYRUdKN0RkttWtMrZbShCLNl3Dx
M1WCZsvINkNCu2RkTP1jWvvDhB8OWhI16VKpwfPJccaC+VjAjdl8bUVbLF2F9Xg+
Y5mFCJaH/lPHI4OCJPNGwnK5fYd983HR8MV+jVgKlHfQF3y9JMR9aC8kjqjjzMfu
jNEDLiZ5mx0aFpBAUCY0Rf+qvTKzUcaEarchr24AmrzjxPgsZIVbiEot/8/OPxpa
QpWtJMQnwCaNklx6L8ulRi6a8iAuMFZxeJhjfkqNmMl3AR8qZUNs1hcPOiSd49Nh
8y5ky5xT7DAIe2yExr2ItFeNBgJKpgttZLa6XMIPvZDD/8beOEEKOncI/MZl4C/u
H/fE5TEMynW2kaCTz+k5hbt2llnYM+IS/9p1cF49f8JaehSyVl1u0p4Ol4zcMBZj
AVRgdnNydsc1jzqVTzGcwQ/gAovsLAI8/GJGVOIFmp/f0auptwMoRmX52LRhsRfI
oI3kZ7i7Sz7tTSm1WN6ZYbTSo5KPE2WOV7Rvz8Dn1N3UxRHivOJVy+MKwbrJKD3R
u7ll6K9eZjYoCd6a4destMIUf2zmtccxzQ1XiI5ClZY5eezb0nDeBThKQ8YAPPJw
xO7WijvNdIXoSS3SkIdtu3HxDKeA95z+eMtIpuDAJ1Yln477+oFs89o7JwM2SU9B
BQHUSRzp/luAGYXrdjNwuDnUaEWZmN5AP3f6Kqbfpm4rhFNgM0fSMbaeuy3y+K4P
5rDa1k+ZixXXv7QElIlsvKfLnTAASxBpYJmHRDmES8iwSC2a23gS3KffcxevZ3Yl
gm9mZCicVLrV7KxPqFZ6/AtY/r/QgUuV52mYbC0i3SiwfN6rClQXKxHBEb5oKd3I
k1cRXf+XlId75h2C4nFJgwOSAO439jXVBmD3yp0wxw0LxBCqesAlzD8a71voR/AC
duCsyg0JbeOvXZs7qOluN2QAXMmJPCaS78zXGbuNwKvpokbV7lDE3oPdIprDSdl5
UNRo1Yw7nGrecpaD7VGbifGuOVBbpkoIndMeJGFh6u7iG6xsRKi4wA7RozFqqCof
ITc2aFARHZZRx1fsbTDMuc7K5RR1yfcq1wmBmVu1CXjGI/mfCwP8yNIITsJgjPMh
wfTxeDBroRivdHuJA8LaW3Xm0tpil/vcxfmJU0e/H4rRY/annEZLhPSZk6iLZftu
XwKsaM8cq8BuIVGN4++WIZlhpURKGX2P5RSRPnCqZsArqLiEuyyzIatwoOAYRO2R
as+qDHLcasbTyvj5UCsVMIPiszE8sDZYDgkd3DZumEuagKCO8D5Qm9Tm0BtBef0Y
1kHmPRzDZxPK9jTIeGtexiLoM0itEv/N7HyZOHNN6gYp8DejReStM2DTieE4h3er
5hhGKZq/+np659qG7BLL7hwqkz/91IlvCb7wQE2EFre8hiXHqhhPIiZ0KNAA6PRz
ui8deBQacX7DloZzOILY/BjWH3ayGFXfsHqd7lYu3MVE9LwfKCh10/hBgI/EpJeB
OqaHZaHekmBQOmOPa1XJMeM8ruQG7YU8HQshlP8NzpseHjrLoBsLDcE9gMscCAHC
OLGOpkLSN0bBvB8f+29wQ4ulX329FbOYP+5fLowDmY6WNFmpCF4wC7SQteyoaHFE
Aew3jRIfx8lh19ER7wdzzYCDSuGJWqwnrBONpQSYnzIIx5LNWCkIwLzif9JW66Gh
OidKNLMFb7Wgfv9e4DDE9bsufpcDTBFktj4SkoKPsh7X5f5aFgQri2vYa0tSUzQ4
ePNoNUF7sdJgYTcX+NFeLo4YdcpKWPeulCNuw9NC0kr852z79ZSwdyEKVJpE0wFX
ExOaK71DDw2fuwrsTqp88uyPQ5v+bxJCw5jCzuUdxSdODXyqfe6qm7pKH0+8YUSZ
iBzmNxpnf3yfeclP9p+Xl/5iQp2PswXqLmjwSoO4lMAua1/Ek2Ika8vRqNQvl6Yf
cMN+p2gJBj2+7CfvkeLAVZuSK7wwslBvIWkRp3y2bggFU9U1VVTUwk/heaAEi4Vh
PxUCjhqLWuTqyu8DQ9wYDD7U4J5GE4jFsxEVsYlIFSNxt7JHHEibkKbnzjsd5C9F
T2/kc/cf81QJCTp82PV5X4aZ5At+eUZBBYLsNLKXgIIkUpq0BWXN6muOENclZB4j
5RHRTyNwg0FaVRox+add8x2NyniXpGtwWR7xErRElaTzWYImZ8tduABjpRTbx1Kx
fGePHRaYkDy8Lg/7j0WfejLB389zU+Mg2cfQ32Msdj8lb7IAbpkcQEbWbp+V2yxI
6B7oM4lXgxWDlOVXXGnGpQUSdxhahRqMXUBfSPt3tljpiWCze6QXXOx0SxqasY+2
2PgzHpeZfAJ1uACtx/sVCo86IaDA73rx7V8RaPb33IlIWDrRMKx/Aegz65EnOaX4
C5fKADjgd0jINCq3dD3o/z5QF53mYmBgdrN6QbHDUw0cPRxJwr1gMTIZVvHWPPMH
n7S//qYQKL9bbvc7E9OzEFIEVA5R2FQ/UMdAXAJeE0j4/uNXJmN3dsB+KsPYsSRn
MmTZn26XUdhXAE9h3tj4mT5siGSEPt5MSfmv/Pj+nD0t7KOiyBMOyvJ2huBVj/tE
SitWKmBsD8eHwO4it42E0cVuz6BR/ZaOpoUxTtLMBKy2L5oEp9N1C6HhdV9o/4Tz
yqUoSSSLK5VZG/c7VPHRMabcDXcm/ODjtYDLlmLMqfGtz/8WmUOp9TvvpkbHjnqD
LByqYjptcK2wUH8wlaZSBrOa+/zAUZJ9xDez/mvXVQadsuYDH1LTjKOlK4gRVog0
EZ+iL4AD7rPFq4vzIipsWjaIyoI4bEgJUnNIHAdyQGqbTFPaozEnzMbnVBybaq+s
1qpjnCOx44symZSNHHIneAdbuKtV3cDvMH4gqsdjRFxYQhHG1rADAC9dN9Znb1Gn
f4rkKcIxKqIIC09SWxIVqIdXPS0im8VmyRCfatWPtCRh1FyVub+BBGT7XQJJoPEU
xKY+DWmJCSOfR1815/TpBL8Mi8gmPyJMqeV1aVfwKcKTrepmQAPTQ7VAaBQrJsPv
JMeiRB/dqIWm1e3Us04B4+WtilXxF0cT5mm9CIRWw7HjX6xJfVp1tfnGAVcVoiYr
YZOnjrk6jNxF91uPmvU4+uKOqRt4J1JgA8aFMUY2u1VI/BymbXRtwyPdFf9abHRt
TSXeyF+yy74VPL1g4z2xUFmnWPislP8e0tY85xXkgQkr4sS55woBrSlfeoLNdoyZ
MXtuiQgzZUIZq7frF5Q0CPVnzVQAiI9DntPXzSnEnxoIpyxvC904TAzH1tfijBeF
cG+UAXlj05G9+TGB7ZmjmS+zjc/XQkr5HhkRslamF4zjC4tOI9ZdJQ4U6QDgCzqd
TjmKM+G2fuQoVIezd35+KTEGI8AXXTWsAELXz6H+e0+vfNQlHORFiP0OnMkzSS1L
sWibYaVYxlJLw5KBdz0LzzGou48fPwWIQ11faUBIChfH+gPcnTYqF3fV6f2qv+KL
RJMt4Xa24Bu+MMwI/kA5Yu0D4+OzjgLze6bEuBPGgGH6X91B2JNGmTR4Sv0WC3Xk
4ITIVUmcnpBH5YllmUWPzPrc9I63n3RtlAaGQaUx2GAJdL+61kg9mJzrxEmD85HZ
YD1fFgYcZ6RShTVvvsgK7BpW5Yewrzy/esH6aOhX0DgU1vUdNvBm92nJWMOR+cY4
t5hgwmLGmHfOT0idXMwCgfU0D5kgdK/uYUmfBCo6w2Y2GN2BlKCQGEmsNT1QcTKg
wxfE/4dA8MpMDL9/uuZhNdm81hykl1OyyKl2j/rAdpWgp0ABIqmQEtF4Bd+r7mDG
US8bbfri4ic4Ez2LceS0Jz6F2Lw3ntv93vuB7X+TO2Goe7+ZhAzP4sheGI47wO4/
BsN5IXk/yO/BjCStX99lssOxst0PZVwTqG9/X2qEJmywXX5WuhBdXRJXPp3xWIq+
zCM3exDIAHsiYUAG57TPwAIn3aEeeSjANca+Ud5ky3B7h0TH7Df126MS1mDWTQA2
ffeknImhIc9rQnXQfjH1Huimm0AbnPPRcYUndHwAe9VZTsKc1TGBKLNgm4fUeg7S
twici/JgB4iOnvVfl8SWJpMALIdNhhOAE/4pB+SAsqWksnigSNLOxigkLgoP2rG0
SU+a/1bTd415bAZiicGqDirbwjI82eXkdQXb4v0Hi2NmG/isG4JsW3GKODAUjZhV
q27cb52k22Fk3Prdd08WRSKp1qVqdJc2AeL54WwfwUNm1imkeyCrNHZGpYWPdPfz
ZHZNG4Q843XQyu76A4dSPwUfAs1GZb3sxuDVOTTJXiTVGS307wW5fJwXhri4n1G3
zZwiMNTCwYYaDE5a8pcoMeEmEGrfLXn5MD9h5gd5KFqrtXImgFxUyxhns+Zy7CdL
R/J8xnxBiIhQf1WVBLWZwdoM0nJgDTgoy8pshOVFfLUFyOMOtF6dVwJ8b4PbRZ8K
KlZK7nVlSdKpyye1Hr6d9dYueVhWPNNwS1k7JonRODfqzTK0Tz+tb0ZicnjaQejX
joRVeXXZDTz/6Yxhjk8b3JywjN/Tck/daaUvAKlnaleSCsUJRW18xEU+9dszvt0z
zoCgh7KdDEkS/3t8NqJGvSErMYX8HwGhHeXGdmBv5DBcyeoLlpQpw0Yi3X76Qald
xbTvbH3YLPAvZhQR47m/mp7RjyaAOScgR75SpkFu2VBmiLPiO7lrTtdGNe5lyB4P
HlLRGFrvG8bC+VC3YVVq9HHztcGGGuvxWHAYDLfbZ3Hy3S5kXCQSMOP72kBU50DO
FKZYiWIyL+R/iJC7y+f0dOqJqJfhHvP8HzIW/5ttfArzruk6yKMCXslZNjcxRhOx
7KddLaeg+pqEeeXrnLB3cyaju506l71arXo5YQ8Fsiqa00BHIxzWoJFDnnqeXWeD
T0A0Cg4D8GaS7Ab6Z+9S5apXCJLr4CaIhcapdeWkjiOY9qZdzHAAGquPultkLc7Q
1YWdsbQXfaB4rjlfVuYB4Pj0xcFRjG87ZfIXvfzfusAE+qNkNjEa4PRWGp+QlDSj
aXzcC7gDUVr7BM9i9TvCQUD9KaA2SoYhSTZf6QUkj/01Wp1UZibDmkULw69fW9Su
xsVr/eL7rcyASJZhZd+LtRFRxeJ2YHEfSYy/93t2TZicKMa5PI+nFszE/fGS2I10
ljovi9/6lQz9f6rOkdSihgTKacdbQJKLfG6X2dLDk8IR2j4UcRbgiQuQRfloF+LB
M4CS0TJHk1UhSygXBiojYLtf2VaXjW46Qy2Lez4gMMtbNtyjoucy/QLT8t+O45W9
bxlochsjk6Tq7J1TkbtZ0cHvIF58NFEjDwzoJ7BbvYfOD4a/XelIo4Y+p+qXUrJK
Z2kr3kNjmvrHxMa1rz8PoClunPr/bObKoZ2fjjdOCx6+pXR9Zlralylk9nLiMFBe
cRBi06+3x041+DyKtNEvad/pQ6jQMTdpyW+U/Y0u6pOMtx6caMFCP38wCzkElqCV
IOR7nFfLhGVqbhuie7jwLYX2ZOAaFrNpwyWiYi3zG0xBz7jM9SMtt5HPpqTkQHt+
fo+XVlM54BMSUEr3Y9xE1lpy53iBr4kMBu9lszf+LKyYixwuVCjnYtWU/LPi5hUR
+Pg14Oulvprbeoz/VcnA+aTsjnRY9+wiYRTjCmz7R+7YnGesKgBE2+tlJArdxfKo
KcQN0F2SUOigQ2YaoH9ITF1o1P6jS2Mdfett/+XRUp2wf7rGoAhaJsTqBqvqkzre
dN0Q86AWNDg6FeaIs/gXBm7SVAnQqw256abYpm7LynXBvQMH5zOkTZOqYLMa6VtS
f6GGHyaR+15NrPz1zc2NeeUCm6r/GXUE1vZh3/CXmRISkPxOPOOeJlYw13sdPrIm
zEEEkOFO0nYT7gzZSqVAfx9UoJt6IXrmVNMoFG9AmSuGJUFvNgNqGNWxNy65tDRW
5LSuL5Eqi+lH8JKdpEaNaX3zlTbbhkPkMNV28BHglZS8x5MJchPVo9RFIbUGnyQd
AZ/PzMoYPdgodAmgCPaZ2Q8gU9eoM1iDNMdMVpPnfwZTnAUjMFDiPqTSKyyAfrq6
90CHzflAsbp5eJf7HFD2ea4WBtW9ALQE/b8UzwxXgtnqkYi6UGQnivxqrbtZvZ/X
RtZ+dyYsCqVVWgT9LLgRwmd9D+uJjN3nCzACN17GLaVh5v04CJUlTSmtjeMqDfPi
ENZZ+qYu9dZbbK6IEk6uXz6Mu3g6oSnYF9QIXPxrWrBlhYwZnjt8X9PIAgesJN4a
dCvo1KOzCbOu2SUNCCHYKwQDXqSKeXMkwvrbwxYop25kmKPn4r5XiSdiy2TaFkQ7
6HxL9hkq0hu47NeTc3GXZe/gwsth9o2WgzlAPnnQiVGukJM0L5mcFmMfZeQIWvXU
keGO6JEmuvnDXLJQbApU4idwuiNVpRCk83Hs49uon9s5CuBRxinqsmGEwdg0aXju
9fkH58IJycn0G3ilM88mYlPwVv6/cZGLNPh8s3gyOQ+Ajk6l3MCnR/TeFxLBhCK8
L55eflDSLcVRSW/+tjAIZLtkALmZGKHtY3kg0idw0iC+S7S0se0HMT0Tg+oj6xDk
wUHtzJxXlmqQKYyZa6NRywLab6rMGGrAeKwZkVEyHvG+WEDUV+uuy6rEBmoKbZR/
DBjoJD2ep8CFVSzzcQLDzh/JJ/ELzZG0vd2vWH2gVyivWVdj/FDkmsormf72gLM+
YiLqEeVBFIoGqG2GbdPGi6nEz+DELV24vMFRkw5g77fIVGoPT0zIslecrPJ+i6YL
6fRjiVH0svN6U2v+VF5wXTwc2I7RAYPj5eYfeQ94fmogwHteDQGAIWdytx77XaHr
vSMK50aLsYJar9Bg5jCp7i9/W3Z/WUEY78wJm8U2jCBTE3jpP+eqRQaEi6SqfHLc
rSz8BVYz+ruTrc3wrOcON9/FnGi7uI+CU3gcykxKJsIrAsE8HzWz2vclNBex/v5L
cTx9ENi54+Pr3bHHVHKMYA6tpguXB18c0D5+USukLSltvnGEBZZuLRjWh5EPb4A3
RpaiFDdb/w0JFHJ1ZDcnAmEW74fKlZwtmG2s7vRgTk/wJxWXpGzwMOrTsi0BIxz8
qD9QkVy9pNMSe/7szgOo5maWnge5f33u1ev0sQqICev1q2y9CqatLPO9XhjKW7m1
SksrndUnITznXKxreJ/1Npxdaz+Y3yFJUc1K8C2K4DG9f1084WC7oq6bfK1qTKZ6
+9+0JMgfSbeIyToVl6eg9MlhfrOZ9rwIndJJKXPNNn35U21UXnJ2eLmpSoadopWH
XKZQJvG4RjHXuHYgOSFtZm4smy4u1ymYLjyQ8hvd2YY5SNhpCTJqPcRku+MpbVIE
AXxcWruPzAVCw81v+URsZGKQlHmX/QuHwxp5QfixU+Tc/zQBZn/JIgaOxK2LbK/T
WnuxDISUHr15kkvMESCf9x8zRpSrV8Mrmfonfx4VpOsXHJ9+8CwAsiLD+idNoqSy
lLhxV4HxpUzIXdscDiG17ZTNTZ/qVgshWswq0jycdqgJFDKqHjGMNlfbEHSmeP1N
QwRNAYEn6rFd088zUuXI9z3R3A8LhkaKlLmlgO9JgUquZGYOy9gZn7zxhxdX6yFf
ntDFAfQ0N7fxroCqceIsBTrddHDUdyDV4fg/1fdFuqhW04bofLM5kN3rQTjGshJh
SfMs1vVszLUIgWerSt8h29dK3qFMfWsF7h8dfIeeywXptGYUr0vx8gWyXQ7gpXm2
0iyr1Uka4yKUd7jNc7gAyuMoNW1EBettUUATzim13ytthEZbXpd8aKTIVble8QXb
DOrIJZAV+zq7aKpBf6unkL2ev1J0Caxpe0ggZ1+EOkIC36ArpOjeT8aVYmYLoHCB
bbg0EWtFKGI//m2I511WlKHY54W1hSIoWz0uDH7AJr/pqPVBlkDXuhIv54DFRMCG
cMQXmjSsS+vJW+avZboCVY8zB0K4obzqvEKDPq/y+VMlznm+Z3ipjsYcfavfgx9q
Zz1kuZ/ea5o2un/FhpZPz0FoVl0f89MVEGfKuPOwEdju7mhGBmSWCfIytwp0iQUi
FG4NJpkBWviNFrZuC6cqlIAnqVMBnU1gRFK36ySes9PAjIEMqrmZ6IkTESF4oLv/
KQd7e/4UUqTbV/b1gjUTSBA/2uKBquoz87LdFv+jxJbJd5cVQc4eEcxrwB3IW91l
gVGwHyHFXgihsUa31xEIDhpHTh+RFCqhy+huef5KRz1D/eZWoCxzdChbI/RBxsYq
F5vow4j5oDIr3rqHGzKuUvHbbDEHg+R51Nk5PeXr8SDObfylvJUP+7QchhO1Duvt
ESuQiWGe/NbqPxjEzcSyXtfLAVGFWHjT/F9wKoHG7p6unZsTXTVncj1NZp8IvbU6
nlPIRQsH6BHs53wBXPtT/zRUGZB7fJYHchOokMBtyTvNOpRsqGn9Yv/e8KT/JlsS
UzflKdqpXrqxDXZ9WAx7ax39365CXSD0h/nw/4xel1AA3lVcH5pPV5Ax5yNLDDWy
o7jvdIst+0rXqMNGNe43QqRLYHTlBIwXRET6q9BUQ4D+h7Y9INKJfK9xqWFEjOEt
wGF4w9Mqbp3dAdg/TpPr1lupdxvG8CzsI/DGe8eKzs2GU3Vol5M+R822xerWry31
tIgcrzocsmIUBXIZv3/WIzUmRS9XcNiFgXQukVhW1yNbVAniRWfUQZyRyxpbtLms
Jnzl/kUDClU7dRIWkbyC/rLC+lNKX6S1CsIwKDyy9HUeSP5yCB7twizfyY18GLav
PugIBVwTZq9PtWs1r38920pnQOMfuH4IJgIO3ZH4kx6w9rGMD6hFm+HJxUMHjWui
MnN1GknjNwdIfGW3tGqsn0S0R6JiC+Ky2xotg1/qUFzQ0O/rqDwHPnD22c2noVAu
pjpho+NvIrdwdVBRo3kF402/v/dHMxiFk9RVh6DcDgzHEi9vZHTC1lDgTckT6ee9
bYVvOWZbYDCqCGUdfXagktmxhLgGDTaSVD8Oo6RbOToN428W3Vv19i9cJA/8e0hJ
REmv/KerjpqpET2yqBfizahS0LSzsjCluhtrAs7xQ47Z2OSt2kfUjub34ggaCTKT
NAU3NCnNoVdL+6pYyWuaHdpCbxAZoE5QH86E3TzmPNR9dCKj1EWhD3oZDtyodA+i
3GDrFiBSLmyT2ZKg75QWyhblnW76nqjkiv3w67e4BMj3bcFb1HjiVG+afylIt1m2
LiorBc0NOtxiGunNUSy8rp+IEAXtHvnmQSAnfzo8MbxAulhARIDmgCem+q0ok6tN
skbLD1Mubn5PY3PBhLO4UpN9vQXB9EyVkmZZdzz1nUO/ZsQFifmiymDEyQyIyAB8
kgERT3YbUAS1o3VRwCOswzfdd3vNuW8IpVzD/7us1pmijq/LIy7cgsOI3b7OJVbA
QMfKbe1MPb8fCfkuWKB0kDrj7JPOGhKMKtrG2jNrtw4SueR+Ahm5zoIX/c4c+7oP
6e7y3MABLaiu5FCQkM12sPwDl7yjKUDGb7O4f1n5/4Vz/Msxhix3Bvdnl7krI6mQ
WirPyPaW1e+TueVameyI80Q8yJo5vHyJ/QFOclbEfgQjoja6PlwYZBqmeOzFWTj5
AIBoE6oiRKW7OIcG4OGNouo3Zj5bQXdXgAIfGLKEfuIF+t8yrURzX8EBDU8w0USc
ADQWEZ2OW9DzEGkmRhGniHY/wtvkXlpS0hcShJBY405kygGa5XtpBDQuiGjelL1M
Upu/y1w7+nlTKFRtOftIhRL3PTTwZm8taNumLVgjntihNCW6qve2wEnarLrKfqg/
vLworOjFp6noBfdP0MDSzLv9q/pESRMJsBkFl6Odihn3veBbXJJ19nEXSascwQVm
AuuHsCeKaF2jC9GAhUIZ2AXMhFxB2p5cForQ7SUDgn84QqDCJmQQkg44pL8hvIYX
q3Z5h5zZBKgIehj1nugdPmfc32YcIYwDHrue01hNrfznZsNsK37OfVq6QQSS5Dsf
wdZNlV/U+iuvG6e13L2MN91ZHiCnc/kBwLmQP2TVbAYFBgQs13X+t6r8RWSHQiBD
dE6m8PYiqV64Z2jeJeZp3DIP3R5VCyLsPH2JEbpEwodQlUYNm2lXIGPzy/VW1bvH
e6IYVGL/j3uvJnykxzM94Gmfy8RtS5T32VhO2watxO2ZV9qyVshDvRRUKRI5ps1/
6+umvQwGU64D7OZWx7myb6g5Vb+Nn+YJNaEgY8gXMDTOVPT63mzS+3sJIw1HEvkO
FN3CnYDBYDKdAMpXl0qoXnXPBiPY3oSqKDmqPyvqhF0zOuS/TqSQcIJuFbfW/qmh
Z2rVjDj67jJqNhIwn9jP5cf6FcFpRG4fao6LK+qpi4Y0uanXwydOkcj1Z71H5z+W
UZ4tRfn9JKE/Xgsy29KJLpdVcIhTsuQvz/ww/UWY0tGc3Zc4B/umPINAbCaPe6ZI
VrbTInKQmZvj3VsJwixIFLA8ozrlhsU1SSV0NBtdqk/3u0RxaqgHVzn8JYR0iH54
X79E1NLAdKBc+tnCOE6NZUWSbYM/DIkJoqqmDRDKVmpUa72OF0WpvOThJmmkC+PL
ks9Bp/jEPWC8py2QCJ5gmirhWJNPV1HAh5Ch1lg5DoxbOWiCU9IEcfWOyZd+mgIB
rX4v0r+HCdM6ibLoODx2sLJ36jvWkZEzZTINOs2D3mhqK6a1JBxcnVdHqkNW6AMq
hdmO8H1qXBlee5eSXA/dcg5tDj5eoPR1OgbPlYTL5AyrKpSDSwcc8rlA4fbXZygE
StHeXV/I881fF5rfDUTX4+xnmIQ7cjbK052bz3XFFpqABG0AxFOOj/eAN1t+uJF5
F7Q2WbZjSolCzQ7IWs+k8msBi8voafHLM/yrQBHUdxhW83esRkEi0VXBkQvOI3OS
NMC4zN/b4GwFFM6Vao+e6qMUiJdJ7KPc9CIoYqfuewmzIfchfIeRyE5cnszN5u4/
zIOZ3Nu0kxpVOsJuhC4YbIjDtrONibHyFxG88KJi6i2LyATFOtlVSMNqLrL/PudN
9EabQH736arcp7GTVEgQ/Fn2MaI3dThzTDK6Ug32eg82TWxXxwXxIKjKozlkB3pK
0DI6SGGqbcdJ6B8opnHXIR4Wffw0elQqbdef+B2ni6q5Ca2E2kUwdqANOyTC5pKp
1cjLIBddvUUc2wfMVfgeJDQjhgDwE7kf+ggAx7YyUP8=
`pragma protect end_protected
