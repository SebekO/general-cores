// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LIMt4jKxuN/WtrmLIiFutllCB2/h84wNdogKp8Pm0Zwk1ukyYNu/Hp9tSwr8ZgxI
LKiiVV3h1l2za/7sLGpRu5Be/qZ4DOJx7KfRkaG1VYHtuHRDEFe9T56TAC/hBZYf
u9pEtlG91dGvP4c4ZpHpNvQPu9NpsDYbnvkoOr3pzFA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749632)
JDCpzEOnoHlSvcCcDbeu0ooPJaw7XzbTVr3r4ucDOklUtBKxdpICiWQyEPPx9G5r
ETMwaP5htiLdX5Xhy8KyefM23nPtzwir04R1tanI1hhWDrZZhUpX8NzM96Tc4BwP
IkkEOh4ddM4gGZKg8Uqli4dNcqNZuuOXJLAsFeJa3Gg6ICEYd0BFNxvcrD3zaQSF
jibvgiMbQo24lc0AF+r/L/Lpw+T0QV2aYxDNKa/6/zxM04+UsCjo/a/WzSar6QQ5
oZwQC24Ngx5JXUrrP97lZ/s7KSd5Lz1IpQ927dUaEBFlPgHCS91wy6Wnvb7QKKu8
xpFTwKYtGRfqmsSbJYWP2jblcQdnBV9MiGlvHvQTaVxm6jpe2La3mUXQOCkHWmZE
K7SUGtnQ+Q/CMgVPm/qy+mQmi9Yehxc/kkNOGOCcLpLHPMMcdAuo9m0DIweZ7g2G
8vJVUMy2rFRLSRcKMHr5nxkWL/f4bnWOyDmbjQIs1v6SL75x8+pL2EcrObHrIECU
oL3GJEwf+bRmithlOTU5kk4MDQmo2dj3olxPoSOK4ySs4U+QSSIRNQsAQSb6zAvq
Lr7JwnIoW6sVJ1swiTDYZQDLSw6MsnIxkf9bJHSzAvs0mOCMOR0XCcS1OXFJhjiq
We68ONjfaBvMs0QE0ppWSeN0P5RBKnSOMZCcxhZP0PdCk+Ued2AgS7TQVPmsSYb+
S9Wt839zBFQZahXAYN5Q+eGIsnNxIOwgRD65Lc80rKNSYVTkah3D9X5yql/zz3ym
/qNNqpUhOEzY6Syod6WYYXBTAp2Q7++NnUCuuPORGrN90L5jFXFwqlYbZ7i8PThC
gjYOO0wRFNHispw786N5j6/YqyNkCOLvZsmYkPyd1xrFHd3RkjpLk33CuN5UxXwO
+W5072HMGHarLUC71Vpw0TIsJoNYQYln4uaOtpxzakRL9xH0BDgVV7YEElzcdLgY
7ND16dvV+F+vgYa6YGAbcsbv8CfzikdwHb5EMsfvwIOhxTgah4YOZtrHhHELQfw8
mPe73QAaa+HJJYTb9z1YMHC+nUPCG+AUwCFfSvxH2R02kw8hPSMgZoz5y7IprWa1
UPTD9A0DFgNYIGPCAp4bINi+PCfet5oNY7VuqoEYhjbado0qu2UkTBKTRPNaBOba
sb08RwlRduoKhExgDlGswaioQf0TChe6bbN3/eu3wX+W06nzoS4ngmcI4KKxTUA/
fJX/OFo0EaFjLc3lAziJ2tJlKa0PkgdsylkiucD0FU/aFtUJi/L33osdj/VuEfPV
6hIXWeXs/YKlVLBoAtVvl55SJpOnXht3l1DxnT7xznM0otPwvSAYxhF1lV2dxkBc
OEAHRHCjrUKgAkrad/4Nm+mbTmD4pIRvR4CKZrmne2hWHMhdmanrkww9+JZFUEN7
NZjmjnp1l+zEX+VIfCDofoqZ1dKNzMIEbB33jXawechFIStQJ7D7fBc3YKVxqbVH
0zZjZLYStEYLfiIxoRWpRHNrOKwdhYY2jB1HbQ2D54gChq5fnncpOofJR6Nfm6aN
Wo7UN+JrwzMI2a+RHwyJM4ZR6pa2u8qjRd3SAFSg+4Hk28UpIuGvkIe8D6Uqibyi
0qAty7GuEi8UgYwJuNl80F/nYJDhix8GYThxDN1lHObjqRibyPAZZAD7eJ6Eyi/l
3PEkxtvLH8P5ViKH7tLCKrEbn23+pN/NPql2+tbPBcO5zVfvM0G3aR+cvUiqGj+i
u7RW5hyb31IsVhmqKZhS9yG/dR29yd9dTgAvVTPLS0P4l//vwoNBJjtS60WRNmTG
3e8x+OGON3PjFKA1ohQnzHl2Jua99b9IUnLcExNBmP9SzujEZHaFlxlXCAwl0Djm
rFvA4raV68sNoWYwJ6NtKTW+5fu4ObLXXDqD5rP/W8kR23jcPZKPXensB22Glcj+
wSaag3or0pTa0HZqnm6IPX/R9lBFezLKRbPNVD9Prmu92GMdcbnVhWZu/VHKd89B
xUBjtqPe/DkXki9HX4YK8pPplk2he+CPBMcnxKMOSQIj93vaXnDxJ2A03mhCxkRm
ckhhO4tpw/BQOshfnXqn4EsHk9yqpdT9rFbSqZE48vu8ziZOhKWoteZZXywcj6UX
mz4PT3ccFSyAzqW+GvysDC/DkgxyIghhpexQsORVnkt/nAkZE5LX4mI4JV9qjDj3
knBIaUwoo3XGWlfGS59KN50CDNbYG6iwTKGxv9QcB7PG6GAjl+EuWdBApYyKIIK7
wtGUNEANr8EjY0IkzeOEHQYAVDciS6YRm6GBkEKL3Ed4S6dRr1u8QtSbMZmgICu/
ax9nlcHyPCvoA/VbS2WwupahLgykj6mXcpIJNO7D2p+65Ps+vhytmlcrX7f1zpue
vYYY5k2FIuiMs7yoiqOtn5OXiF5xUlqc00sa0zSzqpH1eEW51nh1q44j5V9rkQ6j
8xN5UMlrVM24ow+TTqdVvYQu5yyF88eoZvh0JpAPTtR66pboPKSkFP8gZQOvZOQb
HYQKLqRlbOe0/cDlacZqfIvawmAH9Co4lS+GIhnCkpxAnZM535dF3HiY0oBxy27V
JrQSU+IXPMZd0kPXsPayftELFhRGfuQ25I9m0+9AnUBx/+1TxRLJBo5GUB7wcjLj
wW2mAO4D7pJNEOSqs4LSJwQtQMU+NW2JjrvTv56dV61UwgH+28HxfgCh1OowZF6p
5nAkGtwC0sss+lketxXiQOSsBqYe7EPrqbfCfeeQ7AMHr3GLNVEpzdm0nAlqOato
rQAxlEatVPjf8Fv7W2mPbs0tOK1mWrUAY5mG16UK8AXctDWa2++P7wAaSQhWLDHo
fwHC9w38Wac8AFYbKoPSPxejrxNS8OekP/ZB50tEDNHlyiGcrFWArdKZ1+f2LWqU
ftYkXnNrvAo/GAcNHK2eWc8JVOHupD1YPxRq+rlNbDkXzL/It+xpcRV5sQPmJQ8u
Q1RlclTLhbulw92v21XCX0EzP67cwbzXIg0cdqUJvlul+phLlK5UNxd5/I9ajHwX
aWVek9JLk/4NkaHI1Vy/mPZgK5UOg8RiIf4tVDuwNYHKm+ZtHo+LOjoBH0ctnm6k
8aGuMWnuLk2MOHSNVt51aiNO4edsLb7Xdyp532D5gb64Mf6xdRPSixjC9i18wxnE
e7Irx7pv7JE8RDzrO2QiDUSbVgoG2EGlfobnaX+J6mpsJL36p9nNcjZcypVq6v4b
OKBouzw/ucuUt8dqCfz7qJV6FzQ9xqV2iShfidWDy0Iq1/5708I+hwXZQDdRmTw4
S3FuxeJ6ET1Is83j6OanyCxD86bpItYlKwsLsAWvG9U/Y8KpcnZUxVUnK6Z7hue0
C9HphW/t4zbf0jAUpHMxfFjfuvzuAz3MWhEBmzXmFTpBjToofVWUq+Hff+oxE7Hb
Ijz1cUK75Bzq9zRQ5cXe1HHrLbY4D7zfCwdQLhl4Tg+Z9Kg19Lp0K3YUwBr6rSKC
fG6mq768u46OU5+kzCQbvbl3wyZVQ8e0oAphLmGJVTsme0yndqyb6u1HyDTKZxrN
FAVvHIkteXNXdsDJSh1JBM2N/yjtk8paIlquXeGmqbIhht3v8/3dY2GNtKWN5cf4
csZQKHxTqUTTApoKPJGj96UOPS7qPehDWlXXWrcs9/CzMwj/4AFJPeOokR/2NNet
pL7NpsQLDGOjq2YOVAV/pdrkkaVViOXR4H+kK1xDVzQ35Qu/rm9RCOLeshpAMmrj
tJ+gHO5LpADziL+LgHGzx+uxPfNdVN4kjNfRAa5K0pFSQ2wMojmeFbtJwMPwz3lD
vqC+NPAq+c2ZMiAUhraG1yrM/VdlD8qdBX8CYUKl9tzJjEd6TbavWceq9qg80tPz
sz00FA/RPZNZoQGfN7UzbZ0D2heWUfiX9qP790X47U7BYQDheejk1iPXdEVXu5nq
EeUVB4f03TjC6kqbdleUUFksWhc0iCvucEnesxfo6PTnfY9uXqbWotW2LjpJ5vsT
JCIpkm/9w14W/MQ0jDw2kIBadGurHeEApH8PU424A/F28PZ0lDP0T9bbOCiBs/EA
lAVm4F36DNH3mroDLMZg4JZDkeb9VtENlBnRfoBQxDa2OuJIso3uLzxKht0/olhG
OxK4twETqVxt7Cw1GYd0++NuBJ8w6hgUxty1n9e1dbeABNx2Q99iBuKyAWfhZ+CT
aIFwE9hO7cMv76qj/ZUhy+Oc2NomRyotFsJbjtVJgsKBtliJmedSQFbvr/Kf8CQb
oWSS22YC8UoySlzwl1yjlpLDJakb/2jUcwSjNOgNMLHNO5GV0wOTdWbGWdfCV5sJ
J+0+10srcmve0bjFDI1fSTN2E+W5EJEciECb9NpZkup3ZXuLQvHfx6sZkiF/ZcCU
dyiLLfeS+I1UUEuPW7bOOcZwxNH8k1Ws+i55CWxQNOBW/aDLjWBOjq62fPdOiPcx
H1f3JhY/EHgBiw3CAkdlha2cKyfmKiOBjBmOt1uRN+kiA8RZaJwJL+V0CCDRdIMY
6qV9VRtxFwV8wruyvWXLB4/aglSk53nlS6ckAriVagf/f39H5W/ZQsLgNSdl3YBD
/BuPM0nlHNUsmLEizRCsBMyhf/ioCiOz1r30OT26TRekc8MSY9XZleCmeIlgFvW9
ADTBdNuPqUvHQHENUM7d5yX7ZL5S2Fkyb6tJpE1+V/gpQNv9yzpYaOVauvt8di5t
Id71AX5mOiIXsSV1S/E6udrQx0lIxdEwwsbawV785C0wDjk+RtmOIlQjH6tIjPkn
3zVRsBNuMaRZ2u+PhiOxBLzTtUUjXJHlxF95RPxQMRcEw51s90edavS2ZP/Y0lVl
vg+4Hs5ihbPpi2/389xpJbs8p6Ag6RpT28x5s+xsWKrGoQiIPz/JEHaxPTF+DBGo
UO3HCokOGBdGTyWUDmUjgOUhmUNYz8LoYmu6U1QEgZ05B9gQp+C2p4/tRSFAVQe5
mQkAKopndYIVzCgnTFTh1Fe4BxpiJcSvL3LLeO7fmnf9RL0gLfpBDeMRXIkZaRQw
ULXxq9mgs2jOM2KYrKKAnuK51ftpUbOaqVuNfTg9hzlwwCPY+7nYdgp2XQJdPuOM
ds6eOeT2dunhUenuN4HfJUQF+Rmk0orZNwNmaFm0cNaQAn49H0L0HDbqV0lwJJr0
d83gQS4kmG5u95G5nVLVkcq+KiHfV5dxdsb0Z+GgSezCxJT0ddxmBMgjL8eosmZ6
s/bO2fSHPaugcbAYBq4ncNyyIp4PntvMn3DBULOe0XipxT+gEd1w4Y9yYolVqg8k
0WsSkocSYI7J9plcBcdAAPEX2gg11xv5JhoPXkIYg3F6Ww8JORjoel6WTUZk4o4K
p62dHH3YjSHIrdGIXYLWhsyKVT3rqA6XiNHxyeEf20iT7qe0Vu4ph+kZO7yj7fFB
9qv0siL9jC5SLICx5FvhjAfMIH9jQnwexZvYfNztoKKTCMYfGM6OVAOKHJcRgEvC
geMyTdP+rwqs2F+WYP6/LHNXjJUrhY/Q7tA1pPUVJ+b3SQTsCSha4PBpWIsGSUqb
oiwlXNq/T67jhomnqwBLtPdPXGWTgVQ4XQ4puU4B1Xo4kPRCcEQD1piNtcR6ulBG
fKj2yGntGtJTGt8CSRX/kE9EE3jMprECdirs8Z3OKnfCT1i28x8Dj2irNJOCE8vy
E2dZceeJ4QUeKMmX+9EAZ8JpP34zkMkOM4/bXcNaJD+wdsLNroKZSlFepQQVUVSz
OuncIZbhbdslZTmlGta0g6IXHsWDa9OeaiHT1jUoSl58TDYiiQopoDNggzzJ+z6u
wGNFw24/8sQMjIsasu0ADSMnOFRHNNNoqYTaC/2l28/qmKbPDP94sYTv9R7gP40Z
F4bwH1c1fI9dmetAqUerM26CjS9nMopkseGvvD77OGpaEa/D2eAT16GGJwo5QZ16
P07etPL2K+XKW/GJW2k++Ljyv6T8q5io+AMOw54YnrXr5wVeEg0l9fdLgatwow8g
AylbVFGvUC47xaAdguPX+IfsFPc/X+ZMMMxpVviktJ3B9F9RvixLB876wi2XivHi
n72LK7xscouKCbwXs0jiPX9Ys9/4I6ZKoZjgPwagnDsfuioYyswLZbxFpbFydptt
KwoHFmODxG3UsRHHXoA+T1BsMkvFwvix+Ti89lkSgQ71OUsTCv83ryQYh43fuudC
n+TEyUlQ4brUIytBzruy9WXSXA4keHRZHN1a3m0ye9nVRwvjUgM5GXqDgrc0KqXE
XNSpk1et8UYzvR+Ggdfkxt3AeoSYWtIfmIzwd4IQT7PT9CICaed0YiD1dV0GRkUK
2Hw8yem7Z0awuunMeqmJcXRl00YV7mO+AVMlC1KjKTUHevRLysPQAcQQr+mHXuBO
hLIdgJvplR5UA/CHa8WJEkl6jft/y4icOcReO3u1lohR+T3vDHdju/7kX6hx95Ku
+RxrJ06TGcONiRzDtaDTxkLhMSE83fWnVXNAUr3eGZZWt2XDPtLVKr51nr0mhtAu
Kq2cd/tJwDz0ZMXeqrXKzPx5STJPIwuR1Bd3a2LamOQq3F2c2Mn8VPSUeLOpKG4m
GTwvrr07ANKDeVlnz0Q4nwN5NspBbWQBXLWuptK2z7bQeQEMWcD00iPQcMFyBL5j
4elMeC4x/Yc94YOKtiZu1wgGHK3P3tlOYuiYv+nlZvWlkmAy/ljJcuF8fz45L8Dk
6dSSdA9MVT5XG8EjECCFzZiRILgqVrkwRkAjpss6NJr1q9Q3dPH/j/D700b3kyJv
h4cXusWdCnHxqTUWcO3eeSIzSrnZrURvaPK2dREwXXNljz4K36CGef2YIcbs8Tyi
o4IhXEl1ZQOHtDrXFgTlEXRMZLPiAqRdW340IzAkQGNf/Po1Z8q5upXkbxSnmkhY
Zss0AI1p6G9M+Y4SV8LlXd04wNdscC73odxBTbp7KvLB3v/uSWeljheNGAhPRq95
02bR+ZOysk7zPMLapMr3HQ3aW8tHr1tG7agZIB9El5TDnGQ+Vx0yj1KDcOSbehYU
G3grk2nwOpzRFamM/DjrKW1qgXrVj4h8ZQEP/nEWTWZ+F0KR5NoOrh2N6tuEIK2+
76UAgDSVGTK7DA2utqYglpzKIAJMar20Hiy20ebvZe7iyuIOlelvcmORwKLtP+BZ
y9MzgNar2dV2vBrzy+WN9a9UOQAV8bbsEYjJDmiALrqMAgCtVd7bXbWRocm9Nfhf
xsP/y1bRc+uLnFO/wKa2IiEQP+AfbK2pihpRJwtSaTj8v3KpEsB0TEXMP9NXWhAE
8R45lquEG2W8QprJ2CwLual/EYo4nywJhXDoUo3w1YywUiphTxSQ3QoyusoKLe7G
acra9l1/A/JGVQQ4rYePkUooCzCsMELgqHR5OiDHX0nAv4YZFDU6Z37CJjNzE6iW
4ef4UfuH9SD9x4kKoJTTSVwyK2YscxseIpDikge+wjJ6Ibf/TzSKn2Qe4SnELBOV
/3RsX9v1Obn1i0rXaO4qrMQx2iZx2TbzhapZNJ0p8E5hwQOs5W8c+B5YhZikdPuH
WLEuq0J/SfV4XguUE1P+vagZPIWcEbaWnAuRdNRD3DZskGQI4GPhx4v4nReIAjCJ
2HfnMxLtfBHYmvotFChqyzqhbySASVSqFljYeBybX1ICPMJZvlVdq2U/q3kfw37I
q82tQK6hW4V6hytAcJpoFgUIgOyzY0F+HWaPKlnPKruaRiUOZOhXjeoBaBsNZ7cr
S0B7JXVbZQagU4Yss7WOE4c7RCedsm7MT/fZw6ZI4s6iO/I9Btl9cJ2vHfEIjeFJ
49gd7oAxSk8mgP39vzR4u9sL9UaZSrZhIIrsqiiYWatJbHqhRPrS7yC6bBVFsE79
1oEyepTwMFvZyNFuAOuhVL0QF+5mxkjcQOXQ8t2XlNU4dJAl185jr5u6DJ5F2L+k
4XxZ8+VOjv1sDDG6c0ITlh6o+kaZWjDG7OdD46LrDKsPLoyKFSUcpdStV7iNT+nU
7wlPxcgxu+uKHPhGb0SZOXj8T4AqE4aqu2zPiRwl55xq+HBbdyYXuIPP0ddQshHY
Fp0wEZ8a7tZLitAbuLjcnfI+ouvaBLJqNiM2dzID1I0Srg4xSaWMDo1QlO9pVjZM
TS3tAGchQNHdCafqYkRgcd2CeCuCTFwtFwm/fBpleoPjJIKpGl+08OYXyWtOvXms
SAO/DBcY+91lQQAvtccS2LnG8BpSmlfWy6itpzyu061qm/iqNvLEemJ2uCI+/8Ce
pMWu9nJ+lscjRvPaGflJsim5PLdF0mKMvIQjy1XnybEREv+2aEe7d/j1YcdmOYxB
P8VSPzvQ/1RL3PbJGSpFoi37c4XYtxACHpXFddpf9jG6/qlibZNd4I/8qdc+NIgj
qdVMnQnRf+cosbcqx3iICYkQbdH424fHzX608HJxM+vbOP4s9L60TiHnMKucv7sB
eR3W7Yfu02dB+VclwxOEsNBrMhQ9RDotcpMwFetXb66v1wIU4ppqkjp8/oC5ynW4
mdA6KpsxDQeY4k3TAyDU0Wo2u2DT+J1kgo8p1McIVsm8ZjO2DJrdpwpqs5HDUyyV
KR9zPa1xYxFwD9kpywwBKGNEkDM98pKN8nBnKxegkzEdbQkchpWbzUf3WauSvrX9
uw5hgEAeRYHUIEojp91Y7oXtbpUejH/wzael0edUlw4MHKPYC9UAVpq+fWM+vJJZ
6NEOuT3vfpfPdnok1JFAs876rPA2L2/J5IU+D10UjdvgfWiLuC89FOhM9U1Dtia/
NmRyFwq/++VUR9XR3poBMidVw0InoGCXFlSYzi201VSwy6doNiO03GZ0Dl2G3WyP
nPYE03zGkxxopUQvwdIJkL3ZRTdOhQp+Yj1lP3IRLINITOaM9hZPygVl/nclBcnu
WJFzHRqHFy6J+I3EJD2Q+8R0mj4D+MUmDB1X/5u8n4tt1++Ptyb3Byeomj5fv8s8
S/Zcowf9tyoPCLhA+KEKyHCDv6gxlITdoBoZSBBqZPL224VnuUnBIq5B8IGqBKjU
UH3NDDXzTTC5+0+QsTEw1gB7jb0ni7igHCMjqiFJIc494x0DjSjXAJ/emdyichZ1
qmR6u+EJ695VBfpZW2kPkluHo7wRFoCCg4lJ/H84D1RtCaUFau9UR5ZsTe8BdTIe
E97zOqGP+/4xp6aYBICSwrELoqmjB39OWow2LJcaguX+1l7hocoHjt5DLS/Ctn83
VBC+yVnqWGy6VtOZYWOFlsZPFaKYxrM7ovZzJGABN5m9LaZWFlgkXQcr2rksoWrO
+7MZB0G/MNRWZRrlBDehqHnrPMRjB0LovY4pReZPd/2e1uHSgWAqWFonEYweIMKI
d/N4SKApcKK77UwdpbGesKGKoBaoIUNOGpKYIKCZdPcVtSoNGA9kcA6X4fQQnbP/
q2wnNQYB4lAVFYMY5zYTjRJbrJQvyFt2YidCd9s/Fxm8hNh7Z8Mpk4Mk49fV4stp
WYZmEQGlWtN58t4FMz+N13jt0Z02SbdPc58vyht6vsCw1BTGOiN+TeJogcTcg57N
Lm2H4CX1cpoJPDhfvO/ZJFw9aY0dLmdxZQVc9LzsBwsSO5Ggb/eS1JxG1HENuQmJ
4Bu8oP0Jr06m4ByX9xMT9m0wEX14QNYRfdVPFqjqiDmHByHXEBKzfCMMUPtfjcWm
2j2oo8XAgOj1u+PetPC+w2eo0F8fd3WKW9FHS/DmNVU9W+jlXROaQBqv5BBXh6F5
CH3ig2tQHSswiO1nTRxOBUfcKv5uglf9zAGihrMHX6w1F1Rj/NmGE0amjhuj11c5
QYVuH9/w31A7/93pvaCJkByF7EhagSOs5d1Pgq2BfAenxziHFbsqFOoaCIn2X3V5
T6m3hkVlFlJap4q3IpMVnk6lAhiUw9Chlj/ucUt1Utf/qr3hDgHC0TsTWxP5s1yc
jrvXVBJTwlNU31EV9hQhT3IMCCdylH/gqRXl1DnoGBUBEDEEoIfO2aTS4VpGgNmW
uw9uus3uB4oCgXdBgQF3x/+856B99u6KyBuKE4YUvW+GMxM4R9C11++2w0uWVXUG
aR1maF2NkQKhwGKqAmAPImKtmKQ5kFZcBy/hYDGEhyTR59b2w32evcmGpfpAtUhY
uSVt/bKSFE5SMJ6MnruSXzBiTK9fZkSMn9Ows7odlmEzMsom8RZffIC9qrmz+NbF
PPUc8MaZys/IvsHk5ZVbX9lgNSmj+ihc2Z+7BmV9FQoKf6UgY03irqymhB4mYojv
UYlKi96S2cxhIbdIlSpoQ2+Eoq/qYX7LXStTYum1axVtq9JNIuKKQXvCjhwVGnn1
XJMrIwBrkxCHWlu1Hf6P+HIRJpkdCcDNzdVAUmZUcY+8kjN0k73OrUqdTcg0vCQQ
JIDvF3hzzMHLubHXL0aYk60v3LNZQgAUEColA8MVBhHACjuDLvQJMX3qGoJ2kjGs
YfclGJNnO69QDbr0x+CyrUad1fOAO12+B6/NojGRtU9g8ujObe9e0mG8WxU7IYos
Tzby5lkdMHPK9RLLMbsk9f4ekKyENCtGjCJ4lDT15+f62VQPnH0I2YwX3qXOk5gR
OHRn3oONsOtHLaTztrVVmUdvbCjCUHwK03EWhxMZcx0NdAEe2xoz/tovIhKzPpbz
UvB4ln+QtKFutxPw0Q3SdH/KxCx9wxIeSQyzfVrTO6Dfj8KZEB2phudqqVROcGGz
fNR+9U6P0dDZK76VNj2M5Q8eVGT1gCh5T04VuXoCgcbovAu2pV57Wuxe3UtZ57W+
DjR0vyBNMEX+1u3O44lQlTDzFPXOJ/qm7Fo/EV+gEnaCIxaU5L5MYL23NEPoMems
qwBw8jl5bXk+b3k52jfQRjncDx30MTOQhqeOi0zjoK4dwWm85JGAN1qfVEwa6DTY
AulUq2EFYoknZ9LkByJMhO0/NnVG9gEExu2sx3cU4hMd4RVDb+7yi+YlMbMKN777
Dt40KpwUzYrdCvrMfpKdGoeJgW07LlpIe0rM7VOyuUuDlmg++vvJfbWwX0GAnKBu
JIKqsFolqvcxVv+qZGfs0aiHFcjj7ZVLtJFJhNyezl6eJAUzO9+bI2ggyJ1CgX/q
SblZt+NopzYYvHjT6dC57s+k8JTn2yrsTpdMtyREzBUfkzdWft8RwEo8JrPhfaVK
XaNOJoPQAU0cm373uwaoqHVQCmnFWq8A3s/0cjx92zwcbTYHkVY3oQ/rWDTuCEOZ
1wFLX/G4ErLGeDfaPBdvVg/YUjx4TlDkhMW4LUDLNC8M0PweZJG0liA3KOiDxWJ0
378KnKL21KOvA8CBSpKwKELwQpGgKRlvUJfCzr6o2TsDh0OixEnQtl1+Js5nkepD
v+xvbLiKaT7DV44rRb5gNUoCyiyUSz/0/JMOpBW2tPuEXVgsBWXlCkV3WieI4Y/x
Aki9JBgNkXDZUGKB/+VOxDNt8QXxh1KC7ovl4j2GjajmL1KBIubU4aQQiyNtjiID
i4wIZUPfrWA7X7Lht9Q4a/s3ew4OI1d5TFp87VY5F33dqwLtlENPrD/T1fRzbZS3
pEIB8wKO3PBctSMcWZWLza3xyZJYr4qS7lku/UtUUT0B0W2BAm1Qvku5k7RTIm4x
q5BLjyw2wGB3zbVvFtevYB7oL7jN5dozPOtIo1cJz2mQlIwhNOb9jffezubd2aNT
iLQBhSeHwPo14bjRUIZft9MJGvvgnEu10MCVp6N7vdzkoeHFF9JYmfkrfONChPFp
RDB2W775pJwQ3wfzTrWNDAl3uDx9T98NNYCoUz8Zo9ydCI4UuHJ4pqlUo5cyxtPL
2k1tVlBXxP06bbv/4QXs7seV95ZzMNrqj+zxdLF0Pi8xYPqK8AyJSZ9kj8VD27C3
AKE8pNL2FPdKcCBgsYwjrx3omAofEj6Kbtt6s6w9ZgDJpKS63WYoGVnFSfSGm3bR
spD3T7hd77fLZvMh3J79cauJ/U3P9hAEwbfROLNHN6ZlIgnqkPeeOFmEcnbAVau1
ImJGTpb+ONtf/WCZVtoGa4j9YS4WSJ6Bk89fwpZg4gkemKiUkvs011Fw/kgdnrdH
rggzrYk+h+1Kip9u11w/drLd25+siC8cyEITSDP2R3ZIhbduR13pidYVPahGUuXg
8ZesKvB+6Gu0mv3njSwHeotmfXYUpDYULotZtN4/OPpzOeSTNxYTRlY2iRyijwaB
cHJapyVYUsLvRYo/e8pNzk/VnUYNycxHZsZnucgdnjB7YSzCHh/B6RuPm0E5/gdf
1Dr7S9o0kJCYx9JPh5TZl4FaB0QiG4wtBedgQwj7+8NCimxyul2OhyhcFsCXvfuF
WeTIYe5DzqQPBnhgy1Ze1Lb4ucgbZPKnZEfNuxpeX8seyBGpyURfRwpUBkQCIH5h
PTxBizfQLvMbtKL1EWq542YunxWSHWOu7xnNA+HCOnolA1JROMQ7SvjJOHdDxZZy
ETMPxyuguF9YS3vM76wA9gALKx5BO6OGi1/JHNPAj96RfofYFG8ic8ECfpQShtcY
aDFcb1s+Al7YT7uQ6UY8iQ/WA3mGgX9PJkICLGv3hexzkmmDpM4Ky0j0EkyxapqG
vUFqce2K3Ca8CiBPaeBtCrHqs1oPuCecwmPyKeOi+RdUEj9BKsaku7ofWhqCcUbs
1wJKyDcGvYwaNWAoo+mz6qk9e24n29dhDltofq8NzkT52VNKmkAPil28ODDPT6YV
ODDN8lW7XnTeNYrqgvLJmyXrtESuKncinpjrq7UkBbNlhxpmFA0S55EZDbaeJaMP
OetbiqspNyXDObt30tj3L7Y2v6sIIoOBSUb2D+9dMxETLAi8G6rS5HuLG6vISF/Y
NODzvT0Yc/hbU5Ga1M+cEkdRXJIBCfZ0by30vEY5v5HZYf2ab6cLgWwMwFK9ltU3
3BPZ6kpfNMf4gI62SJWG2+2p5sZpub5IogMOZRLOJMKvQ3Dyjpa5jGhboM6UeOa1
oid8VdJIdvQSR4nq8G7akA9oJLU4toiue5ejwq65sdre5dnMqft77wk9TsAMTvka
ow3brXCbPsvM1TP7l1uJyaTXIS4CnyPSghvsJjYowiWf3XocVuEQCyDk+5ZCi8Xy
tNn56b+QyXVY50Xl6QuQ9m6GAnPSlf73eV3qAslO9nFDJAyo1TiogOYNVFQhNSJ7
SaY8572U/+7okR4BOvs7yy0Xw74n52SCed0bL5T1hzQdyG5PfUJJs5w1zRYIDRZD
YiyFL1u2Swxl7WK2iso/jO9W3BaXAabgwmJvz6KTeC6MZ5CklBnXE83/3iXxuhNp
C5G/cLZdVKwweHO5JeZQARZuKVKEY5yud3UVyOh4q4BdD/zsRP/9XZQNn64h8eS/
ps2Cetabj9RSX0Ud04LxvrjNNeVr8YpHsurStvwAMv6z6Sb91jUuP3G4DVNSZwgz
WLct/WyzVFjC4RKh5PxIUOt8gk3Yyogx7LvyiL+bd0eJRib2/xA1LFtIbgiIn+x/
lfTYI5GdGckGv+DAEa4Nc6RY95ZcSeg0jdCejnX+H9+8immGkxbGpTNqBNEPVqKK
LS6ub3AmIMe+xg43XKn7JOQGQoxD8hXhgUgkLPYrCATuAHycL4DsiHvlNkXxj1Jw
xpFdvFi3akaapaNy8GFUima26uWWptYR5Ng64UXYKpyExIlKR5ePvOYja91rOSiz
Edk8A0EsW+HbcZxS/nfebx+9146yVQaqk6heyYlj7cF/lPKEg3qYxL2sywariKRd
xkNwTlgoFKgZw/LdxsToI7pHC4ku4Get47LOuaNA8TfOyw93YC/UzeKI/N3zRDke
tcZPoj0aC/6EVhnIaNChMFdFRlbWo/bNC7bYq2lh5huihQtV8ooS6M4MLErP/Meq
2hZTuulyBqGDXRplPp6zxJXsPEN1/CRcCO/b/m9TdSu0rhqYxeoQuHc594pPIbAA
ZsiZHt0HlZk3Ikp47EzEIZUFg2fYlvKcKkA/DFYoEXx1aT1uuX+YjzcypD2MIpJ6
Om3n+QxurN+KQxfR5u5J2pW7NY4KWxLZRVl++j1tmt2sERpqmfYkN5SxMZ/MyqXi
3c0fj/mFHvO5kApjQD88gmWpPpAVcOTrp2GMU4wI0Jn9kyrexgDZCZELThCtvD4Q
09iPgjVqWHMQNb0WNY9bPMjHE/N7XF0un9nDM3kskLT0FLBMIIRZlnjUw/0kuA6W
UfL8G+HlZb2VRwqRz6q4+bDnVKaqRG/g+XWLA43bnW85oOUtbkM08GyDwldkDio6
DmDI/voQe8AP0rrEEfKUK5BAvTxtjGHWmP2l8X2jf7HtS1T+WcJQ9B/lTvH25vzo
AFI6P+XyNfNCfg45ULIhu09s2pqTPyqjOl8US/eWmQrukxvKsl61p1VJiw7B7plF
/DLPT62T6lj8tWvBYggk2z032M+2YCIwu3m3OvhJkKktdLVr/k1qTASuqw+sidgV
5lP6e4D2ip+FKOKrh5epCR+KEDLCZSRsg049jJuocCfvHpFvg9mNtXQhw0Z55XG6
BdfLO57TKMu/oPJZDl0PCZCvhSinUnnJBGtLZ7Rt2j7VwI3INocHQIuv9yIN5SKB
qfM+U3J6gYk3d3NmZr7rALsOQDgxM+iQBWk+i64/x7qFFA5SNFxoYEewrmULroJ1
8hqYbt5mq6cN+hIY22FKnZhqZT7RhmFMSdESzY5UIuktqfDyJv690BYi8lMoQcFy
jSOvCHBmUEniV1BYiYZ7cthIE0WbO9Oj488pLoIKFDnLCE9rQMAboy4iIGl8Qj+f
JKORXHSvCGJVcGD9GTAg9vgTeto+jNR5eOkKb7g2mnXOzWXUeRpZYXD+dgEE9A57
LNQ2C5+4Q/gKvlbULZili1Vy3XAFPIvJgXYP5ZKHzBkupucvcqS6fyUr10UU/MxP
An39UYtkKZoiGfV5gT5WRQCyPj8wryYihUHNyDuMeV+PirvRdV/BTL68lGhQkDrc
BKOn3uDqqHhwfjw1cF+ywHIhi8cnL1SIxoO88tCTmLRlzsGSbQVzO47RVyt6mCC/
lHVJct2QZEfQqu3EMmXTuGuALpZGbPnkRQEDWI6IgWPFAo+vlnJZ+HRu+oN95d59
MzN07PWFCWHx0l/ZcQhroRiUACaef70gOEIYf60oqTJJQxxZNhKgYS0abY2xzYT3
/mEKCB5P2WYarZx2nZTRXHEtPPoiyrjNqsaJEcOjVOZNywf5c/tBt8859vH5Xf4X
bZeg8MLaSL4E56Kw8cf0nT0PkrchMaQtEoFyFCUu95U144jx91Syyu+mohLs5N7L
s8bFoVmg13H304RJAtm8RJpZ6U+Cjl3Tl42OnoPevFmG10LOq7y8eaS3Us5aIcDN
gkQwNkTzgJlgpHSwfIiSD1Dr4cyGTw9Y8Q5+UR5t2Rx0/xEImL4Ccn/QGubOzzvq
tMPRFobDnov0YC/rk0tHieckPwyhfLJrF9xW4/FLt5RbP+g3wVgRwH1WJumTTI75
q3/0bM7nh9Na0gER08WkWCwynDUyxXK1dtHXtemxFNFt8UbKtLDF3ehC3IYHi3qD
P5eLXyqGQmsi2dmDxP9Rx4wk84yuSRx/DWcblREdDEivnPS4YWMWpZ/CRm+Ox3FK
6oT0uF/LGGs2Q90zS+zGXa6pm3+BXF7iGJSUcl06xRuo9Cfi/lW2JvlvzinVydcf
cxOVNq1R1R+7mnehm4cNQ3AMn3lqGEQJGjgQcwuaYLvg/BJ71k0e1QQbQeGVxLfG
JaJvag9b2kCeKx+EH7GYVVK2ucv6WmvIiLAg6rOMosPNfYFqcN8nE+3ctK3zmsFl
dfIyWFyYSPepInJUtxF7/sifIoxstRKzxzBdxZIip14EhY4FfRGpnrZL6fPJQY19
IzCifzZ9VywuGpSHk7wAr1513y6jL4R3V/F+0VWJWZPREYW+W83+zvzzEsjB4fdv
fSA37xMoqqEhX57D1oJmdmKMRe+WusWqWdaFGdzO4rEIh/RmHlMQjnDRChhqWAe9
R09NFqytqE8UuS1Zf+iagKzqRYyLsM4VDrFYZBdDb/+fPxKG3NmNuQt6YyGaPiF/
wNFBVuicNkO3YZGc2AUZ0Zd31BiCwThUUbbFBnHjf8nFQxzL+8IwfRGaMKmky59c
qVPB4ej3f0um87azGsnzmyXM2/eXZThZzd6fNuYriPbOJAm0i4ZXrqtlE2dxLcHT
dYZq96mhh+FmCA1NMJSr5UqZOc7fNXOm56urddtPgVxp8l7QumaTI6KoIUl7vtNb
bMMKwkuFF4wqZ0qDn2lvBpKj5eVmqey+LVPL1omzg+KbKQcNmlmS7Erj4qu+DEyF
Kq/PJM9VQmH2jjgbBD40Lk/wvRdjG9xz8yOxTTtLFDpj5cog4ameO2UIR9JIyDMQ
t8pkuG6NxJ7Fk+9vfld11e0Lh/ixBtbnTQaEPJYuNuE5MmXwCH7Qgn6RvqubHBlh
V9ZjruYJkAhgFMjhiC1Utc0V6KvAbZtKF+3N4uxY+/Jw3+YYxavNZqxpl3JaqHMg
NEEP7htnyWDSOxbVCoKnuNQZoT2JNCBcBRUr7oeFUggSis6VfsFvU56FYG/lq8IG
tHPGm4wM1flanKdrU74qHUSW4fgvfVkszSdTs5zUaOr7ngf7GKIKHM2zrOm6az1q
VrjgTOw/AX8shpq7uHW9oh38ZeFHi+JzpmPE4CNbAlvU7HEhkWpmeHb9CM6vg4ym
4lQhdKunb1oqtuK5t2UdjhxvAz8WgSMMeNbtr3PvgXfFBBRJzbI6hdfKn16auGaP
vQkOjImuB56RqXPIPmWT1VpU/w3AL+jKVdYLT8/POMf6Qbyf5qRwZBewcxDcJJSc
26PVulbfxbRaDudzXU7l+ybVpxNfFosfD2fWvCDfgAVwnNmLXf30U/VQTfa0+ImC
2yiYSPYWrHu1aWaQvrXxMeE1RqAgJj40iX03nSiMUbW8qKJA9Np3TcNp1iCV7kYS
kGfAs3UAY1KcGyVfjQn5978lV4BQ2q6kF2Dm1swjyN3Gkjbtm6s4uIUOATv/zeRV
nIn3Rj6klHPyAjKaU5+HsSDdfkQfXst+BCJQq+q18Qu6/rEQbK+P//BvxXwCWvSy
qS/Jx5Wh4qTzNSlCXdnZwosHY6Xyqtr6dZqPE4PLLvYmKhD5x2TEBN2CCCDeH+QF
0Lk2AZ2pI2vMPRD0/zn1rBAIbJqdQAqSjysmrb9uSJ4txjV69CVVz7/W5hU7jl9N
ShZs2Dqku6fOlL22QMuhX+j/QwQB9ybW2pMfma+ZLdflm//jlEu0KWthaXFKLVUh
+4WMuU6KSA/+RTZLTlTgv+r+n2/o/i+uycVj9QLsWeGnCRYHqZwuzgvsspHMUKSj
k4bb0b6SquUB+RYKuzkcyZxrJzRuXHJeGRrJ39jdnix2lRXzHfHBqLMRaLWYDqKB
tFNmPkx71im+2GiJ/YTc/5/VEQDFRqNw4a/tFR6wQ9fTy44GkOXWmD5Wh26HpS3K
/FufSqsAVchxALWYQKztkQKyBUGAGowGsmQJEO02YPi0cIJDFgssH8J81hrFfwv/
dx47I1YHFmjsUdop1dHembVmbPtlI8LmQspgBCRaoS3htnoxEkw+rJvm+RrlI/0c
eNYnnlT3c/eIVz5czvhogecyHJsm710/4ZTbm8D9/FcBgTX+M9kBHaGg0rP8wPIK
DHdW08Ny6Ybf+svtyD01azknJM/RTubNGqnw5YB2zsoKrtxadmi30/JESLtwj07e
mEUOpCHYndC42HxqdrD4JJsP5vG2kvV0POcvYsp6OKKlsk0ArLjJBs1cUzTPegzw
meXWrkm2TNuwxhFYLGcRNHgSiPzMChpbBsOr6BQXd2KxhcJWNfJQiTZ6eINvsuYh
Qeog7ffgnoflnR56403qhWRps3ZhD8hGFuc2S8WZgKO5M3Zz8CXNcw16z+nhYztp
DSsCz709NSGDGokP1Pcz4n/IdmQQTB66AEbwkPmeHqeHoEVsLCjvAL4KeP/Fj+Lv
Dktpe1XGYj10B5iQUdHf+nSNRZW9tx1RtzGhGZRHCAfOojOpstwWpO3dWDKSPNtj
bxiMO5ZAH5z0lH5VfE0+Meq3D7bYRhWsTCD1o76v3kvU6inpCjLY+LlLtBP1ucU4
R8ogCLF2ZlAFJjhydT1CKsS5V6OYackYfj1Z2N6A5yLaAkXouYJFH54ZDmITdBZK
0aUa25vZ4dga8TyUlFv3YR091FNNpsnINhMsbqySqSc75fZSV2U54ZP/ZT00MAu3
nEsKN1/cAiYdJ+OSn3bNRNKchBIMthtk6ZhiW938+fJQNq6si/uXidvKUziio1Hw
RB3z+r7K0HJtb9VqTRDrLXctzTqI2n7XmHO6JcSl/4wbOZ88CnHckjnorrT9dXe7
bUN5pM7/qa+DllyFkalbKx6OhNy4/y9JM3+MURMUJ1sLFgkibSR4RjkptH9HVPQl
Un+4USqg1J91XM437g4/JHSyMipXk7jptyFDJGa/XJZRr2fCy1NHzxpUheh7FkjI
DLe6GOp6LZG2I+gfbwF/QXqRXMkmZ9hiH+YdSL2uo97k9OVVyvv357dbhRIPEZvb
GSYLsoQuMrz0FlcafgmYFfCFI3QLWgo64th17B8eU+UWvPv1E3TksMhT/i7VgD5t
Mx5tQtEUIMA/OiBqziaIOgoYqjzpl+TfxTbpzc97drqy4zz2l/HhfRDvK5XQHHlc
ODlrVg4cCVMfg6cQcxj291fJOhzAa4HpEB/auo7Ov1L1db6+ZKjFwpOOiTXXRSGB
H87xEiZb2lyeZB/5VgKEuEghKb/bwaZ6l0G4XK97x0HTJ9uz1th/tuW6xonWd3+T
k/aEcSfHuwHpDfg4Zc2Cr0qoC6B5apxP/WVzi0mbhHupywZxi7Kd0LTfaI5d8Zl5
3ZkD9n0YC7L944TPdqhmwZeJ22VH6+6qA9rjoU5nHFWDQ1sKpkLIjmMeArsEaqN9
wbSp280UuTSx1adqtnC5kXuc3JpI1yW5ZCzGsKKIt4NS81UhlaR8PPEAKcegQrYJ
QWTEUDivSlMjlP6J9tKpfZ0RTrwJQcY2Y9rvlp9wHxqhJ90cu5BwDyHrR/TlY5Lk
L6YP2V1GO4PbjW+7fCDp2QzNxW05AKJay9aDfS6/VMnAbGuFDXhvRfK3MSjja/OZ
sQ+1wuytDWxMQ9s3jSgCCxUzI9zKx8Y74lqoHaQSQgvn1wf+/13pCMV6Q3a7ObKd
TQ6b23hXa1AUNV4qurV+pacrRtszUa1fVr214c4FxuZ6GbeJ/WsrhjF4DJykXyhq
TzxF/dsw3jkZEQwsv1kQ3its2hdXHKO5KmU/3hThmvWXYMAgF3ta51fy0EqJPZR4
d9FsX8S79rKuAjpTlG5RkpIypp1ameff8SvEpxYRt7HZ9s+WE8ehjl2z9gnpTev6
VL17zinPgUvbPU9emWQFPnXN0CCcmW+P9KyiNWSTHtA5iTBn+I0qay3VngxI+S2Z
SIKHA836XxOjpMA4nJPJRFFVKDGv7QTaWwd48EPwkx2yq6hgLk1/RYfW4wOxvVUk
7sS17GCxtdvhj7Qq/yzC/d3URKa8VNp0BVYfwyBlF4iMm/10qcArl3ZLc30DrVD0
feid87Yt3aQh/C+7AZFQH7DrRsf2Hv1rSGllxe35l0l5cbNjsnQA36+OXOZQD90H
OEs35aweJfovzwmOHywHBuP+EKXI2WcYHkaT5v5V/aA0Ko6f108Swul6mJFa3Xx9
DClcvvvE6lMxEevrwkLOACNwOhWP/tPJLYV5+SK3pTwDrY3Gss2xXjTdBkq4eTOo
h+hwo+VT4/f7OmtKQsk7cgsPe6Bh58KRt/zfyJHvOSvZu4+if1SFD0cioDSZvQVg
DKP+ua/ju1pTXJMKCj5Oon4DnrHtTMisGXBHbJxNvM7VMyeHjItzZO1vsQTdM0Y9
0c0fDrDwXwGt1/Ft5gslcrEMGLVM5DKwcPLaFthiVgdIOeyIzI2pfi8OTREDRNC+
5W4lTud5cEsmlvbMv8/xtuUj7R3JQO9b04b/TWTp5hucA/jcHQpkDHwRRLzR1XIm
Teg4hudNU0p09f39uz6m4TlM+NJk++1f8UHDFJd0FtIH850XQBchiq1CM7q8MkHu
6QpPgVHx2jTPo8CpGFwYfwnnXooNDAmKSCPt30hVKyO/VSSJEWoCbNC60o6AxLER
kjtz3AwL+VgE561gb7FKVXCQiZjtARYRLo97srm1NueUay4xeQ8KilCZwyHbP4UC
HTtuOg6gXSRjLDQCxw8lU3C3i1twN50sfv8ziv8uKm3xSV35gWTQxhWaTwG/m6nB
oLFryTbj5WgsZYiWofrJjQq/fgTo9o+aBTU2t6dQ9X51GgzFHgQtr3iGOL3GnF1n
zTv8Hyo/c70LiJU7jpLELrIJsROA0Nrzo186hKeRPJQ4tvzUlgrd9pjhse2F2wYd
ZezLHuJ4pF1wHTrU8vmDq45buhpFz/ddrGdmnUJt4x+I303mnHCz7j9wuzRyWlTN
6XeQjjEDF9RwaDpf4I7xrISk/TyLIn9B7X8PFrFR0m/DoGhl4DDBZhHt1TyOGv21
SVP9iMP1l7RvBe9G7vbZ+5KqEIRZs/5cJIY59EIVUZxyvGQwhbk+95Tkh2b+V3dY
KzptYfqHVyJbUwnVRiU1DTHo03ZYsTyMknNMgDH+2YApigiv6h8EEJbdBEzQJnWy
GCDXrU4zaV4NbwpjMre54r1hTM1Uordv+goRx716xqe/25jDN+ez0Ok4ekhRpImJ
qepJNSLcHt5oJEa1BMWW0i8tApLXeEEtkbF1O/0r5Mt02KNH6i1Z8Mu+pldf193R
BGh3hwGvT0ui6J2Qkt48z2jvLuhPSzprHBUkfKSpe8+evrXklGThL7uAO4xyLxwB
F02MhmRQPc2dg8R5e/LVHmvcq1PzUF3/i+92j7YeSDD7PYt01L/8jYNjF4BbxIzR
qfyuC6ErQV3n/XXlOu7EEd1nksNwS45dD5aQRaI0GIsiFtn7w/Jd5WKl1sm8vQd1
4RE/qNMs13KOSCuqB8DDzIE2MKLQuXzNKe/rTCG6ezJCij9lfm9yK9wQcC7mV01F
J7Pl2wy2KCSNbZV0mnO0xDcMKefPUEHUYL22LtRi9FykE+vSkFsJLNGiI9uWbsPH
QGnZGRgrzjPl2dfRATUneLBaRMXwJcooBeu3PANKxBXmZNKGjMM87kECerEu+Ptz
/7EQj5jtzlIHRQRK8VcNWuqyYYahPqRy8kNmzlUd2fNAyItfzGmS0rHlhAiJm3M0
T6WQPqDz2jRuMcSW6zugzOEPJT9GXBzOIdxu3fn5dwUOSGV669iJSwmRLCY7nlLB
Lzfx+GWojIZe+S1Z0AyiTth5sbLjwe/5tOoCI18zQZuWCMxLhXW2LmLtN0LMUTnD
C3skzFQ7FRcxifXsGQD4tpr/4kW3u00Rs5q0KaBT8V3GL6boRcwuGvmOPoq8HAl1
5z5fRgCMPkWOjnPWTnEOT/6BZtH4nJ/EUoXy322u95zvaAYtKSde7QwnOQRq9wul
WK+ca5fMlzBBeMGG31v2XXrJIaOCd4L1N3D+JszWUNqUL6pGnD/78bQK3fQBwO+U
cjfv57e14fjx/EjnwDh49ZztVXZ/7wKu6bvuDUqFYlN47WQUBal2LeOzZgm/hgF/
QDlKHzQWke75/3qUWji4vQf0gPyhsE7tbH/GNJ4AMSz0UR/3O8IXXpeBEgBAtKVI
bAOFnaPkMuP3XQX/w4wlx6UM7uKN3PvewFnlHBHReFDkoi+kohmSgRI/MeehvSIe
/7Tb+U4KMagzSPgreRT7JGPCY1P/O1y+8oS+f4Z3iwDI/f4DE+IwSSb6pULI3Y5A
dSu2Plcv4IBC57YBjivktTYujEaRDyCfxRSSM/OHiYX1iWzHcGgDTvD8Rz4Md4ML
Ijlpx06MA9fAdWBKH6Cw7ni27B8pRez2ai6fmDYxvVfO4xtZzgpoDAIIpXTGkzwt
gZU1v/2DO2f/GQRbHqKK+LxfCTb2hZC/P/2/yIlcjVf/rEdkB0DEWCkF/tgpOckg
J4SfmkyAAACQBWiKjMLM2crTkRhmO6Ke8Eikbik5T4wQdrbAvmBMoNTd9TFgQ/Kb
VVAfdI9RTcyV8rvGrxTLtDLxwIFsQv3+qaRAfNQ8nPa/6ADLfPb2Nwz/+Lq++SUu
UpIo6nEYAGWVuEs8eC7aVqGtJJ5rEvsA3nkaf6IGMweX9DGjDvlJtbhrD3HlfO1h
GSrI+FbbSpwHz6QezvaM3+8cX/8BcIOCcQktqbz7LQppGcS2dq0wid925+BA1lW9
IEtsfnA+SL0DHT936Qal0BvARbGCAc/x5PFEdefkcQWkBcND7x/dRbTjGgBKF8OB
L+8XiMsjHIMA0G2mzoA8SC1297ZiAIF6ByiW7N3Gfsfim9Ie5c0uYdOH5hmGcMC7
iqWYW/aYbityt+LBmLqtQ/hbF1OiCLrJ4YRPtiRPu3uVhO72F68yM0FHuWA3mKSy
wU6t6eWjKFNvfHvtJdfjOEjsNKEGYD0kNnmMZaYBJuOXkzjRGP4ZOdz3OF3KQYS+
BYnA1ap/wAM8mioFQ1LAQuNnscgYlOEOP2H3vue6Yz8F6hc8rF9i9i1SbTH79MyW
4/xJ9hA/sr2K2Nsne3OHF8SGDes82J7Bpd2RVP7A0IowYMm1ZgexshXVk8+gtdWC
WTZ7n6LFT/V6wU5xomBGSp2YKBKyQDtqOmJHr5xz4bEv17DgKxWVUrwmqu7oL9k8
QMX1zX9J7sJoQNGMKaQAhhde9/PDsSNMKeXw9zVeInKxeROZN+fnechbRqrEy3/v
xtSYBjwAzrGaQQwrD9ffjoSESwri2F71v1vF+Fj3rycrR4G8mlf0/AqphvBBkHaX
IBBJgTfxbG4PqAYuwJnQdhWkDvtSQtUJiOtrnR09Fv3OrbjbjuAbMCfP3ZfA/t0J
EG7zXXa+EgoMZPHk3fc6LPXrxdN6zT86q8vGXfLmmosbPUcWKh5KF+9nSkUlfygq
fc+ZKEMcCVvf3jPZYfr3RdkFCoKKA50m9mEr8H6g35QHMM2QP7sVNSMz35Vj7uOb
IWt6KDxiB2dov2tdmskrl/v2Xu+rBLP8dFTCP2e5V0MwYVJnRWTpOH4Nh0FDiPe/
dyPt8r+Du2/VdinntU6SLTnf6RHmt72gjH0/8SpfxirnRdUq/IeUqBd2d3scFb2t
iFCFYsMPBnH/QyVXwhX+33FxwUhjCz9h7tn6dm4TPD6aam+DB/YbLrXdxLNowyCW
iy9XBUpT1zir00t48jRV30uu/aluOcmZ3TPo2pCENr5RhQySfFJ3wfuxnAoOQlL/
YhQ+512gFRrlg1/hBgDIvyQSJZOpdcaBK6KLPdzZ6cvSPhw45VsREkXWBS6qray5
Lk+AYMLZxzEEs1AjwQSQdA1+5Q6ENs5cFFcRqvjOlFo0T1PghNhI2y9/MR+F/aDm
iGIwdv1wgP7VueasSu59R6e29U1oukOjJ7bLRsWam3OVMl7dmy1j1m5XRz5Bi/Jj
eefFgSrKtK/7gaJyS36ZN6evRkYL/P7m2YGsMrUxRlbAOdVCxzd5e7acvjsnNiQd
8vlSTtaQ8Kda/KLjA4CNePr5OSQNgkjazd7svwT178XWqdOJHP0+AWa04Yx2zE0J
jqMknd4Q/cVLheDC1Qitix6IbsSSZmYzOO5Xi656oPysV+l1M5zG/ZWoh+iyGd4D
3Slru1rFpMR57g2pPJ3Zoh9BoEK6JBiDK36qhyoHyV9aTmN8I2qEJAI5FdnOXU+x
FlkVGQa+yRk+u2c4Wp9MGy+POqnIkl8RWG60Xv0po0dvu/tdxVnbTVwyNFYyFSFE
vISs+30lgY5FGKnJNV+XUbGvkrrGn5tGUJDy1/xXk7rEB4JIZpFOj0xuCRZzAyDh
hbq+xxoddSRKGkpjLOEJ0muErEz+3UWXqilo3xXCahXxFgJrQQ/Lcp3WpgEBb5/E
IZ8OpC+YvaaxtlgV8WuLUmN0RhbV3i8N0ry+2r/uyoNHZIJZo+LnpcQ1INlb1+W6
K8EVc936gLuWT5Bgf/81odB9tXInvGkzXJPKInwalhcjeCMjce3FWoAm5DVA+9IY
zlrOEQd8GnsAvtaVQHgTtENukyVAHV9PG48OJ11fB9mXVkSIV9ozd+N00UfvxvKi
9AW1oAnSprTm8eC76RzwNx+KfeBeouFzqPdiXxHkNjQJJuu5rzSx+5iv32YQbag1
VG1YDmdcozj6PQ7ANqNAkvP+LQa1B8PBPX8AzqwLDaCi5lqdO8cWsqOD06dZ5ax/
8nRaM6IiguoPte4SqZj7Nasu4nS07Kny6na3dy9fGj80uZ3f5cOtxOEQUPQfB825
fYrbXYvXl/Tld46R839+9WxzpoFuYM+lrOve6G0ITqw3lPZbqoGqoLRMvLceIUR3
TvV/7kNfLyKYJ/nIWDXP4guz7YjWkzucapyM5g5b0786o+B2NbLtcwK0H4JkBDF3
80zZztmVb/ObJP5IhOlX/r7ZZdu2aQeYGVapsob6qP5tU45eSsWTH7rTnYW/P2Eo
kWaQF8bGWbbJ3SiIbsHompmg+QzhqMWpglkcGlr8dEoGUAaagzoM6e5daRqVYl8L
irstncf6iqGqBtKRbohAKiE8Ll/tRvTLllZVLEIcogsGDulD7ZTAGiImeCfXP6cd
qaeaclB0YojiW4677ypnZNmwDwl/3NUf1eeyJorF3amNC3shl1M9+KubzgtutNIY
90kc7mlZeXX7gRGVSPFi2kyRP/5haBBMZIYb4amar0+BBGs9PZm7VReR1puAfeNT
DSPXn9q8gu3RJaEpCuDRKAzv/cYT/jEg1ZzipkhfBItRkFNA7Kc1Oqw9fLkgy7L8
SNdod/xoScr17YxZfkMPmHTFGrjndsoPtyHDalvio17xHi6pgKAw1K1EQGaGkPCd
fUs+KPEgTCbHjc7q+WqrAiY8EKnvqbBpXvtkTbqD0E6lMTCHHANnhjmnZkq1ZEvv
OMH5+tk+eJ0rSQDiEyEs3y5F09GM+V3HRE5E/DhJ0EceIoe8TnE2Hv7T9vtMcwd3
U590JRGyrknek57l5vL7KuQqT8gJ/v556Sg2gaI+zVDmun/jTYJAWziHt9Kga8sP
oChq4i1i7sb1hqQx7MHQbiH4viJ33ye0hyHoBznGPvmTmqWo7sXdhZbdTa8ckgLz
5O7Uln/Cz7HLSDqV2elci7AeL3psEyXCTShP1zsx+0PbhMgn8SffBWteD6/obJW5
MTttC2oC0RATdgcWafEkVpKcANhE1p8Ncql3Y9q3vXZVogBSggk0B3KX6CoBpK4b
1E2KnelDKXrE4P1wFVH1qZEa9EcLXayNgCNDpbRBes6R87EbNaGqcUCd3kZ7NHKe
Xiasz8Nuz4ziCZGbhPDkSrPxxi+4WHkbCtgnfYgZgt7ZxjT/jimOvUmAfHF8o517
phsUGrUr8kutx2gI//ZIv9O8F+pbRcwiju20seSNWDDXQBNihnYeYfWKiDbc4mGL
brOX/E7Q3X45H63votAme4DVGI5n0Z8z+ErVNEBMlQXup+dNNC2pjyVePGMGCfKv
zP5izfSGmLKnoFprX//jLWck1SWN4GawVFqqorESc5KEn84dDHfyh+5nefPHEmER
lIcS7CYPm5bKKX9hcTmCVAUJ61llbc5bNTkzr5DTuTKCt7gwZOF3lRHRE+hnAyKA
lkvLbxHYLxRh2ZaLbuqT/oVzVY6eAszbQXfLKXeP3RYnoczxUwMy9xg0cu3BaL+D
9/hd4YfyBRooooRXwnKyLjkzkN/dXYnQ3ygvFBrOHl45aOvgUvwq0OOiKxIe3EYU
08DZUafFLJheL9+uIE23/48uukyyJWdgpR4nRnD2ehzrM1VXueHhxGhTQzXh95bY
ThYXSEuMjavQ7La4n4TIAh6ncpq6FhDbhp7/0MOUCC5ZyZsRizNhtBrSY6Z5qIZC
lxO0Ip1y0k0T5KbWRH0LpLROveteZqLMf0x8jeBgkuMJKeuGwUybMQmmKETJhQ3A
c/OZLWuJsyYb8R2Tk9ugNRqPikVcLItZ5C+kPDC00FXa1fb/W/iowsECz2pey55B
5MJS93VWUmS5kO7LV7INNvn5oRYuY9xHOaJdTeIWzc7GvDY7d9G5flM35H1KluSs
+5hdco9xPWLzsM8TeMdf1ctz5tK4L/oemk6VZvZQ3Gsw/vzkGWPcHQg8IwJqeJrq
Jpx4iaCd0EhmkljygsDOB5iZpCLMYFewb/DJuyrvXvmMoYdZrDbBr2Z+yhJd5cMD
lKFqHUIensBRA512mrgetzU17fneGyrTkEeTMd7e1Y67sHdWOmmj9CuCbM5b902x
0b1GIZ79fXY1Hx8KIPd+yILnXGKi4Ynefntq2w+iGoS0HwQu4bBOMPWz9f5MX+ct
zNcZImFHD3YpmFklhtpEdP5oTQPFnZAUtcKNB+46klW5OWsmz4WiSF8isNEcw39M
WXV00BipXy0hPLXauvJooDECe+7PyHG/zP5Na3HKLW0WcfG4Vyxy+cUmovDEnORV
Rt84MchZOJNUui9P+zDvli0teDbpPcHV5m2LDS82yWKM3Q6gkbLzzN7VXGEEY2RX
MHkXK+6jpLE98SqwtBWGELqGAwpr9UK6YBl8Yimk2pPjg8kFGLuFM06c5eeLLZBG
u25UsKBdfJvaViYr8KAhn1DNLu/xFd6AAiDroWlz5TsVlMUddJS0Eirbru5kVQNL
1V3tYy8ae7TZ/AwOGIHyQAl58bHYA0U7s6kQdQInwqMTVJYOZKIUWb5yn4L/UdDA
3u9Rogbgwce/UiR+qW3IwDc5XVrSaUqnL2gXce0Bi/6UqQb25rcasqZTeAczp97H
u76ntdDSFgeR8E2g+iU3RXAMcj8rYbTWPeFEPX6dPPVd0tft6ngKLgnW8qMh0Z6y
NxWCIm24KMEikDYMw0u+uNnaLwH+TSJoa74vaytQjjLue+zOSaIBnklevm8AgtnT
gMTtBoChgd2FfxJXqdTF9lxwBGnTYSBpqYTxDJ/OhQTSM07tYSHqDzUUSKiOi5e1
Vq5IenqSWuIhQPCrmz6CrQf2mgb45DAUIvy3XM5alldZFWFS02ChiVwmYmTfI8Cm
TR81DX5tWplhynUVqrxiF+NGskYyZvh1CazTD0AhKY2IeMv6+ljXF6W991+uwapQ
Is5lfwxhOpHXhJi2GLr3JOXWRF7JgIEzdsuj2XIGZe0OYOR3g/TvLSxtStKcjbPX
OV1ZO0qqsN9gJYPZ4WmD9aZG9z1YIOGFDCvF5BLwAMN8bH6UigcVwkrhznHyG/Vz
fP12HRkHpnAdSvSCUXG6wS4TQOSEjzBdasY4u+BykEXVmfhzNi50sNFozeNMbhRh
koP2Y5qDJhcUJfTO/H+gQC/YJnRrwTY94caQ1Tie9666fxinBBmQzRZUqYL4O2mt
3ioXDvsmmWcc64aTz99tw5HsNxaWk+Q7jF4SAVjJmWeJ9FD/9nfgWMdNwqXx7hQF
DytlUDs+G7HbiPWOsDNdqaDkNbhtTWnfqw0OXa+bqCcry0KDJRlyr9mNPrJkwVVu
NU27ZycptRmHkFVPV+HYFMegD0Yg036U0rzTaXIBKKzhFI/I0KVZXLWj4vEscHBC
+48tj15w1qSMO2fVnQyITX3PpUuxnYwKGujbMJEMSQyedvUM9XwlH4Lam2L5rLgl
1iVE6uNHkHJMEDxI3QB7iyBxcdDQEPJ9SRFKMS8ILdjW/jdszgFI3YxciAOg4VS5
DF9zURe3LAQLNzt8olJgTVPgDJvniD77eMNGYNk7sKgUleKiqzShLGFIFp2b08OJ
IEHrjL1q5YFOYwDhr1qs7Kh5S0YDybsjYsF8P8YXdrko8Oy7VTZGfrWytBTQXbW7
IrMy7jkwqCAcN9b+cFYtC0ilUFOhSsBCJ0kG25rxqqxZ+8GPfuaoba5AabG5bBM0
I7xFK2+R+3g+w2jobHjVtFlv6z7zWJC6a+Al+200TFtuATls7EBGwfhjxydLBgpa
+MQTZow5zUn3aFlyfTo3K6t/IuUcgwcQmySAUNzRIB0X9jRZtshrybeh84pBYFls
QaNqLKpZ4VLfUBS+srkRSCk9jkD93MO00YchYlctnciQhNtgHQ/+EE+VdwmAZUjw
XaagP8WfW0ufGKhbAGRosBR7T0UFU10FcJ665Srh/mg/6BQPzuv2aXeE9LssGIxn
nbZdJJfXGqfIsDk/NRxlkKYbFcbFehuPP8etHMje8BwQJj/uE39TvaZBLq3/fyuR
wms3GWfUgxKQimdVKcApvCOcEIv1LTmbgsP45Lnyz0+GbCMsVTUzQnzI+mHn0zTZ
tw8Fk6KKKYWuVUni8CFM+fElXFxpdDDyhjOhngi5Nwsh+OlLFt+yKYokFa1aoBbZ
21EcG9QE2vYw8Q7iMqhUFzHcgGYxJOkb1IqRHn04fOtW81hxw6rymka5aygsAXZc
IivfCwr3i1VcOohWY9Q/GAIsJfQSGxlpVAeCihaaQzO6zUAkLwDgbv3Yf4vDPHvJ
hHtMQC4CYq9vx4k2HABgOLmEakqx+NcMm7fQQoUMNL+GUDVJWRPTU1GDVtKJcm8P
2+veMF9fQgHFqe6Y3v0y+DraWlfjuhDCRI8gGUbDB9qZOZOMpaGAlJqZVB5vDcG2
dGWrnCAX9QmMi9oayQ5OZApDA8/aLumrv9eg4TDonz+jzGG9CoRDsL73hXb9pgZU
L7hSug1mHPyVp91e1eZoA+CIeDRkNp0xQJ3gTmIg2EJeWNpUSCsrAv5Mvg8oZ3Gm
bAWMy/yCNKsguNbNywCL1kwb7ZKDyuXw4ahqYHD9NfKhcvBKw3HCzJ8SClmPpmfo
/ipfAtrQ7gZRW8x76CcD5+1H7L+xR3xz+ibtdffJBMlG8Iv8Iohm0gtWWCtLTtrw
hUFWSMltS01tqqjKvOYZAWubml1cCsZDo7kYpsyTvF1qy4CL4yDYRY0RL/GCHlQv
VnReWFFgvuXtLdxGYIOEmG9kia0DHxkXbO9xIYUd67zH2IvQtr2/BvhIzVphoLry
jj09YQzCB13eyf4g8N+VYUvRyYovjGJUk5kxlGNOPKd/8YOgMfXzc6nkFz6K0K8B
NSxsr6rAmu/vl6r5WKAhbsJcoj7ceX+nPFwLj4TKm7s3aVJYUWuUaOZ9bFhsrH7R
sIjsUD7PB5i756o76PbzxbBjMugvdobftloNkqZE5kmZMl4CkOss9Pp0LDZylptc
rGrA7MHeBqAR7NeCEE858S/j5x3T5Nmc5Wdn8h1/qxIVOn6T9blQ1RK8gFwDPf3d
vVdLX/bqemNJMV8tQX9fycQC6AcYeW+CFsdQD+3m5nmTTkUJctPQY8QYEmwl5Fmj
pfPh0OW42AaQlnd72gXkISRhBHLAgMbQs/NeVH753vgDaeNJu45DPj2fEWXmt7ZP
unHEcPTLoQilYJCdBGcHCOOq+6dBwsD0LYY70GBVDKu/lC7LGpp210824/680gMq
h9sIC2T974v9WtnMO9Z2Z2DzTWPiVYmmtDBXnzMo0QxzVgPJcCSoteFXapCML7Tv
W+PJ6A3Yp47TF4qHO0+mdVMx85c8hFkWalGMn+6NTXJi4SJsJSb+gAWvEtIdVvsA
aAPNB9KhkjWFnOys/C1LMaxIHlQVNDI1mqmBm1yhDupDhlCqWs3JIGUqQhyl0ce2
oM8iqvsd0J23MTv3iwrq/FFY0Univafl1QJ7yZovJ2ZZfrx+/t/60uS7gZAcmYwE
4HNzM7S8zF5yXo57k5A33RqgmkRuBlC27n84f1uoKXwtPgFPvR4LOIfe7F8y6S3X
JXn1+kbh/UZd2uKhaH8sy+xcgkr64K9KKw332DknzdNmYXao0M9JQxTUvJC1Cypt
t1HIhfBtDnpxFIL6iCZo3JtFW+iH/AiNlMJIc05gdWh/fzSyO5MKJv69fyo+PRWJ
9NGjs80XV6TfIMuxqk1XRtyRdL2+Y3ef8PTkBebbVnJhViRxFnrsdI2YiwymkS9t
q/Dpu/rjY29KL9lCwrksFd5i2qchgBdQnOwGRSZeElK7qC8gyb6djlD2R3FKY1Yc
v3TykQ/d9InPQE7+9oWlQy/8JTX0ux+ZD6+D+YB0zEKA3aJMck+fBpt1ZwXbTCh6
1+FttToJXc6Q5nGF9N/T3sajqUyrox6zp7mX3yPqAGskUTX5xqwfB8i1vBD8oK45
eodhzW6ro+ie12NBno+AvHZaztLGmebnc+QRMuhz2ck1MwuoyTSreRDcPnFzJqef
ICRRYHhg8d8Zv/l/8+RmfqUk8kccXlDugPAo/IkLKo+TER8BSnrXBWwmLpwagCPQ
y0pjv8nnWmhs4KnObqZ+QTVKSxXgBBQ/g15ci5IuOx6nOfOfALP7oac07/PymOjK
PDkq22NhJOrq8tJHy7FRkk+0Io6VeforKZS/CZzIbEt7HX1puUclFsxIvHiYZUYu
ZPY+nx4HhdR0NNtEnbnr9d5uLumE2lRnFahTCSoIJH1Y5wAQs9WpOl6iWnhSr0s5
CiSixJP5eRrdWVX96tyGzyJQj2FDskEQkFawiUjf7ceGPiAVM4P4eae/vEARRBiC
SWj5u3ehAHtjzCqJW0cFcsyTm4HzPtvDU5zIb0JvrViB/ymH223nmjeluugDGORD
IffH0qp/brx3Vr0fiLmAbn0aAeF5owk7ma0lEL5V0X2b92UvVEAF5mhgPd6nnwJZ
AeEVLqrewbzSlhfwLpLkMq2/vOW/OjxHgGhE1OMnGGDp8lEzcnElVKDn5gZRjgCz
19WsEvh3AhkspRki0gT2TLzhw1cyYxK5GtdZHk5+cU3y7viAJyxfI7PVbRT8ZfHv
btHkTAyHxI1dYGrP/sQQiIEQwDYqbIb6UBTEA7pZeG9+a4Cw3DyySkqPmoiTGd6x
BK96kVXq1V2DUVEbt8nlpGiAzlhvs2BRGGKg5zsAwjYmJ2kQQ0m1nBDB2Q4LbzDz
ntVqx4Lg024rOh+bIxQrb5ziuhLJo18ZGJeDOi5yl4jq1GZkkWEdQvaqkGUcauHo
qefOgApWDXfjHqb3IvUk7roO4StJMJ5nk4uzMZ9GFcnwUxsWGJ6O72chZbtJMauL
67G5AyklqF8mEzItzAYpCNK8DF6Vz+4nX6QIVcaOt91uBkZ0HVodAZa+LuldK1Sh
VZfjod7nMQITc/8t/3Kk0Sx+UTf8OrP2UKLyJpUjwWbSuAAxwaYvh0K+aN4ypbGB
VkgbGCL9F4ACfYtW0zdB4kOFtLYwWUc3wd20fXuxSg9ATUAh4Kb3F+7YtaTuL3h2
ra0zv9UWxDO+vmvRypkRcPamtBTNevG5HgmavCJOlmR2EePIQd2r+RVyJPoAVege
3R2BKMjSI7/zkGDUKWP9gEnSlah3XDRuYsFe59mPY8oYXszosAXyOL3ZWIQPeTHg
LEYRD5nMm/SNrjLwyZ5SWleyrMx4D0av/qRr5Z2D+fvVyIydqBb7e4wk+AxjhwX1
4TgrKNkqmgQLozvcRWwUFsKYppqXIk3B4LNiw8jvQn9s+FxY/PXIruEDVQa5PAa4
FF4FurabZRei3jTxbPUABSOjFLzJo1Dr/1y71yBug/CpioX4R/L9FdDZKbB6WyPI
md/Q05RAkYcnYng6JW1F5/o4uO3nkSE8Rej3XS0IrmHfncvDp6rcxv3+x5YjAwI6
LjvMDT59zDIIUSkPKOOory6/q7zfQ4QrLWz/0dTjBVqLNRYzhm0ng3TfSw6n3gm7
2xQBEs0cD0IhxL381Am9yXqahPWI/1V6StGApAYhZFl+AwIcST9azhoayZ1Rxge+
pDKJYSbO66TVGTTZGmT/lwlshFw+QruAtZf8zaFb1JpRihwoXp/3DvXCm8k+HDRS
8VE/ooYDBd4L+8v5n8Ba4j/0bwyb/dgqgAuyroMi7BkaZI0wg6d8EFWnVVXLLA4b
RRM3wow7wsQx1CtQYet+xlfL7d6ekFbWTCTIza5jceEIM2311OwfxLwldHhHle91
tzgHdWtyQkoLIMLl/XAbEcbWAyMVsi2MrSCxnEjiE+tblUFRMW1yuzZCtEDxf587
JfOgS4T1L/Dm/PiLeAM6cShYxwITjCtxZVkl6uEPRDGb9rjS2BWaUyH/bR06yrPg
aEEtuMJPmhHHs1T8xcUV4zeHBXIscbAmdMMEUiuCNJwvrO17OedL2Wet1OaLygOO
k7JDaC51Dl/6uHeFAEpbYezmB8JZH9+PsupmUWMeyfQQzY0GO0X3JyzrBH5gWdWw
h3EspVDNQ+L3V/eu9iDp0veflwUYRrQ4YGvGS3jyTxrg5dl3p0NOKUw/CAmF2S71
OsqIslVEDfYcEX3peocWAxda8P0cwapaSX9yW+rUtxbWivu9OKaCZa824Cek2G1s
wZUjw10PNSfu74qwkClc+Gwp8cjNGZPTLkYGBHUoQZBvTNSj1I0vWLwJWfjKb9mh
vb70MzCta/tRZ7Cyera+P9OFRNnH3TuXcIKW4Qb1YRmYsX59fHrdZKws3EenfV0s
EdLxZEmUwp0Ld7CG5qclVz+innFoFs3NvSvmhu+RcSpkd0O5sd1MIPSugzH5IPjM
3aj+4gi0piQiwDWUtF6S/LFiSXISypP/hKJS3fKxVR2tDP0eexKUVe9G7JRdasGZ
p15BD+S//RZrSAkIdI88f8DduiAw3FNbkCVWxnND6c7yu5X78lScnDnt1oBjH9Zn
HUQe4pm0S1z4D9C3bBBz/A1i99amyepGuYEfKK1BRAk10KfZ8s0sQKSW8eaTEXda
5KTSP1mLkWjR+L70ebr9Sz2v3nlNpSzEIesEqly8HEcJQ8eUwGzVCBE1wzKfYSC/
Q3lTLEpeBnw4tddwx2lgmUlnleXLLD3F9vHyVU4D3NZpX2l+unAYtCFW4Z7+rWCk
AJkwfbOACHF0T0qSh43cL8k5u5NP91SXoBWU71bm4GP6oCZBPkJquz3kWzIw21zd
KRZ/LHqWIoC33RHPdVUYAcaQpU/Dpsp1fpCsdjrBGy1WDTX/cAPOIWmj5wbqq8B3
HGq/5Du6MuXIBMB9lgFH1c79O7Kkra1Xpk6wPIsz8tC2l4spiXTk/qBQuDnNdh67
IDFMI8fW2ss65fkpbV3FAiDafKg7/rf71zfDtr7u1QMInT7lud62cD1LOW8FE70U
+kD4LCKx18jO+XzyWbEkKFdCX132BLx6G9trHUYYqG7BbZtYFKAvef+iC6l44fPu
+Nwled+zhT2ZHRxEWw/XwhF80FH6VVyCXe3i7QH33X9Z6zTeKJv9leYLWBpe4zur
Ki4agTwx/FC5AzD5DgY4bh2ZK5GlK7rLZ8WGadNb9fUmorPON42q/i0E1jlJ7ktS
YIE8yclyLH7gBulMmpdSaUsdKncoEr85rI0xxZmZ7tzoF10Y8Sxz/UC0Kf5lSmg3
PFus3/PfhDNtgZWk0d4zK9+MIcTZ4lVxEJv6doNJKuy0M/7iyziyvCyuiOaK7+t8
EzvwnyPzsfetcJTaudu3ygcQIIL7bM6hz4bJGVSoTc9/pmOll89WsNTam2E3sNMN
S/XFQkXSB2unBec+UaD4PXb1nGKP3PfxEgBBXyalA7VX2fm3/pxAirhjLI8YsECT
yaYkPP+2NVkf973lX6nMoXotFjQyWgCmwfZ8lddSXx6hvRPeexLYWdXjUky1z5nv
QFtXKEpePZcdluk5UVKxnMM+XpNs2QJtwHiEG5B/q8FSwoUYCUo6ulXGMf6xOI9E
Isnqbs2UvfnXiI53LwyoX9/raidPd8z/GMq6wdjwnn9HzHjJwKu3O6mzBKLn5UT0
0u4uO3ya5M2NGt3aIpJGrWh+dBDeG8arp/0oLLyMnE9Q4Xp7Afy/QquzOgu443E4
pfa4EuWHPonbNriqOmuf9cpfLTiULrwA2W7LSAA2uMzVaJO2K2cIYG9bpLRYSOxc
IXLelzwyi792h2YSpAuFsj4xwdjbLYmOw8JU0eAZfOC17TWvJwjeTiSph3/+WPq+
kH2BtkqE9CCnR0eOELKGbS3JR9E5STCTlHb0lsqsssOV+yQ+zfsFQD02ekasXVuJ
VeqWuQbT1NsNeiRqWfDMZyvXUviPCPrdseknrLDH4i5tGRjdsFUQbVUZsCp7/lg1
hD+XtkZq0EgYysUW+1dWypN29iZP8G5i+Wpx2MJeLkNFzQNknZddMOH4qaOpBXKG
Ur5M+1rTa+I+3aRyb+cwHxYsErWcVraDVbZSVSWOl0bueB6j3yUdrOJHQ/u35JWH
d0KP1LOd0WoA+QZiI8bFDwjjegTN/S+Avkkp13RERs20VCpuLaTs9Id4pIhmjTHx
eND2nGCow7azkiFZjeI2cl1p/db1vWTq4jv1XB5IT521pVAk95gZYg6XoTig5gIn
iAsawjIQvJh5Ykyoyfa/H2rZtEiXrSUXS818U6qbk2e+8aIuVdew99lYjtq0RJ1x
9F35D87B33RR9dsfBu2OTJxa1XiMpZ0xU0yDsNPtGI5riciJPkidOy8mGL39fJWz
40+GNHJjRT2j9k5xOjgADq1kiaTosjKNfcAYgmhaOTCXsS8RdhDV8sv1BTT6xUtX
9UJBVXSN+Y4Xxlcv1YeoD5RJJJX2el+Y1o/PIOsHo2Z8P+n3sS7QCPwUyCjlfF4d
MDwzfgBNVOJOGGctiUGm9ezy6bYzMZ8x6NxCGIy4m+O36nv/tLLxDf/bSWwrusY6
30a9bpSg9iKLXsYhJg75iPcN5LtxUCsnuSggidHvcTCPYDyG89eouWDkRVmXTONs
ufAGx8L4/rPTwebmBVGgSpgBHrwUcYw6tkMWDb/SzkmnpM87Q0H7RC/E2QoCOqCm
sAuoP+9d83KlvWzTnwgMrymLCd5Etac9r7NKdsmyrwCPAIptOBhS377+znutITBV
y4vs/RUNJPNYJ0k4Hkqy+2X/8Kpardz4bs6EDNLLIHQhtlTiACGUTf0NNfn4dFW2
wf96is6w4UHsv6K6/N8t1JuiZumxO9BXCVVxnK7779zTsSqBcM/E8elgh7bEpodc
DK0hBvbXJBDpEPQLMFiNTETMRfaB+XSXKu9vWWrghPqpAPVBmYAuQJwwPPbwmGd4
+wm+qYThFoIlFfBNOluzqZfaSuc5fvgqMzQ8uXIH5vSrzkn3HW4qTkYxQZg2kvHm
0MLxo3geVpULHwx/ke/91C4zZr9NslAh6cdy+GucBRjr0q5mc6RZMudiEHm3M6IB
1Ylj8AFYLQubfSAOK692ZzQebAiaB7/NX9c+bdfy6b771BP5zxBsCe6ZgOXSmq2r
YRIx4H/BgVdFOGH2158uQ2SE0TfXr9ncC+k8mzdZq1+hAR6eUTTL4XWi/6uJYyaT
Egwnqv7LNNBFozvLAmyeMTgI5ILb4515vI/hhs0BknLESSzOiQMwlByGNb7ogzhf
3eV33G7qY5nkGMv9e9HflMy/uehGke13MqHdnLyd6II7+lL4cOH5iU2nUHZWULSh
SFL4gYOcx20WfiLOlqZcbkzH8iHVxQAgUXdklpAS+lHUBmtUR/1VlAyQH70X19YI
phBXi3X5MG/4ZivbaGKVA+AcIo7y9LpSuLR/x9YHgT+MdoKhEs2U0VBZQK/GSvOY
RqImp/tWARZonR5Ocvd9aaVXcLOThYK3qi+wvrjLcryOAiFACoqMPaIKaGDOETGS
X+ZQr8xWCWqPHbDeT/4Kf860I1kq0fiFIDjpOnCyVFAdIWGXdvm9ejx+mCU/sChY
qECF32O5dDOlSFxXVSJQFJmtj6oLFU/A1h4Mwleqs+fID8YfwkpM1r/sxaNCSnJP
pxs8y83M/b0K4MmVRi7u1rzh7YPexm4/YG80heum1txqFyqA1EdtDvOehBryqUso
s2l1ldVZgI98nHomMXnlXC2m8Jiyk2nMM91V216ikqtKb0psm/T5V5I1iy2vMhgX
QhlfI22NBti4NJMnEBw0NP4FQFowtiHeCaWH2AwoTD2wkfkNsJKvbxsayE3w0DqO
q/dmH0EwhdiZaIpz7CI00HLQlY+RJDqpL6nvOsBxQ1zz+R8ps2qm1mjCC3D+XuTq
t7TJHw6VYoTEn8owMbys5Bvl/540D0MyZbGOe0i7TuGwrnRCM7Raw6Wx67BkZKfh
4GwFh9o+OlWxIwu1ZaM72h9ahM7VKfHkxmYoMKwosOsEBZsOKxGMGan1SoFPQr2x
d5DRzPlbcl9LdGzsUfVwZ7gVJYFbuq6bOYf/SN0DWnLPDpN8A/p96NhlIqZmKvaY
gYZE8UezyBguw0cwQmYJ6ijxgg+k8TKBLXQlK8N9uY237JSF72pkrEaQSmdbwPlu
vyPbYOHpxGK/4/rLgHFDyC+XaIhxijnlAquDZruyQh/nAOZdQHo8fCailHSetU9W
Oo9ijb7NwIp1bMW8mkmHETZ0b9/dXlkVlJO2PRGXuOQiBg9Jy+UH4gFkVBeD87IY
vrsUw5EMWCrKuoCwQ03QykF4G8FJKrjDnTuoEtxHBVPlBSsfP47VmUlEvDBCrXyg
0St9LKLkr1yEi15gyrLxHJ5SAJO6ouELR8/t+Y7Gxts09fABnDMdWDukWLxr/5lR
nsWY5YLWn8hyph/0vTuUrB2nDLtiyPc8FjkGOxCaQ6H8iyODvNMkKoyPquTeaLe8
2SC+mygOH7HGCzlyTlgRNGIcgOb3F44Dh1RlTMbsgJyMcCKRly4GfuXZGqp2GgjJ
YCEvssfUHcTQGcU3kIgz2Z+3PjI7VxAYP+ZOo6lfOnOwPbi6ePwXPoKdZERRenja
QffPNVf1AeSRMwLlBAUV9urna/Rp9PjEPloGSabXzR8fVWsDpwrFTqgCebclpnY7
sw8bsJnoreczWY5227RhGygRmeZy23xUFA+5tkrvnzgTr4wibRwBuS9CmbYFCtqp
TMnj5mMuKNm2TeUMmbmQ8LNwCJMCq9OP76lpYxitmboLUhBqa9REACqqqVkW08bK
/JQ+yQP5hdnZpniyWEjSCc/cs3KlPNPJ68kr9VbfcTiYpqLMOr7/JyPmK2/5H40E
z98z0TApfYIzNdTG9gXPkXqLlfWYALk+tN//uJYoRpVJ8KZJxKYOmqvgY9VfmkhA
lmJq2KNM7O/L4vS69qf7wXeprLF4NTRsgKR0vkK188yCndNpzyNtQoNMmkzf/6y0
WGVdHf3X71DlnH+96nNAkn9tRjxGz9WHr8BiM4suave/jZ3K2KqmmUQiHLeiCl6R
jOc4eZ+vZDgPJ5dOybH0gRZJh1/j20hNUrc4s0CDLFwNlSHmmUBea1qBIOpcETqm
mvtbKSAXBnWSab1gHTkvgG99x7KpMuoD7vwluVUxO/QWwirWCCHEtp1PN4FpEf4g
90jCzl8iotdKAizFdC9STonm9G8wjyFiF913CL9yERKfn9uiFtwpAIoLm+nVe7QU
ZEk9ndc817qCUEKH7yz84A5gqaxdIkBvtOnpapxfgvJfmWoMgXfnaVtp6SZ4HwBG
weWLfyLP4NVqy/9QS683T/GUJc+J2UzB9mDN66mwMxKGGR/vuUZP+RP8bTx8tVnF
KI29BDm68iSjgvsttPXZM7fu06NwJ6Olt5Y7Tz78hL9hw4xEg4S+HtUMaF2roPO5
wkv1sdBAt2Irk0an/0fOEjMtY/5N+eBbRpkDE9+TgcTOAmK5N6O+Wk49Ggbo4ReB
I3scpQVbcrczAChpCDaPaHc9R1vZIUPIj+/Jc+cP0HVbKMOH0Op8HdGee03Mf4YF
lCYrXK/edT2P5BmKyVR05VMuq2lTmbXcLEH12sxPmYZ3tKE+btsh0DyDVVj3VtyZ
4axNXzNHYIZR7ZdN0XrfT+83qJI0JN8sHlkiYOGXNs1J5oqZE1TEp5F1GJ/4m7iT
n+tO3HdYoi8MY7KP2gmMhVovxPys3pl44UPp5uGrifqBMC2vruLBybqy6F2TkUMj
8T2IG1fiV2ukc0hVmVu6xD9SxPUvzDyXSubeaGiiYl4tMHX7moq5zJ8+6jBfntMn
s66+NStO+eunDX8ha4e7Q7UytS/kFmk71AaK8GjxlcuhWB0Xo5hBDOpJGgfIFgPv
llluUfD4kt1CxkfDbGeg5f5Fx4SN2EH6g5pwkfkGqbC42gObbXPq2ZTnEHRKqq2f
aEmAnTgCL+jJWBxP/+Q/dwKMYD2T5wvuW9kaEpN4tdon/qFrkfl9Qf1JrmSHLtmp
fSbVKc+KjLI2up297Z2zooh4ghk6zb/6yRqszAceV6O7fkaHbPBJay/OjwbYah0o
j8Hr0y0/isZmtKhs9h+b7tBKx9UJSKF7Blns+2SVMZjiXa0BYfTsH0P18EDZS++d
IsL3KVWRwOII713Ve9z5XqxpG5xvYu0mnyGNfFe2ih8/OEqF3Mi/tn55eFsUFzwf
JQvadQ1RxhwhbwYMRk9/S70JIDiEG2eteYJuDnNOpOFH5kSS2wMDXjV5cdZNaUar
1mRFc+zFyklHvAXsgzV92SgoALq1a7jkG7/tMapk0WQetLPgZenpOKDykFeP96qQ
PNwhjdgbTN41phUoXTqYLahOqFyVd2mG1r/oJQXx8eZCdICtaMUvmc2Y1dt5xn/g
QtTABy/jt6k99oMDbwixrYUurv14Aq1upGb5Iz8ObjZD1QJ4p/QDRorMlc10w7a6
DGNiwFauZIYrM19KMMfoAbCxG1uIFDIAG6DaG2rH2JVHThCs0Vw8yg/sBA4sGLAw
iu5becjPpb5i5Dp8VtEWdNDuttfFK1+adaYoDiUNXAdA2JMDWzd5UVEhDbHjNGgS
kto4GzMtXuuFLGe8FVoyE8fp3LVZ5AS3nhL98ph1MDfy+Nx0t9d+KgRdNLfpm/kf
K/ZcwOHNS0Uu9BNbAhVeIUho1XOagDP0OrlJd7Uz3Kl/B/h0lSCmF5iLRHcNZrAy
gKwTQbYRh54m+bjtqnlwPmP0C6EeMLbyZhhVUZrcpT12gMZPtCLqrHZeaTDSHN7o
9OICnKkdqMx9XfsutvAwed5iaCPmIPHVYJa+C7YRgptn2IJ2Egw6s/H2fNukwQQy
5WIICC3AYWcgy+yvg/eSCP0qrSH/SORwDkZx+mYgO2hWbBvkO9FptmRU3tgWaVLw
xFyH5by2nO5NjSla7ChNXFdDWXBQ+wxuaV+fwjUilkwzjbjl5HfunGI7mgunCqyV
dcp1nxWVlYMwh48l824f9OmRKKJxeslFWrHKnxDzC5AjIwpSabdMk72nW1ufCBvU
IbYNpkMcJL9tYyuo4UbF5AT9P0b/Zfr2MTGoWsDMn5ocxr8OblkZQJ6PPVlL2Hfi
W1GvsfuRu5acKTNEu5K2MRPfmJbsQNsD74BUUW+LAanEJ+LOZ3lIxmynIdE1fQ+I
xpCae0lkrXTkARcnFc3+HCUEWYJ/wKER5ah8/jeGg9RKjGRFMUzjZZpR9Fp6fqPe
PHteGL67+zwW5SQAOKB0Y3A9cxC0Zqpb45xvuw3iPWzOhduAdBk1TfMvEguEnKoT
dZzPwt0rTRlHbMclLN4+XvnvVLEXSpPSBZBywvCtnetcdLm1h85JmZ/gz0tS3Z6Q
GoTLubxKVGZlSuaO4BRWfUn+gKuGgnX/vRJa8V6YaHEZ1rM5b+7AFf92u5SyZnK6
hY7RB2YZOLl8/GUTpSzUsmIw86YZISEI3KamIjfi8kqjgclASjlTOvwTB9QwEXcC
+LPml1vp6r7OkpyjI4fgRH/HQY3BiWNQZt85e22aZVkCJTtbiFx3DpDyrgr4EQKc
+9G7oKSSk8EiBug3fyZEyAa08hXBnjHlsFt6CjzVufxlN27+dVf546RM0pagAHdV
Lj4bZqhKd0w7LtYP3ly7FwrCjQqPtvmBVs/xJLXUZPciliOap/uED85qfHMaDcwh
SJDgYhiisoXa7EUfZYqccKK6ZVmjfuu5vhcyI4FCIsUddiI7Onxz/eT5k04/Adze
EVXMODUvLcBs2cdmbybbrdaExq6Nh+zlON22eyOn38YNclvHzLdt3zdsHD4+th2U
Fv/EaM+5r7Xk58meOAhlctY705Ytnp0iPZovwPkXT6hTVQ+CwzhMy3magOlF7hx/
v4CbT84UWUQDC8UB8HPw4Kj7sDmqymzPdcnw0+gRYZaoT7u+m0PDqgtlgmUlIrrC
2q1WRqKRIFSSu3+ZPNBdW92QPR4evkqheA88DSzjCClJfdDTD5C2ha4Mk3JugtKd
4eAvyNz63qlO3tvnc8d6q2jf5PyaRdOq8/dXCja7qrMwxe3hvQTm+ehUI3cMKvE0
pOEhRnjjBt2fo6yHEdgIQ2Z+DyOROsHrvc+t6hFxtb1ee5aUDxZ5c9KlOS+VQl2x
A1QMErz7vJSUJ5I/oZMvriTed+eEIv8864qEux/BG50tdFr7D05YPEP+NqYSiUwt
rREeRRV//2mAb9x4V9wfEZDIsTykxkN9XalvAHwalKYjYLzS+nRqJoJNd6QWPxgD
xktjfd2Wwbi/CeriQaqtTwunZ3smub9KQw4Saau+45IkxrUje+lbRH0FY6uL98hH
EBJWgK9ghlcxGOw8Clf0uge5mxB/WN5A/J1COTS6s67ki3OgleaHrk28e3Ne4Wfi
24W385tTawWQ/Uav+Pd7YQT3YWZn2K2Qx+nkoWszm/QIKwqBtWPyS7dBlvXfyeh4
8v1cZvHmjiEpqutFYLPqSEfD0BS9ydE/rWirtjg3KMo0fTz6xJxTrZSxi/zJaKuy
8f6bqw1hlryG/nz6wTX6XiKz1FQaIK1BB5SbPTLqeCYBLa4IbztZYTEBrTB38PM9
uuk+B9NNh3LyIjCpJVWEr/BlkDjAsJgPT/3Mk5BXzohcCzfKvNl2qR6nuVVDPccb
XB6ws1gTNhvO6Sfl+QV/TfMiHilUaESZXRlTod3vKwSVydMwmrHv0fZFcGs2wg9h
A/KKvsArjZ9kbTFuzHk/TlSTuMwezMEfN/X9VhaWMclGZT9tHab0h46rY3iFjx8G
Q1DlPM9NTy5gTQB9gs+Tx/O4ou0yoTc2NSKQOaR2r1kV0wQVH0zTJvKrGyE7i4KN
88T6VdaGPhOoZrs+K4Sk1nZKXTxWwNuIyPdNQkv6thXg8Z+FH1XeGA2E0DrNcB9m
6mjt2QfPoh0d+9DTq6vHFa+0Pp6GoUryO9nmuVu4v1OoQkzS1g9xf6R1jZutyW74
Tb39dSHlumv+nl8eN5pPljCOJ3E25hFd0jZrSuqD+pJa0TaVcs3uRm6j7/fqCT7D
be+Mm9/mwDbnKVy2DAM3RZCxVhCD5cXBnCwxXbLbggKdp12MGTOZCxWlpaWYx4Tn
FZDKIguCfpq88629pTqjLYccs3VU+/nvh7OO3Sb9timUTIGizN0vfYeHdrhQ9tiS
hTwF7tuWiZsYszeUy5AyjKAHUD7nYkZLCYjh4D86OT6C1qsBe6Hh+7KxdskYfozz
AGFPwJZ4QqMjfZnNMtZrvHCGxznugtdaLA3PLbdy5J/ImzTzhX9NH8HbSG5fnL3K
eWQLJ944mDvQrWcnB/Wk59Qy9cSg9Odctrv4umI3oNkUgr+mD6mmJ4s6qAHP19IK
1YZmI2ThiZSmeDG9YtRmBiZZjYym+ryL+z7hQnSWewDoLyL4/PrLCnOSaG575IQX
ImtN7ybKy+AW+UAwclKZt27RC+KGCbbe3jarjio2cGSorLOoPKgm58eBqNk/n32i
GUyUxllHHGfB/nWeKYb6cH/SYwAIdHSl+MCp6I9cQZrG08ztI6HcrjgKm1Jh+euH
nKSkI0AtIqX8UsrdYBFudmq908SAiP2X1o6agdNOrrYEcZSRppvNq0K0Zzx7m2Tb
+ErBmyGVRxDffAEq2ak4dJXYKaCCzcy2lRwtZrzJA+EQaxzu56pcG6F1IwR4Gek8
63J20v61yJ9L9sktQ+xXOMziKQ7VEu/AN1oNCe7cJ5udEOT+lDb9bjWRaRVeiKJ6
bEzWXzIMu0T6xuwNAp+YUTybRdkfQ6mdOg5TmdVot2w96uGVg9VgGEX33sr91H4s
UUO0g/ZHcQTu+CJGRu6JZsvSU1OrKXTzCWe0vVt9HIU32+2ZRhNc5xCMLyIcv8bc
yzonpuBMefKAPUhGQe2jqXMpVLD8Z7i59F9M3Qex8/5saUcpNrZrLE8MNYy/xA/W
DM/ga1E74i7inrqJS6nmUQHRG3qYGtM/2K7qNE1IHddvxI2PyfHyUDNcJZPdrdqS
QhJyn77TAy4hAGOinkydA9Drb1zhUoDK1f8L9Abimp73fJsVD8YGvwWOcvKJGkR1
prv0ZEOpaCM//qdHeZJn2X8w+ze9tiLR35JbPmzX8aCtZoxgiXY1bW5LPK7chh8d
Kin2oU27J2EUW5KtZIlmz2CbJOGAtMG3DuzfT1XD6nNsZcPwIsJVuia1ufW+yEDa
uOo216Ijil3eMNcW/TkBdoieqmWTsIAiuDpnGtIXI0gP/dZ9A0KpSbxDBMfKwWM/
TFXN3ZULh9Q13hK06QMonnVDzvp2VJDeCG/8+g/xRbqoOnFVnYDSNJzXi7JHLpuK
+t6P3vR7WXHPf0b/207EglCJKSoKSrZYT3uQFeqci2mmsT2Bn+Un9yaa+McqIEYc
ki8smJfw5ov+bqOHCunKW9KPs9RIiBw5k3Xr8gE62qSiwbGnvbQNc3spc0nNJj37
QjAAFvlauU8NSzSqYcdiK2j+XCRoSEYSuaotdodmpn5l20BN46HScfke6alLae2y
abEMbjICJ71MRHjr6CejWEMsyeiuvHNodMsWKxpwUPGYtg/cvPnBYCcAdtPgqC8H
vmIEKL3+QUIhPPyDMECptOsux8LZJWNyg4YBIDCA5r8mJlP+2bDBc1UlLKKWJUuA
3tDnm4eynIrLLU6CU41LatzJzymOaP/7Itjqp+QlIrqjNVUFcL9Mhl4wez/hV+x2
bGcX82s/H3Z3MSjUF7zqht8Mvt6C7GtkRs10VdaL5lMSTLOML/16Off1movWwqCK
4FBragijv84txZgt5TgIapYu6kqqHlHsKN9f80XRZkAUQAp0I4twxSIaOKOSbU9/
zao5oLIuBHDaRFRPJCcRH7AsAFwbxhAep6uEE7/SZrgkj8Y6f+ngOcHmo58qVOcC
Bbc/qzt4iJGuwp1s6zVy4fh0j8PJ3+mbwaBqWuunXfqhltGPkk2PrExry9e9uOtu
AUjxoRR/8ZxeTxjx5VM7I5DlzgOY2Js41wjbYYcSlZY7+Yf0YptMsejMyIzSH/k8
kWfZ9+Hs6J6FAk+HfKa791wWISBxotUOxA7x/ePHx3Ti839kqlhg0t9Cak4dy2dk
BRBDl7OkJkWHDQnoH1wZ6AD/DkTQwG7PHZ5DOgJKFFp1XjWsyQSoHBNuUYWiJYkf
LM6oXOdbI4sJd3ERH/C/5hCHXj2GQ5yTwVt9y3lIIZuLJS2kTQHw7cx5TwkGWclZ
HR4HsaOhuGpZHWp12omX7UnmqSTKLlJNiRfc6q/lgxvvrWzjJbTEqrcIYD8I9eEC
EKIQfdqXVGk/G1huTBQfOVsYA7Nz3DZcTi0YaqTYuribXjRjcbalifN1IpZy3hHB
f4EJWac7o3X8xWEF57K/mIio9M7FzZlpAPCJZ8e2fvJioGuZGpjw1ND9vQ8ZIYf3
V9cw8tEYAqz5rfgxU82LYmd+cAng39TK3w2/JGnOpl0Pn+CTH3XKJTBmPYZbcEVf
b/WePoG/o2aN8XbdUZoP/gT6G/y92Yfz/VuzQFQQGOs8sHnuTVRWcb8KBZsOpVl/
2KHM1/ie3dVCbu+h9J4EcQYypIh7fnjxO17NHD2RFoe0AoGv3xGAD/Kr+2noWNFf
inV9TZN/ZdMRtVGavJ2ZoZMPCogoWSZqka3d5fEYdqyHb1LgwbnTtmKwDJy0HQwO
/toIJ7VwvjNTG0CxgTXaXkOvnLjOp0ZRAqp/AdTQfJ2bU7IXOYRmJMLlg7esLHQf
KFeVkF2L59RoyHb64O972q6iZ9iz2sAINZ3d9LnzLJDPV8JJq/WI1yMXMrbfucWI
afSGBjQdFE32Y4O5dYUXQAEwqGaVrigzEkCPVmzx0uV6as/4hZmSMDosthSpteZJ
Lm6QqNJKr4jcMTJ/AMliM5UYHJpljA92xMrMgoRas5FXsieaoczU3QUX2E+3BKIu
8vHBAe6V6GtExCp4GpuG7tZ8OOOXrdadsHitpb2QhPud923HMtR7/0XOZ5BYvEwL
2Opcu0YcsRVM8Xefh3AncxhNhDD9744NcT8wUYDe2a0tjGmQSQTyDYiIB3Ox/C0g
VOhQ42wdFUWrqK5L57z2r68bwM9ky8rVdSFj0Gf0iRjCbhetYNoWBReBjdDI/4z0
L4rtzJxUzVyXHRncnS2b6xKZa5Z2FJfG4r6B+RN6RJISUXgcDXHU50A5qIAjy5lr
8v0F2cgNp0qPsaDjS4eNo1+ubWGG6aZ/qwByrqmEG7uytj+erFX91iPFn7kLJjAD
dWqyGRJoG8/TiEKCLBjqY4jpqziR78ZdRUJRSOeUWJ2q7On6cX+904l6qbpc+Ck+
1P+Nz8HZ7SfJ0XNHWPFA59MVD5ePh8/j6W/G/xpwJY4T/BWJyXmYyLX9Jo3OWR1b
AwDYuC7OmLi3kLHQoX/Q2zrIyf1dO+h413tJvkYBRnIkaSkMuAZ6ckM1HIJUizQx
pls2dAXdtN8NG46Ibcwb5nfU3L8I9Tde+/uyl5O2tskLyNolBzkpMJb6EN2i2L3q
i3e6MTC2gBzHsTR/eqR+vEPLi94YZsdswhNtLoWBQovYRhuGaqppOjQaMCw7rIGr
8jpKnvkjrHpCEcz0v5TU3bYkisgStOLhl1wQAYX/4ouaOBIJaFQQkyWEjkZDP6OK
yA5I3XbZNsiUwz1Bw/FaX3aqZ8KvotME67lerYUckooZN1HfNcLAggdiHJPup/Sd
B2fbOsr13uY+uZKR9jpY1BXwd7l0EduNsMaPu4crkqcV6AW+Wop4gpc1FI4JlF/F
VrgTIc31XqXA95xAoGDw/EuYwVrMa6rov2+YUwXWjvKU7+ICBP5FORTd5FJPIsja
xhXXzomJkz/JgDHp1L7kmWY5SAv+RouP+JCCrEaK6Af9pletXGYvmV8xk2Zo/m/u
wz5XYoD8un5ReX5kyq7Q3I6Y3JIosiLroHU/gPh7By0xLHDpH67eqgwXDQlKwACc
nKlo/p1q0DJAY8cfVMxv0GpPyjP0+a0LYWO4MDWZPxy/hjJlwpYFkJkJAbZkdg7W
OhRz6agt9wB2WLhN6RpkFlc3Qw6Rbe5j/oVi8EgCVNCHlGqpEcaCzpLRnwWaMgK7
/3wP6pnRL+2PSC4Zl/kT/lc1R3XGBUjY5qxQiShnD7keJ8C1bixtjfqjQ93FD1eH
wIxypbkZ/zUtIal2kkYN6X52sYz64NjaeieazB4Byn8ZD9VZ8I/D1GEBv7ULhQHQ
NEjVuLI9Qrw8C3kN6Qi0nbf18cjGCbLlMXCLRPC8fjFiLGfN9QYAlzqqvjhHfUAh
164XsqDfR8xZpXTFp+H7wuaB/XWF7vNURJQQojCT583PoP84cq7tTqFlP4ehokFg
2LP6x3bdhdGeNbrFaxNZfeKmELk78Qj0uGi7nXvpAUsIVgx0hwpnhvH0ZlBPPx48
qWSk6r3l4lA1doE5blcXZ1Nu33L+uUFr/3ekSXf0906sfkliFMnDrg2Yq2ECvEFY
wNE/myek174yHdRG6FiJf7iYSpKiOaOQLhXLC/UTflQ6F3LDJktMaSiRPCrJBbYB
QZlP2riMTRWiuf97nh3ItLadpPEqsFudq6hyqM9x1FEUIiP33ENHWA653Ge1+33A
p5Jr9RWYe13alHg9KnBH0AW8kHKg0weWJjLG1dKznDLbVdrXmq4I1gupLMlfiB6R
4X+6UPhdCKa4ULyk42a92aqlikk1ERMW9J9eonzVvBSDTuZgA7v5StTOKa8rq8m1
qbqulyDIVLksDnnuRnz0k4cBqg/tg4fTl3RnnEhTC1PeYGAb/60ruyEOcCUEQhpr
c2t0/Bc2SCiUY+HoAvQB/JM7CLv0dFSboRrMlv9psOEpCVP6kyEirTWasVigqGtK
OdfDxnUMyIjLWheMD/DGPhJ6aoDXT+HdyC4e4CMLOfLq6kNdzHbPNhfxp7IPwsqn
JsDwAyjEXANtZiZDQC5i9zNad3X/6LFPpLDFziGR18PUajG0pjN1N6CZhIAKE83K
ec9aGz1+vYBBtdhb5KtTIgsSLTEl+mam114MJP1vJExQu7qKrtuYMu11UQYO6rkH
w3dUnE7hWSTKyJTfD9K0XaWVJWcZUG8t8bCGNTtE6w/mGe6/Hm+Li0jHiXCLOmAZ
ucIPtK3wWTFMIG2eDIEj8T/cF9AbKX4OY9sUWe3jCKvq+DiQpvZ+/6i/Df5sAjzJ
dCPX0Ju/YpyIjX0tolgbFgsW5RbrdTQvDcwMGkzGazlxDueeKxNeSrBwpXbgFAJF
xq34qebm+9w4ST+LYNWHT0M0cw75BBZdvDSNTiy1EVU7KD7yptt08RALlUnngoIK
M4Zp+ZFGIPDKGQju+zehrUFb0gyzNYQ782SVLQVHAY3nphlNHWX98bhiseN2mkVL
X98U5FS7mivHxT4Y+/NpwVHeu+IV+O+GatXy5jCcimGpMl3MYi95nojXwREW2brx
XZ4uN4v/RMhG0UUiuMFCVJ0LfEwR8NwkmW8+P2YxuZY3htxY4nhH3Yqnxn1QlAcH
9T3wr8iMxDAEUZY4FRUclBUCb95uRi3p3ek9ILHtvK52HOEPSJK8zqaZHUetT0t6
geM/cDIPNw4QCao8z9pAD2hVdatzXJl+jAXlTTiB2umnrDDe6Gbtye2lltI4bqir
c5kGNwbPr8kUV6IDQB0JpuhYUaLRAWW0JiyqtbIzeyaMMz03ybfVAwZ3ySifH5Cp
EWxJCyy3/bEjIegkZjUT83LQXnIqi7NoaNI/Y43Vb5k5ceNoQaFpljAp4HR4b/wz
yGVHzz4eJT8+W/znCzxdBwtOLI3QFpmoDHoEHJkIeomKcuztLklZALDLJoAe3yiN
8wWBR7oKpoGFD91hswkXz2ayzE4G/Fp6tWUFh386k5qf6ppyZfeZmXFF2eKfQgXW
BqAy0Rw5gHhkbXOvvhmFe6ht/Q/joFNY6ZRwXHBuE9Wx6nMtpUCrBX7CgzM2CDDH
3FqHYDlWFLqeB4VV0lz6/3zRKPH1C8nNveQdqBDcTXGOub+4kgDdJ6NeaMjLY1cq
DnsVWXfotTKGvLgXmBSPK2BGvp1Dncx/LGbjHzwkO3doSos9DKHnTkO7Vh33/NDj
abyG7z8VfXe26a/nEO/HFX4bDxjvCNEVSShMfmRwiLzf4m7jAakIRfBaGaO5R+S8
9cScUQHRw441OLTD16t9JQt5V2urgccedgekBAx+sYP57Vwe7ezxEtkYNl4iFpiV
XK5XaVk6/hCsaMQdUUEbcv6CQ+2eQxeRjChbsgIklqQApx+zb/6VQvjD8YC2Ntdy
j2Zthgf/n5ialnm7DZV8O+Gh6Zn/zURHfd0KuieL1U5W1HlEiO11L9TS1JKBcGH7
AN1fnvKdCn3WMajQwcT1wDkrP0rwdzkKB+C2Ub8ihUOwTVfOa+JDf+DVrQS4idT+
08PiRbFg6IKIHo0rptCv0ZTs7XGqwF/w9BFVlCIQ3GUBLmgDjfIGEdY+CCrcX1JG
o+c9ADHRiGgj0GNWgjBFkLn2DPA1EpSggZsv4+Hq3bfgHzsFcq9YAkC4ImeKW4DT
4G9UvkyCzBc3RjXtcIWSPvu/5VirYfutk8THioO+DT/LkQqRP0XX20KgAQP1pWrQ
C5hxOWYfCHvnJKBWytYRMoJalUmNP8RZrP8LfpZn4EVendieqLhrqbYp5Qt7JDeg
gbhENIDD5/QqnK9FjEBj4i4aNvJdBB1kvayerclHkrNuy1iTBBrcJY937KTAH0zf
wUVp9edgSDprFGCzasw4fW0zPe6PWaqmTyXJzJdBQTe+i+oMq11YjO4YwFvdih8f
auDLDH+p+ivQowMT5utsdsWbz7KIQLwB/F/B9CfMTAih1vBJYN9KAdcdaKbzRbQ1
SznH1gCzSMh5LKNnU6sZCQ9XUoCP0aHYVU7btQuVuIDJjgatTUiWiB4n8tIfRyzs
+eyY7MLE8GpAr5Sw6X41n44n4OINOvu882LPnZxQ+z0uUj20ZjsPxq0oFETQlAia
D7+jPfMFqqlnmdbMnCCY8USS5KAsExdCxDlF7n0D8H8A4HR66210XPZ4/Jpjgqzi
fWDfBwX/T8Fz68e6nk1JUo6U1CX5vf/4bpLKhjWej2nCZtw2J4A8jfmdvNiE7bXz
Brrh+hLMsMEtfEuGJlBJH0Y3u0Fd3trxVzTe3LsIQWi2dhC1NbNuwyzpF/oEp8s0
sWy7orRBat8JODwlWihElxPCJT6UaD6E+EJTlVtPOBQW8EfOPrVKyHkJROYVO/dt
wCUCgoB2uw3nTT72ko4KXNLHWBD84egySl0jC5rGciNpB6joph/842mslRkH6YBr
ZJ/tLfKo94lJG4OSmNGy4XsVxErxJy0rn9t46zeLVFwbTthUMZtuPCbPqcjseKiN
HIsnoZ36OvbKidHHQdU8jJrHV/zpyzTYGZes7jBKkgRmP5p3tmZ+FO19aO0zvYeU
v7voxCnQTt8jWkLZ4kW5Jws1pbIb14pErgfZ0pdKS08ryXhUqCyaX9FrmhtcELuU
WYdQcGXOtAvQdKe865o1sX+j847qmT9nQe+3L7GGx7Tnpd5dbsesZK1yrXCNpmK8
Lq6nwibJ1DpCcX9tplZajQ+3xL4QtkCPp1UfBjW7A6xGo+bS2a6GN7IoTIX5/Ffy
2+V9s0rHTUslHYvhjZxgJR3oWPeHPUaulm9y5H3a4/hSTqwQq9vIOwJlo4gSpyS9
U7cPk5meIsN0w0xPavNyM71qR8iNhz5FCmBnrSXbR3eaquH3LuZXid9xIzUvZPQl
1zgJoZoy+rdU9w1vX0l3zA1RwTadrIESytz7nMB7WXQIwXjSddleJht2lmfAcxv0
IBDTNZy0Qyi+hWbFA7Cv0DQ0SARaZrCLsB2r4ifusDxWDs3dm2jkcrKIBUDjnh0m
z432X/EJYb/Feijip34o/7Raq//srcpf+VS5LRn2l9FKcCN7UeYQLLvmtymBUlMK
UyjrbJz3fZilgf/L3ga+Pa39sCWWIx5ZTg8Y/LM5WqTy4gPOgY3/cWi/Q9gdcCCU
fxkPLCIrqoDgRyessL7BZ8TVOJnhSPArL/IeLAX4QmEUVa/CxpXtgC9f4rEgQZac
hRKIdKg7VxlkEOTFyUTe39C+Je83KA4zOj+iqPTMmIaL0njekGyAIXPujHBjj5lF
XFBThJviExevBVy9YJ0ekIWZFnEe7nYW5I68lj9E1DC9Pn8brnEbN62vlfz/6E/l
pzPRGJSCsp25Io23ZQP+QHjpnUO1VTr/A3oPub5hEYmibh7eRjbbgRf6JLpuNuXW
S8qYDj/fGCxrdHLpJ3/9Bz0F/evO0R5SlgmkDoUkc1YiCZrnU91APust/USDcUkr
6iZgdHX//lGkUl8m3bAu8QkvgRA2JcNbSD+WN/+ynRwY9Q22tGTNXg8HJbD0otEC
luQo3JDG5+K6dySuP+J9Y6duFlfSAme/hAgjqnX9k6I3IfKA1olfNTPDi15ZkwTY
f7MbKcQk8Fwgg/G8O2C9y77FrtB+pa/a/8JKWesNUrksdf5CGFaLOjsNXGlp7gQQ
4IOncjUGGSE61/BBmxje4ASJnMSqb0DGB/fG1gxeJjT4Z11rQgWcyU42UtTO23mm
whlN11ajCjf11P5xkQcCvdT3xAV+9AF6qqBAVuUAeyJZOrByupWd6oFo8Oi3H2X3
5nzLSarEvcfruTF0YZZMxvAB68bbJDLwKglncUngYiKIHgKwQF1nJAqpFXv6vMOT
aY4ow2uMCExIE3ELEm1LGNCLCPxpl808IbNRF4fcb6glbuAB7e4lA3c6fc4lNtF3
lL0De05CZfQkHlye4uF0lEg5idQCqHjLMoh3YxORiyp5jbcb1Xey5rKcJ9bRYiup
xJgurkC1e9ajtclYI9S9ku/kMqoTPFOfeNIppvb8SlcwVmzFHqmgWanFrH6zlQLI
58OWIkrxSusyN81pMy3zuf2diYAmOsWYFxCY4eeNAYDrFSXbcSvVnJooIhgDQeIp
VqfGFSalklQ6fKipVf/gMfKK2zRncrhXwqBLUNm+dqPewUgy0vd/9e/WirOke0//
Qz2ZSZLQ57L+Uf+zhoqThbMAuHJG3HvgRpgg38y0hj4qS4XltfTkYlaWqQT2vB+u
Q+IeO+LW4EnD10wxm3Sj+4A5gO3FQ5+H5Y7VqYnCiw1pNRuqh1twqQM4W8MU6F9h
ZZg7O/9T9UVU2ullBo9n5sF3mjni0QIvH9DBiywWH5Jt1b31oL8ayzKOsFgSbOSk
iemwo0uOKuv+6t5c8ufVdSHjYyQMsaXTz25dLbeDRzIVjzpoK7VTeupWIHYkbzH7
TrA56SuI8wx7MRAIinyHTAVioVTAN9md8HybcOO1Ha+b2wJIEoFznH7TvtmDIyGU
zke9/GHdC1y5fGUYV4acezNYac80LyI68EW0R+ig0QTD4h17hiIFaXKstJz6Zzcd
2fzgG0mVpwe0EtysAbLKrAjL7Vv2aZQr0UIatelsMyyMqOJ1NG7d4irSuaDULzkf
miSiI2TVE1gV+DPp2zNdMV49ML3c+Pq7XWY4DPF5SS8FLywrEzgP1qKTe3ysitGw
uG1E07Xl06y2blvOoQBcoCT/yE0j8Ly49tGTsssl/nVt06KhcysF2xnE9qnL0xgr
If0LhIKR1QtpqJeXhmgniyEt5zN9GZclpH8PwY0IS3aVuhPvEHgagYmHbf2r7Yy5
bEk9t1U/VLF59EIcoCpAkZKGkW9BRvBSekdPUdMuFtxxEQGzbgXGo3DGMgfK41di
UdATLKg9YXokkwVTn0vi8+ecyBbuXd+mLicujFUv1W51HhBJ73Jif7MgyfRQPtqI
3z85xuXvjRdG2YVhaA/fDbi+mLp21EVMvzB7ewfjvkwdrIv6bnu0zaj+8KEJiLCf
Ni9T3QnWySWMS9MSP6EkJ+z6T14Kg/wnwJ1lkykdf0y5ihB0zegQLfv+ezTe0p7+
GmW4rGmzQwzyfCTVcmwG1g5aZgwO2qrvOqMk27DC51waxCaepJr8mNHLCMbeP0Rk
7JwV3HbYdjfTYPRUIWjge67mHMU57N+zfOQOFgduUsAhnoeY7PiuNwqR6cugRYYB
EPVynWmQQAKQlah/VBXwoMUBfru/7xCGH02a3rYbzfsKben0czWCsJkd3huCu3aP
yhLcsA4+aRIyMNReP41pU+CTRLQLYmPA4qWb6djVOMoRTHYD3qvJUSsUNbJ+ZCmv
v6lIgPBtnXOtCgYfBtaZEM+Jt34P0jJo6u9FDEWDns4Ep2nXidknlHGRl2lXW/Jo
sk1Q+lpA9KO+uza+R/X6Ba4bAxBejrVdI8PXZ4VDjZl5KnLnyvG8T/s2QclbD4Rl
QhdhQzOAoCi+JcvZVLg9tMaPpGXiB6ZX8cO7XAD6VUNrpOQIuAmKfPvLijo6LknH
eRu95U2TCx2BjrW+UeZV1TRoWOe+bpX/EPwsoihfecXSoK/cQHvq6TqVfTOjvzMD
Qwr+NxMdQ8jFa0GP1tjcmrCQe50w88D3H+jVl284E/ORDazcVznXf+AdABtficqB
vX658Nb1kxFQ6q9IYEMpfyMohxk///K1bQoE+ooFaIvwjgMupYlwfw7iZkla+bPk
S6HkGFGZyeU95ZznQWC0BKDeIXWINL8OSZuTvpZCwxpiIJtPQ+T9pMv9+boH4Irm
Hl2ALq177xbKw9krEZdS2SgwNgE7Z0G45fphy4u7OW2jhJi6A1ers3ITdW4OchZT
DcSPTiUUcVe5WG3Plwa7bhFlnOR9eBl97S8fDay049NutoP6MDowu2H+uozWuceL
SI+8lLrGrTI20GSmn8rlryOfgUc66VZX4hieA4lMPfPpIppH+yG6SdiM9qlqSvCP
cf4zz6Fw6Net5k0ObCBYPWRvi1VfhfO3IrRgMRRSBmKDWsw3JN82C8xUasKs8846
th5WBXCK9QqpgPOVoKUBAfPHhQYzEKjm5HHoyVqcwvgsDuDcsxuPILsWI3OQFWjO
SBhKxxxJFy9WCBnHSYOBWyBk8QCxRB0NhREBAgO283FugMxysy99NUqLUnNUCnUs
l4Or2410H7s8QmuT0+5lTmqP1IPT4wju0lnxwLRpw6E6oWzXQrF1B4ztcB7vdLHL
qXjiGwhpMU8UCdudANkKYE5c/DnilSixlTfDfMcfUfzt+AS2aDmNvIRbGkpjaX3H
Kfl5HhyhnYhVzEYCCHS8SF+rJzh7AcCemUJY4kTF+K6Ti+b575IhZ/28SYEO7JLY
qH7fR1H/BiY5xRPfCOF/nfut1EDYrc5LFKoNkaQOhGJgYxTk6FfGOVh43Rm/fCEj
5dOmwLgZ4B5UzG0rxy0i5dx++L1K6yyz8ot7fcnV0aOtVMv7+1wjMgk3GNA4cvZX
xKEOLjePlOiddMA+nkwWmSqTAayCwneihl2sV3IK1P+62jGzDPdpKkbjBGuVRS7X
jttQpovw+PFW1KGRaWSOausPzFeNC4kKkSzCPrypFs2EeGAfD9Rx425xjYEJVFPo
WJMrpYJ2GNS7ZSwIAecNnKGUBdroS4hzFwPsUw3ZaGPpX7ISyTta/YrjE1sOYo9q
sPGv9fzxSCH1IKIcuZwGqQ7MDDaGZM8VFW9+UQ3r9zuNuOqyIQzMEKPrtBEqpIDX
F/W2Nb5PutGShG9ESpwv1zPNFB+LZYhFRdeVCqED2GLvUXjwLtBAtn0tQ4TGc7n+
gaJ2KfnBmtz67EnPDVnIv1uHYSmgFZdHaYPJR5p5Ald5aX3LrV03G7QJhwZUKKaH
Uw9WZGvDwzmF5wvg/UpjCHFLHH3lLu4e+tkq3At0odryKzk6zZSZ/afgQu1fW0HM
6u36fjdLvpomkhMRO1DCfeiKAnTw+q1+xQZDYtVNNMEIkFVWK3TuaMtKfgGD+yds
ZFoVK6FdG8atC/b50m02JTW0j5n+hzRD1fugtCDUkjdhC6LjwLmJo4oA4o9U4P9A
MJXUHjC7d/j2p9MMUVkAchN3K7DlW3If+rgmkhFuNFx4eMjZmcXlDRo9Dc6FXyQt
5QEPCIJhg+QTl0+yONQJwe65SkgwoW/7Pr6v957W9Twj7OyOucZAjzZGlkI/nELQ
hKaijh3QddPe9VQm1uWDCdHE5I5BFqu0tba9JIB5CbZSGqhcG4BsOYVovkkjdR7i
DbCL9m7iIJg2gy0PqCYqqwDHqzyqzokaEcFphPnb0f4menf4eyn/MvW+0fl72Chb
Omfg3kKirzdP1ou6uWK5OJLoJlHTgiu/c+qlCFE+Tr0dJEnY4pdaVYuGjp0dN4fX
WfEJK3qsSuwK8pvfIc9x5rWhk6fAJ1eGXmV1rd0qPVjXeHMwFKLHeXb/E3fVV77J
WEchOXZjIzR21qYk+QoMszHAZDGjTF/uHUy/QS/6IcG/10hz7gsHDPRbjig04yb7
PY5uj73dZVUjqDEsAvp61cZkMsgTxkjqf/Cc3aKrRJiNI9GmNWycXw8GRYlW/Al8
02gTGDB5X7ELEEeWeJqPalN1V9yyGp8yMhfocZTaD479rsJbCWRtQSHLl8ViYkW+
pk/IuUPEyoYEIciS+/xfChnfcI5ltTJE2jtVSA8/JgEpAwVwgzZOzKrMoiaaVL2P
3XKiwmUC6tSCrS/RQdfGLlZe1fuPbvdkNtQRD2HXDuhLWiDHc3qXLdHyJ1f+9NrW
hwf7ahcQO0J8uxkLLetQTTq9kPB8LgJfFBjYgOccPNw6aLhMarY1czesvFEh+fRl
VtEgdUtWnZ35bS97Dv1otb+mTapWj3V3BtHZSyk7/VTkMKkHx/579l4Bu6dquZFb
EPW7Y0qOaMt7oJp/UEmzdKETKvBuiTkQgDlzVzv8ZxK5aNP3zGoicB8FEDSanCOz
juIxSNJMCIWB/68tbqwhKOUzaCxUN7fVW7P7Y8VedDVlP06L26D2HMFUHqYJ6NkT
UZMMr23MrxmJbXFPDNz6kaf2RZxJ1NumeAuBoy5Lbmam7mGknigSrx3WWLdPORFv
Gaad9w0MmnQJ8nGmEzqWidzM8C8yonz5OSRkb8r2469wPC1Lg42ywuT/h3aXgDRH
tRmUgxYjOdNOVi+SqYsyCbZkoPs8vCZVdynR+Tb0evNwWO228hPH4UZLUezagqpv
4M1ysNjAhf9E0hR2PqIMokD4VhEl39udlShNVaU2Hf6hKeZzEiK9d72LFIFqw/k7
YFskW8d969X46qGU9uhx+TwTy+WPx2Tq9Nptst0EtVuioi27heQPXn9jxOddwxlZ
M+X6ZbzITnAj9BEfewE8d69XPHfjp+xm+/hzl3Wz3I1Nq6DsknreWH2IUQnP5XM6
6c/CUB7XzUwMHL1ZYfl+asD4Y+NcOgetR7oxyNz00afmBtRB9LV8xFyEFVtwJ3Tv
El77MueOoJDXSY1MIbTAmALjeCBnNOz3Y7GK/56og6caN2WHyaK98eNxmS8/lxpm
fVYHQXP1Xpd1Py50ccdQFOqQNxgP/XSzttV0MhwUk94A+Avzfgj2DRjFJxTgcuoI
9Xx0nsr9WAT/c0A+OS0H/V6WuhVb2wnteBXKDPEo5OBQRCCUNNmwjWrCfOLmYYr0
34RwyADJVpcV/6fM3v84X7xQBOMyEj4+5LLXwd2Bj1ReZIN61pIGESlQ15D1LwHt
nvvwD2ovzQfz98PAycNkZ1WD4js/A5olf6+S5owEE1TLkW4jfMZTzt1iqLTauCTb
6vbBFefDGZo8Zxttdxcjg9uH+6nLRIHTUWUmhMOLoSUmv5oSfx9g6IUjKQumaMmc
CWN36IbKlOhuuGBbZOGm1SSodTrCElwG06pr25VRDFhDEoiPzAhtqQJ4pJtg26nx
Ybw0V9jRH4/xkvc3mtZ47n4s7uwFidTP1YobA7UXAJey1JpzYa8JTS7lJ6DJbHIz
rbMKMzAeY8lOgnEsYS1vapCxgitZBJiGJda6PlUgKe42PP6JvavUHTUyjcqtMWt7
aJUt1LFwdzsKMA+uhLA9uca1ce86vlEi883d6goiDjLOxkDSphgQOd2cCJeVKN4W
XOSN/LNYSFX5zfAAWO4tEIEESI3e1i/P1nGuiSh9V9IJk3+JfWHaPO0l6FB0hPLp
2BnDu/CPQd6nZumrYc3DNaqAf8T5GNFBUFSETLnrm2NfjEv6N225puTHYr1xJfIc
jmMZnluwr4gOLfxxQNObgYrGqikjCMbkXhzVc/XGmqOCnEA6MwxJEY60NcrqkzLV
6NUhWobsyXwY1+NBu/0TzR0+edODzyLExYfJrT+8WFWmr9grmYhKGgopN1Jw4aD8
liSkw4U9zHZmhAi59IfS9KiQQXhnuoYeK0h1SDSRzSuEk2KrLQlDwExkL1taC2q2
el89ztu/GYnuhnaTe8F6+7fiApOMH00aQNGEz7R4LA5TaCYjC1UiWlArwCWAv+tN
CYhBEc7s3X/fgINrF8QZlWJ2rjy+VpQhXClKakWkFoqx1K4sWrta0W6EAyXxV+p0
2UOQOPhDmQj/GTHteD9euA0mGl3WxevnfwYUTEWh9P6xfSa2jhfvNpbnVopBQXS6
4yd/0jUj8irqbon2rdVhN/LfIXK0GwT3+xmzYZYLYM1ODVIg5dqTyD31wqTGW43A
DMcErnBP2yQq92jGh+pNHhLTlaKVA7cC4182OK2mHGEEmF+woHTSMXJ6mVKoBCXu
uIrT0hzLgbOyqnY12Z7FJJ0Ht58jsgIxk6BPUrK3JLWan8af3y5AKfB5E7Jk0vrC
mbXU+bV9z6Btaq4AE7fKYS10zJle/q8Zbkr0FaiLUxBap2BysjmYcqf8PDlo93Ml
zwPW/+SumCNr+Pm3Mwtp3T2G61ydYNY+Wo7X3/4dnPy1Rqtf260bUlUK4CYDU0u3
8I2R5uHjhTCICLwwVT8pSuJEQcbW0VuLO3y38KPQSMpaItPJnBPt2wFBfvfjFDBl
UFxPuVi7VB2js8eCcURfhVP8dd63cuFDP89VNOkeW09kcrOQnyLoGgkEcVdSEby5
Aq/3/HAvaMZ5VUnDf1QkeYY+HU6EexWxJzvJqmydqZeX4Hl+2lp9cx0a5Ns51CRx
Gv4L83izslF8BE07UWdWewFrnyLhejWfujOolIMAsfp33fMKT7kaTyICczSiadti
IWBHb+G0z5M2rbKm56FbRFgEAXPxD6NF4bDhEfPb7oDOU7kZRid3MlFFo/Efsawd
QaaFqLKaZJjVErLoRQD7qSCszxMvOmziM5ZCCXlbu4qGyuH+1rnIsMPrE2qdLbs4
njUfuZp/bs6Ru/R25BNoeAO78Q67dXBsT/RAGorknn0ccP1sflr6Z9QOKK/2R8AL
MZ4r9ud6ncIH2kutOy6jJeyUgTzhv5nqjyk2PR+J/vM8A5CkrJKd4iM1lqt1vM/G
ZXuW+6l5+GPohaF+fBjexhIXRDx4iTeoZyfXDoJE9fyJ5kMkTyJbNjcFl4lN3Pvk
OjxUIRs+kNx8REa8EXexo9hnKrlCRY1iMgGSbu9MBQfd0t3W7C6459I9SS2vqzEF
FBoysL2dzo0sVqCg4C+r3LB78h1/EWVSR6YbrJjfdbbRJ/htXNmh4bzNyLCy0J9K
XL2pco7lzCnfXOJRlhXXghtdrUORBlKDc0nRRd250bY3QQGOS9SCse+k7dxcgATh
z7b8iPmcvaOUrQ3FmrMcizuWejcaPHj0MJvrFXkFYcoLmeb5SjDny8YAC99V/bD2
SSc/Vz+fR9YSy+l7d80RDpyf9eEaD7Jbgduk3yrH8B64w+D7ovWklQrFN79QbK6o
zYRZq8wtGc/lQW5rGzZM5CeYJ8LA6YkBY4oygqAeM14tyUFGMQwQyps8KOAjhnSO
5sCKNsZsgBkcYrT20eVkFcogrdIvgpzs77JB+JJ0NVqWNsJ7VyMl+1wFIXncOMaX
l4xMcqBUqEckKd6MKhQrUfl46HHLLNbCIwCKC8PmPziEy+twIqeLHIw/ABa7xSPR
ttlyYo5gcdIB75SgvLqdobBI8X8Mw2bWELNXJwnxQ1KndknixDzTqBMYy6hgoWOR
NDTAUJHOrcBcb9XhHD/r7oej45LTFZKCnZMIMSgKzTEwYCnnrvjKMY5MIbcfkkjQ
4PiEDwMxe1ITj27IpW7afiQrAAdbLcM0QtR1TkdaceFikDeRyEVt4B4ZNcMlcHwU
kg6H5b1yMbsgu/V7BNIpKpoMuhitYJi1eLq9UaH7F5BhMIYYrqPDLQAOujoYJ7Q7
0sptZQl1b6cZxsX/tuyWWnx1j/X7NaXclIGDpeyciIlyI983IZodTaIn8VTdtyOH
5LQzdkHooueCcmbf1BgzjN0pcuMIKnETQSt95mwJesHEbX/AjpMD3WFwiC/udWmt
EpBBYxfDDtdFBMclv5uQZJeiNSqzOr7kjb4IgCbxKxcEkrmmLgDBU7e+7yCNrTm6
JijAGu1L+7ISGlegBTPOt7UX+iBwXO0R0UktROQ4Rp0ea+3qAh4kn25XOtgv6Fqb
B8sdltUO/S+Qt+X6rDed1665BG9oIy3yP6pHTFRsRsHywbTb9xQIGUMH/LoVsj39
ywTPgeVxe2Cec49rX0Wjff1rVtnOSGxBqkGucvUGNm7LvYaZ1NWSFDVNUS7Ryazt
IpEsLghJ5oRxpObd0Mp8S0Bg8mtMwlT14d9e4FdHiAI6LdUXHH5xUJfpqpxWq6K7
caEzatPm5Jq8J61TTJ1jGsyHVMtX9KHdpG4oagr64AZ+sZiMmeS3JSeP9BXuZrSD
jlb2wI/yEdHrYZMdlRuXtsORJcx/9y70JcV3Gf9N0Cq6SErwvUVycvH9w+x0aTF7
rLRIzTrBA+wR2rm0mN5kB1w4OxvH7N/Q6sgO5e/h9rnr2tSCDD0Z5QIFXSNva9bR
mgtuRUo5eHFgPcySlfeUOfLMv+P6k98v7pR/rnRUFNRMknR4Yl+tnOgf2pQHE+UW
5eCo8GZ4ROxLhen6duVcjllwX9whwYbn3fh7/7CYGO9xbYA4mkfEwU/qAo1m9PRt
jjd9Bdb7lku+JRQX4yb0v6R4g/iIT9Ry3Q5yBdrjY2lRaykfS7zy2GCZgWIqFNey
ED75x04tf/3wjETBY3x8rm5skP1KZa366pNLO4aGECujgIug0m5+NrWtqa6dPUpe
bAEz8um1PWBeBG5ectNmZceFWkwIK28AXKG8qP/aQ52JwuKDZPvChqcXsWnH6cne
2IYNMN18FpCeioBDyQjgAGCatwz2/CzSHaI/3UZV0BI6XYwj4CMltk9/B/7ubqqg
hZVQNG9LAmA+Gngs7EiLwbhtIfyHhtSkpZsDiTjsVVMyUnCi+bYFWtYzL5Qtlj24
N0omfC7Zll7E7zUULDsVj+VTwK1mpr7pMbkuIk6RIo/G9KwxzpGyfEyT23sKeDdg
OFjIa1jzd92pgKH215Yo0dszcGHB1dCPCpIk7kOOHuRTyGg0AYgeDQuzCXo7FFVt
ct/HvAofHt8OHTIJrB4AEMlpcpm6nYDmSoTj1vDfzwqpie5ZQr/gwVR3cGIGm8zP
lOdoNW+xAjarI/38WcztqHT/pRdLEhsr9T/WL0UcasCVNmeVxOTjjPO8JbajYclm
sHzWVy6zIycgz84uEzc8lUpHL2W7d+tS10itm/QbEYf7VqtdxAimKb+78CywEjd+
5NO5JLQXxMzx9RYzSsCbSkODA/VVy3pusmIRJMsJebyF5haO7EIHwveGs9G79U7T
D5PUKX2mBt1TmT0gjxfg5GYLPe86mEQZDjRdNpvk5e+/mtoXPY3SZCYmAAGTXKkH
mIigTipLGk/2exttpQXiJYtov6gz9xpkE1ba+akbzMdTEgJ5odwcFJEMnTtiRTjs
n2gF7Tv3+25kGPgs3Wg+3YRDduDyzonnzsd9pJ3pSSmzvrUdi3hYYduxA5OgqgYd
YEH1ylb3eHza0WLLFscDq0dfPbrOAkYZ/aZlnOVdTK9PHVKYKZ9xch/f3htzOMLh
nOWMUOgE9ztZ6Ll4h5aXdkn43p1NYqp98dnGjbjmoLp2zOQblj1ETVCcg6kMHSLT
4kTtPqNer8omsJOHXzPAeffAxZp8sOAtEODWwRIKkQGyB9lNLInc/BkZW31DSSwh
BlKbZBRPGxsZncjvd1AzvHcAOu5TvE5HIQfLrFc+jbu7vjB2NEZh/9YncnvZl8LS
+4MjS1GnT+YX9OqnLoUh/+nX8uDUxrta3TMdDSOuZ3pwLPhEjmGN257JSemaWrE2
0+NWP36+9/dxp/vXNg2+N6TxQJ1fTjDJ/RoupDib3zCd30wkeOlWd40hM3xYx+D8
hpjESvdrlVp1ok3aiU8UVVsHemkr+q64LrECgaDgNW5A/1curPl41WdvH6CJC7rN
9ke4vizeJFPDp9DLuGYH7XOUg+/CQzYWfCaPaUh8K3YyNeeEeOWcxl4CzMa3K44U
i8eWNHHhzv2QrcR17uXB4UF8/bxsQ3Y+nS7RAJRXhQLwvxcunMgYJxXhlxdx9GqT
nUSnGZsZh74zfnT0Qz+9gnW2IeqMyTy7HdUsKxG0KsiCB77SKa2CcTakyqX3HX75
qn8oDnIEB3ijwcjjHjXvS5z2hxcVome/5LxUShbWodF52Qd7EHlbXi3PYTEb7Bdi
VV3m2sHQk1yO275uT1Kd7RKvJi9NknhSBGd6N3I3v+BbqFTVwwLAwC85HNYi2jKR
njkkHaPQkj3IPlRx3yk/0GI9ZqQMhak15ApAlD+JRvfgWnAn7C7+PQloAC/ikOH1
Pci9AaxCsGM8+T2SaIVA/7pWSLneiQ5O9DxYdCOuk38itWs1lnrHd+3EcOPCMFCB
yFODBX/iLip6J945Q1ZoWrAODI89k64LzLx7EIZz82wxs8jXMNEKy+3I7Mryl9Iu
Cf8hWVSEXNSNfSg6+lpm2Mb2f6gKwlvZlU0kMaLIiRaAk4nZ/tHypT5yR1k80xFy
cmpx/2OOohPQDPilsahmL+ElgPxZdVV7NQru3cXm6IrCnf3cDMR8tXGp4bgePuoy
94OKBDugGboIE4dY0f6k+MKBnZy11r4ZY4ebzS4+7R1lRtGfUb4KGGrMyLMLfoej
vo6A5zh//Bg/xxA261j4uiySQ94Z3VOdLO9O41JqrpxXpITV7xU3qHYoGJ73xUdJ
1KMYKx2MCgTu0ZpGA9YCn4sky2RlQRxoh2uEbyRIbe+DKj6HfnsEM3AJsc9gzn6Y
px0bx/A40JvJVNLqlVI6fcsSiE9JTKEnpRAdSZUzgw19Ksf8N1sw0NxQ3xip29+2
GDV23NLUlatC4prOycRChcUNiZU1TCLV8c2e7YS6lHvoIX4Kqzs14aghyQp/k37y
vPAkIFVIz3IsL+CJxv0PsOLNxiVP8B56+LqECvNqXmtpUpyfSSPjrzlb7L6gnJ1L
RTiJgfzdhKaJZaWfW0DIsxSDCbm8yBQ7n4M/jzlf3oZo4ucj4/ho84TRF7fE5HWW
BFB/TL/jZa1ku5ZyOY/nv0W/z4f5FiVrNhfWgDOCpY2VLF+p8OTAUbMSCWv6gsb2
1gnLhf9ckvFCJa4acZqvsA3DfOh6YuNrNkTzyT9lrl48P+zKWOJUJPOHWnI714uK
WxVfO+X3bK82ZR21aqQ0r+3OzYgpziWdyOdqWbZRZ36z7sv6IeiaR7aLXhoaa2i3
HL78xfSG0K6+6WW46tcUvr2bO6AC4Ku5oJtyiHLB9KZy+N+33U56lMVlq/kitg6d
MF2CvmsB7TUi9Ro2SqNWuCH7/nh2Cekj2o3YSey5cKaCI6J44VhUk5QTN1ASUF65
3nrIzE2pbnY3eU36qhN/qmJMJcbrT/i5iFMizGQTAQ4DaVou5IqDQZumAeEVGIV3
sO46j+EEpdEjAm+nhOCopmX/mp0UBIXoOBMW5xz05AUwIN26cto4dvxiZOf63hyh
xfCpCcU/1ANW9clWIU9GDtIwm7BFF9foUIzXkoJdSwQEkXQGki2DEPyvtMytcN7J
3umtKFlo63Q90bhY3wF/vFP4J4X42aEjOmGTCH1tGZ7hdSd8dS19BQdmSpZTYXpy
FTNh6Ce/GJSC+rxvhzcPVVEN8FemuLEoV4rLj/3TnIlfiP6odcFiWfvfZf6cHqCj
OscqfNa5JYiXf2vlGEkzeke1/sk822EOYV0qKu8VXKdfJh6RuTXIbv77654dABOa
FC6ocSUx02SxzTq+UUJkNY5D33j3aJx+f/7qVUDRZxxjNZ5ig3sY1bu/cTY+RXHD
LtkF1s69Llz1Xpps4FPSSCCvdk/vNzX31n0DwyjBj8Br6qFHdITEbrlZgdQ5/6Mk
+Z7nQ9eIF0BGYnD9H9FgMEr7ODhD/MxE8NHqodXy7S8g/lNytSJPI77d2IXSTKwx
ZF51/BCUJfKhp6y5xTFq4DEx0hL3Mq+kNc8jHAbF4HmMFREGNPDWGkoM3XQTLCFy
aWUKlxPT5xS9SYvdN5EYNz/Is51GjMblVp+Uq4YW6GgeevVBfdaZDnKZjiqmT1Mo
DDBDDPsHT5AqvhlGWBIzo7cW+/wnWlP/tYMh7NnTCUjppWQs5HV4Mom8IJw5RoNS
pJdxhUx1TzZsP8qDhjw42wR8/1H938kmmvctV7ytY5S9ervrxbiKazi+Yfi1GGEk
lvvtRBn1RGgPMLHKVBzsbciG6+TgHqBaGh7oXpz5WAsD5GHBUkHenjpN9ksHtd7k
2FYBV+MjfLzb/9Xa9VV37pz31Zv1XS1wfPkMCBWtgCcaLj5E51AZZPcDNgD16DxD
IObR99C4qIF5gbGSZkPBTvmpv2ilLP96dBA9mkLV/rge71WeC1Bcmdy0hiW/Bi+m
u0VAaCrUdo/4BE9oTpASq3kptMqMBIrQ3tz1ZLQ+1BM1kTPiAkxngE0eHHv6SX+v
fG8dJXUGmnv+LT8WocgY6PLAEV0clBTuXpIcJ9ZBj0sDDXmxAAEY1PuhSSdL67Fn
nx64AaQxR/4KrsF4yd1HRTrJ9OoN4Hl5WtK8XuHUcYrVS0joIRbtKuQeoPZsr/r6
p0lThCr0GJuHpfTXdRQ4VCHN3i2qOKiWFaSFGgmV9uCdUoifGmasonbxgpEanyNz
2/rTPSROO8vDEwmVpo33MPjJ8SnloKyDOVXpxp46Lg/lmdVox90LilxoJAq5rM+X
xoILD1OXzelj2VtxNuMcHTGRODq7ez2CMR65exfHh/9XnTm4zeRzL/0e/2BIT/2n
HXgy+yE+iI5N04mzbEjZYFeiOSn6SVcF8XoE1BRXL6XbNgujif40paNa38dLZS1W
1RdBGfhLIdjLxxfd6vVxYtC4UAzieus+HMIbxaOZRNxus0b9Yba+Uw+MlrwWMu44
OiF+X7kCeV0isy41wMJujejWTuMsU38ylOYPvnIVax7/eh+Rfl63i3JNSBXz2jNO
IuR5gNhxAu18NwWMMA4v+kUv0SPC7iog1n2uSJQ1PQ/R8ipxppgplQGXE1wMumIr
4RFUpmhyZVwfI+UDzgvfGBgrqQY3/8mC0Sz4HQzAuUSCDbmLL3uzsriR170vyPMk
up2QI1TK5EynukV90wen5C6mKFmno7D+Z6kPobyRF8LdMdrVLRC2mUV+EMvPEg1v
fT0anQisie3wevrRVtPEpHl5bvabAmIJYadXIalYY8oV6MLNekdJWM4wmGXaR2cJ
mdvkZofbW5ccga0Es+tO1i+sAQlhVOHvcn1X09vCTHBEtUJsqSBw7UcQFMGlFW5A
kLZOR6gGItoHe2bAucnOmIPaOElLamRDC24k9M6A1LblI3GzZ8u+C2m2qH3qe7As
sniadlPBJ3HPw6JNu5d6wJzedHslCza0jYSTPpzFMNt9jBMHCW6rEtohi1AWTPfb
pgGYZV92MxVpEqopFlurD22qfewyKU/++t84dua0CqMNR6xGko8kSnyrTFJSVKaB
30+Ak5pTyscIqJhvZCZCcc74SjqWcba7ISFnWJkPiHIQBN/Br0b+35jEI17qbFQh
jyR8n6SX+jUyO+fvM0asZIQGnlz02JFMhdmD4wYlHjkHRYf2dYWK8jT6OjqalbvH
UkyjtyOsl26q9/BMcsUqDszqYvNMNHQS6U59uRbU3ogUSyE8AbqPV5XrykErP3ec
eeZCi/jHjGwXBhB7T8B7eAm71ajFaquSOM2dOFak6h8/FTf3WLskiSN7OpZ/qP3n
wEw7SAOPKgUxdGXOG2W0J3WUEpcNw9REF1NYQz70kutbbEX2ZRxJrbC8e1W9Xnl1
J0YANuSG6mJJSGF+YRknaaXKBw9VyfkIxjaBKUHw2tTfbb/iUXfeB0LO40hmEfzA
efkoRtSpeHgIlWP5jMNUmfZtFHGQt51G4uAdGfmAxGllrgel3J/8wgARS39yjC96
smeRwqmUm9EGm619W5/sClmESNSAkE3WlkTe1UGMvMQ/dL6FwjLdX59p47Xljmoz
huAdXt8fY1KsK3N8hSNZk8Z5Fj399M8CeVNyr0xDroqrelJNpvvF2ogA7+XRFv48
tFEPLValWM5jbpWmCC8Lw/d8L2F/y9A/hiYCevn85KFPXTSGkKWNR+D7a/wcjnbv
HAWJw9/aHlGkPS5mxZrsegG5iLazz2ZTdnt5M+15Dt+LeT33JoPYGrdD9B3A8nfm
L/a6toh0I9DIIAL7Zy/X+drTLmInDNuaqLvypWbQCyZ+pZ2iqHJgtT2ovKW8BC6k
NwQu9mLftbRibtdqjcQytMaL9RlGrJHrgYFAaUOiFXdHwMC8B62LGL7biMr8oepN
YxDD8JxtqOHbtjopoABC/+sVyDVL7n0UPysNpjcFnbPrgnwQlahySS61C6wI3Gni
S1Fhkim57Qa+xw+RBLtakZnj2/PmblMqhmf37OoYaqa1CS8oic/IvrxE5LYry449
7cqiZ6n5KiCPKMgyRQM69rJHXMrDeh0CrEci1LlDRFcfOXbwMPrkNr3kujhiKC6B
CVofEDYjOaQltE6tcF/qamvXaHpFyG36QwREgiHo1X+2O0eD1d9XkkqWnIecJfI3
ZeTyPp5ywFLILOHlfIzZqP/2dIdPLr9qrvuC17XJjUCz+nfs+L5mSV2rWSOABW/r
4AyZMdQ0pgJliXiDXLb8r35MmPWMS7CN0FdsNiDNWegAXam4tu+12ZxuK3T1chmp
+VR1Gbod3CIRv9i7g/G8IO8H87jqTv5JJmvkW5RzBlPdLo9pHlOAuiLdIU5BpCCz
n0t/Grkcl1Q4iJhzYN0E7lh8RZsQHfRO6tnkcJ03cre8T2Kdyvx8UHUcIkgdjjJ5
SmLvj76/Sg1j/IdrJqF3kyO9S30m41zjERqa4rDtKLve8L+0ThEzW4s9iQYW3Itr
WFiKNupahYin5OVxgNC6j6OUmCvY9shNGVgitsMINFMsG3Xn+lNgpsi9jOa7jSHB
DAAmObRbJC4u3tqqINcPCnC++0TIKZ4rr3hOllUbQDaWk9yrUliZDXPE0Asx6LFR
gh+c7Q3svo01mlG194NyYf2OcJBn5jvDWtnBHajaX8yjqwz+qX5ETEMz8krfGIAU
xASPiZh8O2ovW9oNhmWIba/B4SaEvXUrIThsRoBTEGAmbcT84XmEGYo0OoZwfJ/L
G5xsKYvdKJ2RsKUPrMebkZJkTvLTFkdFCr+uRxSChPEwkovhUSHH6BJZX+/DUBIj
WGEF2z+uxsOfneZEFzmQhU+c4YsmSFI2Uk3Vvg1aSIltZ/chbbiA50PpPuxthGTQ
8Tu+Idr20B+7UeVV82vO9ECOSg8BW6IIfrFFz2ygxu0D96Op5AspaupvYnkXqp8e
MrcjG1rG3/5EI9rvQwRoQd55mUzke8UwkrwJeojqdUPhMvOOhnd6V4ukWCXEBsOs
/+6muT4NsTWlO7fs3dB8IreAaOsoqIsDgFM61MZ6OjvLcRa3wbZbwpVn1BLe5bCt
VQabJss6zrrNNNxVgss0Xck5XW9ZI7IGR+6cjbGzoA/+3TUnAfDqgvGUtT9TnDz9
Gdnia0J3btpwQgGB9tVOQYJs76ZMkmWcVhSUdxwu2CvMi3qiTCW7u3+mHpOFSJRj
2BNel2df/C5cqoCWjiROA5gH7vv+bD86SWCX3y/nriSWij/NXhUMWwJfMKBN1BqQ
33TZnrtFC7TMNYDywGw/xK4xqfNtA/Z0iyXVbxwoSvsTf/LArDUEf+hLjAcuXPju
OsY4Z5T3SIKqmtJyu6XbWmESQtgLo7zSBefZH1knUhN2JWK5jCQYlVL+x2USE4Mp
blNUS8pkJXpOJnwaIoGgh2EhoTEF1tdsgNjV8pIv9QwA6m96CdIrYOpq62xhWsev
9GQ8Kgk1xF9GRc9Js/m33dAiEBo5RV15b4kIufFkATFU3yPFTvbLKpbK6njRnbTP
YHtAnLL3K+AckGUuAoQlfXtU5XtUsFRQ0daBXhJnptrXRp9laND++vrAt5RAKTmW
XdV+7Uce9yiluJw1LJTTV+bIFISJ9SYjywqDkeIBQqk1r+r0GI+ipTZJOqDCF9PP
bHUVyDfWt/c1vqingUjLhg9JaHlb2cyrCKbYtlxbKcsGEOGvOhin8GInbYt6ei5p
NvTsdhUYRb24JjfAyAOZL3BGNyP9UvWyHUt/88TrGl29vDG3inadRAEg71xEkVpB
krPfzeaPoNs1fQ2Su78pxmX+tm7imNj2hNxg8tF05igJJsPkrZBiQqFA5ECb3sZ7
CgI7djTsEx65t2uE3+cFKbVXeoxceJIGgcw/DoU33LrjP5asMh8ps9KN0JheQPkH
ievUUCzkZIFbQPf+AHMg6uYXEfDig7CXqrkox8Glf+QY0NMPeiQIqBQMejthxmiY
D1DIhol2FWXmJ6j/+KMfiwKGmak4vlVr9/2oSsT5jFFbNPV69CBevVFC+uoBwRpJ
PjLjPLvQzSkply1JmsO3mW38EyMZRHoinwx+PXo77nN8MMzoezTUIos30MJiUqHl
DsvxPhSyuIuLreyYFso6hL5+A8q3MrcTB6XgNdGpP+FTlYI5eJXSlobWl1mlzIb1
x66/LL/YWHqxOjO6a5R1u9seEwlwoOiPTUV63jQMTltmsnwDfjYvqCrX6iLpqJw3
0f8m67bJoAL5xKXNdY9mjuevb9W950eix3T22Po0lcEuztdniiGDPHcUQM41owHe
26b76nl7+BgK/6mb1JO/0joOAa/cJjLd6x2ODfsps6U+6AViJ2i5rtKxHuu71Dj4
l8NgrWhcR7ylSwRyjFNV7VoV9NEP75T0MHo4icv9JdYfNwfr7HNsJQ40Bva/mzrn
LMYqB6ly0copMjZ5FV6TPicgHlosUG39wZfwMHNzIz5yeMJwCW90WFqw6U3HDEcD
0o2Vmo5cPkuHiiWZRA2xidzxz4hKZlSoZhOWmhi55nuDtte8hMhiLOjebd8GS8V3
/O/LATJoZag4LbtLCeNe7R5/upguNs1mpdBGJKCVPu+jYSamVq3XpXVtTXNOPt5z
FfBdjLg2ijO/RIgugkYPblC4ZWiHsYNTXKOIPaCveu2TBwonJsDRgxKiRX+r+dA+
tki+02/BqKo7DuBnqHwFIYyOfoGyT/kQ2jEmCl3zBTTY2mpeNHVHs29qGrC7CMVr
n7DJk44Qdtay1VsFNdqH3+LoNLVS8EPnbmoZZdyRlJM1lAVkYP7O8oIqxKR/K0v9
kELS/TfBdJgB4jBLrQWYjzTGKB0FGR28G2zOFsF2DbKxdxMS/1vDddfNvmYrIcvo
4egAbEQLQPd7DS1rC5mxESkvjIwPsXoxjHslpR6v3YcYjjiaApfmKmAw88KiQOk9
Z5ZBOAqh9c4nVWGhNjB8lvujo4XhtXdLHcUMSTNnNepRpAX73whnuC6ho8w8MJUF
yp+2/SIGhCvA9wbrVpB9vUliT37tGaHKEy5ASLZcNimaGdwYJgyomGR8DqlCTwMg
bKrJdxwWuYf2jMJggko160YR0eSVAZyE9HXqTk+z7rnk/0mFmI+Q3mM2zXdIIDiI
a2wgTwONJyA66K47Q5PAb0ho0sgiZgzKTj33z0Dl4vlKbSYd2CiDUhTK9jDM4EF4
DiXKy51pHMVJfWScUqbveZcnNbj14oP28JqfSdko08JcrOcMGkQsZJzcvcP+I7ZC
XPuTDkUsCEXlZkmt0A5D0zhOuSUKvxd7TFrAV/f/FH4nWEH3riBMWc5nlR/XsZns
Pr1tV7J4St0uK1rKmkFxlMq8/HTO46xdexKO82x6DRanYePwKEFFw2C2NzmzKrZh
4BKgNN5y+Re2vpDFwRDI2AIdl0FtOMIayLqhYUXHs3hSVGaZcoOMCQ/20mqwt29S
2VEjqrEuK5jpcaNSli3P/pAu0kzNUHWPxSSJH9vwVcaMunRmuOhydt+RAY3P5QLQ
tHcvihhBPxHh8Xl1OfZBqOPzNAt3Sj1X+2eZoqUsB7ybJ3oOx8h+FEyQ0uVujoMF
y0VSRWVqSZL9LzX2Fwl/7vjjmOc/tRVCwIJz1KNWK77DtSNXyjtc2pWsvzGmyP2k
ze7Ai/4WrnnYNZwqr4Q3gcguxB0m0wjsb8euYjpOCk3kdq8+uewKeK35O4A6383C
BsvJsdeBhXj4IIb8NS15qVx/ZM1k7720WZ3PFUu7FQ0y62FruJsDMTY3DT0KrmHq
i+7y/d8A7v8LEt3YeJ/IuvF0fXJnRj7vJ23I8GtndVOLs5G7gLJGTRcbrWbJhlzH
0ZXZYJCO/RuD8xfcpKawOW3KvM/aXqUVecupbgEw/P28lB+62FO0HnL9Y7uOA2a5
1nGWur34oUQUmf4FOpSAmB//j0ZDoNZPe8Mfb8h00ofRpw/mkIfo3jLIwho64qgm
ZHicFMctRTwh8sNeiTHalpIyYOSYxlq0/8fqDrsxqJTebGBrFz0TuW+4Qngu1wRJ
zYqArT9534h5W1c4F9jzoPGIbHJSVsp3eNZNyBkfPKjykdntmSonA1kO7q5GF0V1
nhc3VZQjmKLlSc5Uas6Vt2dgPhraX1th006q6pLFJP22+5NZs5ebEPcfchxxerFn
4bNmAw+NiEsOJs1pUj1oYukF7fPd/FbBWvuQXi9vMV2tN7TFIgeia2TLeZmOSgJb
UUcSHjUpvI4gnw19aPVu/qCnHZMKLG8ozVGdJqrvvSSPnN5Bqc1jpWQB6uGA52NY
Ny9IVUckwy9NOK0yF5zBUo/HUN4hgtT3vfn53vrAyoosaJBzi3952ydBwf36Ptwz
NxStkNFpV16ehlrz6LCOtLAUz5OAnlUa8JsRUouynDj53MxIFRULXg9U5sW4b08b
L8SuGQEI0qh93g2a2/q3LbbYiRlTGLq2Yov7+TcA/r9CHFyGNPewhnx7UKyKG3cv
GWnW9FJTmEty8CdxCGZFSfq990EKuQ4kLqKqoICLICeTf11n0bj61MaKbRc2TUvQ
CQm6HeeHitMSaIOPf74Pc8dD0OPgkxmJPhgqU4/5AouYHFyt1MWzposGStNupoaW
Lfx3AmxQWUmc6pBrVo3Dw2KKV99vnzKCHp9IFcak56CKM8R8vmtzJiJW9dw9lXC7
oSZmhhSJFL3IvtNMfQopigFLoV5Nn3J2NR7hog4Tl959SjqKp6A3E5gDUGvzR7lG
66p2oOEsrXxR7HZ+vhcIrfoZ7ALmeffTvlPNvKnYfApki4wLJ2qyV1Ymf3gnIltz
rNLOB6XwWi+1aax7xIdcbM+01avupcmdvsDtnRUfpSs2pJpdCFdUTqt5xkO6oRVv
Zc0aGJV3TNS9edg2qMfpMj8NIejnQv1fIR5bbhwxoveh/Os1Y8RM7BTlYggHUtGF
NJ8s+YKc2fzkCBKY/iLy6G0Tb+GW4E0uBWdx2CT06MGoeQz2BizJsS0+Gu77NIRo
T69o8uMMi6tu7PVCjrpzG1AUOW4SetHFKg0mON8HGPphilS3Cxryh9STr4lJe/GR
0S73Mb4k83CaIlod5+YtpdR7N5zBb/0oPs/UqA6D6pQn2wJamOVedHBYYfB1HOjs
69VVlNM8vvf/+iCvp9OE9bxBhimEQ3jJKEDuuaJi4QldeII/7eIH3Hj+GmpxQ7OA
r+1XF+DTVJPt/Ly+5IUGx12WmY7NvlKSLqgxUFM3po3OsVVbi13S24sacJJyPaeq
YW1AsU9Kjr7abIwy5JRJce89M7z0VlkXBF43apy+bTIRLhUnSxzhSlDYo29Fi1BC
GsNgSZKsQ3CGpVAjfrh5Tte7v6S48Xj+BFEbydwsXBj5YWWQ3Li0bOwCgKaNJtP9
LoiL3M/SFAEJF2tIVEwR3zvUUuuqyKqJ/+jbl5kzjYZ+WvqT7hEADdbyX8Y6Vmne
CoCmNk+Cpwh45x59Yf/zX5LLUMNxG+lR7Z96wuV/Aqb4bAnA9tjkusdQMHANfRAK
ReBLDLMfhDhU93jeqb/IdJ9zlKlyCwABE4cWSvocXGlWS26259GkE9QTa3r01tfV
TiFlOEsbW+vv3Mj+5ANG5IAzSC5LCC3C4+7PrIcfaEuBdt85wkR2CMy4x2wQA8pa
VQp/g/8paKPcqqL3GW4zGaX1qrZwa9aQaAnUAK0rjVCyoy0PT7uUpRfeqK4eYAtx
oK0H2sNkMljjS1zLfxaprfyj+sKO3GCInp9wa9m9BoKphhHYtTPDnmHi3Rp6JVph
hFiFChpvFpyXeZiR46NCat+qpO+AhamqmzSdDzcLZ12O695G8EduWn4gEi7X35IG
tgoJAcYg934+0A7V48MU9JrGOpNUChQP09kS+pyuZKyyoS2uQ0qlFklBfwVJ71ig
XagKz6RkHNHVEf1k+dgD0XGq0el6thEc8/UcX0z2zXELcVT24Jj/yftqKYhq0Al2
lUgxoFOT7k7/nPExkOySVhE0aDK59k5xAHuZSnLK8WpI40XjfMM3ZTdaO1Y6Tq73
tlEXpQunqpMdaPD82AcL6rCtBbCZxFlonktVN9zk/Om7/DVMhJRRSP4m69xPMRXP
fxdO0qkpYTVH9KXlAElI9ApeFEGxzDGNW6sMiuWR3TPVTPJntNPKeJMDiw70LTMD
ggJzxOMS+idUUD3j5k/ThQQLOb4KDZVuPoMK+ouaOUQN37YA9oBb14dAd2G7PvaS
pdjNJE4vmKxZTS1iAQcog9QKm2XD92w5LX/3+rpJUPC9kZmycmE8+JKoF2H4N7Ab
pKEiOBr8KaXrKh0S5tYKqSJGXd78NrN6OyywASUwTrUHKtDUwnCc0M9DnCs5lWlM
Zmg4Yx31GvK9zRJoTuT1+9b3YwCV9Vi8IzfCNxZoKZgz7IzWfj0wz2XjaSWHxWo/
H8dgqb61zloYVXMnOxaGzVWDmApmyNQlWQr9Iq13uuY67G72CDWpSnh5fOa+wXzG
3CljqaPGVDK5VK7sPkXos/4KVtPkEbROyHs5xjt83YM5zmciBo1DckaORcCSx02N
Lx7KK1Fiw+kVTG0v0Lvx/yvgkQHBI7mVqn82WIJtN8TTLpLRRZXjpzfld7vQoyRZ
wQBon2dJzMP+/bHWJoKcvvjjVRSwuZ8u7KBZACKNASNsuFYEmApcJpVjlt3GXUVZ
70HMOrsJ7ejdKU1k8zVgcRhotrzbzd4AG32DgdNiOVho0NYZ1CvQakUVvoPKwyWg
cAt1Mq5a+ik6IVl4RCZWm/gn5pwCedqJvhe5DMX8xVFjA8vKYGqhkHYewl4bfmlD
6s8ySTFzYwLvfPauZpQrw65+jNbyAEZjPlKSUHuC0mGaUj29ZdvEut3wOlZZxvw5
ey7vVDNPwq2p0ztxUdL7NeTP7FNINKxSPff6+/G/6sfPjQqb/YJN5OWyW1ymm5Kg
0EXDQVTbjfWS9EXC6AAodbghdOuY7f2PVTnluncu7pyNubRi0NRdo7XIo0Df/BfL
kQ1XYaTgEMbf9rHVcC05Djdc5R8aO9KV9LCLdCJYkGDc+msCOz4XANGqeqhvJg6B
qJdMJkq5bRyjPpGg4qAsF9tweJMoBVR7fHlJIuSu+qjhRK0i3hT7qeF3huxxqPTU
DAjN2rTe9Kl0Ax7i8ybY1ecNN2P8KLraLAjEGFrtOubhUtdqxNuvU4jSYfqmEQNJ
y6ViAUY0IOsaLq+fcIPDRl+c8MZbMFSgm/xoUnjmk5d3UnS//Ryqkm9xcIBf4R+k
dbKNLBMcJ5un7j/3apRo8KE04ArzaUguKmttBPjpSRM7jbJh6Qz84Uq+ksv/ArGB
VUpBwKmY193Z+MNZwHntKBD6IgfNr37gQFIQxSihduHQd4v7iI9Gp2yHe29Ri77F
okebEu48/sG92U6D0LImbrEEYh5tnCTvTu+ZFHP8sYnn2gllQsF5Tmjskfb5lMKN
Ae/DNLUkXlx1WvDc7lUO6Sn2eGx7Cdcr6WZpWjc3s490XVyLqM3wY1vDUz4IwAh2
gueHRdbuYRaJkaTjGF5zDUMe4GDTgYZMkhj5R31j4HFMywAyW8NU3Jpj5fvswwzk
4TEnxHwlla865VLzEoZzX8MVcW2EdHuxcG4YsisszV5iwnTWS7athMH2DdBSp5pu
C8JDmEzSM83S0ZpGd5gebW+kNVCbhlJd2129HnFxEImqh52s2fn3iY8p6wh81Phb
RTQm2CiKITfvNL/fdX3viLmA+CX043lrEbZVdDokqgmWeFQMJL9uqBiCrPA5D3BU
neaJvZ5O114z7W0RKNyjrZ9INQEnHwKJHzuIVlyBowg8Ka/5Q3tO6W6wLL5rK8Rx
FDPMWMeV+yXOv7GBlENvjf0tTJef9Sw4P1njEUk8yDMEA/r1yJ8U8Nne78lkm0Jh
NzbjrNDKctcTlfnnaI1YKr1o2zwCenMVaEN5jHTcl279f/9M3Fb1zcKboti0cgWI
z+LEY/WEdDI7cqbEOfrMyZJ2QQYZ44sS3GmVpQVSpEW7Mi4Swk6hG3NohCvFXTy3
NHG6GqhrJ77JalOPfUvvF2BiqaZjLztXijgxhVchnaQDze9X3CdN1YE71GozCVKp
WTZtZT7pBjhShjaAdkhZ3PD2/FTQp/oX+IiSh3G0rh/ERaHo7vpL8RzIh0n1qLPM
kMWacZVTVpvgXJPqU4DUTXwjBdDiSzIeGJKT8l5R8p1E1Im558nL/ESW4vsbfhLu
8Jog/EOw1oIvxKRPj09iBGC5h2CcE8luyDG0hhQDUpCNe+LgDhM1YwnlUo5WImwe
SC8hZ2Vgop/RvVgUGyrcMahHdEi+BdF5LKwD0ZB2c7ePhrbwZEP+q4OkzXBwuZ0U
A9fOtF5DWBIqPVH3Jo7vPnAxjtBfbJ1A3iUd1oBY8rzxDzhckO7cOKOzT9s2ARl9
BIV/1xdSxShc7uzkVzgWlanm8OJg3cmM4gxjt2N7VYlnEG+qQbW9avkugNvmxZj3
yGUX9lVD8dWX0hsKLKi0WFY3/Eb3jlwX6wzzIEIrgM2s83C5KjdfH8oXUWDUE6fi
G5O3Xj2NMZTamyyhZRefBEtOhFwAFYZgE6d6G4QM+1UYHMJAJFfVCFFLIldTa8Al
J6aOldxNE+Wh/AjgDoTsUjZX7BYc6SX/DfSqEBW3S7+S9opYPJmqDATQabsTQPyH
ve6ZHv6BXxmj/8HBi83qwsWrhX2VrBUrTY6sA9yQ47ZVOwVwOLuIL/33vdnQIt3o
khXJLoE7VpoC1exidpgLZl5QYXuvo8jJVTJuj3PwMO5pVje/ufR78Y8YDJQY7BI/
yxlAFMpcD7EIoFsxZ7PH/zs0bMkKx3vVAlETR3jmsa6Wt6jlxHVEgIgLu8K/1/cc
EdL2l49li6PFcW+MTOOE+Fn2E3xle7Ode+wIuUOpA5Way5zroQwvpJKjgxeGtCRC
TyARpEOZD8pAE8KFZ3kyC9C28AHdXhzAI0Ss9fyfygK7MOAyYmhh9h4qNS1uJWPW
ZnhqsswcoX+X63TF3yi9a67BLDpCWj6E4L3m2UW5i9bdkjaVztpODJuVYmGDrGfD
92tKWVL4GVY2lQykwr73RWtqSBJ3WvCzZ9jg8iuCqJcBMEKk6ksA/BYKR0ncSyMn
2yChIrdf5Na0RDeLluHHFCUoVwoEuhzJpsG2wdDMdJZt1ntnRYmCnn8wvTaQvIzQ
E1YH/m3KgwobuuOe4GWDltbWa6mWaQapDnnTtAkCRiB0JpQR7vx/QrPIhpJiToK5
gfHHfPdGY3LJCg+nHI18PSlF7atzZecWwb2zBY2tjkZ/AsIuNrp0VKG0kPrKGXsI
uq2RLS1vJuhQIViDM5H1G51yCkTDfQNFZpdkzPXNMLJ5FELdXQOOVp4Y99SgwBtR
GAiWazUNKWw0+FjpvpM4d6M+qdglmY51HPjphAzybOdpIQ0SCoIPap4wdY05oJa8
tZWd9IQ01wOjZvIeXfxHvpvg9IUOcNCsFQq/dBWto3B/I/agqUdSq18bAUr+/w41
uvXIbS7wESm4cBTXBz43UC+2Ku6zI9T0UqoIqZqwb9Wp+rFPLRCIFSLo3FhyxNzH
b0Mabl6akjxXPR9AWF4/ILPicjMhCvzvfKFyvurfiej+qNs2c8NouR7Zp+dOUsEb
EoTCj7QoRdSRZaalf3ys8dWpWIzWJOEAl4NYje9Q9N2esi6wQ/lcA+eUwx2AAYY/
c1HnIIu3UegtfEbCpUZmm5XFfsXDtKWT4zXL+y3XEA0oMJaTwZTz5KxI3jD0/bTz
49aGDnqeAORkoci5NNQrerUUNTP8lvoYRrPPR/Y4PwkKPAg/jiLwZPtW1YhrFndg
PZJBtJv6D+0U4sfl3W5TqqVNrF3tA3ye2j10qn2losKGp3Z/mZ4lEBqY5c8PaqVf
YnZ+v3Fs5aO7B+rT06S9JSGYnDK4NOtOr3m08IMcW0oBabYCTbm7CH+UoFSAI5UD
T2JsHlGnhZ67NZriMjzzoJAtmoOvwrwHS06mmarlDQkBC7oDiMIlXmxVH7YWix3u
C6Iv6sNyc4VSrsnTmpiGI4GN+zFCadrg3iVPNbx2EYglpSS478tCuZVf5dm+o8Un
v1HS9C3BHK301Umj2OLk6u4ICpvmvRBUjAH4xME1xf2YOKzBhe47GVntvCRWIUDA
TaIwviuT4qLJRVmdJnmUsHRrrREVy4vRE7YbD3GEGoSN40ngVRSn/Ig6djK3EadY
QTRhBIzJTAbLp+Y6n9sIlFSWFpBCKaFMobDycyeS1KupXh6WMJTJTEhnM3BW7/91
jTh3b1CF6+VS8kQuyTpbSsnCukPuR6CSGjJTPtfSUOXT5KHE30UfBG4Gn68oMM/o
8XsiuaniibRLm/f2ZJ3+li/pLl1XwgggnoJhpfJ3cetrHcUAKdzwimyj4dLpfpfx
Hvz7pIzUt+V7n2IcjJWtbGn7LplDOWFhuB8yBO8F84lIIwlqJHE7qd6UJOxSn72d
Kc+OSYbtFRQC29pf4RN7/PqHbk1wOqkuOYoaUCFFEe6vZ//bCKSwRrE4sZiuZY1e
Q7kL6YHsmoiCBq0rYO1vJ70UByWpXl5J2voWY6Uz02uwBzYdDT15srxeazWSrUD5
Dj4U6KVvKCuDjxvcWLyEguY94DS4oSvmL69PjhfAd7jigtGeLHbDLTs4RbnQdde1
v6DhBzX3FLngrUQm/bohoc8EX1GDeGDq3SnpIhIiQNg7LLOzIWhj55v7d9iLtMSp
DTK0CQjg/TCmztFllAGpKT3nTnYEQA23tvIm+XAtXNpkI/YKtHNJVAU96aVvJmn9
n+pj16LmrC3W2984tL9T43ufuqn+SxDS1KyRmhLLGdeV2iUug9js1ypVrAWtGVTz
kgBZLvrmq/lJhnxaw1VgivTSxZPYtNPF/mWBke0ZJLqt2ydzb3iPscR/MUVJ9zlK
tg8Nv2/+AeA+4h/W1D/UPd4MjULLsHig8YhCpYxmNWkYZ310/137BGATzalUy1Yz
+SK+p5kKs5PASqOAWjMpF/seCPfxmZDd9MfezYwLnBAMTCqilhuMAaCyjHHRj6aZ
7VxsG2giPnAqHtjVcLCgO3Or2z7M8d3y0dcn8sBvF7pGH0Nmk1v6mU8O819G3BrS
tZrGdTfpgfgoFcNRg5+mq90CyT0VCNJYc47I17NJCVpT92zeFl2wyh7erDeFEfx6
S6lyaAc3o8F71FfwxhLJEUiD6mzvRwLXiHBEV/YOaxgchmVfYJxMPGCg42Y4uyy0
kMEWkf2JQIGs53KY9yu60zaSq48nQcockW8eK7UsV3n7c7yDROzi6PRi4n95jbY4
YMQZNRGrgbbhhCgHtT3RKP51mKhlsdwfINVZjhAbGpl4sCjeZEfQFMCMSiTm8EU5
batM1kzIuYTTpxDCQ5/BG/JyOBfOV/V3NzKmLPGy7iVp0KTYHSeh3jday6meQvM3
tSU9oJIcEaY2cwZPW8ImysoCBu+KMWcpXCE8uOUO7J6/uVGEd/Pyli7gEnjCh7Gi
0TmUh8XOJUNdk80VUBkhi0GfMp8lcu6iSaQgFt5czEjQtVkn/kN5kmWp9N2RQgCP
mpDfoj0YzPreAzOUe12L/rn6lvRtzIPKJqOmuOVhZPZU2dTfhZI6vlaRMsH/inuS
giOr2PZ2YNmWA0ht4umqwh2vLiFyVVfpBLpyzA3WgD9Zi/UQRcoBurXTF8zFQtcR
QvCqcWSEDpki9p7GZGJugv85ULfqGpbDxf8bDlwXZt+oqQ1fi+sbmBmdgkybeIMw
2fc0l5wFr9Tu/oS0rKiTQyPIBqLciduM52UbGtxssd8xrvI3ww4zme9Ny21OWm64
SDA0EIskakpyxalv5LB6vB2JGw01/UEXvJuS6ij53va3ak6gwtHL8GURMJMAZtDV
CUx3sl2cVjDtr12/xrDUsy0f52WP8MUFI9/ANpPWOtzEa+lfTdVvbp4BKmFIm1pq
oQ6lsENmfhb9IoQ1Cl7/zweX3q0sx6GPphdpkVPfKYdaE0nIms2ExTPaD77DULRY
JpKkD5Ws5hsWALSK3xSMjCF6neAqvdmQTxXkTBoAtB25hD86TGxgYSVw7TXLirOT
PYdtxk+FPMpr+j8CyBiSY82Cgv7Dl2q14cyjn1QJFsNAXlikgVAnz7CSPIWa3k/R
nnzxqjpQgg5EWJBybOlfjstisr38DQc54L9giO8QvXzeRtYqAxXB7cD9OCyMR8ii
o0g2OGYuF/N7gwRBwSSfOmEu3jJzAGe1j7srl8sr68mWmGxZVNIAwGxm7oYzAdTf
Hy28wVx4Z6dtLLmCRdyvY0YUbNyzXZ0xsxdlCKRN+56nslpKUCMitvQLCX+Tfi68
dcgxPZR8DTZUXbmoR0LUo+O3P2Vz8jldX9GXFOekyDFuXjDQsJX94KLASjMr90kw
Ryb6KSR8p1ZS+gvvbtI6e0EJLNsJfTw38sYT8KMNGJTi9RC9VVHoF0XCyy9wURqW
oSueFmu91XPSNW5O/ElRN/CCfIk4peh1ku7W0pBBfv2c+BohYI0ewyaut2EGvCAp
nLb4zdtHEg9pkHh0JerYiKjLBJIJnNlln8rD9nM4JVFXfvCFr6wb8WtBdrUMpLMt
Us4+O7ef56QJ2AcEFCkID/MgmfAVM3q5V4IcWpTZqm7HC3EDiC0La4cMF31JJKF+
+W0HWvWDhbVV8eSHoqGYNpn6KYiQsAVrkLkWZDye12icWf+eo8e5euvNsidpB/ap
T68rDwONCagpazV/kQUu5Csxt67T5pktfDqcxvXpf27Gnptkcmm+65jS71aOLWKc
T4nhR21mHffyJ9K4yYz03UdIBGCcgM/h1spk3OxXnxIHXuWCGNqw/p4kg0MNDZIW
4nmNhHVkdD7khkdbilEfza/oWRVpGZedrwP6oigaNdZZP+3riz7iEYpRBGPVB310
wrYvyTetj5wPZjJ07KO/9YlMtvQjmOiHln6kSHv8DQcDKwtDPX3aJeQGUrk7ivBH
LVaJIDGUERsPy5Sc8NUFmR2xkejRiy44miyhqbCB4KgkzJiCGwGwx6ODUZNiwfFh
tFQGiBzVgOmM+IEBPcmwudVHhLcvaPfPLUT0xxpOxHj6ceRSjWsTormhVN/lQ1nx
5acYtSWvlC1myO0RXXZi0blPgqQaDiV+bDjQpeng6w96gqBcMMk2wHzDEyy5Jvbg
3RLi/KcAX0ng5X7BL+mzC0RVw5XF6FycbgL7D0GVnuHXY9hgbI1T2Cy9KH0ny4qb
V0a9MqQ8MxeDNRewcDVrkI0f9wJVbUMR8a/nLWMeYvQ6fshlvRB+ZoelA4xqcT0f
bzv/MmczB1oqL3952zH2rHdgTHbZV2Pe69Ia8Ry7gw1Kf4z8xH5kEDfB3ZHGYKZl
W4Q1VJVF9Dfi9YNogQCREQTmYODFmQV+e82PgwgoQclzl+Zbaqw4KKFXL6KNaiwI
qsOxiWZ4SJ2XwYyjOQk6AAihmmmwdNN+FskOD/H28S1W3YtpOglUHlezQVyA4zNV
zStvgNJLZRq0YVqWrCs9oeExT/KedK1WwRGgIwRZmRZKWiKTKjAnMEqgnoAqrzgj
ptNSpOmcxbKpPU2S/wDBpkbKoansoySEHhuilzwltWLjSCZgNPmvqNljuRCLUTVP
jneZG+NpimvW0VrtJpsfGRZ3AqELxZQpNk4ZwHJkom3I8roNcD3r72vWjUCVlLw+
r83MKJ3mgsMhMsC1XASKxODDvHq5fNHr45pKFg0rJsidQFj1o1ray3s/B43bZjxW
q985NzBZQMlUY9NKtqBMZMdBLddqyEK/qyJ1NBpsTDS9sfakKxPGaq23A3DUj9i+
voA8F4dfGNbKWjzquxBbrJYBzEAePdubqKBebQgc0d2siNFOWfK4wfvFK0blw0RX
3EUYS9X5A+LZTyZ8Kuy2oxrFXzKgKlSGGGiHPMFRxkzR4fheDoULt5HLyd+JVmT9
bbSbLaGR6iSErQqUbbruUhWZ+zgKXppsyW/aWNIK1xwQbXMWflQWNN+hkQ0FCFjr
1gjC3UmgjNNCtZW8VcsMbcCV+uFk0PUDQzt4Xx9mBdnZFbRE1ItqCDQEkDvSBgJw
KCysjG0wls7nRK/1wmQkTEU4mv5IlT4bZIbturtriIbavJrgCRgiKVDYLgJZX9yO
K6JRhjyYMKwOKCaYknrvleVq2O40FeTRi6I+TdDsKiYhg54YaJeSayhiDLtlXlkW
WjehCPZcdoq+GSDTLMTb+VgEGdBxb73lne79kHfFbQk/n9dRK8P1BhEsYdY782QF
GK5koU+wUN3gFOVa9haKyU9Q+vMnIqe39oa6BgdaMkptGJs9UgvYO/bGYjsbsB1z
aFeLc+c6ExRmwy+l3QxLSweQyzpvn4aywNvo0CWyexkgQmDUOcAw1yt6m4kl40s3
/BywoJodkjbk91Ck+tliH6Wz9Bzr8iSXKFBD3+o3PTbm020VTDye2kBE1PqMCV11
bxYOF3jPIcNG6LnZ5arqZOyrRfD8i2Y3hAi9/xNEeFxdp7b2gFukzhaBuIlh9D/9
y5Y6W+UVfwAzwOadpR4oTTI491udyGCua1Hpq4J4knJuA+SZJwqBWGLbYTG3uewy
JtgihFTy+fuHgY4iu5LaMC1gKXrAgcjYHPTy6wXKt5q2cCvJQtS3rOKX1rMCLthQ
pvod6u8jtf+QVc9vkiNPTSwo66C1jJK/81nDFt+Uv591/33NkFuT+J2Pcv8UX5ry
qiM5w+GvT8rAA8sNiXkQ1jbvSxWcCCQPjVaqCLKOlvZ03DwNhz9vYiYmZ6tKjeFx
NGlgAsBCodlkq8y6Vn/pGLS0G4g1tOLjuMfIhtiukt0C85wA7uox4/P8AP3jzZ34
oaPcfgg9lA70aXX6jO3wXpB82wiFldV8Tkl2ImxK+dJViK5IgxPmdh7BmlM0MFt/
ZRkFZKyJTyn4OI9/tH1GdP4tWdcjbDjPpx63K5pYPRGxlOTXBzT2ggkmcxIP31OJ
s1vw3jUP5lGKDH0JnEmv/1BquZ8djZE6CR4xu3v1ZwqbErUO4x4+M/XuQGQvd4h0
V9RnCdsI2r6swuqIJUHFHMO3B1s/KKh+G/3LLL/t4/3FNTRQEWLQF8FJ1sHi3BsG
qcJUQ/55etakV8osh01HpYTJY7m3jXBfFfSg2SuSdk9ehgNWHwWuTdptpgPGiI03
Fu6C7TVEIm0tr2Lj9Vn97MPyayj8lcC61RKxcaXN7I0sYdLcgn238eD0NcKrrZQQ
aqPHW5mY43SZzuRYW5v5XmeNWlSD89MsOTcZes9qWrB3SfabF1SkUaTXhasLHHYq
slR+psT72ySDv++m5qZRRWuM5q8h8WbUjAYBZXiN4MXvHxvLoQGZhsH75dR/KD1i
Lqe1W6tOBY/XJseRUj6sGQ2P6bonqrkzd1HvDzTw3fcoRDirM0QWs5icTV+UwpWi
fFNulMbn5+Dzh1B5243aFr2lvoOhTr30wcNhdSZS+MAMmrBRTVzopT1Xh3Eigyc/
gqp9kG4TYTMVbFj2eJ8U+eV0cnwmLh8w06RwOPY2huDcViLzt1chWkitE0c+4RLE
s7t3EN5aYjA72bcfZBlGEOYj+wX7zDTzi620/aszbCEcrCjLfxQETBFsyzjgts5A
JatBIqndO4J5wQkNF1olxq3hn/d2MyTzhQEWRf7VecSP3/z9/4ajsxr0IsSH4MoP
X5AFPJWygXPmhHttNqXtuGvsnLt8pk3BpQsH50TkXgfQ/U83B690C/Tembxr14AX
F69AaxENj9Z+zG4wK+FDvcMHhyCVC1TUNs07d4L+g8107YOIqKjs/2/IOGfBOe2h
JY5YgvLWUq8m8rZ9LidOA+URW5RGSNnQiX+IO/RasdZV+7IxNvf+S+k9uzK0Ua5D
LR8fo5x/oHX8E3tV0Xe7tzA7ht1Ffdv9sS4atFuOXyG4hAd4WLWc0/6KFRLuNUtA
SfrrTA6+mIXxBvJ3QCRmaLK4HW4uzMmy6mUSkxgOLpgoE+fe97BlXrOrauWUjKAE
7aDCJuu+1dZyfGbV6sKGyTVzI9Nqxw9Zdv9n6PXxwSfD8lSeUOik9nC6Oglm73X8
s+zKm8mFzLQR6fC5KkANAy+hOX109kMMTC+dqqZ6llCw1tkcZvJXsboGJRdAGa1C
mFr2m9Tdmc4eQ6lNjfGQu60D+LBbQbFikO80QVJulNiei4lyJX7qFtwJoyKvq5H6
pOAfFWCYJFtNHe4saym3dWf5M3t/vAy+/j4LC8D3cHI+RsfqcLc051escqZuGG/T
uiiZm4/Y2twRWa1yi1sznl3WqKmZw1jtSE4fkKMhy6CtKVLoJJmlQ9i72dQvRx5u
rDG1+W3yhtKv0kmtjrx9wlgcQqzkbQgzXQbn+rSLDz3cCR8gggwv7tz0Ppgcd7RL
d/ekfD1+VzqbRwl8trCEbjLC+X6X19CXvhs+nbvts0sVowQjv2POm8jmmzRBY4CQ
YQHYnQsJCwJnZmjWtK8oERMwyxuR0dvriRY8rc4W4ozOLAv7N4Zxn2fTBABtcD12
jZz369ul9PBDCU+EvvCy2tZkp9RQRyzF2vzoAYaSeSHzks1xmCYpjOoHVHd0l2Lh
ScAq0xg0GFfPEFxfXdmAHv8dUGfbaQTaTLjTrPyu9+V69VV1wGEMl4fqvf0oEsBb
XJRTvT2D7YuFGVW8Olrgtbd+ldbJV+sUa+zxfJh1w4+1kRzZrCZwnzEpFzh+2Mp4
RAIX41LQw6iMsDcRcfD0S+fZ4C1rDeIO7qPfsOX+MWpsp906HO+GVHpr+u9FoUPt
TRq8pAGWcZWUhNfo+a2Ji0K5wx8XmLrwH2QMa5CEf6VrQV/qFWoCoGVe2pgmle8r
TB8YNzkKmZEgejryihvu01r55mkibSdwwt6D0Mo3ntmNfI2xcUa+VKd9LS004JeE
ev5Vfh6Qwzh2Bni3C0plRRvwdhaQaK5NM1xv4KBEh+E82Y92piTlx1cWxpWUS6yh
kvAzRhsp13Vy1b8vWXDpogQeoow1SnxAgcVVGyxRBlWfNKGt6p3IvhPR9lc5xelh
2nbspnTMb/uBuShCxaBOQxhh7+x93r1jMZj9Ky/RLnb1HSq0z26s9NuMyElS/0gI
Q2X/Z+K3Lg9Z2Ox7HZUdJq7Yo2GmoR3c/WhhR5x0G42KGs8hYp80s2/3RViyrD/L
hIGqczy45+vms7COzhaMCTvoW3nOb9zc5fo47MfviKmgPdePi29pgaGonxd/oFe7
qfzltMDeKYAT68fSXb8nGZHUx6naC/iGVcZWifD6sG5RUQUkbZ6jnGlu34SsAO4K
Qv61xe0/l/RRX79fiux9rWw9WRp+CQsGL5pC4CC+qHGvVsHB3c7YNl/DhIFjCVtt
MRN/KJjQWNdSnxMavTDhVAa6Tejp81wjl3XNHAQ3nixJjh/OpZ+n94uLCZkTO1hS
dFMvodx8k03D7x/v/XN5xQRaawmsFCb1PoYnkYJP17StuTXoi1v3DHkvH6AAxrsj
mmNcdXcv6SRJh7PDxqgnoKN2ppnjAOXiT5jqIOkVrYdSrgxJY67axFWlMPCj2O1i
zhzpiL1kjCbW/tB39hTZvybtCSy5wfhtt+BSb09fyPAEqQwchpEt+WuJraT1vyjF
jSOKjJXIqVCp4girCae405ZRq1oGAX81iBjagGOgExBRG3/dvt88+63Rt7pCfeK3
PZPErfYt/f5XljbN0EE/bQw7JkpTK7LhaLqD7AW9U9HVjWAf2YbGuDSkr39e/0Ug
e+iyIvlgsnRJViIlu/yZTPxGlgfCZi53ev3djd1NfsTsRA1vwQkriewicaJdeAgh
WXRH+vKRzlog0Xs4yMFkOZURou188hikZQ/7SEcVTefm28PLgDXvN3fsFTsmsG9c
Cl6im769FZ2jTIPYodu4jdxTqO+apUxsZ54rUdx1k6uYgcvUi9RcPQlbB9LiLmtL
eHw3TdKFzfomGJXNtoTnV8ZWjM0PrZZm3Pi5piuYMUOIFupoS6dgYfALhItuVLfS
ot0oq1bANew3zpG+YTqc1rrKvPH+XOXM+HcwM0kubaDhD9OCzweKTYPtOThCcWhO
oYJo8YkBhUjb2BGH7L3Rv165OV49O1cKWRaIfXGV9ZvM9xybeBzW4DNUDm/DfB79
I9t2VTwHuIA2OyjfGjCl9QIs7jbbmECz53hlswzSy5zx6zg/S/Mvx+2xDtT4mqj8
nPpzzZ5yxtIx9jUSBFzxBGPQtonL1UTmuXDBbarcrlYIeUe71MSkOyu7qpOm+CSG
ynAZuHU27zH9H7mtyvQt74lYD82jtDD8Z6dwjn9PIQe9qlApHUTyNyZxvQEfJgDj
WSk/vdY+Vc/U2S2aySfYSGDwLPx1QMs8NghM/cjeMK6a8kf0EyiuQXtPj2tmvowL
OYUfdy+zPR01vYY8oXUKfSxh9tUwkAqSJjspWxFyoDjnIMSTBJuepj9bM3TSix0b
+AsVa709AgjSWYBOfzYji8y3hxnmn9JSQUsMZLZmAs86C3XjxvKDgq4NC7duqTbE
gQ1U6TfNKnJuL/ujokwM4Q3DdIRwEIiP3SeMElIu2lr9ED90APGptbx3BfoOGoZN
+KUn/GKlkOci8+c0FM2xQsLXjJ+QmCf4KzdjaTgorj11ts5CMv7+a82o93lxJog4
++IxQl3iBLsS0sRkqR4kkAT9HxpLYbTo4yJzvcTgWoni/dE4G2Llrqb25a052FLU
lGNjie5SMDLii3D9XXn7o8HMqUOVlWBitVagtNH/WAZ5CjzirvImqyM6z3PY7AUl
cr5gCZDkwf4sutQBahTjuqTdE5ZE1WUvmOl4ZJ8vpybbbqHsQpfj2ER1laYzFlmp
R1DDUtMlEoGf0aanqJ9vdfnMdwcg2rByJxC8mJyWG+Xh0TQPJn/c47ldTkGniaq+
ZA9PTsVg1gMG+T8r6nmxF24AdsCKVv14hf3VfbkSDyGyuG8OjIDClEc4vD1qc2vJ
3wWhA9usWqf/cRXr6UHn8utQ2XpINLUO6DWX8je5BQLNUAagQG8oU8tIAK8/nSAj
dlEqkPaUAGUG9JDHGYaDTnscGjvmbEspFG3/inSn1PkrzVfpu2j9U/vfsZkkZCGG
0TkX0elAq7x89/nahmzjuW740C1MaRcMUDGNSNJwaDM49bbQ57oa3fgrCPiXYvKv
qHggye4AdD9S5xzV7JhjZR+3Pw1Uh9y28ROC+StucTBngs2gmFklwIfmXxwYbsQ4
XHu24JQmr9vjwsl8OAycSY+KW18umKQDCLjJObd5nbWutpvyhSpae0SDjxIq7MpB
z6CAJHIa/BdYB+Tz+vSILWsq4SfDmoJI7hztJKWs8QRtV+41HRn9qXHJHkIYnfv4
yfibZ6erbjFn3/Me1wekSyASQ+XRSkFFlzmsFtqiBALZM6m5goKbblyLISmvMyva
fVB/PIJJtnMz+CPExfk4mLT0Yk9QcoeLhkc09LjaUf4K4McLkfscKRVNku/yhOUt
lmiMRQvkq3lLOuiM7X8b8nzoD9VU/n2LBOANEjbx4SCGFtqjDg806zj3KSXUP+xW
tjMT9NVdrZgc1ePz5a5pzBzpvLgN/qLAhZaqKVwQvB/urzB3p+9xwUkV90L29Hi/
uzZnNsbAfvEB/7E0pkNJIiMbOHqa2SjnoloNQqdTd+l7BmUHxetvv8uEbnO+A/Ha
5gI8WdPogVu4FvWgyaRtcBIRyvGxgjePt52kpiVDI/yVFbBwdcNVY5VSxzM/8wTe
6knQSRijMspVcOE4cl3MCGpf5WNurSRAkK1PDE1MX9nUEDtRZsmmiOWnzuUHcQW3
K9lG0qzZD6XSAAMHKDmDbTlcKtB0a8a0EGIf6LtTF6C30ecxdUFFip+lGrrPFA9+
XsoYcTIomgbc2ft/IXhS1Th/Q4A321v8ueJ+2JbT1tMH4PqRyfsvl0Z7PI4pbCgS
iOjcgBY6qf8R8vR5Huv7YBSDoEGy6PDRNB2aGaaUWKeQUYtywS/6IMiXIxKs1Eyf
mgWmUbtBFqqPopiZDJ5HWasojPNZl40Ok5Mlyk2aylQ6oQ/Qvky+SNWTdMVtJZ6P
rCYEzWRRLCu3ML4ppuZrctMVcORIPOA+z8pv5jR/R6C5NsfTqBGJGSia/zhPO6YI
xrEmnvoix8I1pqLwS/809Gq/Gf6tzwU6NaaOwRyoj15JIU4Y0nW03ecph9v27RgG
+MW5g1nLcl8p4ZbMep0Lin2PoWfDtZrfdtUnSVFlYOZm9r1BvsIE7fj0+mAwV6yl
B5MZuHUIozg0CcbXMa84c5LU+CaXB0rhUN8xf8M2PNLB5MV0D7i315a3b1+n5Wrw
D6wAg1bv/Sb0pmmPIcTXHvHXit9RjxpgConfXLkVRrA9Uhzhd2WWlKd8DnPCaEoV
3i1rGMc/FGZze6e6nE3OGB9rV3JVneuJCaLwz1gq7rAo9a8cV/i5iLndqHqlkWO3
o9FPNSkf2KzjSqskYNpFAmUPLN49LCJrdd5bMs6gla2sTnOJUwesJtSytHqpFpM6
Jr2EhpzHTpRnkwhYlUWylA6GJ14ioD6wA92FOetxCOAdolqrr1lFL4KkxN3VYvm8
Jm+ToIqcyF8BhQqavXUR9/e0FkhVS1LuO2D7OPmkFcUY60aSnoKeU7KMqrfl8/PK
XrNcBheonmk2wrq6BOfN5mFk1frPK+qhaLfG4m8Qoi6GeMToxmWNGxUuyVkWnE0f
w07BL0ux8h4psqe/f1kfyjLQ5kN1DNqL+1c37+LERUiOg/sDuo3Ul4rfg3pD2YQD
dYvM6xfp08aNlkUmHquXx5m7N4BimffRdBqM4MazKO6qah784CneKCwks/SS67gT
zneen8oR/WERqf/LiPGbqe+XPcBWWFtQ1uhD1ukDCS40+cRNYUG+JldqklOiwGaw
z60jnMe8AC6DKIlNfD/9bVnvRNd2lZu9gwaMxi0U2caZi2u9me3xZl7hEaGJHfEE
oxNtH85JHyvbV8QBPDjaqWZJ3t+HlTqy+0L5soD7ih7XanKGy2uuDPSCp9JuuyO9
mJNgydYNX8UeklxoNti6aHpTaDlwRs6frv0SmFnA0OT/YKRQLg6FQ249qRv06vl/
luf7biPi1kHlZUjLX1IWrRXuwV4s+TE1ouyHBQlheRXkcBfL+UQL9ShOs3mZMht8
gnpcY4WUyIfToDhabl330gPQEzOBiU6rDPwd0hXEPfeVMme24xTCKjhtvug70z34
5YsqqvSSe+03t/hM0Q/sUPQ2Mik/g+2crNPkPeM8SmTRykzmsxLMfowmhffbuCvg
9lbs1ugATMCWJiZEVDnTeUZAXDBbG4CORKXnieKaKVm9oMhr8wLUVwtKcIraFqOp
I6HRqSwNNyTVO7l/ZdikgLX3HBNOVTfwgxOjmYMFtuwMFM2dAhFbukcyz65mLxGS
+FKttQHLir0H0oUYjHQSfx4IwTlkG6i7n665whv/l0ILOr4vLASJjbIbF99rs3m8
VoNKgMlOs3wIcC0xRtBv++Sgee0/fSA3ZiLp5C9b56NsURdkv86FMHhazB7mg+Xa
pq0ugIsYVdYkVNRHIwP1PTQQLlTSBzSp9oHCda9civOl9m6FHFEHShOBBrrmtY1/
Pfd4WdwPDY0J5ODQ08uK+alM5QnPfz5+jpdfXspa8v/Tiw8PYhMZROatsWAOrtlx
6gm6gJPgHz6J6popC41hEdv01eCKHn+zQbCwPyw/MzyrmvK88gyBqkH5K+OE+ind
sqyBAosutk0g0vjBkoHWJ59ogYaFyAbCwHN/FOjQK+TXGhgZ3sFQiqZ/7iXEkSw3
JJk0zU0Kyjx6GtUpENUoeoo6NSVSEvCO1PZLvc5yIx7IlBxbkvY+9cki5MfWWDXY
UbfIMGy2xooeehTo7aEVH+OAIcUFH90x5WVmohYOqws+zgS/jFwsvEBwGJ+1vQLL
jNv0/yuBpwmt9jcZQx06EjwBI1wUl4HnCvHz8bhNh3KbGzF+Tn6wKX4N9w59rRUO
8543JryHQdUt024a6Vwkmp9sC9Et0Y+9Uf6xfohrMyBzPNysJeLb5R4MOB9UWbCM
TFb0k2gv8z9Ic9sNppspyzIthqH9xCaan6DiYKc91uLhMGOzNhcFqZ5qFk+dx/s7
CzZL007bkwHGHfdLrq/G+KCkeYsXwlFt2YhquARJGIaMb2yzFyV4EAb/73+DH88S
hc0BYaPOpSvwWAmRdk/HNe6132sf+7cbZRlO+RNXfnvqMO4UIwNoapMKPSziMWvG
IIYgfW1ia0P6ibF+wyKqs0lYk404Snx1NqjO+K9/pgjRDK0FnHlVbFToSg/A5F+u
l07urjTZQOM5u+y5SfB9JD0Z0Ro42CRrXV3nK1oWcygOeNalEbgpZawcrc/ftxdz
osHy7R5+OdRD63GqvZuzGuQDhN5fkJTT63BTPRfkZoSaGnAi9eolGxNta07smNF1
z+Wv1md9Ve3lVW9SxyxoZ6Psg/yknLWZtDeGXgachgc++m4gkDMWOdA7mgh+21Tw
41kA+nzPsnST25BUH2S2A2G0nxh0Hu2P1F4opdCud6aHoQ4X1IebW2BRT18tZuV1
MpoY2tuVktlj9s0TgjYAco2AomLGeYHN4K45/vxNX8RRwpTHungOdzUNsua1JXeg
fAvQKxdS5u0lBZN5hLlXZ94wYoP2Bplsuqmlceaa/mW4jcy7X074gU1N3+QnaHR1
EruqxyNOIWdDAZyCnYFmhowE5P0QMDH4FhopiREGtxQnKD7B9ByMszBC2kTJmHsC
8pUBV4zu4jD6JXyqzYdEsB6Y70tv/mc6ddXkzkVgDqNaBqyqaKhtFOz5I5CoSfWX
ssXkbaozzCYj1u8xJFKUC/MFK70nyC4aFCn8rjb7eazjPN7WlIZ2p4C9noQc3BLS
05txlj1U258sDbUAQ9m2FR8OVyJMxxaEJBktCEdk91hrGSDugL4gubLFuZhkN5g5
bgyKkw1vr1FWkheJUstmhssbD9AG2yiv86R7ve6Yq/KhsCijMrp5Y3vXAqKkok5n
vmu1ZRErHvXZ+Xyoc/utp7/mWjMa/1cQRN0ZbOFjU/E+JLqqL5gZxSFl4wFpqLzT
/Bmdwp+GftTHCvhdjC34IsKgJfTCzj/ecdnPiMrtAwzPkPfwIcwP/re/ijQBBxQq
DPNUBVY2O3b3mVikwFYpeIOLCatOAONpKP40SsAoKX08uVUFySZN0KfD7Jpl4kvz
N5yJexFtPlX2xxHqTvdzvPAt/2dZdD3jXHjk0ZqM1wG31eLGGOuttU9RtFqaUoxX
IqXzGcliGEwdOHzu0xXgfBY1nf8hSd2YJbqrU86sAQlgRK6n+8pfN4CeVFWQec3x
QlHD8TG78KyxHtuoj+cifkhSkKOUCrybxNeVtqR0Ck9D8Q2TwlNmpEWyWurjll/U
Hm3A/HQwTniH3N9YWEtz5fBIezHdiaSfEuUqhlqqXk2RtvxswzYPVZbYL0TXavRA
g8gIXRRQefphsdM4/9zLca2caCM7UyicQ2tK7udI5PUOsO27C63TONGN6kKh2EL6
L1Gg1IXOsdtnUjfzSY1S3nx4xfip1aSxmYNy4cu6I6Kzfh+YVt4/ERNgKGAxdZ5H
Y0DSO2xIsEf38vXn/pt52mxmmqpNFozCsqXjUqrYEZCT1pM80tq3lLKe9NcxuHyq
0s9Mq0BlaMF5vluCpSZXiyjT1fPienKdWcwlIF53spUhctPSj9FZQVaZjPbvTs0d
Rauo+aSsXJRgMUMqq5rhlE//zY6i0CwLBehZLqZf+g5OaS2oveLxliUbiQ+RB1xx
5H2kDMgA0blrftU/Oo8EBcfKfK5+D7IypYH0JAJbgNN4WIL4j1c/DFfNHDhd8GPC
jxLAnYt0zWs1OWJtQoJQZF3Ra4HF3fwtV9WYJ+Hg+CEQ0qeO0QqU1VDcHzSW/NsW
upsBtnwaMqrKCtI+nw/GqPt1Iea7C89wOhjr/hTlFw32R4sKreHhMdIaCFMlFMfZ
pshVx7J4DYTZa6JOsxooRdDUPmZCf1OVBkeVE1otyzUFWnbujvZg1aUGs7GO7U4h
W9TS+EiSPV37PM2q1o8MIcG71IEhL3/eF5I8/gf+/7X8y/8bEKsDCWFrapHcWi7r
nDRiEE+U1QYx11D/BnDiwZcRz29IcO2fAvNpCUvR2yVfBsXnrO4FiNIWKfmF9Fb2
fJxJQT0Exo0tz/eL5XlxgzlUcAnpIpUGB4ku3MlLdt2jJwFcFURQXduyPfrK10kR
xh9wVR/9UKCqU+SKuqSdzQfGKQQcdOiZMG7rOgRXNuXccNVM2N8ViIlyWwb4u7QN
aunU107bPyMhJGlriHYQv92LVUFGqssI+gC3jIcyVa+Jxxs4i9ghWJ/U6mdQJehV
w13TrLwZX7PvSQMQgQDHAVVlf5ekfAwOQpi8ZdmzxuQXlLxHZOS99i24yyaVkMkU
Lh+Ps8HmIVBCGdUp2QEstyh1LgKIRt6zvE9Q216RGVfSzImupbNUK8BniP3x5yiV
AVod/lNgEM7VBeXMrtxPkpjOdGKLh6HY/OT7B5VqQfus4TlUg/U2q76hFOFUzA7Y
4LiGsVAvS2TTEkMmE+snajmHKb+ykRzcdp+X/LTBc8vYC8RYiAhsmcPXCgypEz6u
0Vj0X6Viyv1BhkrZn2YC/tPqoRjaKStOpGblTnB6Bc5QJLJXmqLA4X9HnclSehI0
OrBb9CjXFH9z1Q1+JXi6AIQWAvipxsrN/uMRmByHeqZHOiwrYz1fCbTs7LLyEI2I
WBmiyrHy8Wa/MLX063Pk989GhQXak1C4dCxos7TYw11kheeeyu3osrWA77bQtrnS
Y08T0sUULXRBSm1e4Ktew1XseaphcOgP/Pi3jhsKJOJM789S8POfbEzRBjMLe5IV
ei1NTPaTYqUji2OS9L+/PfwZu/NLiJsQbslCZ6U8hiBPK83eBEE3NQcP7MC1dOUn
pl2ZUELuVNd8C2BqqPuUGj3y2CzYanCYCgBjspGvYvh5+h4er80neo7iF5WsX2VY
M+yLMNx5tqUdK4o+UT13w02W0CDAAlJIOIZ34g6OH126ICcyO8nSI4yTvnGva9UR
pQi3UFPBD6Lwjfj0on2SEAzJ4Pu2ygtC3vi3j5pZbwgXnpyiNSAlYHDl6WsxZn4Q
ATT6rmwyopKBdMFF7tZ+KuUTr2xWMV5ajFiLWYWgyVFVYv0uv+0YFKXBsvGZNT4o
CR+eAOSuwsQDufl6Yyi8VEND1q6qPJtJOmejFPQhgMIWw0CGem/ir5sJm6as0Xg+
Vgx5RJISP3VYsfv7rFXxjRpZTmo6ZirKZxUS5+aJZd1FFGrvVfy97m+cvyDOyfHr
FOAT6mEa8Mj2Geu3Ro8Uq2edcsW9pxDRLva9JnovOcAAGcKMlaA627bv+CeAVaIF
tzFbRiEyu7lgSJlrIpJKO6H47tOWIuoZUOxr7HbyO96PDzbbO/evJFeNRfTJ20T3
XfGgX/jA4hmPs0GpaY/cYRdgtYQJayOW2iVaewFrdjseOmAScPEXjCBjZb9L3/0r
96NAvUKFdQWBDjTNI6NbYB9cxyZWj6Snp1TeUJ1NAsrdD54PDCX4q/Sryck6vy8r
ayCY/LWflCYsPAOuDWG4dw7xSJHcdmVM+2qtKpwDHCdlOR0cag1RjtYTqwOd3R6X
1p2I2u8BmHTL3l4BvjHSni/2GHXXI90Qr4Y9fgTOIltorSP1jnrKWsm9J14sZgMl
7VRvzoej7ozPBgks8q+RRUxgreT1fpxto968MQZLh2LbBSPMw7aYBzQouEVwZkoX
cLkkOiQIBzZaAEHWZPR6pI30n5jn7BUk/aV1kf4xHsjY5a3AVKQnxwvJbb/QVf7n
ZVohZvaR9fra6opxeRJl9FcxkPsKCtV1eI8qdY+7As6r/J8DYaaFLq5M6UdwcsCZ
gvILRlimVn+HV9OE0lh05lZQxsM0nSyBkS+IIgI2ItRkVeNeLknwE5B0B1DzwR2s
Exc1acOWiaaj0JwOA3N82zsHt6iMrSiw7FMrT2oQsPpC9Y32TK8SSbAsO0S1bgrg
Q1p3rMoN7VSgeuQzFx9TtMEc4nMvy5s+m3SEpDdr0kC8eBUsYTSL+W9YPYTnVooZ
/eebes7bnYge9LkfUShTBvTXq8fIzO+QDfmwdtX+ZPnZ4ya3BvkuJ894qFM1sw+0
Xa/IDibfHW2EYmB++azr04sYDEA6uaBa0ry/oz6ufjtIW5A+h92Q84JeW2df7qDe
MRkMCJZFJ8hHX9keErOn+gZ5S8ByYR6WZstZCXml23+fN8GBJj9VSgHYq3HyBQQ5
hnyuBgBZKLvhUqNkOD5D+MbCZaHvru3DZSJzo/a7Dy6ShKgM1EKdPqzy+9jUI2ah
fIqcTsKeqL7LFKG0Db6JpgPfIHhoYm9LTiw5ExAI6FKFBlOqlYKTRTb912STcPAS
uyc16hao9JLcBohXqDLegC3fsLgiSHiEicnmmLkaaOXDb/AfJqjA28ESQsg3lvX6
DIu1z8vBqv0zTiZnNePjma2kQlJuhL5qbeR40mSxeOLkaZ5dkBsLBJBuShR5CW/p
/9wmebUiBXRgDUq5to9fhHeoC47eFjfUPW1KXuXq8YEawXGgibA+5YM4BQ2vfhsV
Cb+61sixWTykOWMnyUEhVR0v4LoD/5I3czo4ERxYpxHtXquXiFvegc2UIQuvy6oq
gVrnqGrPgIU+2k8vnCWhSntW+rYXrBNgrCXgklNYkRJ83xXchQ5ra4Fuui3LtClO
1QEU/RC5XcivYVyiKALVRJ6fx5K7lE4Cql18QdrCFifTmKh+AFSlovOVFxvOm0Xt
O2jOhT1YWeqZZtaeDdDVQmHqg8V43rK6qtWlWhzMsWzdvQyQmwRirC068QjyJ1oH
bFFyZ5iEOXWAuaYUOKrQHcgtVHqDnTxfTIjoSKeK0xuAiwPXMX+VFqeoNoWgE4u9
S4YAsNuhHD/eThnvWodTl36Ve+TwjI+QmSTW8jDvJgArZjWeBMHrN0XUfY++k+Lp
FTgCQmNvjcasjtD8QJqzA3p32gLqpjc8z+ljSb320YwYH0wnty7RGKsvDf4fpb8v
LLinZ7wr8tL4xhu17y0WsVy7r0d4A5fNlTBXSJZaefoHs6Sdp0zEYr0CTC44gCJP
rypWyIlD/18tG57i7urxI3v+MoE4CQaQbzTjHST6ttbN9Ijx/eSYEc+wvEwh/7cE
e3lsj3RqgrSBMFzDMLq/8a0n7B/373HcGWYUbwEG2AWSC4dgyajc1Zu3vThveKlf
Eo+OUpYtB3ValFCLnenSn6VDov7yiebAgVKsjZKEmDeI+PAewPYE2WsUjAHV6YP3
qMmLJUSXoO80UNdlSNRb4M44dnwUMyGNBg+7homErd97rAe8IdPnhIwLXEAxiUTE
uBDsXFvdHkzvlS0m+vThthkjiOH1D1qIz04KhYGG0KwJtTfRPPgWdfFGCOYTcGs/
CO4grptXvs1Ngzo8UYVG5bWQGHCNlWEtJTZb0tituSMWun1kAv3hYEq3313ICxh0
fiJqIIICdgpdNRITzJ9VphnncpbcwGmzCrUKPGDzJnntI276L9VWqlGDsr93e8pj
8cJdlpSN/QhN76rXMaRrmxJBZNvv3VaAZSSsM/8p9KTVsPnokdldMBshzju+1z7c
xEK670L7CZDFXUfjFEwoVCE7289JdzOOPXxMyBkiO9n2UW8ymwnkTAPIU1QWxyiR
L0naVNd7J6pREYzv1d8tu/dxywd/Ft4OyI4J3RKHJXLpLy38EAfYmj+uDHYb88oL
UUZj2yNs9T9enfUxUlXfO4R2NJWkktz9VsKvgLqXIt9SsC+rnXaBD+8qnIEEzshJ
GPpDMnQnerYJ8ILqCS95g4goDjLWhF4Ssj5szbdYd1T4NCBDpTMDbVY9friVqE37
NTpwZE+j3zni6S6k8GbVZ8+fL4Z5ivcbxFNeddvg1+dhUf2bZZ3v0Imt4Mple5fh
dL9iPXRxQPYTi2NPQxbivjhMs7XngBMnH3AYDUYQ1EYmbnDWPOMxhiYtc4jHLSgl
9DB8ae/M+N7JjzPgGlPy9CsHAB4DMNnBJUm+263HhhbWFYeFkehY3xzDb129djly
67Sd/fXaB+2PE/CgGZJ5kWfMYQLcvdqH6xNgAGDAoyQdqSKhMinyZ5Lv+8oRjq6F
CQ4+sRsPjZlQwkJNnv36eoN5B9p9DhbI28xv6L6JLNGxj4uSiKdb/jOHyLTMlJOK
1f3WWyLGEb9kWLIyBf+8RbeZpTlhisJOPtExg6rB5Fc8TGRyb7tI05HmuTrC8UD6
UUk1o6G87ehna/0HAwyqU0x2No5T91YI7mBC8JgtagbVbleZH7ev0Qf2yLB1VMoy
5DL7S67zQpBusIZwrMbnzb1oRa5kA7p8E6yR5mVWstP3XRlVRAIADS9GHn6Rfz1k
kywaCmF+RsNdkvVtV8ea/r1QIT9q7YEe1F0AcaSxByL02Mkj+QNJZX1zuMusrjWG
pcWG9VkmCk87huHw2sADZAPsM/kypFG0bHyM8G7ygmkndKjU+CAOaN37a62Q8oY6
SZ8ozFR8ioaE6z1TvERZ9J8LTAasgvaPUusQT+ebyUWcD/IRzvtg1fAgCpZwPru3
TfetOu3ZtZ6dK8nbhI5WhPS0k2tT3aafIPWdcSAQypmJjmQK1ig0gsdBQWy70DFE
gx2ujAczc0+Ub3Z+BsySg7n4mzp/hzW6BWRyPyfsVbRSa2DLMJkngjIWE7elyTPN
36BOhSmqTV4YxZ+WhOkn7y/5HxCo7VcbH4IKaaA15GXVGJ3XSL7wHZ/3iRWmLU/T
GKFVn3cYaKIQIhdAn5QTTcXRu7oS4A5RQBMDDv0WidB24b+WSpMjO/i3Ey8jIr7u
eKcKyFPQgLO9krsjXC/e9fTwA8HKNGnsCO02nYkB12pyJqdHAkH0WCy+VEcpz4ok
MfJUanYIhvlZsonTcUwiGghrTxX44kMO+FvaH8cFWkvNC6q/hf7kNjLof5R4a9ns
Pz+kSIp2cdeXz3136i6kowlSUGXEFCwzPaLajiC4QB5zcxiu3qmCTzR1dJKqD4vU
1GcI6s8fg/S0csso4HsOODLYnPtUXb6S8qHmzuJzBBC+UqVMeia4LL8DfbJ0gdG0
MdFSKW/CzUOhJNikcDU/KQcNCEnCzcPZx2j138r3MYmAgSI8BE911ReIwEuQI88J
+zvMghvzcXAfM/eAF+Fhwd1Z71NrhssTIXD1S/4R+iCg3x9ydMa/s91XZDMMLpsx
3c7KCYEaUcNA3tQMgmsU5yNGv2n8njCZfzZF4ja7oejQhW3DDAJbtmULJVD2UpGF
iCIahkyWkejdV8/sk5O3Xkn66lCrj66zTWSGOb8DGwSG3nkW/fsmN0HM4jF6PpFB
pJxKc7Vv4E89BfWvcQcdZo558CesmBCo60aIqOqxgnamwvrCIub8fRUVEZLJlsSl
M1VjNOFjAGCNDGAMlryxY2NGB89zovA2XIseDZo9P4hIHnoQ+sM6kViyXcSdZxRD
hLj/jyp0CTVgjaGPdxYeXBcqt46tgr2Oy2oHJ34fsiTwvZgCvttYNdid2+FIBnWV
YaolWYHIbgtsXiDJWMNjzRmYwsaHfald0lOit4mlkALeNv7pdcXSR7bYLmHS/oyU
9r9SEeTjyqfgRsbVV+xwJUOkUU5pVnvu7A0hSKHEW060cvvSMyVDJF4ML9Uwta7c
ly1Inc+OAVqoIt/I0F3ryWoheAonFcmFz52Xwh15usqFImozq5tRZN3YckW+bKUp
qlkFa+tZ0j2UomJZHl121MXZxNWcPFq1E+OzR7cxwa5D0MxvtAZnMml86ASqf1H8
jRDox9DwYA5JAJIt8UAPlew7kajI/I0Nl6Md/UQEsZeft8X5TTWrXW3Onau1O6T9
nWw0MsmcyVIG6yzl/v+d0lHxiZctAB8SIz9biae0EzztcudU4b4sESk7YWRXLora
kDbF+NiAb+iLuTb4I6tO37E2r5lxtxcl/PWGv0YPqMOcZ7xeN9JbT/2fZmjaWRdA
uxTrwbsQPJ8v7mVWAjExiBwXh+dVh8V75H4d6ItA2jK4eVBP1cwOKa8uxYpftG3X
UY1pXWzwK5GduSPrqAB5k3SzDMO+qc/+a+K8JY5VyiTT5cnXHNubZuD7rHurhN05
CvIe3ZdMQOWNIdY6AFCiYzVH5quoVl9mE88oHkNsOFN2uzl7aJem/FWW4eyBdiCc
tipanz57nmOusHuJqr7BPIuPMQFIMZxxXWRjcBgKP2CI4DZqhMgiPIa2gL8czCn6
7WSMZybmfgmE19Waflzu+l5w7n+v6T22gz42fDQ+UTvrZv6Vwvl/w9u8OfFviZMM
e3KqeJWHrqZsEMIDjyyUvy/1ccsbaCUJ8Sz/Syl/ZYOTxAE285CIBFI4VEPth5gb
syiX+tthvpNsx4zLRnbXUtbaiaPVLx3/t3880IMqtoaDwOeCNDG73lTsJC7Sixlm
gY6FqmoE8yIH7usmEHQl3cyhiE0QKbHgmb/CkM1fIp0ZbfkQ3qTZN7se/YznUPh5
hyEKqsUu1/AeGGtFxC5DXHvS+5OlLB+Dqna2LhINBctOwI5pr1kf2IXWw8nOZpxh
w0hsMUkQpNnTlVKgWOTT3b3eSm5OA6AEipYEdWFKCnjRWZlQ6dNFCgtPMv66Nh/4
1KuxkiPoV5cisWN5my3mgiu/N4Qp/4B65w6A7yqqufonlcEbLpc0iwqXvI4jYUwf
TYpGHepBkFPtz0sY8Px/geSVQM9P+PpO7OS/xTnSf/ME+jyh4qN4TqPyE4Yhjnkk
2Ky7IwMP5SYvks3lK4Gr98g8cAQ1mA9WP6V27uRlTsG/IkWK6OmkOYDTdVYivvGr
dTPYooZtvC8mwgCNYWxRUeW4XEGass5WG8r2xJKQAuJ+gr+F6LkwYx/NTUVXeZD+
mLdbjmFWMjI28dDSQpNIG092PaWChnddvGy16U1xKOLaAtIMpCxCt9ft70cVBLN+
nHbAxVwLMyze+YTIcmWaSvzV4mOwEpG1ESLtvx9oGINXWZBWW+wUTNfc2odptktM
EPCS78srNlXQ0QPIK9m/ziZLK6Ubw/sYCDmdbStbTSkmHE04wQFXu9nDSIuiHIGu
5cvueEa58IMDcyZxHJS9TaRxUFrlkAc51hCZBG/T834CtOcHJ6JZJvhVux6XpmeY
uWi131BF2mXAVL7K9ytDi3GzCJ2FwgwZ9RzlJqGRTd8c3u5xWvrFgs3WFPVbHrMo
OXYU2VUB5S5/30E2XurLSsJEo1UH+zumaX3JxFIuAaIBawQkCnp+qW7h85J5UWq2
L6U9GlV8YSnnGFlUYv1Z+OcMZTfrthDDwwJY6MadRn4BgTLymnDC6JyKm8lWv/rE
gSfSZBzYKbnmssLMRiKlncHgy3wxbJEF3Uoo+lZcycAuEdoU47s4E15zuzuH3kla
Tuc153UANyi3J9BzXz4oZP/bxcF+1oyZ42Xkti58SgXiHpbh1BN9StxBITv6LLB5
m5GFJhU/PBEi6S1NjXAd6AuCptBfG7kXEkZpfyE4pakQUvYWj4lDllEUQrrQspk4
V3W9kIDUBu6st51OeI79B87tvFcyRFfiiVH464NDdmdXzmmmbF3C4R+OYnkRyzZR
zSu/b943I/ICPdcnMrkwNvxfnJJLZ+96X7bl85hZlSHIqRytvJFYc3FsDoxjX5gc
6W8n+NiRC0JIdiMDRWoIP2Wovrko4T70bHUlkPgLQFjXx3sLuyL1H4RPVY3CH7p6
oBRvkwMZjbLGMpmXDtHzYvgo/Y9bXJARPsiChu+07bOz7BfkiEZ5NOeggeVrk8Ql
paW7HNgad4DQF7CVskX9F6ji8r/NC1QPo3JrmZrXLbVvJIvvnDS4FUEx5WN1UE+w
S4QEzKNwS5Dll8aPoTR8/B91niZdz3pJqTa7PZMwGmNG2rVTi0HZvUhKkF1LPw3R
iaTyCCqx2gMQWmB++97k+DykOgFxJKBZsKLHqQy+UcSwrvvH32AEL476mz0nag3q
+F8HUWJMwDlejt+5hy7hsZX7nnR4UzNqwWNzouaPV1CWw5LW+gKmS2tLdFW/m37c
o0jMLT6RCM/2T8Xucc9oVIf3VKLguZZ4d47fI9vYzJAfq8ngWxOkA7ntKI0dXcVD
qykHojPwvi0B/AWy3pHn8SI61smFGusBrwId4RrwushrZ1fQF3VYoXCBRLZ0TZpZ
qZ9lawSDuvQTkdgmPLSNnxiLtzvJTTFgv/tfhkXLbZchhYHzuG5/X7eTTmgNLE/b
LLtTo67shtG/GNNOQD6vzjg4lNKD9fO70GBcX4dMBhKD/XeuOOLLvsAeezo4SvJS
OlT3w4ISfVHWzgXbxSlYSVXknVNYnh//lXwrWOg9IVa/gYkWjtX1t9T1BZJtzkwm
brGsbfr6N81naOK8XBvPQPGsWid1ojgbNAIUM+nzdU0pvr5b7VPRXAwk+k3Xd0/7
EC6tMWNRvbZQOGCApuVfSfxxTRTUn20vRRChz9MiAU7MkH5suLwasH/8jvHPI3cO
N+a+EaopL3agRzyLfDCrIRK+2qG7X4V+Fmacq9vXChm4ZaFGDMr39JXJQ+iqdxU7
egBhcgzigwFhKctwYrOtgtAq+MBKv1riGT5sHMNAepcosazfJk0o005qK2yLnaid
Oz8ZufgUxmrBgJVy4h2uevdhB9GZUrbS3b/WFqjB5/mVYyIf+xfYn/GlQFjdZSvD
1M9d2NVsoa5usqHLd4W+Iz6dFBWlOG9t2R1T+1g+xl9dzUhgFElxcYCdFBEP8ve6
6vCQKyP5Vvt4PoPe0infkpfFD4Kt4ZGsFYKIa19y0nauprpGgKNh3jWnz1orML9C
kZ8hLaZm21BRfApysRl79EB86goTHkO93faWQ4MMLFf+3Y3ysQQwEOtB2PAo4kHk
6rcSOYntK8TM7iidzHg4FgKtuqXuI+hJa4hmFIQ6UOJFRLDnA5Cb3lhywr8B8ueO
V7ExO0Ecv+tI+Jz1mM2jlyU1/rrJFdVTT7YYlRwFHGYdmnZStykBzNt3Z+QwW9Xy
2+wuba5Iu6zGvLjF22QSKhSx/xRlNmVMG3X50HCt+OnFgzr3KEWtZusIY2mNGn5b
Sm4Gpfo+qtNfU+r3pyX+tU/zjUYh0/BvF6Wd61NHm1YCnmzoAyN/iIj4DT72R4BV
r6CyG+RdT54uGPQnq2+XqzCpH+zlcLmbwQR783gxh25oHgRebC+xjzXfnSFDOLmn
6VQCJGOxa47tIqCGrKj/B3aJQtTEFn2afExNEcWqNe0dg7kc7lOvqAmJQO1xuUeR
fVooWuuYPG6zeqXSPOgvFa8JDE1Cyg/HJ7yEVrB9kSdSYo1xz8TNe6skkxmDG+My
+IRYngWcrIOfOr9tLdtaHec6b0ENNbJ9fjiEjKC0lAS/tDckIWyRh/Ic10hBFeBo
xZJBw0QMVhmYnNmOheZfePf4E0hHYnFK+pDhddItnZKkH1ot9qYC1hGSwh6PYD3+
2uk/BYO3bMmeWU3YxYXuk/kWJjuM/kWyj8FimuYIAXQrH7oKO9FQTpqZUQf+MckZ
HZWIHTX9gmvTZSQfTXPwXUAtGQIMrJ3JLzJFF6Q6k0SngYn3H0cehb3+8hjrS8sT
PowwwNe3u9xWexkNcyCS9LqEqlzxZ07dzugvEzNyHKvG80I+nKBTucPs2ly7xNd0
KJczXnk7bQoE1pwo5DgyPy/33WYDHV1eV+CuOWk60uif6AxTNDVbVcleS7Vm97AQ
vN17/XGydXWso6kr9N5bD2Y5c27ChKH42C3jMsYwXP1Z1MQW9ibqopozPyaC1itg
0VG9uC7KGqFiS7EbwgggnCFsr8JTXr4WDgIL094CtMY0CO6GrAOQET3PutoH4+3J
tCF5SZrzCihjKeIkZ0RijQYFmLyzEgfdGyN85yY9H1YvqvoW4P6p9feFMjMSigyL
u+FfQZyLWQfy2KP2fYOxSzLkh3J6IHct3NbcjnS1Y3fyeA9CNX7LRFzsQeEySZKz
pvDob1/XD4TXZPEA9WPRH/DFMg83w9G5lRwPRm41TGiaEdbU756bjN1BwL7+CYLK
En9T5nZrcMe7mAtGM7M3Q+BAYMuU19zoE6uKm7TyQDjhT5x9mKblw8eVYAdkrcwO
3XpFa12/MV5ggs3jGZiky8OBcRbVdC77kXmf8mo2fbOJ9p61FyhG/kM1FziPubpP
uUs2NAfelaIbhqGxtexKP8Ggiv5mAT/jPzIazXsGCW+9Ll7xf/2srGqDmotN5JtD
pDvQ8gG7SxajSpej9umCpViHyNxCyYJEBWOzhCQvrx1WdXimsk4DGWKc/bDjava2
69ncfEaErMD0WpreLECwZDIuPS/LhkyG1lxQnxwgi5YV0B8wY35vSpDQelrULn8h
z5M1Ovi7Fc8QdDbLdkUtbTLVT33gpgYrTyIQPNXHiA8gKj30EC7z3Hk5teTa7z9R
dgxeP7YATpqnROqpa1oNkt8q+rEocTFxb50cM6Gi4kt30PHU1XFCe8eC5+hf6oWN
E9WWKdIwO9kB2XVYvQw2fS5jCeyK/+i11gND8snfChr1J27ZOYGWxCR5pR0efeSH
AUU3SyQYyR0Q5Z74oZxn9/NQsyjj72W5bScpZCaxnyX+Cl0tFGpPI6C/Bdm/r726
HEmZANcu0bf/Di9hXjeTpeLlRL9CQHRp8gbnjxY+ftw6/180HTjKb9h+1fVzKa8r
xxXdQ3UUJve/f7LpEkShfQrnkrVXF7F4Xfluobdq1XP86upo9KUyRVkjIbBXiImi
SDwqfjWRqTCG//TD5cVrKNucMVehspxVIhj0aybLcAOyeQq6Fn1F0nJNXwyBY2bC
qcYnkxbuxCHFM7oEO0qkrZpDOdLjhItSj8tbddUly1NiCXQmaSG6B80qBVV7wffA
qPho/d4bsNSKdG52l6OOUVNohV2sI6fkiV3VQJ2H9ajP3OGawdrJNC4rzIRrWI+Q
clymMbnJ7YtT5X51KB262U8mYOR3JsbJns6mFSbus0rsK7su7+lD9I3PnizIrFUq
yLIvITc3ITJCrkTqSr1n6AN8YccpKSgqRV5Jj7hErWQ6PgzpQvTmTGaKnZYbIs+4
8XODL3tviG3j+iIKtGVP/08rzLWxTlHC/XmJCYOL70TV2CZlHcJk9DFXAZXBoBUp
338GDfn9qugbovGUxwHoE2xeyCZbF+rE6t8CGlMyMEjMQJ0gpDluOJ5U22qG5bpW
7oA+Hk8YYl2cAa9L54cAtJc4/RE55LWKesiD71J3JWpxdBBnRfj05z9UDrkAdmtx
8AYMIyvPypqyi5f/LQV84qZC77jQP3XiSNfK+EB3myHz8Vn3QJVMBq1Vk74MK0jE
rSGzazqkI2eTxuc76BN7gSYCB4eOpLRnsoWIrUoUZdku1SAsZpelup84Mrv1PuG2
uBPYuzVE8qyie9Q3j5gNifSRYyouJFnfMI0FCeVcOXTmb1PwHbuA+CPJDG/bvxnO
pxtYweXUXTfYqomC0Txf1Jw40LUFIExFlbbRU92SWyT0RKp3uHE8mZmZaGR+Pglo
d0XmjxUuUwDWPaHdFRR+mz/WmK3WMc5UCGFNNR47R1FIzk+yKJkahu0lIWCS78u8
FdFUY0r/e5pfqeOb3jXOWybY2rvN1q2CFUtxg0QC4Hh2MZsXHOsxfPclR/ozK3jO
QGh+OpZuCm7UrGLN6YOYScT4RXCnA6dQSTCJ35+mBSgbM70PnmuXuqjZaKJbzM2J
TdAoKQLfpqBj984TNntDTOeDU7RO+flLSaBCLMe4vTzs+pAHE3kn6Knr3q5KgH1h
jLELAg+Uzqmn9Y8OQ9vzq/x30v3wbXmlynQwkf0WK+GnntgtdpWbIC8X0pBS100D
9nauqrWc3Wz5x62pwsvlx2Mn42YbXEAwcmhd8NUKEPBiStDzxQfqt9mfH9CUZwcO
1aQdwcKYvVGLTj87egsSPr1qrHGOCcjqFJWYhYhiqEavUC42qxBnMnh4dGizqnXg
tSgL5kKqS8rxhR4dPkr8HAWGRGErD5gL4IU/cW4CA2+qNKtUHbJziZZe7rGMCjHQ
vCFZbeTtNE/29CfKE9hLVL89ZZlpJlv06vFhc6ZhRUymTb+k8MSGPtBUh26Qvp3d
g8wfbW5kkPyoM90ahU7MSka5hwHWDoxoV+ClqfXV8GZ6UGyVuWzWb33jqFWcGq3E
PWHkECRpyVeukuBK9tA+Pf0LRfuzvul/3BDTZTE/JI9O0oRDQAjcpIWi7P7BxBMv
PDwGHQNZFy6TtagLJptt0ghFQ7OgTHRGl4VRH1Siqa08D2Bj2qP60t5s6TtAyfgX
WuSs0Z9og6uW9X2HkgVuAqXAnT1UR9fuZA4/I5bg0EGxmrqbJES8fFcNxhWT4xqk
hboegb5SEZo2kSj+5SArL9JuIYWwlzHO1JkxrQFddQwreWPsyl8S4I5NYF4cBxxv
5zcl1TLaYb9wHCjBCQ9VygwiSehfLVQJc2c5i1qtN17+tsVHJs3h3z/RHZpc5Wkh
l2ilK1mq4OapCVC6vlTF4YEb4Ne3uR/Kz3K32VqIz57HhYUZgtere9VCDemWohmM
r2ts/qXnWo/u1KV7GgY3/zvBqEEGcr+QsPd7U272Heil6b+jtji7zOM/uEyy/kby
QIoafh60MVuyfU2elQA/KCb1LamNdG8/1voTWlD03MLfEKDDGmsivNN5sCnNzWJS
I86phtforzhgRlmeHhhAGE2NU+SDCrlnyT5OHpHrAD0sfGKaUz0VpRCWXm8K4eVa
hS/dVO9RzvkVTltxTDy/iGMCP31zQ+5lQIHwbRAfdjv6AL6J7fc8rhAJcQJiPhwl
IxgsY7AAAP9cpref3Hl1HGIuFvM/XApP3PQBU05zVbibyuE6QPOs3YHfIHeHEpXh
d4bLZbtWywkarwdPrSA+tYIwo7Jg/uqMC9TL1d04H7aSlWf9v5nnX7qbvvM9gWZa
hpyYELp41ddyqquZzvrOb/yV7AfojeJOu9UV5hsTLX1/12i+Qe4qn39sMcsixVeB
w52sTzl+QB2a6GSu0e5hCY/uIxUR/ygy7zJu1s6QWJtrlZxRoSlWqMbm/F290vlT
NDZNErge4DkOv/dzEvkEwFrDm6XceOTuT+vcAtvKM+qEBriuh64Egs7QvEJohpaU
C9SjJV9BedS8vHmtBLl1kxdgzvRmC0UXq2bQf+apHddyosXX8JoxuaI+mLLEKv0x
u8uJoqGsSclVlNrWLYqUrtOMXj7ipxYLrCG8gi1NYInkuCkiZ5CW6zxcx1UFWWYC
5miPXfJMnlWlYo7orqVFqXXMXpcfblmRxTf/PI+qVd5mVql4SrnLxiSkz8zDo9+X
rVXWODxluZjyHj+npnMTxAyxrzLehWZEm8Msoj7UedqHVd2K2V4g1muNUJU5Jbs1
n5rJ7gFowYzSaZHV0a76bn9rtVAMmIjgJ6soHpmXJJCWTIpgR2CdeoVztI/brS91
YaOy9TNYLFD82FzDGL5xqN3bPc40Pbpn448bnUUSSoEeVwEsN7gEciBZfSxRFXqs
Cyl67M6tKpnvmddwQVmrwhcEs7wDevcyqB2/+3cBv6KESl2MsHnn2aWuH2I9W50k
Z0WtcSmk3ulM0mZdEfPMs9BqnZKNSDCf8+USsnT0pFSKEpbyEAsZubvAtKFwcFA5
JVPCTjXORoG9LC3f9PO0cLM/SZYqgomrB+w1FTKowmSbAH6150unbwydN+AsuqJw
si15EzHJ0m5fx4bS5HaRzB+XijoX/jmsci/GUFSfygZIftB/EitXMxh+LibciXtH
U1mQ7w8w9pCbHQxwqLgcr48x4FgjGG5uwfWBEehKjMhAgenwITVpm8d0DMs/pZtt
dbtJbJqMpp7h7ipXu/as+Dlmj+1qh9aNIrwzb3b8mhFpfhRWXPeCd+yPdDXrRHJa
zG1rUinr0WZWXAO4zlt2WnV21RMo8eVh/xHVVg8PKbJ9fB1uAawr+1ohFFhfbW2G
OAor1GZxXKtlwxYoY4xxFrZVCMaHfAzSNm0XMOUecuBnHDAnHoO7cHz/5KBGaIuY
TysSAqrMTZQEk1qn+Zr22pldlrCt8RMYLHamncjFOHkPLleE47G98WNnq0+m2Akk
8fPn0UxGZ90bq+XJIo/uVcZUGQu3OdPclCRviFdQn05izpCfL+vc9wg2ofkCNbrP
7PwXCY4xFoS2NP+iPKoUH2CtwPU06Gd590FGRrUWVbfvLvukvbpcEpkywozJT8Gz
6JmEkWK25unCxI10XtZQ2jYZ5v1rvOxu6AJhsVxViHwCW6zD3PHFn23ydRQm6DtA
gQ56iJRcNEnR9dN+NcfEYesCNWxsW3qnsOnd74H7O4C+49YDMgKvSzv6Qz5BiXCR
VFNwcLdsGuikktmiCAuFd1c2gcMq499LYzvmOt7WO8uFGKJvF4A/Q+aJ7URcCdKS
sYSGYOsquWskFDOCCEEEgf2gjLm7yi0f6B3LuBGH82zpSvrkOTswQRSTIhzRLcYT
4nPwwOwQMNTtrDfKJ8ypstU3hqidq1/0WgcLkOe79rwpRq+uS8zWAbSi/7z1u009
X+ybBw7NruFzWB9qPL/AV0e/XP51VPK022WW0oRE/S+9etdXUAOcl7Mx1+hzEHsN
ZrBeoWCiM70/89YC8HBC7iaGj1A/VYbgBuvcSnTcfDiC2/uitBBwFrQWR3qWRNq/
I8xBiEWIRw2wFdqciXbdiPzcrtCpAf12SG8Rsx8YzhF92uZO860PF8qVKKdezjGg
rm9HyLfeG7VuP8nyrFCzTg9RJHH+JHGcUVSmH5IEvfY/LdAnU1DD3O2bEmaUxsbk
kxumKfAbZ0CGnv1TgoAJcS9bk+EDpGfFAjPpSA9OU2Qd6pzUGyN1hy/FDi1K03kG
RFUySjRkga6hmArrXc7ElPPjDXzPJ2aBi7t/JAJbVIt4IF9REUNmyKWMT1XfO4wZ
RBXlqmpbn4QohGTAAxU0WSii3qgfKVI3HcCQ604QSjrzF1Bnfkt4OBX1f3xmksu6
EMP2nAR/tnJiakNnJ6X+XtU8ujAnOFnGu4CpU6KcHywcZfC55NwTDX/0TDCzEHTs
wBwHNzTp+ViyOLO7e8pZvlieI59h1b+T28MGM0NOs4LtS9bY4j6yxurQZQ+QpN8f
jk+Cx71tA6zpE2v762IixRTeUaGo53Ea+BYfZFYiA6zC7KkVbjLfev6dw8kAAaP9
IlxdpAj94XYz36QC2ebazPqGUoBjr4i06OqHTaiNHCxqYVdno8fZz84IdjjB3j7/
+75cqgfasq5U5yXCV8ohmrWM+VnHFMJTPRLCamzTYoh6rzUoG3ylqtFrMjNWFJ4N
SqkHEg52nWNRL7JM/IgGiriFZ128tpgZzBun7MVeNdzzP+E4ImfeF7j+rwUPlr5Q
yRcauCdJg1h6FK42Tn6lG8SU6usK1mTOtztZ2szglspc0xlvT33KgLswHf8WhxMh
wrXgp2+ePnxkycLnofFm5x1vqGtTm5RYHflDYMM/HDmcxWfXXdAWC9IlpyqRvoeM
8R2WNv0CO0ndxN/ilGY6CrJbysItKQcnfennIbri4mydd0Ohq8Jpw1/p9qiDLHBL
4Sur70QPZb0gSn8fFg04YCIZ5LKFa8isZlBZu/8w5bvrWxOUf2IWEKGlvd0SYq+V
7Nj2+97O7Chq06CFIrxks1d3BEhfcfp2497WrhlxOGtaOLjQ2Zan9/8xVRa9CGAa
dt9DpvMiURM2JS5BgMBYd+IBvsu8v/+6kkHKQgVjBrg/eiaRs2YoF5RAXUoSDo/Q
/QvZC+wOv15NW7nvWo0EHrCNCdf6vRT1WB/MU+16Qd5VwV6WLjSCT3Ki5C/iTBPj
MYr+FFVwUhnpxVI4ToSWatgn4ZaxlTNJuIK9+qBsVxDUIPJcUJWBxtzOuB61Q+0s
StMC3JTetjvx5YsZ4MyKYRZ/lH2SZ+gXbku5/CnXAso1DONEQS8fwa+HaUBaTGZV
YAVeoXIUan31epC97z66ibBYAkee86Ph6oETBAXLjfNm6p9T6wtIGc49hawdSIdn
lrPCm9EVp1ynobiU6x3LbhHOFAFJ3tmLETDOcFSty5gf009cwOcc2c/qdw7QkJbI
fCpvFX+HtOSApC5hVoVxdmiHCNjsrkhbcTTHFcDfPp5fYXXRTVFQJ72l+s7h0ebT
Vcdehgk/6yjgvbw4G1xG1BNB5fS5+VulBj7WbOKdbrc3/5+y74AB4QpK4Af9dnhU
tDblK/A8XqYfSAiP7VxyA+VTh/GZKYZ3eSi4CXQMVxkAW9di0w5MO8Ha9eY0rS16
rv70kVD8hxJBZztAiKvzpMOp8b11iSciGkAjBgUoWv0stZ3Y3KvfIKp+tt8nDQKi
EXy8mgxubjDyYPGn9vwIrAgfmDmYj8pcebv/GkeMUuBBosIidX8WQbvrj8TEnFhg
qHlNNbo26Jz7J0Ea9bZJVvxNI0ffjdFU/KPyZz+irqoWl9+MlKx7NXLieNK0HEbX
c4ZSabC02Bj+Z09KYzdjYUmqcLSdMwrRsaZAIMk/gdWmXP7qD4D38Dh7+xdDR1/t
PmHKHxT902jwwkBw6K0OphBHc8nI2iOzzFG/vOdQTevHTvbjc9EmYbdz+CAZrmJn
V+mlOGEWyb1jIck6uK6bA+hE88O8JaYMJv7G1bflcgtSHXSBf0vYAGdv24mCVMXA
rTMvlXyF9l6XIEqZWSwDQ25GaFl3W29/cxx4KcPSrbOdgkpg4ruJohLp5URuhkeA
05QIr3XTQbJpT5gGRMoeGcZu4/OkpXAy+OnIHiOTzmnExntbs3ov/AZCGtHivl49
czNaOG/spWIehCIpphyol1suq33J+iTLicfDiF/dCx56l9PM2Fk0LCSkqCj98RjS
neukOoDoO5QVbfoHpDMe4oDYafXxPHBD/vM7WekJrtZiROuGw1Tv+DKVKep9iWBb
DmpqWFPmK0qpqDVzDtBu5OoFXtI1L/YiN1WUElBDHzdIYvQvSQin+toOsuxnElC9
PDNg29GuoxmDuHGvItpdqrcefpObiHz61g6A4GqIh6ywxRrfoCufnJeY3C6z6EVY
iCnj66J+UcML8coQJDCabaXrFWQoEYrl3r5NcOPfs3VI0HzxUkM4tGQHzel5rRPk
3ZXfxZNuvKJk3MsTiPGE71ZpUGS4mHZyQAnHmGaOCPfpy17shYSxJ3wXXclLW4Ne
BJ2IyKXiOBKDOTyj/WE1oNr6j1xCTrBCg1EaMTGU/177HgFeJKKjNQXTNlbDed4f
c9i5g9EcOxPuvBEn05FkLPeX6787AFT4JI8u3ceic1nqxaeSWxs3nntFid0At5kJ
IcydF1ayTMrl3/XBlFBNLT1hgQeTBns4msFRraI3OmNMLgPRn6HInC5AiIoCqGjB
VhOgq6kFK2kUkKcMLnnU1repZG+s22rBGUHXyiGYBLXcyAX4LGxNfCGwWP7ACLEv
VAPnzq1pg8cFOH6FvIxEkFmNjaw8ViXXATLYFCZ0gmr8aC9D3q+p9DV6umui45mI
WyKmttDwM9PQSVdJj8QRQ6RlDolT+tVjjhzC4INf2DWsNuB4ldRrx4en9DV/KFn6
6uORhBEnlQU5pN9I2bDzKVm+/q5FAo24UHdRJVeDTfTxk6IyQssPM6BYpaspkbru
CB6xiJUzfAwzHD7IfAOAxtNNV2nc4wp0He0+lNETZG6ZJ3Ua9YnoADF6+PJ8rFaa
5UWwp+zzbLqM6ebcr/ehC3vy4TCYxVReIFvPi2v0a8QXo6PwgQ2MbEgxZ0eUECJ1
nFSP30tJfhDVZHf4g0/tpP803G1fLpoe3rAm9NLWmrMa5jDQU5YaWoEFonDIX7UV
60OcKPwnZVw5Z6+KFNQzvlQ3ri/vCdt3Lqjh/7I7hv+AgXmOSyUgzHwCYDxrBFPq
/P+aKyd2pfnCJ4fb2zoTmkOYxcaWnaGgPU3d2Pg3iIZzmkn039q7PjZyOCdbbpxD
r27i4xlVC3TipXxp4P2vmGSe7insK5xq0hPYUeIUjeDX+RROvyw596AQEIQBrT7G
Ip8KtQkgoilL/Hjf5gvNMwPQe8QTPlKDnXznOZRjeByzjf1rhOo5acZ9iA9GYHZR
CWJzv7sjqY62cdbfj+weKNSjQXxeUFun1uHhRqZCjbSOhAyLjF1xU1FDu+e5bGua
Y3wAAWNR5tScwPnizfgp40/gaFc+ejFLlt1kM4F5BoJxkzpu+PwAztVAg4u0Bb4i
WSXdw1KCYG4zTGCON/GqVdvH27oTs15f0ye4be51pKM00Xq8UNvkHulhO/yQDi2x
biqcNK5nrEYN9bSxyOHt6D0mql0O/LO9ihyHJA6cNGw3X6yqcQ3/YLMGXJNY7R5f
QbD8/1dT/qBT4Wyad9AL6gGVq2HOZiOQLZbr0MU+rTMzSiyVyjJYjehE2v/2hjPh
CUZoTNQ5c3hwaIRplh5bNLXPctu91OlLc7hLP0BULT/PluL0BCmD6iqLXJnFoHou
yz9XG/1tDgjE2wmByTakRv/1CvD8ZK/oZ4gnRTSMRNHqZ+v6jsiNAvBH9ac2S/4d
H75NL640KatHia6lClE5CiEmai7/TIDxGEKouF/MZXC9MUtwlMTcG0i4XYcqtHJZ
fMVBRAUfpak9ubjBHb5I4/LwxvkQCLxnDQOKGzROWHj9nhUAwSqsoLJay1utBdK+
ErESMrAlP1ZEQCgp19hqNvtN4tcpvQv7E/XAwYjqx0huTYSwo+GNdNweBk/MtrSj
0DEVaxsgBJ0c7lnze6bqVC4lAAabJU5hCT1PNyueoWUVAFGDmC8FITTGkw7OUZfr
2gNXKzrx+PVovu6xsmYcLx2XDJu57P5/SYfweAGdcTKSVX9J/2BzV8R+bPrMzUON
kOOayf62k7ak3oCFkwOr97xznPktrDwDZr7tk/IDQLbXF244fofk8O5c2h8JVrcU
YXKFOK8XPICv7Vf9vqWL7IgYXrZd6Hi/QMULtiNdfudYY4dBprWGNAUWiI0w1YUj
amRug24t2V1fFEBJuqPfBGXn7AC0bsqvrrIiiOvt2LmikNh8zidmSBn1qJd1VyPd
RGOmNw9RYQN9yj9ZvDSN28p3pD3RPvGY+Wj2UdoLGSpyUC/3ePiqGSFsLucgnYDF
haXnIQSj9jRaQ4s3BiIxITq9fVDru7d5cu7U3riaCnRjW6q8DpMAm4If5SFqMME8
dcQWL+JSXevTGaptssfsTdaL3TEK7YKWyXWVWWq8JqruKO7tqf75R2ZNFZ4YRxXZ
SO/D4NacqpagqNHeXZiTwLhAEaX/UsvsXA7NsLpkeB4TbHI2UK6CQ+A+SIT1X8F2
fxZ7rilLwPahlDbgjIOhq+mv+O664D4jIGAM9klHC0N9fAUuMXW92HBTMNJXO1zc
qt6lhasM+f4qg7KqLlp2aik1kuPfvu4CiKZP1WXaY64RXxU3zpIcV2AbIJJE1rL1
t+ohD/U8gyU4zxhBcJc+v5uwXZ0V++H75g3hqVRvi4/NuCrIFSuR5Rgqs0+k2IqM
XT3yNlmQfao/2wYkv7IWNSRrWmhJCZcLwb27vybhEadsBh1XjVV5r7UZCWM5Whmv
HNlIMN0coUk1iLJHppjQ7qMDMlKAoBsdRXf48BejUYorQhP7UXssYgoua/JfbpJ5
SJAHwh7VpRJDPuqdvpYgMUvraqKA0R8ShMhpZJ+HgbsNeJgamHaPqaamiGNzAivv
F8XEfUWQJmTemltGLiX7p1qyjh5qCJFjc2uZ+10552oj8P+cOonh/n0HZipDpVCC
XjW8nzL4nXkTJujZ3jTTgRCDQwZRqc+eKB9I9zllKuhuSKYj/j0HuN23pYDicIEz
592uF4/GA287Q2sJwseSriqLrkPyJIQufQqrTEVItkNNpq9+dbQCeJX4Y0wisUeU
Fix5WK9ntAThr7sZHfJLE6b5zz+KnkBwCg6LR5+P9K8Z9V+rJhED9fFnYXJEQmoY
f1XTadDsv+QIjBw1vyO/n7jhhF7sQwooRkJFnStMtUgGmFK4bapIjW65QH1e2x53
b1X3Np6U6PjUXlQWCB5ld1Omue68JkGh4N9HHHBdU5HJnKVnE+mXvSQxKFQhu9u7
ZSZK5JttY2e8vT4z8e2AkYjr2/OrpPpgFRzNXQb2qr0E3DX4FSWrtFAIG+RhDe1u
dFHz+QLMuhIS8HEhXDrI+cyRcjRwifdI5/Sla1VUtBf7v7FFQ9wALdd9EwYY3MId
vbPYMU2Mbh2H3vaPPA0Xez6Vqsh25AyXvHseEwlUie60+s3trfeoBPjIumjVRnDt
fzK/X250WM4DOMNLcKa0W6bOxc58lS+wkV/Pt4TeS0gkkUPkP6vhCCygrkn/LsHG
kSHHnZEO94EFL7ZDIiclwhzBnj8W93njkm1GXsuf8kVbMB6/C8zYuzT8qYfvy6pZ
xbGQH1PeLiDw4Rad/Rx8BCrezLNT0AEjxWBVoZopBsAWCP9RAMlQb4OgFi9V0nAy
h2FmbHrGFAUXeBxBGNGvDGYZ2Uohzr70ri3c8/nedlrun4l7kOx8Id6Wn68KPxXD
+zYb86cBB8OFdTtnRk0li49FBYg/VXyUsPUIzwjWqgkI9HbxiIl9L/dmGk8Hpvx2
DNMl4cIAwnusS5Tv++v1G3/54Sa4gyf7HbcQqQVeqZZHm6AUw3uU5Y4YBh1c+VqI
XmlzAqqf/V68kBQu2zFXna/fe2WmvihMxhbLULWDivK7Fx8J+1oVcj47ZXRWXu6r
32929jFMhoBLIcM8liovbPPUIT9PJb/lLgTvlOQ7ie7ZNkgjRDEeDhk46aerLwmp
kN2o3uM8zJjTC3bYqWrr+ud57hfpv/TCVWpmpe2H9UVhVeSkwEsiBzkDvqNqu8yx
9dmeWyLkavrPOjEaa8y2IdY075pf0oNC1OPr7G5jvYZHVlyCZNr21hr1ZP39O4hp
lpMTA8vJbh5vuc5+/fz68n9U74DYzg4513G0IdjSCONwVNOtW/bDUl2tO3fKLpIH
u6hKYZ9Cen6H8sOcpI+ugI4reosjbGEsd8dkTo9axIwThyn8yYufhrX4Nfo6qxw8
xyh2CtP/4n4wRpZc3HSnHnf28N3kz/0BZunLvVwimFlKS+upOr5o7vpyY5Dm0Z7/
ih/eNWTwInq+2d1o1ncdggqduA0Ert/7LvF+lgrcm3M2iUJl6aYMMoldJMuYDV7t
oprmjm/e5yRGXgnG0G62zX4P91QHHxoXXwWgRGo7gQARd6oiB8eXLTRTQLPpNyLg
9Gx44n5t+WdYbcCJE+beV/I/flfmnMik/qkulrKghVEgI0f1QMwHyXVzGF5E0pRO
Pd4XVTEs/JczHDYNDCDfRjd3QEZktzD/+3haq9bIT5EMq/ZMVB1XsL5fU7oWG8bM
m2nB2acX9Q6tUXX6rbtBkjNyERaj1ecC1fB5xtD5NynuP1wsajbfOIkQN4tOnQLM
a00otw37pI6+ZWggD6Hh+lQHzf+r4S7iFwwlLJdUQvk0RBMPqrAMNRed1MZfJ4mo
2MP87KkRGixT3zdXMCh4Zn+N/M2R0qnzlEa+AxhfLsOaDJQhlh7+dMeYlbTg5pEi
tpHBZ0rVwYjLk393/CDlKmnvYsgkysyKGu/pjg8da8T9LoI9UG/29bYMC5773ogs
kKQ4cXNjtRT7RHUvbyeRejQNVuBvoCY85fZ245dJ8FhoNu08xceRuSDHQWGO8QbH
lkDbvfwd1vvYellIbqhs/prp8Iefk1Ipiu07TIiwtODrkC4Rg3Kc0GcZreqc9qbu
LEO6J6cmlyHhc5tgn4kvyvZDoeVJNfDADfNB3hYCJcWDu137VJnsWoQv1+HtuhtQ
7aZZBGXNHB956kaK4LmgLpqLHjJJOmb2zNlDoeYQQxi7Hseeck4ncYPJ5Fmpo8qZ
VHjPPcv2IPUjzlAX35HeRtzjKcGJXXPv5S507rsLKJsQ5hsQIQWRth2SWTvuCLQb
g9xjYpKpb++7Jy7yqiDU2WZSbDKfNQhKzFbmDTy4tH3AK3XXCkkXyub9WAFNjgV6
YAd+/qqiexMi1rfkZU6xNtdVx7c5exJHpHkDmAf3wFdkiqMJhsGYL4ZTlvYjq4Hy
/fsYfRYy/++TMepmYcLXIfvbJqTg4BDQp6zJ1R67Co11YNxBs3biLPqhGsO2yFEO
yuUoaCctm9+asljXA5Votdx9muqdzfWscSh7kxYbIlmZggqB4Nrk8DE+vkUfY/k6
A4IHXtRsuCSeOfJT+ZBV7JgcjAkrNUtUjGyQfHOz8qaaqkLTwniOz1c7De4FuFuU
beRwUQDqsW86XyIKREZbXaIB/Pi+NdnoPeOyPwjS14/jLDF86Ls9ZdkHPriHFCiA
dq+Unyx+ZR4+HPdfAs4I0xKsa3ebWvq0I317KEBn5eNLS7Wgz45mdekDUKuuuZvY
cJW/dzMBYzxX0OLcDVzNdlyRzxqXlLXseaF9zQxBtKiQCKI7rv8nKDCQfl17Xv+t
Gzhai/gaXaggnQ0jpC0GbJmZjVCmBTyDVWoX+1+wFJQALlpO1L1bKJrRDt3rb3tK
5kZKf9u1cGu7XHwBmaM02RWjziIAeYVT3Oelcp2e+34CL+FpIxKz+MrSeDEikbr1
p7QYJr2fCC+1BU3w1K34Rrdkz3D3YC8qvuIjkW2h+MjRNjo21bXmn1Qc/GuYbWiv
G/HV+pCSedmFL4Irn7VmwqHHz9me2cp2PifjIi7bxean9ht7rYlmXOwSH2SzNMdR
PsQPn6dj3jncX6HfJSsSV8iebwe5vskU90Dwuqip97z35/iG44XBAEz6pz8v0hn5
E2iVR15hqWpoYfO/Z1BMjZkLlfKbZvq+jD33+iPrztPKblYeB7c96kL3ubUFstkA
JIufTpFo8gYGyXjZqU9FyK68sexMmc/7ksxLQ7xG+jW9dtw0BQDAu1+OZRCCXvB7
+QTa+ZQ3IM7LkxxIjTFt1Py8Usa4st5WOPlOABivzdsdIPJosY+daEHwZUm2ZGC1
Y7/FyH+/RdSJq2/bwcwZAz+8YTlBD/0s9QjQ5md37qoknzN9PZwldeturdetzHSM
Actlgr8Txph1hbx1p2BPabV+6WnamRdu5NL/vLfWx7/R/08k+CtZvcAXZz6CdRYn
4rNkOxTyjD46jR6bcZrakpekR3ka95Rnrdk0Lqh/+ywU3FnHmvmIN0k6axAwdhLF
jALv/byYdrulXvWT7oTRTlIHsZFdukIcchqt3TmGbp0H8GsbJHXhqadelk5rvXhl
CK5a1sDFS9+Z8yoTYcqB5mrOdbDZdV3cJvjKK12WNwOuplstkASzMtFyYqrz/7XH
ycpqehT7K+qDuUFe3SJaQ7lxCxUSSdH+pgC7dQOG9pUKguQX3gUedUuoIPuC7uD8
pABK+CRKoEOE+x9PvM/Nwpq8/gKdqWw1tzPPEwWoKdT6ptNoYzBgzXBoTJfRYavn
r14Hcr1n6Ay9VPFwO0nQRC+6k0MiNi7FuNa3ggu6IUVNAA3wavhv1KU2yHk4sPYT
zPY7l/2c5zcx8bKiqAWwk3YYh3rGR/bS/VUvlTVdWIGL8pL+cx46F+yU5iCTEGCn
ISc9m0hRQTTtakpteY6y8QeI7j7GT6PFTw6u7aLfJJfvpzumK5TztNWu+rII+tKd
eck/TqRKc4S5R5oPrPJlz7y3J5oNG6nMLuh3A8asw+T/+kMzKf66bCq3kUL5kWs4
pB8U84CDx/bAOrnKCtGE3EBInxTQx0I/+NpJNte+ZTRb2NbP9WXVRI/LauUcUQiW
Dtb6KtUG74aEhS4K7KAHyb2iKcBPuwBykUNS+OlFZUVSOKdoL8l4qsNKhdwv2V94
KyKxvH52qdyUzZvnMF43jpHIjU+RfYdRufvhC+k0VM6zCL2lcJQHngwKzuNfbr3e
2VewYkujV1hLrGeqMdpy8Uut3DXABv0txT7YyrXnRdYOVsWLs6gJS59+yMOFZyOF
BkRJ/lXCiiGXS075djuWhcndg9ThMDpcy3PMGvOtVpEM1V33jCrkoL9b/g5VAMci
2zhigD5NQZVJWl6Y8cv2vVIj6BW8xufh700yyxnaRjJdhrnwG5eVhj3hZiJB654q
P3HPqBxjgh6TJC7l+awN27cdp5iuvm7v+mYGgGa+w5o6398jV0tHIWUCF3DuVUNH
kARtjWDEcLa8Ib6ke70ajvoLjhqnkHm/zqss0UUH4i1dntSbUXo2txQX3PBgGPLw
0j6tNhpZPMFnKdRPBdxZw9UM1KHBpZFuuayLLhhOo5aFYSLRMw2n3QKnkvsN33QL
rBI+5xWVSaDJ4L1KQet9led86cv/V8oyUixBV9hcwidm27usFsrNkelQw3t8/Fhm
MRWUEQs4WY1l2s4Q5otB6VgLFNhPWw2VA3+3N+B6k762+LJsqcKzcqpJYjt4tU/r
dESy31EbQGIK5ohWI/ZPgAkccIRr60OE9LwpBAJEslC4iUUuoASZSS8xeVPI7Uye
ZWmxjDpfntUC+JKdZIzw/0maiIH1PLolFMWYfYsp4ukyrY3wKpG45JvIjfX5unzw
5xcYe8lmCEWFug3A2OmOLcgGpv/Br0YLO3JH1OsEFnwltIiryT0OmzHi0/10Dr4N
OIIvMHpn/sAw1WglJ+DCwVEFvNiwt+gGFOADZhnSvq65rM4mqI6UnjrX+c+ZLzAw
w6TmbkuUDRRuBsY4RVdVIlRBS/LZXvEezzkWjIhVwjmT/EXoaQMhNSRdr6VZBmsc
3071mDmGVGMvAhJxjUuoHunIJ3eVeynxhTBHukMqWPFayooo7GXSiJfySg1tjqox
eD0v6sVO2LXox/p6Sc+GZJxc/Kbz/Xyq/dOvjJ+V6z6Vykbup6pTITvmXv6zdQmK
2lweoJI/SUfZl3uXvTQbEqPBe4kepGQPd+76AhlD7z24HU60j9chmVO1vTAarapa
5mSfe+SabZG+5ChdFOHXeTojzwVmePrp3XcI7U4UUhz+Abx/tuSGKA5aF5bKonQt
a6bCGY8xLwunp9HxnlygLiPravFm02dKpcb7P41QQbxOWA+koYXcJZR0KAI0fPfV
Pr6lM5G6WzSBTxxofh60yq8nhwE1TnCprz/lFzAKGqssWU0L0mwOkHoiMgijCekj
qbaYbjdQEfrKCHiJ8jwz7RmFsISmUf6Nv77Je6BQ08g6eTmYe6bCY83RpxeV/2eh
oto9KTdjKTcv6NdWQwh+UwIYBPpOQ+dsoNhXM3w7wCZH97PhN+tNYrxx2psBiv/p
nQ+ma3u25MWqgxfPsSErIQG9J6PX7Wihk+PJGcX1n3rTiLaAK5ipmoP+71blygWx
cwp1+G1kNTXSm+c3PUklSKGs1mMxMaJnh5oYmq5kx5ENxKw2RA3uDGp81LRSRTuY
e8frm+f0PhEu01trJcC+y3HhaWP+E0FtUo1H/Wwp+5Lv+Cxgg6GMt5GMsxh0wiM6
Lyu0JysCYiyDuU79e1A52WEktTifkOtVSSA4SIplyz79WSD2EGxG7MBn8sgF1PJA
BD99HIImKIIWONN9mhEmaUHHvzZmsVSznJZvvAAW2OQuFi9MiYV7tZbajfX46jzO
Jtp9KVYtIZWqiZODHeLSQeFS1sMx1jR6cKedV4MyWEGmnETmnmVm3275OQ3GY2jR
VGukbTGUlxUWjOtNnTBPghW8OMC5Us89rRJXkWXEoIhgpULdkHjsk0gUx0xxd3GZ
VSp3Ax0xkDIoKdRusKkIxO0tYsVs9b8E+y3kt3tuXLo4xgSu/MftHqfGb4Kba93X
k2uE7T6HQUCQ+83kIyWx3lTcH/lJGokN2D9e8DvEKLiLfPHHSEMJFohvjZKBhXRg
aduvl5xBTqSA35/4y5NSTjepVQqAJCphLHRA7Jd2kfRoaGcfBSceQrPf1/R6Zd/V
6RnK+xds13nrQ2LlT36+R+psfJj4oXQuRc5XNPxD5aWRK/9CXI2uU4wheE3evaMN
I6XT/XxLcl1xLcuBj/xbBDmDtt0T0NJ1dhf+RBriQlMSVculpVgRtqQ87hgEQH6u
9SZ+zYyu4ldoiuRmOWzGseoOA6zv9t27nTBFF8HeQ5zgvgS5/imo0UHXYEnUpbpV
biU/LeLEeTzE3oQk1TWYxL78fMFR9g4XW44khStn/GRkwZ2hz6AmUHrHd7zqoDdD
0G5lAvr01TAkwsqlcAt7eyp2WT72uXI7btVnzLx/O9bADW98lsRHz5GzCt3dnKbo
WQlUZMDR2eyva9zRNHr0uIQ8Y/SgCiaXFp5ryKNT2XRH0B/XhhGOlv6EvizeP5gV
wr9gOlPrZLeSvTNoUX3p6Spdnbta39lZhHhN6cb/mu9cNh3QDJ2x6U0KVzzxbBmq
KR+2/8OC70gx6f6G+1S07eNgsxTOee+Ouhr602CX4cVSwvuwZctiEeoSiGvOm7F0
vBSvERma8TO9mPq8qzEmZa7dFRyW8cEVbxJxlhn54hwOQI/DwuKqa3fRc4l40kUF
nFh+bID/LslCUhrw7jv9Urd/fvzC/DZuvh85kLhThd/X0oG8F7Dqr8dFsjyPCleT
KKgFzrtTVMIno3v4lJnXZ2LVdIOTXp9aCq4CuRso/XpicqmZZbFTog0sXIXcrghA
vM8SUKUVCstWVDtJmz0HQ8YRFMcB1f4SuvYUqvXXOtyzRZCzdFjCmfvFiwYw+ZM5
upnnJPhXWTfFsXrl0z/fMR3VrY2TnC3b7sPWdy8GoFHzB86/ol6IZZT65KL1JeMB
885ybpipYr6NUHbBVC8Ze8j6y1WV7nWSgUrzSSG5jULBqCEhpyMba7xHL6V+mAST
GdsJ590Ouf929+avPOBX/7lMMeKOyeaKsxJ+i0NwelwdaH+qcZZ8vqGHUPZaGMo4
SmEkkSlWDcO5A2XmapyI0OQhZE0icCtSutsWy2fPfzpjR1WJdTnFGRD65C5VZWYx
iwXOV3elJAuT2pVopuGnefxVfoIRjXLa814ODpf3TcwbLeBElXa85Nl4aRnyv2Fi
JWIyp8cB/gD0a9UPTAi2LhVUvEmPvWvo2YJ8DqIaaIBAQNLYnqFJqade24xJHxZQ
+bXgkJiYiISolEq1p0i9eTbXofoqB4ZsMZstFRfwaL1RlAJvZOpLVdvPVVYeEla0
q1W3vJgDnzSs/KxDlD8QaT/7J4xmfQyi50E7H1wYuuIVpm1evmgXddS60hvg8IYQ
c280eiDlROaF14a+GAhm6B+JqZ/4G4Gv6QR02c+iayRVmca8k8G/0G6N43pVCaCt
Jo3o4EOLLZQ4rPwKDXQlZrh6+dvWVSUqO0LUXaTQ+Ca9GiwnF4gNtLNFHKsHI+mf
ddC4wyTzWmwCSxsBU3v7CoewWSpneW0rqpEYtfQgek1DmG6DX7eIJcUSa7r9/YoA
hqHihzBUQrF8LJBXPEiCGfKWUqG6Ut+Y/DhJOuXFAqeVl2ep8+6crabLkzNmFfuL
msKOhpbHMIk3PehdP43LIKPKKHq3dBPie1J0cn+cjepLebxHPIaMvX47W9ugZYyr
/tWRAnBGeDSyVcQAXC+qRMOUhO+IMjdndit9KccnN4cVwrc22T64mMpOgWS6KqhY
uveOdrJaWwlPWeUxC6KQH9WH2TrSAlayPNlSCmCB9jr1kjCycpmsCdaSHC39yuNu
GNZvZt8lPhhlTElnf6TGQ1YKcO/N8g56T0rEFujz1eyjWYOaj7hOBa+iNGJnkcKA
P8ruNR5iX3TascXw1avFYFPWz6OjhnYE4fvHLen6qctZukL//psnTqGeZoF2vlLK
UHrEKg789bCcyDLHjbhRmxfwtSAX+5GsyC+tggL9kIn33UXRnOmk/G+0wACZLYji
huJPjG2IP/7HpeVjE0rPd77H0U9G8F3qU4ARd06a0lP06wVza/bkkPnTkTiKpSLw
IFwONVUKwZS+WQ9iBxuwVSlcY11ekt+JF5wLdDnsQ23+dsWDqs+ameWBekWCusFf
KBa7lwR3TOXTOJ7KwqYLBaQNsuq50FFOip7pJVzAPOusDCPfWC4R32Pe76LUpiGr
4TeNzwynoN4+dt18pSM4iaOT4pAEPdGfrvnja7f0XG4p+cuAdPPo7MBIrO9vh6LC
S/YAq30FBsrOKkInopqUQwuOseBHrOLLf+VWvzuv/lcAih27/H/2gaiNopKu7En8
cX1oKeUO19oz/60Jrd47y2x/R2Vk0FbVyWtHKLiCJFdp7ao6sEiWuHvg0/njPiUO
RUKry4Stwxaj0+sxZ4SyH0TKleMCbmK1jfSY8Fc324pUs5wdECkqDD3VnPvog2EY
Z8OGwtUcte+9QNY4Brf3OokSlpspYeUSvCcqxeVv7YhxK7AMdOOB9n/Oy/d4/B9w
0HvN0EgceYvn9Zu9Brm309dgSWyw364PvGcLFT5GoIsgvKn8vzskjAiUVGVLf7tq
rpIcklOK9MpPksnxHswWllTE3Oxs0gDuvLpsTZD7COxn8UOtsPKUqxEMidK5k8KS
ziZZ6azswZVadwasg+C/sz6RVQvVmIFxZ6vVwo+792rmTCKo0D/kbjmIPCs5Z0it
qyjKzmhHFwEH92EGeeVd+1Sr+qDhN+OrJ/l2Po9kUCVNdzciGyqOSE4X7XTRQBEh
vhOY+xBhh2gtp8likD5F0U1hmgYH5qxwdN6mtqVkGGwuquJlrDtlDvqfg8axSV6+
ZwNhzq58zSDO1K0yNHcE458fEjuDubFtRMI1l9BkElkkRou5VRa7Hwv7Mi3OLN01
bX/52kOJwlaVQPKdK1fVU+Elw0cQKNxYHrdMaInGdteAzqazeiaP968jvvPpWVix
1n+KzlWuXZvoJi/Jbd56g/yLA6v9WnHxXvJae58OPMVN+QyHxvcI2/8OnY/3M+w8
uSOgVY80ph9WZREAkmbeENbU7ACztVGpgYTNdUNNG4b9zHEy4+cPSJEcQkrFchKG
+HecMIjKm8SiuEElYuSs3XAXprl/S2uiB0z7FLAp7VbecZAaZ0fET3FrpZfHQfTn
IFnl63xWro9age0cSiO3puRyjOSNBBxXzRmnwt9EgYUXaDZSr3sJd9U5LuYi1P9O
8EYYmPdY5/ZwwBWkAhaeNYQuAt/pP4YxpaRYR/pWoOPL/Fi3qaEJbblAwO+1NlmK
MMlSoiANmvXv/xg733uY2pD/AeZs152RqSxOK4FzdhXITd2cL25gI5mJPLVIT5TY
VQ4cK058Ts6KAsnk8Zr2HHeM4ql/fmgM35vsSyp7yCSzHUFrPeLZmFAnRQbhpXJA
XOscfZOnBxMr/ycwM7hqsYOY3MdlkzU0vMvaULeqVk6bMsW8IOn7PBjveUZspw84
I2FwwbN+GqWCKjo6YsWXfP/k58evGs2YbJbErAgWuAsRtfBTJz09Kb9NIUWmX+BT
/IJgK4hTTwU8f6DPNQyO5fzB4XdFy1NkfovomdWo0zpUCUrzKe3Iybo6JM3NsV+Y
zbeKzdQAAPI1gwDfGPbwX5C66hCxSEqEQeUuPFkuXUpH91kvR+SceGTbYvwN2/J7
qQlD3j4tu+pAqje+5utyCC10edGl/M0d7/8mFiz1unpNN4RkH2TZA2OSJ6Zo+yUp
4BSiL4YgM+/N1Su0GG3ZAZtIBlSGC1V8JKpCvDAH8MmLWTEdAqIowYeHjRYtXWo3
VeMF97dLM3FebXbgyxq8sNrfjFk1eRKlK5cgNxHBQPXJ7n2bIvAVU9rmDT1L8nyv
gOeMp1808laSN9zfJGEdVH71UI6GHAsG2cYz1cmCHbt8O/lKxxZpUrvDF4PyJh1D
69LHJSuFfVyy1gBRJa/ntVx/p+Gw5SH8nz5aMVa+3IDxDYvtYSq8MdUx9dN7F0lj
4sNjvKDADDQPKvWMdsq1vPp94/YJP+w2YZtyUtMz6W3X5o8lnt/49AqV+ExV14kv
e2UJ5T9RBPEjdaYZ4KpzM/MKEe4hhC6NJraZpYxfI5dKQHHFjZp9sx4sgw9DL5e7
1OIqO+LsfcEKD13efpP28d4zv3wx/qu/CV9W/fo6vqtf9v7P+30uwSILu0nRqakl
Vtq9RWDnDZHd9ZD3IXqRw2rqFSvHFAlDEs+Ae0HhFwv8ATId/iONPIXrQOMDQppN
Gw7lj/KbDUmIXIHZPhOk2xknM/E+H+3bNkEAyGH+YOkbQFonirC/RpdOwr3W9kB1
hWUAK8bLp2tUmYIT0KpACccGkdXJU0abv0Uo8CU6bZSs9HukboRAQSCLg5zSKBSM
oynrkJPnV2EsDWJvbb74GTciElLEbTr0UY9i3757DDQd2HPpAVqaDsGQVnRnfzZE
1xIFe1X3DYH2cirruWp0QRUcg0szrdA43YiYYOrjZa6w2N9qfVlKV4wRx6vSEDxw
yT1wcqm5pY8NCAvfZZJEWpPWx/WPjVB6In3Mss0WYujTLkrRB2gT7jJGLP4wc7q2
r6Pjk+q9mUQzhfOJCxSlQffymMC7qy4YF0yey6CErLnxZX8v3RoNggUC+nD2lJF2
+hLWpHBYG3THaQ/2VxztApt+clYmjWJ4LqO3LDwZ6l5SWB54Wi52NJAFsSBrvMbp
A2F+ig3Ij030NlpCEhwU3VPbx7Kj48L8Ygix8wua7UnYUHnpjndYf5gL5iPe6b5u
/t79a8kRAFIFuPzmAba4E5/uAeJwSyT5t1RwAWlLkpxQDNgOxSV+9D8oGqcyuLMS
UlMIH2M2Sbyx83CkbyYQpNBmOuq9AqxiwHwhHNcv6gC3eMoMfO2dTpO7bQJnOeSg
DUG25IzUVKa2/1lD6zJlgk1BvEMz6B7R7zJ2tS7I47Ve7lUiR0eJFmIvti1FW7O/
3xSNoBVvVqjz9E6NElPmScSXmnmAVI/OfEcR90SdInZKEgQssseKexPLp+TCY87l
AcLkYFMOuV2hxSNYeBz343qjae6RI/AnaaZLH709kcgTeLRgaPZb2jOeNDRrZ72W
rFigwqt8L9FGnrEiRW67GcKnDyTJuDeGb/jtvEGxZSNR5OISH1EnZxsrID8nsA5+
Bovt6kB/W+PD7vszI9fgtuehtDgZ+WseUIq84jqKkNOaFxlNVIGJOiaH1KTXfbtr
YwQD83m4nTyGvRFqRH2ZO17GEBoKCUvIxGVkTgMetcBBT3kHlNHlHj47Iu7XvoKW
5Ajvr+8ju9EAfweTXLZILTNvYoRGIGHUN95YzGCP8UogAmzUbHhhd2MWCKnZ/ZNb
BGfK/22qZ38mhsvdA2JD98fk1xdz8iMF/UmALjYjJDcpaALkUkxwqugCqnpOPIW8
jhCI5elGaqUHqPNQ+hrg4a3nST7vjPuAmNeBieZw5i2o1NMt1arbXNQ28xhCXjE+
ae6z1L7tk/GxNcOKLvT8cYxD+ky95E6rz8J5Ybd965wTFZmWZZj+B+PlFAl5PXto
zFNh1UUJn9ZSNsq3h0fOawTOIjeQQoukfgWFlcx8UKEE/PB2U2R4l0wvlb8Uwt6r
lLQaoBdK84t1ht0Sw1xFRUxG7fj5YEypGEXihX/2mtYFeTLKqdYxpOEgb5ITCm5e
qyKtyNKHyPLRpIHIfLF/nVjKp8xS5ap0n4RdtRsBprLT4crxMjriKFlrQkNm7kab
VtKPv3bdrzd0uBwB+EJQyiSCyVpjOOZ3PfP0XkNpe1WZao2hl40aPErFwSHdwfTi
epHCr0Hhgm9qaXEP2hbuEpW6HG0lHj66eTIDh9Vv2ZcLOeRwx9ufeFQ3UkuBovWj
QuChfsEH+CVIHimQMU9EbkT5zyHIj/nw1Lm4zC8rwvZcnXtTq/Ne9kScBiKiAI1O
tp243WsAok3tQWyn8DoeSeP0YUkfKEwOWj0ZurWehYb2XE2BbT++bxmJnJqCULa7
6UIc8ryh2kV8fktZhkrqvA8/v3CBFrZIeRELqjTyYJpPWc/zRQ/oJnqVVICLpkBV
FcP8uo/jo2nk/XDgZl0d0K/NJkYblhLghZP3bQoC/6BD7yENvZWT1xuPDNdw6nrk
3eDD4zrvR9XAAdaEPJ1aJkpAotHmAVDrcrn+ZFdY9o86aJcXbV9lC7sso46ABVMW
sQC03ORzpwcdPscIC0NAtQ2g5riPPyXE5/2Z5ychdmEWie1Wb8Z/NRJnt+Tb8GRW
L39eIHEK+sz3KfMU02Q8QeB9Ri5555qPp6Ld0wWq29aOfyGUoKeSAc77MPBWQdk3
JkCWaYqjCH+260XiG6P2d0rSQR27hB3spHoRyl4LjTxOT1OUVdT3N72agatUrzn1
Gg4foeoJtPMqVw0nEk0Ys6XiR7s9bUpdI/7dwAI7P/lmiqkhj5YbcdF6yCZzCD4Z
ftpd03cx4S9KnplOHYXiaHJ3GQSI6HDQx39Xm0OdOj0JhTChBbGq0die/gF+OPcH
mV2A+t28/3FCpzhVzF81y9K3iXPAsWvgRZBxmlFFt1aXNX/3hwFYiSx9T8g6LCs0
uJiiO9KOxzdAq9W/Te4YVZ8GLQcpBAu48HOlmZHyrHPi0Uc/JIokwEa5xruIsRgC
BPizjaCb4XM9arn4B7YWASnjOiwhgrpbncRAz4d2QION6STDVlGVwwMeFmMT4Tbp
oboxrCVg60RXc6sI+ZKXFmAbzQsBpbB0kA+w4ad6kY6FLTVUt7tsyYWNmgW+Yhxr
moWeYZd494yVnE3T8Y2kJHXjLhW0byyA1Ji0HdkTtbxUB4DxuQ/GXEBmOseuSOY8
ySlZCh1wIPGFGHo1fFrjMxx/ro+SnM2DIXFOxK4oCVnV3TYdSUwO1wfMywp1f5Kd
4fnPKJSLVzl0p5AuU5JJwnLMv7M8Vp3PlPgdwweQvx/nLRg/Lx4XQEOoxJ4w/Nxk
lkZwzW1hoMPvnxyoYPnFQy2J5/RLQJiVjLfmOtNyJ8YvjJK/CvjQvg4YJ38fVzLi
ycy6HNdNaJjH/IqjzXieJmq2SivEGIhe3mBCUDKpMXX0PRj+ZCXHZTjhnU1SjjO1
tsQbOqY5+PtaWYvX8wPKtKaXMWGCUIh+CihC5yj4s3RoHl2XPA2pyDMoLwNB+sdE
AjaiDXjHo8qUGmSRWjH8Qpf8KZzRcO5UUFPaL05/6xLichfbMZ4IdDeQMG8ZtSZa
Etik8M1juXxfMXFAgK3rWTCuOM1W6fWDZjwK9627vVopYboKR31WC+QYpgBu5h3/
Qc9Jcm186U0bzIPh2G88PA3uR4anClMLzhGfcD0Ft46SUdtXmyoWUD3Tqc/Smc/G
Hy6+wqgyRK3zXJ6JbzBqhXA3ifTxPEjxcKuR24t9d2aex8Gp5MtOZ8s9BzuWDit/
tIu1JvQalX3V7H8j0UtoZaHGSo2Pdc/ZvGOylpys0BvuOSpvdoGdBG+oY+WJHPPJ
a2gv4JOo97sRwcHhTZZMf1EEs4Uc0gPOpE6A4TMybpx9HMcVQnlabBjTqsJLvZPK
IMKU7VokyJFVCUG7JLj/Ggp4wCOTqw26biy2z44daH4MZEj2APxGmFJrqM+MdITJ
13j/MU87C4406iFzIib/j+cbYhj2bjvimNp7ZwsC+R5wNsPWZ1Z0f11emm1EeMUQ
4PWeG2s6qNV/HuPKvisR+IX1quEJ5t6PLbbLveZPEJoch3EP4ZbTFeu65dsOBuKv
0c4yWnF57bdA2CsiXuMRKX69HDSTN1DdlIrE2+zxtLIkyTwm2FIYXnt0LAstD6It
Pn9rPR4xojCj8tZ5UTJnogGCOgRyXjK/NgVdXkMyU5JG7bSf+0MCr26ddQLQXwvb
V7EnE04RBN42xJYzaGm9PB2Kdj3P2pTIy9PiQJ1c/qwi32Vnz/kw54ts4RiOJLqd
gUr073njJAl7X71LcbXXdHOyesfBNMtBlNn/JKiHayF4pJhgFSOMHaXxiTojCCJZ
mRxu1peiGniQQwgs7S65foJ9LmzMZ6ztfDQ4kj4tPVSjmMe0Zaos2B2EhIEClM4I
VaZA6nrIjCLQ0yMD9igjzvBLsBDdD4Wo2hDsOmjxvxqaRmDZiBPIK59PtXd2Ew9C
Jy1tg4sfz4YOKHbyzz+AAQi9NJKNsZLXrZVJ/laf8qCSlEY7ao1H67ACilg29gWT
RC0pjcjvPM4/Opc/OY31+eXP9r30+W2g3NcJWQu/Y045/aqQvTPVskQC5/n9DtET
7P91CXC65RnZXScZk4AkyGfq5+4tGKl8QitjgEo9lEc51QX05W9f94hzU0BgTmG0
00m9XJqpiyZlq8sLbXPRx92BxhkiKYPozJYIBGo42Nl+AgbmG/mF+EWa37/JXNN5
INt1yWnvJvMLkzALY6BWVG8Ox1/iJSmBko68zgF0sxIVbvTPh0YvWsJdR5PSVUvT
yn28tuCFy0qMX6E43BpP8B77j1PYE830ABhdYkuU//2FdFYbGgEcc27tM0kdfDeu
SVBIZUMJ6zjb/OQ7j6jJUo4lTSUp6p02SOpLRM83dKQzUrQlA9QC8DtPxQGSHHVD
89tp2SfmA8NNf2LnaepgbSd6jQTS5+06RbXl7nvBMCBCmI3hHaQvY1F/l0kVQKAj
oOuPkhclnKl4JiFz+Nwu8U8FrBUPMfBSxQgSmwXpachtuJN1hV6YegJcLFwCGnfW
Cwbw/cuMHcrm/kGvPNuo8c4GgZZR0iMC1xdIZ/URy0h5XJuapSr8+mxwgjydx1j/
G47V57f2zPA0Va7DLm9xc13SVIBy2g5EwH8RhzplciM7k2Ftq8QAx2EnawddY1RX
snbdaDaQ7hW/ECZqKtiDa/WFO1NBRNi8V7iv+MXpv6tHctb2VWpIene8+67m3uYv
2PyfqMRdgKMxHdN5mtWAW1zp2mfqpSAuzKCQEIF3FK0w5iLpIfMCh9jp/VQ/pT2Y
PQQl7OnKEvMF4oib9KlNyjlSZ4tr6UGU3TOJ2TpK3hVTKwzLRRqte9Dhm/5x5D+k
8XFF+QyQeWXr4iKeOlnsm+rl0oEmvXwfylQ69A2SJ6BPasK5aCYIKyrbwDUrM+1w
vdSz2gkWCJ8RicUe2h7aNp+nxtvItSUWqL7Aw8YHm7dfMEJvj6gVaSwpVj8sU3zx
xAz0MI6Q2yRG4H7UYcsnl7gEc6BspQkTtg0z1ZCtyBm1PUwCm2EqGNqb8rnGG9Tu
94pXDo6mZoKwZfTl5zK+wD2Yponto3Bo8cb2VIegzPKj79QzKl9HAlfnF1ha5RS3
OTinbSJTlpJbX4epGxeC8XkClKXIjjJRGKYogSm2+2jyfX8Ayp+0EGjV8n8qkTFD
71VX79ZyT5IcqE3tDTMiy5ce25rA1xfD+Fpzq12i67sSYFgJBFoBx7AlATL9xJU+
ytUiw+iwiNZ79viKpwdDfTa8eYGLwL1j6XJPokJNiymmvP4w57QFMmTMi54Y+86i
FjtRd4n/5/pV49g1NCzdcBJ/HoeJA/vY1NThswp4VpFreFb6nhhgxsyKk6CFMrES
zsSKMUripAoYhXJDNtjrGvAJtX66jWKGLcTl1bIjnBFONYNY3tXTKTZj1Bbf7epl
q/NSDVvC7gYyRKLOA1Kq6QJnpJyonBSwC5F0wo/E+PWeRm6UqCvMCIY6T50ax579
dlKcIzPraMrSsWAdMrcHgEQ0IzuaqBzBBVYTJyQXS1GztLP/qFqUqSSapdJ5Da43
Z6OWtaa/fWIFuLa+BqMsNo8Z/gw/pvaOz6bsLqGP6mbdVrhjWtZdH/NHRnRvHMG0
gkuh14mohY7TKy9/zOYnWGK4UDb77cZtsl/bl5+7X2pluxCARG9r5fP7rKasw7cE
YgRkDFghgxPNlDIZvH0DXbHJiBgS4q+n+8uELsv/4EUurJghTOBtxZsAGUstxQE5
cvNeM8lbKyevE1vMHPTH4SuwztZyDiUhreZctRRcFCqHHTeHD3/LcZCN+r0b+qFL
WJEsksb7B2aE2W/tIupG1051KxxgIYk8g3xrnoDW0S0KVq09qoBrnZNZy3gP6NPb
/HZMvr4SNe6HIQDtuIq9ETVIDDD1anNinQ7QM+iuWFFbn8biJl6ybgiroe0L94qI
xDLvAPY+rs9K/SDY4T6cstP16NO0GJQFbMTj2ax3jkResoxkZzZ9VeBAkZCeEAga
5sE78iFIs6zDGeTGU8CmZpPVIAakDrJcv/yR1LtKQGFM84NHQFqEEgC6EDdeqACU
b6mLHOkfaaeilopXsJjqky3w/UWXN3CLg4z0nC6C5byJeL+O/I//eaCxZZuOTz/S
dhTBNieuJXNwsjxeIfITyhmnCyO1avsREL1PFwO9t1hzzTD7LFBLVDH9gm9cVhFN
IASCYLZW/HkUAO1oLFaTHHGhJip/gZGPBavQ3NCt12Fd8ogcQWJmdXgOvmwZKJSf
IlrA9PQoBOCs42E6jeC4X6WkK7VT5ccO1KejEc9uwDf9M39V2GjknAP35StyDU2C
QDGUjJtoZshe86xI6iG6K2BDqNsIiaxwH9YfT6amSOlsqduVZnjUMeynVTgtx4Nd
t3xoJ9bWUTEYMe0igBmB3pQQ888QhbDyOtCK9WFZ0+qn2VPPNRrNJ4rJwXRiQaPQ
DCCroOiT/FstvXUnwEotw5foqlKkMCROxAmcmhuRdKSRQ309nzpH8NVA2E3jyQXu
CTz5u7sGfQTGOvyLEC4ObBvMOJ4239GTLtTy+hq2roK47VLSPcTNncL+Sx0fOY+w
mDePbVcp+BNrIcL3I/wZgOsJSEozAnUz/vfnGBrB5DXwziM6MXawWneTooIBwxqm
fU8zy1VLMnZ7vC96b9W89CVQ6C4Fhc29CCaJoSA1lkPuWJ3+uUPhNRT7N5at02hL
EhgDSpbQ+coNedELExFn2AUDqnDLJyJexuGtmPq4CFwOIFVhMtr4GGVlahanszA1
V4i3uzEHJTx5ZRXL5ZRhqE3zGLdATU+0S4GFh8lmH3PjbDc3Y9fKnZz2jqO2/Jd+
OhnqwsEqF0RZY3ZvCNtarjvH+OU7Q6cUMq9ILkPpCP9IJzvJ1PcdSpx9m4UEOdju
R7tO1BeWDESwLMrJAu8JuzpSlFY84mpAO+bqnbmno30WWdpCxAftBRgYjfNTgsaO
++lIvlgcPiTcGcWruDCuDQmU0k0oheOqhIoVzzySqO48YuFA0aPhiy+cblcfLv8X
HmnzIDKVloF1Nbai4mZVDWbhbKrV+Gzacl77pwCCKYc+LA4ZLT67fPcc6umfE/cM
dgU+B+/cY6uCJS8ROpyWiESkidMZ9Zz66L2N5OqDbpBYz/LC3QUPlW2bOj0BV5T/
NcZtvHswXvhxN3ats8585J0d7sKWSbWLariOCZXTZpNpmpcAmG+u1z/rKl4F2Mm/
x0aM/8QmOtSnZdlZjJDsHaDK5p5ek4I14A4J2Cs0sOV3R4yGruug/S85AWMnELz0
Hw8r3lyqmXE3xk0ww9Nt1N00eET08uxEZWdItvbR47JtEHtH3VZ7T51I+Z0sRMLZ
LPrnuZQzwqHqJmT9Q05EdwhUJnEQI0JckjrRn9evR63YK6rB9ZXsMHUukuivf0sC
wXDQKEiZ0XderWJAjsZfdyKIrIDmGK4AY7v75nr9QFDGlBFEAR+yTspY46ZhCKUd
TBLy+ELBUrtLO3J0IJobHWXAAa6jXgb6/ZRYMyqlMARJrrvCV5S1EImL35UXWmOc
yLXNaqNtpsxA0qTjDMQiYyEZSBpEA9cMqdlwgiCmu2Y4uLeZAJ1DOC4LyVNVZNuF
jRpy1cKmDRDVQIN2YhaPMHEOf23DfLufix1/uo9vAv+pmUcsptpYpoYanTmJ+VtD
iHWk2m6a6BrXI9qKQj2Dv9XME2mHTBlca0NonOq8tqmsrPdA6Nz/OXj1bUtnYQbB
TMMI6uhNQyt4OwvTPuhrdOef6oHAfjEdg5McGUaqwR6CVXE9IoxV8hMkPs2jATon
O3sBMrneyfPj2BM+3WV/kpFpfPsSoACgDyb2kD/MFgbeJe63IHHF1yJkuCAD3drT
QqlgyZ3pcnYwu9CS3IjxVWmvpZeynvGhD9ZErHsrDI0voPowQPtwUaT4mCZ18SEV
Kjqb//OGzIiia/wUaG4ZTctK7wALNRiprvncmdiRMYtam5HX4c7TRGFroCVWlX7u
O056jZtGAn3w2rYPQmo3vNpLOXsJQxou2pjV+qOcyyXhHzc2AU0TpdWnJD8ouUu+
rhhGhxtDXUKm9vKTr55m0ZUYBFDxawunk00uhp5bXbSezrKGOlL1X6iaGJBF6EoE
269goO9bVQpCzHBt27BTmrG9pD6d4HoXy5du81ff07JPhUa9u1RF+09JRfSyNUHW
x/NsdNYrYJIEQkwjetdAuYbN+xpxwOL1qSlIFicLa8BlPvtrN2ycsBocqipb1h5r
NZBCEUhabD3GfxXcTQgEDSXTq5/etftlZqRSQQbAqDbxXR40xq5xh7/Zr8z3I4vH
XCTN1F2xjRl/jFDZ48cGG7Vv2a58xnD/LacUkeJoJW8smQj123oYIKAc8hs+qOKJ
9rdeuxuTm5QOFS7AxbA4/1dL5NciIxNknerd2sErByAHnnxi0DwttDdekVvtqJ1K
cNU/+t8C05Y4xMWSM0fz4VdEwWWRV82mAPNo+rnVh7eLpgbkeyqp3faM3ScaT7V9
w1t1icXYvO4aFMGqMN+sh2ZKxk+GJBnt+QX6adQfzCR0n4S8WPpIwowrX82lmPsI
wFP4p1qyUwhRg6DzW35zptZ2Vtw/Sem10xNvC65Q/U/fD17nig3shRXCazKQFXM8
iZFUv2/qrVi1IviwAdFT2q7rqNohiiuyWpeYMk8+kDRRZPYhFTbllmKmp+vrYRPL
+pErxgDpZeowbWG36iPOK52jdWTmjpY2abJW72FpI8mI1A/Cm1GTlOF2ZJw1o9li
tzKeviBW7FUZaLcj1qpjqGAe51TVvX/ORyaQuqxqAUnJIPrx3jbqv8O2XPVDTNW2
6h2J7BiG80eqOJN8iBtCx1lcA0ARIuW3mGN8tOsbovl1WR9O0lKKowybE+c0yYqU
Y/e5InJAAxlwuLzdn/TmullR4q7JfHi636PbVpBLpZsZZ6CxCkXvp4B/ECVukhdu
8SoCgkzYz/hU5LESdRDAnBVtg0so6p4KrmJV0hnKVxkFVbeGcMRTwTl3TsVi5Pow
X/DX/w1iETXDwNO+v/vVk0l2nl7QN+XRA2blFEkOicrYedXOPomZ5w4sweZgM5PX
FMRBQC3v532AELwAOTp4wJTPrsjsBuiHinNWcUoYQ5I+N1D5Pgvzt2WJWrT8zfP7
/oGtRHqyVGN3o1esjKnZYVk9LCqgGLNmUZEP/wketAxbksA7X89d8a52avX96ldW
3uNHMA5I5MjESfMz24htCY+DE/OWZif+9ZwmSdGAOrV7gDrgc3H9UJoY1izOCrNw
tPO919tnMbIGcf/KTvSl8+V69LEV9wcZ8waLILmy0HlHr++z8qw4KpNIulDwWGCo
uDdyfPEtX580dK1OwZzNulSxyr+QO519KBNDO245TAbO1PT26iNtEdflmjDUW0Hm
shT9t5SucP/gYrkEmYeUJYb01KUmT0RAQcoA5cWIOBuH3tmdasacSZ/dvXc/EPnp
VO96+/Kooe5JPOhPJPm0LIW/I2RONoB5+/LZ98cXXP80+iwcRVMQyktLEbDHRAMa
nFQCy++GPsMI6QzQYAIA1K0/nCkk80IjC2n6ST4Qf+y989JRV4beQRrhluSnMdh5
r7tRdtpmMweDJ1Fsmjlk8yEZhx6ItAEKZe5iHCYGi7JGZ8Nqso9fJwkKzqfmd+/z
ahK6RGuZUgU50P6vVUOoxvuavViYifpc1isdGcIyoq9VwQwjRnsQ5bUD0UjJI71X
IHXlvGi0q34wMpS+7aOK7suMg+w66HgZT8aSkeOgQfQTZbWW0YIL/etoTewKygHR
RAd7emNqXUZQtTIGdeXfbecyosHT2WVjUOJ78kvt5L6MDo8iHn/xZQjE3Qvap4oK
ABYcaMa+1ynssnMsybnITKTWUg2pfXtcnpre+BVzDkkJF9VTaTCg8OGP6BAl16AN
zA0+fKaB7fjPBiKdINdujtJ7ZXS+8bIQoA2J30yxDz8VEppxCe5+vEqcMsih4TaO
H2TErwYUr8Yckn+MIQ0FCXB5bK7fWp+kueVkulFCRjkZWJMk29qk9tvjr5/m8zBY
t7bNwTwgaAYr6oRgBNtQxZoz+oNqbZ0bOTRDhry/FE6PmwrOoB0zD0NsWI3P5poA
bIdwu/Axlwu66H2RwhM64YPe+sMjtD4OSRLRuM1sSWMR1IKLSbjw03fB1ZhtRA2q
oz1cF81CjRfbVELRhx04zIJ7hLkBBjbHJZ8qMD1OPVpTkKKYmquKj0y/lXk0G6wA
8ncA6IatvOUy/GL24tYTYsVWERaHhx4ZprnpWyiV6SbZoq2oCav9albZCiK/LO71
2MpAmrIXja7keS4sa/veVZ4gXkvMK3siF4dYTmy7SGwfdL2CY9WJ8PL+VJHWoGC/
TnAFFKprsLpg7qcfhclT6ln8bRgKlFXD+bub5Ke7VPnK54jmtCBl1R+XPghLPlmG
sycITUp0IKqNw4vhuSRUbEEMLUjaLrh0ldk6qPfxcv7YENPr4oO2QluMWf43MOv5
fjsY+mENpFzG/arAvtf41hS12PF3C3t1p1mRaESHo9W2fA2KrFwcovo7nnHb7YSw
LbYD9m+njw4ulGzWYjBfffLjyfWgBtXH4rT1bISrzmkUj5naBIXOwHEzHgLm8V/f
akp3PNm214X455gMJcRDorA5ai5ePJBIP5rRbXRo+Ol5PYN8+WKayG15i6Ff6j5C
qaUmTS0FMwL+BOtc4CLYBsng7lLNQsnUaUOMfhUOtjLDs7wbbh03PuDQ1QaobXq3
d1uugAZF4jcSyRSav1k4g8u+uyp9y5tDyPzbVPq1e+pNwHygMteFVTNifdATp9tQ
Jvi+ymaniac/e70jCoKnvYTdO8aBg8KjwwqepTToL9afF7nKYQTayWtp0aYkPtok
m8xV/UG9VZuZqa+1QHD9PGN7pFY+1i2er91kW2ZJw6QwVkyf3hwGtmpyGX50xNvy
LcZCmwqVU3kXpLvI1iwCMqPodHN+Uf7c4BjAgRDH6GrmWDcndMd6Hfjsrs3ntnyr
GOm46aEJMnvmbynLhcrx/SilACuFhNX5N925SDx/WwKexCSdU5mLiC4GTI0uHe3Z
i3PxH2sBqxMezqS2QQn6U5M5Ww4oqk2KqMN0vZHD7MyzNfSDoV9zMEfL4F7mwySs
JilZ2f6xhQUr8Hjgrcep/WiNA9OSHeQ30Ins//136Joa3Z/zS043Kw3tjz5HMfGA
mmc86wG2lbwAZB6++QfnaK5Nd1cZsJDjJwny9AzsyOVsKKaAW8lvbM/RW6YH6/DI
wIo4luqLRWnXnHFz9quyY7U+i+qEIciVMPnAi6V0HQvoPkjO+lXts5eNm97VQOMN
G14iOyEJR1jCfls+XM1Nvk/zX7c2mcjmvm9qr95HNrol54H1NR4HmQfSHTtvWNuD
pn/YREDBULcGlVnFhmRjrcw2JOSRcuTGX4SRaBSTs2jtaMeNVzcx7y67HIaVQWEC
pZAUlKT2jfA+fmrjN2b297zx1rd696rTnqYmiT8I0VBN8CvvyXPyFzOe5+XQldiT
q6Q3Czfk7c9kUzZrlAPWnaZERWYpYvCTrw4mK7YfVX4QZhjs5vzE9C+iP/CVBZU1
WJHS1gp1jSnVP9ZbZsjQ5RVgJoM59n8jpoBDJHj9kIUGa5kGmn8mZfXPufFkhQtG
NGB8CId8XBCnCxxNM1pFe8juI0sdQVoZ27lytXJmxvgbcHE9iyjp8Gj2bHC7EVId
CtW3NA1kRBfXDf2mK83MljUsDeWGhsFtBu72KSb0jfiOSOgLjBPhbH3Mbg/uq7rB
Yp3/v9kQWW8GhGw+tLCIdSYz4DekZE7mlg0LOw6LqqGbFaY1k6GaAzoKREiyzVqQ
4zGhvlAPAgOp5D84FHFs2jCMOAo8IqjCQvs4v32eE8kipdfUyQqC0YCSFyB/HIM/
dIfrjw9lGQTOVzVkdkqzxYUkQD5l4/Rt67GT6S/We1I4m++DMNKzDCIO3BrATwT/
B6O5k6+PNrhQ9HjJWpb3HC9Z1y1KCRdtWjiQIPNuiYQK7J9QvfqojvYs3fd+TxHP
1DSzCEqt+gbBEBEPoZ0WoOGDUYcPsVB/qcjR7fdhROLVXRu/1etxQZwAs+YBOYye
QnTCfOP/5Bue0q5iZ3ZE9ZQQKzRBleaDhcf5IZVTKy6XVTk01ZlGDQFa6dzbzuhz
OJdxSc+IpYy7gZaoAGHFuZqdJZMO8okpzfVENz21yhMjQGDSpjkQ4deeKCE8585u
WnTSNDfABkBo/mWe9psTpExxlUC/ssf/7pzW+y+3dcuOuE+RC9CCaV9n9tzit0y3
YYKScEYXVOfZSnKij3JGiy5HOnwYd3SNwg/MGnig8+/rXVu6n9K8K5lWp73iq3Q5
6LD4W+AW/rQ3Ds/n4e9Il+SxFhS93inrgJcFSJAyoqeMO37QI7D6OUakv90O4BqR
RMXEip8grlzAaRX7ZR2mgau3kXCi1qSdgVcyXCkANNZNV5BrAT/MhH5oPfJ4UHzv
jKBxLnrkWt8CEL2NiSwb0sY1W5pIE4eLpYKWvmSjXYKadeD01qqj/wdccA0ntD7O
gEAoYMoFS9v/c56qPt/jMMldPRxfb88eA1DVckluEVhdaCi/Tbh071SARs4suygy
6FSDNWdQY1xXpkL7Q31OQKhwyZpT/kIQ5BfMwm47P5WvCyALx+7p6DeSONq8jsjC
C4d+7gcofU9Nq+iI8AGBZB3mvMyiMk4tyDciX3msinVFdKXWicmSXcG5n1Uj4mm1
SqFWrE5zC5T1v7Xv9u35X7MCRM3azjCSo6gVgWcppr3BakfqsZyZyeX1x++W8vxc
B94Y9gP8x+25JrmpX2kU4qFIRnUNk6z49vagRa9Au2QvhFJwkkSPXiIIfcrt0fgr
Ve+/yKFKwHCzP6C8mBD/Gr5Jbw0qbRONUBMvj3kosjoeqvm41XfGGYgg7QL91Vgx
HSoOVLTQoN+kK1oxIdUFHyXZdnpRlYzHZJSoHzPibRIw73+2h55jUjdqbWPlkUzs
hWJgTYPazjMA/62lV8pa+qyOUsXwaQ2+4J3UKmSiMODrr+R2J8eH2FzAV8p3ec5l
iZcsCM4dhhNECyAVfVn09EuGnr9ACzz/7850SzW2TB0fqw/8tGDeTNBvhqGKk5dR
SDfW05aBKqTgjjV4cCQHhPc2Vcz8TAvGfQJqxwqrTyXf61sQ7pq2p9c1tn+JbcpG
Qb4UMgEqFBwiPbHa5HVtS+L2daW0sBZd02/iyRkIaINOBs5v7ZnKUsZCHKTXHNCN
nUwIKxZ2r9Iy7do/pOWqu8FbuHCVMrmV7yoRQ4LZqW8V29AGUgAedoVQzsBN0xVv
b7A6x9+9Wrg40oHe+IN42opD0YDCUbVL2CysSp9cUjfk4T2wJ8R3FhITkAGG+o7y
7ga5NkhZj+1JBOmsGpdMQIVe5Yymm5N1FCW16XA+q+s9Y/etNEeE7z5su6x4wjWQ
xuxSd8LZyhVZPFPuSpStXaJnjypM/vwHIEJpplzjbqxXTbS/XI23C5zX25APj0zg
qv1jht/2y3YPXo6DrKGjAvRL+tki8u/VLXjtx/+rlS9NrWJxFzT3vWtGeeX5HP6K
pWEBsjux2YEYPjODPCJht7Z/5wjobZzhWSwYOuvJzghnvKjAL0yATQZh6uM9VIpa
m35ExqpWP8CTjnyRZ4WKpgZTS2wzsNxaqsaKO4e9WHlR4ugs2GYHk9O4+FFQiCuu
6ZaWo94b9wDdboxunuBQer3eaVgBv05zJqp2iusXirAKErb5zZwtGjj7jovzgo1h
Aldl1/eLby5hCFWWDUzY4Dmdp8/r0YOnUz9TzlOkrkJYUKW6d9RzG1RpTzSnFcyp
+mX96RB/3DvFtvNhQyUQvsF1snbBm6Iibeq7OLpnVFwKMYhod1/Qer6gUwbv17qU
mT4vbufvhQ6wmI19d4ybMUUkjlLFaWHa88gydinPG2s6S9TGvD3Iq5KvFYtyb1Fk
+FqLKW2MIUkqe9GHjMay45cx7D9jvxBiA5M14w/lBoRp11GagIlcfiLrBVSOgTCg
rx3ZdoGyVYObDSag/+IOCVR64UY6iG7BAg1w0BrFhyLOQ04F6u5tTfE5Vqgd/DGq
oXbGpe8PVqU27GZ5gOuNYhh/4v9bsZj9wQVcIPUHQg9YrecXAw2W8ehLJWAU3OyH
y8D4rkeAfgk2T3SrAS1CcGCw9siaGT3oiLOgdL5MahOYqephQfFPs+xMu6gtboVl
EOM3TuIodQ0I8tcXosoO4SMwfeM6qlvPKOG7qZXeDI5pl+F/NnEVBCfpZGhX0DmO
ULRXr2a5SbGiqIsbtPFvIRY59Sh42X9iXB8ueuVS9PzPrNoSBBIK2f3RX65wo1Sh
xVVazXAJhfs8Ok0G7tSau9/0GTVDPGvV05tVG/9uXNSGhn165fEUVSLBDX1dRrbC
67ErjJDhN1e1FPssK2/34qM8Wyx/9VfxanMP3h86oWdu/6YeqXVshOJRllUIrWX9
TshXXdsZE/MJZ66R8twDH/kW2d71KnlpAog6lLoz54a4HOgyNWUUbQuJfMpZf5ul
aelS0sXnMtISw+LVAfDG6Iz006gvN7UwQv1yNpzlAxdyYFXl9SukvhfzlHDDCs9n
OiwNYEZ7dyRqX6E/RckNwmpFwlXlM+Wv9heXFnXjDE8v2vVEGwtX6n0yasf2crxs
mDStSdAn1ggiFt+Ozn1CySHILtA8KgcxQNvBWeb8SjJNF9W4asDg98DuNCEdPJvm
/A7sU1qxqSN9dEqi7MkwD4zSBP/Bz8VnD4KG61q9CZN1OPsXb6Cw4va9Jvdbowpj
Hp9Zxj4Td7o/E5aViI2b7IZknpefQLq0Rym2yg/mbGQsO90o8dv8lqVDSDOpHu+s
+3rcEw547iPgReiYrGhttKK7kJxuFZJ8LmYKh7Aes1ns2ju8/2GsBBjnam5iYPd8
YKVFGKaS2l4ICEFyHPSN/bHhBMiOeY5cMYGU7HyEZyCHmVJz6DvlTAkbh6lw8R2Y
Vs/hzc81oUvbgtCSNxEv1gaAzUXzZvNkAq7WzTNQtSutyu306bI9zAWfZn3YcdQ+
YD35Uub20Y9dDuNnXAomLFuyyX6XVguJh2oN9t0EWErvLSpJsK2GrvUX6jz54Bzx
XtxyYy3PUB3jyBOyXc0xeEwrwjg1izsTeDyYmxvslq73G3tBPUsROl/68qMxobNP
Qn2+ENBivQBzj68FvAbMZ38dACQD0s+/NHt2jkT49GJWVxdkpglvCG6XPzQr/3fU
QfC04JwOdDTNEdzq/lIaQms0BLYrLU24xSqso7IbnF6N5X43+dkyTwzquzQf9RhX
5FTLb5tGQlsA4+62jKkjz7fla/UjxQU6Km6kEBT9mLrAM0zWH0k4BlKAyRh5LjG9
CWB+TSYZsdzTYKanCKNk2UPfrgzoS8s4r/NAk1mjwnc3l60LZ3VbX0QJO3msSfjU
ddcY4HCu5ltu2TdDfFUj/U+UqLGmD7enpV0MrODE54FcQTtS4Z7HpTzk3joUDIEZ
3TW6zvHJeZQkGHmKHw/RGgZ/JQFUcR5eqGzuSI8RCJ9CmKKEXLm7IFzwP0VJio7Q
A72tei3YtZTgBEOdvzBTJJaw2pH3DmOLkPAz9hBQunmYTlwCOryFcOGTNicGA/vg
KTWODiw0/EsQwj0Gsu6DZdwGp/yEN/39HCHpMgmFiomDeTVAssovvOZYPiAoJR+s
OaF6DDV7TETq+miatRY00Xf2PALqs6/W7/1P5RmveWcDZMOrXVk5RRymWHaClDWn
qzswf4MWjucdyhxv2zjCkBSbqTupldtglw5WUafjf2AMbGvpMHRiG9AvuGqLC0JD
ObCWcYtADBTEAb1sHElaM9zOIXDR6RDoSDby7s8Eetlb6zcgZdDQGyiy8jhhvexl
ggxbAEdx1ei6M5NIMTi6cNmP2ODhG5lNBBBaeOrwqopQMu9PmEeuQTpal0UynKf1
2Tz1x4lZ1ffc/dxz2YsMmxvuPj5kLmw58qR84Y7MANUz/RV0tIaLWXyC39OL7V2S
wAB+kLQXM3VtIulVyK97V3reQ/b9tq5B/K7WHgVp93+cCFo5McN6+UdeEzP0zN1/
DCsr8cq7i8ju1PECIwuQ0PhWI7IiY8kkpIFawRVU4DY+cVtYtUFLz38snzhxLcpk
YEBKSunsMG/JowlEV+YgzK54QEmHUi6uerCxsPfa21ACoGlSRreCo9Lh4Svpzocy
8GdWdv+uhPIAx5Xgv/VFRX8NbG373RXeg4VLog1Ibtm2OJVXw/KLCWidxbHxRogS
AC+jus5ja6EFSkA1NvtNvFVsOX+jy6qFD8OBLSKzZAfnLpNqQRQ8nx6f5lbcIBzc
wFmcRaq3JeQdGj0Fz5PMakm1Vp8VCXJYGpzmeny4ZrZC1MlPjspWhdgAjdxrC6GH
c4uXKMJ7PlvOwoHNfnsU5Zjk0QnNO3FkoOaPadcUnfy7nB0iGXj8HLGPFvuDxoRB
bXqVuIURuHJ5wDC2iCHkbZ5euwXjm8qTa077ko/RrUqB6YD3n1ngpHKAn6n/Cwwo
neC8sqwjQ9B3zHmmCdyIfhavTLG/PXc997xLo9N3/GyaieSqVjjsrdZ6W47U5hJl
Iv592w42m0AcDLCi/qHvUs6yy/kR9/JZHeIqkY4l93R7rN3zNScxc5KmwF+OU7BV
nbeubwaCjjUMjrKVveskcRNy7kDGj/mgtpDksIeNAsmMv5vEpDt8rDQWgbyYGQb8
mSvxtNmsjbluyh2U3hMqsWmWAu2n8aCbX12/1y/dcNKeTw+2Ht2Q8yXmkZYPLSDZ
tPI2xXhkLpPRQD1qhapz+ARaYFIIijf4EuLtpvHpZZEY/s7ESygM+YNXdlNjkNlh
jiUvBQd8iRH/Dt9arX3gRBwCyLFkeNvZe3jNH8S5c/+ZgtHxi2FsRYE+YgjSnq/0
9n9TUXvcu/JmsFBfXDRl5SC/hUWGmjIOoGjo7lPbq1/r3D905flsJQQElkLlteZV
yC6jAmvGF/vIDNEZD1D3jyLC9Ar3ImUCWpgVcc/PGsGWOzjVqWjbZAndDd6tDp/M
UxRrVjuxgeLYRwYlX9XtlzC90UIOHs9fYs9N7+Vr9dEb38cHY86yyZbp5w51oFUt
QdSWMBXZDx7j5y1HeYUbTKfd7la+2pABx2JbFSm1l1lXR2XbeEyVz+Q40k20u64C
9HXThEIqbENQRYsh66M/SdyWWxOgWDula+C5IvnBpxVy+4wpZaCyIiI6Y9e89gfk
7mE2f2vGbhnwCt4Lt7ZMdMfFNe6GmCN8WhWlhKq4p/s5XLrSNODRwYdnih6KBjoU
gwrIa/fEnrW9H375uVa7skWnNmVxmXsV1wZTQUtx6LYhEgDqjsCYhkBam6GtpRWY
gSKyGLeQJiIf4G/G3gIE9qzL5AM14Mc2w5B/w8Ea7hGPXiarAevGbc/ChFdUUB6q
V0zkbllXWAexsDjt96HlWH1rsElPGGa0EL529H4x6CD+X4oj2r/ENS5sNmgiM19y
X/OmsRUm1bWgmLBDAlF0eywWVQrk8Ggfd/gepYjFM5/XCOzHq3rO9r68B7zpc+J/
7eLjBepTd/I6TVH9kNXGWAtQ9QPfiwOc1CnC3XL8QXuHuJ0hLQp3MY49zuy4aAkA
txS1cQzt0Nu/y6tWIrffr/FN0htvAaiYlkBxLvNj3WsP89OZ0eRL6WYeNUyPm9Fu
yZozZPWlwWspRwBFiM1Yj445zu28v4KmOyyLM1MdqTN1MeSKlWJW/G9LFJe2zdD7
BEwZcwWDLT4J0nzOB4dny4b+Xbnn5djTZVNzdxCF1ZKS+tWkEXAq0rfy9PXdmsmq
6nY/4874BG4aqO+0ytQZ/mWSno9VWaHapuirHTZyom9gDLgO7GTFh7AxNaV79wAR
gTC/qRqT0lDPommIwd9bG7jrisRuHdtVXVEz9i351kXixIrIbKnAXjLbI0O2Iv7o
J9qoAj3Tl+HuuRx3OySiiLdl+7WqU27j71V8cw5GxQdzj714r+tFIryhEFAdNXPR
vveM+waFOCwJgCwZhkeiuZJeXX6v9igw0QGLiU2ecIPYwCux97pzZyA6tczBQluL
DjZ3QpiCVTBqKANw4APGegA77+X84ciDQZMJ59gqOT3qnGnzQ8zGFRvMOQOOvYlV
3pMWr8RgLeL2K/slTB2uNIVj6WNQTuKXMUSGXUN2o4v0Vaq2l+l5epocg5ylgbO2
UT4aLSVjwMwK4uL7zxSTuiAnIiZs4RthS5Fg2wBrnERFiEMWoFOcHMFjxV+l0tXX
xnvJqF0CLBt3kZeAaE/iIAxEpltJAeO5tHbUfhxQca2K8AMWyOeLrrN9v6LPicMm
3czsBlruOKNUEyLe8RzMY/8g2adHUo1Dv2CdAeMllF5g/z63lhR9DuYejWXK/hhC
oZuTPx8m20oFSSSLeN40fNKffE7VjjTxrfU1nNhHTIJ/FfZe0rLo6Vd96Oc4AqkO
SSMUabwFhwL2YA12P5ff3mLBAAhlwbJyjk7gi670fSNt8iQNREHpOjo0V89yM9O5
4TAAImS+563vmlkx7w0LS12X+7upNq4AMYWChzuVl1RxV8D9N+ABzGR+039oSH8k
xGHsJsns2uNINo8yHqwYoKdzxUT4TA80PEdM+XWdqKct+uyEh2u5i3QXeLaoM1da
fOKEDbsYiAwrMhKaPSImwi8O3fw5BTpJDQ1qtppGevGo0K0iyV7xXXHXmEHYCveg
ZxuV0Usa4ghFbJF33w5eQu0Fk/7jMkN+KrX4BADf3LWD5sguz8JdntnVyeXCnOo4
awkG4M4iO2cRJrurmU0WBfBYrcDFZQciTxN0Y+284dP3g3TIwYCnRtTJcqirGqlP
G6ghL2cp0MWja+veV3XgojtIhHOsmlKPaF4uGNJFG/aSYAEUZnMvkRw7Iuu7BDdf
HkeaJbatmopsu59ls2Ibw7t9/5MUtoJZeO6qh5cpSkKTPlPRBjnB4Rt2Dm2nUwYd
ckd0KoNehd6eb6h5pi+bFCBWOK0SLQBFKeG78wzp6iNtARRs/mgZRJAdvlCMxuJc
1YpxIuHLP9IYLR9eTo/WdmIyEuZZE00GOzWoFV2VvPi/hbNsB7H7aWFHZgqUREij
ZQ5wVV8AbIgvpKAr2doNIwFmdJMByPTGBN11VrdYhS94zqSCxiGoDdh2T2ks+L00
Eq6nxVQOJcdTfKA3qakbbDDrvYCsOz/4EM1BEsUvdFw/RSWip0NDa4LqsfxeUfRu
ZqLgWcleXcwbh3C560Xu/0stv5FFrdMwTpPvP48KQ846sKEzhyxxpO9aK/syMWNe
yYY0UqD8IuSDups/Kfbdjm1xbL0BmzwSbOzMi4yRDtdr7EcS1+EtS/V1/U6skn/D
qBhsx12icKNFlnuLwXwPqtExPr/KEVc8J24LUuBJOKzZpa7VIwc2rqsrMffAD3HH
5NRuURCTJTxSkipftJOjMXC6tKSKE3iuuj8NQ4csvG2+B2qHMZPjADWSjQbw6hog
LQLsKC+gcOW8qzan1nkICl/uN1nd3EoaBfjFFkOhrp4OREOylucTUBqM6WpkAHUv
y7qnM600RnG9irlPuQOaFZiznXZ2jxzMgeUsY+b0zyEpX412UOGhrg4hNUeCbIcN
p9uPVC73xtMg+NRYOkH/QUf5Cjkl6rw4jfNwN0T/QVnfgVvdgzHlzdgdaArE+CnN
xJhdRENjYkyqRnfch2Q//Tx0Uzfn/BHTms1kMiGSSyw0xszbWpWGe9xz8t2NKeiV
mLR/GiHnL9NzM22gW8lDvvma7NvHhQSmmxlaLR0OojuPMeJu0638QNra4xGiGTzL
Fp1bRgEHn07ssWW5RFapnf+jTsxg0WVWdxmVg7eQgpf9Hqm+MwIpIvoM7EOLQw3C
i8+VkHuCsSqQsUyueOCbk8QzBie/2XJ7KswQX6tK3VFJcmFExhmGYTLdC8lGa57w
Yi2YFpnjRU2lFzguvFLkZcdDc0dUqkJbKMSh5cZy5yUOGe3bUb5m0ACu1isqkE0p
eCJJynrJQbqC2S1MegLbodrHRGpm+CTkSV5zqU6NEvrT5UlymRhg2JPipxnDhG/N
lTe4cXcRCKhkAP3UvcKup3K3f6vbjW5OH16NFwx4Fj9q42+dcqMx8EFYICE7E/5v
/IhC1V6S+0wdFFUz4izlGVArSg4AyftlPQZfS2taqdERo/OWkwmbo4PDPnWaAacg
LXhUvDSiHfFn2ptXuo1kikvN8864xiRLIwKCoNxiS2UXcZ0A0gIaL7wg2oYb/uE9
44QHMxRPzdaEGAYfViwnJwxeAuAxG9eZ1ZLltXWhJZ4RlvRMPiLmT4TA1OLFKabB
ZL9BiMFStfUcEsC1MECIZ+gFoAuVDImgb6EztBaLSsw5PHIl5rQOA6kDeoAIPt3E
2cQWF56VtjC24wDDpXme8/b+22g8KsFQk1dH7pHgBazRB9Im0t9RBPhptIiw0jSN
9N+FavynHA3yFpkfHMrXvUDSgTp3U+3JGDLR7NLuhXg9bIkfX5ermtOPRc9Vj+Kx
MK3TmUWI19GQ4nzQKqZLsdVRBT0wL5wOYn8FaRjYIK8uUWYURyu/lLip5WPAgtyC
TyI6y7zsKHWodmRpIGUb2EC1FRgrp/5ZCGaYIspWM2gLTRkOVDUeBJ06yJOYNgn+
TtQfs92wWVcY/v9t3d1E9+G9edGT2Llrtnknu11yvZlUL3D1TX1XuVp4OnCpiP1j
WSkSWVujtgcQjqsJY0+5CNu8tXjwCsXYyBZ21baBvy16kBYqjmUOKI+EsnwDGtic
F1726KGZj4S6c2QS5/WBUPkPYugAkGQ7WIp1bOuWP+61Y+BG0KRzSGgfDDlL/lM7
euJhJW0ukldH6zALljUdV+7uZbSqvTll+ZlT6XFLM/mthG1KlDBZDGaT25i5swdM
YhnDGRxOU+DC7Mp6JIFumqRKK3Ab6P5HVywF7nSZRMrtNc9cvdc73B2Zloqy69DP
1fDh1QZGMzCyPdg/Pd3ImckPg4pxNUKm3oXk+HpNmDaYGTzO+WS3nyuXoisHJW0J
6JdKR7/hN6M9y0dgMgHUy58c2233Bn8x7Dg1gmKFgoSB/1waKPoMWN016sMVLf6j
0DQvDpL9mKyJyiv3NdwOE1DiPPC6RWfgMpv7B1A2cMrf3N1CkPB2K9/ihoTWiXCL
PKp1p2R8v9ns5ICI1ALSE+apdp+vCt9RFOtwjfzKlvuTwlPgzF5cy0ehWUcuKcBu
VfFLigAc8pqDuzotunbDEW+3awMEPepZ+10sL9KqCK7cAmn3fPjNowkQRK+eRN4U
4voPtQIC0CsTkvaHQ/bzLUEdzxS7zntnrKAnpCDrmgL2fpYizuFoP3+W3/demDDj
BZTw/QuU9VnfkJ99kI06DVytsbPZdfOA+dXy7d5BomXcPViui64THK89JhlBM9vZ
bXyCGNmsuL6xNxSKEX8PML7W4Qvr62aNe6Y97RAWkYy+6MwsDrxi6sGidD6dMb6M
w5hismv0nwZadeegoo1i5d8modXUECDDwJkD8+pIsoZUSfsW2fAhoh2NO0J7Xpuh
oa6boeX9E7ZCtkWlJyM0cUHVn5ZaU9uNbpmZ3yI+0PufFl6onDTLV9VoJAQOmshn
NJG4lHPUehVJy7MVEYZFB2CyC+X6jHCwUO/UHI0dEfDeAduI3GZT8nif1A6bklnn
i3gSXxLW7fGxJHTtVGwRA8sCv/bgVaarI2jHnxt0lmdztYK6W+AVKm6TuuFNZpc4
ywKh8yVA6qSbY8LkO1N02LBbgDfwNbZNvHsm9UpfAusi+SBaRe5NAmcpFeVdFzks
/efVbvVgP/6pJRx3wdR+J0u38xnR0ubOK34MsiUJmr5hbxHvhGL6FkF03iPRxcLX
FjhYHXxUN42lCZ3LAMP5L2HUzBBxP6atMJPa4i5pp4VJqb2AqM5VIWXYtIFZZLQw
QiI4v7dbL1rbWRdX5+j0G/HFiACl8qhd9aO+Mj/Rsa3bnfVYB8BGXg6eA8J0G0Qu
Qqy1jIQFaYxcXEYEZezloyVc4gKAwAvd2OHxOopg5U0IRDaXvJIhEsTpRL9ZrBwE
QbgQHugcFGWrK6cRH2bpdEPP9OMr3OCnV3T4Dx8iQcPa7O/SO1SuHsajbR8povuK
RJhFrjTKIe6olWJEcvi0XUgN9h7+jhoCzFCXr+WDxTCq4p17oEMXKsXZShNvvQIP
b4NGBPKQBbxuHy3DKregYH+hJqtpALLmJ/LepIlYcmIUBa98D9rEoH1AUh/FNcAD
85G/VgovxRwrxXp4fnNdw9uUsuxsg90dXpFiEF5qzW68V8Zu50hRjYlEQyv2wDzP
9WX7XxQw/0QdWCn2LKJNVGXzzsThMHx81k9Y+Jn05Go05BV0stPY6vSL9DVITL8c
cidiBwmOmgaO61Y//zHXMu4k484/h23cGRp+zhI9EYjGxo2DZFTIY32Xiovxd7kp
t01Hw2GNa35AEaHWSWQVbIHtpqbWPIAeTJiLluJSljmajQKqlWZYdRL23Z0FjgNc
xi3uX4j72RPD6Htfqb1pMol5Duh2PxN5dDSXcRPOx6siIdqZtO+rd6RUF3iKgufy
cPr8xB9NLXl+2iL52LbwjhZx9lw4rTft+qi612ebjc6UW9yFfcCYKkOaic1a2/1s
k0pisTjoeWX3eBGeAMUocK6FYv8dHUuTAR5Bah0X00Dt/yMV1B1Lw5GCBak9/93F
o14m/sucu1I9eVa5rPags+/Krdu2GZvXI2aUk6dSJVb7FmUN4FPvg7gXXGWJicpk
rtGaWMZgKzx3756jiZ+aEsSrCE4ftBUMHdB4iV86Uaa1Fp1r/nzl6PgfiLf1yOhL
yFptjw9gB1C7vtOVrI9+zx2Xm9eOJbLtrmRBivWTYYDtGvmBKa9namgY4lQl7lxz
7oIvXZAEMpCQQSnzszvQFQMZ2KRaH+I+oMCMgf8UOUbKR1HEWB75JmJqEVoGND5h
tIH45bmgtk/vOdOs9mB+3OuhBe6a7FpT5yyz+u3bMkkDcFbL9QtySyQBKUT+9ijU
3AfGmAfy5RsCrBMwV3I5QIYEd5swJ0NIkLNjmmOJ6gFgPdwcEJRTK/h3W7y//Wmh
zC/7H6OZnLn9Q6sY3sHO+o+f46TcQKtyTna+0pwC4Vuoeh6VsYUlhWVu5G/F5lRK
R/yK3SliXaYPND7ipkzxNbfOHlsPDLaSIS+ebZtd+GZh0OdaTORnNhH+6rv77CoU
DykfjBQCfVbhUEk3j4mG+d7aLo2iW9XhNDW/4zNSi2rgNB78bif59544+6KFx9WL
75LufAjCGcbT8ZB/wZKYM1yip4mJgebuySMcdy/rM6ALd5X6Vz3HA6QaELdys7nc
9vjMiGGcRFtG7WmPK4BbplD0DOWNa0uLAK3njG/oHNDYBnQXp0mcZY2ctDJ3AaJ0
SNxLFP9CmxFbaP+f0EW/PWEiC8lD30VbWyAjlRlepCd4ccZ3ElZ8uvAw99KOQ2S9
FTEMLSXrY3Gi5x5VYYDa8+YUWqTKvVALuoNDQoUBz4yt9jNJGBcAw8AZDafIUdOd
ptv9l4Ya3v3d0LR34/RK69IDTN5lsR5EczNjFSngxAam5eJ4xrg3VptDrRCrcDJ9
pPKXZ2/4kIflc2uJRoqkEO4R5yCB9o4pUAqcfY9rr0tBXX6wc0TQEcYrot/FmYaz
8iJkunOo+c0/psFjrXfqXIDJTBTiNC8TZ5eGXqJ8deRQQLV25RL0JRbsZObdgwYM
Z+24OCsjGv09PmcWK1YbH1UkgR4dLhNdNIKZ6kiPVHqIGRH4YNjJWvaZVAshcOX2
W3fzNLs3aLyEgV5IU4l2utyQQBLr/i9qhkEs1gYz3kGZJ8Ssa6CO2qOg/fWZnXg0
44d1BNY5yIwZH95wu0zN4/MTrUXJds90uAnF0RxUdxQtIbkVFuz1VbM8/uPkDJN+
v9zOomthF8e7kn93XXT/VGiIXrKbrqEbd6LM5y5IDiKGEJnIIq3w1MGsaV2o9AQV
9rAaQepQGBjyxUsdQfbPt5PFFrbTzgAiOFTJqMDSTVCf16uf2sBXMcmx6nwaN6+m
WFtSc/orUDcvBZdK7FP5GXuEXBNMSwarxYONZgrC8mRuabYi3Lwu677IQJtayhpS
P+vgQ23rZw2h5uoxrw+Pf2DUwplnOtp7gHuPw2sbxO8l9R6KMJpDGi07wUwUJnuA
ZGGfxriOEUKDLkw6GJNqTC5lwukCTSehqkmg9STUW5hhqe7LaqobO2y+rrtp7D5h
ZIs0N+q4DoTQCHP3wmEXLLziZYVdrrrV8pDTf64QHxk8NOA4Zp6haRlhJmL7DxOu
WC+r13+Q5xi6kUMfdgtGWIsNg+4UFBeGx7GWo9o+I3bbuVOclGoRoKL99f76Kksj
GWVNHUs2CRRQLCAk/lssc+YxCBUAcKVuRYhaXxrHpTcc4Y41g/kzWdVtYF4Zhx1U
IpwQcyBxDnNrRP0ygAMt4G/14TX2DX9OFjItECd8JC7yLiX7IZz+QEsRzyKNL0Eb
ISS4pfthGcfaU5sIlPB+vE3V0fAdfAsboD2PGbnmYfrIoAyclWSjcWiERxh2Bp6A
Xgpexypr6J6yrriDsSy0g48Ik6aVmiX1AUqg5Jxm92kw7Y4wVWKThOqZSmTmYFgG
L0kUHV7oWPV4p/uThqI1gAt19FV/gRtNuFs03W018J9hJIiAHW/TJDchioTjOMTu
2eL12LsBPGEGsfombS18laxMkmYsYOEryqzNfikg2HtTV8wpgri3ZYqYVIukIvzw
wISiSvN5b5HlCz/jKxQ3mpyKtDhvDYbpbkw3pmSKqNkLzhtgLeeFlEl/8bok2vHk
KKw3WOY7x8Zn3Rp580uUalo3mfku3PIpCqTiUh1iIJ3IiCxRECxy+jrEDgBrNzMB
KdVjGjqvwZEIZ7o+GfAhxM7zqTJryK+Jk6lIpbZS9NNlLtMtNSwGLP5XgbVHRhXZ
H/y0Vx9BKA+TN0qr16JquqmMq9Yd+GP5fCdVNEiQf6VjW9THedhm82ERpKf2qHsZ
2AY4KLWBWCGg1EB0y8JlHEMlzPJs2TOxc3Bgnu81uqtRwNVlLcUeVZYvalmVB7Fx
bgRJvE2MCtzLvfOYJcw8toNZCBQTkKQ32VJDI9+UTgoZmnXSf9xOBB1as2VZ2cKD
LdXF7texOdQ2duckh7LvivpW7EElE8opCnoBuvrXLztzYQgG5rpT1wFRQMxCKq0u
UmE9zmN5fWwiT4n+oaYS37YopFPYNTl3xCS7CryC72iPxHcnDtn5SWJXmZCrR4AH
T3jxYUFMy71G2OqcUtwvaQUIIpPZ822NQ0+97/CCGbwlbdvy4JYkuJt+G9F3oWtT
V3FKWJpII/FJAcv+qF6wQnL5Rp08C1StZzqJWflAexw52NRij9pkcH3PA/j51leL
iLd4J1yoafQOWLxWUMeCb2WMTpli2Bi2RQb0xq5hC8s7od8wUJrcK2gzpzcZuErX
MOEJTJ8oIQf6tqbIfOAintQMSIY+ULai6q8OW2g2itmpmxa0kGe8robQf/CW2jHf
WO1U1Th+tzUKq6+dv7yi3EXHoeT9xMvznOa1XHYdmFGyAhuZib2cET+mKYFCaumH
VoFbDFY2iTm90qyYQDepk4mkThSjl6ZXGBK3SbGKwaSCh/oyaqlpW9VSAzyxrwH7
lUcfYlR46xsEago8OmHpSkaOG6cj1sRI1ij6V8Mh7B/cG21ie+dYhcyboWY3hbkW
PMOGaSslKGr8iRx0nctBHQXtnvAzBO0tUaPbW6SJyVtDSzdLhUlERX+e5UKJJg5b
l8BQTOMgpidBvWBxVbgwkAodkQ/eYipnID3zkxnMxH4CJg4E5pjW9Dl5CyG9gK/G
T0Yw81UtAK0wJi/bNzdwfIi6HF5Ah1NcpV8a0Hp3B3ZEXLXG6R/sYakWmCJjMIFD
+20tGcHFSxuGpX1k56k3Qfgco9o+Uap/JjP72vFzcmHS9exo41OR9srkdZUBi17G
R04LHdWs1UGnDgCvX0dHOcsW/xo8V9yZXOpD0mDg4nTJ44uv//Cxbkz6nvqwnsei
oqYtO8DB+ywPp3B8YUqlJKSDg2MK5hBC7cEeZodbGl7LNAIcz4rT3ybnx2yfEjkC
aBJ3sHQN1fo+fhhKlQkedEUayU+gN9UOfcICYMKNlQLIGR9PKRLVLsia+jX2OREo
2IKWPM5XJ1N0/kNdoAK5qMmWSCQAjg5KT7uo7BJCcbSLwMD8djm/Rs0THIXZlMGQ
NSfocDruaDJd83GzACtZFpOqrjrsNHzkV1Ej7jDpygTxOBsYCOuQP2VRDgU9q282
feSbrlquYlcwzZX3JECI4qsSOuGZgCdlddP11G48mmHRuJYep92AhRYOwXgpB9Gf
+0I8Ky8gqqeeW9cFyKadb9xcdwZqUkRtRjwoPlyFHjiJJJGI1ABkayL5w83NXfpm
aZSLBBQDI7lktu3cotq6yQI1RBc6qeNNSPP7OYcDzNeTkIGgbd1TsiD6/tRGB0zF
dug0aLc1iz7MhSpC61/w2tC4afekrMlAMnAJtsmHUzfUmdw9qPvht+1xRgSCIK4l
3T4Opl+gmmTuwdzxO+aZdpH5vYKsqYkbnliowAGiSUs7eS3Ww7wCN0lEBLY67N9c
8xAN+2HaQXRp/7rubJ/6p2DVUttK4PRv2Mh3r4veqmGkWX5PxkZZ3bxNM0pBraSm
8nfJ8W8zyOtTRBCSFJu6XiR2vxNj6JtiqtOBbuPxxAA3yX02OkfuJP9yBDjBj4Ue
rPTHI1Q9PM3LSUT/oi18W14IlkLP7fN5qiJe61i/r92lX4TyVdsW4MxCj8dH7RcX
oSje9bTeWZpYxsxz4k+3kKHhWoctjL5wnFwtyojzEEAN6p1VfTqyfGaR0NcMPttK
h73dL7KdQRjO/GdUyH33vmrRuaMLc5sQSMNnPQFJB1535iUO8Qo7sCySKUKFI0YH
cbLg23pl2G791xmMhJsvgTTbh+fXNtb9wGWtzuP4grKKC9dBTmckwJ7GZPQ0U2Qz
cZvJTQWUHf8zRG/X6In4gDIqjeUA8heaQKnyG7q6nzY8V6rleeOje9KF1X41IfrW
+LXtDRMUpJZs3UDxnpOrCAtfmz4EPwyVxH2PVitfHHt3HTr5nY6iHAyLi8HmbR0y
QulOMec6fZMCM/PZ5Vw938upymHMJ2DmhoNkA81KWLUqFBIJTLG62XNK1qNNyYRA
eVt3t5GcUZ4uYGREuDqtRIUPYUreOzXZpw9F1p4yv7O5AVXB9+lj/hNVqUJYKMHE
MIf5tUeR7O51F5XsPQ38TmWqMQpWP5EnGo2riHOpCsy1rEMeXVGlhqutBGwEfCJi
LH/4Ej0QIyVM4gJNkwbdDyvfnSRhpbl5uo0rjgvarUMoFFWWw9aw7MQfb3q9ApWq
XLPdzhKoFWS9Rdyx2mQpPU1O8PdDPLP5u2H8L4OG/w8NV5q+zfqLNuXaRj/kJl5Q
a9zkOSIU0kqS031s5V1N0Ud+K/H9Jm7dmjEpaoEPqQtt6mPPsIrc8vCKyP8Tz4Au
s4F0XU4o8UrL4OL2B594AvDZTtzbXKgXXbJtg7M9oIXSA1Kil6TjmIyLR6TpW74e
JyjhIq9MdIxK1iDPP77NgPbUiUysZPo+h75mMaEfAhG0+Jh+kF2wIqBWKDidWZMa
CDxbRBZIexu1xX7CThTlF61gGdnmSR0ysfoYQybh2+MjJbJ65DSB4N/7f+O12S+C
Jcf2Q0N6MI3sSR2qMR9dLpGg1Fs8T7o6ZQEW2Rz205VyIdbWSbArRjFUsyJPhXWz
bYhPa5w41MSlUZBLxjyzas2Vx6Kodvq52zt2Q1F2xvpXgmv4jvnTNtAhpvpYhslS
ZaNTH+HEx6MU186ZDg+BWRQRxPqSGF4M8vJcWu3bf3dvWX8qBqncU21Z4nuKm+fM
wnzGk1+oSxsPOUsVqMPAxbYWqvIT//Vl2ZJxXf/yc0ACEdh7XiQ29YjAjWH1+LFW
B5smjhu3m2b0SrYcBwAKjiM8ImIb6iK7OGKY7aHgldDMoO+uX6naNyIbsDizAUAi
hr91UMufaAVsj5pccEOS/rffcsCjMu8FEExunUd3WMPKPVX0DlAO7uoSQ80XM8/g
iW7dz7S4iQ/O/CiRJcXjgovpGvVohuCrtM72CKGtdBcAbYgu//C8G/G5izkVMBdQ
WPCzSGMTWF5Tsj4O+xtyYs3Mj8aQItqJ7UhK1Ozs2ao9YRHPPfc5Awr49/a4KV04
zg+HMh4oY7SgcxOeJ22hTaI7PRJA2RNHQtmi9CRT6XhDl/x0NjsBfqQ/UBNjttmr
P7YR8z/lNjotLu/zKvAU0DOiTthjnmGXbXYfP0/oH8+0BC+MXBz/3r7dJNn2HBSi
4tLGEntY4Qz8KZ+1xEjVLPSBABDdpi5+zT9iuUsnME6UJNxgK7FDGWZrRzwkQcqD
yRhl/kV8zYkLCKAh9RfE0D36yCapHhZ9gMnYWYSk9iaXNFAxzFhcpew2DzPW/0iW
U8qe5MpDue/StBQrUMLFsPY50Dy03bSiKOzkSfWhkxrv6F0QVC8ZnCC8+xFpoWrN
yTo2z4D/dEfhZW16GJyzFeHA3uHBh8pgh8IBcdehBVeKpo5ugbdtCdnJoVtNJUD1
tmu5/WqRqL89LXLHK1mqukLNQ7oem0Gylb/KWIT+kFGHGILs/fqa5Bbei/WHuk+d
vgjUAntirHBAC6uGboSiL35cVlrV2v32kspfqiIo0uWs4UihEtVnVqekBD2NCE0g
zfX54KGh3q/VK5l09IS56tYI/nZqYd9NA3dHzyBIofl0jaUwmIIQjJz22kmyRkWs
NU9t9tTNPhFzkJ9dxcutaZODNJFSWG3+nEx+Jk4sn3ymbS3LWfnSxNu2SEj3p/16
hyjjq6ymruzSHAHRRtMiLTnzdr5aSpNjZO7oAc1nV2YGtTVE4rB7bXLyG7xetzI6
xg3DbAuq+ylFUa2uYOyVApyyxDQbWBoK1m1xe4ci7SqRdMiHcZONC0TSzDJvmVvF
dVZD5WVOQB7inVLLdojyXI/GXpPi/UW8BLH9L2X/DIO7w3q//5RchVN68Jt43YYU
51gn2rFl+3rBUMpnyAufamkebeCkiC5eoHnol3hyXHU/qYgckDz1ujd29gKCXE2x
M5OcsZdvLCdwu/Fewsu5Xq9N1Oh5QvBxGbgr7X1niVFB2PosXN7PE7j29oaapPir
gUUBEv4v4JWHn4v1jldJmXuKWFVigrsyZx5x39RMbNad9r4BV1K5qxVD3iIlvtJ+
a6KQJ6X8g5xCfC9LhSNeG7YRU5WQUAYU8Se5bE69H4GiedfIVkHT74ne5i6XOj/X
N4S4TSXYjeHxReYY6/wxhOXGJyBv2Kh/BpOXF3fhvob3tz5fV4RbxlUud1whmxPV
a9RhdJuBdGr65I+AiqFdvtkO+COVMRkK/L/WDCld0BH/JSBwZLz830AS3r1XIpED
DzsiJg6ZHJPfVVOFxNc2Xe+qhghjNNOI6b9/2dt2NeRIhDkmhlzoQvZut1DMz4nX
+BPjGRUiUlWblNW2c60BdiBi+U8gVyHMoZY1l6U826bXUina7yFw2C+S1kEOCVMQ
909K+sw4VZHoGaowLrQZLtA4rvBYp/zMtaFxCrS5hoCyZRqcxNeI9bAHGiYqxMBA
LfQKr/aaQG7WYYqh7P7HX9YqhyufCa2ZlcXrtHRFWt7teJRHOu6I3tNaT3dm159h
kMv/GGNNdSGya1gJKR0kljH3i7By/GOIo6ywZZfijspGYYBTmkFCCAvd3lgq+wIG
pPja1Q5x/fWfvCSjq8y3gfM66W0VM3BQ1OX0nvJbYj37CaRQzjRUKgz0KRwbxcOI
4Qt/VvpQgZKdi6c1KImiLMu48iTBSzpftAeP8MB9qq1+82HlBhX2LV0CVYWde2Do
y6Ec1U3MVof6OeIDP59gekmOQ7mLSgBYfM+ttVXVA2Eey2J2CWdZlqhNa6WlPh5D
2CIYP8TqlxTmPsv6LBsgBAR0IVDGVN0EoCMWdELvtjDMOM/at838kQC2a+b30L18
KzCo9uQWIb/pu0+YFIRv2XtRoInohaWJ4KTSTNk16BvUwEQWUe277SQW8A5CJDPs
2BEBquWjSS2jcAjlZTlQHDBS9rWwUJIeMHcCiy8BIjoZOkwKhTM+m5X/iJ6ly5/r
4uYf2fG0Sely6EFN0YmNgHlFGB3qCwPESivX/oS3dhXesU6/3LN6soSGHgg7O24/
yPSdDBiyEQelwdOtdgImkgBOb3LwmsaqIQxjzExavcsCVBayuIVWCm8sKelAq/qN
uFAjZHQtRse0zFNEOG3HeRxDnuMAf7NCA4v5fzlplSbJXq8uRRcdVQqI5/jLYx3+
yo9WFy/oKgRIlzaw/lXLjbZ635pGXf7AXtEaDge3flZVMSfzUrErq6yyA/l9E9Zb
6qT4Y6HgMqW7oOdfh3AuXz9F02SN/q7AaE6slayr/6fySHarwFhXQm/cHPGbfWfB
8fbuj3QMWlXCqoFPvHP/accb9DNjX+T/aM3+S+P388KGOmtzgSYlyOhwNBgY97ks
qslP21ckEjYAaQkJTZKqVkbm8tGlfInMsZXO9Ex9AHZ+oRsoUtRXXO6xjeWkiN4/
R+LxfVDePFzeI3qDWlIq23yqG7WGRbBqszqRNbDTBAYOXoHxA8tr8h4IDlWk86rn
nIMEIN24lT8+FwMRBqQC8TlG5GHhi1nAbsJH6BNfBglnGMJKaaC0K2d5nvQzGqYI
lYb97oXMYkt4YCD1uQ0zKlHcIuDHSOdKAaz96wpm2xmGF8XKlwAd2ue/JEjiWFh3
rpVqup4vCia4sslAWmLCZAOtNKpo8INOqnayJNJcy1BTvuz1qY9F3cvU9RqPSWeA
XZdMnyJmJkbA22TxOX6NLvUywkZA53qpGxmQ3gQPYkvmhtu9WePIIYhJcERVsvqZ
INDEjdwJ0dbgWZ+JoueAmz/aB2FiToe0a6MnSedBhUKdWkOdtm+1fvtOOG7bMQdE
VFgZyS+8RPo3+t6n4ezMVg+SZfyu2DVGnDnuvRvkGtXwZC5xCQXn+VE10vvGcmN9
Qj8UDb8VJ7bfx98h0Udvti7d9he6fhZrQSAUp54kyQai8t9T0IVeNWWcQnGfSRK0
JMS6537iSF3cy75ieZjDnlkrPTrZI2sNSwrnVnyGmOOhu6wet/vT9uCqvBswWdln
p+3Z+7jkQvMuROeoK0MHPO9xfkMa40ytMEnjhUEwgzjFV2s1ZEKfKU2x/Lp9/KeM
AELeEqBJ1l8O40P9tql9gmff//PVcwCbFLfcvLealy9/+iMrVUVXjCoDmIGYRC5T
/fWRtRN6NaUGsln67bhZJxytskd5FLjVXyO3HobTyIejBJKXrxkOzskTztDJ3BIH
w945Cx6ao/w6cRo/WYW4qiQY3XV15xF09kY/5YkBYuqzP3ysvM5NaqtHWvjvyRvd
w+x7v1pJep9Tg1PiWDRf7I+zd6n64K8uM/bjdguCmmK7Jm7EwmkPi8VrNC2rdUqO
GXCOtwcxAmkZoGoi1MsAtZr2fijKb07ZlB7qXk95PMgjRml2CC7zzvw7mvnC8UDs
U5YEq0RL6ucYT8rCrVf18+KCweOYWUrnzeaR/FGeJE4foSRRUxG9MhFoBsfa6W/K
B7Zv0wgO8nh+5E5hBPxsPHW6RQi3znJQzKbIDXRpmEg5qaF9nLrkmFAijHxAckHo
4wbRu3bS5jTfquyCUPSvB6dRaoukJmUNX3bEoIXJNFUHBdLAVNEsDSSrQtwMw6Zp
3KKKkTp6VWn04V0HcYfaIG3Or7qQXutYLo1APrAaWsajThMou8OeQ5pTn6siMl2y
FXG6MDRPQYvlIiHIlREV4MH2wRZWrJubFYUGzMa4Jrk4pfflEO1S4Ug3KTJiKwqu
eu4Z4jtiRoLyeCNBD2VL4vRohrXxCmxtK79P8SamCR+RedrXTdOiRZxBPtYujOss
6hU2N2aNMXHCTE6Zw/Ypv217nwBUmpYTxv05xl21h18iGvpOKWwZnobFW8pTHLum
zOqaAjJ+eR3Wn9LRrF35k/FnbdcZC5ozR8lNMp7wI1YLx8LfJSpOmKCg8txhMs3f
gMznVVIKidxXqIc8gcUqp8XaC5uGYKbQmTk2mWwuKBsODexnzGCgP4ZBebvB5lHp
C76UXxfnHEUJJAzgcABejCUG0Tv8SGqIGog/MMnXQYRGbLX+5sKjRcXYXbAxFzxK
HpKuVrxHaTneKnPl3AMGhZZNA7t/ZKExdsM8wTiFgRKxL4dgSi5ZlZYCT5YsMu9B
jnEIgDkcXZ56ionvWUsLbcVowYXphUm+gtU4K5YeL6nYKHt6R1cfBqUiwKAUD509
/cukaJPyiFccJ4D6qFHUEeS+rA0lPsPaoirywOXR4BfWLyMLIQogywVCWGaH7EWM
librchpLj90QwiNsiUWFBw3aP+PantQS8rLBuExeJNp7OpMCeGFMHmOqYp2uIhW7
P0mLFp0gzC7z4n7ZR/Y4gq7p4+Z4aNrzQdMP6eRVyIgiugoezemHd+GRvXE5KqQz
rk5hP105puiFJUGsGAOJD9Ib2y4W9YusboHSm9tD1llmLtwV/BQueBg1lr9l5cYq
GjrffGrdRfwbHaCGy0Up+FmH1MCgn6570WmbzZzsxO/bjnOUHmKu2rvxhnGSKnQc
/lQzIiScDuU67gVoTupkCqsx1pcdHslK9zA8sTR9WbsqhQElJI4ZDiCVzNEvQp8K
UT6Cpr7wOvmW3NtwmiQ1set3qiVYOet8bYdyQPe977/P/HnC39rWIyrhEa/8TJc8
sQ/XbObNKXWJEW3iqqgPt8FcHlS7+4jWTLk2/LJSjEEgIdSWAGvwUBj6GEp9Sw5E
t6gnoJuLPm1N0/ka8yA9Z88lc1jvLPd3TUPsKu71fHwvsiR7vW7gt8hNPW9EXA/Z
P6JT0sjcfv79fAWlvE8TSPR3ajvXHnEavP4tId1QGY3MzL7qMWFyLM2S6GmE5M7P
HcgHYuGSEOJ+YVqWBLiuXcURkRKSsF6VcceUvDxryR1hri0pz5zt4AEkHshSxerg
50GtLznQLEkGuMgG6vXirMrilOHg+SbhIFyn60opk2bh/lseLVEFGBjG0vHbIjwX
tRwEgaz6Uh0u9jD9mRDWARTb3k2Ve4NxuGORAL3DJedgHo7NUMkbWT7MtwFCFz6w
WvfQb5lKXDjlv3KJlrPyGyV41iHBK+djbsZhlNLDOpDrkeA7dlAw3WrWLQeeDA6V
H0nxQDvpcoVhnn23B4TrnR6N0qryMOeYtYeNuFAmD6TnP353WkuWRkoZVt1Bmr8N
XTXWwDC47FS1bvCFfkH7KxFDLoZoJHm16DDQL/Dkw8CDHml+BJUJ5r14LHrxwGD3
X3n/5CCl0HiINquw2etz+fsQDxKYU0WkQc86//ieSHYiJlDA7w1Oh1UFqMnuImbW
8p+np47FNllz8NcsNvHqocZwz0HR7qZ7WEy3sk/txbwHjMf6arYYZb9JZbdYMAgy
yw7Z11W29vLjIZXcA9GjkUjG09+1GjaPvHwwFV0xmlZH8Iox6MecRzqldjGL2b2p
zBYRtfnTVhi1DJHsrzL/WdDOD9mVhvEAuU0lRbVA2eXFPzQRCOcZSx0NQg4ZQnNi
pRYKl72DbypoHQ5GuTlJ8+IkGJQ09/UPa/fUh8+S8joqnX1y5tI8DDh2vQkSlg2E
slyZc5gqlflbThEBAD7epiZFmkOO57eA06t6O+hpS6ddElcLQJYf/ilnS7Gp29q6
prSnUy1oC4BOulD1xtbwESpG86Pz4arzm8mx77ldpSjfgko3+2zPoOg9rq8UUhLD
e+e1X3LasjxegbSUqZ1L8IIsEdAzIAmBj79t17+Hn5DMvXQFciSrBYC/A7VkPXI2
AcoHYWxg7wXpT0rX47E6RdtJlfJQQqS1vg36Ajc+rYGoCndB8xQqQ6CC8ziBiwZJ
CsiLxJk6ZRqxkK0rLdRiEnFFHNG3dqfZNm6NwfFy/UKVUZc6ezsxxZ5/ch6d7gyn
G8TBMZ0SR7uUo7g07617Upcwayb9IGlGe8t2Mf6lpSNv2sgZ3Z/D9SkWvTJ8SuEG
bf3OrShR5hGE32b6uFa6gOzbDRrcVVBagrvV+Ag6dsoB2tEIMFzZvWqFJtktSd+W
4Gw0d6lHjf9NNs1o6oXxKi6seXFp9B8EXwKO4KOx+HEUMkOv60su08PmyYfPMDgf
m+LSMkeRvb/t4RVRiyz5TcAYRz4iWT88W3nzu/UWvI5wl5kswbussbdQDq9aUuW9
IbrmLoBTK8IWUjPLL35E9aiGG4h2s2RX26tVVsf5MzXcfdFX4lCoaoIA3jyvy9IW
2rNEmIC8BiW8mK9CTHoCO7xqKXbBE6btcWTDdDmB39hSA4OGCFiwSrCYs5mQ//Oo
RC+/qJg6UviuX9RjaWN4LXIMmT6zTBGU3knOp0z9l89FXKnmZutTDGu9A9hlOvnu
jQl7uNEEHG7FgTmhAzkeWwIQBi2hx8hYjDKmryIAwAe52McqrwmB/7dVdHdSS9Pa
bXVwuDQi5ReFxDnD6GPluTG8KgB15mRT1qbTX5SiuBdkCSn2/QbmdfzS0aOpUUIe
IG3u3codvVfL6jRA0lquv7d3wPcZ68MlYKho2Tt6JASxQibbzwS0MUigNgzdE1kz
CSwQKReBhtkzQNmDsx1hReT+HC3b025GhNS/+oJzlMuiFusffAZwIHXluHgZAFMh
xTKjSmYcB7VeUrLqgJ0UHguG7xEiwi4PXdCX2Fo/++icPV3zoLTSxxylUvXhsa/1
49AFMxpj1RlTkjkUpEe4rSJBGCD/s+8YU6NpGQ9lqmlifpaYxQNKZVYnsoScq+c4
A+spPQCLYvx1MCJS4J+YDobw+Ar72WgaarATs6R/CsEOWroICmEiTVZrAj4CNh2n
bTNgatz8iJhCF3fp98a2Q6X1ZNfFo8hzNUe/MLjf9F6Wreyuxkxasss61il60ta0
O9Qqo9WP8d0Fr8/wPPKUY7aY7JSjddBI+RvKNzDIB9rNJ9m8Y0ARIA2BrtZ768RT
doS3Kxu7QdIvjM054Rb1YnKNkALVJzBNqlVZE8R79boJQTmETtMjXtZbwke39H2t
r120HHDElnRkKtXXNM6tq2E2g/bYu1Epl/3GSs/BEpqHd7pnQUAfFY41M5pLpjyS
8lS4OpPvnwhPSKB/2kN+38uOJm5eidYspSt1+/NTaYuJOAmeuf1D750oTCuLsalC
L1NFhc8irXpXGOj6oH06y7K65iyt4mGFBjHThPHI4YQBDyKCDKCZJwsR3n4TENGR
YolA3vh/KsvaFAnIegbOAC5jHuQfG6VMPUr9TzVmpYgjThAQsuHSV/wAxN+38b+q
S/ks8PfKtL70cmV1UqpAgWM5w9pAk6MJ6GgAshqBS8yw8YCRzvnbzp67DJE/3gS7
moBEqVRQGfZaGOShdiOOjraSUdXcKTuEzXjOhXbKqT68Nx8AGdeFaSZLGpj7pnJ8
jjTk2LkwmYyfkfr+Vo1czW7cr8vqsKCaxAA2ls75zPNKAMHmdt1aQ62XT0DbCQXN
F+0RQ+xkaepHqzcl9CkTwvdvQ1V7VSN2eBSwle4RC2abTgCs5/w6ku1zizShFUcT
gYSmGns4///KXxkO/7ZVG7vWeC4SMmhFXl2nq0CKHWQjNKl7nSa1sjqOAJ9hR0Un
ukSxsP9dFwtaTaulO2wSZypY6lgJGzdSMLlZzghG6aOIwTztnEIQrH5F7Z8WPyyv
1diMkCU4VQBda+l8F0EWeyU+jz55+9BZQ+5bKcIBlGp5yqFs8QOffSiON/rCMNi4
SNTW6wAlKODWtgljVp4J0kAiGNNI1zbQDTCkSBxvAukkX08BNqPMKxXqA4h31wzh
HfQXWi5Lzst40vgPNzQ0aSQUmcTyq4MbDxHV1VDiovNXaIIFeDJrvdO8Kv90uaaW
1QNJic/CXecJX0CXH7he8/Eegd443lF99sORpy0SezzvmzKvbsQZ7IJo6gmm2OSb
Qaf1P+b2axUYmGpdf3FNMSsrbV2Sp6zyDVGYppwAEj1cxxmvzfOBiCVKFSQv6a9V
/LNkgrAemcffvOAgJtbMQdPb4ONytgyKObjcJ+1XI3RFE8z1wmcHCF2id/vSzdlY
Eeyk/2dw/dWuOdQU8By2Jr2nFDps4MJfpYzfcc3xO62EUiVUnQ/3MqL5lgdj6F8B
wjYgC4wLfalru1ByryJdxc92tRvlrPAMKOPqPqCw17JByDkOFdGyShsg5nb4LKGC
+7NPNrYFVWxDj3d7xlskxZTJZ6QPZ+gHlWMUalHfTMWrkK60mQI4ULQC6TwTx/+X
NDoMFj05A9wqf9Nkx7E/Tr1T0xMPgneXcQxlACMXdM01XQEcKiUCG1mX8yu3aLmW
a39B9RdhvmrD1ieTUXJRbpxp7yK+TJqU6To1y01W9xqtOkoayuFbQTuTPKhRK4L3
WscVEBesCF0DjPy0rIJRc4nAA8MVN4eC44IurOR8ClRuvR2y9J++zDFmJanAaxrJ
7dl0cqtX0MshJWI0WLj8HmtH1lhKiUbeWaHbyrnKgT3L70Y8gDkms483QADRoqXj
arYrKUkt51iUXAm6HDZ7Fq7ALRImqPNS029q8Yrz5Sa53O97Nvxiq18OQRsdSm6f
ta6RxjPC226GeKcBvEiYggcmKmVQ9bj6yO5yBoV46j+/Umxs7yy92ya7/0Pd9gM/
r+1CultUs5IZ0F+x0ExR7mf27rv1i5bjNOZhb+a5LIgjn7ie4DfKiWZ85Yf1vVlE
vWrlqxSTrsHpQ3E/7OBA6ui8gwDJJcAbQdImaFf8R35MRll94fvEivkCcg85DlaR
RL38J49vS0QE9CY3RBl0PJ+i3y0nyeoZD0rZnA/HZ1NY48+Y5R7/BZQeaKjfbgbt
DobH0y728ouDeojJChbxlcQ+rCnLgWdlkGz+WfHIt7fUVlb7zJiiAsg0aZlfkLac
3ober3AUEidAC9oVwg2obugbA/CTVndJYiQaxR6/lASBC4hr3WaXnk4JWIgDgH1D
k/RUqocSWbPzyGDd+zTxvK9ovYRc+e6hk8dYvueKW+aesGoONarUnRPprOa3+3qL
K9/arh7LIWtZdJu3/6SHW9WAbFPjfDXou6+rjacHW1052LNKR0ZccAtH2dGSgflu
lE5+4p24xIoNb9/q+TjVR35MFL/+4sKOaIwT7UnqLAi20elFISW+zDkjAlbky+aG
raOV+GTrEhDdmP9X4wp2d6SKokUFpCASACuUCIt5zg59F7pap6xOScVtDh4C3FgU
Smd265emp9DTevI5BMXkHmdZfNamPSAw8oO9w4RUl5buWwfI4UowqyWryrdMQ1iM
6yBZzq+9/pHOtPF7ZWlAJ+4MWZwQNFNIyn5BcF1wZ9kA7X/z+Yvq/pVPgW+LFmVc
JuzJeAKdJnXsIWe8jX0zzsdDzbxkIAXmRLuyU/CquUSr/Tp2VfE8duXdzWEDXpyj
1LXKikOGMSJ9MAefoIicfGZQqtEOzt46HOFbUNvyx/RuGmGxdBaWvii66puG0F+6
KJKiM0Ic9EYHtOtMZmahZR0LAaOgBfciWSm/dTf4jScWoTZsO9TUJGYCP0SZ4/78
SZ6zBwHiCcYCyyqTsuQznbVA7yyS7WxyeULJ39jocIh/7EQyDBLKpI6koPp7QrW7
VS1qiZyjAJq/3GvWyLnHcUIY2cPVAvc+/ssni2k/8mPbM/eTxVdlhX1zWQJvuJs9
tgiYIdQC/s9TA1hLj3bkFmFc6oDy7vAMk6Cat69a4tF+ijMzbselUjseMqgRALqm
qYyNYvHWa511pQilgXVl0CH7ZCTdRR4HCq4WqxJAHhAHIsbCGpJ3yOlrYsb4w33t
qDOXLACSQQxdjo1hwqSogxtISWIDP/QUNYITcAsCHO6hxKjQ210TG8Qpv2ga0SpZ
jJZPuFKgll3PWHJcJ72t/RQsKO+3mCEvw9RC/EnHwq2934decbTnZ3OBCne6aSa6
BC5aqM+LxnOs8Hzc+GnGsIN/ZCszD8V+CQ0iwuT1Mq8bwpjprM/P6sSvWW7rFnnQ
7E58+zLRleOkO3WCI7B+vNNXpbCsJp0kbDu2Wx7hlyFmnSnnPYJxVQqMfINBEan3
3AyPmaxtazVe1kZWngcAMJC3ucdOUvDpMNEeRQiQN4bb+pz1RrDnACd6oW41yz2d
PD64g2H/S4a2CTBGAJGikFMSbHU4HxeRRgdGHKKWHPZI/68P4QqdYi5x/+g5eF+l
rK57CbxLyBLzrNx86uQkOHSJtecuwjCCxbiyPlsEDiJLOt+Z4n90YKpyymG4xvs9
RwbedkVj9t6lCvHNWYWKloji2beiyMWwom+u/4sEK/AD1hyXTqGFYNLnXOwguXbE
pW6nsc+KigzpNfO3BmyNidlBcWV683ATIMyiFdQBQDKkbTQyeOU2A8Dor7pnn6hV
wG1SewSjwhyK+89heKobG7ue2BsrW3+ZiDagTok/xjDXMEMT3DbaAFqrStfiszbg
yKYLJvOkqkmAhRf7s6uRg+QbDtAWhKSIapuA3P6M2pj7Muh0GpChPM+9RgZ1xkQv
ADFlGWPxe5Vbf+8DNK61+s8xlWXnjRKzT/apZs36eQjFtQKyUyr0ZKFvpnsLJmCx
YrVXWKUIFUkU2YOg1jHZKJPpPDnxcgx2ulZdrdvzNeCgkiyIsb2EBUqXsB4DnZjI
MK500kqia1wXofJKeaiRhaeHwOA9tUn8Tx04txrDoJbUmT7V+UFMeRhopKrvyKER
NjJvI3yxXpAWvRBuJGcPJz/EoEnVaXQPtZXzsR9ME0zSOrovjPzOnBl9IyC3HhdV
+tTW0H09bYsZid3XIUcvf2ocRuraHiqMXCG/uNKYRGpi3lQ+Cxx4nlNEd0Y62p/q
F73v7kMcxdk5nDZVhuvOVL+71UPujsx1lgZgrSUC2Taonha+vPVzzf+9ossMzxE7
XWL5GqOuWMHzU0OnAXlczMG7oxfxRRk+LQsVCow/EVxYEQHEM1HWJVYtiDQEytAe
mrM6oUm+joN2qMAepUIzWw0LFa1iyY4tr61CBtxKNTz22wh/Fk354qaJh2MjSXHr
4DXH0fQ1Gc95NL7kLTlTVmLB6LOIfBCGwvb7K/cW3NRVcax/ZEQ4zzg93OTTsGtz
a7EkKMbi/ltKTtf23E8LB90r6LE+HkgiKNiumd3/vVkx8gWcCON7n5lHNL+OjtMc
YV07a1mQZ09EZk3zhAw21gK+W0oPKmS6V+ysQ8aXMD7OE5hyz6FjyJtGiOPSYYpW
YEalS4WRc9JMYlS7BY0/y4h6u210lq+UfcwJ1EjNQfk0DZxiSQqhchoBUhOEzvdS
4SdWAH9RmCDVBZx9H/uo41VylBVYGC0k8NWFHjbIm4tKbSUtubdOdSZkSAhQPzpy
x5MhVXpnradF9UY00Zk98TtQw51RI4mnpuGL8KFlRTM6OQ8QEHV6s9319wHEf8n9
HwmkUQVQMeMqaNnuofxCxwgtGtZBl+WFif5L5Acu7OjrdWW3vvFBhrRd+5/C3ocB
K7BjI57tpAHs1YJu7UbDWRp3BEUqa5OZBMgWyzFD6iXZudDc6MYyd6e+svnKfrYp
STO6IU0l8tAOUHPm9ljv6u1nxExr0rwdhb8EJDychj55hyeRKpiTOUDwNNV3yARp
jIq1SIMtccj1Xj4qw5D7KSe8M37Pa7tmkTN6VAaNQMgPyrWuWoxhUoM8TUqCDQcZ
UAhwpjtNWpSnQO/u0yhSzh1RdHICXZIedq3h/6CVeF0nzuUdi9qtKSHJs9MH/Hat
3q5s4Jotn7vef566UcyjEuxi9vZbceEh9UIRtT0y7ia7p5e72gESELS0m7JG03UA
ni33YRL3PUzLlfn6G+p6rxl5NH9Vya0aWQQl5J1z8eQADjmi/073GSZAp/2s3ps8
TmmLbEJnScGh9dMT18oDUlAVgGyBcq8VbeuEKbx3S5rXNY9ijz5xS4QcLJM0TA9C
rT1wwiQAG0IWUQ2MqxW2ibA7EtD9VwlSRy2g3pG5Z4Y5NEBxZBt11kmiXxAVSXUe
KxD0diwqENf9dEU5Bj1Zw0OPBdiLPg+U/UktaYarTBq7QbZ+fkwE9N3IXTHL6YhX
Ml+B4TWN/cS+dpZcxpXYrI1ZnCNNuLywgCGarI+o2jjMWo7tlQGvTpd084i0n0qX
hp9xLHTRSo/WwjYYE4jPws7/0QLwACLeIWooMNot3c+CgH9Hhq+LlNM5KPEDN8o9
QhRb7va/mdJuirRRU+ZJyUX/H1Zjy2OnRnFhLbIOs+ANzOf85on8hbNdd7PThyuA
5A8hU4dnYd7DBBtWLujz4WJrQpR7eSd9JdWZuUIuYvzTe+2DthBKraKdsbQw4li8
n6aZ5WKCHulFXATUpNi0Wc8J1yJdRmTgD2dLmj8IgIgcvTEWtyumVuqdA+KA3ZhF
5YigpAhMCP0dfxsCLLAdwZaCwpT9zD7vL62unP3TLrAHRGlJnAyeNCvP5Gy2XPXP
cS4SvXRYJTDi46GlrN43ZjSHhg58fkGg7pxc8coEXxzLYQSLWsWcYXurY9NxO4Pf
25Q0W5QYfgSUJC8Y9y8k3wLzv7uONmghjMvUFlVtWMWF+1vXRqvvTKDtMG0qSUsd
OEDkiszeAQbdV4l/dlDmckOd8aJSL4A45NjlKrkpFkDLBNEeRept1XQPsxDnC+OA
/3T2TPkjdRIf3ZlF42R026ciIZb2v9644KZ7UvseJx0I2qgXJ8puHLJGssIYaTdH
+KSOQkDDb+AOav1yBa0t+zEr/SQxG2XDOrrxU2bXbQEQ2la/J/uFDOSvb2UDKBXI
Vm7rXEXs0uQTwb3pTyk2QxbjwvAblpvFt/+yrEzUYabqp8gXQvkWPzC8QSjsgpRH
Ex7WOBfbyHJPt9XPUiUgDsBzxI6qzC3Z5zw6ngkA9/kreFcTD+qpL5Mts2g4mxeQ
SrWPdSTYC7xX3Ez2h+iBU2ogmUI/Q5U1a8lCmeFfkr03pcQChqfvHP19853hamaB
0zp+PYjNEfq7osTVDF99bYIHLsujDnTvrQrClY5qcNfK9zw4TB5AUsMW/Jmm+Hah
hr6FvXVa8RLnYDBmZ0Ajl/bDRBKvmcdVqic6iHfzx/ULkDE4/QVLKknlnhPYq/5U
VTNRxcquuCW0BdjEsNFtXAWSr7ewZ2NvxjAAFuTADOAu76erUXGMdsZ9M4v9EZuY
bl4GEhpCqMSjOpTzZBSYL26fhMGXKTA5sdbtXjCBfmdrX3reT1he05a0WjC3tJmz
rl+kTtlzTIzA8G+N2ZYwy4cB5bB/ooEI6OJGISBaD4wjVF0tNC5JXB8ZlD6ZC7VM
+/fK4RM2GjlUTDxPJc7QRjlgfk0IAHkyJcgxbHagw3/cVPZP0QY+BH5MFpkHHfw2
G7WDuyGiZX4zIBIQsDhG9aONgpVD9pKJye2OqV6Jm6PuZ/m4XpvWb44ZM3kP+R4g
bghG4HBWh3ZwL4h1dcpSvHP7ruddXjOOntYQSUlNRoDNqB35v+84n34az6cq4bky
fczzK/9D0AJSg8nUHcopM8JlvyjbTLYO8BcOb3/95pD3/obINQEdgQExnEi1Qepv
6KJQGci/OpP6rJNbJuGwl816C2zkHyXXgwaqXxrH8ryjGE8+6GnmrKFoWH5egmxZ
X6sS05OjhUUcZt/GexjdrtJRtcFCrzZWzkiiCyCN9QTuRGPS+YQf/2Hyt/RDow7g
wS3Cjru2CMJK0rQhmAHt2ydaxIZLsxwh3xtr4XwA6K5GTSeW410rrWZnkwivo8z6
vQANBENVd7iHpycxCDcmI7fcDHOQzQ9+kkiGj1uWxLQLBSlewAmgKLoM1To7rAQ1
sAM8f8dhrJE5v6wEzklh/zf7ZNJd+BGlzTcq4amKiQ4VOWLkkGkS8ok6c5eJwtia
ZAFuu3OZC3tb6j1duCao3i7nTrxBomYja4k3NEu3ORdGHc1KJarBi5IsbQsgp1gg
y6ERWg2NVvN+YGxy2hqFCwFoivhsSkAMCNZFXdHZOp/bAfhwOMfW9SZF/rg4tuu3
RbUu+PXSc7bWo0yGekTFaiLoENb6PYklx/vWaoZ0epw9NRuz6V989yJtAd1NzGfI
bcVWFtGhyVWurx/7+9O8uuKpGiy+ykLXsqOObdRnPaJwdDHz9jRue41XFvW3FZX+
iIF/vrX66NjjfUzDYQgwJMz8SArRbE8BWY+FCvi5uscSEvCdfXTjXmttxegvU8tS
oFUHvFeNUt8WPsOPLM7hNCO3YTIdqyFQp+TKlLVdlPMXW4kNOBuegtxluWdNlNGT
gobyhQjqs7JsIVod6gZq0ULianMScQjagtEg1fPlFoTyH4TuU4VtOqdTVjl/KAsg
SIKyN24Xt2z/pA6Fbv4gWaeQcNNLzcdrmW6K3ci7Sukcdbe0tV4dCjc1hLb54AhB
NFTxaOjm+jcPZzG9mHMgTzXNCDBiJyTxNJaxmP1hArqttdsOzOfU5pHycQS0FSJ7
DQoqBn+QwYoJ5S67rhR02stYP14xfoFyh6aAhOe33BlBOVF/gALAUphs57MXM1wS
sQP1eQ+MBjM0wBfeYucYZmdK8EQZqIywZNOevGlslJHW48DzwG5iJ9zakptOp67k
WB/M21gEEXNtW7XEYxAsfesDK6ap4VT0CY2OHtLMZd1vnXFyAgN1JGWWzvdNR1Pn
DfdK9grzXUHbfuWGwElDgY4P0VvUq81DJEQZR4mQiCvUaM8PpqPZAL9swdFdD0Sk
65XZwnZ3Sx2O5N34RjtR4eb8veflF9Zo+Di+R7AYmusNDnDr4pBMUgzkpDCXU1OL
cFdorpoMjTpYTCr760f+xvrjX8DAwiVWhMFvnL08IME9Yv7VriRkbR8InXNwVtIX
4c05Oi9t2W0MDELajBfKOBbhbmr85FNZQPJ3Mk6zaDx1d0TTWoWmJeRqt2Zrauso
RKoRIP8OJNk/veOS6s81qAMn0NmhBGNqjiT3tMZhid/nA0yY5DWSI9UbIcI46aVU
rCB/3BKC0CQRfnxV/s58pIgmPjdcH2IZL7R6uJF1WasyQH1bsCyhnPJY3fhghCRX
pLBK8rP0+10lpdKCtJjlkYljKzt2ohbXlNe9iSNMrsVnG0rhuXT0LMBn9IM43z+g
ExJqSzs4uf7OH1bTVB8PTlzU+u2UfuWs+HgxFgeQZsB70/pO86hf8fTUcI2Vhx4K
QZh/cqjplTWh3ck+mhKjSHbRvndDdIIp6Jk6GhWo67lpPrFMXnUa0/4dQZhwJ9Pk
OMJ83lfNFli/kmEtoMn7uYByfHPdCl/GsxNa0hElRG1QDMwv1y2b+sztFFz/oe7X
ju1lkh/ccNqmCWFb6+UE5+gw0bV1iksc+RafCgwPL7Lv/yXOUQsRVK4Xpi4h8Ato
8OnczMlXkIOZng/sRKs3ST35eWT7M+V0kNI9KOmtVUC7/tPvgEwBPe9S9BSWwkyl
aO9LyKgZjLjg8OsTs9RaDQ+2gFFWfhoJTlTqFpVtM48bWwHrlCUg5PX6ENshjAhp
Z8YH7pJZ/tRPxiG5VGak6dhJEtMQm47L/bZflwYBkEampZwcIm9oszpOXr3MDZI8
KCuuq64gg5BTnTuS8lz7dD0cpKnNkO6bjpPj5Z2AdHVg2SQ9g5Gf9+20U6xbKwaY
WRIUyfKpAoTrTeyc0vc0asEOmWeRDulSHyZUH3XgkbVd86sSDLvNk98scgOUyRci
07bZRBI8QDpClLxY1wLPStmYdJU3Q+694U9ZWzDKh1xgVoLDzleCnogkQyqNqjTR
gQ+DcwXZx7eD5+JSRUb4Vbx9wQYSFAasHPlmGEtkpz4QeX7tVrTnnr/P1xRmMcL2
JaiOEUcMpCPwf3piQvH9YLbZ43KAUjzVYNBADsMKR5LmYVOfSgH08BZBGV40YMg/
Uq3dZAOHjavYKxwDRRxGKkxQMytMAUmgMKOwYQGF5g3xZJlGfLgd62miuaEWNfh2
udR0W0J6bBigDWvEfAzHq+iPrC8T0VZgMkDfUpWXqG3qgo/F4F7ePt0vVGOG9mcQ
bZChiFMlDhX3RV0OtZx1o426ELL73MpR9NUJ9Sgeolz7pxmHraXwI1/4+83L4wnO
flrkJMipcIGhXJPq3umwCiRXz/efcZZq0zTQ8bsngqyfgM4d2AemArg0yIyqlSyu
wqX3i8qjEt8nRVk2cS/Ol2xPkau2opWUF0SH3TDmPUtA6U+l58e3wrxrnVWmw/rL
y+/VDC5ipARCx+Mm+uAH4Ugvn5aSodyTsHIN0O+NcJnEeRxFWeELBY76rJeHuHVr
S+K5GoA3L9pFki5pxluQKlSmBlxRcPECr0F/3W/p3+hXG0uiApk04vlgHFQzd+Q0
6wJdvkJ2OqkonF0Ol/tcFgfrcEmacIggMezzbtVY77OhgJdCGOo09XJk8S+tSrf5
eNwFM0Ho7Bc11BGQSSAps7dbVzpIvv5ypVU9Mj6fAtSG+BzTBoMoRjCRXUiZfQ2o
bWimSpGtqhi8bLfFBnKSIyp17kRwhZcJRMlZJyw5Jzaynl3bsBua2Foa8EfMkOi7
tC8psiWKZEBwB75tDxgUTEWlARRW+tZ9MVHpOPrnmV6b66Ir+D3cuzWdyTpe/I+x
ppD9PpCEFvdwKsu947kRHKEnuatTdDcW2RtC8CSwfnS61Dbopwg6/vZhJFOZg06W
hTx0IHdafS9GCuSnB86oq3K520fBF1zUlv6aRgWuVuY0nWfAEj2mFzxw2B7sEecc
olXb3BnMC9Q2bjq0lEWoQWAbRgCxOlh7grIJ9XptBUXPpybGuJWSb+2ujVZ9qG3U
cwA8EBEPrJGaUEP4KNsGgQ9WyoF/WrFlqzcyhnzIS7McyblyQ7NRYg3NxZ0E0D4/
yOtgXMTBjeSvQcOEyUOUwbDW/zthvaEGsGad4GnpC/utXR4yd22l+ux9CZ0XvghM
p9DAipF46ogV1oWu51SLG1mRLfsaWLmMhMGElOw7jRo+3V4vED4VWFwYlCJIHhrs
q74fuHPkdw2fGnMeea7Rclc1bZoaLxMIvXnCnV/55ekBz7fT+n+JtovbHnBCGnUa
xEem9vcFlk8kcvJS+bj3ttlt9DXDvXXjHmN3fiHxpleNVitAhngTePZzF10uhozS
FrpxOzzTMUZE1KObxTWLzAtuLj3veHowcTMwIKT53IdN3JNviuqC8pv7r9mrIKrn
p+89S7r8SyULw2VXxbejS9v/aLJNcTbyErwrN+SEP/4D9aroPN0AZHjV1dvo2Olt
GlCBbfs8MKieb+q13sSZQB+sEmA09pLUeYtrMksvTiwJB3aSSkkNQu1EyOuYJrvi
OK0QzTt/2LNw3q1iOuqNOAP497KOXu+z6NnZf0m8aGaNS1I1UTkG8FuPpGEBaBD+
jeiPtymwdV82q6B/7rh1moRRWYVgLDLZoOQhvjbZFeloXymxso07fmkeDt65R+zk
nE2eYgx7KMg6xDCwe307DH+hrWFNmQibiZOPhscI//D4Z0JcgTSQGhTsP8Ymiy2i
uPS6teJIh66ijjAsRqibcsXrKaUciSpckNAu6k9sQ96EodTuXq6kupwsFKvF4EPU
/NGuGuQRQafWHwGFeJIH433YXHY1VHzFD39E7hFseiDunvtkP06t7Aio0z5+vkVB
OavLCx4A0azm7fcWnH1UrxJLTM8vA8nhCBjmExdOLnyj1q8boH1XRT6MniAv6oCx
Kx0E6X2xV6VzS2X7A/BjjcQiSyfI1tuFWTD1cyB6LUpb4lwxqnJ/03kURJbruNJP
eIbB5a6nU0koR85TLGjlwiV7h1jc/QEtzcHe2ZSv5oKuX9BYZzyN6YocBO6bpQtZ
HfRlofJx7xDHKGzkPeEQ2GGK7CEUe0em83MB+ZD2py410fPFh2rgDoFyOj/VsZtX
o2Sw9AWRExi7vjP2QrYRxPbqhVjY8BvRoJrttBLkGbMjOxAUWSoQMg5swWiBw6n1
GR4zVwg0xWRS0ajUjw/lFBNrFnrMdR6pgsWdi0WuOVwNURjGCAbdJHg0dmNQjk1U
f0qk7A/Uzd6MbQM2oX8p8qfTM2RMp13eShKyzJtrOGtDC42EU3SDADOAZ5pjNN2A
tZtebSrpHS31oa9JyVR3yDtP4DQcI5Kzot/vugnUZYQ+ITqVqog5law1iW2FxUuZ
C2S/UrchmuP6WH68cq0kBx9HZrN+VcIdbE9NdMbUOQznmcwb2YMu2pDEfBVkMOfX
UiEPN3Vg4ng8KIKzEvuZwCv5X16U5fE12O0Ytby46JeVcXKpRqWh6HWnftqjcutN
VfHimNswE05o3l2/mP5NCB6VyfTujufhmMdPBK5NBArtz8jtrt7DhQsHB0awPUgF
JtcS6COGd8fVFIejE5U9+VkVSNU0ddcdPMeHyLiFYWTupbTSBkXJFUT/WTOZB/G2
DX0E+p5q/lHt9vtu1MudtinebvnHa7WpCfQUlXf2wX5cRPESQI+ZpzWS9kYDIqd8
G468odY1dqihLqKtiM7QESoLP51IpJUbBz++NdNYFcnOLARNFLwm8fuXkDo8xEdm
hTjkRmGQcF+9324Qwk1z3n3g0xQNmMdiyDDRb34Nfvp9NH3Xs8fkFOcG6HSApf2u
WSo+9j/0RqrK8se+xSuBy5Lq5ADMBBJQ9+P84KOINjuM0YZWSr0SNUHO1W6DMkjR
lChiMqJ87CrCysFHZJcI4kgF+eELpMM7OdChNFA3RdYu29+zmXPcRtSnPqCuC7PR
p5ZKIt5HJ9T83RQbOE96uQTiNFfRBbzGTWHBA6+2erVpWsL8D5R3Oxhnu7Fyx7D8
zk9GiZ+msGg3cVdRTswPTFoZPCYzZR4cIJ3kS1Z3kMa8yqX3uyXqjRDXKpqk1JJv
EaFnoPGGfrBHXFIri00i6D99bJkgNLibt5fVUY0A85TqNrG7urj/tBm5GDvIBzil
GQWoVN8wyR+FVn0LILByWQtsuVDR5Hf6ICac7fEKAbMqVp8+sGHH04jNyuCYLHac
dpwX4mcsOX2OQVjGq1bN0W1IQa/2CyWSqVMF1QCVkv7bRYr/7AjhpMPUKxk3wfDo
XDljjAhgBWZEQrrjFBhsZTR++UiVIISjUvb1uT7wtqVBXonbIj8U/Z7Np80D6x/U
uVHlotXHXnxQoFMbN+eXIy6jTpLNfoZmpWbBdnMkCnD5glOcEij9RqSPCtHG5y9f
xqCKk34P9FEJyoHYftHl4Wo2K9XhCnDVtC0IUTjRFtvcg+NvOzyoDwHUnBJUoT8X
7dmarePkHoTlPrIiLKWxn05KZxaIXfc7llkpAers3rr50XBxK1zweVFn3lM8wi3d
/kkgyE+v8q8S6RoiAibPVP4ejYzjlA22ZeOtSdjp2NEwz7pm+RDtFwGwjjhILG75
qpU7siACqOufRGd7aHwaK1R4bY6aRpPU+RNfTk2pRaMuzpKGVcyDkbjvWXdLk7o9
V2tKHo6IERoOMouqAPoqirYWD87axKvzQOX1WQNPIGRbemC13X+zKRamopCcTPxi
LIVCM1jYepUQjiB0sQOnP+ag2qjPYmtZmgYTTOWuazQxpSVZqP938AUbwyVTMBwP
14gdRbfGBljAZjGnjjTFMfF6MQQdARAIv5AjkZDNPY/74f1aTDLasP/GMJUeHNFQ
dWFSCZeb6/i1RIhddkzAfwxeMH1wxi3jbxsggrgieYl6rtCsoF8pBpbm+ZuxNfr+
2XOnjxrNyjjHQEOVRQqb//NrmHexwTG+webSIJCUUiJUEACax7XoAvkQPsXOAbq+
hq0qOC77+CsfttaQUIF+w2KYFoWqs3qIsgza7GplPt879mFO11a2FjLN9W5NopfY
LGk8Bk2MI0SWBHGH4c8U8xLBmGYgnHH47S4dVbmjWZZTpywjUFhxcX7iHxVEqING
vl+ArYZsEwSO0NCFc2gWucKkJum0OQQNS4Lq2fCdkFERA5oNcdyPXvy+6Pql+ZDd
/1g8vLhoN6azQTHhPJPLigDiM0JyH1lXwQnF9zZmy3e8uohpN+wpsZPo0+Dhqfk0
5sNfiFMP2wQaOMeaSgvxJJowAAmxH2EzTYz7s3n6NE4eEf4uFQ/PYy0yXZsTUd6/
8kj16zs55b/RFJt1XUVkXRt1wuu3Mc261/L1AU6iVfeuZPCZzZDphmoO36+Gkm5n
txw9PuWg7dxtjS9PrXa80mD9PG9tFkB6hw3ewWLFhv9ukvRT0RyZkNrde+Zt5N9x
ABzsKDZsVF8F/Mt4Q4isbN8XwlkyKuMlTJcMRjTrdTETczJE70Nsx13rM/dRCY4R
c3foI7STkGFn3NQ+YEl4zc5Ita50/Yhqf85VfpMoiVqgcD3WJ3mezu4M4J7Leh3u
iPZ1fhcV7CEuqaFI48n5KViiWdTsWdTqf2DC0VzN5NzA7tboEsv3J1KX4yksnthG
J8UXq9YSoFtuqqr9AKsvoOz2KA2yiLXqO8eJfm2rV4dFOsONRWT5jWhRk6xjkIeX
WZFNdHiIuCgSkFWmjOQy/K6VOK3/3BvhiEiofwNUdC7a8mDG79fct3mOtFpWqK1D
IKttHEwpplbpOXv1nwNgvaVGQ11PmOGtPHGdJ63H4r/IdkNpUZtb9Iz7Bpoi8Xv8
OdlByxruNzMjDFwbTOci5HhI3V+5Tf/zSpz44c6Eu+zf/cG/rTuuTYIE6sU1jD3U
1z0ib4P5aM5oqnP4Y0To8l4FGaLgjYORzuZDP+CMprD8URaOaPq92XjT1/FNJd4p
pWvHbiCbDC3iaAy3A1aP3O8PA7s71pftR0etHrbgclo0fRzeT2neMLe7f03EXYV5
bpDL8Mo8Sxq7/jIEUt4olbK64QCcSarEvqQRQjB+zuFbVoV+cySg58NHKwl9HEG6
yOX1clUXKnjXUwliaIkVc9D9UdczjcxIt7xaPKOz3qTg3mijXdO3Cdja8584x5nl
j3cKqRAja8RdrDiZZ0TATE1Lym2m2Z8Qn3Cmc6cGKFNfjZBk9+2iPAtLRVCeSRMn
rGRodDNkQy+VGjHVARAQUZFkiwAyJEh6ZmCOZ8Pxpj9iS0P1wRiwS9FsCyethEg8
M+b1FFaY+e47+eadZfY24CkTzATEQcsImVmlRYWyzwnGKHEHWZ2UrTUIGOiEYTXf
FBnc0Gdunmz5qhtRoGJpE265TqqRITS6VJPrqAoNspS4/Lvh9np9jC6TQTfznJ7p
ZEs3IfnqfnuCaWw7xdICJ9H6OIEmcfNoNL/QT8h9n3qnkz8wS4xaNiOcmLpXEZMx
S9T32a4axc34AJbwGejiXAyCMIqun6ph8X/wOy3Qv0tNS2xCPyqLenvBBbyP3uqA
l+bhSooS180UbG6VPmhjGeqfRs2eT6AEoHKmg9PQK/GiZpJXruVkv2CgzCJOnQun
a9xuNrtjrFFHt45OEHCq3m1QvW0RM3UbABCE5QCw46MXG0ARNCQ2TL6PU8nZY/q2
8nBD78P3V39ZMocpCfOt7i948YN5bWpbbCoDtvc9cnviGDo5M/MBTb+mF1ncuknC
LaO140iWfDDSgjxW54XDlnzYPLGufH9Rjn6/SbltIvb5hUWVHkYDj0jLSDWwWA43
ir3Oo698parJTIBtWkBrHC3K7slcz1X6H8hA4TTpYFJ4ps85CfB9EvRnklC2vZDA
tesvoLq/cERGCc1hV0N2bRaJDeUnZVO/W0978tLWgOJd8a8eA1P6oWn3VMZWymea
27ZB7d1cBJ9jeJaSgWP6L0OSNorDg0lSoKB44jLc5wrUkS0UZHfq/3FpobiK/uxI
BHqSaqCjo0rWLtjPNcrYwsHB7P4FjFqJVi5XnStFIRbaW3sRDPokXn0uLwG80qAn
zrI2LfYt5qgxDKzY2L40yE0OO72WstA/gOLQgJfgvD78RG/Rb5HJfQT12xaHjaPh
g5P6zR0kzwSRRzsNGzgFIm+g3gC+fsaEjdaBJiWYimozytibpaR3sM/11JpJoOIr
JxIpp2l1UYgwMJHFBIBPwdr2//pqvVJvatOHY7//kgyN9oGEoy//wHYa9UB8h+3l
6Jy250GPDLKtnyxlQ2cpq6/Fhd7V/lGta3YEmunagNARXRK0ZKg7TNNpMZB2C3/x
yJ1rgakZXPdRs4I57WX5dLVRLhlQVQ764bKdD7iUsMzUydqME5QQMCUdjnmeKVz7
zsk/HPgu5TXsSxZtNQ7ARk5xLuSQ/+flOwf86wDVsWK3Xjox7WEQjkAIhrJdMC9d
qBzGZ+M+dssLUaYYdXAAGtr9k1wNexpprehkY6rRArzxwo6JBnmwHzprxb8hXUPn
23qarkzMsh3dRRRZ1dRghGg73ww7QT2HkPNh70ndfAhAGiKdzrW4+di04xRgnV3R
bd2cpZL8kflRIN9j0g0tXEK7+V/GMZWT575eVDpfKz6kF2XRH74cCGJ64ThSH0+0
jJPQ9znWXEs4sKErxtzwrTCw7r6lzPKlDq7GuB2GA2F9ocrxHRk4AzLOJi+Xo4Ci
54WkayL/LRJ/Lk3YsWmB4SI6yclVBebD9OUsvcxDz0yL6q/tUi/xGl+riqjazvsh
/n5D4O/RjSI5G4kNt62t5hEE2NS1CTNqJy5Vat3r2b8WU3rsGkQsJOdhFD70/KqK
SWYsgt5Zalx8SRHLfXqfyVpn5Zakp9CPRGe2DcLBzn5l98UlE1ww6zevZebtbihI
21i0+rM5G6eNTlhASrXeygGJngfOBD810U/p/imcyFku71YhVNAu/GBuTVyOYis8
oCbxa81bS6mCpF46bYiFrj4HC7vT61ayLPgPbvITf1HCkFvinGRUuDNjjBmLhr1K
oQ+XAwkktTMyH6y+nlVVSDxkL8nTyzlDINMfj2ddMcckRuIxRMdwT2C3c4Q9PKMC
pd3s2QHekMyd0Rkdq67vnDmjM+YJ6sn/52ywF6gWImjGJ6dhOXb7x/SIycXIP8NT
7i7rn2tFblFZLXLD0qlKB0Lo4cp+51UfX5MhMSDilGqhufiWF1T8aaBVgPKcZXj4
QVkcAWUn/cpXDgRSsvqQ2Pzuost9/R7VMr62YxnXIYV/18bxKrU+j8rjT+7IsneV
HfLiPbrqlr/3QP09TJCM88M5YjLebgymr9UowXRhb82CNVBk3P0gr9cnmmSoCVTe
ccY4p9JNIOM9e4b/A5zj6c1movsWlAdAgFY4EK7CD0IJ3iQKiOYXD0B+/iYffeEZ
Zv427NfTIqJ3dYaAdLtDcuGesw/1aoi5RVqxJP7PACu4p1WmAb4omu1eRzWdwy+e
AaZQRD1DN2/LjtJx4sKx2x/uY+73/v0v1iyHelC+W2zEoKHPK+e6EmQcpv0nGBTL
ergCoIEvhTlw4rWBWEfslM53tEnQYzADN0bkyCKh5xNUwTF/Q/wHDsu30TVpfElu
4G01LlWoP47h6wfaOcKphKyoY996iMEmzddAXIT855feztALbJoJEXjmXet1/Ezq
X3U2gSj9A6WrWfz2zReo/Q5I8CXnUA5t/cOeMFGsXqDPsjcpyCWUV8DpCGVFdAKT
tWzB0ZhrS4KZPOAIXW4rlsC9WySJ9CW6HUNbSCxknI4oaOPlySnbgKdvInc3EaDK
/5fRQk4reP0r4JQ5DKNi4iuTTSeG/lq4AtPzVcFEATsEE7W0Qldugii5w/LEJm5Y
w/3iuD39wVhTAdMas+uL42bqScGoiRz8AFqtpZ35t7F9v9Rgddj2wkQ6mQJ8hrB4
hbjTQBjCF7eHVLgPamTNik0+xQBN1WtBOgJziMYQlnKZ1gq4BJCUmOmHr1fdq/jp
xl1w78hxdPk0AqyFk06yghOrJtTeFvhpVtb/dmrUvCdap/ppq/VewX7JcmFwutzC
T8J24vhZyTzdf+NbJdKYoJ4LGXGmqm4lILUYbjghNEqvNQ+GZZRVfWF1pPvwfWlF
ssBVshBAhR3+bZsqby8otKkqn4aK+m1e5hWYYkVAYAdgXN0ftgmwYxQpqCJ9k/7q
a5IusAaRrxXr/EHewjsMuPXKGxjGoz4KdHbQFPxo6+jnKvelKdB+Z09eX3NHle5T
mgeOGBLCipflD46MG9gDLK6GRp3JQoeuS0aIBDHgh3PcrwSmbVVTIVOyyuAjorbg
RIjJN3OSNEEyCt2bva+5N5kmY8ZGJvUkQ7SHu4P2LVOx8hzMy8IPsd38zi/oRVnB
AAv+QXPMtzmDb0+vOleLUFvUKsEb7/W3Z0yK91Iw5rfyaVYmdD0XemEki4Aveas5
4RW3Tj1ArdS4zY58Y65S2h3YY0uQFWno9rJR+ISWeG0mu+aHzT3WkiMxl55OA+L7
lf/EONn4+pSeU2BYZGhhHc1QaAeyCmicokldpRxbdnp/4G1AGAIjGiFXPQwi3Iap
pU1PlwVYnfeoqQWYLIfr6c1/YeJfncqTPhyxc7VKTlUR50RPT9Df0a6F8Hf8v7J2
lY0INsSF2DO3gHOwHSP+hFF8IcOVmS7xvMbVhntpgprLJ3PrJuwE4ult+Sv2mkTp
d40/xugUMnKzdi6vYdWDb2FAYG15Z4caYgW8562fW8nlHsK4TjHernC+cE30bZ1q
9NLrchg50lNLFQWWT/53ni3aaRrROXpzKvMnH5IKebfzP3avsUufGgyNw6S0Ep/b
Cmxn270kZkTYL5jFzfqhpt+WsgjDDpkjAzUD8DqLNfMASZb0q9uQsIw3o3fFq3o+
2kxX2lFxbnqle9mKbeVcA1FuWf3ZpLWu7amO2ushPNRK583yZPtK6NMTGMT3y5Mg
OvsJegFBj5483ZXlePtgBM9BGUkBYJ8GDVblGqAS8vn464dl8lsiK/9XQChgvQY1
4SjdyGvI4Ubt9+lUs3KyzVTAx9eYV0lFiS7NfKkPb4OfiX1FSEP9PyszmfdKfATf
eqWNklFbAMsmPJMILsC/L3iiQ8lLAcGjkd072/YmJiQXi46tghYdKqxVHV+IidRt
bc/gJsQE6lHlpkavJ00vVr49JkYjdvuCMOse6xIUpdHg+ilvqvMW2xo524lDAA6d
SNCHXwd6IrAj2xzvYbmdxZBmdbfjnxWkQwJwTDvLdG5VBCBMoe730+7UxGh/5aIi
FtmdlyNjgFIaH1uGAf3AoOJcUd7UcLsG0h5jmbuZxlP2XCzFqzL9B5goCHK2npPq
zvLc/OPhpqv3jcYX2pHodgunDHoinJpECVoS5QnDpml5/b7VwITRp/q7HAKG7e2I
6aDRRVcL3h5s4eApWR9WDNkAUburhJhQe6xYMUUYOrhdtxAgd4kStINOZRVHBpqh
JATxVfjvC6QcR5HFrWBT724aiWvkXdT0NrvPnR/eXwub/ygifbs0zXyyGm5RYVVy
v8meWPmyx7MIR5v0ZvMK5E86c31tV/odGP64int3f5WFjAvMIXgiWcQ8lFsYvuRw
zpc/fklh+C7XJfyuyndP6s2Dy6e8LI0kKVaLxW2buK4gapaaS9UmAbT+pxp3RuVp
AMqTZR2T5sKCHHWdg2D+H61DJn4h8waBhwLC7z2TwUhWa3/hXYAN+t0q/WXxI29i
RkzVakEsOy6DekrSehHoWNmX409J3l3t6lP9g8brlRJICgysxwhkRBv5rfQtchib
Az4sKd6Cy2Ihy5klJ1UDHDJzuhL4ZbJVrzC/IhP8Wc5ysuDtxCPHkYlGk0XDXZoK
E2r1r6gVmqZNwexAqBAqdo3E/AnHxi3Gv1mreP5iNwBJJF8cA1evx62ECb/MUaeM
IwWdDeXel25WVNzeSMS0veomTnGd7C+jgFBHfudmRoZaM4BvlLJV6Ylunz7SXqeV
Z0rk3ycAiVj3LpO4IW3oYMCzFu7xhWmu+PR3u6AnJux9tO4Bd9GaG2lLGOVjVoRp
B54hcDKoFsuYFPXKLweXCP3yrAleYGWMVhiEtefYcZeoc9NSc8jT9ejpKYcMhtXn
o/iQT6HCHZ1psvGPugn8qdE7YPdCn7hCT85Z/iWTfJMGDnPZTv2zfI8lp0pvhQaN
tqrsDIY5VmGEKIjFtfGCePgifnm0FYrSiUkI7mrXr8WTuYAYlYJ8psnocmCFIxfZ
iljpNOAKlxsSAUKZKPeiwPZvQbZF7tzboWK0mjTNkWjjKg0556+0U2JrSoQErp7B
8EUN2GArlVX/KirC/SqEwy0Q6BEnWCqgiI7XHlDZG6qv5oBU/JlRMRwuLvQ5WKZJ
b9HXa0/reg0ZHHTI6EypzznO0pkDi5S6A1iBfWyeXub1qoGfwNte3E+o57HurQ6S
Htaa0xXjDqU0T4oJk3tb/hwE2RarfKzpL158cHzd0/JuevRnRh35n3+MDf3vnw42
y78IyD3ZdSjJK4bmbF8MmkijC73WFFmRztrc2NGY3JASo24q1Y1gb6FkEDgnwgWb
bMNw7lJS/Szm1xntv+kP+pLYMOGKtiDFJ5fZU/7mUYJvdAzj+1URU0ZVCDsEmwdw
kAEV4pxXiQ5yQdxmJh3UNbNdpq0N8bcvgcbW7TNIdw0OCE5+f+9i3h0a30D+vAG6
5Dl6inAFMBUQTNMMvPD6zVNe+F/cfZZNxIA+i8Yqw0wSwpN9mJitcXRizk3EtxWq
XNvN4pug2W/CMWD8PG2sT/EJUmjaVGBzadmKv2GW4OI7DrBqhCVfgSfXKrQuHiSn
igBRV9xXzMi0Q/6yYD9MNtazwtSjRIXspBbxxa3j82yEMT9qoOdX3wpluvcJOIYd
YTsXXlrKySuox2916t5eBen8hfJomMTrKIdhPGrjas7HgOhfsSjKr8wZ+7nEqY/z
qSh7SMJWvaN5wI+siI+QIoqjpZ06DV1K+9jdJ6Z/wWSJN30U1VrbRtCztp2feHz/
11vocpJDuKA8ACJ8rDqILm9ZDq3RJTUJ2fSpok0n6MfVNwHMjUH/qRw03ZPmp58u
QsQv8dZq/tK9eQvRB/n7vXWksAQ1ZNeak3m+9SwrBVJ8LL9WYywx6665Nv/LGIuf
1SMuAe4QPEgHIwp11/fdGuQjhKuye1pWAZMJcU6CK10vUyH1SoBxUh/Q2BZTSLBo
QwZ/g0V6PCvwDtgTdF2ECIx7G38wPPBJa0YQ87ASm7aC6AaYfUKLJdYmV0mGMjUs
uCOY+KAIEWHozMw8JTY0420WCu/v9VhbxvlYTd0d6xcSRrH6OTl14c7IkPPamNa7
yk0CANl4yIMLD9cIbdf1/eNYkKUdmRkirMwKZxN77umY/zoxIHJb1Q8Hdi1uAsr9
89DLZIEdK3Kkyf4p8osgQsNHuJGKKx/DV02uk1SVQXNUnTBdme9Nwb+/lxtxwfou
wSFnMgeHS1Pk6HJilWE0gs3u87jQcdKvMiKB/yDS33IwAXmoHXFtDNQCDuGa9tol
uulfjUautR9Lfi2AvMfNw1i5fAURkTdwkyrXzJrQax5gnUU/mDgCrec3LFf0flvO
Gi2YUSXlISDyZE8aZ7Mgkdgf+EwE2q5Wd/Dh3Tdcr0zhCogrp6slu+uh9SYZUHPh
PXiuRvNN4efA8WRpu96E68Vddr8B3ejr1GbJbh/ExMfFojyc311O9qlpDOVOZaW8
e7miyUdfAdnIjz9KjCpUjT1aBk4XZtd4wVN2Xqb889mcmje0yf5zGNEsahkVy4Kc
dosX05qy8TT9iK1g22lEyf+dpd/o2Y1A7Jd+HOEyMYtYNApNG9VPjJhdXJiIXcsN
cddNmp806GsI4KTB+2JQT96vMYlJ4/H5Z0qgGGSzGmqDvQSradNncVuikspnUWJd
RerIqzlOQTKMq58Y+6/2uMnoNGVwCwGSZWQig+QlMiuOtKpqhkfuzq3FVPx84BEd
TCVvI6Ez47MJIYQ+4Xak5V7Uj4HbRzSldImnTY8oCX54gyvmFl3kfI09IzjXo+sI
XpVFOYw6wS9UvgBcDujXtJ0S3Ru+7HkQsJYEJN8naQpgTqjCZLPJo1yNAWL5PtBk
MNt6k7OypYAqhEcIDzRqZ6C1H31xm1a3WsladmmcLiLDRUgXdzdfDb4HYIkjEgvs
2fDkFsRiUy6kAfqIYQydPsrMjwYnaJzTmHGCw7rN8J03wH3fjOlcoipQalAC9FoY
xtIDPz+pbfO+QIM9OWfQdz38o5PBzBIEXbBRHD0l/WyzSkMae0SfPfQo2MgNpdEx
2c9HmcQ8/C3yid15PDddyTfC/yc0PgjeLu8EypFLf24xQxuwqp+frIAC6Un0afAY
8YGHM+EF6qqeTrXIPA8ScfCx8KfQluIEuT02ChqG0fXt0pYDqC9YzSZGhI2wgK6N
AU9Zb01EpH5hOu6OvZnCME5+5SRFeC1qYGDm1L21N9g6u3xanbMH39TJ8jpbB+P8
MCBebm1UqviCP5lCLW+rYJ+Qw+AmTD+LEy7ZHM8mIxiRzlEdjudWrDKFw87VLeWv
J3MdhDIrY5TCFIJdbuT03v64sAlbsLVfR5jP7orKHXu+X7SMIGLKldDZ9z2lmFcS
STWVeMeqz5u3DCHB65Fz/uSh7bpi7Imv9Q72VQtdPJny0aSnYCOBSHk5PqdcFep+
/REu34v2WBSj8a5OjXbjBR0eQ4EekeT8l1F+hA8crTJPYHkbOe+HX3ZbjoMYkxtK
ERDXcb8O0T96g77dqjrLKanZSam0HGRlAai6M4SH1difd+W9PvRbDyjHiTnrWAPo
f/ZTOYPqWRZS6n/GZuifAefLmr/8NeR7STlFhbGVQHHovyDsh+5zmM7VW5mShIoP
tiAyiwHPXg0iuULmUrgTlllrOxeir7CE5mH18UCLh1/rpHulWtdbezHh1h0GE03T
aur14qV9HJ84RSqizZOdvkRQpy9C4WSod0X0vacHbx7DsRDgCiPe11271J46s8DR
Gx+FCQBK3QFWbpKYEZEDSSk7OOJE8gI6VxQue6Vb9YWinnSpq/661mq8kBR4J5Aw
xivONj8873axWD21ITWBa9CHuujAbt9Fqla2VpyPyVBI9VhTGQVRlHajbVFf6IBj
5yrNKufSxcyrDB1RBOBpLck7vUL7mKH4HvGgEkIzYt9/nKaldBcalI10atGMUOy9
o0DAo6c9c6at3a4EYxKU8oQmRW3KHj6+aFPfZ3eS5QdD4eEW9y6WyfDV1SU/BgIs
BDLvnqY4gN0+JlzxyozU3Y9xD3pQ8SxsiTFfqIybW3PoALTgdiV0xOXN6qCW6Gwc
ZOJOpV8RZ9nhSlGbzHQ+yfWpNuEEx4gfMsxCth8n5d+o3m5HTa+KZOv+1+o0eSHJ
gFeRMyAqXIt9qmoluKaMyH7XPhWSv7oiATrMD1/X2fvzn4MCKy9jwSjVvT7Cu4sL
+IHpM5nRw1FxpAKjiO4GoavdHCuOWzpGheGLSffc5KT3RsxxotrzapxW1kgzHRfV
Rt9i6RlmX4D2QdkiOjirwwDbTEexw/kMJuk+YSEpDwRvmhGKyQn1ARASxCCjambu
EHb8jmei95w7tDG/AiR+7PvM6w4ShQrYOFxTpC7hlYCqfblqET46DqiJ/VzAdJ9O
SCH5sxzrh5y/8sWRdmtvJX6Q8WD0azqKlNXtZmbjIl2WH5IFec9my5VPA2k1kKJH
nZW46CDCZ+4JiKV7bWqhLmk1Scy3EUzC1egPxJ3KwO3zCICx3xnEe9Zn+5Q6B7dq
AJlME29g+/7rTScBJGJXbXSdOVk/ZjqeKhPyYZAHz6FgL/oRVJNX3XYILXRlxOkm
wglgjvbk/mv/M7TR/6VbDNnk0LyiXXsR6F9u8CzbFaLBAaoBzK5N+wOVcg5y9pwV
2Ra3rdUfW8csMHtPOXImF6rdtBb9KCZJB4VTMJXXerkJRYwHH8nAxK2ovQhBu/SE
WuNccHp4IBWVEuH6pt5KLwv4J/8IC85/Y8aqJJNVNjx5c9cuHg2Y4aHKo2vQ9Qnh
4orxUx1+PKlJ81z+7SUAXq68WwTtDJZY8xKYNYIuH2a83/H4qcz70Npn4uhPokru
2ypw34pCsbIZv7SLqXJBb/FslrtKjyWSVJKYsF3GpRUwu3KimNCP/uq5ILwH4tFO
hj21e/su1VOpgwgdG3tRY5C4EZyUzPyGzIlu8QIZASploxenwmzV+97lvNHRe3SM
+MZ87AeQu/8UpMusHLtSII+KphVHEXRRvHBUPmkU03O5PoUkKPkTd9yK45VGrZea
HxUzKR7sFuJQCWKXlFcNu9Uir3iJ5xcNYzfKT62j0JuglfVySfJ5oqoX1V10BlMN
CPjkLisiKQSwEeFn3EhBMOLJ1308Gwi4qGHiQGPE8jUVqkBZ2nw0jK5PmxSYG17/
8uhQGM0fBxcM1yWY/+GkQZsd+NTNzGv3+T+oaVkqgDoYoAsxDf/heeUEF18ikHLy
oVyv5atu0z3iOkRpO/VLiSDGfUtdBbSxCVivd/2rSAW5Kj604ZhLyGYXTmussGhO
vtxobwCIR+Cx+rnKVAgVYgGWFWuuPOUEwZftcSWGf7cBWqdQScmSoUJOn91vs7bq
BJxDdoSv9I/8V/eo2j5XhI/RtxI+GfLO6cYHrkm4Ay1wDZZeOVXRcg61Nt6RDA9d
eUQ3JhhGeIL4btBtRwWS3rGHqzHgnm4QDU+EMHcxueg+tYimEDYrontYdVM60D+N
4botiZRCgnONf+3nq6NIDBFcvhEuJbAaf+6LgWijtO4L2PQfZieqVE6kPCdhR3RN
7pfRvJE0iRQwIIhlPCUR7LS/WM4vgcv3XxjIXAUVau3YSYTZGwZTsnXhTLzY//u/
p2xG3L4FjrPUmK54KMTa4uBqcKooZLZsjezdLbTDMa2uUHL/cpbWnl/Nam11FHTm
P4VGgCWRhvp5DKGy/X7ykjV0UirOvZT0ym6iO6l56Om0icA0e57vOmnhP2aYrWDJ
6nTyXAOFo/Nya5X05cX0FmhI1K+R44xTnA7AD00Mg3k1A1pX0F3dF/GE0zuff9Le
CddKANxbAFJBNHxBp5mA2WErOvqeW+C7cshKY4y8BHDjCQ4zpwz5ewdz2YspOvZE
b2wWB746sWzik4nv8X0yDvbMlpka8Hox2mDJp09SsvGnHui6zkQyt00+cEF+BzX7
IN1eqMg3oLPLm5xqiYZpAQ0MVd7jfIDX2/nj3Q5olLAKt7WJNNBy5yVuHMsd2RpU
AfmcigvokZesaPijPU9DXxSGLdOhnheo9UKZlryVEO8hWkAfIk8CI136kJAqL/xf
XdxeOgIkJoJMF8MwTTBfRHQKBupm6pJzYlMVh+wIs5hfac5MEbse7hC61CRwf/Q6
1awDyq17NfZLz3j6obk7uwhTbOifQfp2RhvZKstXMnVK3AwHiRNK+y+VKro4ikUw
aWcqeXjWC31cCShqEZtWYqgi2tOVw2YWAY2Y5yjBNJ1hseN9+BsZbTaXKt+zg67V
7X8b46ZtjNdeNWvy02brmygfHFdfr8ZdEsaaOjG0V9Zj0Gg72HWdkwrY8jPaKj6N
w4XCeUxxKJmjxzs0a58aR+ATiq0I0PoqVQlOQsLk+j08eInAPe0KqcnDIAdZ9sjx
Guui2DLGjXVAtex/KtGiBwpzbTo9T8LP4kXsxMNQ5FsnJ8JK1PsjjthpdBIv3nTw
gw99cj7MQkPoyvoz98Befu7vuFTutL5fls6dSaqD2XgMnJmLJ3yjYlHpjT4Gx1AK
FYEK/Whj2uPEWMccX3AAmSkLmm55V78t3bY+S4cPS2NtenXViXe9ekNEq8z3rx9R
Q953XM3wXbfJn/9equoRXBid58ifIKhU4c+mlcEY+M690bF6pHN09yjVUiyLJijP
eStCrVCfmySxIvjvG2WTfg34Y5C7ZPu4/kO0lCrK8CbENDEZLI0jp2AXp6Zx2Nv2
vAeBJTExdrIkYKNs4SVCalQpQrfJcNFtksh80+rxETiGFP/3EsUlhYXjJePC8cHO
1vGUqjSi2LczJgeTskzGALR6f8Ig5/TXpJTtIVaMZP+KFEJlnf79PRqaPGzXt0wI
h5V+6GJXiiWjNzPqO7+9hRU5G9SMbMSBHIJNUR4k0Gi9Hph01ljiHWx78a4y3tZ8
/5NOUjh7LIrQ1OmEljHSIaUkpY6t7HKnSpSbCxXNRBOOr9ow0UhHDKpZliJh1tcA
6PgePNYhLtMjeYPpp/7yWnnHQhGSBJc06EfIkhYkAGhZCvMM3iOf8qF2FBH4YM10
0FVK0epuQC1XnPOabSV+q8IXwFPkUvtP9bUis2NSqb9CkrLJaUiEuIE0QPBWfNsO
Gc9tcr//ZWcUjyDd6A+xzYvhFkwIBmUCe2wltikA2jB4KLhiNnK7e0lbwUSL1m0e
fhtUHP/nA7Y2y2MFKN5/b4fr/tyTMjGsJmmXFb65ms+B09Cw1RRmoHDUhrU72OI9
vE1e9Q8qlTjsT1Vhdduu7A9hJENGvBt1wufVV6OxHh3G8vZ1ruEAs+PwhBHR7RLs
qnUqTkC2BBYKKChP1ZFOEPptarkAXJ14LJRG86EFCnL9MKG6Cam0XBDxNsYLfqym
3h/k9ZrsYdxVDauavxX5VI6NwRHLMYuz/7ICBgtHc0f1Flb3iFFhpKaoWCfml+us
TkYkCOX12vdf7t3UkfedTOuq4L4MF4wV60mMpL7zmGwTqD/eb8ck188nC7+76Vn8
pnJUhQiasmf9PusIv3KD3GIoyx4uf9BqjuAH3diqlCoRWpu0a/rJAKYt57JQB73w
+kL89BYamfeIx+909EhmRq6NFbmpLRVbn6otsTMR8P24fQQxqhLa4IPoOdPEzURT
qUj4pdKUETQbjLFdz51LF8zz8MPyWwSnGpc4Z91DjlvElGF2D09pJ293d2AAJ8Db
rteea8b5hwolttJ3lYJ+rzf/NSv6k4V+yd0PJ3Uda299+Wm62ldFTQUH1z6Czrdy
Q1nErjmGpkgRcE/+aJjMAdUVNeTNTf2cXS8wPaUJPvRl23M/SpgPJYJtMCKY8lY8
gzcH/A8xM2ibP1WoMDtxg6pCwSkIYx5R4+3+MNGu8uRHTIO5UOoSAV8FDlCi9HX7
YMdXThv4TN5f2rMm38gzXQFC2oIdj3GMuMX2t75tQgGkOGIYLIBr7twKpFXbFd/i
LrC3jpZWeiVMKwruZO7RXmVDqcvjWPubYGQT8YioIryEsDiYq2gGagJOyHBmYTW+
9PqJ8oU90mVeJnNIJisYKwz6qerA0Jpo8AipC3FLj1HJQTi1O6k8gYZnhH55S2vl
TNoXD2EUDbMXO+KqeJZxsX/cuqlP3Kui653jVV4VMgEUwy4XwCCaSXiAeQJcmHfw
08CmNYT5Ly4+9Bjezl9reTOHPf2C3Gt4Ijx+WIaXogTpbiFhmX2kFiu4OVhZfNgv
eGTDtK6qAg86upkLUmOylSN4BrTvJUgEdez5yMjTDDcQRObCnM8dcMhL0hQ7CiPm
NNGFWQEvDeIYrqiVDWCmoQPMHAlWdcXF0iRZez2Q/0DgbfQLHvKwZNlBWMyaQF+C
JRsLwQmrMjF0ftv6SQxl8ZNfLPcQX4IobeP1Y6DGNXH6uWCfgFjjNYunGtxFO9NY
V9McpekPqPteDH6rnk/UsCJDqPTn342SGV/3ZQYNGrUNBX2CTxTKyDjiNhxnw2MC
D2X/cRkwkB1i87lYebDNLZ5tpndpPYKyQMmQjP3ETwjxMF2YNZEBz8ucMjKkqSsa
8C4FFp3Jq9QD/YLUBznss/G1tAcngnlYWLD1eRJd9czxHDm908z3FBvAIfMDfSjO
WulicuaeVz8AbO/bORH4S5pN05niwrMsvdZ/4397jyY0bmTlHV7bn00LL2no+kBB
+2L8LmKcBuWX6an9lFl/tvcyuzxUrSLgEKGCqaOda5RQrZUYE50D7Uc2oNaigcr0
zxVzvsHbP0OYsnHimb1Y63RtlesJufMAdPlGXRuqe9pAx7CB2VT1HMA1J3leCGYv
51aJUlmhFP1Uc97BYg+TUHkVRmJHINGTQdESVKMjcMFmBSZCB8G1qIGZBrfJ5FUw
SF1HycNF1yxnhu5kWpN59Lrl1Vk9U6YJmY+dpUbjqIOTiU0QYCaMQyJ+qhcxPZy4
gqRsP6vdJoxWF1nqrugQMZc278+mEu8Cj/JxzHtd0iPEcP/oecBlW1ru4y/nMhZC
oyI7qkytHnr2lAEPBjWwM6lg54uFV1KfA5W6DJ1HkQm+PZN7ObYhKXJlm+RXua0t
5kns5Meo0HqG2c/gF/0mPoVgWL/AIJpYfK9JnyTBt4pLtEOkG9FPq7qJ7GyF9939
L1PEyZLXtr166fu2xWWYTU8lwRKJWr4Ic7axrwAXxPfrAW4IU/Ic3xOwWCJo+9IS
swtUzL1KjaaheZgMPDdH1sFiTdORKkBBGIs+q7JEDv1pKM7+nyA6K8AO344gMcdQ
N4cGAWzDwUz8yfHYf0lLC8U2NNjFhPaESUTE3osa6R6Ti/LVKDp/8312Z828a6qJ
JDMYaCV9hap37zlN9dyVuSTJurEciwZKADi22BJdSbG5R/LIcuMTq+TPYiXprAvK
n/YcoRwnphfm1d8GRS4AS10OTGmCn+cg/E7Jf66MHYaKTS3fcNkpJ3dEqrz7iunv
pBTHZZspR0ILwr6ceBhiCBgc1jtBbRXUBR2Q5DrpBX3WiMamCQ0+7dlIK9IvwrI8
ep9vB14g3VtQ9ClL1PIJtu4Wy06tSgaMZrb/3v3ZGBH68JBEdCBmCwHAlYouvOqB
CB2tprRvuUOVfUZkhnmaq4f/mDIAaPDUK01Mn0JLmZvZ5ovsDdf65Fm9Pjd+AuKp
SqGSRklqdsMx7mhzAXdtB5hnD6J0lvey90G4vj9ejA/utCm0dqk1hmLmgmUukvB5
3uk3pIQ9gH13xOXGdAPJOvWfeglx0t1+48Fag3xHRg0fpNDtDQRXnKQLWduW/QPy
u0ob3+4kuFK4FoxYZt+IcVLjhT8euARHHC7MbkLkfHGHPbm26Sv09c8vk9W779mU
3vDmpHruARAnvCwYaq27y1ljmGVrmdO0k5kehuE9xfkqQ7ABxdCiAnsYqDu+W5dN
s9g0rxbp949ioisKb5raDxkDhy5dJSMnePDDBXVjf4fpsHqGxXCSoWkwiGgixK7V
q/eO7F1Fo68keHsNUkYpMy35x9zapQ7XOpjGfyfuwTJX67Tjj5qKSyrM22HvWw8L
qAbHmK36HxD1wTt+9vyGOfSURcRXxkC5C8jh/5+8Q70KZ6YWElMPyQzGH0R1yx/z
Eu116/vtE0KG6ZJqDVt51wSNW2IteF27HyXeVS/3MzrtBj77wPFxpgqAq4e4WRoF
yG3SWYeDtpua5MSi8pJUee/N3TGxuwq0AJQUVV/C0naxGBFHP/i3UgCKWdYpxTvd
uOXVanmKYN7rnLkje+Eknyy4p+qArni9ppIXmzYN++6F5D/vQ5RfqRrddm7IFnYB
fqzpb6ORXZlsnzJxObGDc6p+53qQgGW69iThOIUtpmszfMrcSWbBwSxlcEhyb993
e9hvw5qdmWaF7bAZ9F56b+4Pdcjm54yZzF4simMaGg5tlCjqqeLIY7XId/MendcH
SkBaSrKp43+DNedcmTgzfv93hqqrDV7mn94DvdmteMkWDrLO3XJ10wKD5elSVbaf
5KjO9dEpcC5SqEYgIQOSJgaWRu6ZCd9gDv90biQRd5My0DMP8LEfMzyynkcdpDPE
yBV81jwPdfuB5hwZ0nSE3rzf55iz2CrdJrffL752uGMHvzU3UtNHazCzGbCFFZQV
1dGAQ4Mt+ytQy9tiJSg+/Rxq7g12X/UbkXa7qx/3LLsNYkLG0/V/nEhr+peu7dAz
c+ajEm97WHQlYpW9ONU+CGKQZuHuGiUNg/76s0gKRyBphby3Qg+TyYYX5fmzOpqT
bd6YzEYXUodp7H+ZROU8Q8GEDIVTRiJi+Ycpn693qw7nUbtKq9nR2TMhUX9kaCsd
H8cm1n+IhyZv5C4OGzQ/cbQynU9KsZBSxfswUUxmfS+mxm81lbn2HBB1bAE5nGmJ
LM3XyWH3PvcBVjHlze/mH6aNNUudlH5sG9ySyaO5OpT9KifQpU7q6hyqIToA2sDD
Ye+n4TKJWhu7FJ+0Gc9wY/7MiFcd6O6QuOMHwI/Q1M5XbzxTZ9p4fEurJJa4UIhi
3xAz+Iof1tHB0yxUK3rSehyrHmVuuxS9vKgD+P7lK1mgY0Vk7gLLCk07ux0fvukU
HAa6UQQEDsJH5PDIxmDdI6TiNnANPSaWGkkWz9pGykzQC5bs+QwhU5kxsXVeKRvK
y4K4dXehGzx2ATZJPFEMkcfSCTsWM2ToPMKBcziCWnXhoI42ZX6sA1GIdIC0A2cr
lXJwwTDi9KMAPnIo0FHo2N2CaMcCWqvhAATNeNKoYVu+vWeofC7IzadFcu90hIpy
ZEgEy0wzr9txSeHviF42GB8otfFcQXdh7h2H/ZZDewXbNq+TNVmsQckG9/EHshDb
qRGFGZwH4FLnJm4uPKSRO1Hn4M7FbI38aLLbPJ6b6CEkQeWb3VfDwljJ406vtxoY
IllIqZfSa81nv4K7XDnQywlNc9riJAZ5NUpCtaRGQvLE9rnpSXmyCfP2sntvkryu
9uPX/jNuc7VdtFSMPNpxlDthR7dMvZAkIejcYWpBtueB19YeHF2RHw61AtS5QxP2
fgQZrAxca/zF9t5eza7N1C2UOES8rUI9IJ19+bZExwQLCqaOvz1eULeSI/bsqbTM
mA2tjztRnOjO7Fq1xc0ZWFLbjcwKDz/wixF2lkMd1mzgtJCfCYP3eL5tUqwMdbL8
+NvaW11qZ6A2BVs61sV294AuOKMIf0anx7HIRcVvFBHBGgC1xIPep5XTk4M+9Kc5
tIvctbv41XlcEBswpFurEbUsOC5FjYFCeC+diqIKKjJCL37JDFoyzNmQwYbELVv3
KxV9FgvIy2D5pOGoKaVdIn6s8Kb5NAzwRRHeUVosKL42uTWpglo1UTk1Z/AmUu8j
n7O9jaErSUGj6I/c+40e7yoqCOMvHsTJwXAcQsAZzoLGpTJ7uLyQnXS3pkdvxBFZ
E9GQ0L2HQIgxSBIK6BtoGR83OooyoYSn/L4yJzEhWREYkQIJJz5Rm911g+oXjmE7
KGnY1xeOtL9KJlNuy0lQwVoqnQMwaKbjH2a58AtTqdRDL07jiZpRNRtJPcklLKQ0
Q1NZCfeBXCfjigoGlIl4fihCS98hwKjEMglYe6ENVu2gl16ymIJQ22E9EOw6Z1eV
ImvU3aVxW+68pnn0B5uULEbc0yNzBjOIWReYMoNsa1C2X6o8y7aZ22vSemUrZClD
rDCytRQ6exxFhJ0tOFZz0nNwTHvRky4vzWENZraKbuBoLvsrpUCmhUc5FuXMI7id
o++guaopl+x2X6bp6SDLj3Dl3vNt2u9cU2m4kqHBkOlwJ3MVeQoyLDLw9ksTbACz
pHjNa7oEgDjUWQwRZCZjiQDkOu59hzMAFIDzzgeiswp7upCHDSoyZK5XZuK9Hs2x
AyMDTgtGhgIJFk34OpVY8jBNlLF6Sf6foeY7mOYW17jkZuhOmOHiB6chBCo5+Mec
IQ6oTuAXt+KyLbr0Bncq/hDOLIaCx1oB+S73CACl+sQ2eGUxN8einhumI9d3A/Dc
aM/7PQaHgsMXMb3BxMBxQV6pSJUZd09V0rGsD9GMqvtsVWz3luLPrkVXngUVcZx7
tNi70ztqGQEKQSX7cqHlWyKAxI7xVXqS5dyGoxhVqBpSPkA1apusm94phHzeYI1B
a+o4Ozfz05VEnPQVGBQVgc4Rz5Vt91h9EE3M8q/ZwUllGwoDHX/ltO3psv8nFwnh
0CXo+h9fx3NW/PSr0BYjd9QbircjCGMEY0XEnjtVH/ICsessBhzOrLwkfLbiTaW8
L1wjUIaebrvtZ8YpRd5+GrAWzeWl1Sv+Cmx1+NY7saXx5ylOxGBtxURRMXrRMQd4
4opGNj+CpsNMylZ/IIN8u42/UzJYYnoFW2y5fLTENBxMl84YhsFkj8gI3cq33Bxi
urmWfKIupAYI0Qsf0P8YoiaQdGL4J9hMa2BktBaqCYdh8bmAHEzf1p4hJIbaKx61
82bcghd2BR2dqvLQJh/OGVGsnVBRXoGild8ZhAWgWStbO9eWWFwMyIK3qRSB4/QN
4QUeIp+ArWqDPsZs8WNPggDDjaobK4oPkJn/cwXxdBMYEjFXb+uvO2/iN1gESaiD
U9g57nSNzyThKyIYiyIBJ/Sls4V+bf++GKvPSxxGcZkVjC3tsD+VKbBDDev3ECl4
VMKF5AaiQwAIHKvJNVhCyq8uw/gVwY+oVHi5RjxqkELOdzelRKYwneZTGrdJmyeP
bIiXjn3SrKhzCZDRgJszr+p6MPLBzPko/BVGhcMhUCHD2y3ugj4mGZVPcuhFSvzn
BbbD2g6OEXHV0NvCEzo8exzRKktrPWM7htV452XtlPKbWOyPGUXSXLus4iJHf1In
xsmXGZCgu71iIyAQuZ7l7RSO42fxNy3i9/6MHEGCzcuBq9huH7jhzexh45Nz7Igu
i0Q2P8uCqRVLtvaCJYcb1fXXk0pyK24/LCVcdFUVN7oivhmvVYjI7s3nLOairyCh
G84D3yicGd6fx1AyDLLt2tZAjE4UvGBinVuOW9fTRgYaD6JDRNH4L+ke978pEGL1
rnu3FGUw6+OlGpFqAhRg2JOVClf65Gvpye0aArJHgTJVJUIC1katBDUrVYALhnEt
fVDg655rKUwNk7lMIpTPE8TrCBM0bOeqZXrWzdb6StE34+p2Yy+b3pZmXmgiHHkE
tfUI1Bd6VJZyDWvrVLqpVn7X/eFxv5Xd9uehExmlRwBWJ+mbW6s/UqKVsOhpY0Wi
Q1vvJKzf+T8VTJuLEcN8XC52vOXBQud55Z3hVOq+xBAXjcMItChFD1l9AraL/+IR
17/hgM/acklQXjQhE8dW2il9um96qBoehlgFaln00f1iRPl6RceboCjOw91xKS69
tBcjS9D9O8scEF5ca62CBg2R22agtFQFMRmZeLb8++Jn5mBxFfy8B+tVjKQz1ZsR
wnMj/wD5jI0WcXN55MrdzIF76p2s1pwfCVUyjRq9ODoiFNGoUaEGCWWYeetjvGYK
yPis5/bdjkUbj1xZCxMKGn13HtQMudQ8/9k7yfQ9FwCdu0VuYMPO0kqOgxZGXQpu
+4MTI2MMN6yDnnQC2lBiNjosjwJp9sf1agX61wLB5iF6GvghMxD8xY1vSGZaJTuX
bmwbrMD0ahK3z/Y6vPkVv7b0ykFDgwjN8CD/YI/+793q478vxJoPHreokGci/J0u
H3tjRxKRbH2fdo94NlBlxb24o86Hc+s3YOHQeYlicHxYVc+pZqjTlFTIUcq2l+xf
xSwNtnKy0HQ4QZtTNCyz8499uYw8twVlmO6KysCSoY0tfEm3hzFGxqfr48TzPFTw
ed1q9fyWo0RVPQwB/2RplDfTbnRtYWd2O/39D03VTGY7nDzNma5Lfb0ur4L/99Yn
RoCL+6tYihs3BNWqhMhEe5wcF5SQzDQfg7MtjDEPXcOYJ1szXzZGddnoZqtesr3u
O74YLi0pfT72KOP4/tcnKYWJe9yqS9fUjZ65srmkq5R/9kvT9T5UiMHph/s5mIeK
1jAMVfJjeqVkxLokIZGO5w/ecf6B41OYrP6nk+CaLQPcmTJsXcz3c0qGRwsypCzM
x3t2twVGEcFjT6Q65XtBzULBt998ojmn87RuahJ+4yvPGeqgDrmen12tNnBpoiDG
HrzWRMCwtRIx5lUC6oup4fuffjFTZCugkyLxCDwG4cYGy/J7UeasgL740y3Lq9bJ
Jz4Nyi+dQae7WSMfOBVKCcK643D+iVxTWNA8MrW7S5lPIN0NtooAu7v28lOQU5zT
RMu6S4yZBf9G96qJsXx+ACy4vlel1rOtyMjfFst2M6kryz9XSE2zGJuFAedi3vaZ
yKgFhzksGXBVdYZBymZUDcHTxIP8qNys8xa8JrXVgb7yyxQEtAXgeVjAwOChsmcJ
6fM2VsL0smPFmRYDV4HIq9vpI4vl+wSst2PwBchyeD5PWUwTA+TyJ6qf1g2VWsEq
602sQmsZ1AkEw+1/SmTpTH8OppZk6NBjVHO3iWOk+nNYkqgAnrkzvskqAYfzfMgK
qSBBxKGEu64H8EfX5/AUc3Pt4H+8ZQRoROvn7aWOmhDagaunFxjFcKoe9E5oCWTC
ivqTn4VgGYfKGmdYBTD6aW28AC72spPKRNq+DeJ+n+v/N6wCXAPB2Fyp9ILs5Q8j
7evYxxiB3uP4bFl75/rcUZssnaGOLMte3nAjZ72QwiCfHt7LwbhGikyhr5ffgI+H
Yf64lmAbkgCxWnMiipej2OFVk65wl/52csrpcgW2frqLEYWawm37tdcpmbnWAP8+
ZKPwxe968Gmlo0+3ZO4UnmqobEnrXyxh0T2Dgryio6XqbAgxqpP4DGe3L8/K65AE
8o6s9eBf0lBinJ/MaQdYTwXLDxXlhYSIC7kyym3ag5nAenj6N++pDn3GrxOT15fZ
uzdZEayRylALuWiUv7V99e8tVqeFnTav5KMOaAFn8Z9AnScCcR4+NXPLwB6prkMH
FiLEfl92D5vnAMsAyN5WFc75NTcbVjo5Ao84YTeqzRKk2pRDrHvf3qckv6iBw57G
4Qe8t5zXbvoE/CFy3KL6MzMKeysYZ2YCZtN1FvxiZxwYSlqy9qfJle/QKO7EONXx
D3D/FxvBCkSe4FcsaZi4MsRR+eAPNrC/NKs6kkIUUBI/U0h3NZc99lypScD8f3bO
og5LQUFMWNaLZyF0tNOBj23S1X4Enmw8f+f0NJ2f2Yog1mxbM+r1FztYwNtFyX55
J3V2ZnEEUaKg/DEEs72BJjs2beFsGJ8H4OzNT7uyiii4eKURPq/Hbdc+QQ/V1oku
nQZQEUqjjzNk740sfXviT8uCotIzKQtegpWF7v3FPttaX8R4e2Azec+GWY8CEDS5
j4D7bFE6UvGShR203LZAaRoHEG0QQaO+lWFSNnKXjFyN2kC1rYLJ/atCKltQOMvQ
F6FdFO+VPUlPf8N3U7L8sCvK4YtqEGRz3+vYQjuP8rPBNFloPsDVF2gtGMKUccIy
brdZr5nrvQhlzFiAdrfPVwbjc61HMBQMVMV1Wvhxujbqy8yu2FZn48O8i9Zp4FT1
gio1QpBgscTviMueIYyiMtF339qx3DqbjcZdX4ssxDUue8B0CxCpdXfA7L6hcLoD
NHwcxdBnJ3OlxuiRH4/Kj09i0BKOWFl6Ssw+dtnuAP5OmJXxftsiArLW2Z3qt+E1
YnCBXxePOvaZX2bPc/1fWgIl/OoyBiEWDoPrKaYJ2vL/sr9oCx5AKVtlnl/wT3CB
21wUtvVMzy8ul/q22554I38ZlbROpZCYl0t/fXRLvTnKU98F9ITkpniYwAnY6XNc
SPh9YfwtVrjiuO1zFH0JeSC41gCEXgUMH5PUXvPCOHIUAdg28JpZsD+FZ48v59wy
IL0jfiBCGarHejQY4y6PSqDt4KM1/OeB0gB7OFmdNbRv3iGf/biMq0BKq0jB17+q
EeA5+vPkAX8MpVeJlJfH5BFI8XkEysXY8GO2EP4I088eDASvEwFFMTLq//XqGexk
2xqED4okE2bRUjw6xMxDNettpLQVVHBAYu35cIZeLrZJa6/LcPMijx4KJn3z7kBR
Zw2vvbpeca4dM6epbqlT/3t9NToEgIhqhNLUYfrAnTYUpuTCtieHUhvKQZ85J83K
dv7ZzhOf51duIc04UGGqTmsF5Vd1DlVWSRN1M9+okf+NyhxDe/2tc1pWpFkQgksi
AyfCZ1nijEPyLvO2VrwvtEO1PzHgU5WN2u+3D37IvGXlUcBgGc4FTQ4cQYwdyZNj
9/ZJiP1d/C001IjYL/9JMxGf3VVJmpWxrmIWu1M9UCkTyC6bLl7BkUVPIrtlcf+R
rilT6RLAcXh7Zbw2y0i0zmrJXEpUCsNx8iCJ9a+IoFuFe7WAU4qpGGyHAx6lxvJW
Y2U1gfqlUWWiZlC5MdfmGhqzd4kHo/uSkBPql61o/0c5iWDvIDkSzT+lpoWXh9C0
WpOudwaSARDN0LQ1/ZUqp6NXPZleYVFbjKxdksJDbLrgdcpi69JokH8WWMWV/gqD
gFmNj/UGo2a54nbxDsQ534+Bc3rFmqSNtzSsUy0uxRE3WrbYPRE+iobqDxfoX+1e
6n8YcUnn4aO8oj+ZD9iO2aqqpEGo0I1PY9kb5ar4WYmlcX5BeekHWhlsGhHPh2aQ
3Aa5fto1+d620VsqjlOXiJpP98q+x0ox+mJv1RtOM82L39n+Po2FaBgnQsUGo5PO
OO+s7TKcV7pH+Nmt26rVGJ7x/uPr9xn7bAgifgK/BSTbkLtWpsT2hHxBH+FjPvwP
NsbCxVQ7k4vHyrlgHqc/VqlCVgRvbZue46yomVCz1NZupk+Hu9uw9xj9oT9k4ECV
+F34hYl2hkacFBazpWiPrkUFe7/ZMMK+LcD29uI/SwOVv8/AsfCOAW4adev//LjX
RaLV7W8nnQQDkhl6PY/LDu9xVQL9NnuKZ6wX2EhA3yaHAjwUOkWCsJUuyMjzY9Ez
q9L+ufakW7/WUSBZHYUTXAyMknjAfn4sfGUff2LUyaV291lU6p7q5V2YNh0fWhtH
a0d8NNLnbieEy0zEO66KdZ1aWrhQ8uTCwYZYGVwOJOciAfPK2ZRA6Ip03Y5NBAz6
zu1MjNEhc6NIQ9EkGYfj6yQmF0qIiMH0ezWQYyZCR60N3OwjTy9l4t1EJE7treOJ
1Xbk87yDF5R6qom4rZO8E+Tv5vPUMKmUr1tJRM7tkPjqHzYWkoo7xQQ4nKA7uut/
Ei3B/4xCYmxFlEFwq7lZJ4exQgF4pGE4wMDjAxmnz1KtLwY96mZnmbvnnNylIBP2
dTVlQ+oDJ3AZ070CQDxW9dCTc0whTYdPJmhIsJXKSNxPz2Z4b5NicLYaL4RYs19I
oHZtEZpxGaHIUXX14Lx3Is7a3NyZLVW0KuBubiXRCiLJt5FuKRqz1xKz+lyXg9ks
hbZ2hx8UperoDnRrt2HnEsRkm9PY+lHOIj4eFVXJ7ZqUUSPJiO/GFV2JT8/IgO+q
ApoBpftie82ezuX6mN9H4clH/xLcZ/UbBYeKMgMJbNY+BCDNCYGKTp4WhdVPuU1C
mqBP2SnTbqOUWJdcZl60IpVxEyk3A7rSGj0kirA4TDpMWDnh/Gx5671P2HyA0VxY
3MhZgg4egP1ZWyNTxdvF/TCp4hhKyIpyUp2QfTVydnGUoDv0OwfPIqIqWDD7epsJ
JCQHXOoSWZ9QG/IU86bKK6GnDvrO8MqiORqCEJyNJMiDxSQQVwCxZ9fHQdl0AtEF
vm44/W2VbalLK8lykjFg2I8V4qEfBtciaOggmoNmdZ7pruLzHUHwSvaSW+N5GIvn
Wv5g7lsWqAhmUm+wI6CCEFdlt9xopW1AhH1BDHrBSzTYJru807XufL+9K8CpU9le
DPJGYHDSlNiwF3GrMizGgDdf7hDEEvAlWxroyUixNJeiGFRWFJxzUD6M6tNdaHPX
chjK0rJDJTEI7NxuQp1lCvOPkXJ2UkpVOvNQz1myaV9CpJ8gGF6GRYbGCLWml5i0
WaQSe3ZJcp01UEhBKebJp1yW8ilLpooawdcm0IezF+SI3UM6iCvRCoAL/BjfsqKz
cUmA4Je4h/b+IPv2IbmmIFkdDRyNKOsCmFCNFXCafSTukJF62UM8vX1DM7POBvZ2
KsHofiflnNxE30aQIltTq+lKtgaP58QumIYfNc0BkxxqqtFTRDmxZFotetBLVBGi
xcjFxAyDD5XWmyI8lux+tCLFMzT//6k6D7EmbLI5e3pGXylc+8tI0MgrFf7hMBBU
X6+ream2vox5i7NgID9s+J82CO1QNvD+wvHelB9iyPpSEGgP6p8zF8E0mm6mVMBW
hVi9ZaMdCVIcM0vFuul5oALVOsik9T1SqjTtiMhBmDUm/nptGj4G5ACWZIpOFmj1
EO2iY2mcvOle1Ie+t8sZTM3hTl9gMNLvkso6CYVbmsm76/RKVe7H3zbClbEbpdWE
IFRq6zM1rb3zi1drDOT/9Ft2T7g74zaJxRdmxEgP7xGL7+zLwpMNdMo3gfZW0EtE
/39ET8GlWQiXfjDdfX7B3eCTNc2G9h1Gi4Qy36l8FHf1VyfKJL51T83/fxVUbqtc
0c18s7itaz5sdFsld/mqSm89TsrAIT4ucYOPTgApW/FErq+pN7l2ZdcgZsrL5kK2
kSKfCVDzLgaOWetQKFiQVVarzj9GkiFDJp+Ez/uGuk7gVW0BTUo1hJrY0iFNNRpz
hmhT6DIB4WiZ31O5CH7aRjsB89Ft3a4q6lhPruE/QfMcKhhpJpWaopvZ8n+WaJy/
0gr8W1aSsCRQ4j540Y3L+niMYIQfEbqfYDUSPhgak4Rp96HfgabIsCPaokOH5FaO
24LGyC21TZScElEWK4qmPEeANGyW0Lgbvsp/daF0iez88FFZTW61ps4p44EHR9NT
r3Cpa9ijvbVNPKql60/rn8MFntZy4u4NePrdQbolnHSDlLQpwWfpnU7PekFAiTPA
gPgrpzPefsNF6xfgP94zAoZAIn9uza07yWmeflIMTMSM3nQj2SFb36T+kJPxMYpT
qOwaf58H+meFh9XVxbAAtpRpx64PsuxQvAXJUTrN6GzYHhCIrok7wlNpTiwvFDOu
InzMfhApQXiVzyzCeao1uZz5kSHzjRsO/Fq0bQYN3VK2OJEKLgCETQ/bwlgPk8/v
4ChHJ6tCVbUZ7bC4D9R1XK1HHj9I41cKOZKMb2E+CgrkT2O3P+v8bwJfzS2jzmB4
Dhp1tyXoHbow64g/vna4x3STAz/mLkbDKZXJLHZwNhrdyqe54ucqVf6dum0IMLCe
QozDlvvKdMswNHWPIrFnPmXtSAXlxb8VwTbSCF1Gan+B94gK3XrbrcRXYOlPrLhe
wr+paHtSBBH5nN59cds8tZTNlyZvLLbJOYO5RDA8gND1dyg+tvJ3HL5gBFFS1uLk
aU1zeMtnyVM/UxJdMsgA+f0Mns9i//fCKLVbC0JpUMF3vghY2Jlk+Hm4VA+4aue5
/SBJNiWxG6K44u5cy3NifGOqYB8E0XDQVs5mFxqSYQNy3bRUHPyy+KeVK4m5KRrc
AqB+vwUZJbLhojGUsZZcYAkjtqo3A8KBgTyEiOp+YNR48b2FtE5jamZY++cy5g09
2H8gc3+cfxZ5EgIJr5mYVAb5l1BpPZuFYyJhuDao8A7OpNTGBeQtT7tMfuVp6xSQ
u8wBptKBxGHuqaalpmmsVwHy4Wf9AQpxhnymi8R3V2A84xSCNEeBXPWRtABJJmsq
68vz4QRIpZzVAsad/wrN7jpms7OfD4fcUNfYYRDU7zHR/mDoa1nlq/7Lh7zwKD2x
5cOQR5YC4eefZJKov9x5pm6C758NdI+xOV2U2LgQUGucpnwyWgYBNK8livup774p
w/f4REhhdRYyATNZZPeHDzy/Pi6yD/5jFIAiWSI0syyGXFFCBcF2M8HDbtkW+s9i
JMwmIhcE9oiWPMLYegSpXkQ2MO96gsh0cSrpsLgh65PxhNr29kOObbuSmovZTkmg
gV5aO15mcBMktWuIH6XPgExnSJti3oL2BJrdFtsDFt3JNQm/vY3+A9G9klHh1AbH
T3pMYnHGxHre2CaX73oj8rRJQ9xVbv9igC5/5qG8JsXZwXgnK58/TPvp6BcR8yqy
Gkm8s3xFhZUk3fBxM2QRSN3FWNvvQi7qecbtzuiXHAw0zlGI0+LnKpk5RlDT4Uzv
e3kzPLb9xcO2cxkumwySglhMyaa1X2b1RbaDz4S5cMb2pKdmaAe9CD4UxSJFFFx+
pChEuyM9Lp6oVGEP1AMRKSR+Qls6yKCjhFzs5Ag/vnN9n08IhMqZMwPWUEMCeHGR
KzWAK6k8IF0PyQPJeSUbpjdLTaxnA3vb900EAnHK7iKBI6NTIK3EdTAXBkGTZHHb
lxG+yFaYOdkr8GRCV6kSIxZXfnlALXsnkwS8SxsIVIPHvdxVZ8DwxMDimoQ+avV9
qcsmJnrncdKqf9z2qdDHN7DoXpvNipDeOkvugtMKEmmnGs18KK2DW50eiNQzSJga
Htr00gPMn04flGHx0YYiZgOsRNPpMX9hXa08nvpXN3lhsoPFkZpnns8HBwFg4XYP
MFXZ1jb7GaKS9R7NBrDo4Ipkix5MJvZhWNcn+MRBKVHR2hJocIK7OcfjMJNBOZri
LUR0kIly1QRK1xyAEgRoBGWsWYNHrZ5XDSU0VQs0KvfVCw9d1yFrmrqCS9MBrc/6
dxx428DL/M/Jx4LiScsiNBToFWn1YmDcuAd39XYqiobMofF+KejZBmX2QDRgjdUf
h33+zahI5d6sSLTw4Ql0+HexymwD4uDf70Zi/htvsB5Hda018cTpTy4/Evg+XgYO
Ngj+CMVkJONNPucbX8z7rYMwbvZRfAOOy3F6YBkvUZ72Dh2dRTu3DIi9pDIAl7zK
a4qtzQLYlZDAZoy+7kSkFo0XKXwXfZPj8WFBNUuqillgKW/b77RammMo24m7CZVB
lR8K0Uu62QL+IA1Rvptg+M7dWkt+oHDWTqPKEtSoXZ+6k9SPs5kmTOWYlByHoMPf
TxXP6Tk54dU73zPDUXJJPNYXVo6pIh3isXfydLp/lXhtK85Zrxp9f68jHeiaS7ZX
Ca6fuEQJ2RVLDa3mouPRjpOnRyHsRGhm+T2gQxNfzcJOlbYpBUguqoAK89BCsgZ5
I9COkmPG3fC3tOQnTFGBShbPZuDfDvJlht9l0+7vogcqK17S1QfUFWM3D8cdl1t1
nKBtP9y4xqh7JCD3w6yVk0C2nc6U7LuqoRDRfgQ00iaW0FyUcKeGFnNuX5JHQwcG
aAHQKfTP61DT3cDFP4Ak53hNNl9fGsgE+Y5z3uYaiVqvnH676ry3PJVmkaC0oDw2
uK+hhJ2L4ECJHffr0GHC86L9jKdlKKMx1oIqYLBIbm5CwUnsMr17pf4kVAboE1FD
ul9qR9/JZLZpieNHvBTUSZqkFrUZUp41Hh4ZEmfB4VpW3z8kkqBPZNaKeMhl8t4L
J8Zo8fjk4potMnLkP9G7lWbLGnSB8zh2KC8yAAOrPQx+c9ZH0a3qKGlzB5gxM6hX
fcCfMXmaIslffMcMFENq3zJNCdc35aBZICLWdD3nJ9KJUFdgPiYteZS0qr8DuQe3
f7G8Sua+sI35qWMK4owI2IFNcNuzfXrl/YZ6mveGi9x9nm2hLGzQWf+pTbEnjicv
DlWfmf9LRxuBLnmbgo5zf8AIMIRiXF/1AEffgCOC6iuvWWs3A5bS6KtldD5kea0q
p0DRP1kZ+yNy0d5s8XT8P0KFQT4Sc6LFbWLVbX+8caz5Phy6PANTavfmqKN7T4ks
GbZnP55rn5K2HLHoiTiwdFTPSi0qxYrMYNqex7PPHXkv1hScSg89X50+Cke+S6Vb
zJ5u55t2CR+7RVmsnMIVa1U11eES1oEbojZqPoCzZ9QESHTmg2uoSIfZt7b8IxvM
5eEWx10G6rRn+W0m/Gj+jKWCd5n3jlNleukCflZ27ysnoESC99G+HtKbKNPwQaMQ
fPv8Sp02XUA5FYqwWzh/+ZVYZxVDxEhUYHqglVe+acm48PkWuHj/7m+rxW0iaNaU
NgrxG6L+IZYyk4Qy+YoH8wdMoaYBV6C0qcDDZUfY+f8KywIr+3nsSU4wccL8MIgn
7ZYzHGsyP5ASXSXzCgzY0e21OVv+NslXe3+qJ0Y806+x4CLBMMFN1EQmfnbT/8Yc
VrqD9RVR7wSoibkFe4RMPvT2QZDL2ns1vsidYWWLdguNSCGwxh0sqoOnwm4epEp7
95kV4xrFz60vvsYsS1/Mq0JIAGxuLamlPxOEtQkGWiPxH5eSZhSnVviEh5KATKN9
gg+sF2vcXbPAGDy0vUQc5etlvhVhYM/Gr7AuI8DcRSEeNDJRKxY+0+Sic2fSsFIo
NI+4ZvVLsLrGjYHNZtt7BY7TfXW7yQsrT6/lZtNbZwWQtOJskzrYydtF3idGgcbf
921gk5ygYY2uoYx1AXXuOL3RuRcauotdb2XMe3Y8SS+S+v8Diu+NeBTjoPTf6G2F
PYx1/8t5i6kGv7M2hjQ04kZyRJcGMjEDRTwxB3nLx5HK9KNANffS9jI2fmRpllfA
kgBP+/YHfo2Kb9h4bOb52SwNr7GYJwmphFXVzU9nfeYpoIGSUe1ZuNlvlYMGCaMV
TX9BRqM94X3zh4lLPWY7Y0BZ+jlyZjjLpbEXQmvetp7HTbKc9M/cpjmP+rfoRf6C
YB9WVRAjCCwEv5DR5dwkUQZaU8BgBdHxSky/aoo+EsM9WdgE78Mj8DWX5K/rPXBJ
GB9P2csZLI4lGRIGt6Z/uLMXA8mIrHUMRGav7SU2lPC9v9Q8B4MBY0X6HSpaA6oN
rjd8m6cgt3Y6RAZOyj492RMQs4g1CxHb3ZIdyz/J1Sy067aBvPAadYZLufBNyScU
FRh5OzvFW4WgxR6OC0Ko5FwFs2hmLRkzIze8IiO5jA+1QJN1bxSZR6lFowrHRmbe
x9K3FUGX4C9sm5N8YiVhe7wvWY94t+tN+3V7UpYQqU333ispp4K6AwGHIj6DW1gd
be0wvLj8H18yQj+75txhcownbEnqjHVjRx+v4mN7oSYb41kXhaPb7qwzNxQBx+aZ
g9vh2N7oyny4A5fJ6OHBlR7cEQEf+e4NvQeDHe30op/fC2lC25M5DYS1kDFYmGmr
BYlzPJ9R4BFabYeC//VrBLy0pVHdBEAhz0841r1BrqFtm76bRuSZu8J+9z11Fi+K
CjpqQMZ9Ce2GRfytbnFmxSVE/5oiPQ6Bu4HFwRPompCN+JeIL4WHZ4DwVXxXSAUG
YQiZDzkTye7n2V+Ix9bWffhhl6fedVw0SAMNGk7xxp4LLzFlws+WX2V66Xt/KWFy
NGDKalAS7KK1gZFABpuC2Q1kGCCSB9YY0pol73xYBeZJu4W7u2aiJEOp9F+5dttU
g/RfXoTF9sIk+Nf7MWN5Jbob3Gfd1Iu7dyBjMDdnWZudvM763uT/bFICez57kfbj
ZCdRWCs4Zwa2eDmxhADYkVyoDQjgzffdMMwZSv4T0JpwfgK/0VNB55qFXFqX6L+3
yUio5v2dPCwMezuMylDIL7+SpXV0W35E2ovYsUu/S5RtGApzUULauPlATNZK2/xE
N3sEbHP/Jw32ZzeyJlopWiQkaCMyd50wh9zF+hDeETxEz79110bqO8Ju51U80QTc
7Aor+KJMMHbgVms+EVV0yTNUDDNtRJbBv7CnjNhcT470eGXItrxj5e5O+muddDos
FRsmMmVWqaiE6qLw2m/ROTC7M2stUVXd+QVkIzEiLso1x+0EfO4682w/RHlrskId
P+7WiD8ZhIndeVPVk9cUCfZmhalO3L6sAxv5booAbhWxK+XT6RRyRTU53ZMMDDzk
vX1MDcQbie1LgVcNIsw/kDGqtIUUpVOs4u9tSnF/MdrZ6d9xYLBlPGntQuJm6QIB
3pDZvJpiR6WrwLyVxCO5xjxXv/9yeNknn6hR+nowXJksCAXfRWC7pSeuCduCQYdw
LPCGB9dBkdKHQeaAAOYDKX12gDccTe0M1tLwBDRthAf3fhlw4DVhqFuWjjogjH7j
JdO2z4Eid+i8M94rEaTQw7XWQcdv3zbnIyIoHJmuzEkYSsEih7d/3yb0nPKY4FYN
01QiApE2A5mP9Kj8Pbcy4fI1+ZD+2tCdCtiRd3Wbk9EL/Sq1p/9cUdQvsFKqlO1x
qzN1az6mgTBoSWlaTXjzn1FdTg78eNVr39MNLKdAX2szKn9bh+ulhdoeU6gr1wQ6
e68/swVKl8CvlcNgAGlNbuTlkvvS6RmyUNby6AUNRGfU0HVIuVCmusLiYgF6nmfQ
zr3Ix2OQS+msl0+qvMNoD4k0Zv5It6Y4mHEicnletnv5MsFnxyB7eRoDYSBG7DvA
/XijEq6zw9wuHZ8MvFqXYmcOvn91nAIwpjSIa7GD9DWUXqxs1Y2iZ8J2F82PjSZw
KT5XWYryPZjztMvr2Dau6cjf97HVw4daGtT4lbO6ZGsDXDA8n5FuiibzgE3cclIf
3X7zWI8ie8b2tSQzaBdThCDfS7ER8E6xn+MWEhGOuWnq2jo0uEtPZhIvrFW6y+vY
wNvNqbuGUUDaOCqNQ2rhyUvvqF4iJJyO16MyeORYdexOluFS2YbLgkvRaNJ7F6gq
0yurIJKw1GnYQy9WVKn5R7juHV5veOe2emTalvTwhrywuZP1+WVejc2CcU6xeUsQ
jlfzS05dDnY9nPsstYG8FdPDLF0gVpqmp3UyXRVXrqwF0Gs/Gv7uEPRBj6K3ukeg
JwjCYOcfRxbgr0/Ok343bYX7swWsunibWLVUzqZGBadXsclsSKgy4FJ2F6XqVPHh
l+ZjqjT+eo063KQm/7slKE6XmPXKgv+HJBbDBsxvTnRWTCvwvhG4S5IKxFL3IOTT
3pstxwVZmSzuyTP4g8Ul6cAZYY17Ke2YFdACfkPFlPx2FQc/wHbglBwnm6iL16Of
xZYhA8tlRD3FKVCzviCTDVqsurCfvpp4L6VmRm29cZIXqDqjR61bLtyc5Nr+09Zc
4gQ5369STPryrJ4N2aJXRJIan0JLR5ptUdYaf2I8Hj5fTOlVeJA5l8HNu0Uf/rRk
c/E/InhoZhKN3sglTMICPGYy9MKz8PmESttk7ThLD1k33dlOZfQiO7uwoXWHrknC
opWlzMw3D/d4Q7kBpwlM4aXb3Y0YN8SD8C3VE4kZeUMwxLgd72nHBKXTGNFlLedO
jhkpaD311jAd9dzwOA1P8rkjels+Int9yoDFR+JFgLChSM/dcJt44L+kMhDkDQSE
B44Foa9yYNwhAePD9LJ8Em4ZXV5ULVXfI9vPD3jjfc/uanZ+JBosSPQ86ox5HYYl
v0QEuuuc9ifts3PWwi1N0Nq7j5IhFTT2Zzt5VniC/v+IxKkA+DuK3v4/uD0ck+rq
+5eX3fVCB5twyvVjM0/EZJ80PPFDTdmdl2eVAO7g7JE/JzcV13Ur5/0r9rRdXn5D
Dg8k5cBsd/g5Pa5IrpHACcEQGOrUaUKMK67O9Z0VKy/GbGmFevRVL41aGj0r/3AI
1nodjNJvwHxqoFStoKVJCEvAA7a7tRaIkvL6eAvbpVRrGGdlxEQI3ayYDc/6G2u3
Agaw6SDl0gUikhD8n1Hf7zO0+8fgoPvMkvWARrtiVRm8DOD0JragGX1BW0nwJLcL
ivDbzpLnDShjRxqGvMwHxIHHSFCLUEcZI1mQ1X+gb1Vi18vxb1rjUPB1FK4qKi9T
X3vYS7zvrdj2S8qqP7U1pGG5B5S24s6fHfzAdcafktsg+XhGHSvcUIoAHu0OqnW0
MP9gmkjusvBzG0khWzqLdLKvKOpvntN3UETJPcnUUm8qksRN0hMBlYmJic8mqc/W
YtetKU3RzMqJwC3/3q+B9Tlnct8hftDE74SGEtuFZ4b4F4tx85uli1DWBKZtnZXE
1l/3um5vkWUZz3FGGchi93lpQIwFniOCd0ZU7vcWEa2V/zzGPOpkN3lAQfry/K9W
98D3PhQhCy3Ptm/11BSw9BgS/mn+UB4NLv4Hp7Jb9giEPVQxNLu7sJFMohN2Sk45
WwgrVev0ktIGOGllOW2ZN8VU1bWBevhp0kQRRf4cekNR7RfT/ERkef/PHYfbTd1O
AmeYjaaJJL5jdDWiru9+sf/L3NE53v4mF/p4hJqN8bRa7X4xTwZRe/qMiEeu1sfl
VDtwgruKFjTuygsacQMtZ9W9nOG7Stv13IAXIj5dNiHLCT9WfBi619c969NachXU
B+/ENkwNDXtLJI5BbLIclWjm0b9Gil/Loo0DGMjSYU8KZ6g2RojaZVuntoji7NV7
nZmU4VDkzu2bTaCTWiSXkj6CgnE0QfY5aUF+ZooexS9JM6eYkrrU/RitREGpE1Ie
IBY5MDsVemUOsdHs6LBLPFkBTbBk6qQsGYFA7pfbBhic6Yw6DbsNox0j+yBm6hqU
9UFsOhFKfbX+iE0f4nLQO0+tGrugUny1BKMRQFMOtUEqW0YSVRQIbH+ZJ6d1yHOz
Xt+s8wg0T/M2G6TWHRn5njWCsS+E1ewgMqyikiFDjhRnSk65IiEXX6s6TGHNjPr6
KYD2TPW2xQ66acbcxtRT2x0H15LNDYP+cDeHD6vbwKKCKRT1L3qg9MhYgeOodnxN
VFvMZm6bqnDBF7vJP0i+gwNLVwvBNhdGBEhvZJcDBLkgTsAtgJm2cp7fP3fTMyw4
fE02k2YSaGpAW+qS4M6shV1Mw0fCLBKVIm+CAtuFoPPMkeRl0QL0hQOIxGfCqRFw
OW4PQSY/JDCZ/ZQX3iyGtDByhbGxPPQnC67CKbyMKXhKbU/AzaPf6p9ftBZWSBcQ
rRhvTlxlqQww/GApYtvmhYWIuciohjanN8wVjvdnx+qATKkGUTmtlkCOjeJznPre
M01l5AaLgjPQQoau8gjy78/TgKZ+nv8Q2S59uvFatN2QCnIGf3JCw9mdZ+6/QKXg
Xtb4rYEUBv4m/kYiD0Jx/dN2Hop2mwuunMCAHxgs9DcXf9vA1fC+2D/qp9K8pFGY
3Dji+JOgSCdeEmrrRx+S6o8w4poVdhEUbQtl5sivisxJETk9K1fLGc/tkcjA07dZ
2TUh+7gxOZlwI2nSIk7MYTFJieLzJ+VsNP+Usv4DHVq0jEmSxeUbwtEKKN/8aRoX
M+I/86pCaCacHC4MADteC1IKj2zroSievbLn1xroAPJ8PzBNiI7hPXAEtGJgRHqk
SwLuZvaGNhMVDENBMHk35S7paNAdlIurujSo6QBvaR8JvebwXbXcKHkxNC5X12OV
tRAacTBLD3ndot5HwcduatCSsS3Aeci6PPILUcHqHwROqUDc40niepoyN92OBHph
QJzae6lADTsAT9iw3IH1YtB/aba575ZYaxnBLMJMemuRG22zxnxsWrtLdeuyStMm
T5X3aDjiZay0UFJbaoUcKZ+OubbNn008guh4cUYf4ajGeK7z0yzdZ+xrxOzhf4ru
etyUJSkZ3R0zj8MTCIrDd1kNqxv5CqOrgWDcX5O1sZM9KB76+2Uhg/mQ/CIswk6b
x190Ul2F0SDpRXLv4Wmzhw0DzEOXrIAgTkfDbxfpi1PKW96KCUqc2S8JK2i4sLzn
3VMo6WivayBAhOb/Y9jODkKMH1lS3zOwLNNrtzSuBtyAQQyDP1CnWDX+fPskHAsi
osL7Dp+udF19CSio+oQBENc+4FmnKJwjEBpjjujQnytfrGQRLzzX9EBVr6ylvzdM
LeHZBp5AAY5sMsPhwDJq/vVbOJyqiGl6MyfEsaI7gWJocUFtWJjMIDa6oQByd4Ld
pGdVgF4Ws2FlrUFRmFdjcsiaey9q/sZS/bsm/f/Qyk0SLHEA8syFTTbDz+HwJa+8
zEgX9LminRmy8nX6p0SorRylqTa4xgNZEj5hKMruX4yfCUoyufaARL9hSionNMD6
YEKpJ/2rsned9rO90cUGqc7Aor1enGyuH9tk9404ybdB1hvbY1lL7DMP+T714gci
B4gTQ7uXLmFRr/2SBwpdYi+LwgSoxTqjRSzlJeH+r6WMEKBGv0GWZhADE3mM49ZH
6mb8yUrh6SHRAPIcqsbNk5R2LBsLXSMpib71ABMM+wOwYRHIUZpKUqjypg5V/nF0
U6fBw4tMIln2z9dGXnM6gEQorF8eAdG1ZHzk1D/gwRIVYZnGasJZ8RCdi7DBRwk1
WqDU/qi/f2EwRN7NM4+69ApBIg8cs+mmukXG8GDlbOXYGvgr8S4AiFJUx8WBQiq5
REv3iTNgErWDPU1c61KdT+CouThs9icUhcypcKeS2XRFKLmlfzWedQm5VrpyZW8p
XoygcWDOlBBXRHhvr6wgCS6z+YFutF5yvUj7v5xjsljzrzNK7jTRqvoyZpQ0RJgJ
75WyFLFjO9gH8qOfSbkS10pYNFXOJv3h8hUMm9+bxLRjeD5uy7OvByJQQYP2zgav
9SOPwS+qLQ+PhiW+oxBHrERzQfDeK6OpUSZE/OBBGCB6cHSzxes50bLzucFoktys
bmcyveiXOeNGl5mEPmR0zdC3dVEJcVe5Rh5hnF/KPjXdkEtJvgUGxFscybfUY16B
yhGAn6qYrno7nN3f5/HFjVb5jwJ8+Neoa9OiXW68o48htJN6P6jdtzk9sUWGTyVL
0MsbKcKBOanZ9uTn5Yp5VnRO1YsZQZx1a7xfBcE/hMmTNqDdWMGBFJaVp83w0RAv
USEcIE1vqDHYv2FfQJpWTpqTmuwHIg4AhTjwiFMddDTMX2rXVcIwrH3hYvqnZNn2
ymszb42pFqUVjYb+V32Yo0qkRSwCIqXLud1T8AZJuYn3ek3l9RkT6EOxG5knvx0D
zQrmt3wX3q+drNlwve9qr2jnZoQ7ZqbHXH1bG7HhTJnVYfq6DCcFDChKI4ncuu64
ltGt+USJppOmh0Dzc506RaGMl3cePs6rR6RprFNkJujb9dWtAhxecnHCKJlhPxRz
ydNRF1svTvxws0RhKl4sA/0hoKon/eQBrPUlm40cVVJFbNCy36lxUlDR9TxLuOgy
pFtzvsKm+UnB95Ydtv5LQGumAbH1tgk/PavuONTTbD+C8HaPvNcrX/nt16QxGSSC
GPzqQXujG/1Q4KIGg8WM8aLr0Jl4JcHZp+CaXJ9KARxyqWE2L/UZnTZ0kUK5UyVe
ZkNbBWZcnk86rMVwSAqZFlSsS3ZloWW3RYVABsh3TruKIDE7qaOUfJZkj4IEym13
X8stAU6OoR9P73Ss1V76hPdjMcun3jHp53gekPxzTtyTfaxBx4G0eMGqf5LFYiY9
orGJLf0zV2ThFxdkc+pTXnEfdyR71S8cfbyAI6VmfKWAwPn0T4f9jmoNrnOODQ1T
WFp9/lnpr4a3kScJLAAjUZfAMHL0uCOfFj70fiIHfoD33Gu67kQGdTZS6BtU0Hbs
9MvvUxF8Y81X9/mylMqqG0rqsU1AtHJgvajSQmBL7tx/1jwkt8mvaVdO9RQqRNto
Acrip3st9XdbN/MUN1UOOqAuVSMX6G09j0rnOKeOZkbR5voKRrKT8SeevR9/J0E5
zuOB77bg/vP1YdzDQouMxmQBojOwyp5rRUoYhpRD6Jo6RnNlouxTLe4ufKGXbWxV
P5Nar5zTgqDG7TyGONa6Dpe1dBWbHKyrzUCguADaCULF2huw6mP8j4hyABsFiBGY
ThQu0zVmeyIcLL6cuqCE3EPPy1H26spV/2IAPXapi6+xNIYxHFB4sWghom00x+pe
DGsG1gmDs+hkwaS9yhSou1Q/r7+8ota9Y0fnIEe6K9uZuunVtiZUUNlXLiR1mHh2
MflnLPI3n8dEeS/jLQzXPxwXOxpheV8hTIlCRGMAcfLHWBk0nqn55J/8f6tGP5AO
trOq5tsle1ZfNT3wpoYRqRIlTVHxtIxHBixCNqnAaa7PkhEacswNutI3wPqcXN3D
sRfOeSGIdY9i9kz3qg/a2FWcZlbo0CG0kZTy536OqGdVzo851ghVzHYYAhqtnFE3
CXKbzmzwLmV9IKtpoQK2cDDsWD2R7TR+EeVpoEVTBQ1z3RGk6hU06d38YodJySAH
RTNlAhj85Wp//xw4Rlm1qy2RU7XIRjIq8waCWxAv6qOOof5JubvUorvw6Y95OB/8
iuZhUfQ88Y6uuTe9OEAjTI1kN7sQNpqc3VXZKeZobz8RGgo+HgyQxr85Z8byQUmb
0g0PozK3icii26Uq8KEMl4K+S3cApkLZH3XJOgONjroTGW/OsFPD9nMY3y4hD2xh
OCbSnT538OGgcU1gfPkyT4CIlzAKu8eVxgWFQCHkhxfdF/Apk8Pyjbzv9GBf7/Fl
OxrY/FMrbCNUumJ6BTrO57u7vfOFfVe3fLSFOL4jHKR8hijjfhJBa+ZLZXswNBKl
LjtjFCj1rAubRFr7PvCq/tVosotZMKfXM4HcTQE/fEcJlwdBCjoxIfZ3yBJ5NE0O
xh6ARpu2169OygCSsX/Agr2d3IMyJcsqekGlDy0dSvimQjH4QPoeG3urhi7AD1i+
qLEOrfd3OYApQaCGDgCk/7DuT93w7KPq4fy0eguC70Jo0kLmcNkT8JW0i28fHpkP
m2bAqzTx8AoXtvA9NsMatQeTefxVK5hcbFsbKHny9Eikg/6Md6qO/U7pwqzvzB0m
Dy0n34UwLbTD4sHP7QR7/mvIB6/40ZJT18v2TFT5bWB20yKhCT3FJfevmJs5Xq/S
daYjRsSK/dISh4ajZB0wXDyB3fxBLGwW6dW8k3XzpzMRiSxzo3GmpcOSZCnw0Hkn
RKMOh1J77yT1LraFD3gQzLjlk7fl8TSSwPpaA81fy8gJPHs+xfY1tUNjgA4RUX1/
EgDpHUXo7HwSgSi0UDlDnfCsdwiLcZyzfMKBC2B4XTsgV8ZSzcVN+4eNjazalD/D
TlOcKDcGBULdRinvVjzS7Qu9GV7k1/yu+sngIHCAMoJC+4TJV6xQXO9jTFMK+0Fq
twzmc22UNC0kPCm1DdDCF5daKcVnjQskxWV5j1Ils5uh9e+h78jtY7rkVhXnkbG/
67uV/eCS79BLn8PKDMl6V9z9hsdt4sD9GfavFwasv1csoEYeRGL1x9IHGZ7Wx1vk
rSosaoVlwNZCmK/8mmT1Rw4AhBM72dhtYTfy0NmdPOY7wI2zFPYQWeX3DMo3kq9r
cpVXvHF1K8M/4bmpAwiBwgMGH89iW0AZoA/XoiT0vuaBp0vBN79zMiUzITFnmcUB
DEzn38R0AjD7g5Fxgag01QyeRrHhUGnmKR0rz3ndVGyRShBxiLpG9InIjJtAT5VW
dn9N462AUq2xvn8K+cVvPZPdLv1GvjyXnxAxCBdlUkESD+qussrt9wGefLOTi4eK
4QCJzUrUDH8huE8g7cr9DqaYboW9RtgNM4RwvcUUucEklfV/8doc5rubSHrZHnGq
OKMYAKTrBwMRHCL3lLQ476yaZPR8FNqFv7VXb48m0FM9XOrhTP6UxWd2qpQHbiHd
rcO/Mv55+LcTtrXQHBI8nswK1DJsFiLXOXiUvi/5gT+8YHR42zutSXpWdHCjI4R9
y7IXXLObVRydeS1Tf9Qta8KjooLSEELrmfP6KNQkJ46x4yQ9aNyFdMeIZibnsrT8
8pyOhWV3444z1C2gNM3y7wmpFsbAfs53u5ipwC/0B/pepNP9rCzaW0P1BPIrddQ8
dw+YbxNpfZSczijf2CumPtDRpMHZqLmt+d/+poU+WtCUk41ou2iYlXAc8vqrz63z
7TV+zFU+HqARHuILwKh/302BzGBlg4AH0IUFm1YcDXKsg6YWuwIibQy24A+WTmVu
L4U3S1wlk/q8q/UJ0wr5U9FzITT27t9AsTkzKbZh+YAHWkMO1FPDMF3XlWiF+fAf
GJpUvmWh0GBIdCTRL1mtrrc0BrUauUASli7nLiV5+73ifmfPJqHZTY+Loi15rbaz
KFbF2nCnUgUeNWfXyRChEV0VmlGbycype7fQSei7JsOxpE2yOb5io0S2xy4rNS/6
qOxMvQQKcgPxvOmv8IIqYFmfXp+mP2nGtHrE/Cog8eUuMvgZ00tlfU6d8qOcmibK
IHoddnGtqUGvhLg6G4APIFy/o4MbSwihcCBojKDIMqZk19+lO6uyHJC/PAcKhg8Q
PrE/zZKryWmvYoAv0kdNbIXgn19LJ82aWnbfyrVJo33gG4cHAZtRw26yDHsIbd0M
Mt1Dny7JUiJWNbUdwoM8j+hkUda4ZMONxtIfWnyKkBFPbjVv7oJdskBkZSl7p2uR
0jUDjy5Jcf0sQ/UfkX/mtvghmADWVItnOE1ICeFSARciqjs8aUcAp0m3fl5TkyK1
Erv1rRTSRa/S3iWGvziY8qh3soH6SOj+fbeJnvE8oI6AP7+WUb0vRIX3UTTy3Yhh
2OmKAUwDnKPAHuWutOxxwMMzVFQ67VffThzUnY+8BmNZBkd0cf/2YXn11DeuSKHA
qxDPJvWA/PLHs17qJEYKIlvOdUFx0B2MKqsSsI64GX24Fxi2mk6zgSt7pnCL4IBh
8/7MmKboFOwIhMA2pRdOmec/Eppybu8jHoKURSY8h9jEAc15M3AqfqcZH223uo8X
8O08qxzOZJs8k5raz088MMToCNiEdeq0tPQaEgcP6VnJ+OsHIdz7JsEYlwSzDNmP
zeH7SeMQQUdRIphBwFQkXJdOw7cWIaTWDfS9saKMnPW9FhnW0WRXC+0LBlBCMnuF
JXuNVCe/0sq1gKTN33iHoROjL9CBP+JWx5JdWBr/Kv9XZq2jBZeu8YOrZDVQETYS
YuP3rm/tEMzC+E+OJh3NFqbJ6UiW/mj/0xgIMqG6aEvPS3l+UHeyrikJyRIcNNsJ
Ou9PC8l/M7EFqkEc6Q4u5uNW1J6yoNtiwYxONYe3VlTp2FUzd2wo84g0wRq95ry4
zHnvzAQ+snm60hIjczOEOR5B8hYDHuEHdlqQ6q/YNcGiaAOzyCvHt6QE3OFN4kGP
a8nhUXslTcHI9V/ni2SRFoBNN6Qd3GnUbUyZ/JlrvgOe5XLpRkUF7vsdBz2JkP0l
qSe11lN5XyC+EHLBYeoaJdUgN8MsY6NQbv5w4m5EYm0sotudoapzgcDxkTUVCHEP
cZ99M9DDQaTBFjSZmHj6QFBBKxeLBEmsqIinjpaSV37zLOPbD8GS4865YYKbcBmH
dWQDv2++5ivYe8Pi2imY/gnA9kp7jjwcVGrMyNI0GxjdafodWhvCahsp7pqgLQYU
YsV/iJe+6pRLIXPWUc2CblDtVmmengKjuRTrrwwShZhXJQqJVicXQzYXbmCer+CS
deAzDWOaHCl9l6XqFScJ8lZKr2jZjLSjzQL184advHVmhE18yS4PWo67wcm/uyL4
2daqoQSVd5OAGlNqZf/Wp6xnKMngL2NqRHymHUpP9KsqW/kQ3Jjl+2cziRgGLUUy
TjcrNUaTv+Wj8n4qqRDBqEyUjvnYowxX/B0/9Mqc5pTWSPgXfjGNrANE9kHsGrqz
SNSCFDoH/AJu/rCMry1qaZMZUsJE8lynrm/czPJzMDLHqh9bRLVTy0A+dMqQr7++
BYKUnJDd/0js+6ID+clMg56Jh5lNzB/V2z4PWYfKVTs7pJMJ9p+HXEJSq7/I6Dzb
zXb2/2ZtEe+dknZu0FeT5NrdJpX4lnf3FkkMi4rdN3z6rFrSSlcq5+qgHJH7lRTe
qlZebgajYZbSauhYGkM4mdUyenMQUK/0Yd0YznnOfTb8UuhaNPzL/BtWEN7fPhU5
w1aOUyknyNOsaED3AvsElXXamw/c+wGMXDbI4hHBb0goWCiAzZRnV8y2uQsJWYtv
KW9un3dpcNgMBU18f8OQWks4uJpK0GxIdNGGUTZH/rWihUCdOg7PuU/c5Say/uCA
mKyrDQ3NALWfZz/9e5ShnLZHZSq4KEDWgll3MBtMzDSmsXgyNmYbLqAgBCdmuZYy
FbJSrHCsOlT/9wLboyvpjvDeFCugzy1lwZokTvdqfQANppz/i1myiox3+XucBD2y
HnlRvoHyMOfF6TXOme0ueTcTlgHA5s8VXbwxglzOrHAIw2aoYZ8tUgGYuBYx73Cm
tRSSG3aFZAVzKwxY99UifDoTtGYgfxGasqz1ytlVcZuUSs+hW8uxE+dw1xdfCVpl
YNkUUKFEUtZ/MO5+1C4YkayAk/ZJlVYB0S+PEJPp8fE/EoQx5U/z+UnU61MwbQo3
Bihus8H6hoipNaGIlBDXuT2Msk5ye358nfj4uKd3IPTrl3kyOMcN4b2mYLrdRynF
cLRld3sN22nyNjgpFftWQdeN3OoUj8hiU2S1siGnLMZkgU8qNny04aPeqEPI+R+Q
Hbqy5oStiLdbzHAz8d/QFPYi3sR6U5ZUyWbP44PTIuLLRMyAcqPo1Fc3kpT7ijt3
pmo6f8K7DXkvoumq9YFZ+UdOLQ/9Fc9B/I2Ho14r0Sz8kXyOpNbx8yQFw5vQbtkN
N9ohQu019Dhg/Eu0e0Bf/R3uR/afdPqFpf+L3JOBxyF1UT7uoEb4YHM+Uye0p+Lb
8iCYt/QEQz4FwvCMe9rRfivptoMoPSHwUFxRhoe8OnnQMifiAEfqGd9gU6qFvvn2
rE9n6KhICl13d3kg4Cck35aydY/1F+lZbFCu5YPnx86lzFULk6V1vIoImRIB4eVT
NlW3qiymrxwK6Twr1ZIVbdyb69U2zKTlVeNokQrANLvwpk/sTL1DFIRIV3gbCHX3
SCLclG/CnMphUytQtapx8cGlGCUjm91zumq06uOJF40/sbhQk5szt+XAzOkXH3T+
WgEDLx4ZdaD/+WATz9R4+ZYaL8PDpuMseUbNUJABd6oKf5SGLjAFAO2lEMLlXnBu
LjLmTtuqguPIFFvc1voWkwJALtU7YqDNFENNo6pIpyvdNgXsRZ4vmbRUnaBFvQCi
jV4cuTst1VKWRs89u0ar7L4Y286t9T0ZarCl8dWIh4lTD3RAlMSKRBrtqALJDhXY
TJYTzk+mdWBq9wtUSy3iikfHKRBgrIls21VgJ18hVKOonN5lR61Iwa/xfaJUDV8F
HX+cBTj9jOjziugjk3RtqcSiNW4jzZ1aymjx4Xadnd5A7Hxpix5dn7kK9TCoJqdZ
m+T2/EGOOIFUzMHPLdEj7pQQ7E9L36BgBkkic+V2Ap68dHcUUDmTTY3n0jkNCDYw
IIFE3KFPJz+rg98p8TrOW9/RohsV26lu9QY3dFW/GClFBgu2ODjuXob3QHCWLOvi
xwMSFe4dbEt130WXOfqhCUfM8qhdmCATYAKKvoR8POR/+cxuMIZ+N0LpZw/yMiPn
LeXlGNirlG8hQA5HpDcoxGSuxN+GEshU/HW8rAX32Ck2kcPRd/psdkqteOK7tWuk
zZDk8o1z0nJGbPmBriSqxvbzgtpXdmgEe3gykzun3yO0hev/3unGmbJcDrFOeJsL
xq7XgRNATuvdcAUdTc7O6pkR0zNB3+FZnpa2qLKdcBnsXcY/FQhls6Ik7/bQOmxe
OsBeaLlE1+p+PMyLTgI9BAbaVd9WZTYQIGT81dYSGJ0MqG02nWPtESjATlq/v9Cr
Rbo1QQPw8JGKhzLjsDk8HlldwkRYjEo+2O5KgN6ZuBIgQRNpt+V5MDnwCCvzomER
Wo5rmiPxF1ryh8/iZIp4AKcR6f1L3fQ2uMZFBLHQYZ/OTdT02vJgSYSXLRTgU4rp
3VatTbj/a0ofUrYMO+EkQQ11ZdXDb6mYyryBKNhlGAO7YSbufFt/rumce+KlXPXY
9qW6NPJKL2XRxM7pGO4UHT/7se4ysacNG1CqaHOiUYrkM35A8Whlt/rROgwOaiaD
ng1ti3o9vS6zwPQLzJH828z+sNPVHU3n6fXHHhT8bMVZzE/IvEmc/4Gw33GYhLOz
Q1xE/5Xitx49qRJO9id/eaA2XSQnzdSeQkNeD3bOjl+in2fEG0dvngwdzIZmEuFj
3Hxs1EtJRbqI1n1zXSQQTEoottzHCJBy2mbmo4/0Fq55zRrr8339fk31/47loUqQ
fEQrU4AWSjZtLvzeb4lFpekLNakojd78t3VYVOVlvtaftX3fw5CGpTb1UikKJLcq
EqzAwUzCvZfhptr9QUJIgjENtrzlKsghAQy1VJU7LNwgmpTEb9MIi9dnyzBnEc6v
GGfvBhq0bJOoX0Nf0A+pRFCgB0YsEbh2ANb+P5kwtU+ql+57h1K2ryYMh6cLv7ja
FNwz5f1KNSRtC3jY0MiLStNeYhjC0MhES/lhQ6MyvTzDWvKuvSnEDordyAhz3HI/
HgvyeXGCu0NRoE9+k/5fITSicPL3cbTZ6CUXVHu00XL/VKqw/b1smyAhUyth8l75
A3BVSzPipFbt8+tnI7BttmhLBepVzhllckhr6/Uabw0Gq9Jp3aDg8l5QmxJ9aTrH
tdwqwMWc5ISVCfFzR2/n5IjDXt3eEDOlvlimvtxWQ5AXGwZZ+6tNuDnKrIYC59zn
42Qqnnjq4/37ZxdpPI9WxrP5MGWe7GUijl0MlcfYSECsXqrK6mbODR6ViuN4eJwP
EjqHplwSXa7F2r311aDIYwIBAh7Bq8Yrm6epGNMKqdFqsYqC9RPO52FQixCgFNkN
LBLVWGaMeJiQFG7l3/WpnijgEAEs2zmdDKk9x73uYa7u4PRuHhheRlySY+nF/E3b
gSpOqS2wD/M7nIhMagfQ4dBoLSprHpToPIvDYZDTiOq0iatf0si3od4pZb6/sOVf
EurP82HHsIaMq1xIhimGelRpaPfBYPj7fU4UsXZyGZnjoODErOef9I/43JomeVpd
l+w8L+UOgqt2i+04We26+6HLYsI2f00x0dZKt0hpXC6Y5dpeZO2fhMgeuVg0W7qz
0ZheVM4P5kqglMkSvvWeL7QLMtaPmrdL6zP4w+RJ0jMw5TGf9K7+xOLqmobTi/0m
74Wg/xqPD/bhzYctUsMyXzKy4wRP8Ktovq8QCCuZWQ8s6Wi4FJ9KT8Iav9dK5ALg
ezI7BViIm03YifPRoV3fDzyY/bzsN19XKqj9jsj82fABMomtFybUFyNIqRfjEqq6
5ZUKEgHi8rn3aOBqjzv8Emltj76Ahve5KiEu6Fm4VLO/9Q/b079z2XNNZ0cmnPf4
ZpXajjvUGv4dv4+ABaGTNuHc79pDDuBBf3rMD1pjSzxZWS6h+qKPg3zZxoSoUior
SXFl+X7qVx4p9n6lqpu6g4fSZKWxPY83MTZT4yFqrG1H6jfdjKvFi5qL1rHBByKn
A3c05D9cfQbf3n9xABPW7liDP5o1Y4ygS/kRliDS5oTAMja3zyA7ZAmMhIuKlH/A
4HRm5jbWEOadY8BOt28JPdtORgAsU4TkSDf3vTLLAyXWfrGhjDisNwfxgyNXT7Sd
2YFb1OsbmPtDVGYlGrjE0/mO+ImeCL0rBRTG2cl3YVB7Jl7OKEqFxEWhmQAllhk3
8BLJeGmYxToxYtxwfdcuzUEQe0sxPKZu1GCp7/sNVciSxPSCSot8Tg47fKippfZ+
bzaQ6wBa6ZPIjfQrYuIGmyNX9z5lReM6bH6usFzDVsmoJBiwgw/4bgHI0ewQ3tHq
gsA02silIBuqLoZFnCS0JfJMA3YJxqMTP06yGjPOhvXhKepwCvdOemdup6mevZC7
Fv09BAThvGmflChSiWzy9GL1knINs+1bvwAoUdmMCP+/um7FN0IMG0um8s8yrUUd
RF7pINHAs55IEhKPG2b3nP+QZjk6NLTqXsLnYychhC1pC8nbioEQUB8YGCjekfgu
/k6uS8yBocqeG4PnHaTVSV+T5Tvhhe/bdteyApkbRfqmKJa1FYmlx84qlxnRJPes
b9Iqo79WitJWT+b2q6c1BnrirXEsAtg4ZLP2xaySFzhkyWqeQi+63XZakx8pwUsH
riRPDxHkytAecWA9v7ekWAYtjpQ7KNymWWOURUdA07H177GfO9NPYbI48i8NJW3M
8PaObiCHfjUdZQfjAPuDJprA7ui6wCVrM2ylo/ZSsxYnt56KbyxvqEDDVdS0o0xJ
V95So6ZqYmJ5DFuoGCFWzJmug5e0ETWoH5P6DW6LxSjZI9ldi+oG5LpbsFuGsZSK
03M3MYFIoL1OZqwsJn0z6vrEGgNj/wQt0Lf7LAEIsYUjY8Mje/zBXmljscP6NEXe
GwGv+9R8s5hLGvXDqZ24Ic/qSKZ4V9aShct58h9tjlNCx/KK/bsspyoy+9KTfKSw
psLHJRkwOsWshKVW51aYmTtL2TS6LYtr+QfMuIcAbh4HNbLFgPZN78O0cIXxAKyG
hGJSRQAjHKr01X9qN6pTklSfmY9LtaGoAin+k+L0UnObJgJ0qPk19cEARDBanUTh
TJn+ma1mFhWNidB9c/4i5yBazhb2d+jVfeC71pFQr2GiyD4B9frxFzS3CrdehtA8
ABD1pwo5j8lrwnE940Ifq+6vwKULuhpYNmtDTTb6qZQ/0vErAHR3m1RQ0INa/ONx
CLx8kV4BfKsMr9N5hktGsmQbUCKPbwQwTAix5YHxKXORkCjVlbuzCZxJqTd21cy6
wuCXUcFzurQfIynsbuxQg83WIEfMhYvdKFmeJ6RPaiKk/xRcdJanGyfUHm2HCaaP
PSEsKIsyajS+2iofgXUMp1bRuTTBl8cZXQitehuex+fhRapFWz2sI1gY7Hht0L4A
HVcmcDQomgIREEEqKQFE/Av3rmxQEZMPHuGnd/nwsjE5CzcsVzIBZ6TMgfwPSlXH
F97VxlzuEnjFa9zy3NJ06hH/zAlLo0sYz43F8XwfxGNcye5lqy+RkHengWBBim2h
EonIgJ/7kFGH4cPuiJiuTd6iCbXVsD0Rp2TbEkvojokSNgHKijngCV7U0LCocJS/
AXOFLsLjnJ/6mSI6P07dpxpyQBt7eH7iAFzeA4kip1hP4NdPqYF+wp6q4FGCVoFu
wd+nTJLITMrZwEDyRI5iFcP9ukIBDyEgvITp7lp5vLFv374YAA4O/k1MDybDnvpo
7w6i2biFZfrmcyPF6NBE2aVEOmGOeiNscr6dTqFD7lKD9Kh7fjeyLh905WTaT4iq
6/kCpL+SmLWRmkRReaWeWJLydZ4pRVCKrmN12IKIUnBry3BcVmXzt/XCSpYEX9J0
t+3QtaQB5qLdNp8tGdORCinIfLRiZ73rIkJ6eZzeqphUWiaVimFCOEzJQ5IowNG1
4pxq8kd3mik+xPbj2pDM/epf2JJRl+7q0OdEQTOYkHbKRobecrYzao485qau2F1v
hF2I32SriI+Axx14Qp3uVRwCFfCgCDE3t57eVr2ccEl4+DzSpHwxXWxnBpTP4W6V
578CFjL/1rU9erNR6rq3FIuSIEd8nFLzOOrE+vDtm4RkFo50JZLfxr3adYrTMsjW
Do2/cIetp7Y309bz0zfNjnC6z68c94B6NJ/OrFURUDVP2I54wOds+v/IUvboXg/d
hYk94Pto8zVXVR7CjBplbZEPdYehBZFEJrkI4lzt+2KTQtDkk7yee1OIYIGrCbTM
Uf46SP483MJhF9as+ezMXLeKbSRwJu9YWy/zsE5IofjXkfK+VUWFS8/NWi3vh90Z
ZSgwf1tdE2F8sh43l6iJX+iu5MmW9pFvp7Q4zW+tCS82S1UwAMFM/M9BLULFfhyr
P/1x75B7IJmKuTveAchoHIBzCFCiODDggK/gnUuoGAgp7z4DXp9896G/BlQIbSaS
mS/oOgmVlCfQwPsdj0XZSqrPgL8wGGfMHPknGCqyCmrbKVxzSz37JwIvL1dNKp+R
YjLbYP6yUN7CC4hSGpxDdZSU4wh3q2ir7c4wLPwYikI5USOVBdp9896wGYazk2ok
Jte90uXFmo+Tk+9iE2aa1rrr2LGkXjV+Xkinf4OlltICke47ntKUYBTuYc2j9QXv
9vYsblH6mbKFdG/yItmJNuSYVbsYVgc0eHCBuC4cvSH+XF15vZU0VmBBNZeDrdRJ
2p8PZj0xW0ZcvIwSrEQAbUzXpcRezTrku01CCZvSEG6sYO+/RDPwZ9EkSkbRnbJk
xmRXrmTxJ45UlZCVABHiVn3QoLABKy9ByswTiKLsm4v8/1jsvBYW1OgjwrON+86v
fl1OpbzwOWQhBKSZScRk9MfhKQ5w9SfL5ksBosBjb8IN5HktwSoYJ25BBmn23nXM
aJsWhM7mW2jHMevkaVWDaTRGtJhpE0WhH13cmF9rMHn7+rglEqkeP3qbJEj3l6K5
NaQ8NgZrKuCp8o2BikV67BDhdrD60Mm+wrntdP/yxjUpabS0Ur2zHenW/S8moODh
yKDXwLckNh9vFBu2HdtCpXEEn6DknRa5yG5Xvg8q3kIdgWrz00E6vqFuNnldt2Zj
7ZZAL9gys1PL0Q+eK+TmW2TLafYUkVHw+uqs0ppup/vOf7a1TOBMhl3lgXeL4i5c
shW3RvEk3iRTTGhDymFP1jylhuRuhcZYQbjwJl1zIjT8WOd2cDk5V7S5r+rVPHng
OTFxiqWnm+m0maEf7vDDZgKRa7Ze0y2FdHOoBJ5+6G8/UqUFQlDXGU/bNU6mxcEA
5AZrx8ZWKCBuUTp1N1f4Tzyg0O6WbNPTFi6SLmi8GeT4h7B0vKpxuf7ZV6rdT0/n
ScYT/DEw9uWlpB0P89O+WAkaZlpcFc7mVi/I6nlWeqMA+EXt2GRLIB7qomk9JY61
4KRpjl1eQA8qhty7C8Hbu5mkUMVS/UW2n/yn6HpmkLKtP3ZsQAr+7E5HuI3nxqf1
EfdpMJA/QfCdMrllsSpA15QSNtd8O86hpsRbZsWmKeh9w1Ka+tClrWm/mLRBz92X
+60q24+DjWihF7QLfN07Eju1j5qme+8kK2sK4jGYIQFm5fwuRUtx4xq+qzIBJaLG
m2MOXuQO6YqPHH7MqMqplenhc+Qx7ho2d+wGIWdKUB7ofLmCvfCv0hQnMD3MND6f
sc0Q6ZlkZZ6KNwm5wUmz1uBnczSLVlzk+jlcZg2OVZSo1RJOJo31+6NSYjHDeidm
WP3Vg9Lfm3aCrS0vPFbVwM/uZWTemVpS/L7WxQAw+tvS5wIMjVekqqbYtfPIiaXQ
8oLyFu0OSJu++yoyX980gnOEUgIBy67ckdF1HB8Ln1xSElsyxcpZcCN21ddam7j0
2VbMV38vIJMe+Ec8388hGVfewR9q1Mls835UsXuueTepqwu7WQckWWSdRn7E8KrU
0vWFPMcOisHofcJt5V/A2AtTE5pL/1FMZ3d+yfNSSMeAiUMnBsTCd4eDFOFcw9Wx
a/0pc8EZQ8GYf5G/a62RK/JUXMDy0ajj1g6U3acVYSzTmv98W6KEhKZqvi8iEWTx
I8xFJh+g05qzj4iOE2/9bXvrzqMvkImp7cilS3z1QYPHwDkZ+IsOW4kPtgC8h5cs
jvCtw2Qo/ZdWI+MGmDtC1wISt0ZQBzBp4mDD523VztJp2U1XlgKsQnaC9zBD3HLV
QCYVO7+iY/YuqA+fATvUlU8LnCu0cblWmd0pzGtX5TjRpJR5ZeEdyKAVObMqudYk
R7ZpmsJnN4zUfHQ/Nxz2kYx6ezgEqEjfu7GUZfDR868vjss/fzVFw/ZogJKLks+r
dqdwZNonArUehfq0j7LA28oZo79saXKT/vY3fQZRcqWH3s0AhCcOJOP1P3FJlGpX
Yshqzb+LoUQCJV7wb2eEPyEfCZmBJVlsyaItdcVjF5+YXY3xoNHwuQobAy4CV0SH
zvZKYoelkeAEHZcJCg5EJvvDWBVWaRLOgzCp5iHMKjYd4ZJG8DO+lZ4Zq82XxgP0
lSEGlfbcCMWzYUiPC6F/zftn/LhtLW5oCmyQSjAScAG4xkG+DUlYj/fO3KhPrXxu
BkTpVw/o5NUMwzmTzcaXy5fZ+pKlQo6z/DQZFsmu5GVOaGFT1QjUWRVZkeHfTFOX
EjSstuwymUkwsdrW9DbPvOAhK71a1fpbARfN/i4wr7Oafz2SBi83DG2gUk4Xbk0O
xCIzs2NdZqt5f+DdbAFZF24O4GUqFT8+237NRkyCwnDks+Bb2/VRgevGsIjjb6hX
7IrJ4JRSblDM5Q96hRpIXCh5PCJJ7Tr237uKs32rXssc8wHoVtNMsAbxvUhOx49C
PqygP9SxZR7626gxjcKWLJWFq3W1+49p7f06gW17XQgGQL+atO4Oh7PmUvY3frRC
IvZn6+ffWN2sySAv5SO/W7VWzkQHcGue2JnuHQM4G9xhKUNfLVPJ4XskqF0xGcLv
mp3lmNelNCWkHdyN2vbeyUCHU+Mp+REbeeRkc0+otMvsR8YkNDF37fxQdI+IuMLu
a1p7L2I45d0R/ABMEvENFCH1gtNHOqbn9RIHV9NSsRY4AeHwDfHDbTYc5o016//z
wsBjkqJMt4Hcp1KnBq2dFr93bE18Dn0t5Z5ZwQ3OEgy27jjxxCpSTl1sCqXhnfDA
QZVa16M4B/7O4X8fcOwIrZSLv9FUiplMYugSRpK12F6hWH7dWUlK7qSTxm6NerqE
Qs54mmTA+L2EO3vJXBPDZd8Axp7/MMC7oc4Ul5XjUZ7VJbzqqpSPw9lFK8aM5MlK
q6XsPTbGn4lP6upyJKSBeHzO91t5GCZ0A0i/Fe5B73Dz3kVPpSbbyaOWtU9ljYTo
2E22wbyB7ojDptwTRCR+BCnpLGpe0vsOkz183nt16cfwrwyF+Z0PsZnbZCDt9/Vz
aZqYzyLqR5xRWowezNqVkUlyKYaOaF6EpJ2JTqdWJS27ajBIWvvQ/lZEh1C8UyGp
PQgxyDr30B0nBFBJAFvyDUiNNAXPaRx/DFV9Rr+OmtQ7AB3Io48ucAYp0JI0wInZ
Op0qzIQLGZ0EyutS8OS1eVc24PBP7T75APGbSZnBonNCfHJBsGNLYYFJDSsw0z2G
5p9dqy/BnM7MlyEotog9yzKKrkwgeWatjz3cYOrkJm+JO1OBKM0wXtN5IXPIlHbA
B0BQrfLc4PhCy+mBvmQzxtBaJOuftCojUYpSP89IvDXVXDvI3RQ2nPP3ldvd5E0x
r8jQFtMXVYfQOplq1hKTVRxqmHA9NSEQLoR2jsu/I+568Xp5tn5oZUz8mQBHbbzE
66bX7qemp9bWu31CzeDi6HBSL6tx56JnXHnvXH7f6PevituO0JQULU/nPR0rvz6K
8c6D+oEqTK3gIRzIihGyTVCs4vAeTgLoN1Xt1ZD5NsawQ0z9vpSC8v+R2o57+kXj
umF2/0b4nWIYxqxca2724Z7uHN0rxY4jywcjIyVdBod9TnZEf0S9w/hA0i7KVRae
Snavv7awJeIYgsKJh97Y4Stv5/D/k8HS3RRNmEDfvi1VS8+Q3qaUFQ+ykj2PORbX
e/3yb/cZyegOgu9gDhPlSUIDmM/p3tDUCUUK3kehB7ZdjZSRyRygorm0scHj0uNv
9U5BOXdrE72p3Hh4gACXTxEozkLePJd6mcw61wsniGydWjb+78MWf/uFkjkICVHN
gpikLDEjnXcroRgGqcb4lMeCfrWihy2gnlaDFDb9oaQv36i+++AOESfrjRBKTdQj
jxZIgEIBLtBbJkYClC0zBZzgbuuHvWsqkE++vWmUJ7uQUIx8+c5rHyd3h0xkZGkY
zM7l/H537jUZjCAVA7QWd0CJNxLyiyE7EBr50Hd0gVSs5+AWbxTeM9dqs2yrnyD6
fwDjonaXSFcjCZFezgKvoO5bpiQdfAWrfz9EH8Hro15eTJdFLv2iL/b0tHdSyetq
k1s6V7EWgzF3yDzNqrVe/cIpXKjvgcblI0LM44LhqPzlQjLYcy0sc43OF3wCt1UC
/oA0hASGpmdfvs2odudRR6M6rs8gHjXBbjYLXHLUEk2bFfKebg+ZiSJrbh+MdSMC
S5P+c1L/KrwxApb9RoC2Rm8c6vdeckAdLYgjIuKcKzCJ0nwexIWH+TNxk6izzhLI
Ywjhkvy9uCypWWb4FjAo3Zta1+RcCmG1ysqu1sWOWiIx0QbUFGwceKLx9I8cIMae
gM4DQd/rYTnu7gY7zQgoELEbh/OhWQ8rsPZSbuwZ1jUvh6IgAQYU9S74+8fz4Mbo
vOUtVPBOihZSCx5bEDrVb0WYWie8EeY8tFIaGzXyDX3OlnHH5RXsLDXI7bgc2igR
J0OpctNDh0Q31dejlYan6JiWHY+xWmk5yq2se8vybKngZACC3Fsjj0hmFA5D/ozl
sD31GoBSBsDEVrFXfDGir+c9p2+vOnd9YAKbELtulPoNPvD7DPO+NbjB04MHfSW2
OpcTFCu0wL3EgHzxgv0cvZSSTXdx5j0Z7i0CrgUg+H4A1ZJ6t1jTdFN+IZtzGX8z
PMQEYUj91r4x1ByUUhFqtlj4zcfVFzSew0wagoK0gSnxske3amjyZHMuiJVaNtZF
u8Y6y6FSf+DHhS9tx5AnvmIlPRrK8YrBXP6bcqVuxNe+PPSA2CawSMRokAK3+mGr
u0cuEACSMqZXRcGO5tf6nmrKQMrNvVIhIH6CGtgnJ9Mh8ofrnMUgre9P1GFC8zX/
Rj6r4pRQ9v18oU+78LeVvJAXh2BkSOSShDJHEpH/FTa9pXcBjBXGDoTg2LtnNdMe
qjN+M5E/uVRKRgV7TCsbmHD37ZvNbrPWQltHW4/iYDpHjfEjGXIBenmfg8dnMjF5
Fftsgaf/z3eYkxDgvVSqtHNbRwJq+h7p0kZVjaboN4J5h5iiWMke1+wwUQB1D2eT
8YULQ27saJ/DQQ1iN7Zh+F2b4fr4QSkG6NhKuQXVdECljk2qg812k3GZayzn7T9c
emr1nLaZTebaJrtf2sgtt0K3Hj0UcJLFUF/KVtLWUMPetxJ2L1w8VPr6N3ye499C
nzBMZocmafJLKR+4pnyaqXhFcCI3r1M5eC9GX+J54+Uwl0sd/lodFveFabOZ6U0X
DSFQumpLsVLQp7Xj2r1gZmWvfh537ucuDzMivC5gEkwfi8NHf/qrOp/otHpjN9Aa
Fy7YWi0GFiZHOb2TG98RzaExqz2SbQEg/7i2vFWIiWYebluZiz979kO2v/mH+R4e
jBb67KvG3pSBJ5lUH+9mXyn6wh8N0AV76hRxqaQc2sJiSe4ZQne2NlMtuNhQkVQd
aMuJo28iqeoGwp6A0+Q/BbHzFKrsdvc0AL2+ObMqBExFD46Fa99n5NhuTXu985yF
UAAu/KfTv52eQnN53XgPLjYcg9kOvp4HLvLOgyrtmEnSVRpskEzr8JDHxkzMU8E8
0+LaaRDnu659MaSdvpGUZCYbyGfVYbdzE0UKiOVANr8S+L4h0yJy9aJ83UecZlGz
DFwzHEQU0iXpAW0ShLj2osqUzSKKxdGfKQ8IEp8+GeFeaWBRhayWmWREVKoGHmky
rJL0SxGF3QBWzi+sfIqyvUNp0wsxMs2Q9dC0+nPzJ/8gd+9raROD6ZfEORqpBtBp
5iuiagEiGCSK7/JaOlj9p/SurvVVCXiyfJVZNU8QGN8H2oR3SsZriDktiaVJ3HKL
4JjyU1LOC7h9FXelO1dGkhg7Wzwps3RLsZr31SvnjZr3vWunNuzvEs3AuF6xcLRF
/5q8HUzASW4DFUaleGOJAKu+WZH5f7Na/mL1Q5EryxaV51mNgHtUseAXSFXCcq0F
jLLLGCMhZkDy8dRtzCEqWrNK0k7PPDmJl6RqOoAMRcSG+7gOFCdRfu+6meon2YRL
nImJQlsTo8MmVVG8EONhDSnyLEblycTdIYDGWRM13bSWkq+btyE5gCzNkECyGkR9
+8t3dDALx3CxrmV4xDGDgDTXbphoMQ9k2SCisZp4Hp2NXZeDD2zf/DPQh7ycacGp
+Jx2aSEStigEM1vG8h3eydnEswJxwZvXdMJahfgSRiiezjglWU9bhtdyhfF+EbHI
UbPRGdR65Z7KCUkwoojLAbkMEkqiSU1Y8rABczLg74qKEsg1mVVfq+LVzp74SpCX
F2G0nLVehQZ2NisUQQipCsmqlKMmENib2ayJXUxai0ac6Kp9kUiHuNHGf7d+fqEr
W8GGQWMN7hJ7Ay6AexGJ031I9M97YQv/d2X/lupiwrf3ZQtd6f8Ht8CK4A18Os4L
wyuay9PNmLLYB2FUJBYpYJG24Ud/hP5it5M1Rf4oWUJzcohh8KyJj3SOF/dqj/cO
2Bry6CGEJF6tLHqgM3/pKFDE4flNYOM0PUhZxXV/dOLn/UcDUhqKjrxj686G6iHV
jbeK8cEzIxGggnexmasKursPjt2rIsSfLFOSsUTNSUfLB4SrMFuoUVgVGkpvNUCH
1x7SjxA5lMN93P+If32Q/WDm2RnVOjvb71ClbaOXJjjPK8IDdz5KIkh6+f7/9iU5
Ha8IcN7daqTMs4NpMGNkaOYNyOlWuXfVl54PzezVI1Tv0JO3pVO3sp5iiy531Nkz
mPq48jbp1wjGwiEPQo/OtPnL26601FS4CWPXj/xZiW6Pg034udrVgVDJfpbPhc9V
rrXWssFZzYt0bMQFc+l6Fvr12/MxBbCDLVp8PbJzF2w/m7kA62+oMXl4CxBa9JTP
akJFlEWyDtsoorzdg2x+1V5Hb4Nqv5kwuw2K9p2p8lo8yr1czvb9b/FEk1G0KImp
uBW3RTB27iCb7mvSlbQc7cRy79LLHBknaJHnlT4fcD0YmX++LLVVNTbY7Zz9C0oa
lsjN6PycLH4D8qx8g8z4QcVNuenpPYXmsSrq/djNFPrUDmxo/18dlldwfJmMuWPo
wPJuStH3vNwUU98Y3Iu7Ys1PiaRV+wSo2npw6KS+CP/WOubqSeb0jucuXllT9hSy
cAb2oKKiWD5rzoZxlmXp2YNZsvHKsArj6ieGhKhTty3VZ4pR6yfQG8UHhqjh72kz
2KD0NG9Y+vCJoeAOUGYS7QXYYFEYZtcedc7B5ZB9fZtaXNYA4w0UYGVD6XNRquvK
WPZHdUJAh7XlYj6Ax2XZWfmCDE5VlMl6wFORCyPfguSiLFxIaaH73W/KSJrGVd0j
wbA2wojhUWxMan3omA9D/PbYF82z6ZMr2HBCKdbSaMEL0ioHqfdvLoFr2T3mAiU9
SdVKvxdEVVeNEI5yagMDdlmw1BHEp7983WH1yVE9L70sXLSGbaMflU0x3lDqm1hp
Xi0lcUUj/qBjlXewkX6jfz8ZMRuhKR/N3tP7ZmscJkTwQSMuWewzJwwZA9prbDCD
XP4X1HCd+7uX16/JPcyT2Verya3shTUwHw8wAcddACSIMG/DqSXzVBk4QTOkL0zA
eukdQZvUAPb13vzP0oe7d3X228X7Oz1LJ7ALlXrV8hfxYrH5bJTttrmw6zf1l3X5
jiwieUDJhoX0rfqv2J+KnC/K8OqJtjFcLhREuR4MO02o+Ug455NFpIYIE+w6kM2x
R/XdL/A1tK6ABBAfjFcLpEMOUoyTYsz3iEp/cV1Jc9oVyxKdMBqf4s4e4nZ4ROzK
YqxyFqHvhSMoJTVT1mo9zJhMt3GA91xg2vWe4xh7SwbliLFBVzUa5fxeRvqYlHxs
nCb+5qMb8B+QCV2HoGQNg/Lxc15LOJZONz5FZi+CoUpctFPOxevSfMNr/TjxjC/A
xW6EzSBAZd0dkBzxCfPfUWjF+YMMWoOnm0yYKmpxt1HB+mMz1dqsEL1qM6UhGT3Y
eu4LnW4YfDpQj3uN2q7Pl84j44/AcPVnNB4gXDvtGnQKACgKgp0tEeP7rAJ4EUYX
0roCMabgRn5otEV8Lw6Lb5w1LiHezkKSbaoMj2VxjlFZcgtzNULNpQDZiBL005cg
rcmvXoljncyfSt3F4OzJA/RnBK4dDSgQpYt3d29MPeSiIjajGtHzSqxGd9tl7iLn
kK9oIgksSiXx7GQzMP6ME0ULmQBshonmWkJ8+jM9Trk1Qoff7VBc9oNnRm+dPEp9
Sy7IswApEdOiw4AyCV8qWLc8kYMuj9KmX3wj40Evsz5OTaQmFterMcgzFlhIMDbC
cl83BTMc7YHW6XqE1/P5uMHmxwPrGCE9nghm12J2BOikpHvE8K6qxsWgQ1ZwnWkt
TE4mdiaz6vKDO70l5xAOBN43jsGJ5qwfdC1cheYh6nkVIqMDtZXOijS/VfjT76PX
cmx8+vuVSnKDN8Ef+DZlbCEg1VAofJbqMHUqv4rW376JwaXcoEcdCGMFJnXO70F1
bEKNMfKJYGueQiNhHI0mWkDjIuPxJeEnKtTsgY4d/aqgvrnfMYGjTMhfGhEeJWQi
/gPA8b8OyulpED56KWMN6P62TN6fn1mVpfLR2NuxJxu4utGihlrllACSeYxeapUE
d7+c2q38Ttr63/PYpsUgu5MsWKhYqMme0S9Cv2PIek1I2ZTCZYtO/Dsyab6ajvIh
jjHTL+TIGfTUkNGHY6vX531xlFQB1ja2v4XnjE4FCSgKgk88+su0Woj0MRROdGsV
wydMtgL3BnpPA0YYRtTFRZxAO8tXRVVdRkfezJqcXUNrof3M4HR7sIgHUGBdaFC6
laTxDiD9Koc45KG7OnOxZtmsh7KQ8aCXPIw+VGovq9qKkMGKhfTx1PCu8h2tEWL5
e//aOCtEbzM6lKId0aXCJMV3Qp3o4pZ6uroZfCg41NsOdtXAb7Oq0PpgsYudW3N6
l55vyI6L+b0CWBHfP9yGqLl/vtOA7I2rhNJur5ahmcZs4DzsqCtBhCeUHwrnPii6
CVxDXvIZP1NujVwR4Fp3DNJeMd0DI01xfoFeMt4AIUq6G5fpgLm4eKA6HLUeOfbS
xS/T1MKhFGwTINZ2igFLecNGro1y5HrMB0oL7mD1Paqno2Vpc58kFDDbqqtHI81m
G1JDpn+h1MJ95l9TmvWvapbrMNQAOPuVx3Xghn6LTJgcx3+/fCkBSHerRH7e8Zmw
tex3hmPphMF0eCt/DkmR8AOoV7Dirlh0BYJPXGOypakBuNP4A09gIkKjRBC72g3g
0r7oxDdLZ2Gxb4gVsAbCPd8xJKLASn5spk/9nJtP5sTfGm57J+r20YCrshvAGPdd
sfwriPcYhHnq8UgKKtTT8Y0KKnXP+EorfygOutSk9BXiGeMO9LYbCXyZkGh9LMPX
1FSmC1PLVvFiEk7mAJKJOT4sHP1+94oeMvkDNKIW3+vCXC+35zyzTL1gltuBDZJH
qZnfgZoWN/3hyZD8H558pT6/NIBdVnsObW8tHLkOJ5ALLDncCcWfUnOVjkMASXLq
vtsCh1PtIUqIbXYJR202GcLAFAljQHVqyRJ8iKdFFzM7b8vihLgNYsa92MtvIQed
ss+ULBlzlzTOx+kB8lckrE/qIFF1H3Uo5m7QAFPWpwAKMWnxLt1c0CkKhKqMRJF4
nf+Isu632O/D8XWH+UlR/HWdXYnZa6yrbgvPApmOANn29yO7CM+dqs+ObHcjl9zF
YO3TAa99/4wwGHGMw+vhLAseDcab+MmRlfCwY8nFUEZVulUwlUN950PQ9E5Dd4n3
UASrv3zSMgz2DgDh2ojbZIZc8xsA9bjLcFzW5xCTifoD/WJaxY7OhoCGTsjeJE9y
/M1PGOcx2HSJvelk9PYe4/COawb0j6dGpNR+GJPZBqBulHsMPcHX7EY3bLgCANSN
X7VpsFUP/G+0MAYnTTmFXfdFS7p6JiRF/zc+e1n+JHMByGuGRM6E/CzWIAAmk/uM
wNw9WCmLbz0yHdi4f9K7UKVBYp7BcMffituo+LR+i2KO40zcivseR9QzSjCmmh0Y
Vh8ksqjpbc/iw7N71dDh7UnotbzYHW+Y0392VmeDEAvr20ejuLg+qpx6wKuLWo/K
7L6Qwr75pcxYf/WptIc0MuYFtjPTpdbzdroa/Ve3EAYjQocRzHcP4Qud6TM5Ioyx
WiyZqB6nr3hWQFoOsIw/d3ew4So9m32sW1Vu+mHF1cjwKtC62mO5diiyxK+6cywE
LFyISUGkZWuwfXG95g+uNgOhm38P9DulgaHHXEfacrSzCxpeD29CA1CROfOAuP0f
vyG4wNFbnUA3o2elWsR3fVFhDtHuklYiKSW4lndnRSwYkKSekOIISYcjhUmd4c3v
sE8JHm0tniTSomZ0LkHF2Q7A4jB+AKjW3xUY5SPq3J01IO6omgWQDkfzHTnWfenl
1B/ZJNFJQvNTbuHFm3FhEUdUxFCvZD2MUbgWX262X4gITTk/GqKcweWShOdcphsF
GZb3RvxQ9dIUanZsnD11Q/2eEYCu3IO7vcmuRN0vxKPa8jV/njUsTVNcZ+t/6rc/
q6N/WrpsCfZlneoUsg3BxNXBhHlHkuH+Lu8znAnm6CVZKgf+co/XSjdhlZ9jx1ha
c8xof8G+uq5nUwBmI5kuGbEzRyYuTaVUtDxJZFD5TjVHUP1BAk73332NFK8VRSKM
8VBReB5IYDO5QeRC/D0x735vP+g2t9PXfREZ9Ump+4t7mrtmGXjsQoNy36CnJ9Hf
zJ8oy39iNh1FTRbotV31hRfGVW9GNRBLt8xBDwdhODw8nps6aX5ypAB7HkZkIehc
nLHWWgcq6hw5vvv+QY3pUjfLt/lT0xpakAYYzbXsEcpB+EGjr/mLyNcqi4FOPG5c
lQsb3EKwjsCbXlx2YQfZ0uXZ1nEou/wAv7CTxElMS3TOKpvA7FwHxy6xwIbfA31K
6gLg2UszKPLLCDcChEEB6YcVo7boMKDXll3DiKDf/EJJHmM9kSVjbnhdV0aRE/nZ
kIvP1+klGZnK2NUR8XFFWn53ksRawgclau4Pgb5Yvefut9+47LT2HqMZ90aRiUlo
Lj7gXE71RQcLE2PD5F2Hm5zLHAlvp3vhYIMaHqCjU7c78NdU6F47qr8vyAkv8bvV
lmUd2Re7IWEI4Rm7A5N/r7xTSb7lBO21+uT/r3vOus+LY6F9tE/VMSZBPcoob6Xp
WOBW9xGrc3QtAKKsEdpljAGkr+4bsUwA7Qqk5HZSU35o0OB3jXO9/Y1NMPMrAA2l
bcCiHmrXySYQrkVjBjovAK31Gbe4jLdg9l7YeqyWfMqTWPyfqBWrlnUfDWcz9ioW
7ej+mKol9Li2fLQgE+IOVi2Ovm1t6LffcwX8EX5Aa7KJC1+HQrE+bTgk+GtvXhnN
AgFb1ev92diDxFVutxoJeaFENpljj8svlnhY/06CJ9Sm6NEL9SMVJOE/rjbiZEGG
NJv/eERTlXpiBFPK5/aaj2IxIISjX0gzvUdlhEqAg4s0MBaoCrxW3Ejgj2upUYuA
AD6qPSII7Z1a9GVguGr6fWpbozxCauQ60EIm2hQfNd9YGWo5ZK+1v/Aj9G7GJdaP
+rNoDqZyyYTkRLiHNRrElGKRn8fRJbF1qwEq8hEyq3Ex5nbOo11hjRZ79LNRPATI
IyhY3TaRDeGDIsv9eOoRJtSFb1hV7SkfhCsGXF4/FfdTvN8IzYwb3HGVu4diNjlC
ZtpmwqoKiWGHoKolC13zN2dyDxTyXd604Nzb3UbMkT4cuLPMnhMuwsnNCmSL4slt
KtDG6EMY17GndjNkl5/yiNEIqmK59pYIuLwlpzma1H/wb8T7rjU8HAcRmPYKYflf
F7a9SDCPnSHywuqGw2eQvFWbBlFqOMdPF8r0J4OeZ/ifwSDwHv0GklMgAWWSmXEE
p6spcyB3N2nvD/k5THkIAcxjyFaDraJFELj7sA4Ex0sXPQpHGFGwilTOpAoDyHcH
sr/iwCVUe+pdPV57aFMlfjZDTkY8Jej3QdSBtsUOhQkVNVjsETgOqoisn+NlnWmX
dg6KXw4rpTJJTSegTzY74LRvc+U+hbgEfxQdzzu9aYkJxG+r61j+duhVIoy9+wd5
f1G49fIhvtPCY/StxIw4wHHgUYD8pvAx7mJVPMSkxRj2wwnpxt4/Oze03GmLIJZX
Od/apvxGZLuwzaHHZZN6vtoiLYyGqUC3S+XVW8ePZZSXj/BE3+g5MulNpXgG+Urp
bXU/+PojFeGkTon61eUnWAYmQkgiPL+UDcsp3/wzVMjPDUX9KK//Pmf12C4cWsbh
GoJvfE9TmFINPsO2H1RXlB2u2e8ElmsrRd4kpsebnmymmPoEZwxH9S1tyEUnozLA
/i8ZDuugfDXiiz7KS6eIBZN4fm1Xz9E8j9RjjUKfp0Eg+v33fPcnIiGRmQrgjS/4
8v/zB17dhJtNl+TOAZ38VtqXJbeGz3o8SDfg6Reg/KXk7EseEpB5ySmGQRS3S+64
FI2BpD58kiGPQqdiUCHo8OH7shh7Sfs0F5C2D9MZJuKB+v+YdxuZp8KOQBmHoYf5
DLH6EdWVOUE9l46E++jMTS/iF7Dp9VgVjXXogrPdoWqmXaLUxmFcmu3sAxQCSvnV
yp0o1oVUFhxI2R7RIL8Y1rX5L2uXyBhfKJuTcKaBZQrm2Cp9D6Ifczre0xeKaTPY
LMYcsTv2YCxoVK42CvCvYBkKET/TperWeMiN9n8j/kSEFGQSEPfxZSTdGodrKium
LfV+zcMWBvlGimW3UkCCCxBqgVoiXg4v/4tU3t0QMkRBgwxJjgZ7NSwB0pHeCwPu
ozxls5XE0+CdT0IZa1X/3xcuP+A8E74kFaXtrpbjae3HRzG0eDKct6OZSIUO96Ot
JLz8pDjydLTYUE3TNv0lenm/u3OHxEf3ko05kFGb5QkUBHGc1ayDEq7zx93ZXUdg
WzLLq5HKz2BBFn1UF0i0JDREEHKGNYSyEhjdow/xB/RsO0+gt9MBa/KY8JW0Aujq
rV+Z13wIQ8xw+pPl3+GVUjwYwNpRSDKKfEiHkjy/eYjJrkxlVzjU+sbeVgne2Cru
X4LMwvDFP97GYVfazAAEnQt9cCEBx9joASqmsrdHygLAX4kWSa59RI+HIIozJzOH
KKAZTstz/E3B3JNsijeWKk2fruLr85+fDdHYW7T45Vrvj2bkdBHbqMHoZrDU4f7i
tvKmITkTlTGKF8HORQjcVuzRSj8LC8OH6Vt9lr+VxhZ3cCawxrDMZQNV0QQnRFp6
orsoRMHpf37WUhzz6Lz8aVZBa7jdX6M7pJwlju0azc+N5OWyo61YDRcorPkpm75L
UtyHeVO7cFjsiyaW9xeX1k3uyHVF22C/4Pp5KE61t+wFQgbDOhtvir5ekmx/n0i8
YvhiZ7ol2Hxa/SkMdYJeu4o9hcWAP9YMAhI5qheLeacwpnNU5w7RGcv3IdyxHTd1
hTXF8HgP4fZ3OWnx2QwuvXO2zS0Kb9f0XwuWqKOeXlverlh/0APUFWZU7Q3QSlNS
m3F1QabSXKqeZ38ksrERE7So9yNE25PQqMPWOd/7RzU0oMg9EuPuXVONc0Wq1clX
aeBG64l3OmDFARI2hIQ8VAUkWgi/IdJduKUmzM4EUncwigDzzkC72GDsOr5fl+rF
gzsxefFCDbUD5sKrbJ5Y7WQjqdAHAXzKZm4ai5KrY2V9I+bBlOkEcZe86/mxaS7Z
04MaSBDpgK6KzfSNsEfKWKqADIXvgRx+AQF+G/w2xJd0xYsPNoHEE/q8Sec3qtWU
mVZQ4anl/wgdLtCghT5TvZ4xAQIRs+iv8ysjkeOAG8vhDMD8xn2ayuCFtMuO9jKj
lW3Hxob4Nan6wPiT0xaI76Z5q8Dury6ktraTg29HHes9OhRzTDH9pC6sq3SWKHQO
L1fkqqQAN2ApQAwkAM71Ujfjz4B26P9u3tvxwpoG4CbLUvO359z/2l4pK4OfMuDo
V6xtoc3UUdDUqsmK2Ant78ZRm8xBYqGBnFVaSBFIUrg+pZP8HvgJSi9PqlX2zEzz
12qfrnh5iyX54Lyda5iHQE/QhUBZKfy6h82fT6Nv7/rAQcOkHXjg4tSIYwp3GvcP
UjZc8cOWkIYNSOgkZtSVlyhJpxl4XTZEnsIgBLiJ/hbmhER7GL9PXt8h1HiwvC5k
9D2WCsjdI78By4ixdY3lEWFdLqjjs6HLhejgYBHC0uMvtx89CY0jMj92ToN0YSaE
s729x2071jF01+qxUva/Yyr5yIv6DIxwmh7Bt36smgMu1DwWP+naLTn6pXDCT1Mr
jfGYvI8tZ2ig6zZMSkDU1WURFda3z9c00UQ9f8tRkp+MJSPNsYNr9K9h9y1R0afl
E6RvnIL0NMQzesch+hHV7t6sOS57kTih3wkh6+IbT5QMUsJ1ZYZ4UcPyn72S3HOr
eDrmHOb113cMHVByFcSAtw5hqVVZCGpvoM8QKJZBTAgf/4okzL196cyvcHKhOkJF
Q4UuFT4JPKbhFW2pdiStZbcgRFk1UxgfG5IZPrGZKcb9Tr8d8h6lsJtwvmIWnwCS
6iNrMl5NuObIsjmMHmgEX489NXQEPhdtNtV8JyNY4AAuxOcqScBGkSEiOkh6ZoUy
wpVgEVyawEcVwVQ8aLBVz1YwEuFFcnjW1hzwtcCXDGG+68KduSNRd0X3gK7DS7Cr
H2F//Sq+mEsJkqcoN583N29//fTRrfmmKhvIVlWAIsA7uWL1v1cERWP0xplXspXY
LNrCE4Dw/QgOYqQKQlFxLaKQlEWFGvNBmBlipDVX0OFWoBT/ioFNHg5c4xKW4FUO
m9vFgCQ5sVf/rvylXB70kSZznK2Nv03/4pTpW0eFSgkUrn/cKf868sKsmL1af/Ry
cQXBvAfXXPY7u3TO3aHg45hOA/4avVuTh1vDOT/nl1Ljo4WYJiP4qTV03cHEhMQK
vR336tYll84Vfm9aXBoJNWxmJeNGQo7ULmHtty5Zoucl0U/JwYqKUS/71Tsh7hIO
NtIXUaZSeiu3NSxECc3aTfGd/1nqLYsb1hy8PtKxxca/BnMeEgO/OAIoJvbYmtX7
ba7uMRKlfeXH6Xlx+wKGyiMdAjZDwpUOQYZkRTgcMgPbQnNztKUGY8W5AeCmydiM
IiNVmU1v28PoiRkZ9UlZ8drzDm9mTFZnyMeTsQjXnr0RCLM96sEX5vFZvdYF07tp
lswfOQOIhg8pCPCMCmSyn57omWySTVDi04v8PvuB1c6i36b5yarW27ukrW1qClrb
k+ACQ8sPu5mu4spzB+KHQG5B8jBKpaD+umw3kpCT6lSyVZe5kf5Gu6ZVRw6Gxx/4
sGiTZFZI7iBdi59Wxfxwc/cS3UMLwTBGtebNEvqBDKWo+SJ1XDsoPJhrg+Ks56pl
fXboy6Nv5nex0Q+JXp71NedL7+Wi+e2t3CLLtVI0/fRC8p/e1Nfg6eSNLBZ5rqQ9
7HKnjGAAT8RpRDm+YXBAvALt3T1MIr0+qUImZz5XQ+sHP0mHP7QSvAH6yFD16dSl
7HdxMTo/7uV5WuHOO5PQQFkSkO954pmkuCdXYC2vDaKzrM6Y5hcq0uu8RTyl2XGD
Ek9mLQ471cDPepESliLsqiiOxU1kfgegx0SmN94WYJy5LNnZbWeRWwZlmHuwdzRT
20/Z3LV6tGcQjlr4Yo1FM6Y13BU/lSlR5ZPlwf6R/R6rPdXfwr66Jy6TNjq52kDv
5Tdvs0dQfZrQEqp1QwA5Piz+4mCNuuZ13devkHqElepSb2lYRVxFoQYDTuOfvypJ
uOFPdF/9n5ih6AuSMKMVi4mkUAhkFRySaYFCeV/gaJpI5Y3BjIO858pHaWUAJtj1
ttNvt3ONrfeWXFcS+JJ0OdXZt/Lf1dl81JRwLtEwJDVh92TpmdPyFg8xxEi3pWvE
wLIbN6B2SRGyGd0ArPhbmPVf3fZxRoCODYXYdwozeIaUyxH1+Q+J4QqXG9YcfyU1
FBttTnktfHSr7ZOVDTqwfLEvs8l6712VWeYZqoFpU7Sbhe9nJiyp1zMjdDdX52b1
quQUqic5843LXpQlaF9rHB/Lqxz77LQrLFOH/jzBgQZw563hFqluYyCktyq6ZrQz
Ti2Zxi/clztgneGaemcZesUDbNghXaqnygkRtJV4lEEk1WwnQa/NmgnKqRJnDrJz
mWUd80RB43EM4tgTuzNzugGpaTHFwfYIQzpLCbgpVInPjAa9zucNY/mmTlUC2KMN
6WefkCnH3nvF+nRD8krQdkJn5SUeQv9ojmLWzN6owA0zyGTIJW3f1L5dXOuNBCuj
kjn8zjQx03eFqfPdS+Zr/HReN1KKfHzfI4PzsJjM4D4V4DxdQtewuwBtF/6p9MyC
zeTeM/zTvVHpkyYvpDgdGNO12SUX0H+MUN8OCl/GvcdL4MHofg47xw8c3SpfRUiu
/CtsvWqUPgGKuBbx1RixbDRSsy0PkdHOhbof9paorv4BV9+93Zw/+f83lxzVABBl
PNXTFZQ3qLmlSZk8QFmFVg6SnVM6L74JlbuyjiOF+Sl4Nat9Z5kxOwvw6Ig1TpAu
cefxErctv2LLaNUXn/Wxp3C7lEFWEK0LBAAYtOKxAxX2fluMGY1DXv9H6do32ex1
pWolsRhZerwid5lPaAwJ/gL56SIk/BIzyLS9Lpt9xB1hz7No4FFDLlhkdGhlUqTn
OseSAwWDEkmgsy75IRIt8FTrcACajxMP0kQtye2SiK2nauRmTiJknH7JoqYPE25H
hfH/4ggdFq2dfFIEP7LTLfsTUlk1t8xHZSq7ppBEO8xabCzzYQDPgrBviD1RcsBG
DKrYadjVumOP6pqampz+fRpltsK6o2fZeXwNr1RYTk550tSgY5gowlWFyho3Bikr
TahrwQwcWlXbZK8vkv7dUTGCKr2Ezi/qiuXCuN3/lPjS7PIE/46IJYEOQBZpWoSQ
4fXw8uw1WfwOLbCnOzLF2KyADD4N4mBCkahWPY9Vovcm8lr2r0ZPZNaDo1t0PIv2
SSCDm0MTu8mv6ngdOBWQYdfdJJib702I2Y7/vcJGl27hqpBiQWQtd1s+Xh0zFysx
iRu4ygIfcM0rUQN/dlsWUUSBVuULJBV3bZL7iJmK3T42iGvSI5mVw6jkJJZgXJ+j
yZQcYUjddokqViHaLLIvIzs0JEPaMQbBtZafageO5I0ZtU0fGBd68tNKxSxXvccP
tLyEecbdzvXPQr3CSOsYKbfg5fxkvyjxCx+VJ2IZO2UOuWeAPR7vVtM8lXBCm2xF
aCOvQfciQZ5YHxyVufKr2HIX00qoP64o8ytTOmo0ftAWLGaR5sWBotK8mfYmuwwi
QacqW+ivQzcTrvZzTwi7P2GszlYppl9wpdGUOldP/JVHwioZf0bmaoc+s2TEuuDD
B5cJp2HEYn9S0P26jkyFX/jyRAZr5rr6A33DmeMIq+K2K5uWCYzbwcpipN0A0PFF
WF5mzCk6xyxm2UbGQHvqI1ffx2wgvgEfJ/eMM6g3cJ92C5+o6/EX9JRuri9UAhHA
olnlUVfUY9uQ+j0+dYp2jFd6X12pJjc9hXY0F9Tzdf7mLj9zU7wsmuBrR0WAl2YH
pczzBvTQZFoobKhO77IZSBEaiuGt9W8mapNnZzBks6nvcemW0cgTZqN3TD+07vZ0
ReW3/QQCphUx/BCnEoYVtZvwDWbMO2T0pDFmEKQDJ/ykmij2Xb6ARsQUIvUf5OZD
JkqNSB7ZGLP6LIR7+2I0EkoRo4hMKUKZQ6kVfpsd9KfJ9u+fHANPliOl/oNTdurV
WZt/G//BKjmvfy9G6VnxAheCzi+3gTWYuEkHYfmT8xmYPFpmps8gVfvP+kTofat7
z/kEyHpWG77Ef9FEz4/xZURB6HcLwOpro2xCBfcLFXvIP8I8snY6RAGxRJLhJQea
02wW+ldoYWSf/7YRkLU4eV6uOJftvAPq0zVinGjjjGdCUmfYCfWGrnySx+1WbeJc
nSTtS8Sjud6XC2Lao36OM6Gn/73W/L8/xqZEUmeMGeQU7stc62XxBxK5mhQuZSZU
C5Gq1EUeVlqiqWa7R1bILlhxQ1Icf466kXF7LA+47nBQE2IHUPolE4ae88KoSL1I
0+hgMOj2s9G4wdq+0ohzSuAu6/g6ZxZXkgybenI3bio1V4zOwO/L+QT4z6L4ZHmm
qMh7qmRpJd0jfbylXd0qZeS0/junJTGT8gaxhMSc8AcHaECdPSvhGe2ETzkLsDCG
Gd90/GHZiRVQblx8gqx/ruLpMlXAN/UGplboPg7gOBBw6WPEnmkM8Es8kAdsKaYJ
ul8nt7RaGQVSQ+f0zgMDx2kaQNyG31oZewqqif02ldxpBDKmNGssv4aViTLA1dX6
nNF57H9/p/hiCNfP6Kjy4Mfce9n6IaEDB4C0OX0Ub3dQLGclyIp9XfkFIuYeMFZr
7z9FJxiCG5ep6dhoDNB61Duauz/b1ZwObWoLteKajcTt88GjIFPVKCCYZB7sO4pG
54aBSiQwTmWXnumKOsbY2f++wm54XOGfluPY/MSckQIVkdaqfzu8IOd9gOgTd8UW
c1Wfzev49Bo2aXpswY/EYgbuDhixpw/CRQUfF1oEXZ3NtSXCflQUK8Jd+sRSkUzz
aMdTYzCBmcu4kKi5s+OMD7Ao5rEl4wMdYzCP5VEH4YrkX+5b9tTK8DLdcIajKCX9
wMAEuEJ9tmMUeVQM+OSog8T9m8Liz9QW83NuoXDId7UHwcw8/Ch8XXz+84LWs7XI
u8AWgh8muMNYC7cgYz1+KaRqeQFEvd4sFBXvFsZ3WKgYvClaTjvpjOptkrHFwus1
zWUYMCKh7K0aRhGuFJ4blx+GTzkbtFu6hqywW0GobIKXc5S709lYzIV4AY/2VCxZ
OestbsFHsHSowzAZL1abfEDgt8FFPfD7b/zLx56nvxIEu9hMDR6VWvIv5tewDL7d
4DkuGYfqL0M6krbteNoWOHJnNLPuwK1f9DAx9Ebzp3wxGacWJcLzCascANqAyNzp
b2nkqc5F56hfjF+sWNCie7iWXVQFKYqcICPkl+5Q+1SnGVcHjvMeuoxRInH2Aul/
936aSrwoiUXiAEZqa0bKPlHWeiwk3XJQFnn2P4FMognuccURk6xWW0u23nrNeXW0
KtVnAFg7SmrIzNnE134cQp6Kf9beSOwVsDmb3HOiS3OXc42byQdvV3k1iVNXSsmr
2SN32FRMsc4tTgqXC0Jq3TlRAxTN7wS6U9JZg/5i8p0OrUSsKwnXbY1MEBVWlwr0
WGUKGb+FqURT+LA5oEHz4yFrkHOSLjxP7BD8Tm7UMPYd2U9qz0lMDUQeBtAKMCIj
hRqIK6R15OiKh8jpyEAg1YyNEfvhzy6Rq7N+V5dfwvcy1ebh524nSi6VSf22dreJ
Eo4iZ3iLpqVeAAjDzZgXIXh1K8Lkl3GZ/a0+b60F53dE7lMAYkhrxpjxsWWzUd6g
JQ973/mQMPNBHpnnjVWdvpdR0RGNF8ZKtaXXTZbgO4SxEtUQeQL/oHn5Vxs5+qDr
gBE9aj0hr4brpVhtGZBOBYo6lUjEech1N3TLLQ1bQI+r+KeqYqCr/7KaXP1HN9YI
tSAPhviSwwzox+ez/tgbngprXDS74bBT0latJMToGBGWrKRlFYkjjyqqeSDfpWst
hn9dRw+Pcav+Plg3t9xvkAfTyMupR66hlDiNh7N9mtISURxeI1lXrKbhmsD+vg5J
jBpHKh0ivKYnfJnb7aLSnyb5gNzYHodhqtveM8/rrIg+oxCGeXv9svIKTLzF7S2n
BiWwrBUykzk+eFeK4Wgz8dkd/xIErrek5JNY3Upqz9VDTk8UL7m+Ah+3VdQvzsHT
B+3Szqv48Uxb5Xogz6RsaAhVdJHqZ6+jKdbQPTwcYVcaAEnyZK6FqIEFpUA/XqDR
fV1hjgZqde/R7f6oRgfEJ1MC6KEGBm8t/CX+rr74uISMYard4eK0NehyHkhX0Cwk
TScSljOhYK841LMNR06AKG+r27A45xXb4ajfFUCLrNe4DfyaR5WHL2+X+cU76iv5
I9dWVPGMJroqN4C7c6UmLToQlrRl11jZI6c3QNoIMCfCIi3QA92Cm9gg+tNval8V
uHpct9ScVEAQ/GTPaBDcULfcQ0fEt6eS5uR4i6nPSjVZGt41/IEhVy8qkZFJosfw
SAl4fyFe6hFID2EPwQ+e0y05TVAluY9c7c4DeGqYEv4iAlin0X6HCfaC7XXttwvZ
nnu8fYWPFqs6krYJ2Kh0su9/5SVQChdF2FLcpPpSq6lpZBbN6gRP7dxFVtu9N2uZ
Q+uFWlOG3ug6iK6BirLYXyvjqZpnM8HqsXCSzUH8zqAB8bBjNq8szEHaSmQuGhBE
9z//8yif5f3E+r0oUqLRDC0CzgOsUOEpA7gPOLtQn/bWXOb9vcdo1Vc11uDuHgE1
WCLwYKSKS2VK741b5C1qpApFjBbjqIcit4ASh0oJbieazCtiUJT+rfrup9c1c4ov
J32iBbwGPmeb5VIeMT9eFBe04TIz7CUaX8J/hkUWa75FL5b2hDCxHCas4qQMegtA
VJRLZkzK1+M9QehQSCPNl8apqoxr7cf2zUoBk66PbnD1yR2LeF1MX2m1qD3/tGQk
Mw5bdkNMy52wuB0kFadpuTBl7PJUoKnPp2Gc60XouVpaAMSuXqOEMHg7pzy6rVqV
oIMH/j7o7Yhs23YkEQ4Y+YYf0EFkN6JNySi41HE8rzis9XGxVyOPDqtaR6YtyubO
OdwynLJfkqzSU25kx5tSt3irrPVqGy2AHtUHTVEcLGfNDcvd2B1u6zT6E5jGokCf
AO+sooLe5B/enSF5DafaqMCPHq7eLoM4jMn9QRNUop8HPm1kWiRSkha7vCOT2jrw
KosWynduqfKwcHMeZN04cf7XLrB5PW1fZlm2m4Sripw0KsrkfX2H0cram+YE1Ql6
qeR+2NvSyWCXq9tdqWdGBZZ6bBIlKJYA+I7fuiTWoj5b+jNeMiABPtVzVCH9WJLv
qzk6rzakFf9gZKnA7DMoRL+OdsB33PzJ1ZT4Lj3/2QAKYNO8nLzxeBFnLNtP/GxD
kHUQLlvbf+dUkEOg/MAhVVzJYoOoOcn6Ir9i+fersBFQNlPPkRBcm+vrLf50vv9v
Y57+7WtmXQEsXCO1lTkcxFfdQgEgGMEwvcIulOs6MEs9vYlJ8DToxt5ktG2a4E0F
ITqT08FOmTA2ktSKBGrgYeY2dPgxJJCo+UvLuy6O7YGZVmqNwiXVaf6gvpFAxWBu
Mk1+xToUzfQGzVjubxcA4NU/sky7ujSAM9Bo6jbDBv6vg9LAY/YVDa725KIZrzjm
zf/VGvXQ8XnI/pzSfesd0E6T7E+Hafhx6phPvL2CcFnsTCsqy/5Tmb4L5ohWq7aN
1XMoGQi4He5+7Mvgt6gAqT2JBctLOO9+Pe/cNynMy21bFkJw5JrafmOArq4iaX8I
ffpaU8QVN6PsxB3Udw5jAO1YlP5em15AkR/I4sLujXwjkhTyKyTzDI+VeNuMd8Xz
aMePaEkBnEyxn+huH2W1TKPVeBT6VL8NmWjKjnXQgoiMVosCUT7AcnjvaWw1jnAn
7RX4ssBIL9cqVnTkI7Oq7eeJ0Wtl/9Ft6/ExT3F3+Pm5ZFOWPz/rwZ3PvSNGam9r
kH33J3YJrRazsbecarkngaVr89FdniwCZ8JDxrNcHAFtC0P6LrQwfDcHkzWFLz0t
AnviswSuK/qQD5UCWtlpbXAnvRT1ttKON5XrxbrefOdMm58J7rztnpBuEuY8jx+s
xn3FbPwmUhOrl84FczvY2dZ9FliaPXYG14NG/UD4j4HGjGFNE1xpEvNJauJVXMkc
suaMGVR9GWN3JtOqQJwvsuI+4QxWfosHox0LikhoyJ26O8nLDcrG8oIj0mlm7Xx4
/NrTKvrWW1AT5RbL7MvnN2/PlJ/Oe17bCHx4aJHzRlZYo5mDB/M++9UNPKfxIV53
YZztosy50La9NATOvPm2Ss/hapKgiCeMWEIOFmNUh7qJJiovuMxNiS2hC3OaZfW0
OGbo3MtYJC0XJRmoN5TkiH6rxsDG5XffoqzZwp7uO9TxnjnkaQNNwyqPCcUPShRQ
JaX7Uu3Hlnc0vDI0fYuQjJ9okWb2oJIO5ADRzO/31BxWfJ2LHGOTUVQcyhIlzCZT
jltEpjuN4kxItAJEBp5FtxeD23ly44RWtCuFvZ2wvKb42yoAuaWXOm07Ff+Vw3+0
8/DdYsszF+18S+UMypT9V/KhhdbGnXqCNHAlu0D5J0pIx2ApuBGgEAEbGH5MdpEF
X75yO0HQMsgejcXN1zc+iDfsQCmsfDwSwqHFLVN/m3gPyx/ALqSFJpEODd+dqc82
S9u+RsxZRqEmuacxc5BZik3dfq8nxZvXsAPlpwbDOMBSKylsqUfDjWM4ZxBqBeoj
8P+7oqWKSiKqFcfqzfvcu1f8OW1nM5sZvJM1w6RVfI+atPM77aGodWUZ7uc1lDbV
/7YtzVX+5VyBxoiGTV0WhFg0B+zz15lbNC9dg61p1TK3vsEb3xZ5tWsdxDaA96Gw
DaXQwsUcQArbWWbqWAATQ2MGKvJe9IXUm58e5gt0877lrDyBdbme8hBn79OY9oV0
zMelFKWqS5KWLLFWKlDCzKth9mgMCZxwmRO4nUMTas/GBLfNICAKahqELi0X/XD9
Nui7kvtTLsEMLmmJm1sSFlPGrpy3+u0Q33LJoiKloAq4eP+TL+mDufyb8M8qLY7A
5nW3rhS4/rutCqAFJ9p88iSsth8UWDtjC/qSFkQqtb6FUlkcd8bCSMlL86Dlxl9M
Dwrj3lyf4mlc6WxxyfGDFzHi43QR36X8oqd9jiJZln2yVJrPyDRxyuGuix4daf/Y
o2mY25Zn8jdqujkuvGV61OvEv+OQ5y5JPloWkQV4HamibRUEsvMidFpqmShmO9ZR
QjAEeenHl+zQAW5t9xf1kkfND5SaVIpRf7RKO9NfTuo/URyzowOC5FBRSipNSWQV
cfj9f/rvp5C6qPTBBk4mMWF1w0SJzfwkMgpzOVUK+E1ufdsiskE38Gjlxgw+U78R
GJuK0kzVEPvfInhvk/v0OUeKocKMGeUC7fLOzEnnmg3Yf57i4by7UpMbt8NmL0LJ
65Z7KiEU2riJSnG5a1wgHUQVLYNjx9v+8gmhCHwZDobdwSymXSl83EQ4g8X1GGUL
yv/o7t9vrzLp6Djf8ulD3LF/oQ7W7JnjIo/jLHLetpkuqGU+ZRFRpr+nc9RzVJg0
cSMBYsugeHSio1rLoDfc6RXg8h9f+23o0ACs51fVhaOi5DkHRgCOWAtxicL/ECtn
2O+UN92DFLMZQwE/MjYm38qoMwxKuuOXy7pLKFsV/uOqJRbbhDgyXOP2a+jzo5V6
HKsyPI3vel2aRXtA1pNJdoV6OUMcXIJkFn+3VzYXuo+IT1IBR0EvdPRkYEBTItr7
dqUrO57V0mY4j8DR2F+ABmGcqbTuJeD+EsOS4GYR4JY/xjqbBkw2W5etxd3mJLTV
P9yHXyEQfx11ajWNvkDNt1dYULLxAA/DBNc66ZUAm4sNMLkafdCjkAKqrl4dEKgD
qK8uSeTb3q/XR7ar8BMgyQzp0ClM6R9JLH47qBl/CkYIEUnswKC1GZkVVrdicIXq
mw1rNEZe1EbWpnMjigzB2vI4bOYPDOxpJbgUOwsq9YC5Rm4KopXWkZKoe0Sy/AKu
WS++ThiLve1dlqMXnbXa2wfLVcBkOOsMo++RQXz2iTOQOFKDJ7B8KlAtYsAstc2t
h8KWMl0dWsRxacP71O+YT8UwUYlLHOSZRAZEyhM+cAmPmjXW+CUffyrNaDVSRxSI
jOk556G2puTocMAwScI4EB/gff00+vneT7grhqZM7UEe/yQ9aquFBJNmf1JlxeeJ
9u+JLSuip9fqzdIMLn+esTS4p5OXnl5+Dx8ow1MkpFN3/O6J12zBAHePa+GZa1Iu
TxYbMMTgpT6rLwh2/Fp+HsXuBtCMRwbiNbo9IUW9jcMrPMfxiSewcPLwCf3QYu+U
bnwtEl6GsIpDddj/IB6dOqIUPH10fgrwC5YDVu3Dn8jItR8wPZPkPEliSu3U1DS5
vlcGKRk1nc/+TSTnCyklkO0SQIyu6s7Mfz8n8hjNy51tFc7d3QZpXWdBv3k3dVEj
/z/SR666e7tB/7xK5d58czZotaaFYkJHHEn8xa08zWANwwfxVK7vKPt/CfQa0FGI
HohuyPksWCNNdRfFZnH+n+ofMRTp7UEXuB4OctJtHy2k1bicJwYvBQuCaj8JtZkj
fFVx3UIeEik5ofPz2lnQXO2+DawgX1/2f7zV0XM0OqyqkSN+uSvJ6hrUJG8HGlNY
YkFQJVpgOmlshpb8t1gz9y49zLvEbBy6C0tXK+Vt1Ltcu3gu/Sn9yIcengvEU7X6
dQg5wVUJ4wr5/I0oEpY7E3fS8wrqGWRjtz5cYxCZHnLKXSx/v7Ls6Nn5OJJnZrqP
V0rB3Wl5xXfKNK+ZvPK0Q3xz61KytzYelEqGJUYkEUGKeBLa8T7ls3gCczdmEUni
O4yYy2MN3HwB/hWBz4Oo3QhwykBfJXKZV71U6gE9rlBC55hZQ9XMZ2BVMruEClXm
nqJ8muwtfX9gibe8MfMnJ4Z0MCSLVAhwemf52sQADGQ1pFsp+Ahrz8ywYzhILv+E
YOFCWZGqj0NzFMmVCC0tL7GcH4tUZ5kALtYh/hu9e5YpkPSX/2pU1Jrs4Xv6qTjn
Vwz31ek/vZXJUExhEynKGhntQFPu38iqK5MpzGFM/8XrjpsR461RX3DSSuWtZpjM
yzCFfhFcA1LNjT09QVbjfE5ZjkFr6BJ0lhKJxw9YHXydlOeZ2zrWYiM6eWJHT8kF
eCyrvlJdCJNHqcpZKCDZnYBjkzMtMuwv3bChG4f3AL4Rq0bMVQRXoc5wNZHM/h64
MYu7zKXiLVtkup3eimrsv0t4mSsQHhLTz9NlG/GwbnY5r9b8zhsO60m6Ag21GJGQ
FNujZEhRFY/taNkI2m7x5Q2kMJT00gZHGSC9kEoDg/xMPygL9QAwLCYT5Hqsa2tI
hFF2oLUTp4K6vbDlWLL7SJzm6iSt+JSa8ntvClqzk0VXnWMt6jDNHqmJcSlYt/wP
khDirWBm+fBjxErDTYw0Rwa4WF2NUPS/BAthXEOVgsu+sl/HRf4LWydLwsMwb38H
CC69e3PdA2XNSkidxDDJHY3+O8GKfSDCfq2l0GVK9F/VWeTSxSdOuAdmv06Y8QpT
d8Om9z9LYOX8L38AS92mvk4LxzUuTvgc1EsU0jxt8MnMmGKA+B1oGAkugo5/Ve9Y
s98v4gs9ONpq6+BXD97mfMJx5uEEaK2B6VjpWSG2TPiqQAyQf+uXF8rLAMqwUwL4
wxcEW+NdGolsA5arDkuqg1WZOHpPJp3Zyw3CCzMj1w2C2FJ+CUsCV0GbORVwA/5G
rnZ64vuN29SgU+pTRTtlPPesVANTM1pMFQxFFYLdKiqf76vT4U8sMLAlcxkkEJ2m
Jjj8A9NPv0KP75eSSlDYzAD9hjCjw5mvE5Iq15yzzNXZzRqgT8jSsL29qmaEsCTR
xR7hh0qqwaK17gTnDOqnNo1C33pWPqryR+RIs2w42kF39x9Id8mhuHD8fR9l8dz2
zqT9sFl24sgtYaNW8K1DvhulOEbXjsI8eEchDRCrUvQDxzzQBtdOe7SDo602oTra
iqALdpWCICoS82mdIcxdIzXsk3taquY6TJiIjGpgzX3p5M1ywIp3Ihp2eqmbQtD9
XieVpfNzcCGKqWmlHgfIObomAL8MsKNcu3ejPptn/C+dN34fdGwXsO8sEB/v9YA+
T/v8fVoLc02T4F+Uxy/vW/J2dYHrgCRVG6uuE/1Z6bkr13nsXm6Y6gHjGCcTveT4
Ex7r+ewerkJJc+6lhR9AIbJbGxlFKKzsSCLWPGj0znOIF1rg2VpmyCkNwam6ci2j
UHPVmJkkdRH1qGvj1EpJAeb6KAF5gebuabwenh7wANmc3UsQJ1yNHROHLOPlLfZ5
PGAHt0CChz4r1yCnvyW55NGS+3isRsgWPkfe0oWalsgfhtXMPI9B9epwwmtHzLjT
2Of387xEQEgsQNC1dpbjObnE9F0uR1fJox8akwWFCRh9PwMVS4BdYOzNG4UADAHv
n2B5CkUSMYE5lZHkhpTmPiuxbeCtjPUo2bHyKkAYhWCrNJRHrbLFle6EkTjriS3o
8Fc1Y6RhTfd8akjYoGby1Df9iCclI0j78PtJXLcuuFuvaLSgaEmvTUtV69Qxq0Zi
mz7eHPHSUE+YwIjfMIDnw/yOp/pPYsVrpQMyfFHgq5y12/BiJZmhn6tWlaKbl3Xf
QbtLZ/vEMG0SjV/vbiu5oQULGMFML2PeVjY4MFtg0hRlyNu5tth5C8bJ02fFUH55
BrK67VFE5DWZndZYmB1kSRBZU46z2owVAFE43mQrnbBIv5cX+igaU9y2UrdYojto
3SE6itgXfL9DP1AqMTWKEDIwaXHh9p6Gs0R3Eywf/95epoo6gmXN46Bc8ofw6yAi
w4Os5FaA/Fn878rl9yTbhx4+/1QnZ+eL1N79CsxaJ3AqIx0+mPd/nfVFQQJyBu0l
tFgQGpidqVHu9qnkfJPymYs9As9ilmBQTuFZHyLTPNN3r7yHq30DCl727diw88RC
xSyk4oOaUOMnD9kxAnlLoL6GQrjMKbXi6C0lUiDKxLMNCU3nB87BWiosMOCrhAn9
SAFyU3ljXFB8bTz6f5gPee7X5BqOn8YMBxkoqLq6FOp6BCk3E1QT/UNlNtkfEVcr
74k27Bt3byNxVIhxu6qS9n6P0M8XSMuLanrFsA6t61k1XkTb/gAy3aLFz9VZ8kKI
0I8lnv/FkAX8EwwStmj48I3Np4pjlmdJFUzls6fQlkv4dLRyoq9+RX6QMBB8bbIb
SSY+rHC+skAQ9oCoIGUPeGMOP9mfeJCjYHpxpmYRP7ap50jnpi8efPftE6j3lwu5
rgn6/3bgZnQt9+9tFX6pAiRgg3Jc1+HJw2RUZHoPi3EY1Esa/fimNPvhacM2GlOH
jvMwaPdsP5npbkmbD1ErUtvT+pMNi/Inybdp3o4vmoVOT7gro/tiHdjt/bUx+xzE
d4xqoiXINvqrstjy+IAZmxQkJrPj/moXVuYCMn3tKNODkKTd5Q1CCL4kmJHz4Pxu
vsb7jtcJQZAcSVlTDsrrdWrcal54zfM3PhcGImdQadA1I1k5to5O8jSUua4CU5Mc
Kws3wdo/j095MIKh7Rj7WYIqI4wHkytDSikZWCUL18uszo+3Z58OPE6kNXF1qcZa
OE4tjvgKCpytbSw0x7yNCpe5iTECaQkDxfkMEGXSpuCWtnTY2Ap/F3dswDxmQWem
puz5tlgHPJvmDr5ah68ROX98toh+x3QhLmJWtlRgDIXpTbxE5hBC+K7U81MlfOaG
mquUOZ0oZGGGyYLE8B5HVBlwHosdEq7RIxAaYeWmSSsM8dAyeJnn+3r9HBs+LIMQ
fPW3rPpemnAHqd3jGI0rVbB27JS3USMfMmrRZgRlVfNPxIBubfx7o3TzrWO8LleT
BfsQgDp2uBu896lOv0uNFDGZrRBHdmbqRaCPNHBvT4Hs10x6+Jw+Km01l/5hmcHz
ZImHRUOcG025yhs3h5eDwGO/mifutY1GhdtHcfEWA8+t4xNlCj7hwL2NWgserJ5f
QIoaXhTfvHxLsHjF/0m66WeQUcmHpkbj0keJh3/I2CzN1GjYgKH5si94z5t7jAEE
bCNjAO0rMD3IZiEVgBykshSLuJlL3EWztuZIUJVHd4YuIfIVX3cKLX2ueHI6n2wm
ZZPepA2ImTAVgLXXLVOvh/Bc+oKEcXhHYmhMqHLfwnXD2p/238kyKLswgOsd4/mo
vrHSvH8Wu4LPM0f0vl+AgPBBCMlhzxu0AE1QS5FWqxrIJrKJgi39MpaI+fqrKsp+
ygAm/bIzN8hv3BtiVf2Tisq0/50VSFwGyDXEQpG2Qk3/WemqDosUrjWX+R7n54pp
fB1AbtWe0Iu/dWCMtOWOOIN/hfGVs0AirxAiLCv/tFIbk9B/2f2LzfpdP7p+YwX3
hOYtwvKarj4Rp2vVGRXXzsY0sOwR1S+mRIaOxu/JVBvOG1gliEdN7K8F964QhuRU
XiDHVIYBXlPV0iLErXHSYv6Nm5ojyAYyqI7JdGmsOeZBGlWCGdwVeWV1TyBuhI1y
CAheOZGp5s9J1m+6CTlOof6+vXy56zKpC1XT8uSslaWROEAolofqV1yaFd5l9bW+
ExiW3pGCvCDnFvXxAAup2XqGjnBVOnd0qtIIFI5IpsOoKC6QyImAYcY7+n4gXhRX
iKpaGPHj6m/P83QWxK7gRYzYl7cEeF9Kd3u4SXO1vQDMeuaKc3RmleHCez5D7aiU
gBImZmbs9HpWirpREK6z9G5qlOYCU9S95zJ+bpFBtD0lE8XrEBuTipxLFUfleYVI
7r+n6MxlXIno89Noj3N9W0Ne15sbNoZZtLialkULpRW9o6Elz0OE2XHAc4wA652i
fTwCwce316nI0Sn1uli35vq56g8UGTMsfYdXO+Y9SpLhaFdCWmIIIj02vp0NSjA3
Q6GBqH9TWV/Xh4QM0Lk8x0Al3zZcnQP4p/nXWtRyUMku8u0fqcoR6h5DBayXpbr1
dduDREGlqZjwLc71OmDsEnXKlwKnHBtx2bOTyTm46YehJJJCcN3BXrczAynmmQsE
B+OJHftSKkhsksMYz9sgmvRoXFmaeWq0gWC4VXnygc6rSZvG+SRWZqSAAZAwVgLP
gLuzGi6bs9DdOYDkLNcQtPSt+j4EOXQ9MHEbcwna19gZTakzGVrmmAbR11p+tHnd
31OCyYvqSaoGrwvsGiHm9h17snzSxeZF92jQBw2DXOrhKLJBq+z5Ei3dQn7G8bAz
DzPbf7fjvN6fE4V7ZYVe86w7ogvVvyoYUWFR31/gPk/uBTX9IGGIgnXPB9f0TSpM
LPxwnwEOOkJ6wYQY3UqBLX2M8pZDObrFSiO0ZmdLgmw9adqK0o3W+te/P+Oxp0Sx
ceB5sbHF4TgCqnLFPisUZTTVYhoTjSJqF9qosgGOamYiHTBNjocklwezvGhAVaV8
J6w1i8/hITFzVXtcGuU2gm+7NWE2l97gliimFBZR5H5gYbXxbKRprFZPXAD7jH9V
GL+2jMKK1av+WvHGkrwfKS5ejKdkUtKNh8+nLp0zUF8e0c8xEq7l1xau9lHnCOmi
z+cZbws9MTKQEANdCxSyjGf0kcxq9dNeJJ5bI478gV8w2KllFLkyephpeRqcf7fL
It92rDrV3UvvmYDIOU0MjTzILa1VNwaQzb5sito0Vi8kDSkK9Hn7HvT7E2KWsW+9
kMmHpcZ+yrSaUbeVRCWI25LFO2ILJ5uj/jl+MbqR/Wr8giG6YVQNNm3/rgCxMjMa
aCHo+YvZiihsSfg8keaRPUopgkD4KrWHvp6/kqLb7x3Fc4UrHdpCsMXQQCoWKesF
cxG+QvtvMad2pxZBzJYrbLVJs5A8GGt7EXGvFHG2Z99lLchkJLsbNncbhEXZUOJb
ETpKnaqXYJKC7MFggjj9B57newvKp28UtmKooDNsj1Gu1IH10x83LPzIrms00TRG
u1ZeU8FZwXTul/8BK9V9EhL07BgR3yqrNO+V8/J4luJ/zPOr513zYp/7rDB8c6Id
yIwaSUAUdLUsHWmm9ZxVxE7UxVF643WYFh5HFkYevcv3G8H1Esc0rXhMlbtaa0oj
S2Ec9MJIAwOKjQglKifwDNksdwthjaXYGtHj/tbJfBsSxAH9AGFQRux14dytREpe
Dg5R3hsmKuYL3wBOTaDPYkmdxuOH0jIUR1UuhLAe5GChYtOPhRcl1cVSvf2QkTey
j3fABktdyhvBjhIMVsoEQbiLFLmEZkulBqs5g85d8K0NrySWoSsQMQVPUreMu6VV
saBKqEttW1uU+80ZLwUGtjhG8tjJj9W4tOjpG8tVA4x419K2yeNPWX9y2YPgHWhj
1wrC+Si0MlLp9gVwSLP4Ya/18W3nxPXe/1B5dRQ+DG8FY9QfdVCwH2pHEu5t7kMn
synu/wZ3A1jbvOoujGWB+XMbRhAOUWLK2Nyus32z4mO34poEFAZhbEgAyARcLkYq
3tqWTkAUIVf1IY5CraQdN5ahrSw9xx0Obtoguc55ZlaT42agRHcVrvWSr1LpfC8O
+0DbJHVErkKOKQCmYNFxKY5MZ3nNU1Wr9EAN6mYkvsV/EKNqU5dz3yGyFtPNpUI2
/PC6qTPN0NMBY++GLmlQ0DpqP6Oe0Xfu4RY1rt2vekSRu7e7so5MuRdL4H5e/Nqw
LcUGbpzy9r22RlJyJcVYWrm2pGSmENPXiqY+qoCcfiUNCz1w5I08rkfbNQaor0TL
tyZfh/QbXYBmLuaQas7SKK761fhxTOJxRSHO57R9i80Q3iiKLXQrYpzlZbXmsUyy
RbNIQTws4LA01CieD7lNeE8HL1YWa/G0a+ffY2XqHMseMLPno8+Tfbe9kIdywDJt
TZB4x+dCSZlQdjHzmLrdc8oXk/I6GQmp4gkCIXF5TniS9qoZeVC7ETol35v34uJb
GxuyT5OuUjJGnNXEQhkjbtZFoeOfIVkK3RFGuw0m8xFlnVx7DecMZGaEFqKcG52K
iFrwsg4PhvgtdPoYRlgC+/N+S4/ttYdzJRW8leP+m3iShJJQhfaCZZze17+jTKej
sdwfxj+EyDqCbT8IL800ufPgiVC14gFSCXBc5yeQHxtaj2zM90KX51GwQT+25DC9
WpvyyVSaxnslmEdVdxVCdaFgm8zsB/boyM9yzyVYsIVPjH+wXBRUtbnVvgFo9IYU
u3mdSt2UHHOq8wbaNz6uSz751q66vP9aA6eyh6aIRql+Bf0beKQxNJj+Gbz6zH8q
akV7GGrvuIdm9epf0JSQyycVtzZDXoOlp5z2s984Jeg+JJxFela9w/4v4vC9NX79
OJHchmmakIdCICgNiZgIIet/ErKKD8ylpD0n/ER+puEh7uGAz8N9jGsLMRFdb+Qy
Sge0Wu8WnXduk8F10xSk4klIsB/jZDbWtSCcDpPGJ4toS8BS1otVqoBUWhqwhiQM
sIwHHi//ssNk8wB5C2E2O9e2HKPSbGMTlWn6Hnc0aFCjgl+ikOJ6wqNjzCjD1Rks
qu9glsMcoFCIZroTKfwL49y9mo3BBIUa875X1Th/7tIewHZT/rXrVmfeRxYtWwlg
BCJw/hucsOt9to8rCJXENEkGjBCkLAFIzy64QfZK2Qwdv7X70/sEKCtm2O18B9b3
xoh2dFJJJxDz1JVnBtGPHZpAs4LWy1ivTbKBV9xA9lwgEUVovBQm3oKXaD9ykl7C
4sNcyn214KnuwfnmRz3QLW6OHAx6OFmfk21pw/VNJcbFGqf+dZi2lFZW3g+mGBJx
l7mzhdUii2Lr8BRv47TXhBnrcsGh6bqqWdm53hfT61h0BaH0pkXf2a9OuBgMjBBy
AwLY6EZqQc6Eg4DH9nfgsdvyKL7GTGthwSEv+Zm6zgi3O53frOWTbPczM+7XKZnq
JElBn4f4AjrFVf3bB5AyiqSkWyVbNM/b9pDSUfeDStLAXC4UKTYuz9CtvZMEuRyq
IWJtyXJ18HTuyW9WWM5dmIJxJjixdbkn12kqOoqyAci/GHnKI08WBYd99aifSRIF
BGToS2ZsnTPP7B/YPOnYd4gtZNQJzbCAAKgpuEvUZnv7wsz7VY8QWwyMGcF5DlyB
9L9kyWtQm9L2eVHG+LZksJ9YTLY2uCfQ+P1NQR6jEBj56/aT21yvlz7phZZyWqCt
Bo1Ko3Fo4cf7WMwmyRTen3UnEXNABc3hkahjj9uWf+G1M4PlqLZAWooipHYTdQ+H
tG6f0C1pOevCGnJzIPBa771aOefERKJQtlaf/75ZGsU7e05iAxzIQDIdymgegWBQ
7+QD9pieXTvnVrUkcBNihoKK9lnp5EYcqoczAtmI//7ICoOint9Ios+sNnJQlqv8
Qjxy9GZRpPJ4X92yOD1vAWA0cJpUIW8UkBlJ7i6JVVbOVmV6DgX8tFo415ZVxzKo
oUJH2TYdvQsIZfIldV7ff9oTh/bwxRgGIPbIROFD7eUCvYBZ7rwZpLERdoZ3DbjN
tzkpvdEb0B6CEXHkhjGNdP+OcuWl/sxLlg64qDmZPxxGYeGBCI0PJUnqicEIGgyi
2TKSW1FPKKxhCwaRxrgXRwEAAKo4asyRKeeIuKMqiJe8fkQe3FUsusd4P6NBAnAz
9LKjJFBgWst9j/4yLiIfAZWrwVPzFDhr4/gMJbHW1DLv6SZwZnbCcaXR+lxMTfxI
3tckHRJkXHe6sd1zSEE1uOQBQosnc4JeCzJ1QvJDkKG0LGK0jDXwIyx/ZAQ/ceGt
YC3lavWGqI0rATkoHlhFY5rh5p7Yj4tmUmJQzu/hyNosz174XHyyh9gOZq7oP3Gw
2zKysPQQ60xBoCB7P3zCFymmlB9t39vFX64f/ydzC7Ili7+pw427Me67SH3zBUpN
alNlvL3NmbOWMR9d5Wq2rCvjojvxv8HSGYB9HhEio1KgibSsjVUDfkayTd81RL5+
irm04H6fGvTc2iXXncb41R7kenKhuhTvaIsg5Km/LVg15RlUksuCKNAl7PKwF6Sb
XwVenmxEtMAQM7q23eHnWxzj0hIarMsq4ifIgSKWalQ7axYr3I08s1bwnaQs0TsI
jd2mLPWkY1aj9Rp0sx9H8qfizqxxWXzf2Ahk8VUOPv9pNCjnqZgAMxGda+2mk3Le
w94xngeowlPhJehk6e6rYLhKy5acFN8uwgkMvhIxNDYPf735THa0zB6omtr0A7GF
H0cZ+bkyYhu+aLd8IePWQL2FO3gDv+8ygCjTuYTJrmOX/xayHCoWXgSO3xAU4nd3
S3dNAx3pQAJPQLvTW86qJbpaqmf1KUGoaYzuGauZLaN71j6yoitxPVEc6g8FwEn2
td0GrogU578Lrp2shHdPFwfv536urTkoXIKKo3PCApyNJMeEcXf9l21kWbjP98cl
heDOvgegIKipQ+zqvbBYzZYdKbYBQGyFKlfEviYTzsSDOWb1nXGkQqGSKQu04UKv
ZO2/3LXa7PlwkZMUd53NSLGLZ1JB2BsMJw3ipJ7qt3+MMmyHfcVqsVqxitrGgT+T
y0WQJ6T9qJoNgpR5vYOOkGX4Q+lxvt+mGo7bAw5SeAyjlyjuSWHSJbkf7SzWQuDa
y59KgJPdko+0DV3ULNkChkIlBmafNOYiMST6p6UybShapSDv8tpzjWTTSMrkjFLA
wZf3bVKY8BpLBameAElU4vFIG4qwhV9AcgV+9R42hceAxeIhHZtCY6l4op7iqyqH
X5Lwq4G3eOHCLCjuDdGrBxjiTllf4ecT05d7qdGND3b3J8iBskUGcE8bTWceUgOJ
IgKGmkMxhgOpZ4VenLXv4oNhFrRapNZeqZAP4vy9zVfyuYpS1S6tP/O23n3P2+Hw
gBAWpXKEJYj/GQu6JR54yCNAAoH9Ez2eBXrRx2//kA6madAWPY7MokOTnsCWF9Ss
VRGQ64YxQDUfTyRKPwBfPZDgslj6kCywinTjuTOK27F9aGCAwWuesga/V/roZ7//
phrJpD092At1fDsT51rx54gxuR44TZeiWRCrN/xIVCbJ6rhB/Iy0+kNnlydIitAr
xj9jEMWUFU3XkaePL/FGXoBdEMicEtIFj7w3D4zJwRJKWtrPq4VOrExPVWHCdepA
7CpZhpr1jMnfZUDwWELogBrKhbK+VyeJG9Y0toAExPF0tlA7wy8PEh7YturclcpT
Vm0+e9U5pIVhr948pvARWo7iN7zO/WaDCfeqsHWI8lRCMvDjPPpBUIpHHL/3qSkr
URIgQ/51j1/Wbj5ym3trK6FKskLpUJbJnt3y8Sbt/0ZmOqerkj+In7Mzo6Litj7v
rKDjXnTALjHuhmSlHtTTjvHSR1mSQV/3bORpSyWAGxzloiv3XQpqZmYUjc40T4MK
nXm0g09ZKviPMKBlj8p8gHjvMsEBaOez1HtRewZlAe7hpkZtWkHYGBfTC4YlngBA
L3VD2tvdHL8kF/R26xf2eYoPdiZ09bMMheMQEEJhPjryC0nVa78vKgvJCTMnFD3g
L/+3NyqrXGveCuRuALmSziDNlN+5AF7/7prZjcK/rR614biaykeRiTzBWvZmotM5
OKF4SJd2EsgrPKT9gA6Sef1AMHbetjP5SDwaoerupymYGYoawZfv88N9a9pcGf/v
ARt7qONJ5JVCrwPzDKVcipSGnVq7xxhJe9433qyUmnrgLfzFjVIAa0OkViWsdC5R
6BTzzA4plFjQQV/acbHwEH34oGtTO0YY0usYnxfkZA7pVYlT98CnIuKy3SHeb1WU
EcpNCvJCspvFdIduQXXsMOv1CBMWH7CzUb1B3QkVT7GcuM7PJzJFAhDXCn63loJb
2YN0sOPAUj8KVPZHuE5wdQn6f7QhinvyQgf+Td8MtV/y1Oh7YUWhKnIYk3WnBM6A
A4dKPnYd+WAKRuNMHrUnm3eMq5pEjsYhzeuVcfTrKforGCtuQExaljMvug/onvI5
4MEfIlQ52P3C7R4LE/nxbbR7nbmo1CNLS337nbb7/YKfctc/rvktb1o4i2xb3BaX
q7odSVhnNtNO7KKSsoXwiwzcxTvkJzlV3o+QGalpTDUiwM0q7s3phVN9GAi7Bs8r
iu6N9YoSEnZ8MNgfeR+52lwxYVa/g6NpmAfs5AZn/sO4AnaB7p6clGO15zyHbhPf
y3JLSC4qDKSJsrxqmOLN6VHSXrx5hCr/HvMwuSkec38nQ8uNKYDYpjKo/htE9HRO
t0Fo3HhfL3ryYEylqjkkG5s5ArHTBxMBlyZMmTVhNlVLevdqxPxKsFPttXkVCKjS
pqqSRdrCKK1G76JjhBFt4s0ZuKEO8zgpsoJByD0BHxBWvcqtrdFO7mQEXTf6xyW5
rVEj+J41aObMtrjj6zkR1h4irOddUlcqUP/eAyk3v2AT8AeZW8SBfqevFu9nqHhU
5ELrepy5d6ptbHUZAadrwNm/4Sx5ZCZ5dsw1VHPbCZdN2AEYCWuFBCA92UV/G+5s
IL7BQOfpUgFgxFUZ9UnzVt5fdt9KKy+Iz+tffqpyWjZ3S7Jrqg2H0toyW0Lc/jti
jun2H9Dur2EpMZxFgrQpHK5ssOMtMRrnyhwfbGlJHCetATwMB91lP/LnfQrnPu/s
UuznL69OTu/MxpXVmlQb9yA+redKgQITD50fSdLsKKDMxYbOxiDyZLdjn63BtHwq
ZToZUeMAgpyO/vOZrTTJJfp2pbhGYMETP6uLwabiK40zd/dJfoEDuAf3GvqUpwNW
tUzE0ngn9bGAiReAjiqeA0WBuK40rBx+j0K3h1PlH7vTvf6kxC292l9t9zKoRhcj
GEI4r8CFzkW3+LcMj5ACowa/zkc0R265VK4Bo2CYFYwQ71ItZENImU/TDYobefXk
JTCsjAROKv/zkR4iIq5ERTqfKOtFw1bgiS1b9uEKUyTBTeMMq6pEoqeTbYQDvuZh
Uix3yL91nfyOaFIHUgs1wqyrPkeyxp2na/1jgCKSlT1JXo6tJy+rF3Xl7fHlc9ut
+uvS+Wk3gUQQkLn+sR4rl1DapN9/CZSVxNtqS5RjA2JqNVcYtU4NrvmZ+/sDJONk
Ptj2/eozbEgx/YHkWneOUaes9GsiJEZqQ5hCKSoa6fYoAoMC0dSxfLCfIAlTJQHq
6E5p6qrJhFRwtTikBBI4ENKeKnRhCD7jYoKNXE1vSj/hA0MptYSkvXylFFvNsvdJ
kIC2DL0Ot5/lk1FRk+poMXbhNkoF+TAPa/qNyWKxRHEHwch/FMTgazXbr2RYx+Dn
/jU3gnwZA5eHhd91yGKAO43xRsHcID3ceX0O8l4i2KBFabgHPJvANDGvowD8KD1m
UTxsAlDxRc4/Gzo5ZzSsjq8Gm1UlqgYHRdPOO/IYXg0ymsO56TH8d+q3TX+R6r8U
9vbrQ+hvep1QbpHstA377YjOMKLppQHGJOiLae5sefBqVqspFdl8a5wC96ro5HIT
Y18vIhs/on3phEXhueX5hzPhltunYT1OE87edsHTtkQA5dHBHrq9VEli7KyI01/b
Y9TWcPEemK1quADwsnkoIBxDh4f1KL+7q36zZngWc3l6oInAA/8aLFi+LFqJMgZ1
ebyJoT54ybqzYGfn7rqFKzkC+ZzcPeFYtlMzMsWqei7cje3H4IFg64pOprfKjyDh
UPyF+LIjsjGR8TVpnVp6kUv78tmQrDMSUMCiY1n+B9A660WSlWJgR8/OdwhbuWhs
Mzv/PcRuQ5RM6jk4rZHUdLhK0fXytULSc+qrHAK9IduPVI73KhIfYVP7yrYQmRGW
NTrpPJTOzy9T7pkrCaiKRoKnC3cLlyxvcKTDB+tPhxrIJKGO7x+UkVB0rnk95tMs
N5IQJCBahmYiWjPuxX/uQY2LjCy30eEFLQu1MKNM2xbjjDpQAJQtSNqrYNzdpPfD
P1NWkXltgxP5MFa/axZtkZQDonbqH/JEV5iLZvZZcsEdoOmf+7ADmtxa0taQyezk
6k43VG3XVc4/LDPoDpU1Zg+tJNPotVKxJwtBGmQpOEw/vS58cQfLOdLju3qGEYY7
W+kPNp77fCimVHuTsghKp/RVPzTMvCFPbBSfUupVF0tok+jYcf5K5wqd/bYQWBlv
PMFeIswA/wo830vSlNWDqP8SwZ2Lg4BvYY+VNqQ/rN2HQaKkxmlcB5fBM/Tv8MO0
qR/MrMnMn8UaH9QeBrJqRn6I4ahE5dRbxq79LU03Jof1tKI3b557AG0Ayht887Rt
OfkvoZE3B0nSSpNyMf5lxvKuQnHL3K3JyTdljRaCmBvDmAYxp1T1mSdTjsCM/JoI
+82Jlyn+OYjRXvMM+4mTMkjKD41CfcBJbg6NMh9FBkYnodRkYae8udrNtd7vUcVB
gt42Ap52CW1cgwakxAkFAxkGCuAux2XJY8KUfSD5A7gQXAn44t3oiWarEqJ7swSC
iTu4VP7TQHKbcBuhQ5a5eB3p0sh54UZTujrIZEDJnDgh5QzeWmudw69d2ggvPWLj
dTMKQ9OIb9jIvt6fv+cyWu2Ad7zoF/q+Q8uPKKkJ3Q/F8ZyUu2Q8JKkK2+dn7Dlx
5AjUAu8RPHmwZ15FNFPIY3zzqTKboVIeOoWrWC+Zlq0r3ZWUNqyWBMH3KKrzp0kJ
8n+/Nz+e42wEp6Tj9OzfHl93u1r7QPIdGnOEv4UysxvJMC5VK3SE0s2Qzj9iRaOl
HJ/vzKPBKJMeD6bFZWTBFVn6/RhT9271f5xIXedaZAUaAB82WBEwee32UUedFdYm
n7PgKGcrX9Q2c0PFeu+kDFhq4G/bnDQo7lUQuu2Sv4vTJ6qbMUw4fQnMWD5/77nb
0YWYzMe1gpmAAQSTUAzdyfg0+BKqi5aDnu/308BalPVLCeCq/PawMb/gwT3RthdX
pD1t1CNpT9C1LceLYmbMaKeEIfsHrDkrbfVIqrsfPrLkPLN/s93ZGAIzhPXYnXYn
s7I6fcooNbI9PLe1ecYwuOh3Lp1VX0nqaYH2YEW/qZRaWu2YrLPe7iEnH8m45xHE
jCWGm4ShBIEYasF1CpwxLXAvIKnlFjwGw6gtOIhezKwHIMFJH2Gu8YL52ZQvGici
H3zd9s49Rl5HipZGftMWlcl+BieA85Q954uU33tG2XLhabuij3sIvbjRV85Y5nJo
g/Mlm4APtanhlBcZhT8WKgVOvdV6ZIV0q6HdX6I07fZkSm7+8NdBWhEbxVrKAD+M
txQYTTE0GF4dyc3r08lTeS8crqtdKuDR9i+cX9IluD5dEn6a5/t7qIVysM4B+u8/
W3fKSHWCfdgS2ONuzmKzGbXT1bTbFga3mpt9EyXoQqQSmJ+PpGSbFxZ4ByiX8CXm
6OySd24vOT6fIdLG0g5JZXRNsG9Rcmz3DUGItehuolhLcAlcv+LRcJyp37n1KUkc
BWFubYh/xM7sQHCM4jKQGgYXhw/0J13kqUfpWHebKxKrTaYktv9zrSJI/z6JAKhV
twGP+wVUCry/Ak2/Kd6cXE8aUuHH8wuHCt3vmGFjm9ckP/Wx2mUBP3h8+4j5B1t8
R8QzKtdFmC3BOFdkVW4pBOb2Db1r4pmyh1PSrptzttLW2/nbFgcQRLxGrMTgP/dB
weCtA7wObKnsVfKJIMY3ksBhllo/Dt1d06RopOYgphoUg4quG1mr5V6e1MLo7QH2
m6O+LTcRSOT4/GiLCs09UOogyyjCOFK9S6lBVamau7IK0D1SvOsiNmklJRv0CWN2
Noj30TcpNTYlAOJOc+0orkDQ52mmqvU5gB2ulkZL1GYKCJ3wm+R3t0uazT0md3fJ
XaZBDdvCrVEmuPY2N0U4K3cQqdTlyLPRP4KG/doui22ANsMUWqxzsEYjfdwB0GF6
8267OwGkk4wz2wxwfbHreSPYaApL10iWLFr+1NXf48ujDykNYKJcYe/R7FIjXC/3
70vvIjCwxFaZc642gHz0GpoDjijepGJ4ok3MaI0V7cCK3Xq7DYjc8o9emiBAdC+J
xZYtJtwTR0inEns1NtVyczBAvGDxYEuGvDmGeN2wej6NAp/GiuU8qlbHs/EarlCc
jVwDI8WRe/wlEZPGPRXMT3NQ0v58oh7g/wIbk5Om1da1wORp+rC5kWhuZnVhOfsW
0mMHVKxwfOxeXZnfh5N3U8OqflmoieLUbvP7vD8HoD6SfUlXmEXThCHwWRqNowwC
zvoc/RqSYOjoUU9xKPBY3dEy9rJT9qMzu+RBEbMaXlh1Khys/JpnjnM3UKEGL0IX
INseJnEaGCRMkQ7HTHuKOoTwwiKPJVIk7z541ZAA2KsLxViOgS/6dASIAmHGe6zo
/1vxVfFUZ0Dfa5luYyYQtJ6H4lSAFmvOJPRpvwmmCQKtF9CqP6kZ7qBuPzWsuKPE
6rNs91Ef/FF79U1iqnqcZ/7pA+q19f4vew8wnPogdWZX29HbGFg03cOfiz6iexZV
tXQpcOue1O8SqOFdr5jz1JMgoMQs4F1JN70jzifLWSLk7T1tDVorlE+ussVI2meR
ZI9eYqDwq7lT4TvOrrou3Rolu3tB8M16OombvL89kOZ0afZVN4J7m1zTe2G/lzmq
irnZTcQeYv3x7bOs+G4kcDfd5hckqRdkKy0Q2Iu730VHFq5uOZaaFXr05Wzx3mqN
TjSd7SNwKM15rHechSJufljm0puPeJ9uY8JTPPpKvR8nOks+ghKbuLeFKOqjARC1
zS2mle1PGcUuzlujDJbehgX52nnXANQOGkwg2eHI43TGDMXt/N2Qxvsd+gL2f+v+
oPt8Guvi+GIDxNLdjWL92z1mNPxoAneZ5wKbmnAuD6n2bHP2pfQCb8n/hTKS+O9q
2DM5gLPbEz2uD/xeCpIWAc7a8iI9mlvpmF/INtp0ITRYHEUxDLS0oL2EcHEN5RC3
EPX+UDBl2cIB2qGkOCDEyjxJIa0kE9HYuDU37dtsfy+FS8ehp3fkaZ2N2JAvIewG
NslxyqUW3SU+pLMpRROUfbOk7E5rnprzQPchVx2zGkgUxdRGAthe+VGZEDRiCe8u
y6faXj3UMPqT6fYmti9ClPW7445/P82X78mkNfEr7ZfqfLkiHU5mcscov33vU5Lg
mLqMTAF2ZtEy2a4NrIf4YqF35fqlUWgBqgZB7rNb812VriHwcZFNNJeXKNd/+O0k
tGnk6G8dUOxHABQUmFS4l05lSfitSqY/pnZgxTETD+iASeK+WZqRZvQlnTeZ3rLC
+KRjROMpYG1GdM3ugHwRtKIh6nZymQnYqUNo4udG9A6A9RbkvIGRFP+WSIRFSmkX
owTP6yxnKDJhjdTx5on9Lrb8ulMo2H3ggYK74pCgMhnkNNQBjPbJpUD047axtNuU
kgwkPN5heYYnTCgE0FGCAIt+bzUtI3D9oOXlBXvQ88owsJ91NryzzLo5LGEqWGkg
8SF0y4eWit4m0AUgcZTs7Z0JtPLg1nXLncz0KvxvZL4uVg1sqJw7WWRCkq6jGGAg
FKjoQQdjR3W2hQ5GhOUVfQRsuHuAFOsJthG/k0WC7GYT3K4Pg1Q1YTkL6Z9XWq54
cYrPTit9Ku3WHQNyI+WQEDxWzNJyQKRJx7UFUFcXVycOwZB/zIFTK7INT7dlB3hl
wKcDXSdhZlXKbQOu/sAgxR81iC9S/UbYWuvNcJuSzCOrTYGrzDslJVcUFVI1rBKq
0n1PEmJHOsC1Lwmd/bYdqWOD/YpeXPDK93AKX5XpUqcb1i8KiAZvj4it890YYOf6
507Fli9kVOJgQRkd9osZmxe3obNl+hwIgyxB3rY2NJdUcLudSLkkRrCeM0qn1gnY
wu61CBOr2iavXQwC70whvAyyTL3nyKgL1/0+4IPfLzHBoVBFEyVQkO6/yTdtFoAV
qjgVESWR348v8DpIT7JXVjZtUohY+qxMkKmHLJI789cqJSBrvVQ29PqYJWS/6gjD
DluifLeEmF/yilcmwEBhFW9p/zPcM3nYsW5pNH+170bbSMku0TBBf6QpbPofb93I
mHXbtNfcF6zg6B6eA/A1hHoSx7Dr5rGL1gXcRwhoOI07FdlENL14cpubu3ICvZNq
o9OLxaSqBOBRaMigeYpid18gCCzPojVjdFD6KSj/DVFIwO01W0YW4hqkr06qMSLl
kAK68mlOZXO4VSdwcXSQSudiedl6WQvsaKiZdW8iarQ03i5ImJBAi2JdBE4dAgnV
or+pLcHqRlNeKmZdV0cofrtU9fj41ILHPrzrq5QzEAbRyUMb3WfOAJEXsb8dRdCo
Tsa5g5dazW0oY1U3dIMD3o0jHAtrcq/nk9Te5SsypiRdZJgGWasOttHK3q1CaCcc
OCFKVUgBeMkNQJHODCf6v0osD22wFaLcnt+nNAONvquX/nGDEwMVkvE0dxKgeal/
bWJOgZ7HxMTwL+uvjDmTv1JSwZgtnoq3x4gmOcfxDbSPBOB3wvr3+phSdDC3gcfV
p2iiRMuh0LwyrzbwlCzz9+3m4rTqD5zfi8mbGrtwMUpGD3JfE4b0TyMuIbnYZ6EV
lb/ekX0nt0yWdG2K2eiQT+XsAZyo5Cn73dUsdT/JTFlFlmcAwaSwmDQf0rTZ2efF
jbyooukeaPpUQ9Mk2qvtGNB9FUN0aDS5FedBGM1dwd6zkRkSRpxQOGmHMraUquGw
GZEmTdWF4A0rbdRpyCzx+AW9sFi7UHVqTRIbOAotcDnWyXG7MhleTQqEiKZIMe8x
3dUkDvXPtBywCKhup5PA8mgfzy2omP5nwvG4xDYtCWdunZvZM2kI3R3rsix1Ylxm
dNXQlbjPv8aFoWqVQpBPmPN7b24ts6cLwcliWmDt3+qZyDZfkKqkkjdDa8g/Sgvu
7nmLLtLueSwQDO++fiDOqwAcZKPzksQIfzXi25V4xn36SwklNtKsvWD8IxrfXIw3
+mgyFSNmsZYQ6EnPeH+1dyCVSWAIRqEDYraAZO5JBBxFPhy8fLXJ5m/Jtkz0lFjq
eFIjxbliURI9+JzzfvZxKR1z5jKIkjPSO6wW390dhi1qWgOrBZoV9VdQTreM9Luq
D9BMUzRldYfRCFwLrzYD6EjsPXkIobL4U/RV0ZJrpBEDe4t7XiTMo+fivteUyxT3
h9SC/D5LtkFVwa8wG0R/YgyEvSkNyANlqVtGn8f6aifPcmQBUPhy6im7iaHrQ8PK
bjuPWtN2vlDVPilFwEcSafMBnMsAF6T9OTHFfOGF3W87V9IebNhGb1WEN7OQSqtX
RrixhjyVdz19ROSU0NXWlCGwAc5jd35JiG5UMbYHqfRosPcUbiwW/O9Zr4eRRDox
3c8z8hHXmSf2Ps4DHFmrKsRKo3+1OV7fDh5uTeYm/vzwVrfy5zl3gCbcRwW2Yee0
auK8biJWpblCXM+7WDFyKBsMHjbZLEzWkR+1wiX5HT5rWMyKfnNxaRfVjhBPZ3+H
j069NPR0o9AXHq+fuMapQHKT3mCc73PqKZQt2SOnMW9hEmnWZI6PwvJ3psei1Icl
3RdFzc2dz3uFyWt8dJxbmXtGyQ4ekgII7suanxEXnBRaRu4MoqTluUAxABGzxcYV
szopPyJkzpbiFaJXk4y+awkQnBOeJbDM49L8vtphFMe1TnwboeGST1xo/61d6ZJs
jn17UK1dmrXrHBxmK7jsRA2heD3SUuxq8IROg9NKnkjlh1JxhCMXjidb/IbwUGmd
p9e4Jk9w67y2AfA31/zgU//dngoZdnRR6RIvb8zBAe/4e4/e5TgIfElZjMvAlX5T
bQ963HJusH6COZpAyk4wMGpzRTwU3+QhsNHjzKX9WvV3MSFEYAGyE29S+Ow2SmJ1
RsqhfUwdXx8+sUsUZ4oFBjphLuOhSE03fGX2rk52d8sqKNMgnutVXGjXjA16vE3S
QVrsajkNaM9xPS+ehvrpikksQ6fT5hggPWXJiojlAIUqaHwWgqBFMGKnz1NRH8F4
owCw2wQo52teL90hxYPdX+eIzx2x/XK7M/xp3oH+bevGqHwcbnoPdpdTHlOJHyYN
bkZzWELfs8y6t58yYMnK6Bc4qsEIYKs4zcfd8h9QPNNd1/WDfuXXDFqcyACp1RPJ
FPH+NFV4lDasit+N2DCQt1qiYujLCSGZS12Jwljssf3RnhFDx0K8tN6q0bRqZK4E
JNmb5G9zEFXd1EFmUEN0JLo7nnWUh75Pah8VLnhJ5PuqHauuone1a2UhrfO2vC14
pu+RqLzG/s/RVmrNy2gfKJUydkcQWKDWiu4+ArsoHYmU6OL5zMsm7niXQcZR5dfa
eR9OYFTEyZ+j2vb+er91F5PcHLRh8HFP+1aj1fi2PIM25iTgNCEHtc3LNw9s0KF/
5SmZV4ku1ikjmxR4JkZUEjixG0UVO9njcopfl7mpXiT19IFQEqnxlcp25z0Rwo4a
y1IaWIv6N3A5+E7UBqzGNeoG7iqWB5+y8Tmnzee4ToOfK9OfbLT345gh4kezlJKF
oQpUh+s9+Up1IZGMm6ACYBVMq8H/WLkfQXhQj96eMzcUMLCEHy6Quk8rn2Q7SfJe
Ww75aFhva9XlqtEiVCS7XDx/iCOsig72RMiQssGX8miH6RuDwFVhNv5j+Ljl/6Xs
q3s+ucITNUykvDth6gnOFt/m/pDnQj+80bxy1IfN95g5AA0mvGHAogSBKx3wbBPf
06xezhkFAU/Fh4OsvbmwbwO2nGPsFvZh0ScFcuitWLoU2NzjqJV/lQ84bNPweclx
bmrgjABE0Nhs73oJdmXBnj3fjpJY7ELhP9BLOY1iQIhtRbNCF+RJKW1zEjIVVG/m
YNWWojRAhw7fqaRLsZDq9qQ5xKeMaF+lLKmDNZD3V1+1Fhf6fMqW/Xk86jw0Cv5w
sWvJhFUISCMt59jXh6AVsXdeLgWzp+pn/ZDmXMBExYLr3wuzvYuk47i/bpuBspGV
FtFau0dFSfimG33S6bauV1sDoPtDdUPK6GSX9S0MUW2aUP+ff0iz2xSPnRc084Sl
2hXIhl9jsK+DeWT3VgAo/wDl0f7Nrkh7M0zIQPoC7QnMLv3/ahFrDsGtADGxbtFC
gpVVM0ki4EN2EnTvGDdBfH0xnWozu19IfAjQzY5PmdMg+jQgGh8SeqNWG0phOAbH
xdTJwcU4Y70QZx3lJ98r7UwiUCvFlnss0IWBiMl0rQMwxgIcjkkQft1Z8N3l3sI4
5QVCWIrRyrsbvlfq5vKf35u2/6995OG0yr9tFrnjgSx1IUTUNmRLqFb79/ynovXK
kZTgKrHGYLMzHSEi3FJane15X7p56l3oBEIdi2EnSuX/KphsPSJ9GlZA8KeVQ2Zr
K14HF6Rd4LDgGOykmnDAm4N3beG+6uqbgPPi1Kv/+Jw31FFghtcROQmDaxKmOzcY
hlNWML34IxL2emMOuGAcycrfnV7eppGxoC4q2KpYAGn0aYzFxy8M0NHiOHj5r9D0
0mKFd+xIimSsUIbg7Sh68ew8KvVOB3yKE4GlsGgkMI7aAJNoVle/6hNYETUdGoEN
6cD3sles6TKobjWYcb1MEno1FOXI7wvLab/LzyhP8a//4flju0DoUETWH0uJDkeC
R5rAQbF0pZfPlK7RgLK+lJ4YEKMfzshag4aauvLivmoUIzeiZ84tOWvb7MyZLFgx
y3Th8zAjothooudwYAACp9Hgz2HC++l/zmDYRIQoIuv4GADcq5CWoHXomVi9tTrs
D5+beCeSHA7/QBJgZl/wfCcHZ/41m7l1RmFxz76s3EEIjHrY6SuWmcWEWJnfjfjr
dgMWZQob+sh4iHCxhg+Hm3x4KgGT406tIPvmD+aJtPkNKktcQYsOl4aOUS8UgMVM
NW+KwNuam6iSqRtAFyRilsje8jTOYdy8+1Ao+xTBDZGOE4Wu78ZFOEenbiaFuimu
vOIYi8bTQQE6QGLobt3Eawknn5uFHfodOPbH/ZaZj1ql8VE9tDk69HHCQ8M91JzI
V7MNTsGgXfNUqOFJ8fbjxiDOepYGJDmA20fERztYdwWj8UOaLJ6vkRPTkIlr4IRZ
svqytN5bxSjEuY06bs5+gqc9JdF6i0WtKuRjm5ZAjPTs5aH2OTZWqHgFjWedTysi
/KZmQG+uqNuvQWgnPcdwAiJ0Mli+CVu9xdYn8h96WW8VJfn/itXxr8kmxPlFrXwU
eO6Nr+Z0qNLLBLyeN0tteCmNOwojp8bEN5ej83tDkycZrcrpq1fszieAq38bl3Sb
PRJbKQ8668vtpBgGz8udkTGbV2c22Qdd34tsvkPrr2vtallKLoRsqzF87ttHzrcg
S/9+hBc7J5wBELN9WkEO9vBvhKFF2uVwB+HXI7v3up3Yp8/QkyuYvy8zedqbzkAo
dkUG6YUqhnE2E5/0UedzyH6phVW6/HAL5s7hqzFhgt9Oxe3+IhXk2WSouGbwqmaa
BGw9EhEbxoANlgo1TM+FW7qIvy7xB27IesqSi8ZSaHIRhUmk/0jSOcFdQkrmYTXh
eFxSCHwCganzR2j0LEBrE0iDmMgtrwEhFeRXaiLmcYcOEIaPHCeMCsO313SLRSS7
ZFLbDdAkrPnhpnDldMkRjg9ZPDPyX31DGvR35y8p7lgok9q81nxE95lu2YefXuE3
VCEx/vKLrUHdn8HhMzTbwfAIC4hXEJQdqZLBoE/Qx/BElaIXA63bseFV9W0OFAz1
DXq95daw1/9WT/Ld/aKB+jjNrSvHTSn5DF+NnhukLivYUSM6P1mvw1i6KIqKTEVO
usyr7ZudQPonYJ4ybtI13470ODkJuG+aiRUvI4K2PsogFNk0HKTSLezlgHs4Tq5Y
N/7nCNcA9FFSOHc+6Usuj9lEZlQjTV7lnVBNDehgvM4v2girz3ApTzDVFs9WVM9Q
MtEWIzlFAWBNB7NG1Id1SRS5tvi/VAripX+qctyKBmklfkRzEdbQFKVppa+y3If2
rDzDohODPc2rkau8sXmvj+gHYdcCivvjg3MqWaGYJP1tCPgvY2s2VnWv7H3jxhiI
rLHo2G+I23hAo9/I1APLAOFYYNK8jRm7D12oPei4ekApFY4dlyzyWhCKojVAj/Fz
6JsYLkVuJIS+20DgCIIYWsEulPFaadOIyFUHyweEQ8CVP5N4/gru74dOw6XKkKSg
4g8itDUpTaVPNh4Mloli1fUpsw/C0J4fR7BuxmAK97BuMlQpSjG4cPKbeKj8FL/Z
2rWa73rSniQPRA8O7pjlfPKON+uKRHBrPT97/A4cDk2M+YAHiYPOtJEVYCoAVUJL
jIP8izVerVlKcdLgN3fF12UUOl5wiCnxZ7g7vGFXVqKhp7JBAknIX+bNNxHmQxYZ
WzwYrIAXyfYtRQD3yhzmHwjB/zDT8s1LKqITWRU364wzhvDNJ9xODcDp+eFWPNIn
ikSYBw9cF5SNww/tUYnI2G4xKyCQupEE622ImwnjWRAkfmouOmYPpoY1KBMGyVxT
yIV6j62XKGxshWFWpoKOtdBaaTiho/N5Ev5j3KLudL7ieH14zIXvA0aJ42AKIO7Z
oa1OdpzlEoa3iFqOxrly349PFPRoV81Hpd0riM7jOSvJ2Q5xe74A2s5aT0dVgJw8
x48wZs4EseR5ify8fo2J61/rNcIuC9/l9+xEaDUvjL13NXmY10GnS0k7CFd0Et/L
G0jHLsjkBD5wuC7rdi+iCG26RMR06feFOi274J9NPoMEaNrqlpsHpXIUIrv1zT+i
e+rydC+UNHVB2sL6O38mjnBR0TVLL66hh9wULD589wN6WM0VxLZc3wJu9ECwg6Vb
elL3rZL21iM+EOAymgiZwkp8E19oJmJu3mRqOe9DToN80SY4o487gFHABPTLpnTI
K6oejK7Z6OUIuGVJaldF1LnUjpGqk5wewty2qrOiVWCnJqItbZ/xMXlxiaWGb8UO
5p8+jHmzSEgA2U6ZqSU9khgRLhAQDH4HXwOdw3qfrjhd8uvzmPZIgU9wLBd84f/o
1I7CY/YfbF/r94Kv3YrAO2IL4Xx+ZcMTy4VCnxw10m5AbtP+n+8FF3IhL45oxcxd
LkadNx4++VF9qlQ5noTy2X0lNWykDq/cjj9BRmfd4ZKxFreuB/D9bDDYkhsrpWD2
ksWqPik530tYe7zuSZCBoEfYUoX1XS0frmI1hRTrtDJfsLE63IoT4o2guWquPm0p
GfCCRGbwIERtkmBmvoPinD+qrNujgfWecpEquirHct9xGtIhLlEZZFNqlGDNXN/Z
SwxN0xMQsdtgkI0swUl+Q/JAzT5lsTt2u1blYJlD1yGRchmZaikArQDgQQe4AUNN
NCnqa3cJkurq47eHqV4R4Iwhg8liKGpPUR0zrY6vV3a4ZQoAI4xivBMVfqgfpf9h
hy+m9rMk/c7U9NKRlqHAsYAIKFlIB2254zs38WrrfLz6+aJ3KbKxK+JetpNg1Oyc
Fqtoyjc6RVWPOFHDqYWYi8NN07r5p84ok2xVBanD2M3yotz2Mv+dE3IYBmBhiXUa
xCieABBFORCZ2haCKZKtV++5bqfN1f35fKxTOPNyblH4al4faMHsK827lwk0yaDe
aPqjq0x6y/iTE2+xNoDLu0LzrZYlKuIfmxZ6PKJvZzEy6sXfC9SuvOanJUIFcuQT
8+atWZiun4VBGhCBX+NNJ335BiRnxYgzmtm8D6MwyM1LWBH/8cFHo03jIgZbY6U7
5yxUV2xTvXCgLt0S0X5Ib8mCIo0zIBjl0dqDqHdwFiyZKoa/s11V/wBBYBHGx/D6
Tilb2fFuCtLBn1CLf3S5fBBYvJjjydLwyIAuny4CwrdD1klcnpTaOKTEv7wHYHul
NQB4+GVfF+43HeRLn1L929jkYsC3SvXdNFiJEkNFbIaUBiC+Ia+7l5kYa0M/THhW
ZMzkJSGpv2RLbVfPexxPc5s80SGxV+eKx53Cr53ZW6Ffs0I72qoaHy7NpLL7E9o0
OIMXXUXg+xlDWUF6x4lBsDOJ6tiNFcZ0ScrtHBLWbdus1SsnW+Ib+LIL5BMCLmbj
e5L+4TSKc4CRRZ1X+eO7EcMxl0BSQmgSMcVWbhKC/6tyw4lfPBv0bDKUTPPCy04u
wK8rbKg6eW7D+FYLqnkNqiFO/0xnryCtFM8M/yRaonHf8DH2heY4c7wPx1qqHtoa
uvu0PlfTrGuAJwgVK7Qdg5yq69RpsTC63qAECU53i9XlJEK+tTq9Ooiog3bEJ3Fh
NLx2KMAsc++ZrkRbkLS5CV1pniruedkysq9dm8MYbWKs1KFpe3TBCWCpJx2zX3fL
Fi/EG4abhmfyegnwjA2Hf7Fv4lh2SOv643JLlhKo7hIlHZnuLpvJHGBK04BrKTjF
z0vhytPqe54TnkGMt/9q6XuFEq9lu1sYWFPBmJeBKJImOCEMKke4jVxkWFy9mWjK
dmA3L95omPW/VIvEJ3gGsebxGwjMeSwsbQB17HjziOr0HZgizzopN37M07VhBGYn
oRAwv6gIXhfEID6lVOI1D4KIrrKVYQUkKqHOcDtscEmT8SKwQpmR5GLzeoQ2zhb2
+7bWBSzUW4kTa5y6Q7ZFJD8ovjZCUaAKYGbnMqPKLVaCA2jpAcoKF5Nkzk0xS6Bx
z18KOlZfSXUmZ8Un4RmPAJL8r+v5LwSuJCGTitDdEbzRj9Yx3zHVL0Ejt16j2Zb0
hy67Pg7rXWtS3ZQyAj5a4SmEqQ2dzMnNxhv97ErIuQtGXkhchTAMn7Q9Iodqo1pr
/27ch4F6/1tkTG7Y8NddAX6BLUHVNmsSmUSJuGtiTMAaej/vQiU55v7VjT7BkpIA
25WOCptrXLB8vlJJ9p9BglaHz8e7XCau/w9wwZeCbStz3C44dL8RHU0kOQwNG8Cu
L5S4w4XguENis7zv4UhyfgZ7GnGPtOP5qsU1A2Ys4tliz/Uw5ii5iQnSZyp8D3Vf
gCxmk5xbRzb9kgQEb8DeCEpUwDJy8SAxJPQ4Tye+z7Iji4q0wyfVjMs7q+xLMdU/
xxuHSFLhpCl177VTb7cfvhlCp3G9pqfOtbvAJqn36yN0fZMN5rhQY6RjqleW0fjk
UWSN2kZvjlDd8k+OwD/gQIo4iELO+XhhaEMqyMa7n28H/bNoNfcK6RCIKQRJWccd
2EB29LeMbZzh7OgR+j3kMUvDjGDFdIox/x68ZY2S8yvdXsqZoNdlvtHs4wUM4hok
ZZd6vizDi2x1nlPS9W0xCiyijlj6/W0FOOccKsrq4FD3sf9mfK0BeQjfzkT4/WlE
0rmkCnoN36eNnFFWQRQE4oK9EdtaWndzrMXCAKSFzPr+1dO2WtS0SkuNscewsC2S
ol0oxJC3fTG04ec+eCUnwP1NIS1ntegISgKgx1QF1p5d0ODEOOeoZ8xokoUBoroE
3eqesd82VgRRIs79lmdpIKIDokEBS55hy91ejuRzu29/yjL1kEk+gYD0I1mSZhvG
MWP5yNG4k7CLBhcAmmeI4lWSIBZCpwMFoHaXp7IMWOjZGHOH3k4H6VqK+zueVS9c
lpq2aoVyJ0O1iLMLixhAExGpQr68xcYJHCZqrf+WmxKu1GFn15WyWG7VihQcHCFC
fdMbZ4Y1sPLMvxv9J5haN9CAjAmg3RuslveJbka6+1uDLLNNEdK5BSgmz5vzW8lv
Y4pQd05zlEizY03i3HDxZbBF5fZOc5/ISp+0j5I7nuFkXwI3RQNbyJy/NQ1iOQyM
efLcxVzVyzAo6OB9qPq35MJuYyeGoh1EXubofKKEA3qnZZTbHzpFexfx+1yUGoL1
hBHzu6O9KGw0b4tX27W3fO52nmeWoGZr4o0+nOb/9Vz3CEbI3t+IqqY9Gdm94SyG
ntmUg0gK4fRO/7EMHpAxwjMsYB0zY6kC85Y9FFXFhU8tJEkmjGPwN91n95JVQCHF
6wrT+ddOMrjtMNbP+v9jD2FBq7UwLkJv9a33hKrahL+fSYGehJlxWgNvA44D/iXR
nqcMq63polIDBNFm+YJEv0y3pXQbA9YSlNMDp4cVBrrbkpC8X5PoJc5RxvONjd/q
QiWvizJigDqBekzcOz8IgR4EmYJgIZSzoxzRA9fYslF0klZbsYyTS9UXlcQs/p79
iRkysR/VTOW5aIqq3VQAFfVkqFTXcOtgCzY21tUhDbrocuzlnBnH25gy9c945YHN
G3ODg9M6UbMdSlwRbKne3sR5z0HEpwokUZ2xKehmZEdwTZK7tA9YQFQrGb5DK6Wj
Q/zw/BweHbMztXbnSuKM2a6fnuZXtK4I+90eGsVTXROGTpec9D+QYsmjEBd9Aq8m
vkiib2pN/vMal+7mZbMQlZ56YFoDJSJBPAb3MkDbTJzm2rWaR2TSjym1ZoAC1CBx
Ml4DmGmsrGiriu2VyfCzPEQmjlR6Sp5j6157jZ8dWgzaH9+DT3uMD1/xMBuL8miI
SzMw9nI+e5nwEytMlMlEqsePAP2U0fZVuauPxHF+1zXGdniRC2gcbn+FOOIDF3vr
RYyjgrUdoy8z7uF6CZ/uSqksJ4se0hfRLWhixYFekPrHUVdn9nscqWp97wJahba2
mnt/10zY2dQXAh/ns5PHD7p2Ujf9ZaQAPh78oTmZa9ZJognpW971pmf8Vbab2y5Z
yntyoSrC0R335GDb7TWDk/hZAo9l/ziAcdxgbkV76QWQOD4B6CNc7lc4QxH2PkA7
04rG51Syoq0VTYHhY9H3IpphlIfC5lkoAl90OzJ2fFwS5VilPYiJIJeXqLciVqKr
etrQ1Hl/8l8o4SYGWi6FUTjBEsg9H+wBxOcUN2p7xKvi8NxsV7BVUA3DaKz+rkx4
OsrYz2zZToNswK+unbMz0q3/62/ct9N/JgyD8oIK2NQR1pM+iPZjB5GW8IYWTFlC
nb5A01/eSz/DKXdD7V6dunwW2mGfXJAXyBsntEqDMUGXEeDRoBb1MkhTapTDXdSG
Gmg4Z0OK1CmWbJGVdfKmwhN++jUPEoVpd+8ZyHouH1nDti5phBbNeQ7R48U1BgVL
fLeOOgSWLPY/PVqIdaxwSjW1Nr4EE1CPp2q/dMUjmfQVX+c430JkVjJt+77epUme
rImQpuOgDHq8z5efUm/I9L8Nq+0PMuQBEGVaFpUTjHrXpLhhILxeaz2ZadO25Vfy
pJ8UKi/oZAjXBPTSxHAHDcGihp5amAiZIzLmz+jHL8U7x4VuCiHWq8ktbKqC0uta
HhMVakfMjHetJwoZo9UgEqd63hL0TIcusY2pdypQWbRL/xdLiX9y7LWJwFIbxU6S
2OEQballC+2S2oxeA1mx28xZlbDpfXOrQsGFAr8BUV0OcagK5ibr66SupkKl6eD6
wkZk1fQufqcd6dlkn2XDwNsRCC8h8jwonYfEhC1aW3CwncOwgpkN/2VW3voFEBzI
grLPIl1JACEnsbcIfscKeBpmUc9mwbuq4b8rvqV25Dt7KbD+xzeJFQ48htd0sxKw
8iGSLv3iB4et2NZwdbJ9m2aVq1ZTjHYW0f8DfUy+rtpaT0dCY0yEcmQ18cryWHLr
1U1qaFVUZPjDidm9Lkdetm2Pt70+PnM6KgrFikcqtMcpA0DPICYoPaK+JNbm0T/5
tKsyxcZlPoPvQ6lOdndujQhOzoq5mSa1QH+52jriJmXmZ77o2on0eEp9uPhnwGZb
bxViU5rkRYBJQzU3a1VsvIOYMH4G0OPPnDmTF2f9YAeAtbZJkRSv+BjOHvpXhZpI
tUiVzse9ll4pdoe9OeJgG1TvTUEq3rXoO0K2mWhyErpTemnfBCkCQH3P1bd2tWr9
eXvQwde+F9WjBP+gkzDTJeaoLV+uWzvqiYCRbsRNqu6qiNUeMC2qTQyq1D/PBZx0
UC102lzV1gPKV2PH/6boJbpRbYCPF5dI7pIRp/Ga1PekenXEA81LTM8MUL4yWnpV
dRgqcxW2Uj4kq4nYyysAnwTgjYEHoIJz6DyI7nR8N1OZsyUJ1/V4Y4wZSmELPTVd
ky45sH6mdPSFaYDFpwizUIl4ateIQAPIKFN2X81QM4KQ2WdeceZjHG3qowZnroTq
ywIKgCroPjXRNP25KdJSsy7ERji8gKfUvq7mR3TiIMz7u5RxIIEb5W5WidgbeHhJ
oPAGFcq6rUIHU2o7UD6PGuNWUwrQQvTKcftGr0a5I0D7GcrKBXpWvBcRV7HHYPOI
TGWYUg54fDASVSUr+r5O9v7/yH3CxTg/oj1NSyPIhEpqW3VUlYGy2xGH4NBf9Mdf
r0VbIcTanc9J2i/Z4PSdx8zdHH1XtkXjjK+Q4ZyTbgBWcK25gd27GbnvXUvQ1eiA
MgdhbwHbWjf877EJCKyjYl4+S5hpzXgbV5JgdfHuUT/F6z/vjcz++Ro/wENhKQ/Y
nsX+easTy+B68QpafNov9mlIy3ZIhQI7JfgpU+M7SkAPR+qJ7eowOCDvBKYIq27W
oimj+L/N7aYPtSfpySzqoCeD8xYqFSSBBnf4CxooyvMTBuS83YxhsVZ+8jywcDRS
PfERGXw/ruPj0EnDX199mj4fXxJVSmOocOe+hv31dA3VIq3Ea8oJbKnRcPVvl0nT
Qv4Wrc6GFEUm6SEvd8qHc080GRvS/d8dYVV5ImMSCzE0b2vVIyVMq0zfCOWRUn3X
kxqfiqyHg6WtcvLvYokN9Hpq5FubERJfoutaSM8QWkTcjrheNpA6ftvNf9Z45B8U
xcSNc18sCDSPoF//T00k9ZNortviHljwDm9aQQ/bHiPKgaOB+c4X2fXgeSnIgkrj
WE64mdChNfSoo0vX8qGbEHvea5vjUL6mzuKGLEI5hzNAD8OZMhfcjRKcjU6cBKca
DRNFkkuO+HuiMVefrrEO5V6xeUfdlT0/mmR8Ub84ipyTZoE4NGKVAWamc3H1ILtf
B7H/WSm+8zKHjIEw9+Dc3vcjwxTo4fghn/Cw3XsMR08c6Bpu5aF1tpvGYrYp4BHi
ERQT/NM7XwVzp3r5B6lMo+yjc48n48Gu8HDcdGmRmxBUUZMY2daWNxRZMRj4O+qs
3ZTQH1x2bMXEBSiwvOqeHNZ5MyCk8n5IaP329mrR25OLrGUzJPfBHcqKA/UlQYKF
BB9PcFBGCaHdFrlqTEsOA/C4u/aFyRoWB0hycA7H4teck9964ody1+3VTDGndPNj
VhmYo1wKeej3876yCDGwOyJTh4sduUmpMDebElOkV7jdzzUY3cvB8Z5HQBYpFTpB
w3P1e8rFHZUyjAxA8vrFt3VZ7EAz5e/v0J+52Kolqh/joeJPok9emi/4aQpEEfZz
cU37EvVAQQ8m5akIAaEVbiHFnq0yHR9xVxgjvP1e8Omac38K/Z23YrxVfdb6gnYH
SILVXV/Bswnes0OBZ9xq4Q0dSRwNipFzcN3ar0sC22PNtN9ao4EF7xn99yY8OI6V
YVfrhQao8z+sT0BnodefyqVAK/5MAbF2ybnRJBiO2l7slTs6jSCf1bc/Ll5CPoNI
bPJqQrkWRHEoCn7uFzBt9VAQClElWiWTzMeTavm716ILc6spLBZmRqWQeCQLccpc
OJcAI0VgR4PTtFBDjUpAkDql5zId2ir0xsUF3h3cp79iU6iP+NiQtWbcyMOAPVsN
sviZBMtjp7TrI/o+2oDMH34+kNyfGedMolnVuYMZ26ESq9IVkLvbTET8Xd0CSl52
KkGjIBM6f2v+eI8zEQErkEq8lgRUx78fesgTGHM9VLgbmM4DGUTTfEozDTJamCAC
X81tUHjbfEmbdcQZMVPjmAuK53KyclP+sy81qVIVwtaOmeuWmZVNerfhaJi5/pz1
fMb7zC3Ndepyn8WNCXdiTCrciFs9ad1yV7OwS18zdxhM1WzWzE7im0mt/getuLbT
CxyvBee8OpS6THk2hoTKW1zpgDHGZyGiK/xk6PLt7wQG1aFVQ0VH0Cv9zjVxokHr
soyaOC939yQeyNJKs825xNDwRAtpVgydwD0nxRPLqxcg1MOTBPRaD3RLglN306mx
ZXbCk/XxJMfK8jiKd4UUph9R9BJhuOLvzcbLJHtyYm7d9TfeEsvIMEZuI+NFuY6L
0WzHQBgda0she0U37zd1m+B4b9o+NtOYjwFNaA3XWCqWfYyklzRpfWN/9eX88V+p
7mHOP38HqFtVJ+xYdN7kk9aRKBwNRg0lkrZFBHT6+jokU/MhJ3zfHNcpOC1wUoKF
iZUFlM/i0cEyhONCxqzbX7HWKB2RDDcO5o20tEC+zPeHk0CBOpNZp8zNMp5BY0ea
fd/4laQxAK/YK16IGGn8HjpWNVM08ZsRNwPEvpZPve8ldHA06FyRxvy/TtGjLEyW
NsUbu7pz+h1f/cEFmOYERiMuTHPIo5BTV04ArvDjPJi70V5/Nh5JnyoOfzkrh+cV
NWqhYM+PkOwPoIRvkSWXQId273qfaqCZHe3N03plZpjsN2irupFYDxFduUqxTK9F
XrOeJB+SNcwoxRxXcgRkbe6WhxiR8X7z5od+gOOPbeleeQ6drhAW8sSJfg/zRc8P
53lDc2RFmvolhutnNMljs6WJF3mpLlYxU3WF3ED8nnpl/MxUnIMmM+a3xFs1Y3GU
p1rd4mdRbdnsqm2vMNN9XZCgg/tvyo6eoZYFu/CanR533ClwfnJ67BlHfsDrNBeL
7LYBKa9c4AhfHPCABcANplOxDxDL9itJGRgsNkY38EpYVFGpt2E530ADPAzhvlnw
aBzK/G/e63uvZrXDhrVykRjvxPkPIS2k8f0TGocdnRHrAY6AhsH+erMtHaTVTeHQ
T5gBbMcuCNFCGUhXHa+GpvmeFv43MYO/GkPI+6zat1K80+qxFJXpJ5mbpodQciIv
S9tBqe4EAc7NGKsNE29ffvAVL+mzC2Ejc+BDKWnud5m160qIVvURyMU8R5P9SIXM
/r1tKGJX4/AD6xWmseE1F+zbFSzXYRUD6i1opZmANqP1SPuGDUrV7HgXnlM1wjNv
i1Tph5JDKtanVWMQ0fERpZkzmIFQ9lsipIWL0OSolBBKb/E6FF73f3QCxYBi75f/
OM02m2BuBIfFVJ30TLGj6mV1KWReByIN1wpGtEB7XU1737Rd7IanfxvRoJ25noum
m4+l82Pk6sv5n8Kz0Fc3NEux8rQCiLpyGJNHYSThSAk3A08XCcIzqnyHzvdjPhFy
Y14HcGW82HhtzOp8tvg5LROiluMFbq9gqMP/D1bMlJqlSBLPUid35gbmG7rEZiJm
3ptcT9CO/fyAUPuA7bvkFMRZYg6mdJNt2NzCmxe8cIxiEOo2EQ/0ZQaxxS11MUDQ
9qKvMSgLXyRp216NmnpCZA/lQIC61BwTS4fl6aOYXGOC76Xu3QlIrRoZQswQJH1B
ljzrXFd/+xX0PrQ5cPgvSNOuVcyUTAnHMAxksR+41L+rj9E2JrCGpDtx9GhFpChb
2RKrTDSz6EI4PjL8lKQDVVVjp1N+6j4R9pqKRNHJbFjcHgQYo4kNkz27cwN3esny
RFPH9jGeMdVrUsgMAcVP6bxfkTu9+RVGH/+RTvFXPF9nTnR1VrTSY909Ratt/NkU
FlUmBfvfttkjKaNqF+M8CkVG9cQPKH0EYEQOdw6NUkbQWGZVhpvmIkDVEFCB62y8
jmyzeeX3BpwM2OzLV6eyTcf+vnYL4HTZYZ7YTSG0r/ou/HCsagQkIUvbVBSje7Xt
5/E9X18cy/xkIi/xxd5kR95tTE3u/3W653jr4Fx/fZzChCyYTmA2vT3jKdQ0TsXA
5Luvd6FwRJPKVuSQs5ILDMX6rFFU1tKp1d58D2xsf0KwnJONWIOj4Bfet7MnTZxe
MUvSc1mT7frWqeYDsxGs9npB2z/EOR9ez7qX5UN27oIK1f7WVL68cWeGLMGsC4vx
pyw3Deny7K/rx0ez9343imS1qC9YFxpRJDkp0uSodOQGuEc1+HqHzmezidEilkU0
2PA0PS0GTcnOFxx8qszMFkQ7FRZK3pUADxudZtZjt4/Qy+RkjsPBfieQJi9fbkLr
CpdWyvVTW2aRyOcbfLyy6Jz/JWzocwNtRcC+WegnvrMYU3A9OPzOa0tf7i5l81vg
MxEYTa8s8wj2zET9l/VWeJ5Nc7vuU+moILeohcZ/gklmBxsdXZp3pKN2wATOdn4H
2zaFanYxyO0Qd4OB2R2Lv4k9UwGo3dA/g99x7gb9iXgLiI92RUuN8YBPgdZvG+SR
TfTvNOqo0+LgM70Hn79PnRV94oNLWZ/g4grSNrTPT2wNT7E6UxaSaxcip9suMTTA
OcGAgbzY78tw1RTGndrYzFK/Mzo0kJjTr82FQw010RY9tVd/DBa7YWorQ8ve7jTe
jl1AaB2VkvnVe+KX/ANRabaoWRk6DzBBatfRJPSMpOdgeTnpjmB7aIt0X5+HyJ8w
GEiaUbp/06LNYXV4hUag3LseyDrMCimwIY5R9pXqMXI2ZAHbBJGfmZWK5JThVzT4
Iu9PT0vVnwpfB7kf1ms8YsXtUgi7qrbmPRF/lOD+ajx5/zbTZcSU5EBflfJen4d6
eQYV6FqmzkuZwr/by9fJD3tQL4wYonWBxoweSlzEQKV7fOcv4rUlBTEUyprhqhvt
Xm+B4ar/Iz3zJ4IA3IiwxVJQVT2Qhd68UMqTd7jQy5NF/flK+JD2bJtjxy+KRflJ
U747NpMxm/V8fMHkHW1eHpt/l9atrrrAWihk5+usYUlHoTUIXRh3QIOn4FPc+Rua
Hv+5w8dzzplcvkqFropuzO8U+5XtNjkmY9kQYURFuNL2SQAbc81ZFHozhC6Os52y
SAVC39DOXzzQdIVvChNUvy/vDYeIz95Q/J+WgQrrcqvQ932d1PjstcwkwQO7/T2G
wqdAbged6I3jaSISYXys3p7oFtwjwi9+PO4O0GylJ1szfRl7/BMXTHCWvytrnUAy
R+hZqKqbjIJYXFesfAl+pXW65Gvb5V3VJSMbc7+7hLc3R8upuusbV+P4F+FlPR/a
X6BKen2qFcz45uIo8xAVwZZNTB6lu41iqssqHt970KGxcBKO7oIXsUHdE4hUDRwU
B0n11hS6zEUQQ95FOwg78JevhSgI3Qo8nBRrOQxkqcrty6cl6Xxzdh/z+E1BymYB
S1hQx+FPbNPWIOyWzMYVdphcKaTqCuCSCb4KsqLwCXjJL17G2yuXTYB76EOaKhAj
13O5BrOIYodO1vIUHSjZ2F0mkhBXRXSM9DHY3Q0nAzhxOUPaHDgj2xIQ7fTxsPAr
qKuVPw+25KUpjRjvgRlNodWN4TaQP5SqfqXZMedH9Om5Xs9gLdUIHMMv0Mg2v7aU
MJqtcYyF494fJ2l0amOgDvQ5fTRlqee1gj3zWchgQGIB2nkoOGnNe5PvZXCva8Pp
dC4+MJOuLXqxWqnbErJO964ZzWSKvJ39/ODcPAR0QAv+0vh9gKJxee/NN8J8MxiB
s3jaVFuFupK3nRhKfVRoRZex8TElgo3ig7jUx4uisu5GE6+0/sdIgMXy9dTWqxMR
k06rx3RczT6fsgZ0/Qn4EkOftS1OK+q1Mh3nCyvCFB0gSeQWVB9XbQwMqetjZvbc
EwcyDRaSZOB2lRugI9EcGK2rpubrCXKD5GayKuJ4GmWvzgaBbjlMLGjdTkpm5635
Agr7hLNpnFYGPMTEU4QnAulCy0/2wOQYaUwp3NoNs6csDgun35zJ6vtQwPkxi0SD
pJk/BzVsM9ngB1vaaR/xIF7fSvE7RhyjnLiwTHW6Pq9ivtZT7GVu2TimYlo4vbwZ
hhMkiAnjrI2HaBuadTlt2HWhbVc145LJqyEdBYylM77osC5w1SdILvrzxdetrfbK
WbinVOzNIpiUyQd/+Bk+dxk6aKgZiVhcrTcrv3vN1LzEAj9RvRaFcPE5K91XJzS+
Zqs6thCLBSP/JxeFs3FPorIiExyM8l5NnRRyNRr7vmO6diRXnjswAc1l/a2G8OrX
V4yF0oLTXgsQyfBhVvu95y9XdE6HPKHUbC8hR8ZhVqBfgB/sIp9NeeYgHo96AG5B
7CkPW7nELCzBAaZOSBb8oASWKU32Ljs93lFlgJvhV2uiEBgkd/K4fcpR2cZP4Sh2
n88LdlVDsUtT5p8bzQpr0/3tvzNYCPeUQpDAeREcw1XR1E/Pf7JpjSd/6L8LkvSJ
J+O2NOxDbFOrXS/1FXD+whUG+5psXrGE3ZeGKQKZCO4cXzH+Swi6m2aWyu3yoSc+
IyON+DBQ0CR2ml7zMLIZXVmjA5JCmB6w0j12yw1/rsbYpA8jD/XwZfVadBjE/yDG
dzBRRxWO6aiAd2YapKSlNZkmrWCJ6Ioj0WXRHHqBNI7CngKaZmf65MdrSBZkZ+ma
0QZmJbBO1Yo9vewU+GPqI4bz5uznrDMGzS0chU5JDayh3GszvbJFgbQysgfY9UCe
DINp5IklP9sl4SE7giilJlMRkDxzB+k4XW8TmtwBw1/NZwpHHeFBVDFMMYhIhErp
2a5/NQqLJrVtcep+pBbDpNJsm2JPqoH7krOr+zeazLaBF/IBVfhc7cS0xWDlx+mP
TuACTCtSaaFHpngW9ZWjYYzQ/+v7IoiORYlamsCI29J2vktb04z/4byZrPQz/Fcp
WUxAf3GlIZJ8VkhD1Pi3H7B8az+hfMe+EpdaZutwcBd2IdY+0zDtOa1OEvzX0JuO
+oD+vXaSnp6c3xnENe3fKJuMKWw9JIuow9mFyoa85g2TsZOlFQDjlO6XleMi6x/m
heqM9Rsfif23tFY278CCgE5jukLQwrpMrbv8CTGRyfXxDmqr+WPTJuDwAYXsMO00
Ytr7jQVzTk99CcBbB/c+gqkmsAx+c+FETEDFaHucbDgI52fVzS4xz6Ij5f83/yAi
sVSV4jo6JcQ0Wc0dFwQX4fpXN3bDPhAycBkUzoCUxz8Fh5xxXwo0rxb9cCjkxQpq
dRNW5txyT2ULgBjo7GzY/0J27a7QcGChBRNah3drGZsxH8naU+8ynkR+WmdlaKxg
L1+KeJDDYdyTMZM9xBtacR6VnNctkE22SWrMI3inMFYbXFm/MDtMyqdmN9vtQTZV
3rpI2Ac6NOBxQcf67Q/0PEFkYFJjSR9SYzmAOQAUbeh2Tv3+FHfrEU05TPVoyf7F
bOy8TBRlcebZgk79xnzNkJ1jUO+MkWwjvOpwLrqNAoAcFyr+qwk+LnqSAK8icd2l
DYpWYrHzSxiepocXC4c/m3yXUA8QaWcbYN10vpi+S8A3KPgF7JTMQ8JofKwXshhA
0p35NJcObnREGPzSOSYUU+QGTrIL1zh0MFEHWicWfVDJZSIAZyncV06K3D8KbZY+
U2Stpstf5Sv2UTwCQQADrZA9Tv7i6x5H9lRT4ipFdSRHzCFdQXt63lLo2VCFKm8n
t6ZqXao8Gksj4S7fsdVgmL/2utmAJq5upiODCofSnopDCBXBLpNXoRfnQA6unqvn
ByoRZWrBTTTNxJeqWUI0IakRgeLoxFasVqm+jXgFR08RPfSCrVan64Vtm4Rybjhf
NPYdTo/XfPM9TRnnRNe9TE1v44yg4yrOhgP0uKWTJLci/7skivhYsRAjxDG1fH3Q
Xr5VsqZNwNWT6jDo6GpNkE/olGEXi/Pc9/8ud0DBfz7H6fooZahRsBdRi4hNzp7O
ZJ4+xVZSDIsBc6HdNk87r0WOQ8uc4z9bxQGvszBH4fWtc0rGwij+jr7A73zga1o/
5WjgCRyb++vOM14mk5P2Vqs0xXBYDaCCJUavxd0T7zvhG6VArfM4RiasVkFwUzlc
g9HO+z/8zwpK62eyEnyvTepbk7F8gFf1IoIrYMqsoYq6RaWhM6ggC7ujdkZLSZeH
W3np0vVASi9rpHNkvpGAtE4aYbHGrFyDwjv7VdnPafeJn0sk5qxJHNHWjkfhokKZ
EHKkbPyHtbEisLi1khRPCZYxgRb40Zm/EjcbCcuX7PAdLDcerj0gpqRk5oB7uXd3
7LVeAzoh9Y8aGQG9XGUrO4o+YVC3Y6VeIOWjqIz0Sn8Nkrl0UOSF319mYk9cajgy
w1FZuFnWu0Cb3mUSFfFTNJ3qdkwrczISAXzlIy6fgXa/qFWNmJ/Xal1DuJIlA0Bg
JYQUygkfh3MGCZEUxYbvYzq6CzYkwn6CYScoVAihcv6cK+2xONuJGcVqtR4KmXW9
W/kcGwvoYkeTgO/ORGro/aRuKhUq4wG/vz5wnn2zBxN1VhoJXaz73Ub6zyZ2Htdg
lOW56M//LmgbZyfv/q9vg6CcJ3cCFQHp5p5nycKgpEoGfq+hqJGE5+x0RBpI1Nrr
1Pj6etDZN7FNQlEVJINJYWSdNUPrtPX953X+n/UBuuWqmNhuWwWbC5tfwV2KUSJc
BwazhhWM/7f8vkJlW6s18Z8al1ArMNkCNbIEvPmu4aVAXjxZt7Xn5SH3k4w8IOXy
GgVGZvqPm7hjZB84bdYgBqwpRMEG0jpXCMqOv4RBdBjwSPqc8xVJJqEYKUIcNS9+
UytkyHbs3OEjvFlMqH9sZIcE/yYe2AZYD/vWy4zMVFsMidNUKdqta8Zbyn/chaA8
E4T/39qsZtDiFa2rosANBLnl+pWUHQDX31C+STwVdtU5+vBM3IRTlaD0AAEdPOhZ
dtwdwbQFxZlfExepFKINHJj6otbltrRD8lY6sQjvD8+pxIj+sY5UtvZvr+5axZEn
KS4Wf9uw2aSGu7E+eBQwzc2bumN2XkYzWK/qjmRt8REhAn+2motif1xKJ6kkYNyO
cIm7pYKGfmzxecZtNUvTQe6tigwmOvlQcLiFescIjcQseewkc6MkIv/X1dAFPhtJ
U/7RS+I7xxW+/rjD90RTepexTedeyMqQNCmBbYP3PdWdVjhYyPG2zQCFC3k/7D/C
ENx6+nBLHolA0j6K6qmyJ0lRAiNaGiExVvt2Lydx1y8YO6n+1fgFpjeuaUrCwvzl
/3Jb426OboUkBkDfei03gPvVyqgF7Q6FXOjh/p2+6zbYRCJwRA5kMcMRb6F1tpVY
pVCPuLOdzPmmLg00YW/wLsSoPKiSQwqQ499NjLXltz3BLGx/gigOpTORCm2PhqZM
bmSMRpp6nBv6f16A++67N8yHIDXBnkQ3XEsXZ4z4Xe3Eof6UFn6xDVCFTk6C+vNJ
acofbEa9SCmzMlmcyYQ/OAExFpMi/Ph6DYYeJQu3CHwP+GDtpp5BFdKvKxwyj62Z
yBBXcM0ZuuhEEw4UsH8uMw+1POSyKJ9+Y5pJtQ+RNATDYfZhzrv+z2f+asGgJn5g
JxFbzFMcNfwg5dnLeEXb6PXGqZSmI6NB8dlmMoczAN5OA9EqhzzDLBlt9hf3wQWJ
3edMTSJ6vIB6FFCtmJ/w5f/CTkFWkQBnqeoHKqyyF1D6xIepAD2Xj1/LV1hi+D5A
zy2A5lW97pyKkPZRSDD5SQDYlkHtr/pMxoQmNgxwBkFQd5+Sttk0VA0ETkR0Cpid
vCG9SxeM0wZUWQlyXbiq2WWX0VbvlmcKuIaYunX1/XrwbIO22U+BOz0BLLacRHLa
ydefTZW8TK9Zznl9PsOUd+Mg3mbhXPRLeO2ZxE4uCNlFRV76THTVTa6LaqrsKCCd
2sQjOprPx8sldZePZ82wmzVHenspgmaYVaXOU72lAFU99DVHpvg2VHwQQQFaRxHV
yC26WMSa4MNFoqIkFFyvO3SvJ/FDeedH5rV3+9Xtk3ki3ngTCFuzMXZIZpd5371t
5aabAyYDwQjT5hJr17iLJF4Xejv4TA8aB6AnsvkWUiHkyvQrFwpKBlx/y3AiNMV2
9W1/WrnkDsXzStcdBOBlsbC5IpUa4kc3yZ2HFPfIjl+ldlTXzwxq4Ysh82jkLv93
4gkPYo0hGdKV6vaKl/8IjyqWCMkpxhBNYXiWUPWbCcqSSRka+ahI9LgGvTIT1q7u
a7ctN8B25tVQBQwyoye6RWsHR1PaqnM2Bk4fpgnfl3as0SdZLO6WXmviE3B3i82J
tOsu9b5RAPqL3DupMQCkXQKIUZCQkDMuSCWZcpjREHpRnG9a1b//ZCNRzhn9yjBk
bkhqHQL18Pf9me1QpCDDFwNcMZi5EQ6V9MKiYUMAWfYk9Uz0WueIDZGzCt86eDth
GR/LktwD68V5txCAQWtMhbUhBRVvBIah3TThlPmdr5Cd/Wnyh7cFOCyC0SO5+0+H
HT8A0Z/DTcXrtIRfTGhOogGMF6fYYLfc/O65XNhTY47R/8bsij39w+zhcO5DlGLX
/0ZctsSP5Oks+QzXKlo9c4MuIHMvji2QFm0OpFqm5bmUJ6uSGFe3QZEJCt/sl2JP
VG+JP+Dtk/6KlwP16B4bB9x12XLAKfzXN3Giblu279O5NICxiNfJAstDkg9y5ps6
rngetfJCO8ZWAAkVGjW9+SkSo8czyHAllttfQWjnLEMbgxb6CHr/K3f0sbbrmybL
gZBQRTmGQXQSDoEudxOTC7REHSpHjlw6YsPFIjOgwuziKu1LxNkC9nHZAv4jXC+j
YuvbVEYxljGkGiBfiaRc4eAjdaekDsAH2hNKDmo6wUagAP0s1iC563nzYRxzSE82
/vzX39hmyLjU37b0yTYMDO74UBYrjiouEgnbPt19/D05rUb0Z4AV/dL+9qii45bJ
J/ap+1RzDy4a1DuSlCmgWF57SHXd3DjIZ4e5E98IH8vW/OkXMaf70Dy5TWDDNLEJ
jbCg1KBQXDjdTIWb9bTyjb9Cz++JuR9rEiMJiChdQghNR9Z02h7r5jFNTUafRPqn
D6FPqugxb0TDFucazj7kZo74paMXgRZnt+fR42UBiIudc7FlNwsz5Foj0pDl7NFz
Vkxev69Rfk3VP96RmjLYbLK6S/GNuoOX8CLI5In6QHmzhc/Zj/t+7hRkqtJXLRlK
d9qwLdqLLDFu5PQAjCEVJ/K0I07BOFiJRdu3LxvcX5RbZjHoiMnuGnSIjBricb1i
FHiJq6/jFWHVKdPAIrpGPXzzHJVNJ++FM6iOih8uDuJw+CQHpHy4D82Jp82NCguT
AyyCYvKttWBr55awfRM3kz1MEGy7OP9d0sVodWGWT3TetRlS2E58HGdripNp46cy
TwlzT+CxcWUBRmU/ZVslJ5Co52gRL4nUHFUiYgFsiFpBiZhffuQyKnaX61ow3Q5y
vVWRt7MmFtf+XUizOn2nF2Mz8Ek+WD+L6Wf/3lsFc2cuyQoWIa6cMf0KrNePiNgq
N1aCIw4IxdIajYSFj2BZjlOmDdfiBquWhQNYTuITO7QVnkED40H8YZxUZ0NcsFD+
BXhq0D0D59p268AohAqCnSXvHgsjdfwMGlYbrpVBPeTwesmgQNU9eHYzTcvh79CP
Jcszk2rHLCvUXWOttpP4yPLNmwZS/4mu4YHQg8+bIYUONWESKPZxyfs63gJzn5fN
Xzr+g3mWwvb6iiHONjPQfwfaAczVHCGTaVJUq61Lwp/woZwAUZWyrDMgJf+26nx6
IKauIJVgvYWal2BcyYT9ht4TRqCvqwWZU7j0fL07ugdP71s3PRRimQZPylLrW3NE
GgDoLG3V3HTPxZ2ANOId/S67m9OwfOX39E/VMm3yMB8Pq4uW4Zmg0QU7evI1YLxL
E0vhhpKsiGh1tnzf/iX2HFKF7KL/JZhc6DBvVslAK37FimANB6aNQZCK/E/1uI3E
d/kCZwm0lar7p9z3Q91GtrRqrNXHcLUxBZL2ZlWSdTwfqZOOcXLXjYKJqdqcArJD
vS1WYzaUAv5OV07KiXos9P5pCQ85LgDc8XXvALURBancmPz9+f0Z35JhwQ7Ar2OV
d/UMIZXoNz24sDBdYatcJ0XGHL+NVDtN8olJKots3rEcGCKZbaibhrAvWNPN+xBt
vco9gGQFzPUJD0CQIlJE7b0keWXJ9axJhVilzFN99KschhAEwF3hMjYrbok5qulW
TODwU9czdT0Pvk9mSkWfBSoIxN29+QSVpfAKrpZcI6fQoNLW8vHyidBmIsf0DIZD
VFF6fgxe++RBA7fkZTA8P09rxzHdKwcfy9/rmXG39jrQsAjvybpkbHDohEXP+xGm
mIpzNn3krzHzELeROAaFpaFHZGFY733PRkAtuTilDvZUeptWasOC8oqN77hWpNl2
6Hz84HGX1Sz+572Bbm3Udfwx9dtxN63/5iJjv2FKySsL1MbZBKsZa996lcEMVnai
ylswrKwWpQ6YR0p1E6NGBJRf6wAS2Xtot7PmZ70B3mF1bHdrYl9CIaMVSFxGX4xc
ToakDFkAoAmj4sLS4mlHZFOoLFSSdB5+6n+hZ38eNRA0UXv05h/4vEbPgQGBA7qO
LJHzlBiI/SCz62uoS6LQRXabg9wB0deOrgnE4uWE3ePh+cidZs+lVXCjslCmj/vP
igDxFasUv8qyjMqkBPI/eG7pQm2xuGhO7nEJzxGQugfHf9dTRWbnXRPC3TZlGrsT
PbMJhQkGDYzuKZx4xx6CshirQ6dVj9cqMHVlgMyQJSenHlatSA/5EDJBPz45Fsm8
38J4dl1hm9TpN/BnxuOovqQRphm5wAXByjdX2l4HlafvI1AQ1I8T8HW5SWKyFRdX
7f1ADDkqhJf7aLDrd7z9oPhVXzd/xZ9DH3a1Yn0eVTDNgEXsLpFEGE8GYuTXr9L6
c+REKgHlEDrP22duHCCffWqTlAd6BgJbf0QuISimw8SIX3C+wzwRLlXxolE+WbEU
VE6PoB94ElpE6WUTNdnzIgbdmMpPwOucrPbiy76DSLQ0I/crYOW3VKKBxTnUJlKK
Jeu/Eaxu+9aJDmnWWwkRKgSuScFHrAkvlfit2CYUSeczyY/N9rNTlCbgNR6by5d1
J70vB9mYyQWBEqpPcsWcQSi0kgpo/0wR+L8MS8fPIiHxC04DySPb+ab21XRMI+m+
DPAE8WwpK8HISjCzKoLxGbSSj4aqQTXSf4C82GhwFrJC45VSCKQDNBaaRGLsIC6G
q2K/rBH3xi9VHWWMwnHpsL2B+SXtbFohA9oaA9+n6q5m75yr3D1uHXiqs/2mAqFK
vHUKiSbXkZiu2LsWoHLorNDxXqe15/bzHxQOwp7FO7y/MEUDMWGuckkivepql4MW
dIQC4rDQ//Ljj55zQ/BaISs1laP5yaUTuBvi8pjiy7ZpfpHoLbza5nsQPMO3UQml
Ddifx+tVRTR79z8mIIvQ+yz7/aDLCA3pa1lpKG8OPOJvDfKGWagaiJwwePwBVL9d
lBnGPdCo2GH3t039MNjHQGlnqOpkom3K+YF/BxFYDR9mXGnBsDmkYvudtuPmjzMu
ngOIWBB9WIE+PZBZi0QW52Mk3uFUl44p1BzDBZDYOUrejKjhj83qGziJwFLdrs9y
5k8+ONKjt9lPrlfvKwXSgd0zG3ci9LobfK+GZmE5MBNKYaxcnfQBpGqKBkPQxv+R
TJPIKnzluUsuoeCdjAWZg9ZC+JLTXHTVHPlegxU6i+aIOrfIwxxCTkL9Awar10gr
U4N8FhRBy1k2GFuGIrDfj54UFLnMUiXZwDKfQ280yb4hAWqdQ948Xe03sSCScut/
0F6/4+VIxhGhk89tw5Psqqz35y3WYlNfOuHLqK7WNNqjVBvNONgKIoYR6Bguy7+F
CWjlV2J9D0YRQTOdmxpWtNUbbHzIQe5rOlMjYxdZ7t5L8VJ2+kXdCecg5oSc2HEF
Gwc2SofSHrb670foePgKkqCegjKSafRzNimZ3qY9jjdc2jPE2lLhmHiHDzlKaaLu
3D53uwCHkNZADNRT6qGzuhJ+u1UrJ2OB35Y+PKV1FuwHjPUZZsa55bMYmhH5j6pk
it5RDTwA2vu/t12KUL3IcbvWXoY17F36oP6bhjT0a3lJs23pfNcOZUGRc6HqzraX
XWAjGwAEpUi90oZBNLGNqU++CFAanfdVgTSWwnA26T86mj7lfSERRNeybIhYPOhN
GF8/O8xNKjYJ7lRFXzFwjLH0UbQyRkw7NCz0iXR3nKO/7K9KOW2zKGG1BXYG0DLY
q/G0Lt6dD7JHKubixNG4eF4GFvaI036OcXxJdWRrIjos8fizyXGydxLYeS6NTjxp
nxtO7BILMVf1m3Go30hcJRrwOvh3yhG/OVzR49Zp9UFxJPwRwA/wdColhf3DlBpg
rtY2VeNYten6i+NnDpUMY8aRbD61ddo9uJfUgBQFwZQD7R1zSKtBN4sNgexksbLn
WSfHUeTPEC8Eq6Gj8QJa6Wk+/W/Spbbp8Y6tD/DtOEuYlpq1ukr6UITlV63l3MsY
InjwINqGANaVck3Y7bmtYXwty1NrjCyLevjqRP3oI1rYOhVG/Mvrnndn7rY4dRUU
ZL5sMspNNrLL8wdk7nAyi+S1rpj0DabPqrMJV6aZ0A96mqq0tH0UDXhWmADL5aDH
GxRthVgTR4n+RlyOGX6NWFZCGwmyVpFyAlj3vkypOCABxvvlyrS5tuNn4bHUSsY+
Sfz/sFlfCqzd3tkf2E7I2gRvh8dfTAEsoAPQaqr2GfkEkiV4NpAcafa7mpXyzpLT
9ZgWbz1MHTL6/I6fzFk+eOrB1moRDZMf58zZjKNVJS8osuGyN6LbwOfMFyQYAAfd
nQ5kWv6Pv6FvzRXse1edSnc3fcZW5sr3xRCGHc9FQjs0gKHIkNVhqNc9GmuRdoJF
73sQPcMoZMI7jkuvaw4/ZkVjj+tnT25Wz9Olme0HPa1VjiKDiJbU6iKVOop9Hyh6
ZIbUMzKtyuNUO1swLhwCmDDJxiIb0JVBah8u7edqGDdMb4HAqB+CHavrqZvwVlUF
Nz7yMof7aR0Ljb1Fv0r9TPskf2N7gqeeeXaTgYNIK+p6yFhYZS2faq8VGOnLYN9q
nHIJiCH++/8tTJ5xMCVwTjfBhZ9aoj8eU5622DHa8OIS5hkK/V1hSTh7cPTsWG7C
umQqVmyfZDla2pKVZO3NXpcm8NdNAEBGZQ/K+wmhUxMQDnKXNrUSa0X4O99aXZkO
rutLj8tBzJRdI89MqZ+NXvGU3rA+l7cAm0IKis33cThlCxwx2sgSCoi3pmfohMgX
EieER70NxOshcIMK7mXq9oxocs6NZs1h3X6SF7nNWvq2R1nibwoh8C+IBq+ddBuc
xsMtVqFWCyEbms36L+OVsHkBWqYRI1LE4bHKGpz/5NWK8bWpr47l7+b1sgcl9jmE
L3A/Ql5RvOGT93g8yHG+XCAC3xDJjWEEEpNAqHdodP6SAnKEnyMQr5p2MUHxbsUW
yIbzlHFRhG/5x0kq0ckbEsQKlRQEzCnWXpGgtYOTOKR4nYU7z7hg2CKf0gL1g+Jk
AN8koBrk14bQRANTa5Fx49TJF0ZtgdTyYaz3Yse/5oJZ1jt1t2w9xNlC/LqlVzUg
AMQV3S37F2rxSAPpQdOQ/ew60gKsT9GUNm+rZG3iDcZuwOUlNTL7T18oLd3OsPlp
OZACY2bSBiRV/RJJY1ibWzNlJEAzBR7ufuuBx/L58T/oTewyyY0aRhHP1z2NmJyJ
rriWmB9qeheBsUmfYtm0V4r/QllPNTV2pSTi2Hx2CH+DyWJBOx9AyWW6EiPDAj+7
jUPls82U23A6L6lTuS5AAqSsuaOBINF2zFPGirtijelOkHeaPBtoZLCHowavyFzg
LWm9PZUNOxlzE5H8SlerqwdpMGLn8i/MuR8x1sTERiu++obvb/ge8v3iOp5Mr74S
3XaI0pX9OFSno3uGE71OXE7XkjjqToQ463GnKHhMJ0lUEHEv2saPRO79av06uAFy
HakllK5RKwYBN99CNgqzHErr4kc7gaPi6U/Tm6nLZw4J1qywCM5K9baTqIL16oZG
MdFLy09/zlrIMgPwDzYTutgat4kCsIvrHjRxc9DJnNgKb6rDMT/FTUFyKCttXp4v
xBRYAHVPrD1DO0isavxTwwaN9q8BqHU6FV4eTJaXe2YXtXS+s6NO07xlijFIwkpA
BZ5KEUJSyIlwoL1lyzKQYhNQhmcesAJZEqvFvZ4KqcgDEeEgHydvqS2aPahq183p
G1hYocc4L6PUNevdC7Tt8bG6QKVMo7/A1A88UqsuIfETyQfmDt1Uxn/1wufTh7Au
JUFBhx4SeumDvY7tSRSJ1EP3xkP+KdQ3r0yfIgjBIgd//CEDzMNlKqOjFIYzH8mi
POs73fTgcxnhrXPqJuA4iCG4c16cB5A5sOJbfp9LZvufC1Eoc/RBB/l3uhg6HaTa
mSNxrQgncjMkcZz1PNncLJ1J83NZcb2tIDfspc//yNukN7VEoZl7ZEtN47t+aj8Q
6hEBgG8MOMg+ZEVGjLMcF+GSLwsBwi/+yWTE3vkqARp1CF1kDx9SoAlw4O4fSC02
8ny00koRBXJ8qeM9+vRuAe/oA0cby8lHVyLmuum1jVcObTv9XcY3xC1M+n1nr/Td
/ciRJmw4a8mJhyhX+Dtouhww7GOQRWXeuNrGpfHiAC6QwcsmPqOIwPuLCy+EUIQs
PZxzgokIHoKHstgnIkf+4vYXjSiWNE+adeqOdXxCzHeOmfkpLkwiEbdatPBlnsjB
HTZUuQnoRrq3AB4BCJJz4jG9JrfdK6Tl7H51UD7IP0P3CjsW2FGEzJX+n8C0wW+5
HmeVJ2tMCcbc+xaTEtGwpmYU8iehP3jQoDr8T24CVmz8slE2qTdV603pI80KnXlT
1cFa8mbXRGdPunb6DQ/RM1fF6SB6ep9RmoOM3DICjlWEwX6gRv1AeOyhdmDpatIM
d+mmZzTpHr388vPkg6F1rlWCuJUYchD0pfzpNbm+Oj1z20v735elDHpG7D/Ojbqo
6KzpdgmIEhxDgcVZgjA2SmF4mYG+cpk1pZhn2SMDsZ9mY/LgSbEiPrjPPbIGyxo/
dT7ZcQsLqHbRnbRDKVrjlERiT9zRydAe4Ove9bqgzTG3bWtNccq2MNJv1PTYc82f
DLEgMrZTS6V2m1wgTfw5IDRwY22yQtueFYbm89rpifb5QUcsL6MpGreRNMEW/58Z
TSph7hwzOtZ8QM5C6O/cCXK1grcfTDF0oSgWZmO8fnckeCfVx7PteS9o+WGgEVlj
CJaFetaIK2ANUZj29zwtoF++S70SxlDgXoC27/ry4/05aQNI4zlVnTtMco5PwM2I
bxj9jepcWa9x8watbx4lW1fiA6/Ch+UkyhgTqSKu0obsb8um2PUDmjhDF1+Z6pKd
3O/IP8pGHfTb0xWaVC2w6e0M4JfK89I92GCFJSBbLqcd5S1jMKg2bVrqVio/sY36
pZnLrEecG19mBRcEN6oTyl9QvQwG/bRSDFl7zuOCVJReVyCuSc64Uae9o4at66HV
oaSw2FwlL9MFoMGfh44h10EVEd5ujszSbksE1eoYgH2b/64UDHMcYmwquAhkXq00
hlpX84yOmZoAWVoomRjqcMJYGWCmpyKvTBv0InAernj7Ke++dhQYdxrb+lBS6vkr
leMjZIkXNSm0o8M/D0duE9T26rNZquMVKnwzZMfKNAC6wggUA0NaOJOM6RB6ZcBP
CkYxzX70lfP/SeylQQJJ4s350jaXNXQXV4Io2NSbJFitnUX9PZcwB1F8fFv5pD0Y
va/v6q/MLxoRQXtLeWxExbzhHLkjjFlISJ7PyT7ek1EYxHNBi+xIUitfgj0y6/t5
aXg6vudn9AelyPe9+Jzf8Dp1A0sERG3nuL49aMho7qZzBhcwYZLHpIkO1SEXtkgR
So+02h8/Ur4rGgpNRE37lpCvR0B3P+YFKab1JH1LgEg9rW5XUGmAdnLvzg2RAtz4
ndX5c2GH0kyfGIFtHt859qA0P9hr8tMB/EUP0MzwM09Ke5z1OPEnrNk81GfbdsSV
MKFL7nmG3N6OvZL9Ac8AVs0P4RGXPFBqhKUKL5FDHlojFJqxRKdbx6kMWk026hee
5jE4fPBvcDxInTYGJvC1yoSwRgbidh9Ee63rmYSziFSgYlGjIUe2LJbRCMe3gD1P
upDiVCFoIRYbOp0VPTZsNKCCNyNEq3DDuMIZedGeGIUrj+TIqgEZ1cLFbfUGUyiW
q/DbleiobCc7r7AJQLE98Si2CkjhpAIrSAuEfxbIxItqCZcENkap+GjInRg0MMlB
bi9qllGvyNnUjQbUXLnzHJHLLI6BV5qGDESNL3/r+6H3IHzeXtyy4gfL2KIN7aJG
nVyyH36tKXRi/7tg2nOGhtttFFw7k9XzQLGSgXdN3WVo1NKpzt6QD4OFZBo9PjRC
OLoa7RdN2RNXCqF/Sb+J+6MbKS+MF9QSghjO6hwCDJ8TIKOqrX3C0J9Z9CiKwZiF
wWC5neqp2eXqzKBm+O9R6GViuCJKxr+522gFHGEMXx1BgA9x8mfEpnE4WPkRQVEP
xJpw25UD3pU5eAqUg+DXLn4GqmMW5UuNz8PsatBCDxCdHOEizhB0KrOxQjxxKA9g
WDx2Fx/yEjx7uqyhfI1oUXtgE1dnKhArjOk8ySaVHBszp11FODKsdNNyg08Q1hlj
IbY1UYwLvXKxbTgENAXZO5dSKXiFjfO2vwDsPnaQDxkYKxNqQv2emf0Y6Uw62tcs
nKT0ZJUKixQ5VMrBk566MZSYW8wuX5QF3CSAhj7ts/6fPikHgWQeULnPqiX3WUdI
CbxFhI0ob/xX32LyqRSj1+YH2P2pO66o4JlHPEeMRRN8TDUYNNE5ZEpnFQ1Bi8hR
y7NBJf/2WCRoAjLld1hF/dviy9gy9K3hEhcDwhq+pspNxkZMt0tI92v2N5MAxWqy
lwKv5GLviLYY9i5vtbhEfCyUXDYmefUrJAJiOjeQ1TPBpqKnBORJ20edhR44N9sF
Yq0Yg8P74r0zIvKWCsbCd3QEsK/qOJQUeQV9ycHGUUTPqj/0/S17ZjkAbnrABzKO
w1MQBsS/dxrMs51iKJPIEVpSuDlncvUZjikQ+cXboyJR2gK4SDQMGhN4Dh0D/YrE
wR85Fg763YCxTWSz5wSOYu+r1I8SC+z6m8gJgqyb/wS8OA1PzXm3nZQ+Shc1Esc2
I2MZ48x7bWLaCibYjIwE8VQczMPgk8Z3KEIBFXSjDaMnqP6feyzdMEUsTmTeLXiF
Q1Ahz4Yd9JzDc1b4WWT6K9kfAgrEGf9u9SaFCReulUuE+bBl5wPZ1yRn0L/gr5aN
Uv0mf4lnqOoE999jHWxRTZCzB+gZWxNPZe46l7EkS9CGYF3zUFcYMkwn+sp9YSYo
oK+cQLIIH7/BOnejA9cbjrA17J1t3sa5e/ef6fwWMwbGkNQ4KYIZmWq2CWIsHVb/
0PEUst0A3jfPPO9FS4Eei4Hz42g3+hloGwXzkr7+/XP8hc5+IvuMoidsNvX9U28f
NPi2p6hICrM0+AB/3gu6yVRsmcm6gbczIzZn8p6G3hcGJJktWvDOS4PMaTtp60Fz
/T0fZx5hH4ILUH7VNcbT8y3jP0adIV9qGqTbStDtUcJWBj98NUGqs8lc2z4YzClo
dQwqJL4Ztp8NcqCZV0wrgPBlSQUeOyFkBILC5YtkfVrxsHxt5x8xN9N7QwR4AJIU
RT+W6N2kIs/C2zna9YKSjsqRXPROvgQNHKIuxOO/BPvNl77YVYK3kiAMW3ZSc2qr
+tnB6MpsLv07bTgivaM+P+8Aoy4lrmxIubqt08o/leSe6cJDi7CsTYJHX5v39phx
uoD/bFY7ARF9iMr8yRRZXxCjPcZuSbMbQ2lumP/rgqCPw3pZL7jh404fzRVefhi8
E1Mp8ueLrAAdEUfQkskYcDx4Y1FiqQ4UzcfKro7yB1ImgANjQDYjeG7Ad6/GOGTQ
rSQiQY3lsENetY4BlKGRkY6Wq0WEfyFlkcOcR6eCbYFvxvyLW3O+fFTMYST/RyCt
BYVT/0Nzd7qmCJqDBKahdqd8CdIoEGWW8n5LiZo4U9YqtuIg8UO4cIXO8FUreyFM
EgIsA2Sxni89zu0GDeG2b4ukCcRqUwaPir/k73sJrFSfs1VwyGR16MZcnW6m8LXw
6tWv3k91plOHVPYHKC+hHGg9mbdwxFnV5tDhyK+bNOJ7hOG0vXzxj9PgxMKuDcqM
W3rfoeFn6qomfNWneUA/xA4U+ffc1HydX7KjSNrCbJyRMYHPjlTId9lFBQdyE1GX
IWt7ke6ICMsMxIvJC1DPtki0u42H7KOoikVIt72MZwbcd9xFsxRVjZD450pc0Uq9
A6OsJK36tUhSPGdlopZKv5laLnzBZkpS+JlYcXarPluJPnp+VCO/5laHlKPYV5xT
8bBNgFhyJHnJunRLXoex/RTWJX+cAnYJKZ8JKhd0Os7VsOp6Gf5ET/pIcyihE1oc
YWbJd4UxBU0CIIdz4Wm4M8FasjkDBSKYQAmOvATefl8GoGnzosgcuUVZKgi2PbbN
6eD2B4ja7zRFOS2jtNikStscejOQsiFQTiJH3yNBmscY2oaBjoo7x7x4UjsP6h9B
uWWfP2HBjn9iRtkjRG+Y7Nrg5dT9bFScAuMg0sP58XPcIExBnLokFlLxWqyIAGOx
uFUgUZUMD+I6YRREDFX2uJuwBsiuGtk/45+vrYlRYaglJTCIrXjUe8Ys006/b/GU
FSdOm0VPexLBFNOlHr5dXjaaEQLCtCqgGPAzjJe1swdunz5tOThV5BUSJYIV5O+e
hZ2S5h7smMOpESxiDu5vMToMBPvczPM2tYNfxAjFdq6Dlwa6zb3uWan0mo6SKdNE
7KPA/nkHjxgJaCqGf2A0/8gYM0SVbZKKy9Eb8VDZUTTALa4hJTL45VaQyLILvBWK
+L0X1qmu/96fXX3ItmgrPSB8jKCIND4FvNuMUDWOc7w/yoT+BwOgKncOW9bkwSCt
Y0/P7aE8zwa5DfstTNRtJp4dUmm0CvrA0nJyU3yDGfSpRyYc43IjTZUl5y1NIzr3
OuMmlb5lg4YdZaxqwe2EJTJ/DgKtw+G1Yw0qhXkXh+T0jzBJFPvaWQr7NdFN62ye
74URvJy5pEiM4+Bi30JxmCFTxk477sP9urYMFO+CNLqKEWmApI7YtYijYMEqmNQ6
wDP+YVv/1+iUWgaJmyA59cB9J4peH0VpOAclOlAVinHTAx18eMD4nO1CpaQlE1J+
5fYNUY2LZ8PGZfQIl6dglFvBqu5vAfzyRlUKfviPOpoGJlMwJcotRLdrxWUaqFCF
rYQj2ZKD4icyd7PATYyY06d+DV2W3J/Cup/eqRwdgCkFU2PBqYUsOqtli8YaPW7o
7IZCtplpobzgCTyR6GytTGy0c1T0os0epCFHDdbUgZElzgZdZXYMukuUDNuptyJL
5/ktvQHaoGUEIMKLzICvcqmNPxrKekSRvkWRRo7H8TDo1P4qENpL1zt90Y1MKFZt
zwepkAo5kSF1l2TOU9iSh0Eu8Bsp6o4J6juTyuYuvDuGApB3mm7BLwv70Nvt+48s
powwBXlkkVbdQAvpT6MHFBh5alCWPxAhPmqyeIj4AR4zqjCTv1MWLNAYcLPbxg0/
23uejNOP+NHvQdD0R60VaclBYnz9hmTlw3y6fpZsGovqkAVLm+w3s+ZhxhNLQHI+
XSNW7yti9FgEB6QvLslhz1zQGhELnuQsMrdZ0rzWA8+dTqZDcrc4jtJooGedYw8s
o4Stf04jBy3GmvP6eniaRtNVWo/mWM5sHn/XVWVz7rh52IIirnf29Ur4tkJKWPoK
7OfHdBl6KGqeKy2nw9Z+ywWz4oW6St3BR3nj7ZxSnqvIchPgWXCLMApr+erR9JuZ
t9bY2dEPk1QMXRxwLODmQMAP+RGwCburmODwZd62D5C+ZhvdqiJk8aICRT0HxX1e
U9b71tl3TJSUlvjTTq/FIfSJkTWkP2VMcD4nGRsI2BBt0o5VNYR2US7FC6JtV87I
LbnqIy8ELAA8wVBdAre81XYzQ7yMxcNnvptuXzE7Y+Q0jSfWXtjy5xXBuJ8CghbB
IjMKt5+xYhCHVhdRVQiwQdldXg+2XDnnlT2tesKp0CcTmpNUwSsB1bST7ilbL6cZ
Jjmdj6s3Eetj3q5Z7r/9bpd1ursNNDS1PpsX0+vc32jXvn6iBLffAICdTsYEOqVy
m46Fv8/WL9dyfub3J4MxymRnAunT8f6ytfFI2VJCKcy/9Zgj3YQHA0C8QjQEo/kC
FKIKxK3smsP0TMZNVFWl5OAHzbx7a58TuQI0b/dv2r0fxK/Va6BMcXjSqvmjfyqP
TClrKImZDkU3gb5aqGwK1Qs21MXH/aBvde3NnIK7ft/J17ginM1QCLSPZFDRukDk
OvC7xIbfsRyWm2QAxSi3ncE12HYUzoz/n5nxdRC+QX930PKXd5fxsuLByFsa0vrr
q8BWRdZS+RaNL9FEjr3SqoFIRMSu7JugL4jbUt6s5ev6YDsATSiFisW6lNuJFnrw
sOm2akzB9nfF4nGpCkpmkXwAzKpc0HxjRC0ec6p01VxptO4eNQuObgjbGKLFdDMb
2Si1s+23ANf5sZhBK21diX5oLtbVnp37wmgDXj0/h1GqqTHvc9lLfEpvI4KS6rcq
TVO+RpoUAubvBM6eI4AbTbZTvA76q1WleuZiq6BLI82/O58e5STM5zGo+qwlujj8
y4jNJhiYpQLmkQZkcD6txOCaHRb0R7cHODnBVCDNvphLrEucerfJyICr2/WgTlkJ
sxw0xENJYN5SjH7wm/0TIqgxHuRLPiK/ceSGaciDz3jkQLIPsG8ggrayzS29Fr4y
hfsZXOP/h0WkLr9/DgjPff/L372MKG24RRqAYYNCxNOTxRtqfGCOpXkcXZ8JLbIU
vsf+Tvr5msjtwsXM7YG/iq9p66R9Qa8wnEJbec+QoEXzcLVYkrqpBM5mI4ysKH0h
NLiRIccZCxPGlsH43a78zp0VBZLjh11QnhGbezTThGxurSFHVjX0ii1Rd6Vbsl8L
Xe/WfQo0kEyIgXgUc29ZHaW73bShaHSEHMf75E/mp0WAv36Zo/ChdgHbzZrFG2Ir
xDaJzA8T84e9fhwRJOevrN6unDtiFGYWJX0wuAEh5oIl4aDfKUQuSdBZikSv+mr7
KeR+ig6MdAlccdVR0svLT2ameTM6TNW61uauJQVsr3Jg7rT/X4VGRq+9+bsDI7/B
3IpcrvE0Da/pG8mGnICg1wEziMO0Vj/KLF4Z1X4Linev63/RWntmwcpBY4l9lHHe
aJfXBFRl4IcwMi2Y7s9PJi71PTXhJzJ8B5BNqtewoZHaBA6QM8q6v22ixVtFl77w
qYoYd31wdAT69nI7nMNdgIMoAl+XAHvdWCcAAp6W1k47GHwiXYRsfqusGO0jb1YY
7xhS5HeLVCwz3/CQD/8UK3EQKhT0TtiQgUJLUuHEZ9jYXzd967tbqKBBWjz0O+Sl
IRAoSV7+7poNtvP/TOpXWaQnwNxIS1epr57RJYZTNgCPOI7wvTdtVa5oJToW9cHB
O4yw88+SBuVLnyBn/nt/lV2mSfCxKQ/s0Y14hCOMzKrsYXgs6ca7NRcymgje7o7b
0YTF0s7FJ7Eb5Dhlk5Y59OyiCP1Y18ZtgVHHd6gHGQvYkgkd+MlAibmFjq7TAWHS
dkQlu30mUkEBwFZmbc6G6d/vXhJY0oj4CjB9mHp5/5kku1mhOfWbsOuKZQdxVM/P
sJWGCaaC948tguXYwd5cDM2wOoccqugdc4+v0897w4IugjYl+OyvzuJzyTn4wXhe
WPiOWv/+BpnS2eyTi5C/M0CxrVe2kW/P8jI8qVYooRXmKAjbWiv3o4WVlsCTRBg9
nHpPklmrTlgTJrjfD+g/I3ZuOnSk9jMK64SiweNqtdz26Ag0ag8VwoukxTeTRnf8
9OF+nF9C8nMElEVnfDgwbg49DtmtehlQ8ROggplrRci8Q1Y+nbfVjsRbH+2wxtYi
/9zWnRQJTLlTs8ypp8oFXSeGVezPU9l/VOY6LgUSWB0dI7EoUo55YcrtGFO/bACH
mXLyqBcA8zCEBPv2toLQuTMHLkUzIWlGqBA95rsx+JAsoPibzX74XZxM0thJJoIR
opF8hAQy1DQ3knGjrTRS/rJnJ+ty3OkfA67qc2TYY5hhkf1HubLTgGopyeaMtcv4
R3XDwc0VjMHuFxGufq3rso5lG/+eMnrdEgq+9bncQt7PFXsxWr4Q8kPlbQS9+nOF
+2tFAuqkPa2fEY9rEV/SNY35Cy9m8RFC/ISI8AuTfZxk2msysQ0hILrfhjOWNekD
da8ewcYoaP+QKYddr/diJYPBrJkIsv4CAKcgvXXFkHoHqRTbcXmr8xERFXLCN71d
xLYOSs9dhmfuvQAn6PMBG81airw/dcQTcfAtldNUB4yQecE3iRXK5KEu4Q/pRrkH
wcvXki6UzWiL6+3OUMZQn5dmwtqybj76r+9xKpHhT+R+uyaLOOeXbI/lJKMuaonE
kVm7TA1jigqq8Pq6vxL2CXYXVl9Oj18Fo0cWgEGnjGvuzxuwoTcac4QHmzVKrxEQ
kAaw3ifwnU7kELztVNDe3sJhyolccYpqj6hofwd9So9ZOPn9QvG85nKnT0XcLG6W
eLJy0y44dIQadLKQOTFvMczYjA7hUDdIN8DeDIL2Osadjbibs4ijogFsei/3uXQE
cm7PowIR/ZYMmEI4vJVUYbBYH27bfMiiT07g6GCjzjcYZMILfRACwmm+dM/csKvB
yj+8SyZ71qAyThU1ShnCCOSsxEstKavmM/XN5+nWdXlXGE10hRcANWbbeufQrfed
17K7cs317twBSq8UAyr/tQGVhmtYCWdxGc1LHef3PNeBWEJcJZJHSLrJ3JpQvEhx
s56ISG4j8/02g2zk8HEtB4Q6n6xj8435DjIBfz59EZtWBKjWIXD8E5tUBGFLgDFJ
ZxikMfD2C95KNAmqfPpfjHG26lehTohCA7Fs4vykfpqur2UWH/FDLeFI3jIhagUv
/hEmhwcGsOwz76jOV5HhYqa9Lj7VwVzPxrnrBPObY64RG3tQoJhZLzzpTdZd8MWO
pNovYsk7rMh+uYONUiCDei5zveATFqalPGR40G4rga8lpoQB2zBt5QMtrMYOhp7C
x9jiXKlqjOnnJzIMP2v+z7cJfPrj0zkq11QOI+ehEMEdU+3h68XoRyP063qJny/v
N4FRhEKXBJa0QKdQ8R+0RvxqLOzkUs/uruLNmpQTX4W2j72KBNl5/Leoeht93M1t
Oe/7VpfDe+i6oRUoYQ5qZ4qVRo84XBXDWuj5t6KzJmtUNTMloUUCHB+dXT4SoQuo
pC5yydODztCKFdTW5xocCleL5+qWaW02DFiYCZhuRp0lDiEpI3njpfXM1t2+CBk0
RE4ApKCE5/G65Iv4i1w8xJyJfDDlVOEuy5P74SK39eLEr/btoOFlKk8g4URpvbPH
HHkFF1w3rC92l7bG1mFaoq7Jw5UVabNivTLRaFeSd0Qs1M3jSfhBkbuZuiF/H1Iv
Z79xK8/3XbDYidAb1Zuye/DShR6iyK8D4cxEPZPHcN7pv3Te4+mmoXPoqSNhBF1P
HiWtBs+KjWuHxzuZuv2BVReiDmzyWdmLSoJgx5Jac0to4a3Cd8PdiAR2NbP0qXFZ
fqgTcR8FFt0I9WmvRikvcrK8SgkbiGjMnlSGD7T0A8G1vpkksPGxZOtB/j8WLvKS
U4XAyBAwp31a0gogqq/Iia5x4JFqTS3X/yzdcj6TjLADowEbXL2OTWnbI/WliLVS
W8nhrN5m4VTE0pwYoM6aHFP5+etAMIZJEf7uBMcVU2+rKBkLIRq6SupILPtU2pku
L2958Yo2YbucolT2jiU8qpasbFxJ8pjTr+ZnQQlhkBg/ZQMB7zLypZetoN93Kf8f
rW2wxnr6pmfaF6r7bNF7TVcbZOHXi1R0nJfZhtILx0k3eZhdArG52c4iwSr0socv
sdRhvca8rslt0R4lu8Ew74YXuc+ZLbdZuspRHr0QBf0Rvo9VgDpbPxMmarMTLQ9B
qthESml4ypuuZrd6aOBCTF0nZlSrjYdV3W3+kcdRv5tyP0silhGpeURxqb+8FpPK
oNHK7gJ/psxsYDonmu/gEiSB1dyTx5YnWsOvjQ+wtKgDeZOEGxB/D7FcCI5q1IFU
bKGJMUd7bSWZ4BKayQLi2F3I/C81aR5Y+BSBe5cNjgraly+/NEMjGYXM1JUrw0Ig
p8EhdXOPCLJ5DmKawYujaP5ywyltnzeCrUdG/uSG5GzDa449cftoLCbV/wDbMbJK
XSYyUbnKYLsBP4N8U9DkymwE2ZaaW2SbQcF5EQZaQo5ko5XKPW51S6z3TS0byYOM
z2bXhL/41mfiUjaOCnGc8ZoFIlolRbndaWQPuygNhx9Kb6SVDpA+yt1ZmoWnQZf7
EwbzWvzA+R1ylW3RpjqWRsCPzAa/E7UNNzPenYLnprt8UoWkiq8wf7ooDA2R8Y0v
wwAEJ1sTRfd4bV48l5d7pNuENNEVLQkO7/2kLxXR75XjzllNxA8gdyWZTkRe468r
4WrdYkAAyfne1F1rBNqqltro92ULBALHPnFDL1Ef8P+D2eJ4CrAVuO5OistjAjSD
HjtmeMpbb/7SaRMTHi+g2PiV3QJL7MmsH0Fe8z9XemgIvJ1XfMCyCO+FtBT3Y8Br
OgsFSuYemsci+PE/gKB3l/SkzMDVekGcjr+T49DqtmUZxWzfrrsfy1f4EalftJVN
LlveLBM8kwZUwBsB8tJ2+J35lB5aJtAswPdskMb6E3z4CZ/6t4HBh8aiVI05ncdN
ItPcA9aneWvUROSmgUquXg6ktOzvlNRu0/qAX5G+4OHIcCgFSXIyTx4T0WWStvJh
gK8aULi5aOXd5daAudqZMv8Q6H6u0M9ioXxIPBKY0Fp3BQPKaUD9WKaPZCuKpFVD
Z+FOyeM6L75ZyVTGAZ09pJKuFcAwudUsZ1FM+xQWQeokC13Eo6XgiSnlrt2ZgHDj
VOEmqfN1adSvHXDDUQ+h/NtwhkffbxBrZTBN6wQyFWrKL0izVY+3Dpb65P7BQiuz
NUBF6ArzO2JTtvidJ+E54Z4Q7gxtrrJDGTAnhRVzMl7h8RTQ71mmcTLmESTzWKXC
7Hdhn+BwqrDYxMT7PcJLRkIMZVZz8445R/0s3FeVxSu31lPyHkE9hBgYVuKjyBk/
2ms/1FRt+7YGmK90yGWgkPrUQ8yj0Q4xpPW1XG/29chTXtZ/TRWyhtKmHf+totWp
i33sktCiP/bnFRAitkHtxKPy4TSg2DnvkEJQgRyucog8mSMmZCaAdqarOK8Pnppd
NOrtnjHqYs4NZo/lHH46uttS1EfKbVuejBVfCznq7vDBhZiuspihk0G7aH75nmEL
qBCJB4BSXv2REwgJI4ED4dBed3KDXf+MIB8j2VZNqMVJceMXpi2qjn1wkTDaWIo2
rdozCUJsiPiXWHnpD/MMPVddpZlTj0FA1QpfvMCUueK7Q5+W9I+wOLYB/BwXdHP2
EH1Eq0H6Nt4bJe/avDiZ8uaEOwAEXkAZ/ocfHbEy29rcf/IFLNF/oyln2kOSGsRl
Hc+7qnHeeyTMq/hnZ07BgmJc8ZjqrMCJu6WCQZwVFov5DGI9n1YWV/yDIa/IJslc
y28IWBGgw+Ejh8XVDiQarB7FmG1by5+dvX5YRDmYkY1WQUiPyLvisx+CHWgSURmA
wkbgTRXJCLd33z2dimqb7WTcO3OCXSKQzCVZVA8IO3x7eT+bTMgdkXaa+K8BqSiQ
wpEjiwXJCMWCSkm5jhgQJJgbFXb+2JTP5u7Wnw1VP7NpKg/DAgXlzTELh7ZNgRm/
xdEeEbxMU1jCCxJUMuKKstuAcqOSEibj/30QKFPSdOJc9J2JycIzLNBXnqQnIC8H
NiNpUC0vgab+KX9dDaSpiMcksa0bSB0UcDhLg55g6itGtCodGDL/SBzkUXcWhkYD
NIica5MvP/SJn1lHUzkrgeDaYMD5lBm+ol8fn13Tw4RBx0mTM29RjTW7oXtMTrqL
3PqBUns1mdPRXWGoh54IqW9vppauvXo0veIPXhjiUGlYXdkmZ5mr0JWC53ysCgh4
8ccos+riKaaVaR8+uowEniX819maGW0n/sLqf6HUDlekcCjO1pVGBIVpFsf2Z4Ql
DZ497b7/bOp8c3wIegq6ZXmcRK87+M92WsECFt2Ei9LOJvIXUGuFLWxHFSP54jp0
qUPDSibfHa788FvQMCRN2xsbVQWBWsgyriAto2kiaWxkdTmQy+L3OBsk5t4U4uWj
mxP82/0L9b0zbEG5Dt1Nn0x8jf26DvZjeYrr0b/3HespjyYT9/0b02mARXMbPSSg
M8U5TeFstRlXnYUcwzXp3QodYswwFDn7JfppVdrFNnPDUcMoTYJ9ooeoPgDazZYv
24og3rZqhj4bH1ZUfpwrs6jYmbwkWm1Mt0Vfl9nLmo1h5ys5341aYKVlosCrQlId
r+O306JUQMFveabJCMZJprBqOLIpsn5USwm6ISGtgizT4nEclrtapqZTWTuh8hoF
KMzoqda0OE/rNWhXMQfFUz6lFiu6aApTNpOhfSyNcKpYrpAbQLAsu+wkovgDj0mI
9DF0U7K2yfW11T+Pu1E7AzuAmF6b/fDEW89U39kgFSRqhZgRgoK/zNS/bn2efMBC
dXF4VzUk6tlWKOmLL8TEbY65Nt47jYcNoUb7aEvNjYnAmnsd96Pz0CG0EIl06JpH
4c/HAaSNyjqSpNPvW6lM1O16DF/Q4BIgclZEQe7vszCW1DqvIpjwsZMhYu614wA8
q+82ybqbuNokO3r1l6MaacXr7mCP7qFrczyh1B0JCbsrGjQQXaBmsbBysu7Lo7YB
+di/+fyTLsIb/xPT9IUenXrDOI/qaU7yLyoo3GkWNaUrzMubaGL9Hlu7d7+aWtPs
knfyCMuJavkZoLxRGqekrXyf/EDKG9axdqGViSlqiRo9J1YAvVs05Tgqy7bKEbtk
E/5x3eW2JDzKu0znonLurSe3x6b2NhHiZw9fJwHniBkoWkkp9U2rs8o2sS09tAJ9
h0sOCT6+dsqVUKLDBYXcac/cKvVaGLwzsOhVVzzE7QR1sItidBa3YCYHhWAAZM8C
1vxyzMZVkaWhaAVb3oX1iUBBbhxIPQPeuspVCTqWQLwlNZz5KubR1UrDyMFd1i2k
moIHd11hOF8fg1KbySjuail8DKlXgf60PhgdWtrJZKAkbfpLnTSe8UhBGaAa42zk
WfnKPfAkCVBElAZBVlk/uA+10cXw5TEmUMBpkT1G7PBj+xBdHcb+yIWGeXciTWtG
URSEbioEIUV/gU5qrBrpwHtmvAypYTU4OT0yF2AuW5CVClbnzGBwKzfskAEucd+H
LkccNGsjBohMmtT/aOTFczkkXkKjWzb/FHzLpQ9y6peRM0VVozY260mEz4iB8UG4
98vlZVb2jzsyxMNcpEcS4YZgpkv9jauK76w3ag9WbrhfhdXNkWwML4KAScMsXV+/
OX12SqIRDZaXEkNV+ee6Tni71KWzhDlMDmat0+DFQ9gXAPyc88eUGF2O/rfswe+f
ZDdOBDNvATJpwZ+g/9XhK+j4zL2Ee4jqkx/aMts+g6Pwa1NM3mvhG4UIKqkKiv20
415PzW5T5mfnImn1IMZiPhg8G1lsxG12Xtg9OGbVAEhcwFaxGMHwSAeGWIGyHYJh
aa4eXt+fHbHa+UNfH1B+44xgorENdxoCV6GPxzU918QJLCH5qsrstLVOEQP8XPmS
wSeb72bXN7gIWOwBSQuxPDSVjp3r5al6bQu/Jr7zHg7d8gCw+pBn9Mx49QNuxkRo
4YyzdfbCej9fP/gmQoOQBGoRkvYBuz8UPIdJEBA+bM5Dw6s6UgT+/vGUG1203UKe
A4QNf/nuB7Aep9wxZZpm7vkGiUlpItvoil/6qqVbn8vsWkDgIKDXO9UFQczddk8B
6Jy6BJWRXPvjC1o1HGMUwM+95XLseOv8xvOl+VDA3P2MPI3KtBajSTfRMpURbWXq
O88qkRnILqnnt4YvRIUROzWrOqrw4U90alV5wHrex0In11T4cYZGCpV6pI37pmru
jWNUbXGkR+wk904pXh8fpo65+8GuO5JEy3Y7IbN0a4TDyaR2WbgmYrbm4rKngLG3
0hvzYZbW/nNT8ZX9DSMq7LrNierhKRCusZop4SIZtR48NLh8idIU+j61rixIiRRA
Uw33g0LacaRQlaUnG2H7Wtunjn7tBSM8ESeQnBE/USUPRSiFqOgwdY0yW5oJ+8Rg
27AiZAxCR2IZmNzTUUXqWe2cL7DaaFRkhG/Ajg6aB+NkFdWLlT7lDidaPG39yNP/
CvQyhHWpjniwxboVvsdL+rFQ7LYC7LQ/QN6ycXCik12syAQnsClY0J92s5oerWD4
b01EPJEeE5eY+ZKnuws2ZC3wOjCncwLB4XEpDjVIXV/2EIstX98y9XqLPKNHFU+l
SyV5ZdvbFf8NT+EAPwxEcFkOCE/aOVlL0QKS9H1jMsdZKOgv3cdmbxJmrBiV6aJM
kA2Ps+qKg0ZgE7MR1b6dO5JC124wkT/3Rz9GrxUen+ovzmjKOQMCiG7jyAMDBBer
PRWDboM6GZBM7INgf7kKm+3t9xkSvRURgjBx8MfWjg0/X+pwgODm5sPJcVto3bcR
MOMVQPZZTTLCDssDlrMXxo3vBLYwQiCV33zAFxcfm6CD2IsAaxScsuNCJ8sr0qBi
hZjziypm0GbS5YsazPcvecekUoxzGIgbNkBr3ApI+tJllj/Smwxw1kqVI8Y7jvdT
xXw+WOc/dvSaX+ivcOmrGjmiy5VIfuPkmEmcnVhjpguj50y9Fxz4HLxhnlJE5xDc
nBsxVplqO+QTQKxXhH+uGEIKzYZO1KnPd4rcXQqWVXpfYd2mquqoO60ezOcnRs8K
ulkX1/46++HowqhPP3RNstRBz/AgX9SJknD3IzBf8pvc2SFaDaES9kvjNtEupIBZ
UaTTMjdfONxaS6Bt3iNH26hsIpq9qJXgYTeGkfsV994BRwil1ECUwkXg728LMRhk
aceRxuaz9MT2F0d1c9R2CNRDddY4jkaYmlSCcL5ehjQ0LGofx/oJBAUZ3dM9p17L
NHokti8a/QdD8giUsdPQmN7A5DaWSqZVV/pEgPaa5PtYzF+a0MsvH6UbhwWmnsOD
BLHsMCcs4OAA4FfNsicfRRCek79utWgwPeA+VsdCjL5Y9q0I9fLez3vOhTZk4OMi
ySkZSU+WcipDAtQVgh18s4wxCC33gmL2ErQkG7HLcrfdQEdtjm7Yt8ufVgZWpGvM
uLfDar4KoM4jKRDJNOW9vcbC53fdVxt+tkm9qWpayPTlrbEUsGe0MbGGZFmOuEuQ
COxWYw6thOcwCKKJj9q/WLBDnOjcPqpEvlzeODgYbvfib0VJSwxcMby3S9EU+BqE
kTg5LilgI5yfF7GPd/Xh3KZH2SPUr7nhQRENKArNygpT5/MjJaIeY9+31h4JWJXz
4UisP0snk/ddwwZO1Lr91ZgVTpceGkZCRHYWAoFBYQ2zGxz+VH6xEMQwwyB7cOyG
3IJcG5rxX0g1KIvYDm51TL7A7xcSOJYpVMtNeQJWq0ZtGZ1TajAF5wNAwTel2YyN
gUMEoHxAPoYGUMA7kXFZZTmS3kMJ0KTNlb/77TIjXVJV8Y3N0QUuuMFjfFjyFqQJ
yjCNP5Gr6gbEnMUGks7/+muSSSHJyMmNF/q4zk7zLztHfziQ5PwhiqGkytJtX4MW
hHw1Ui6JUHE97HTCPNsyVlYCoDbvK4wDZTWB+CXT/avtYI4ZZvVgwepLRIJAdN/o
4bgUI78kEKoACGql6ngsmuLZPBzNGr6UqeBUJje1Tiv8BUe8bMjVc5AZ2WRibhGm
ihPaIohDCSzqJ5veWu+OvQhr13pqzyorizsOsL2+uH0ZZDTfEdTGv6nBHoz8CNGp
dx0MjOiBusjeeaJdWTlnWD+LS9iMTGSg5SkQrvXYba+OcLbpu5Ybw6IYEnrLUfgm
iJ5KSowvV4Ztz4l9lquZnOPuS4a/+puDH/u/LADR0ShXOHQ06zaIViIzhDc9Ux0U
yxtr+UPBiCyxgfulEdbOCR9W/BIrP4WW1q9CrBBd/PoCryBv+QLBQ6ZNN7JlSXUv
ybS4mewZcQFjwkvmQzexgQgO0iety7Vnu7wHVs6u1cu7akUE7SWu1vY/uSLl5IVb
+s+ZATMihTpPoaFuFcr4HDN5Jtjaq9sFz1XIglm9pqxTY5llUuxMgEirK6lxe+Xw
Tu3RDai23bkGmDI8emMEkoIlA9VHDnL6Kne4/L2+8NKYfYG51k0NhXzwdDnQcWvl
x7pEz5GR6d1CnmH5Fk5ZID+HZdHKscxyK0QYFqyAu2fYM6kfolO5ZTziVuvaMjYd
EVDeHqXMkmmzSmVPs1S61+5XXTpy529DFg2H/QEEUjQXCXF5AGJ91g0iHmq73OxW
bY4SvoF+NEHhdQNfPkf1pv9kzeZolY+0XVpkAt95K5COJmk5FMPMUsKbvax/dgSP
mKwjZZ5O+7O30GOji26hvlOsjHn2uoppn/2LlJmLy9MZZqWu2QNGghATsFaIukAB
9k0+43NLhWHEJVpYf4p/7UY2rys90CuVs6mYC6N3SNbN+2OZAsRdP+qP9K9E9i2w
JyrSwhrkD+N77DGE5PVIilzDogb2BISurfF4Ag/rsEWt2LZRBnF7m7tI1Hyh/+ys
ADOOoRdeUPJRvyjpwO+mL8ycsDAHh5TYuWG0dVTClOdItNvzLE6YUqunIJrXca/8
DE2bAp8yJklrkWn4p7gC1fkZ4kfXlHA6L4KXDRD8ug4gKxXFs0e1Jf+QcFguliXN
Es9ffZibsFhPlNlH+U4yHHMIYz5fzxQJCSgAONlZnpYIknGVPs5ZE1qm8GuVsc0T
RyOlTuZbvGZktq6uCLtQ1snEMx8z9PfCG9iQP9EQIWkbYg1b6/N1/EC8A+m8T+C8
AM1Bmn9wJDe4pVP01pwPCWTXW6PrU2WnPsbCJ1EOXll3JjBXimJJFxXw7X0jQKag
xPl/UFKFVNbPGv+RyYoCFRaNZ+pFlYpKveyWFlXRmtcwpkWiJ9qU8xUy0C7Z7ldi
xhCrU6TesPB4DGRqobcFnLNsLT1bPHRl94YAL9MOAYJnl5387E710PYdbMs7CQQ9
3tEDei+JI4h5iuMZHQqAw+uQQd6r93gndH1JgiuGMFjuBttWt3ZTJfWw34DKcOJn
9HdQD0sxKSVLykplC2nhSoOSUUMv0niyNP3MTZaffu+82WgPO4MkDnzNhIAVIYdH
SXdUOVbKlyJy4TxGiGkyJt2HuzXYOzkXJVvIBbaf1wOeGeIwSj07Y3u6g3deZMck
p/pOUysCZf0rENfnA2I+0ZAmS5bQzd2PTKwM8lyFiYWdtlQ8t4hMXWCIWmhM2QLg
WXqi6zHNH+oot041/jFDBf48k+pfhfXGCPadigNrS3RO+yl2HBSKQvBrklbnOt3S
B+xTcpRgsIWom/uMZm7Q432wv4TikDS89bubHojBmPXRtbNLhMG6dvp0krOH+Cq+
LimGQ5sFNaZOxqS7iN3YDURBItgMN93NZAdT1n2J8voXI7MClPRP+gs8jJrCdiio
Ssi98Y+yOmKfA/nv/D/IgJK0Ef0RHefBAGQYmbWDYuKoWmRDPuqjx3r2guXXocgJ
ub49a21u0tl8l1oJGO8qUm7As+vP7F2XL7XLQK6z9WwKmrsTvzqmjpqdttKjx9PJ
rZP9vpixiB/PjyqKic+4DUqW5n1Leq5I4fnSHonO+atbcO5SNrR0StuzuwYf3xfB
83Qek7pj9uI9wy0yKMGS/ZUWAKWCDgBUyDFzeqAwyHFneKmPMQl1ZNK5jAuw+Bpe
wS5euT08dyR8SaSFMKz+3OHVeHAx+f/bBx1Ec1Nx1Tl4INpqHrTpjCd3ZTLhv/qK
yB87VFsLhkmyAZTkkb8aAkcw8BCXPEi5Yk+6Ot7kk/dArNnZbYHa/LBaGAmDHAn7
QsD+onLHb3hgkQoEKwzSeSKMmCg1s2Zf9RW+Oub/tK8Cw8iwE2f41vPJbSYR7Ob8
WNCBFK0eq46ruCKin0tDJeWZrXYa6os4STwykdMsl0C6o3hqITLZjMi/3hHRhwBQ
x7ycePfI840Tg+Q0eRHbPfh2HM6aOC0vZofZFFx1b6efjRDG0HJs2+piMcsY+0cr
MI2586tbd24Jy0X+pp0rGN535zh57Z4rpmaK+ClvUp3eV3zrBusilnZxakHVLzx7
Wq0sXGmr/q7oaqSjqx9LE+dLVJtxitd/3v8xni/Dnd/7ZzafDUitbjBUuy04bvOs
zibv+jbZVI6wVNDDsJB/7e+JD6IMQHFWx1txLSI+1RpdtC4uEyNpkQI3oU2xGgKC
4Yhm+GmN1yOYRBntKgXwmiOwEX8IOVPEGbLFrasU9V3t3MYKgrQPKGuz+Cj4yLAp
0FMLwQpzVl65ceBdkaeFBmov+PHUprIbWZjiIBzge+O/WQqFHPOt4O1C8VW7+7Cp
g8EivnJQAQ59pyCaUZKVXI+H0pphk7zd88l44dNSDrTkQlSnBgQWbZbU75ns4hwO
TYzEIksoJFZb9x76zpS/6Oryb9bB93goF+PC2Q5DkRIQJjsfrziqVsQpCEGV6JsS
6T+QqjK/MGGb3WH46QPTyWUJosZ1IY3GkkSDDjZpbo9deihTGs6At3UwBe2iiDyS
8TX5DDbcG6pTCmKdjdOdy7FGK9nX/ZP0QnIc6Eq7jO8LmCkPurVHw/yoKwZIwZ7n
08ElDrzk/K3tlCzgXwPmYHbmYzFya29sTpkzksUX9xQzoWZGdzPwsEfT4tFMDbV5
CJqty+3rVsRWVlSFPplff8L0w1euYz7USHdbSDZptQTjl6H/dt5EooTlNYJT0gPp
9o/V5VzUW1Zn11OpmtMYpg6MbHqhJFZ5QKZf1PaDmTXC2zcgcwJw1/bkFohYOmxs
fKh/EHl0arbczQPNYDDQLUk4IfZJi89TsofyQhSzmjrNEdHKhfNWr+ll6FELfY/x
BwES8h3Zns4CAhyORC2QA64XJVqFgyAvHPrJJaNxTrH8kMSJT5uYKlnUHGU2Q+OK
N+VLfDehNC02s99qj240R0rzHBOUM+FSOilPTU889jWtc6k0NpKZwiZScfpczk+h
iFMDbeFCr+3njEvyQOd1nxDjhFGONH7RMNqPysbroa74qiLNilWHnqRVFf/zCWUh
lYGE9723AstQLz6ejvhGb+FniA3Of+0KJ2YwYgIySAYlN8gxWzcb4RXR5IG+iYcd
AUY4u5nOi73TeHJtoAZ/prtlcUBVvGnLFoDg+creJXb3UUOpBZPD4kwGRLsw0pmk
U8GHWBpyKBW4LBEACTCuzCELPW0Ji/VjKRDfjOw6kGhpnUC8JmhWll+oHRQ354ik
9NT1SqUT6b3txxyiyz+KSr9J3scGfqXQzA/LikzakSfC+VQFjTHIoVky7/21hDT5
A91li95XVNVh+2Rvhlyo2FxY0swbtg0FsR3lWTYMCUl7YMSwYPO6NZ6H5kfKpS0O
OeDMX8ImD7osWjPeDB3jwhUGyGH6zXA8wQCc/OHuzY99kYmG+h7XZ4gNpu3Bo6AQ
SWNsPvrb9hUAFbevUtGU9OBfh/8FbckOCXw8FBrjP+5JNzp4ziJ+nR+xEBZCJXhw
ooucxAbD7BGDWYBJVlDRwZQnS398QMIwg0sQgzZnCXI2U7JAII69taOfhaJ7BVUf
gSXbGtWGzSjlCfUwqwD9bI0lYOQ4VlPbcF5QBRxrjS/lNyDjA/HZP8o8wjyR7+L6
q4BVDdIXiKX70q8iKGLdI3humJ3mOrfvPTliSBwfVmSkA8fQq6Rt8TGYzfHWXnuL
pzWmb48IGjjxdJhKIpHlkbbboo5XKviLtkG1teitDBg1ge1spKxxJwtSgQJ17DvI
Dia6UaZOBkSdcn3oNmnKyZHsLaNch/wLmKjlJ4m7lQ7+/J9T/ZDQfeaGzJmbPXhu
Ev46d9lirjbbZlOWcA62dgScX+pyYzlySaIqK278HuV8k4XPTkawKyuvkc26lHsu
+pzZVavD89KW8zfMHePCkp2LqWW9fDivjXWWEKUW57p8i9eDDuPUP5fvEf074OA5
MfW5Jz6Qudoyj5zuWdBsvMKndDXGuXz2BIWSQpqor/o6xwzMPsW9i4xqirHIsE+X
GOupD9HY+tTh2E7G28hyDlgbGPD5rjvaYGYBLsp3f257McM3kulbFBX23imDd1Ce
vDHixat+8i1Lozyx4A5uZh/Xx4qntIlQ0Itkn4ey2Irx3+DPFT6VYJsmq2YzqC9c
EQ/BIoUItONYbK9cdZ38lTs5NxZATskuehYWlEKDjx6StasDvWwrcQJmfj5pWLkI
5a1zFSAp7qVfyAY/goPxklsIcsp7JD0u2V3VGHyTYA4/KnLAwR7b/NrZ04Sdp8kc
Rb6YJ8plMUIHmDKyWgXFveDlvEp/wagXyU2hWosL/kb8RceaGSzMRDCCZffRPvft
AVK0kI/znIxVi6VgCxGHx212XQbaL7+a/QIqbeaaW+mOOLqFxFpBLzimuPD4ophF
hBkUfeUBQkJJ2MrXjw0HiBFdif+XY6fPDqa2FHYJ6FEwObKciZrTVOxhfbNCUs9G
/Fn6Bej21X2JFtvhzJ1xOySJVszRkXYU9sKJ13o+ZYSOiiASsZ7KCRJiuikwyZkN
u9/1QeFIexQ7uu95goPsLFMQnLSjT6EY/3d7j0VHTCiN0Jsk2WTp3bkD3VEo1WE2
+JZJloI4i5Jeqzx8Ka/bDWNvIiPlVt+l2z9ksXjorvlYex99XzFKdtgSnPTmQ+q4
KlKKq9CzpGlY1iGbn0hU81WFRVGjAU9joS9bgtX+xCoisq6UOJHFm4duFYLhqzeL
jzgkiJ0F7BKhMdlYUX21NITs4yUzEaYxp4JUK7Bfn2yViGJzarxq8MwN7smd+UL9
O8Kl1AUELX4BvccRojqa5XFE5KlYyg14qhRvtLQ1rsoY3nraGxJn3utuUWWXYzpx
0sEsBsULQRM+PjLvTARJvxxHI+Ddx4LESS0fsRxXmq9bd/y4TOVAdr4l4sWiGAu9
PxzTlVSXm7NlwapIHqZLGEWHucZmpM6VkRPPhM98DHXwBgy9sPhEiSL4vSGNmCaD
GFr5ia6mr5J+zLInSwLM0+H/d76fC16cP75xiV9PReJVSzwPQG+7WCgpQvGTStwG
EJtk6peuYu2cUsAhA9CkIURGMqbVS5HXAadwOaqP6btQQeks6cXOU7b1Gq9wm5dc
qSIoa3FA3txoVQh08CUxFjZ6+dnN4TYzfZBG2BcUXGLlHZDg2WjmjPD7so2mdhz+
9T2IPIshyn28ipeK3LYU7fIQ3++pzbstzs4u4N/Xd6s7KNVpeZ/fulaummUapT4w
CG9cLLSQlMi3Cz+YLf9HcY24SFVxQl3jaqI6zraYh6DrlokAwjYdhD3RdkcOxu9t
D89TgB4Jx6bGMT+/4VV9LobQwHx9Mg06htNyUQdV2tDeggCRY3w5Fj2tgc2C92Om
qF8wZlTJ8Bgc9cnCx4T++jqjzZAfyYZu3LQjMJZmxwxv00bVgk39YM9YkRf1WtYK
DafIvDhwIz7JiqmhtMqNPgjDJuv1PkA3qe4c33HySo4t8knHjRn2tlWVDU5Yy36r
N7s1ylxLvdDtie/HJQBeHLKWrz1BDIqnEqpXj34NTUAPoIpwSViiKqj7RUDY/IdG
jfrlHglMyIr3GOys1plOWF+HFKQ/2pfDFr0QOj6dAo7oZcCfJrPHlUcaSOBXa2Fb
QANXa+G8hzCQsK4luYrS+x/AnWVG8bfVKBl5Ig1ePtAxsrAvkBZ9mCkm0PQzXKLv
aI5P9OEjLzZvq3X3aZloJgSGVYz6bNH0TswzpmdLP0pFmtRy3HRifY8drLOUZEMQ
+qcY99k6fFNvHqVs/KO4YGLeS30D+sDtwtkPqiCC0j3F0C8U1VC+i/ZbF/b2NIr2
lXfRJjmDvL32DnCNBonve4Vuq6x7gbY5BHn74gO1o4V/QWEs3bPJsqGB6b6cBbza
c6LtmG9m9jsljyEjN+IFdwojMzRvTPIooYUy0uqi3dLaHUGvXj6t+EcWzTUX1RAZ
jxJIRoVRSW5TijU9x4MdVoHqQXgAa6EQvR0YisJGbV3VvIyckVrhsCbr02fJEXMv
IutnVfhEMrP+z5N0x5weY82ThDo4L4gUcAV1e9R4esV3PQohDJIZeOjDssjpj8Lj
HzQ0xwNVOSaDNzaJWauH0tapgD3AzNrJmgqjE7rKqxmKlHPsZ5h6UIod8C/aJtNq
o4tdnobhPQEz6hF3Eb9awEGJPxrZQRTRlOmKdBceC4huF8lBiZ02vNcC3+9SPVJG
mW4jIcuEdQQ8a9jEyx9tHFXwOHp6tcjNejFmHn314bE+MuR4ZQ9JgHeqSxcaaBU0
utOIwsWN1qBeBaUU+b0x2PVObtIG9SX/BNegOYvzyvCXQKICs4NZA/IieL5rBztK
bLdCOGTF1DCHNN3e4Aup6bYYB1WbV8Gk7TZ+KzMhJpCJbt13+638wFqk8YQtyV88
VyG+94mLWVi1y/sORIV5zPNGlwCLHbsZ022v1EZ+DnCmPs7YONwhVww9dixd7qmE
1sUeS8wzHS47naG8GdHiPCiQib3uYkMPGEmVYt76rrQo3J7sPsMy3de62flggKSI
ZW9j483BqMzTf/GcHgapT30Xtd/jRwaIDJ5u87+xE6NIA3KyCyfLjgZLSddoPZhj
lGsxoIEEiBdoua78XHl5IsSk1C/UQsLckZhZwaX0EtzJGq7Hf7aJGoB9wICLUjWy
RI90Vy1kdsoX+bcgMR364d5fG1wfu4D/6lNztKPgZGiR3bIy+f2raymHm5+INU0U
qMMMnW25ggRuDnYkXgLyngw0RMVokkvDZnOfBpyHRvrUaE0peRlPaJGTjwwJ+8sP
36MNiWRcfRTMd0E/JiEIgXyPazTCYimLpl5NWJFNjPml43co4o+IosuUljmp0wVA
l2YyGxzzU/Jd2yrvxHX6P32tlv4CwgTvYST9MDAmsa8igOaEqMfY19fQdvK8jrHb
ysEvgOkwhspjE5UShhOSk6knCRuzEZ8coJQ7d+2206avj0eMGy8gtDWCD8n6eEnQ
xQcoVY5GdijegGcovFkfHKPJuPgKzdQD8nsfkdCXPL6Nkb9q5kou709GkVjVgQhP
WkU8wgM5GU6oF4kyNX5b609v37Z1yFnsxhsuML6FE5xCRbeMC+9bw3vOViuOQ5rN
poKOj5xHBOLzCHrcFLWeMwqxle6WE5bmG/fXB1c8I91L2rxySHjN98MIjtczZibJ
5+7Rk8iMZm43/f8bQqUwbA2BJpuIw0gYxpikTs3TbE9jesPTRe/ip5y2W2+Z1gJN
fXwp6YbWbAdBYYUm0Dw9fE+NxDEDn2EnbU7ZjG/gkozYtW4shaRza1pls9UNSYd0
Jpm+/WNhRSunlAAfQSrn+Wp8JQdQCpuoQG9ec30z4dTHs89vBy3/VPie3yuJVLL+
rrF9eUq48JXdv3ASKGrNraGgpgiRi/2zNFyvoR7oAuz8BBEh+FoX4KVJod1ufzir
QJ5rRPRKqSA2XHHHJMPFQo3weKts0zKleccaqxAsz7hGBOtebH9klX/368gai0tz
up48NIg9/50vQVMX7txsjhZctk9leQvSWBdf81nX+o1i07tE/S5I2WArxLTQIjGK
vydZH/NH70znexG5Sp+qgmb2Et4Y/zafTOCBlm/lvqMTa5R3ZlBzmDlXNdzjw7Dw
jviB+Mm/cGU4RTGVrPJJ4gL4itfK2YuHlmJjpNMpry3uA9x8kDRkhcBC49a+5h8u
hewAzdH4RVX4gCAinZAcvrE9uVyLtXkvXy4+Ijyj2ZEphGRrLzfCG8DabbE89HWP
m2R1iNmZUseAyN6Q2TyBDTvqUKeWP9ISNoXgk+1JjZsQk/WTfGW4JqmxT27lT94e
EPxJoG8FbWVt+u4QLuubcwCPBuAAnf81tG+YA6cu42MPEipdH6HQ4yR5qZK1hyIg
wRJt56px23Quql8hEFnMZrYphKMbmI9EZj588tJlRq6mpEujaAYe0MDxyshdXUra
9YP2bAGKRcd8Yy/7KN8djtfu0bEsJBfBS1lQY2r4KLuRg6SY/J1hzdbCrs9cGyPo
ed069vgNpc8E71UmdgBIZEP/u5FDQg4BSbkyqL9kQ4NBPgveB55TaJ3Ulh6nKG7Z
uTb0Rl8frIw3I0KVLOALNXMDGnxKSjAuaeZy6mt2fCU3cHC7FXk5Ehf+fEnRsSTU
2M0uM/l0uDX4Ryaj5wujvKxRs9ECNIeuKYw/aHBvKgk+KZEIEal1blI9v3Z5uRAM
/zmK/92TtFfYd4TFqA1fUeHq7xQCsVgHFFalwwS2tZUa9CAGbpZfd8GWNYwINbmL
3DWIAC+lxOdOEPSO+SxWhE1UBugxUmBsWv+Uup+xmR/Vo9lCueulDihykLl/CIhr
a+oy9nvMpwXHcrBHG4TG8L7vwsFLcrzw8UkyZPkG/Tiz50RKbSoNxnmYaW19P+M7
ELJ9DyJrnfwdTm5a+AUf3K9xM3S8Ovl/X3ybgJFVZWK/B6b/2fdSoe9oPCXGCckY
HYBW5+i8RH7iE2m4JrsAzyDuSavXygEpGEjNFGwnYSJeEqr7eLYm0Pg6jRkV7Uq5
2//dmG7NYlu4UjEYEa88XTjThNviKSvyKU7S/XZhLrFC5GZfjvHdDppFQ/fPGY0+
dSEhnRphyzna2uwdy03vh9inFswrpplPO68NRmZJ9Kan68OIZscB4IjvSlKuGBnb
K8UTZuxGXC7+JqZcICj5HgM9gsed0z/43O0b/y9uUU6UAec65qn/zCjNnTbxsAFl
4WPQuXWO+Od+ZzkDcucFLKvtoDGFlacj/5AdNO0ZUtFkDSY/Pm5irguGvKX748oR
QP68s6jkqNB4nCeO8KBL1rcdr+kEUOekuGB/vr1A/yfgVFzbFGP/SYCKdcqxLn0s
XAR2gt6RlYr1Wsi4iLwjz9zlckdfn5mHnNwCoPC2FLsciXkKBs4FuvAtuSd/1r1k
YozBLWpQ4v+7807+soYA2INzgutfzCyjDrRjhGyfdfjaW9veOCDTqvqzViv8ZYAt
AWUDZTlDcLYV9cBWBhrUZNe6Lx3AZ0CisVzIW/hj0icydAyvn9qO01Kwj1o1WulM
3mI9pIDgdOrxxdcpW9xU5B+VklCCLISTad2C/X+JpiWteOTRXqcGFoPotKAM3Od2
NHB1fEFbZ+Yp9crZArfBv8E48CaP4wN5QRl5ZbocN0PRzzSa53Oi85syS0u3L1Zh
Vi5LoIiT8f7/JHxQRTKlR1XG59Va1gstgFm/eheA5aqXN1ZMLNQDyiyZTBmutqLh
Rr0mGAvENmLfgVHV7nDIaXcvZ1K5BVDOokFCcxzdhN0ucv8LvvRKzp3KdFxK/bRK
lQLQOsrEFgDbT4PjeJ1vPH0OYTBkVwfEqd9vmMnm7lvUzKf47Rm+gQgzWIFCw4br
F1a8ioDU1rPYL1sGPJjyBAunD/b0cJAFrVKpi4fkj8THFxpDUWkdEkUmdXLZ4Psp
U4/9hkvgm6oMv5oui83T3deGHnct3t5nO9BBucBQysb+AMA8UUOjgKw992TNxjlE
4J+gjmtkSLijs6AbOk0sjh7CMNA/+/Old96eRxXECRvkIVX2tatj1n3O2DymTb+V
jHHGqpcBPP3h7ABlVEbQc7LdvdMWwcIWDlEEM4hn3uONvGFJhRbe6KrrRyPqvXpJ
afjUkpayCFIpyPjIQX6IRm79+uTX9+BejkbZ7iMWk8LAQ3tLTYz2gefTctzVZXAg
yzJ2Httf1+C3Pzmt1iRjTf5tKl+xaKsl7YrgfYaTdeUOWs+nV0FRe6pvKBLV7XNf
KLj2rdJrzL1YBqrw9yp0G+HLmsYqLYhaED8eLtf6TDtOwvEI/7LGuKzUUuHKigm9
AtEd8pfw7LDkuTw3hlL7XsuQlKUFtIAUQwZ1UCKaeI1RPXX5Xk8nAXj/UbtEC96G
UPnc526h0VthIqhDh7WOZmupWDQyAjPl+qOXdtLjNxpFPJVVjHRkj9IGCRl3K/8F
lCcmYb/C99VkkU3EApStGcyPYlFFoYIrqOJq4fywv6gtpTDMbkoj5LQaoH7nqgYl
sJQzodgRGr/0gMtx4y5o4JgveE6u5W2+RTz5Cuj8ZNYNRnbPm4R6AFO9VP8A+teT
CoMllQ3PGYYuygFKb4p8iQUtMTCwOckFvAftH94w3fY9eXCboEWkvtdL8jHtvcG2
czvkpd22XCTbAkb0nEP4kALPsV7O9kA2qtZyEgu3dIvplMEgAIWDYZ81YxcFVbrm
jOcEWGPbLvipZK2Rnz6fE9ciQ5IErh+F0qWi7R5ATEqNYLaJY6cFU0F3WLIz13Le
OkJsiwx3MerIaCt6/2Jmn9XHxn7OxHtlICMcfYJwRo3LcPcOtRttq/ch/iSM7/d1
+j/FqV2i6yKjelZcPSnfmozsvLvQhVmt/ZlHPoQV1hl6qYN+2lMtjrRsuJybvwE8
BtQy8l2KZo7TdSDVYpZNqhJj4v7m6sAVCHJ/1HkWu1pdIkepk18ETNrwoFn5JIKp
OiRtKmPJ84cZ4gyXj1oN6flK+5Q8Bdenw2S3aukbdo2BSsd8uia0wwh7SQGdtWeY
D/8+A/iF4LcK+2d7imKRAScoLpYFV66QkZmnHM5m9CfR+CilLn9/KZzvXCyW6zx3
o5bUORC9tb9gEs1pZqUYsszC5XEXhIQe+wwzKRiKCr/vJ44o9JHtn9UhPsRAD71o
j62+i8OJ9lWSVEHMqhU340JTPRVpZHqE3e3x+HKZBp2Gh5LwKaQllXhmmxKz84HA
CjqUk5lVRye4o2cr4ebafn83v/c1QtTAoYoTcnXcN/sPQNoH34SUDYPb8aNoN8YU
o1p1EISGXb46PjIsTm5l7rblEOwOPj+1YDwfgtZGrby9h5aF/4U+caCDcuFrhqNm
3KqJWM3cE+YP67nSRzdsYpFXvw85XRSQvIBpAl1On4C/677tDFmQhA6+ej3OP7V6
XsM4R5e97Iky2fkEioyEkpEtd1k6ag80BD2mvX3BqFnl42ThBg82bXP53ZQSXf9H
bfiyc/JEzBGXIBgKccWc0Si0/+USkXEwZdYRtFm2qpQBjl84U1ExaA23ex2hVtnR
IIf2w65KOk1oOkWrnsTEvjZyEefaxjtj6hm1X34LmSb3PqCJuDx7M+1HZixARd8c
J5PO7OpzruX4pgr6SH1AGL0cicPb5/hSTvou9En2nBfCSz0ZVl7eodcV0C7kTseQ
U0sazljSYbmF7JtqPRfg8eKmfPt5xJhD3aG1aKjLG4NIgiQenG0LgYHHTWDhD+3+
/FsihZhxJuurimtEPFBY1PJdK15X+cIwgycP/xFFJQYkoerEPHDlgVG8KiwnerPg
EKifycdbdbQ2mXO832a+8REZnk7WqiXBR6IG54EAKgm4rMVdar1YpVrN/HtspMGu
0dSNztsAezMQUlq4BDs2QXuZSwKEvEnVSkC1KMl8sc9E4G3omoZTfP+fkm8msgtT
aLbAIy+ABrfLbVNbqe9XVFnGIthn8arbepJpPp9Uz9Tz4Hd20R+6QtbnCaHA3C/u
A7+vT22xkR5tsAm0GHwW43PQ+1Gs6fdEHCTlHhWIYSdzt+wuSOhVxdriGSTMHdhh
X5KazvlhPKDKuUGr8rdJPK1th60X349kI6JpY/rwKsLsh0NWE4Z4ZBTXLYjJMdnZ
sgyQwmQGb7VY8SxujNMpJK8UJkyeVVMTIZs5sn9EbRidkXMxwFM3w2xIwVzh+wzv
mdknKAIc+yFa7msISs+HUyx9ljSn68P3ySLL8Jt8V3+txzJWi3sRkwsbXXnK9DR3
wnUxkuzsi7eDWla62ud77/u0Er7VkpN1juvKpwspiyI4SlFt3MIIb5/OPrGc0NqK
qX87MyJr7F/rpRYBuXMyM7ob/hR3tYnGf55z/RvcvVSjRJ6wgBqYkYLMXsoY/Moa
gCYI0g9U6UwmWNtITua9wDACWkyq0iNe1Ucs0KE6w7853BnviI+pygw7iFS2VABZ
0dUKmjGjHpXytYSLzbgBeSUwf8LchJSffaap+WNkYT4XWqSgWzvGQQ0zsfTbUiAt
Cku79xTltfv8/WD7WTT2quN2LvZ/on6uxTziOY73R+PDAvlLFZfSnv3mk/axEfYG
lrQs5klT8XYscdqr67IThWafR11EOfQjbpHUwgMJexP443M3BXxFima1fbrkNI9N
xOBiSACEghkjYX4kE7Ng35UwjnPe96SP1kgnwCwsbSbfopLSja33rR6tbpHhkePq
vu0zIca9AUnF92KvkJ0fNr/jP3PesFEaaC7vbTel2Xje9QsnNada2AJLUBS0SxOx
P8BQZW2Ms8VHx81gvwoXMEW5y+kw5tmlpQaZVOnkNpPt1U7utLGjNX+ruEKuSidB
O19oUeeeQkkF+cOseIW3+icEQNaTdMRwp6THmyhqz4GxUMcwtfBMWL3XwGV84m15
9XreZV9K7MOJL6z/B8sI8iyqrBYOqlGdpd+/viV7tYXmRZ3lLLZ6YaubKpgSznxY
DF3B2ZNmCphh+woiH0YxYH8P113G2EotCDIG0D6a5w7AzVRMXP9pzSlHorP1rKo0
4IofFHuWIGgH4Bw67TfxLHpBlL1qAh767xWmiyx0TMp+coYSXdc5Cvs7YDdBUNzH
rgnPMlAeoUwgCu2GB4GPxzfrxRpU/Q73YtyUdwb0lWp5KuoFhkLpSPCAK0rxKQI6
7om9CBZw0lW8giuYXKJ95O15BFL2oo8oBEUpigmEMJCQ/EiiCKx3yPWnFWYwHkKw
GGbxClQB9eBZZQcBpeazUt6cz3yJmNq0Ehw7RirAlwy8SkGYlxKanjpMdJCb6aO4
lnK6MqDIGUo3m/1JYd8ljvLnGcrIXYzhqJzhNQ09us4o9P+6ql0+0jo4qEoeR/l/
78neZ1JMXjx0vVs/lSgdMnK/n2njZ4YvlG0iABquzrK0lgtfM9OvuLqZXxi7Bkrc
Of4Zy8BN/paN1J7n2XN/j0PGbPdw+sIdj9c65WbXHaZOFWLtw8Knvrh1FCpeimjR
RKGuScxN2bDbgqM3KKrpzkt7iMwUVQU3gUUsNTgynaf5IE2E27/+XgfBVTOcV66o
o5lbL4uqrEyD520QM7jHied8K30t5hvre92jec3Bhd2aLAmDwEBfjKTrdmr+fupM
AQFgLV6R5ByQoVjdIZW4e2tiW+uK5cED5lanpC17frFFQhZu/J1YrS9OtjuLq/jr
JPzG1my3hLbGm/TQ+jAIF4XA0PKyhM1ect8e9R1jFgYVrs56lEcmptZK98fPG1M/
romHP9/k5nRvUAvYj9HtXK0gqU4PPRqAa0ROrpysKa+E1QFxpkhdlHAe20OFz0Ut
VNUiEVJwmXgB7kILtrIJ1TdyLk8M2sL2CnoopWKSop5QAwr/yrHuUd96lTitW1sF
5cML3THGxtFTr9rQRVKYcUQq3Y6Uh4kZDkt1lkHQ6G0BzxoyRkBgwAhPM5ALZ5X1
eeJGjggxtFPSv7mmd5xD6d9XrtPG5ZZ4zvLCP3l6ifaCv3tDe8wMNqbnkF2kPcl1
Tp1h2rmr0fRBwizg3qb3P+oBakcm5k3odQ3kcdU2xKiei0TBBSh6e63tNbbx5lwx
Z13JQ0u5cvgi0zR8joWlLoZBGRTreybQoENLhwZPaJS7nO3y1ORqdj/lIWVjSA/H
Yia2ITaiQmzG7hqiu2Xj7SV4J5J7a7Tp91zThGsE6To1Gx6UJErzRc2k4BO7il9M
cpGQ3IOfQZt/7BEGHzDoqP/ZIf+oYSJEtCLNLXAncsrPANh+35VH5oqYy61JDB6c
wETNU7PYl4mFCMS8gxYk65xrXcOYKdrEAnLjv+FkRKe9DwJXfbUngYIuOZXrhQAM
7tfHbEMG4aYsgZYjziVosHkoLCmvhw0+3GCn+8u2yGzqjWD21gZVyfh0ntUfecdI
xpflc5FTxNy47jOVbZwcxd66adO5giB/5e3HbNy9dtSCECaEsg9+kYHizocNZ45N
ajocuTVKy7U20ztZfg+JMrtg+3fFI25UWos+Ynyi0PXMyZQqMMLVEm76C7Fkovoc
U6hhrSZOaJVv5tewaNXwlM+k+TlvAcTzi/hky2UALEejX/lP4g2sK9bjg4eUwQrJ
jfHVzX43ySyP6x/k3w/emUeNDDNEWzQESgwrdP4v1ZaA5TmtVoiXZmYBRkFDgOl/
8eOCGz8DQl6mdlBoCNuHD5Cn29G0a7+dPrjRrQhRz5B7KCu+ycUaUkXFNcKOE2u5
tjRxaa/Y7daAxgwlLEA1YIi0UPfUnXdtTbX3Bx5ZlKANtBcCxp31WGMgTiQFeWPu
+5Q1cn0npbPJGFta5G1cEAxY6kjvF+pGxUBkZnR6bAHrp64RfsYcrB0uoTN6LmzD
ILaxhjEQ73bDiwas8fRvFfD9S0LYktrogK9kX+MnWXvWC084OhnZQnRrkxh7nVe0
vZDak1EK23q/BtiksQiRw8J+D9tTGy/YqjEzCj22aZCglve9S/8YvEYOKsxtqMBF
L0mqgjGEF09cGxEoGgHSY0l9UngiDcPRMMN5OPznd2rbV++ELTRWmUI5xLFqG1P8
DXd0Yr4rRPy0SQthu1C+QZlA9QshvrMqispf4LgInFtCBxWHfy6vrtmTf2o1aq+f
eQqsSIyGYB8NwXdUdqr6TAONhF5AUpY37y73a33EhXeADlogDvQTwuzhPoETs1pS
NAEWKOvw2VVJWHrr/7HbxJxmed2AERJwzTuWLvrFZ+aZ+mGeDKtxfGFtHG+2BCl7
M9EFmVauHkW05LNkgJBVFE1+sYm5wyRDcFkvt4xQC/bIGRQ7B9Ojzf7HprVG16Tl
OiodeS9HtW5WtoBqDzOK46tym3bkpeRTq/sBAR42vPRNPj4IZgXxkOY3wRLAMwVj
VfoUZ3OU6xmML/aCKW2QC3Jf85gZ5WCmrdPJc3bu5O95d+g/cHBIojR+mmfR7V+e
XotnqlGOUwJxsE6pidD2IXVIoFjrQrUGL0vY4R/bQUfOFQn7K6i0woMQ8TsyWsqC
eeNsHoNrclXeaKJtDksSsdOzuEuVODzwwtQc0ia1Mz18bJKTuH0RTTN8bUQKA/9I
xEC5XQLh0HbQvuq/R7bZggeYFHxSxLo/U0gUelJeY2KBcwtABjgjUILzLquTehcQ
exwxYaauOEtftqFNTYnCEXlpgn8AAgAj8y1aO3J1L/eoLLtWPHRGkayYf6O62nic
KnIE0RhTXsD7M0Ab4nhc+EgDgwoq6g4vWqJ/VAJlqXm4vvae9Tl5UnghGKwqa7bB
uuz8vOq6mEr/UocwWddGrLYIj+wz0REQSAgOMvH2Tdlvt4slD4UNycijeA1uLDd2
Oy0sZ0soCy0FP2g3MRqGgxGxknLnnhSTt7ME6XXPXYThtT5ej0U1eltMbpyvVtA2
Df05xDG9Yb+LUT6PLb+gdTCmwf/I0qkkKLENr8VFCbkro5VsP7UjHCwByjR2pc5N
/FLw6Jb0bSmbUtLpLSw5b/ygPzMXwGfrZ/6ar5P3RSv/NXqpHZhcHfnLvS8mu173
kd8jFcBvAGrSC5NeBOAMqvkvJ4kdoT2ejWaVcKJ9LAWSqYSrILDLaIrny8k1LA8e
qaQjB7s/3qNJZAn0h4okHLEOyq727zmXK46kSoZWJVO+95Oar2amY54F58VY/a/F
KI2qlI8S5pXpo4MMVCWjpOViVJ/C4TOSSN26umqm4Y7N6MlqpGIAw8fbIcwEENTP
5xDslIO7WjgYoUfyATvGqbYIxW7XjCs/AEqcUG7wHiZp0vzJBzcYgPRnN9m6IUg4
Lw/qXM7Nh/0kU9/aAXE1QhwNgd83LlPfko6ul8o20EQtUAyggxmYV3boPdUB1sda
8CdkbWpv51EqxrvvgTje0EN+33+W4MSjB9xiVW+GdjQPs7S375Xj/b72b0C8DZ5d
kimiMViTGZWQdNE7BLBCHkCsPRZl8N9WwyxsmLvdXLRj9/T4uIw5dN0x8xAifYRg
05mck+QW3vc5U23Rj2jX4vtXlT05uamnYrJ0Er18o8LT+pl9nw9vERwl8RBqrmFN
D4iBdrjMkfosnvVjVs63/igHIp3rKtode9i0MhsQmXK0wNTLQANG6lg4qB2k37yg
eVgb0Z3J+z/MHt+t6ujE8igf0+t252E6wrEOSjlZJp1hVUgbdCFA7lw5PUlEj4qI
M7eaQ09IA86LVDfomH1o7vSUNKfD1Uc2sdjmNjf14eIzIAVSQGvSm9GUBbxz+VUu
x9jNV5b1x29nDHJA5Zdj3ze90i+iX3OpMTkcVJHKQ2pNnEc6F6ZiYwh4i9R+r8qw
A9Q+GrSX+iwOKlQMRuSGg2n7UCp/BIcM3KB8ah3sQ5/2CGb4KQ4i20LeGMsr4AOp
a1/LGMD1dvUAvKXBDDN1XM5OR17+nTyv6H+7ZG/em4D9SRvYeP72NWUFKpRo3O8U
CSPvnQozXOkV+lOtsDD8gh9qnoO879O7WJgKd1jKN2C+K83D8xJUJomSGRhf4hg1
bM+Z0/lPWsqUqAXr241YrBowMuf8tXy04CGhluDYGIIO7MHo7j8wX8OD4K6D1bIT
BA35RtQ2dU6ebcs4JWaHZXLXhqdBxxuakf4vnIbLBTuVL2tm9Km5xXJtaDGXNTKy
VsChL4k2uDppHVX7+2tdGShjCiGMvF77FG+vr+ERZzGLjXBxPdn6emVz8OKphXk8
MI6cORvrtLMODWeCNPqmrMboi6GFbaQFcWLsFDvANAU3aL1zKz8trrEpz6FABviu
M6R/nRymIrDn1FGQDRDtgs62TbeMiN6PDDr5+YlrvPUlI97pDa3EvM0Oo2l21T4Y
XWbanQS4KuT1VGYgrl7krgeGzmy4zFtX8/sDBWNrd3ewZEoxq0fKKSO1R5KpTPGC
5kRlS8HCZ9GySlLC5TLXakfunLClvJ9GEWdyWfy3NaiA0xaXhmGeIr30BvcFjaD7
KxB0KsYjMMoJR50M4Hhv4Io07aNzLVLohb76QPtBYkU+wlo4ANiJKgefBYWmTkco
h8VgbYA+5TaOu5wcuqb10PTshnxCI7Gn1I5oyUXB6yELpSVNX2NKDsvCHjQjh/nh
/FcBkGPA6skOFc+kJRflzFlUxXYWHcgIDVwxuhzcYsD6SOWhmnJwEXl3E2Rmx6JL
us/v/h+ZQcQyynGG6s45WkGDSg9hHyArX4GRPUKU9pgd/RoIel7IrtLnUOzUApn0
MPwpxzzIH/WKz988WxlJCwAPz2h9ffynUx16Ldt4n91p6x7ktFhKu8l8u0hiyw/n
I4P4knWKuJG6SrbGLboaWC1fPgy/CZOxsNV41r1FnoJB2e1J6BUz673UBm+OxrnO
+dSiJB04UY9kOUBubc0it17+XxiDF72yIdRoW/o43eO5Bws8/mA0m2FR8FCz3Sex
6TJrOD1x7sDOcpjmKNQfcYyVk6NcBekkMkh0lp7bHc3wfSKtaKIHlZ7VCh/0x2Zw
daEJ97e+LbgUI1NkPs6ZBzoqu9HWycF3EFCV+08AoekJEjk0wrPBb8vYM6YDuaYP
kng7jmEeE0rXx2S8Pv2h+ki11dtm7Ms2DplWtwJSekdPdhlElpo4UhF6YiU8FtND
tX2x7ubGkwG6BKYu3hkzid4TVi9nEew7zJRW/P3/XeHQOyIK7kQxKU65rx2pFLwz
zTRnGeNI5jU08XTVhyvzZMCucXZvT3iTW9NH+tlB9+04WJv0BfXkgBtqI4XlaTa+
2h7EnCGxBryGMuWtatuWW7PEDeJT2BOadGd468jsIHcLfuOQCEMNiF2+WGioDc96
VfoW+XrWN6BJTK2ocYG6pK3V3+K8K7aGakhhVSMebMxiqLqSGtiH5GIC+QNB9hVQ
BWlxJGvaJOZdqYIjAEP0l19XmuzcDWqTmpPbTILJGXs3TzIejKTR1pio+CyjV2VT
Vze2psp0KYTALJyGRcQsgEUGCzNWn6Os3vuSQ3Ystk38I3VEZSgXRunlV0aBy5R1
zyA/WeIHkSvyxbEGNaoX9SfY+mY1INVy1MK5Hv10EgbIt3UqrlIZERyMVKK+pfob
zzncsEJSXFx0HskcQQqZko4AwJ44sU5rKFVPf3pEN/f/PQX+A6TrQKage8QWnDvH
xeN6ro16oaYgPwtzWqPvvg1qgkhLlPFJFcvBnc0pb01OhBqI3ytSUgYTacaMW2Fv
ytBwmwJPHIDoORzxAUfpJQHb53Hg2peoXuamg7MN16AW21oI167d2+gvfx1Vn9ow
G0kRn9gkrHuFbuK+F2jzLJx9yZXQla7ngaTVmSAKzb/+R3oVa7zBbOf0DxXD6CrH
3UZ6iJB902D0+tuHIOvUTiQ9lhgJqpBG2TilzWtNb5fqaHJdDUN9NtfVaYDF2Zrj
pBuVG3Ek3qFEWv+QA94po/Zr06jkJEHCLsw7wWSq0bg3KkDKB32+QJ3uWL9MhQYN
zAbSCFqvVTIn3kIxC6qfEIsX9gvBWB641aU1OvprJP0GMfbZMFsMr6I57aKIQQ9K
7yN4QBmara0gonkAJct2ND2jSKgT5VMQ/jP1qJcDa32pJw57MEu1S5irEW1V1p+r
ay8WGXCYGsn0qF8EX/Ezu4Hq2RfTSgQleOZN8tkOECY83+aTJYuHKNWyPhC9c6Mi
519+MtVei/GdFV7fsmTFPURW3neVbdSDzjeujWGRvoeLeEIKkNWFtlTtlccrjSfg
HW3PWZPY6tnf/X8nvV72SLruCloDEbzDdVx0Qd/QAEysz7hRpcLXpB8NXuAB30YS
JwGkftPS/8m9X/VyNjCfYYjzhYnQ70ib7GCKusMstWTmbJr4tQblo6+LxGGaAs+j
V3kklzq6O42DrIAvFOPiiQ0We/raL9ZviOFvudVjs3IRISdudgDBC0KgLUATBPYI
qZIRBvmlUm68d8i5FY5eENVOHGVnhIgo91S1oo3Qm2FJjd+ut2Kk9N18D2latdho
TYAmbDZt4C4cljTFxBT16pIckdXiV7vfBBVgZamSI0vNdbfeK8XcmtsKG8YqhNcB
XFBPb3rUufSY1t6Q+Axyi7JUPfGq+QbsVEMhXh90iSMAlCFdnMWoH51JXlau4l56
4cHan4xYnVAW16kTt4ZRLXwfKFw50EZQSIXIr9S3KVIEQUdhU5HA55DwdZNaYAXE
0wg8H2KS7MGpyd/AZvN4g0q7FQnm4qt0bJN2IQKnybonaxqWtken+iS/YDVzQ53l
hxoAAzNsriS+xbzSP7K2NgXo/dvbfMI+chNXDaHU+yTOLMjQxuIwpFY+Vdqd5D3b
jk8wZNFfVSdI294CCRGSq2f3mwWVNGxfV7csZhzm2bVMfN0KhnXapZq3isUzmxDO
WkRzlmOogESy+cJI05yuDI6Q2aJ7yN6sRwbgaxBb7nFaMhdT2q8ZWhpRnrjNFGVa
3oHgMldUagK3N+mkQ55oz7ij0jkjUcXYXlR7J2FtiGxTOoA8iZ1COxdGxlEBUjwe
xIUJRUveHSJVDmbB8p6HRTdhlGNqnTOTn8O9rUYOvIp/QoH0majPzAAiqAhhMVGT
VXbDKVqYFxvqoCiftbHhr0VRKL9tCiK+ndm3ZjEUOp/A/lY5sNtQ4C/k9BP0i/Ij
lFv/2MxZSneZ8mZ//kvTy1WTEK9O409X43fdcKNSZ4VkBAdgSoyP1XHXFtt0CVod
ehPG995xC6tGfm1PoiV8kCwvW4aaWIfinxDhELdDPRR+1zehNBK5yvBQ8u2qvNQs
SK9alCaf1dGuS+X87gJiByPwwrFiKhg1sBheMpr4ZYgw3xefMCMfoGZ2e+hO1zlw
QBQS1kak4zGCkyrnyacxzmYnY98S7Fcrt1dwZte9CST7PWP/8PevZe9DkEBwEwQS
+jcPMTT2ybi3xepHFC3HG3Ob4ozkuOR70gB+oIGL1E5ZnVEYFdFr0ZG3svu13M3r
m+peSX4aDkZlSPu+BqtBfjYngLc36r8woGbu3bHoAiPzPgvajThjBFVMl2+Mceqi
Dt+axV5+dLg27XD+F9s1DsFt6hjirCWTn6lpMQ9QiZYEMj1XM8QzwxhWHROJiE8Q
jutkfnMZkOUiABa4Blc8Y1FpwpYzsbll60+0z3mQyOdDSf4uFufudwrCewH2rJdf
M5YKMmo7OCsU6ny7rOr/IxVBKEKfvv4IsGD6VktSDOjwEigX8qtrNwvs+u2CYUzn
L+l6rKuKJ3V0U5Kk0mFAAhKgCjtdSQfVrbnoJGDMhlSaywGUpFgj3cACKYUvpxp/
TaebqHo39MMY2gSR28iphALZqd9zoy/lQZIMvqOCxJP2ykuH0w3ZOLF5t5haWAjW
9Kr5Ycm2Naw9qucYLUJVM6zGESCS5ctuQ8GZvCwgtP8UQ58c5waKk0Hw/hxfa59F
0ohCPLk1RNJyt8hlIfVZc+u16B5EKW+kyGSM8xHhIuu5J5H0kIjShw1pQITUV0wx
LTfBcsdv8jBTDTIrdo4tbu1wxHdWP9RVPrB42kSc0JTNIBLGOeakkbFfqLq6RqEP
VbY2dm3hmWpy6cT1clBU5lDzPvRgwQUUi8yZyBaBZaenII5OWgSnICOxh3mnDx49
z8Gan7ie5ZH7q8jmlxCel4/g83XP6e4rqAjb9SKGMIHFAlAkFd0k4TfZ2Fv7baas
LLfJXAIkb9WKD8c41/HMYa9QHueq4l8M135WoTM4aC6fITQ2aj6MQpbFFzH2bRyF
fkga588Y2aBwYWtXt3SII46KhKcFRLNJ0tSqa9V3PMq0zcZ5+G1REOjqfcj+avQg
r6DGCnCjjxVEOQV2hgbgh8ziO+8xA3sb6eydjafX2UTDUNqoJ4lLrTGEHn39ZEJi
gmYBcGv3yI+b3eyrqdiHjNtZ/c4gitiMDD4w6CXwMP/yMAf+p3hMX82wetSqNpIh
7cSsyoMQHZRVyk3I1CWLguHF5F1/rttKyKRrjxxwilHiMJEz8RjCaeXtdXb5VQgI
0jox7AeotR8yf77U/1fTFDX+66BPvQmiuXCErY1ISCAcTp3wCA1id7QI93uJ37uS
Sb3Lvb0E0smHG5ucagjgWHszs7lboTMTcq+h2C86vcKaFYckK3xvM2fsaCfKeTs7
G41LlKyzlYUHHYMHlON6/7RsVDGzD598deSgkRZzsmzd0Ms6Q88Ig+lT10psI2xt
yBDE84nNZB0BdyMXVVuZwglhnzd3DF3pyOXc5seU4zSSq9/rzqEDh+THAqFonJVn
oHNkTqHiQlcXaYqGpIVYDHuyT6Bvm8Zwq47LkxgkAfr+0sOCB9m6xA2L7b0VcAOL
P008zfIuVQ/fYdo6B+gtRs5LgsDZ5ehCJY9bIPNOr+5fk710FTcraSggkU8kQKKW
9AmVSpiK3a9hJfyRJrOnmUx5Y5zBOJm2vB7qgqmHB34AHDkZivBYsHOPnTHhCtG4
y6f8IEESO966bwwDT4Afv+YS0U8cqyGUPQd6Thn8qr/tg3iFsDD5UWLbzFfNL5qK
y0G5qyQZ6WCec2v11COhaiVkdH+5m2fToZCoY8dmgKMgtLIHGeqP77sJwEufJAr3
U8UNDichSKedPmbTl73Cz0ihxac+OlMmgtxoqTrQqiE2BmSiSKdsS++4goPE+oAZ
hjpWxwdy2/uEn1CMTE/6Vr3Bk8tJkmUmAEftJkWn/URp5YPJ8gKsOv6OJ8ol6e6j
SKL24mLLZvPx7SUdRns5F5Daj+SXCSD7v0rUmri9zGukPEssoZKI9odXHUlvyXO9
0EXfKR1CRmGTl/DT94UHHzHfxwnIP3AMiQQEPXXW/+wRsHACrcKhqFccWMd++Tjr
WLcUlTujyuhlJh20j44RCfpYzX+dgT2sYc1ypc570K1r7bEDc9au7e4zR45kxhr1
2viPo6RpytUD5vYIUJ85hVUjXC2j3aVQzcAfd0YhLIRQBGV03nkZqSDNc5fDwx3b
opJzerDQ85O9hCYVgMlO+YcLwkx1nPrtHpJnfId7K5qnsr6tmEpMC65YM++I2dTQ
4V9NuAHrpDbdy7L290DomfyDBxgU9P2Jk1fUv6dDN5e38ecPef0/aitKz+4FmJvs
SfcLPL9gwwPeQoPOWfABauqhP4+yr22b9HxqvSXIu673RvOo1ys/f0We/WvTWjHq
NiPNxlSXcqhQK2yVSVkwN6gIwxvbIb2OP0pey+iTZ55Q3VhXPN2VqkGkFKndpDCi
cQFDD/d2hm0t+twIqa/Gje+DjKkJt90wF43RM7y4kx8p+YiW+IWvRXkD7wf9kNH6
aN3KwbiWRHLdBimAdWKwn4o10Xfmienm5sg2mVLmuB+KAyMjUxlEw2X/r161w7Te
noABhUn/V683Ufhfo7P0CqJP97oNHZhTYKnE0+AC4tGPkR3qNIceoXAboByBTFOD
fRRyrc5EbjRwi38+I7GWUt9rxVRSPBeCU3tdcIgSPbXGWh3mSeq8OWUadMV72Z2a
5T2s4yZPuhpp4OHXenepYji4oXl0P0uwbjRxURFh7UjtbPRVhKORVtFilezvBmYe
OCzPsTtLJR+KOR3WTkP+9/7AXC4KmmobSBF+j7ACv6X47G8L5p1xcYoljG2qAhjQ
chZSEEvONabSoYGnKEC5eytZhhPLoe/rG9UUwzDiU7mbnCPfuMFYhn9lvpalWLp/
cXYHdVg06k7KuVKfKTu8Ox7lNBMn8N00NbF+TBKW72+1Arfrnx/Lgnlt7iI0/jvU
i9FmJGSH7s182Mrx4OD7j15BJhNN8Hht0HNtjYP+leMZd1Uvx+BGBvmAb99YQR2k
6lxE41J/WNsJZ5Sbhc5nsRFGg8nP4cS7N3K5cWdSwswiepjyOdB+S+AsLtRAzPTP
6j0pfr/k6Fd8z/iTHyaT389etI4eFDsrUcWxcbeF0WL8GV0Rl6ibS3vkPr3z+7x5
o8op2PFcjpmuv2MWodrRlveFH7sKFcT9TbR0vhO5oVpNXAYn/MGp5C81o6MUqmL7
cDqFYFP0hSfidq3743VX9n8TYT/FjYHslssVExiD2l/BL/iRNw8zCTTGd828Gd70
yuwzGYFe+rZX3yaGjJ5u5aClJE/mLxCy43NHx1npghH0aFeO8taa9j8iou3dM5ih
YYUG4uqw2SqmFihGTWwbukNDoOtk4WuPKY8gyeZuMkrThNM25XjYX9Iz3wBu8pPT
qhQMHdzfes/mFyZms0wZpZjWBsdlFUdP4sCyRd++OzieKl2HjM+LF/Lx81fVhPJa
xzULKklYR4jvFacsLxia2I4PLnrRNtOhKMdeglmRgf0LHHN/qK21r9cCNp2PupWg
3S3WNQeTHrLw0sb/DY+16Mpj2oNtzu6s7QZWCpIHM24aNmdi6O+SUNjVjBVVYGpR
QF9VZXE/J2rJsPpGTejhItoY6CQTsSSYk6dcIIuiDbFKUIE768o4hdCviQdPdjgs
C6hpm6MmuVW95psFJyB+10doYBhAktuOPSqNtfw8NpieXoSViQNXlBamsdXxiJS3
/9uT3bXl3VKMQrkxJFpdTfEUE7+bwtXuTWYfhPaniNCbArVJop2AH5c+zajUdPel
wNjOdwvctrvPOWfH9IfP/taMTe10CeGNH2sPGGgNS7P8qww2q3vkvwz0LujYizTW
L3gUiBuJftd6GkHDL11/nWyqkTEj9kDov3/cppKFvTNyJ6btWzi/n+X6fOfUr8dI
OEucICpQ05jlSjke6AVUiBO3Dwt2IxK23pqfBAd4TQ8dOgL4kL5CvsVicSRP904e
QHmkEdH/yudwB3EFo8pTwtIVFX+Y4iKh2qycvOHQJWN0Jhi/v+pIO1zqs/xO6ZW5
kbFGPdzv07LgzFFel0xvytETaDwyzPRvhRr9Hm0FVwYepgeoGDMvvCagpwa1hBby
2xOttfsDIUquzmthy237iDCSzQhbUaxMwGECNQvAvvecUcEps847p9o1XTOsJE4y
UdXgQ7mBf8UlEyVyhIkwqKp20jF9ylg6aQAwPAsuVcAKl+oD00bH48QZ5PIkOtIP
9djJCt/aYFM7R3sD5VQwPa1PHpSZONv34huEWb/zh5HVMLWgXeNnhcbFvItRkun0
/Y/mSLMpPB90Lw5zEChUG7VC/eYhJ1In41c2o/pD8tnHWJtYRgHg5YTc/biPshHc
Vod2Zg6iE9u9MapiyXWKD5BwRucatN2EJCGlvloWuFoNqqQFUWAMtf+8yeWN9zkD
xoq0zqcJr2mb8pE9515rVOQeu4ZI7Qh+f1eDK2h9M8UsHSk1lEHwqony7+zQeNkr
VuuKjpwF+KNuHKw7OPlloAMNER+fqXvHoAKQb4yHFYeeHHi0CfH9Ps6BA00ANCCN
av4dvQzQe1ZtEvUs9JcWATCQD0JJKThdpQQdRbn9G3H6moyQl677GSFSifrDaI2w
aycYpVygB7N/tDsAgkLcagxMTzLDhVLafkFjBCwtrrpYQjd51xyrvMsvFTOHzIg3
ptT2MBywVkga0yyqI04gM2A2gYD5O3s59LIH+Y6oOaZrdgcoXEjCspWzqZEVrZ7K
89uS98Ps0xeAq4phJex6Tq2r3Cyo3A+CRlvhZCSm5qZsScw7u5Y3BIQNhW8ZGk4W
mGXxYV0UwB9ebZQuimWgrI1HsWPbf1QFz0u1PzwusHURNzFs1PDtv/GYTRD9b4mN
ME9izA24Da7ct1Ir4+VPCQgi+ZWt4P/7OxT+YhPQ2t0e73Hv1ikkSNHknPy7KU8E
qbvSReK/4xOI0meH25AOP2k4N5wXK/+RYNQbpZ2TNq+BDP3ywTSkEXwJREw/knSU
z/Vz10OM42iwlSY5o/qV3I9mT2r89IkCAbQWDRiK1+ozFlybSwQX1bJgRhGKlxAH
d6L5DDo+ZATrtNkFTzlQN0+sOOZprrpTC31FA1tUaqkNuvR/OLrPlngDsAIS0l29
6G64sOdyNa5eVmkKmmKzu2sIKp3u5IybLpgK7yDCOmdnIIux4svA4m0hUcLd6iXk
D4t+zPTLfqu/n/AwlYfkHn/Xwr4D/84+Ox8uXDaMFXXlGv4GFcl1NISzt061MMOM
MsTc8jfYuKbwzNZf35vnz/lql6yfzoL07ANvYX8c3axYnFld9fTpQxe9e0i5a8qx
QrlsRntc4rLtKzm5C5msM4USai1+mU7pzRFGM4pWBTl2Vc5nFQyXiOvIbJFYGIrZ
WHI1BIOcVqiK9PrZj0S3DONlUYeCk49vSFlrI64b75sIyfAMNGtD9xgEzgmDMPn0
3EMd3svpgwdC2VqEALRIZVfgMLX2D9vuQqU+Sp7EtnGgCgPOgnIq0eb29DpPfrD7
rPAFrcUe/xfqo3UIY1uNbgEypIcjVwWuLY6ULZORtvN15R+hP1YvhuEwhOqDdbHf
mxtITVJbSvBOosGtspkrpdg+X54Yw8OGZjy9hUo3gHIdY9aPn7LGCxpw9c1Lp2JL
y2RWvUhehoDqDxnmYuJWHMnJyFl9Umw0PeJIiS7+EZOTCk8nBzGuCWJdHRgMsmb+
s7F/8llB7C0sf1Xq5bU8Ymtc1KhixY1KstjEbr4NvAQWDWPV/lbt75pwW4TZSS5j
m+GfqbzhD9vEbyfPp4nZeDCVRNn3PjAHYa3OqKSasLuGDpnp69Av4g/cl0qhZjzi
Ik6D21SaeeeJKQNx2lqe2NudCcamJV9Afm1r5wqNhKhk9XEGFhb7I5cR+kVxMZq/
iWstfcoJ0p3pPsgaqtibpx2pjTq+8lwzg/vXDsTHoa1yMGWJ1e9+mgrnosQ4sHur
RKZVbiD5BhrlCd8gYIMKmR5lVu+8KE/92lHIj9pH6gGNmkkTdtmbG1OFxxHr19Oi
TVFBsbhTD/l7n0XO0HEO3Xw8s5KUqhnQ5svQBUCz79KITN6NLNT7yPRybi+XKegj
wP628R3a0Aj4Ya6Jt8q0/kwvC6S0FMPjtKVKkzeR+DHr0aQA4+RwDb+QwVUyiLX+
pSmuymCnHDjW9gA26Wvkxe02MLBaCJqcudkUlK46PJSAXfDUDI2UmFE9bdRXSNSM
nh6wWLocuJF+9tfB0ObCBK0DwFummvOgb0h1s2X329PLAjcgjv8h58XdoTdUOpHH
KuWrYw0oXkQsdzjhaByHzCpCiSN7TpOxOnvpNuZ2m9y3kmYxU6K73a8bqph0aE9q
d12H6sRnO9t5B+43TO+BpY2M0l51gt78FOjAuAvQtfvUUU44UWOefP0XS79M4A3M
LoRyAjlHJN04J6TpqYskE9pnEhNf/Cy5bWNF0qPdcx3sSFauCZPzMXh47ZqkzI6S
o5RcYFiG2/GwHYk9stUsjuBsro+zhiAVL/W5oSMH65TlaqZ5pVAtKL4ZxhlvB2Da
1eYDXg4NkwXUALdu2pwAA7T8Os8BhJpDCrzBbiq5ASkwCMjhRglJ4El+ga+5Jhki
k5k9+g8p/OWTYY94Thy4vDnwBXuSnQavqcnKLnt8H+jm1XrQy4Kv+mdofdWFypv7
eyff6n+nORavJ7ZbwWUF3dIw5aALatiW79BDnCdq+7MbX7Ifq9cchLeAP1cC09rW
uy6M//UNYMrPdLTjfcBPG+ruTkbumCqEl6x9dvQ8neu8U9lqz6qnzv4dF3r2Reig
ZJyyOdcPeqBFBIR4HPAo/Oe87hktIJe6YtlQX5dNuVqKxb5zgKqn4t4TMicf69TR
WbBQ5IJY4PYtQUmQjwCYbdgFETsWd09VdF4jcYKUTR1aK5pn0JRIhF3rmRE0ACFi
+diBCMpgkByceraWTCMaQlbKvLPd+NmXkEQX/lNoOtLElnbMyA6nBYNvhwvPRVzO
rfupilgkDk8DIcjc+YptN7JUCxY3kr2x3HDFfcZPh5Zict1GYvDLkMLMAPbAQV0g
u+dkpvVBcwwPK+bZiXZMudLfWppH2yAzV59smbcLROgk+2Zd/XX/xFlXQd6PCWFu
w8sUHV/IVyqCWYwQYmrG+sfljldteQTf1vm+X11iqvfieXWpSDGRiOPn8guw5Ruj
PYQPaSvo+9XlMeZqCl5SAi3HO0UikAZNcooTR912wIAGd0UK7TrkTtWh2HpmMGGh
SfgYvGL4Yehe77ONDnla9KiVsYDoLk6FqU06r2MWU6tNgWjnckuimAWU4UPAA9fI
KMZMMPMEt856Z2/TkkpFx/O2guzjiwAk73UGJVdhRvBL9pQvamjU6K9p7Mp8DYm1
uNVAVFxgII2YEDDaLHTYW0ZZF8j0LHDSQipStxDLcVrxRUVOaTzECOhBCSTgwP6v
Bph70ds5HdtRHXmBYgthPNIqYreYZPmWvWOI1FUQzmOymkF3TlDXKDxJAgrKUE9a
yaPmLEuUyTYARRFmy+qoVWPPYQ1wOTGOD0HdqFoLp7/jLI82q99z0mXE0V9Q7HE+
OPxZeb0hei7yXJlZ7OiBggSXv+BXSlG0CRNJ4zhmEYnWgWdBKPtI5RA7CmhKnb4E
qmceZIAvX16Ce10da8Qh3VRD5YcNHj8EMgJ0IlR1Oq2Lb/Jwd+USCZwHprZ8NMt+
KRIQdfyJwVpc4It2QzGm+H8s4NNhv0/zLH6DSZatxGlD5TLOy0+wYtDiKFG8xox6
PGGG5feria9t7XWomDH4OUrK+AfCs6LzVRS3YWr7PMrv3BsxMFCq5FRxG1QKmeJ6
+1A5k3Qiw58SgOMNLMKPUtspBYOJ62XZqmm19Jqx+8EdUTjZDJ+YwgGmNMfNAwGZ
7okcP6pu5A6cvJEwlpiFq4LT4qlzH+4ml1T+laG9RtB5WrtnZJ0Q5zCC1qDV7ZZ4
feW3iweGojNBmjByU2QorP+zgCTyeQeoCN0jXwKp/5g377GEL9aFlt0mTGv8vk/1
BmOu+jMW4DhOuYUhaZhpFoZ8wHNSLzSNOo+d3ZbjzWPriqZx1tE/YOpZTK5fRRMw
KTLMNMF/ncas+E96eHJtD97XNrj+0BfjCvCc7GhcEzKVrzKd0G4bNVQ4lIXk1+Ju
vd5WMLB4iWJs5FD7YEDYXn+PTm2kCEuD31wWpG4SpUYmS00tZwkr2mufpJeCWbrX
AXbiFDTlJvfcuMPh70FN5xARHcHOk4tDHO0bsEhLhPHDO77OBX9Yx4+CiY3zEToD
zIw8Rq+lRP1ASiSx7cRSg6ssLbk7gdumN2f/qbDeC/V6Tw91FWsSLh8ohW3hhJvT
xA5qDKXOAwtundCeN/CG5uQ/b0Q8kAdguYy8RGeeg6GZbAzOK47caSJWTKD6igmN
MrMOa0kaT4cLZ25u0KrOa4Opy5yQSAKEdFFtZ9l40EB+gcUefVYC0JjQXSkD2Aya
iDr9bB5BMLDx+XZTMrKRQvxOi0RP0U0zsJ6GBkfTnUd9lrpII2a92gitbrspZSEf
ZwcEfGFdUcIis1JRfOL1sbRt6GcnLbhXyQVeR5OVqGswePYwmxMXODn2aUjUAVIB
aT9Mkd0QmcI+ZwMSA1C6ZFxeOko37UL9Ibd5xrCsAr9sPo7ID/Xo/NjJfB0k8wo4
76pNsMpKxJj/KpCsoDoJ5Nxid7zqZnFfUweIPkgNPZ2Thxut8GYq4AXqfKe2Esdm
fWT/Q0oSko2pstJDY5NYS4aQLLH01E9Chrhe8u12i4SqT+qI5FYBjpGFufLVzUuS
uK4TrS+5FhAo1nQnfjekFpnTLYbG5dbw3lg2ib/iO2xLDr2TwL3sQRzvusUewvP6
q01oSlS1L3j87WHQQ0W+DA3b+V5Yz4YpOqabGXqasQunkpeeGV+D9FJSLZp2NkJf
HyG1CQwhsyVTWEVpGPmcig0qUeOFFLbcTzc1+mI2ToFY2cVETz4biYoxRdBsT+c/
rrLrx9C6HCPInjB2wZaoW/Xfp4HxaMU5V/z5X7SfvUFPJO/Vkvh+MDLvOw0eQekX
DXI7DnlkMGPLpFFd3GiRxGFIBfH6Smd4W12umH9qAP0O72qZSvtCw8Jv/aNlVbUr
OwNhvbMrueozOLOXb3g9IjJG940rcaPuxpn6NdLeSBpkN/EtUUsXUrnBeFc8NRkg
oL/gWYBe7CsOgJ22eUoTbwP5sYGpOw++8cQsZJvb/6vazfq4NLeLojO30JJVV0pr
DvKisEwoQKo7yu95QNqjA0+/df6RNXXR0P8OxBqb7kUkhFwJ6i/dO2wcU05UX90G
uUmluTOEWzfpHpAWTE0nYz6jNJZDJ7vp5ne0cSdyO8KMdn0EYPQketjAz8oH15d4
/tp+ArIPletY8MxmA3YnUtbVjT4ebMumT0bvGe+Fj7ZHnvoLN0mqzO0wAUJjkByt
wY3HGrxFSrjI7IaZeoIQnxFfYJeqVJb6N6b7J7sY3j+oGYKS7KoJwFG3ckthKmZ8
xzzWZZCtl2Y6br40/7NdkTVMam+oLDpxTX3ApAOayOkpuuK6Tr6tmMfAi9A8aOeq
NK7Z7DbuujTCT1QJhOc9Nx2kiqiuMPBp41sxlnI6LRlSxW37Sr+gSeDV3+e4CC6F
2QuwkTCK7dZeRTYm2Yt1nKH6KqcSDkUVnDj+69ZZZ9mpV6J8l0IOFulPeqvdxOkJ
v8RwDPMuoTx6h1CU0H94EdbS3qxxnNXvMMzwRqDzYUNyxaSS40tQo53h3ShzjBtF
hZwRt6AqrNbTOGpjha3oKGc9jM1R9/lcCo2iS0Einz7wtvjTSta2rSypPbIMFH39
wQy+1pGNHhlnRW/UamOWb5YdSFhU6vhyTApveAhZtUJnmLEcG+h7dL7bOnBgiOwN
sci6L7N4O+lZpZGyh3Sp8nM4VPuHxzotRAQBqN3EFw/ivtZurS7dNjvIQWHlHpd/
fy2WXJfy6FlQ9C8zRHgolj4FQ3YC+BbH9pSUkdgge8K3Ybbm5/q4MbNYds5CbpWz
zIXHDTrAgqWktm+Y2Vv5E/DfM1JVtnhPMuMGdFpRJZwETJXLz7bT3MqYBh3ec5B0
AGoAAMsi0H2FYixjhrkK9f7uh7lLTtsDzMe8hqdGlmDPQDyidfXTSl1NtLFLnny8
C7j5UfFkFwF+8Tae/R76ri/71Vb48C9k5z/9yxzVHSIrRgJ/j5NRmXF1rnbDenVz
j1XZwNqcXa5NUZQDptgiL0abF5D2chXs9LPDlERwY3B+xDZWWEWP2UxDfxNIcWzH
1N6xuAUQRyMrrDH6eDAxZcQ8rdjdvmppcFVaSYw/CLEX0tF2/IEX3Uk393VWeeV5
Mcs+DKDqV5zoIC0EcfESy27oeTCQWwEjYOyD98cONhZEvK0PpnR0Obr2C/H+eBFw
i1+djTQOMwtKpPpUvFtUeCILKBP+k1Z7yrlgn3/QvqPiTjwHXUl/NByK5IJKxe9y
BZhgpZFhwXt8Cl1uqHRu9u+YTzrHRytFXfHKlVOChtuKwV/YPE2xUDX9+AWuevek
zO2msZvOeqbVQWFzWJhe+hIPaEmOxnn11S6SvZQlqg+2luXFQpSfVZ/kvltlyigP
W8e/9GqmeYmw1vfVzAGMF6l+U3faaUvfw5vycJSu0nvFXy1TASnPcc5AXDflkiVp
GIwp7N4K8nXKrRp3zbDegT/UjqwRDbl2YtKh+zO5iw1+7wPNx4YLUx9B5UiGqNZy
m/8o7QNd79Wla/kmMkykqRm5huRTGSgGYdQTzUcqLmn+CHcaI4xF9+hoZeNcs2D/
KRKZ2g294TI5LbI2jz+ET56yJO2cbbXs6KCFmG+cCLu08XZucgMRfUm+X2N7YZKH
ZTUz5lMFvS3AtYka2mjAGon5L3vV+pSsekONdbD2+ywWNDEkdaqSGOByVGGakiGg
veB52gp37t66Te0nyq3Oowi99dIph1+XvN1NTAmPbbO/8NmDP1olQLDmOvM3LUd9
RBJW8Gyxj7lho3cE46oktBvkS3XjlnGr5ZptCFDP2h7dR8rYv1fiKArFw6BuTmVQ
b7cLL8j39zo9GM3Yrhh/8na/vSm2LcSlIHww4rFYezK/qIfp3dZYsQszaz0uinwW
0g7wMjkVl5z/aJ2IaUkJh71pwAOwPriLvm3W6lrg/fiXNTu5iKQQyl791PuV+ExQ
dLtxiZkDxlxnv/YYs3HGuc/t+igNV04HZZNVMPjUlkAlgnj2EgurosiqkIPFM48a
g9Xqlz0WXczxnsVwkBJcxEjGokNIWsemeTfW06lZ8k8dK1zqVdb8X1+pScx9YpC5
Q8M55kk2oVQIYoa7QNQuzbas+4WIE7lw+X+HE8g6t7Or9Is9fIlTe1shg2BS8z9k
42WD8aF9nUKjcddkhjNrbW65gde3gWHSw+vBGSc8Txw99OCQCESiazviubFmCoLW
WDy565gFtEKdU4+sONqIb026XH26R8YoRWOoQL8ad9gtAgZ8DRsQRxHAq44Co59W
gZ+j9XQN/YyL3NSJ7Yvcfe3C/ZfKbMcsxV4VqMyMWoSkeLbXxEJl55u+iIF+VC9K
l7NJcLXQiWjJPCQCh0guZTibENw1ZoJiPkV4qTcmoU7C2l3oqfBVnVg8Ot4bDWhF
WDtm6wy6a6FtTmMPxz2HIOjsvbIM03NxWLTs7sFYxcyheNyzfYGIfe0u04mUW8Hy
b2+/gJZgvgxbFJ2HfKem5fBDvl1duPZmUerVe0hagDKHmR2eDoiEfCQgzXcLW7Wh
NMly3uQDj9RxTWFHvj8fjznJmvoXPxKPtXFJFkbBE7zaPf+nSeYRsFb85Qotyge6
ioO0YJIV9Re6mkn5xFBnjENW473rI4F9C0zUMQFEDZ9+iTy5X6PxgWz3TvcvbUoR
CKZMvNJcschl+5RXpjRYj76Wt+39dNTWdEHriJ9vIOFExfbX0l69C+gUxkvT6NfG
CWwltvEtw7EA0pEoMtrc5PywwzRU4dWDedBYf4nZEy5Bf27FeRRByA5bVYfnuErj
1+rWfWgBO8nXymDnlslJ9d/71VymwSeJdISYv+z1udzP8M+2Fh7xRIIIxG7y2eiO
/i5ab0ldCBqJx6Xue3h5NI04Od/iELDGNbkj4F06saNL5KEZmCApoHojElkmh8OH
SJoeoK1+W+9A1xQzJun0PaXgm38Jnyjd6KD4zIIF+5sLK7GGhpUnlZWHtkSQpeXS
+P04KKikVXFD46M0kZWbv4yuADfqlKxfiJUV7RzrpTnrOPeJWrhFSk6UHFct6TfA
Rn8PHumMQbNfWfOOnAaU+uJzdCWO2maSxQPm+ZPOlEjNiq4BJzZi8xhFiq9chmEC
eiIOwq7JGc7TqANiUQ4rv6SAFl8KkgVAK+q4K9NbP/sZEKax6K/2PripP9u6eLoK
MZmISdaM1O8W8bOB6759UnaaU3W9EyvV/sIFJNoRB4a9S5m2IWV1kpUXFutN9Z9m
rZfanxPSuy9STMYtB7PLq+Qc8dWk5PgomYNIT9bjxMpqIyeCpZeNIhMJ3yXzdaLo
vv07vyN6S0trVMqM9OoPZNqKjTIOCOy8kXa8JLKvtZEnuXUa3xPb7qcyplAEQJvr
jnAJ/F7Ep5nWMxZDWIRQAL5a4HNwieO7vns5+NjLwAFP0odPpMiJS6fzJ4uPmc9f
GHtxO86J++uWDo1o4W6mus+8Z7K7CDtjUMkqgZqGNl9gz36VfPRVUkovoj0bOSZr
Y7G1DfLR9aDpPlP3WH065CaGoYI40pTlhSllrW5P1n12bomOUlW2w82bMv5PBuS9
bnGpCnwpXvDFYfTtt1sJVytYn1dnzJ470NiI6LF8JDodwC5igYvv6/ILyPZsxVnS
WyB53eM6lWD1Rjpa81sw8HLjw1qtXzcmy6l29K0A8fqtswPcGGL0C2sFPjcnbDu7
ScGx+dNr96iBsmQXn2Eg7MNSVNXQ+v/heRecOmhVvKifb0xCF8YJsKzkCWO+UIGA
eC/g4iLgzjOIyvGQ0/43Ykk4YdzbApE/3wgPO3/ecba1ptvuPB7gNIkw3eUv1dVk
gsPu51fzRcfB8TLEAEnW7kI9Lu+Ua3gdILiHzyOrFxOme7Gd37OHFFfwn3Z439BV
j12GbKaS5o3QAMPoE4DUw2nFUdDXE+rzd7fHZtDWOjvz+HwTJL8OftHoeWroeBXG
qxKRFBG6ZunnlO+J1pfwMZjtZbCil19SIgrcXCKpGT62Y00WHABQArhtgKJ1QxNb
zaiVrug6TH3BIOVdGTmxbwpw/o1Miel7j+CHdFIAkPCTEljYpFCXbKlgRoCnOvGl
d07WI+nr8+hXOLdQgRojV43+OguwTDd6h+xzfeCqqB2+/l8fJYsrUiHUQCFfisM0
bIeE+rFOwYQ52e0vlJ3CbAetFDYkhE3ZPaVZT6JaY8JW2arKFNP0EE7SxWTZ2NUX
+LqavKy3HuZ9gkcEywL26jUVbsFWsFXRa+RTKP4KyPVgpxJjJRVxJ0XRX7HbXwWU
inHxdqoyULV6chdGPXMKdJFYTJv499uKrN1Lam61B6YXnuf2l7AjODxbqJRElwDe
TsBvSDHsrjvs4PvsQVyzXjN+QeZBwA/Wx29d3jMjVeiHZ2aBLx4c3rZV0lvZ14sB
U2ih+wKvcXQo1ysgGyZt0hE199RTBpwGZHCGAOeizFdCGVLe0PgMEeHW0ASNtYx0
pO4PS5lod9imYwaPQFg6V47JzEgbQIcplQ3pvVCICzU/fWQ/dy/CDicroRtUoEMq
0bZHXaAJQ+ZwlK6oZ+YwX3IzPmtIst0L9To5pLqs9z/6rAG7bMJA3EoZFDkWxsfn
gL3Wuu7S4IloPkYBMFO1P07MZcMGNzWIAR3rC0oGXfJgJafRCr01KeQ+Z66MTdWE
ObS4q3drTCqnM7lgHkBqvaUl4B9zBkdSoJP18dZoGVTJqUTFEEhKUMAYkXNiXFAS
nzEo0su4BW8pthsIxVt9Xsk+El52NlaxlCryVIFiiP27u6QBKUnbZIYVENOHeX23
y0Tq03PHwoOCN+yZFblFhEkd1Fz6PZxT1O39chqz5Vk20myeG694fwPiHyqvwoUg
Kr67JMxx1ggrdh4Z5OpmmSayV4E1aERXhzsca4ZNeoPIHKoIkWrTwKD2Reym1Gr/
xyHBEUasho9F8ti1tu5su8+811bS0taDuBuQEL3w88E0noEmi+JDoKTu6yHOqyhV
bBzauUbZFFmWOUJqaJbEgWAihDLVZtQEBKwvoyLitz1VwBI62rOLPxQtMMUOs/XE
7X3/ioqg/uOOVcg0x4SRr+mbSqOD7OwWUF9wvcjlDq0vdkZBHs49RsGmzn0I97cN
fK6WyCGKLNvH4cj8mNMavMBLN95hXHZnlbRye7Idqgya4gQpEOfcpUyxce9BOfyJ
6CiKy+fq/HMGpHBBTwuLZ+SMtfxB7pNz+37Sxkl6WrqvNiCwmHvaPQB5PHQMyz81
Hh+aKnPnneX/rQwWFvJkuQIb5cMuB2bTAj++nHcOYPySbhRFPDcQ9JXctlXfQnie
ewsg78nsay7Frfi66QHoLz/Q/4mlo0mK4+jvOYgOLODgwbrp2wX+h2BkVGL+rU60
uBycRydmX6R45gaLIW74W0Krw4B+9CzLRwPV3jFxVLy8mDs0+OLpNtvvYDPrUF/l
9VP6QCUVLNbKYhtZuMb7ZoNEkoxoW5uXJ+Cb29Btyysinq1eu1iT1Nrpir4zxuO0
k2HSEul2xCOUe7L7c31PVBbEYHTmpq0QVtLCktoy81gZHV7HIqn/kWwlEFBnoXzK
uwTIqKW/TTK2dd4aZIogW6gpsUwQ1UG+KE/esJsXr76Qo/ARlTdM/mUS/9mtmI2d
obDtJXDL17jQKIBW9HAz1EiEWZsd+dJrdSp06pO1Clazu1gA+LBFhp0q6yg2HW1z
Z1vjQUOA3SW9j6Vwx8MGgNSWQ7H+H7Dcua4aKQjBwUH3NX4LuwjL6T+eHeio8c2Q
mQPQ475hYb5Fz1LZH+L0C00oav+hX8Tntilu2Fd7VfiCz2ieuLVC9eXe/gKZTqBD
gtqsiHsehBFfqAhvFPPdTaFyy5izj76PJl7vN2HOaJFTrPTgrSuV29JxkWnhb+t5
slSIINeZ3C8X9qWKBu/lffghG6NwftcQjVkjRVb+GdQOqip4mHj9TUV4PkQC2b2s
nfuGFVc91FHBQEGCUks5PChE9eknhaLUxe+3+dQhChKIM/LqiGijhoNmxI6TX1Dw
tRGy/BiTjA0aCkER3tdc85J7dWpUmNYUHrgpfw2Qn5HJbK499MSrV8bZNbZshm60
yi3Kqjxe8i7S1tLTYPVzckBYIS4XAl2OksDChg1zAAbaaha34fVzAEECf4MPl0jX
V8PgvLQ3hbhc7cbBwfUzDc+JNh/R5YpyRgp8Of8A43jvKVaJwvpLkqZaz0MPdYaW
TIuR2CoeXv8uU1j/dNhIL7vBhWzjVwxGzXqT0onpgJsBF2VQM0Ewj7fVxcnB04Xc
GmcoX72KTB4xW9mm3XtO2T4abuuWyo3iRqkHVmZyO/JG6QbWvgHI4r3TGIRJSUDr
3FuumjdVMLP8VrDHRx/g9dOfmRuZ8j6MW9DotR7gthCYe3oEh6t4YtTPqk5x0f+Q
cyPEQ8Svve5WXa1yHCnmCdBx/Ntl05LmkNXs3gdFRelBhQlDtyWXenodySyb1fYl
XI2RXMm3STHGVvfDD5Y9leIgq9rfd9Hw+QtbWjuqeDc2gF93IpjDKVoqYnoMM57L
WQsrmjGxv9MThfxapyVAMioTOhHQWxJr04Vacfoaq9M/4srGQyD5kLTZODNcOqAw
vkLqr9W0P566lQLGgkM7fx0tsXjALJJKKj6kMjqleOT3A5WkVDeTuLuEL0yRzBJV
/TtuuG1LwjA0JSPmQb+Emlghi3sMgdqKHeg95z+JJkAhldoP+2rYSn7Jv0Ulo5P1
A50lzOoYd/M32xR33kuox7Ei7k4epO4pa+mlCXgigEt/ZMrM/Jpk9EyfJMYjDstU
1Hfr809JP7mLEpuYJPF9H0qwgzWYGaABWIDChby4DER0pln8bMWOIfeiF37u03Zb
GpVVg4+4jmdjNgzASKu674e6NPVGbgqAtW2ozxr+toTD8UPeS8u8n2kV9YeV+BfX
bRZV2daYk0kIdJkdeEtI56KvzZrqhZrdBhdX9Bfuy0CciPQJvqteDZgoGR/tY9pv
neZdf3Fmc4JwfuuZZ8LurmWc2rAJ+OAe28xwU1rOHjOKhd8sOCKgOIgal6hxsUDO
sAnqsHWlgI3WvsXU82UNzo8xvUq5Wc+NN/21sfwFiZgOu+KZcnKQ+fUFaMnr6jBM
iKse4vyyMshdGFSlRd3WAdJUWejrimqG+wcTRzuYat0ZWj8MW4UQObsF4YR6BLpI
vqWaWP+RYMmIXCA5r+8Kn06ySoZDDHZlg/LWFeN/mxR08hR/UWF1lJ3M7kqXPZUA
Pyr9qEQ0EuOGi935bBtZkJIgXpVByg31sJ2sFND2oiz1xN/N+rR2NemKxe++N8k6
EmX/pJT7ZHPgZQjy2bxOY8t7eQ/XeiXIBmAcC2lBs3F7XNEBYMqDml1kDFhAgM63
9+dG6NIhZXSWsgmPRXeFkK/g1Db45MzEjZk3pGyF177bMBJBvraEMPluSFWrB6So
nXvlNfmPlIQULw6gZlFXxgx5UmSNVo1DsCB6OaAghmbLZ0lZDyrpu08rJ76scFOP
GZ+vKisaSIPnrrVfOJEXfPNz3hoEmEGEEeI4iDOLQjf8MCwxA/C0XlpI2ZId1Pi1
R0ovTBvIIilD8leAG6tLmOwWdd5HCiXRVhXPVOFlEIdPMagl1YC9onm+ZPteAexc
JO3tuzQXlK2LKy5BU03dxjCkb1oegNlgB4X9j21U1+SV1/SEBCZn5tdTVSKKHgna
T1mDAuxCXh9dVG8o6u6A+8agNya6OEVIUkRf405OuAsnEZH0YXzezhXAYmjTEUpr
JM9YEjrslMOyZ18MvKGtmrUfBh2BBG25bNXxl8aO7kQZ1draKgNo9W2jCKSimOjB
piPQvHNdp+vFgQrY05fyOW/p5GXfN8eM3ElBYU2dYidb2478Qv2d+5jTuBzmYOak
aW93bemY9wRc6YX1+rW9gsxQYq/ZuM7Ghi+o5eWp39j/rVpHhBGTG1wPi71lBLiq
/iqnbCLhGZSOvYOXFQK98y9/LHQed7ZT5Rdy47hY6tc8T1DH6mmdC4D2UGIaYMKC
62f/E5OEuiwOIrJ7n/a7xWj7Wx/813EVADy28wxJ76ZlP/UEtnOD2kZQRj1Q9NbC
PkHQKgSUEU5+XPsgmPqyuviaPsU3E5489H8W3ryFmDoLXdHuajBev5H1+/dAX6ig
bQFBGC4S7yNQmsfBrRqSP4VEOxVqkS3HP7wyhwMIFvSxwOTlJ2TOCR3ZP1oeWQPS
zlBLTAYyX9qum2Wl2VukM759lGzw8QWX4LRwyxptizXpMbiSVpzu/vdTetuocM+i
TU92Ggo9LFRnF4eOKhkO9vIZ5qD8S4lvcuqQiOB6pgF8UsgP24laRvzK/XyMuWn7
YKiJeOIVhsOeoBfs16wxATWFsg0b266/E687HSdy9bjV0xnYLuaY9/ALC98i0ZFW
3CCMtM24pxSFStq8OSxDKKtgI//Ye6uJKMCRHpBtYUiD78tWmiF5mPEo39cd8SYR
cQxIqRAJEt+dVYi+bXu8s/hsjv7FNR17oWVefINCMK18TcuZfkInI++/3mjJOXp/
oF9242z6TD9qHsUv0YUe83WwQvjSOh5+UJiZMe8cj7zoCsVp6bJbTg0U1jgloQif
YsUXnDiVeL449y8Z2VpNn4tHq8ByiN6OllkzqMTziNPQWYLVagoaMZGAwxSES7BH
98XJA7XGyW654jarr5vZki2HMkOjmf53KCTAel8aNaHCi9G3LjlwhFdCIeKlcoUu
q5pkI9saQt16ePf5oipTebjWTwqss3jZfI0KgBkM/v7Lmpit0fbMg0br/GdDT09j
NnfV2rlc88m0Bj99d4TsdAPVzqEnLZu8C7++xsHtxl9VkLkGIPS2RqOVFLmhqQ3n
ZRPkdhTuAyL944yqEJtEaojGf8SdTOLUt3X3INNMdqG4GDKBfjRqoiBiQDEeMX1i
m528dgZ8yBRaTLFi5vJcpXZNBJ3BwqORfvWkPCUxi9+3XBSwLf+jN5opyLv93u6O
mYy40F+pDm5usSfmJhYGUNvEl7ebNxnJCGIlGLR5yZ6KcMHjpHTI+imjojEFFPMH
UNmSbRsHKMUtl4tvPGLUL/1pGgEQEeq1Fz2iEZRntk2sdeX88eBPN+vjJGXaFuW7
a5w9ErNjtQCHDhSrNTm6/WzsiCFMfrD4aFs47Kt9CwmE2B9jzUFEow9qIAx0y6pZ
CeRMErP58PITMfqoXu14Q6WLCIrL1sdDiKoDh+16VrmJORcCJ3LG5C3wVDayjZcO
z66bVXVDF4bAmiWjF+h8PtH7sAStOOFPpfmQUZMSQ8cMEmpasTc7VPXhLiMC93Up
PTPxjpbLaimeEeQL4goT5Q9ccmDYo6li5rBB1rErchu9zGyuodBEfFmqV+a+Qqp9
qWVRewhGV30ZSVyGu0yByySidBojqVhXTfz6P6vMAjqwUqs5ztqwgWSuRMmDyoRt
mngnwrKFEMMQyz8+o9ssNTpdc9b1PY9j5lWPdO+eORf+bvyhUaV0JCYJBTKtrAnZ
AAZKEFKHGuDUdGGlOg8YN3gRMhJR/OGwz8sbObPyUpN+Kdt6Q7DQk8A0HmPtnlOu
i3zj/yIyMBoXoJkjaKkd5za6cUbrybdUF/nw+U/XeRRtMTBXxG+c2E9mWA9b9yYD
kYBFF9lBqXnhcSHGzSMmkAhJ7egeyBg0HtTbY5M4Qgyv5tWh/Bq2O9FN3JBmjRgd
VA+m/vSvuQXd8IFqgPbFJl2p5qqVIrStrIamdosEqoQPvntr2/3brARQlQ+48C4n
W5hfs0VUKPUiOH0U90vp6sVmQkSDcy1DOMca7XsYEvYVvO4YUwzQaplwREaTC5uk
O/jVXPTN/P6lsRaxygUab4S6G1sX+VC/BFhBUpig6GmklmBQoDdS7p8rHbewVFwC
fbNaHyNVmj3bcATzP08mMYhO6B3+UlWXpgFiJDwc94mu1QwxC3fET2mf7OBU5HUF
JCS4KH+7PhP1ly4i8nzrX0RMA6le2f7d/72j5TeyT134Q6NAIMrv/+J5O3AfGW6B
e4ZP92wzuFsHDXAvSN9uosppHXeWgp3mzZ4wEn8GkDA6F1v6O80l2JbvNyfPrD2C
pIw8nT9zMBFwqEPu4r69cmDpsv6EZnUQ+iZOU1ZfimUfGfEbTIOzLfnGrKuQY4/T
O7McMO3ToB1hJdS4q4k+UVkGKMpHVOcnlCOQhN2I1CRVw3pHmGmmadKAZXDaUo/r
9W5IPNnL6PcGXXuZptlzKQe9W5mZLpct9QN5K0rMOnqZ7y8Cv55xYVcl6jJwjJZw
1IOIag6VMGk7pyZic0nercEMWM2K6HqZ6YHfW0JyfezISPycDFoJfUk8wiyxSKu8
liFVdwuPKeqy4qS0loabDu4Qj1U+F2L+b8Uaej70lnf7z2C+Bp7sm8ktRQw8MfAe
JfCKgvInzLu4yKDvdwERMAXPeguvNtjHh/BGfFX+B0JMego4TrA7ogO++o8rI/76
zQZBzWLjIHW5lReUhxeT2aM3kDtgfmJ8FKbH0zlKa77eFphJU7Soh8C9PO70ZvJe
MUwdN6UpEVISmG7+U3Q6byDe2WqYXXUN6NUzNRqLnIXjYrNzABiDjQAtmsPBeHzX
3NXG4MYG40QttCoLb1/J5dF5nHIosE1mNMvmdHASTzxKK2bcBq4khTsP5OtDHYKr
RhX5E0fTWpXgp++QFe14ZOpUqZspziS6y+9wLgSk9bL7d0Rjrr/0FlFoCUgnGEQe
s7x5j7PxFkdZl3zUd0vALprD3HjuVPHW+G7P0yuhNbd8Umh8BKUY24MP12qDAsNU
7VyTreZ9ow42fuIwNRrwkpLl+AoLi+jFbfEjUG/USbGTu2gWYGgjapqItaYMzMBE
+4vzBTmGRuSZa1MqontgpVWDSjkklYoMA8xVICg8dfteNcxLC3V+ot1iMhRRZUrO
+UoLsxhlFXGnGwIO6bXEwZNiXC7/swlISzXm4lqtxambDKG5gd3PiYxgSxIqgsfM
Z5Is1OBC39/geerQeRUoRwi/KwEwGd+g/ikVEj729OwQ3Bs6dcat2YLE9i3N3yNl
3OmWPLLZDimG2i8+JWm51nK58Cpg7xmzl888JKVAhQiFKTy07tzshDppjdcdf+aS
PVh3DIi5WsnKSkMP1KrG0sc95QCwtz9ORm65m5FWJoe8Npklg/9d/uV6bGAmBa6E
FKQ7hLweD0+k8Zb7gKvDlKya+iioi+QJyQTiG2zpoeywEQG3e9DUv8PdMh4Z3+c6
Pr0/0SkCOopnjhY8c5z+WPqiActaG16+oIM1r5e+NlwaLLZPEcVwCPQUW/vLQwwZ
0s2Sfvzw7lCTkgCNzQz4pe3DRLGAZUUZGpOQfw3Kef0teiRDeMiunqtneWHPBY/B
tthxK2DITWgjpdRYCUCV0M/ptqH6QT9eJd4QycCGEWx/sdMPpehDglxMHsqXyRHo
4oECIgllLXrGGAvPtIuo1hgxmIdzc1zlEL7LEow0uDtWVcXUEso5Y7IqrKynlAr4
5bjDRjo4iI24qGptH9rJPlAEJX3n0mDSHdc9KhweJL7DL4SevdkMnTFPEo/S8NsP
+mJKgxgh+Tk5nktHuxUAyxXwwUktg+6T0RWjbnCxGWDgFSBX9udLqw1YXGmvno0i
PUQh8GfitK+v9oUyYRX2wfGroJGg9DbTJlP7zphTbOxwoWE9qP6fHkxtBEazHIFx
auf4J1lJGTzbhOlccbKGi6jn2eN1i+lnIkQfD0LMxRjwiKPTwcZyOipI87zSxzvt
v6xzkHLAIkkehREdzzj/53EXrZHPJ/YYymQCO8VdKAptRn+iEmjUZZC3cbQeHg+X
O30xfTKRzK/UuRDEbJDgvkV/gENfly1V/+0YT/S2jS2WTRmzKwTfokyt7rn18R0F
+iWTPv6XVVlHHEEZrCOd2VcQWLfb1WC3Yy1X3Rf+2k5Z4BSdBU4npu6U20eHvj1l
oU86DKBWFClNsBNgqYqXgmQvvhR5QQCQ+T+yjczrtVl7/lSqhDr19zNT5R8UU58u
0a54qy6RQ2e4vWyVqJ5iPLbLRuynDziz3CNOkLjcAq+8ZKZK3hzpJWjT19qI8oQk
ZN+Xgbd0OrEMnEwkYLYC/x7KKfQKdNo/jWEdByyofILXpQuXmg1knZU/5y5pCzHh
GPH4YOzTQsttZ7/OIVTpN8J1bNqxZboRYwa0RT/9qFhUdFlORstNTcgrpOC0J/L6
8ZZEYG7EzLomD9IZQY0Ejg+wK/QgsBrFKLvbi83BrxhIq9bm+E2Ia15qJsll6LPu
04h7N8whiq422AAdrJQOAR7DFmppFK/CierBxoyAEYqaR8B4Tcb3W1ydxHszgn4I
n1RmCTQRRN/L93bdx+40Ki+1ZO+bxIUX4NZ5E/zs/M/oV2lsvZHGTZz8kfaEIbSx
h2ZL0e5O/hBPuAysyM+FJMc3/miqwANDjD4pAgEWuDVH4apIPIj9z7PIi2lWFYkb
muy8eVnnJIbdehufZTxGc322WfM6kJ9iqN1brWAtbMGB5h7b7xRB/heNg3x4gk8h
m+sU9jwImcUspqgd/Hnd0txUGBHANbj2NdwTBjZGqHXQaWyktZak4VsIu1KAdT/7
pEWuHWMOFzHmUaDL5oDzZI3aksxvJYKpkIhDkLhxmOGvIRS8ze1ULDgDhZYCBkCA
lJUO6c1jsMAhVPozYzMisKU5G0BhGzXMkUOvm+9Ob8RVF4sJF4ShXxIfUy+5JrSB
9GECGAb9vGyH/u2dudhmJwBoD5IPL9mZnYdub6Yp5jsHHN1Lg/8VS4LUhDJGJ3Ae
QXhhD4ZFQ15RfpyOIu8aRQdu9aBT/xkXy+ZsxBYXY7x7jVM85oIPHSD/6905BMQV
hZIjdfN7PH49O/mUvHN8DaR9IFthwA7svmELjsX5vmHQ8w+1weC2QLlK0DdcL0s0
orBSPvEc+tyWRuymHBRHkEmRiQkAmC2pBBAPxO3g209AiGLRxfm22CERYwgtUrsF
K6fzt6Fpr8JS7lT8XIBJxS97dVh8OZw6EZFKjnQk+D7XQKDSrR6XdJJQeSYsFuZN
Lm6ygiGEfYpstHa819Z6Z2xT1Gbky9BhVqhSheds0eK5BbbTOGyL+Sk1niBI9/RO
8fvTyQxNi5ChFb7fWMdNc4OQp9MlUkCaVxX7ClnRHDgtHcVr+4c4T/hhakyXlUW1
fcM7M606axKPwBHgGYe17h4pkF7mnVb2rpZwTnDVzhbPjzlJ3beysUbQdKxurPs3
OAKKe+2usrp53gM0O0doc5n52t2HqE7Fcfvs/hhT2xLRVKj1sF6HYB5lFmudhXQP
Nc75qInBmzlTfmgC+vwlPx7EDl/RqQ7DJwiBP2wozGfTWiZlYlju+cqtzMI8IEL6
zCSvMi5jFB71PwbGkmV39n/rF3VUkb8MxLOWwQysfQ+Xpuvt4yCoUV9oV7A/cdbQ
+2M/Q2qRdZlDJCmPeiM0dMIdoKmCF20Ves8hS9HSlnR0pa44+0BggAOhIDbzAlTj
f470hxHr887zWPvVE/fjPWw0LszMxSZLKFVemCRvivbHOguPHkO/Vyoo66b9EYZe
5foQOwtMr0p/TbeB9kAANGw/p+JCOkPkiBJMSSXBoVnqCnWAfNjMHFl99lB3bwlt
VxH8TJBvLXGQx+ycC33hS32DKDpzIBBuSJuNS3UQ3OFFG6PHF2H7/KK3uYpjUyIO
mlYDixjJ3AG17kOxx3D1p3cVlLqvuRmLYLbE4SYGEsTP6rilt/02iOmBOAA58iew
L2InymzHbsQTWNdRLcQm22JjBLTgv39ggvJG5gkN4lfvprSfSxFZ1wYm5UtOAnZ3
cJu3v3VhVaOWHlmrTMDKxuDKlJjcgAUpeLDwl03AEG7FA0uoHM0IeaE3JC7xGrw0
Ta8D7rl6FfZ+5Y1EIK1fWwMccWxz7F8Vn1x62urMUznd/eNMmmaTCPtBmRbGPVDP
sRiCQisrFBb32Yq55vKQZwRSK4hgnYASQeD028iM1wptXaqCCohhQdaR1FFYmKDT
uyevu39yQyh8D3SL7dul7snRUXXjwfF6YqrJcbWzpgh84sdT0amsB7JDYntPLmYq
Jk7SYjBkPjKsc90t7tG2jqFgvtXR5XnGy4azPH+Py7FGx8cH6thRfDhGUQh4PnO0
GHFq/9EsmvFqnofWEaQDy6B8KmWU7cU36UQ/1QnQNHj+0/KtYRMHH8Jlc2c3Lwbw
pWRSETmB2GfyjmXBemhtS9UCw/Jjqf3LCmYTA8lJKs4aY4kyNwvjsK4qes7tq5Lk
R7VROzwyQwmDqphLnxRzSiYskZsDKxryZGmgp3W9HvtIS37M5lZTg4ZtyVmmsN4C
F5vPnqzWw7m3lQrYbTGSKlNXkuHbYh1KKX1bjgehULqWdOhR42kxBpHRRwCa8p4g
DFxrx4sgO4bu4FbxTSftVF9tR9OqmyCMtx+yGUWaG3wylGRtzTsdUA+hFxgwzxJo
gQe4bDh8qRNruv8A64ZgIY0KtQbgILPDPlgPBxF54MERhhZCDvef3auFG/RAIx5B
IwGNpkZw1nu2MhDsAC0ZOzvYZeyAJRU0FLbOjO8pHcFvY9EZA4TYuMxTGdtrijeU
zQTu5eORSGhQ0oEUTubBk17dEyHWxoJuSlmmjBB2srM4oz4I+PnEt5gENQqg0zJl
oC/IpH9zOvyKPQuyQBW27ahqAusPtL9dc2udvPyU2TLi2toO8XuveN7WJDkJHYge
ASLaRtvJrGGD21vzPXgzzthWBVR3mfeNnioIEYntkM9wde1t0nvrquFY2cRp2VRc
zUZKhqvymr7cZL6HZvdqwmPs4T1auXoRhomcMGcxvfDSbRKOv7gF0Unt9x91Zjv/
LwXaLhziUkbnB42Fwmoh+Jd8Zc4PGfeHa1yJcBRbsUFI7OQKFW5VduOtFhGORfic
BP1mU96dSJkWGwzng9Mv1rPgUdK48oGdW0MPaG6La1ORYs8tEPxo28bNd7sG3aM7
FH/1HJm59nd8ZY18cX1FWijgyllKou8me8AQO5eu0DYSXst5Cczv5i9DFH1u2ClH
UsfW6IDC34BQ773kpdKR3nNxp4D/p/iDBcEw24TDVkPwNRaCn9PpgeqgFaeyfkrk
rpRJTIHOJTsLzFxc7zhOnOwCXd3vw0I9zevMK7jPoF3XqLB7vxwlma8abDSO8lFY
yg1E5yxnw/FTbLHce0hQLwzSmey6C66QGW3qCB/DiT2y26eDWPJZC1R31s5A5vjZ
e7jRYTwHbgh5meND4tg09ageK8z4KRSplkD/0aecIK0KdkUnX/vJCwo6tqjvBOyv
KCxiXoRX4617y5mCrtVpAlkGTMTRpOH0FW5wZsKSJXEXiVz8jo6HxM8o577aKFju
svU6elXS/WFiQy0FnRu+ZUIxq1yx4I43RJsgveSFOux5ya7SiYQglPpB3kLE7pk6
CD+MCNqPOdspF5XacvhBHTFJ0fRmhFIyUgFiKvvLOE4mshRxx05V69YMMMOJ1DU+
7So/l4dzGTuyjBKaYBUjRmJJVg74hY1CKp6wNTjulh/a/hUay6eXgLgsTrPoXTIH
LSvQ+cjjHoIxhYF2Yl/w8KIQ2ddt4lDIXmBh9IZoTuaLhYXRv213+5g2erlKtkeQ
xfsJjYJvfF6eoHK/eoFGR6AistTr7isY5O2tb8Ox8MSHzy1LQl+ccuxYh0S5BagD
Fab7EaF6sp5p2zkNkLvnI//E1pfHQcBykPSsjSGBoa6OGgKQlQDcUiKGvsA1iTm1
acqGXs5DNvoHRsCu9jn0AFVPEBLuZoahHFn2RH97w22/LlJ74ZzXf2wJf4T3n8xI
KqoKHLEVKVjIzRZQtipkMUEC81lN1t8t5XJ8j5qFGxhnAv/aH1ZDlc/ZLz1FgFIe
NQyupd7cQOo8ktFwVFRRD4m9teC1DRf0xi5jCQRT0jVlLMYa5PygKJdqcpmvvL3C
V4rVsMBC1KTyB1GOrVOAm+S6ljdxxWIoOZFKJC1dFN2qGsmVi1NBK07BisOqtM7F
uJAvMEpdvXTN3nEz0nboz19ObYZt/WOUxyotsklGFldG+QSTby0eBO0P9vJgda0m
sqvDWaUL7XV16RgQTFml4a6QgULcbm0VsibB229jBaE2A4AgvjZCsOuDjt+SDECq
zua585SqaweJgEEhR5Zxx+VInx0c/TAGm/7uKEniyREYXmSFYQDoPuUly9a5uND+
XOE9b1eaySzzY4a+cIF8DIDbtzVUZsReFApQcIgA8Z3OwCP6+aKxWPh9nIQ2g11g
Cv5SDOKpRe2TqgO1RVdMTbux/RYHhPONzdW/WOil9Lfmhdnqt2NYKXbgxEaHotAy
wsJkxjCXCQcY3mm6Nk+CnYxEY7YZEOKudgr2EJl3wZaIewmcyc2n9VQc5or2IWl+
Fsyw9gv36+S0Hh0GoltHAT7Owoi5d+p2mGNJrh3WZeykuDPgjAiRirSzAiKL8817
8Nz1viLz+r9QQyF4EoRPJjadiS7M5Gt1GTI9g7qt15mmsA2epBmYHNN0CA2Fvyq5
e4ingg020xhmXB8SuuYTvICpLQ8+aieG10BS0CPh4xWFCz9X9U8wzJ7082jqApll
Ig4P0+xlHOEiMa8Y26i8z/vD99wp1Vd30/tZ7DrjPyD1iiFN/pUl75ShIxH4Iy2P
HloqutfJJXle7J9XYv5jaXeOsmE8MT+MkDaAd9Q2dIzJg1IuxvpVtkARXuE8J25F
duzyiaPEusHr3JfU6r/rG9/Bwp7QQgENIGIjyyCqVpv1c9og7mxeD4LQJShOUYIG
BqhZHIBAjOKEb0kcM/sXK9o0HLM/iIqaKzpi+SgyToNUJqsSoeEwbrADbXmt5YFw
h/1sIcokLwKLyp3r9r4U1N+JIcnfPYXGEV/3/Y02AFNal0068YAOwDSYq0JJLPQ4
RgsgxSAb4dfbFYVzQPeBwlGslREzS0r9SdUhiiMRnfkQa87IjaaVyppHIGx3bgA1
qQWDzjr0nkQaXUU0JfyCyx7361JPYHUF3CssJ7Cgk01ouZiMI0Q78xXzZQsg91cf
GLibteFmOiNh35HOqESRRjiJgpyi3ADujUyCfBNE/RzBgYFaXj12qR63h8mm4BbB
l48jyDnK9lNazNxRlQlaEP48hnIKHMkTohhTG3sDMpLljFStf+3qBwoNZVrrS8UD
p7VyhDON7Ri66bzqejwPB1SDyfS7n48Kxz3mbTiREkd6UAfqM7fiXcVm/P+0ZP6E
5qzl3tfqE2brVE1m6GZJGglsObEGX4+ekTVt4saNdoiW4OrS9bx/i28rim2iT0yD
qr+Fm2ru452NM2FAGDuJyP4PvcwJtCpWdScVK5yizPWkPFgyWKYbBRxNZdmIA05O
+6qNR2niRYf5Kn6UPVVqfD1PT1hugpEbmjaFHvxBV/bkOTjWZB5OLpprKOAczZ22
RZgHg2aZEO8E1nPyypzivsxAq0vG8fRXiWL5DyG53iXusYdpXpQkisO4GG97MADU
gW0N5nYCl5o121w0IkEjubRC+yBEIzsIMwPm2ImtB7bHhZc/FW0Gpey4cExmLJVM
htMXuMxvYiAXnhCQapAL4l3pnt3StBtgnP0TcQXzhvvNc7fd3cb36ukuOk1B3DFk
sh2/aOlds5TSwUXuJ0byBs/qX6hLlVrp7Di5+e7wr/vCgO2x1MQ4vibr2H1wVy/y
h4DIQ2DakjStIKeepgTAV5szCWKVaa48ZcTHiZGtlMBAO0nYB7wXHpqPiWNHACQ9
EXjPps8mpgkYsOZoLbooFFFr+pqEUuazppSS06dsaWF77EUQLTyixVSkUP9EOCyR
HVEkpRsFs+1DTc8lVMI1eYYBFUgLNZOaJQ8C5yvBOWthr2BpArtwa88V7u9vfo2r
VbQlizemQO+F+2IO7L+z4y03iu7xr8bH/F9EWwioEHW0B9PVtuuuSMym80gFHF6V
gHzDZ6KLj/ClJ8i/jbNfixxglfprbqOXXhSAsbf6tjVOXYHLrGzQ1kXE6cuE+3ZJ
jBJmJxkXG2cZ4FBKZkrxOI1wfBWBGhT2VxhWk9SbgahKZndyQJeWFWXB9pepxY7j
JR9wPfDxWFMb8ClolcjFTd8fIya+ua2leyb9kJQcHdDCJOqJxLxAR3xnpomO3GA8
cMCRPb+b+PN8mlVhgPe7GiVNmc4BiunraPoa0BJdy9EMAjmuEfVg0EmdJYMSHCwx
EofgtSd2WQiTta07d4GxI10NcOvkF+Wh2etSYmPGaYuKJry/m0dWHPqzr+M6CzAr
FVnbJGCnV3aZ1rEaLYbI9+1KRH179xUdz5uoEGm9vXe1pK6agFuWFUsxo2br1nyj
OHtKvyFpzfFoDPUFOp1vHNbOaXBki646kwZl39zmEPous/PngUBkwk8gdCTvLcNa
KKu6khfLJmSlcpHBxvHFSvXcif7BOdhkwYXYx/r2fKFxkS72D6oGhBqOrw0fHKfF
mEO0yaWs5CPEa3aBcTnD3Dy1evvfNQKdxApEzxJBXu6ywNo7B8VE/UxevtXyKobw
AaNMhDDjlXSmpnEwjy3XDRdcMsWwk4Ip2sYFlONhMD3Pa10RFVfvlbcy/YU4msuU
XXYfcevazlhbUsUx+p397IjRL5rd2+emqFQV6CcCvKVgyKoBF9rHjNXfLlN5seZA
ryPBHpvBEc9sm5kWaBvcT9O9DCi0Ln2xH1a/SyNNbZlHRi7IWpCKeG7d3XSimmMA
QDxkkK+W35iUxNyrVnSQgjaw5G13fG9liI0xCUzE2RaR3HJVTv3P4lOn5+ZvjikE
pu7T5c/HeQtzidRLKxP2u6x+izoN/a+aWhbLMxBN6A6UmBHTjQnerCiWIR8gxjT8
g1m8qJ24af1YPUurHCiM0biT4LnMJFile6PgOjunKlwfG8QX8cFu2A6aHREpLfKB
eqC+uc2fks5iYAGPFbbVwhWWWv/NX4M3fyInJdGYLWV6oqdxbRTB/zDI542szEkS
Fwe6SZTfR4cMOnGOduVHUXO4UsUSCNZQDP0J5vZQWyoWGwGtu1/rCWjcvN4RpIYF
AF3dKnqShSmUkrdGH1pQEJoZ1mOMliVRTPe7+8DYT9BoNIO2TmlKkuGpRIvV5nUf
i0EU4JkkMwh5oEKWNrOIc+UvvoZ/wqX8b0GmbHzm8ONrnE83iyHLHbED0F9LC3ft
pHwTVwI/RXbnmIwrQ2ZAKBF1lYLbT+1n5uLrR88sTxxLbvpwLd2E6GQiffAodHEn
Lj7JmAz8zQmLq8qKkNyaeMw8NDGRgvcWYXwqYk0Svct3m7fdlH+UguNHut802UKm
x/QZEJRYbMQbDkjkmUk2x/41LKfRC2rWsNBuFX/vLa43QMVFXRIonQ1D7VSLqP5x
bQrZ4FHBybuey3bcWw1qtK4LhlFtWI8SZFxmEd/O2Ca/tC+AId6F/lVa1YhkhAJy
+iFI8KV2bTC8qZYhrZgzRqCQ0LYQPQ2yx9pAN4O/m9UiCB0e3mT+11pCPazaNb5T
nKdR5wniyXjZo5iY1g0F9fbYs/IuMDEjrXchr6QoqglISFnRfzeqAAbJCvtx+U5q
vBGUhRvSMi2Fc488gNpmg/KX/JjYkmkZtOxLLzap/8eih0ZuJfN64+pHuf5RGuW1
yePjZnS4pMiGv0ZPVzk3Gdxe3Fz4iGwK3lPq4+tlkGixo3vzAGX+W6Mb60RB1fkj
3ODpwDxuIlm6n77EE4Wo0SiDbNgEW+LKjX79D/79vxosMNzQO2NjDAYvu9NWk34u
RIyMyazoWL2LZ4e/U8Qi54UC5TpuEjLyGOsk+8278AxIE8+YILJHGg/UOrnBDva6
Rvr7Ka2KmJYVqxlqZ+BJZesehtr+g48HM7hHrWRGelyK83RTHrURwYoXPObFw3cW
udrEiOGJ2EEEHp+GCTjSU4VJxY/UyU4piBMA0Oq7YgB9pgmoieDaPQOn7kQsDNWh
AMwNbemFJsVWNelHmvixkfowfeYmT6OVt1UcfH9kRe0nEeykRxUWpLebHRWB007S
1uvEV/mPAtfxpOmj43N4XFVtxak0biXWGMgQQMtfoY6Ryp3ap28WS/qFjBfKhoT/
tcMoNnv2drfSLQesl3dOlPSF4Gg2JUjLcqP22vnjh4fMhPGG0EMOIa7VJlkRe5Xf
de5QVaTc+IvC8reaiH6GX/2mrcocgHjqGc9qnY1SMn0mkf+xHurY0wh5InNQaQ2P
4MxFowH2z6uow30A4TtkA6Vvx01sr+ByJqQS68ctWq8Z2BoINwzC1dTAIlCkmkz+
+Y92mw4lkPc64jEPRMzklz7veE/yYHVf/w6wwporiNKWxC7HU60DF8j8PyBnFAgM
SaJoXYyuZwSVymNsH2GbJzGj1bgVbRnxhpEa8ZubbJIWTnVr+5D0hKl44NInTJOx
RgRDYg8MeX1a5T+wq1VGF0D/mqkQzwr6MCk8doHWnsb1cm9g9kD+VPDbhZuPRU9p
e6edfdFTP8a2Yf3cxPS00TEfmCG7OsXSCSWApIEENKaUsMNGAHbPz07rkwTFg8FS
j81jLXRpzGJqyDIJRg0T6fEpyY/Eq2j5FlUsdjWC5B3TNIwZlyGOqyf3NzsFjv1Y
Ka/eJynI+4mJJHmtQFtBvYSkewfovZQlPm/df5DRAnPlfjfv0mHEM1RraLoznKrH
kkgWyBifdhFb79UYSDhYabBiyNCH7phIVnywUhuxI35FKb+O6EmqFjPb0p1K2urR
fko24q7V/SY4gQN+NRVqFgpgqNJP5tQk53/S+kSyOi5VjuvXHjXRSGacA9UnzIjj
KLoE6DfHD+2wxViXqj9iOWNnrGv5c9iTdSCMmUj+j2GRyF7nXpnFh/0wqf79Rpx8
h6fPeIQvvKwXg/WbAhetNBNxiMW826Afw7wbo1vncfWuCE5EwumSXe68kCP6M3KJ
qWn5EABp2Jnr+lhp9GYa0f5BJKBVMYaimbXe/Le0b9GbFifDJDZOrcUCeB66uGtO
7TBUcPpckmOlqJbeX87XLE6LscBrz+qWMJ5VU8N/vGrKnC6bu3/UPTgxjAJaav0H
ZFSoXtjahSdzRbqddglcGVHhLEGU8Q8iVrOKUn8yNxbnZmy9Tp3YcDacW4s3xjhj
EHcC207p7dSIiXf7Wkk1o/JBPsOsf6GCyQITjBCcsxlJZnncdsgRibrR2ae254ZH
7vDiRqI90q4dizfrh5CwTtd+Yj7TNqV88qZ0H3wHqrzRmpb5yqkfJDG8R67Jinkt
fE3ZpW+tFg06j5/zj0TuzUpYv7xfTIn3RLy6HsKznbbs5IFaIPMrdJQ7CjwRseUv
R9ytRnpPrV8ADSGWIufHfCf6jAUdXXsGrrOMr27gHlVyDVYjef1ZGnvkcHvBZpWJ
LLkC5fFxmBs73nOGpaON5n3INzkkGFxLQs8Kwt/woHcDNh5gmYX+XLXz7rWqtqBi
8QHw/5J/k8NFV2+j2QTFP5YYfvzFsNKhGhyItg9G2ziVMwHx7/tCvUY8hrG2YnU2
bYtqOCO5RxMTo++4Py6HIdd6KP++t7sbYxWIS5eAr1r+wnV5MEIkZebtquHp7CPm
w8sDmAfAdjJUfRYXexmJgqVsL7ErCTAp3YuPF/xL0ChXH/9+v4COcmEXel0O6vot
Op212TdFAdAYMnUM78WOLWDLKHDd+oW7OMqdL4TowVlbZMN9CW7PBgFeqg893KJe
gI9S/iDqWuV+8QZEQyTihEBJe9lS2OZdTDQ9VRLvmNA5/Utg874erR3cIllqWBJw
Jd4Ts6bm3u1s/mQIan2QhavG4pOrq0rI/9B6L6XsWT8P7SHiIHaAlRdm1ISntIMR
5P1Gq80/tAZpVXTotnFHI7lyo+OAyfLTvwB5yL6ab89UMcGfH/qxX9z6lb32WM+E
ODFuyrwwjdE5B+j+w3BBTZjRec84F66z138f6xLc51JRy421O2NGutkIMLzngX7i
JV5sCsvqz/VT/FrvsXbGafaIq1JPWvyzqmZN6kLSvjzixHxobHtLKCRUfcMnSOrU
IytI6DEBUAu1AgsmKyPbaLlreCbzKLs9bqUXrQzXYjFnmUgZjwx5Ye8JHD0Gm+lX
xIMJ4mnbefzcm+zd0Afyx0P2OaXPSDO73PJyF7c5X7C3uFREico4dD8XJ5tLKtwN
nlISSdnRiaiWBJG1DSSKgXlldEwfrGz8+hsACFt+TQ8NK+8fI28OFeClnC/vY4kj
XB4MiA0Y5U2XXJeSlo/ZIjqxJGtdlbeoOuXU+lpiJoRlR1PoCb8aJlg3N7XWd8l1
PrDEHjWXZ2JxLADoiwzKo2yp1iIPy7te+6sUWfoQVUyt/xOjhwWTVZ3/W1pxunRi
jnVB/J/DbZHisX8J1YXO6gxKYioUubZeG5rP8a0HDu/JaquSI2sGZN07Ar6ABhNh
/+CY21T1/JBm4RFWhq759HfWd6eNj3YwwT/7FuhfiNUMaiavwkFCQ0K3TqlQbFT6
cgaAXunNC/C3lN7Hz2+59TWeWkbKRXwKO8CYB57PQLVforhdunYGVohefX6GbHxW
EZ2lCAl09p6grMZIiagzHaQa4VYa/Rv2XtNUnrT0THkPRFcRPBVOX7vIlkBKNNDU
7RYqGjErOp+viAR480zpDN+m7D6fu+SWz6sOpK/pFO+fKsH4bK3KKL565avLlnhM
3FP3xb1kvv+V/imt0Cb9oLJTroCBtHphTtbYCCCLXusxBDm89nRvu/l1nD+PF/1A
UQOV4u5C33PpaUW7BX9MGsk0ivhC7RoIDAnvIoHmrAExBrI3sTBZvl7hPQLqToPz
PsPGR58SGLCJzdqxG0UemY5l67M3QjFmRpSk7lBOV4KcodtlVOB+kyulgigT4sMZ
pCAlQXJBa3Hmck4fxcaM031uabiXS/sth+JgeaQeEmqifIu96tt5JKDpf3zxKAPX
lhqKKbUSflDda68h6rwWseS4mL2G9zu59FlvoboNZzG9Utdd2r6t7EQIuVdojDFF
CIjwd/G0Lzrz2zz5p3M6ib6PltexoICGPT7A25Im3PaE5UxG+7enxFY2LzW3kVNH
ZJJg80aj/h1N0ad1XD4irJado5/7YXV+Ll5LrxIQA6MCqjpA6k5Wv3evW7syykU9
JMOU5n+RN0adIxM1zPo43yo6AW93XblxyrG5M77+q8JAsc+rC3Pj+hvcURSQfxsS
auTrFaZD+iArMLBpty93VKKyfk7NAb4l94IpD0zsCOrqi0nnS/VIb1c9XQkF7FxV
TQ8Mbf6dlPRzsS1vdwj/kPLNVnCceXksasH2L+lJ0yWiB4Y2mcW/Yl/rs3lH5nTt
zdED9Oz9wxzik3qBLrg6lgXJnBZ82th3sD36GU9GzBs7lbg5BfPp4zYs/67eoJ2g
ecXvv+myHOD4HeZPxDqiRVr2UFgOUID5SkTTUdrOu3VIOjh5c32qZ6BZiN7g1DWH
eljd1bk01x8MzKVyJ2TxBwgJRK0C9yj/DkEbSrgDKPgRnJdkAOw3gl7KY9cfWaF1
4ISCEJTayTFk+UbkG6xEPrSGghn2XGmDk+vgKNyhxu1YgodtzfUB9Qpnoqg/WL4B
QKdwhS9TdxgVHmmJv0l42rUL95+o+2eSAZP09aPIJ1DByV7A2QpyCIvQgtENKwmM
Ajiw4RFoVBNUjXh0Ier/Ay9HwyWBI2BQLHYDcdK0AKK8/VgJbpvHt1nBp0N+TchB
xlNdx+dlTtsi5zGq6lAUEEHtpljD1jfzvcbbij2Pk4VTztjF61oEl7OMT/d9uGja
zzspBVtfGRdmi/Gh6HIvkN4zhdpfj4+7LwwrffMHEDkEpt5r2cdAk2VMwvUZUhJo
NmOIUr89+xZDaP3IBQCryqOhV5iw1L7w1ahVYffDlw2U2mzkDIc5q3cjqWUH7iEW
efIuo9mXWGN4FzYcPlL/3Olo/MQLPIRYI0/b81TaADacr2gg2JFiTKafeS0TrNxj
/aT5/UDp+2Z5Aj+IiRePhXVlx0c4ZpWEOiCtMyhoGdywxBsG8ZpsY8C7hgTqfP+7
V9zB/XPRZOsgs5lM6bS7oNupa2iF+hig8ZBaU9MjCxRe9dfoM21ViibuItK+51v9
yu9joe2Ao/48xujmCYsxWMIG2v9fFuzCwY4TbVnDBKuLfEsaqVLJSN5Rms+o2tsm
cK1DtMIAABehs1zNBIiC4trnk1wmPz98wKHG2N2nFK4Gf1TsjiLGvrb9GUWinE6m
jG46qK5h9ICk/h3qHsWNyJLNi6Wq0MBa18UhweR/ddmMAWSqfFqRmGT7GPkIu7TB
n37c26bAz33Zk6PEIy7kYJvXwL2wkBHOPfrazQFETrke+6w05dtFwGkXoQwGWjvg
/BB1YStjPWQfmv3eUEKTNKQ4OCRXUz0IEAj0V6jzQHDzlbFTnTsJmEW7B0ptoYPR
QD00yiRRZb2cLclaaXiTpFLk+5OQetMlst7i4XIM4xJNjf/iuakM2+x8mXy3lPTu
0LLvGc78BvNZ4xWbNZ+5QnmcMi/vnw4m918KZqfrkpjTP9Pq/6upRybrl8lF5mIG
ggNj2KjG2gJy/9AEkHH2bCgGh6INdIuQlZ7IU0UtcFERbGpOmQO5wKkv0UWDDgGR
qoOnk2WOoiYTslvZuER4vFN+ZervTnmIe9Mmyh7EE5qCfqJOxcemXJw8y8toNQH+
KP0mw8sKKPjvAqRF+ba7n7V1vB3O4gwjtJaf1SJTsUqChy6a+jTDS3p1XGz2vdr7
ZLYOYXXA0teRICMq8pjl5MSEIgyRlhLpsONMxXZd31MjFaQhCUWLZvZO9sC10to6
3+2VdbrjtrV+hI8Qk6wf/rR7dLnIvI5QYcE8M4Z20kvPTbPkqeAvecG6UvtC0hBd
FtiFEzxGJLSrxrUFf8jv177jiQPTd9yppo/WKC6lQI9/Hs7VzLodDYJxWPTol+Pf
peRv39m0shTSBES3I/nW1IUCKEZz7+p+hj46Vt4PoZGDd9f/LLiLmFp2Wm3b7bCg
ULS0Z+ComlI4+BRab9BoLWQjiqi6esDqFOW7Xdg1m2coBeXSxsYxNcqH7A2wS7iw
GTehRx+OK7smmf9d6fO1KUgt+hN7xOm3EkI2OfI4BpoTQsLYR9BJ1Fj6j4x0/rMy
DoY6QpUOlmcwNnpLp7H3QXx3z1OXVdCn2Benaw0WMO+da7QmTsjjWHSbMrIBkOLh
4yKOufAnseFSknMnbtVL5agLPOAE90bEaA6gMavi+SFfMxLSVJJVQWtbrSQK8zbY
wWDSQoL7lZhjlk2HodeVg2x1OOni04ea1PbZFn4lIOHhmnGxlF+hdjjGQD7aCp1X
Amk4Fg5ABxfAqCbah75ehK2lZ2UvvUuXLP8X4Rb8CgSEw9Sbw0nDvt2Qo9OAHeRI
0V20ErRyOZhUhyXFZulNtzxodGxL5dYhwCxgxR44EGoNkw49Ecz+oIbiJb1TWrZk
pidHSK46KuzX/9+x7FaDXUw0++MSz4ClYN2Fu/m/MNvoIL/fxMKVeT23S5KbQWzm
8MAiWAluEbsGF51YxUJJCqLgUk6k2l0Jx/c65emBorH+c4Ud5FA7Vec76KlIiLB6
vUPYBOueoBuyuMHYnDjG+P7U4Y+TZRyOXaTR10Wrj6DokLfNWUBu8nPsxsdsdEE1
xUqYewUjuKgftDi1df91HZvozsa4sEK9YNrcN+YE+tKE/T/GWGht7qzOE+0dAkEN
ryrKggwb/61efhUYvtg3lA26gjswGVWhmFoUZWcCa3p2nloddohKfDs3YNAgEP0K
5dfnuCD9eE4d7S0ypNDzLlKzKiK2FzLBHUmf768ewSt50SNNtZLX1BdU74YaUUD+
d+kWgrJEiUZc8RCt5qJgTDmvisp0dtCV4/tWzcEPl3olj9+tYZTl9McRDcYXEPGY
I7lW5DKk6Z2iCtzORl4fU3JG2ecPmkbn8ocb1ONxqUV6uAUCwGoyIYpLFV8YwZso
gdbCGjhd4NoHgfVIMKF80+LH0jF0Ix5Asi9mFL6a+F05HXFR83GiqxR2oE2svQNf
1tYA3lmyLk0FFTOecW4h5KefzH72Ugv/RlbovI/TjvKZUCmyJ0cOU0lIuW4Yec74
vpWJzmj/5pagFUhhP4Pxe+jl7Xdk8A2xcrcIlt72P3JtcdNrdO5RN9PbipGnTJ06
5g/JFa9NdvdRhEl5ZGGdE+THLqKQI6aH0mzVRo8sZlrPAsRaPDsTnu7GWYQf3xeS
+ApFmU1ls5oR3OXNpD8hhg+sQdeIDsiHGaMZYlxhs6IJ4dCZdNEKWvG1AKwMDEWn
jzauvJwlUvtZxm5ZblHbCdYF4rDQBWYGSGPaaeUlbV2Zgr7FNFPy+vCvPoRnZBHq
skn+P3eZTzYxxg4m0GQzKP3YIuvdaAIO4xFRiZXuzQeGYPYnGHNTUkniO15Rd5pZ
UTD3kWd/gOz7oKjtuuurfqGTnMFSTRd40+m8PgPiv0DKmG/COGrepHONE1+5QNiB
jCJu51UmU5UzPOd2pRKLSLdMz4JN4NTE7AFGlraVgOdOObhp78DATjwFPTPDSB8B
zmFqzzT9+LeMjG5Y/CLGWp+R8sHb1LUcfv74c3WBo/MNkMIIvwIp+iCLhOb7+HSL
hJP+cOxgGqZZVcML8FW4kANci8SxOmgEJiAw3zFuYl0lCdYA8jeHDkTZFUCdlrVQ
5xPisVC/JhHdq+QK+G1tSxd0Kq3cxiGuAhAoTOQM71RBUt/rZ0+st9vK2dxmO16g
a7/32BoKZbRmLNFxkNHIA1uZQC28urRhjv2tpFzWwumKZc2TNppz3lTv3ZPWb7wn
qFgq1LKirIzTYfUqY9wLRt/AsfaoY9R+Ees0Rb+1dTDj//s1eoNcR0m1VgvXNf5I
K9MCTQtdNZLYkLgu8YTfpUpv0HnFEd75xK4GhIzdWSZKIyxLslAPXTmmGFTdai6H
MC8edBMZiKmUdh6Efl+WTAnTSVOmO61Sv7QQnKKAqWJ0NN8bh/OYEgHSVgBUs6ft
PBITbV1PlqmSMdt9krmpSPY42FVsgMq9FB6ZHxvTzauJF1KlEM8HT5tIaFVBYjf+
f75a1W3hX06j2m//Jf2o2Dpd+g7Hob7uSBJa0KYWp8/CIjDwFSUprRaBz43UwIqN
fI4WaXfKaxt0m7TUv8YKJvPsjVXUsx0qQPVszWCnkDABd5tPt15nd/+WygSTlpxF
o76ifbzVXu26maPhvEOuTMfep0fsSwsqjV7G/IwSBAvmnVXIzFchHM0STnWxF2ND
I88XUmoyxsdtytu68t1fO9CHdrOGtm6Pzr+PDuuIzG+GJODkeeAO7O1TNRsqvolj
yvOsnQRmbYujEQFPGzw8S9qyd/UWsTJ+04eF08XfFXZGoTaPFRkpD6TI1+Gen5M5
LO1zVIVDhHi58hOFbTHs9MJACkyI2Jy/uK/KH0+KXqLTlIc4o12I6UYLNxiaVWJS
HH6OO+lJTeVuPIKn1se8ONLPkXroqQ96KvTxNTEcXwwrnGYM63KVxm9F8716UXYI
a38Sc4R/0JiQWesFh39NcDvonoke29JiECxo9VJxhk0G6R7HdqDNlbwkE84Ewsdf
T3kaMAQjH2+xMSngiMD+LIQFEGZ+DXFsSiOFBxVmM0MVVpMy0ZVFxjeDnppLMnIH
9fvSEL666WY1qhu69O7Js7kbYhAVGncWcz+9fd5Q01uKP0so5hAccomU3KZrdS5F
P5Z60CXEgkmPVhSibQ5828nVPzlBRKCP1Px0NKKMX1/RcPMpJQJPSJXujpdbr2BN
rP5nwxD5TampyOYdnH17dtdWW1UAi/s54GQH+0C5IEWWdNf6UN5fQF5Voocyooce
aCb84hyVeC7Cwrl1Jpfz/ZoveE1KR2mh9J4aGHQZ9fOTxuf9yXpcDCSmBgcvVbwN
xQiODTkBF0B+YiWTl/7L0C5eS+mirxxuo+Lk4vw1oGO74f5MwJd0lyQJnDcEnYcw
/qvaM+o+j9LBOcFLAtlJk32JvfKOB68erTzi5fK3eADh75dJ9ZH//eF0hsd0lCbL
buHOszoOdI3UA9nj1xZv3/AsDm+wuxo7FsoYsFVXQN866YX+ekt5BkvMzSIT83hB
cJa46e+lLoM3n/uAhIfqZdpsZregsGa/1ewzQA6it2wtbKuN11LktZjOoYMBM0iG
JeJXDRMBFG3OLjFHoFdcS8L0IOLHX2bi4ytt7SY1U7pd4pu09TlwPTpgQOMFlv9Q
Zo9H+TfhTffwXeMEQrqAeI2QJit1K8ULn2bcgZ+Rwk3oJT1HjuF1Mqkjco5HGmzk
SmLE65DkoK/dLNkcN0JWusLUYxiQK28M8ZrdahOZFRZHPcLk5998/xBkrN+0jOvj
ABJXYlG13/CDBTFj+H4OQhg4cXV7hDVdtgPWlr7b/61HLkpW1bpCifCNKOB4anC0
Kq4s479cK+qAWH/506T46zHWZmCLrI/Wn3ZJkJQvFJugOrVXOX8Lk1xZWfBFhyiY
tC86ZQrA7fEDLBnmZwwjOOg7JFwmy2JW0hYTB3HhudlUCWwHhFm+pWisv10c62pt
fqzuQTrPp9+8ewEXSXIAWn6fGS3fcDgLGc7yla8XWAXTnd8h2fjsUouKwpkIGLEs
yMvasOiIUEsf/ykBiPJjvy1lYShdtMCIAV0zjiNhKErSFE71t7FUOUUEy/5mbEWs
H/aznYxGh3979tyI+lDhP6IhbqZPiLVEj1OA8NZsgODSHgeE9W7V0M6Ok4KeWX8G
Ucknz8jWreXTwA1Ltd0BC3LjyLINIhqLG7LMRy7uuebCX/Exs9BA5hwuS3qf1NVg
Z0q+SZ2mbrRW/vqDGHaW5uk1EkKBhYH6a3lXF3M5HqwBPKtO2oI5p806srOpWU4T
VwK0gvuG6lzgulDNIDMuU4154rtBFQPh3m4RhNCSUhMthD42jQC+tSgnh+LWS9eF
Nah5oZdtdR/I2kTpIei/FrWqVMW3qMQisf2zC2v9Q2wYBRZ5B3AxTki5Mu374s7p
ZljVNSIjjeBiI73ZXKOCvfIu227duqVyRyqrwKhPi5oJEoMeafCs3uz6vB+UW3sL
f4bRb4Egy696sMNbnAfdBPDhju5l+LMNX1YuxZy2lyawule0qyDzqDzcOctdqhHr
vYunM9HR38lsg+zz4utLla7RpOioJhH86OIUAUUoZ7ESiAmuqIqEKtxZO/SWPnUw
tyezLcQ089758qlfilHnI45PTxUVD1CJ7Q77+RIgYjpWBX0saqdUBwhRozQ3mj0t
reO/ezm6brlIBWfB5ICvloMmZh1kibK7XFaxzvXYS58rXJjH1w18HdkAftcqsM7L
IVltFyjQDmU97MK+KfB3KkilT7Qe157EV3Cqq4YP31JG8YOSGE0PoIklcjJ3NC0H
xKQxtBe5Xd2XqwTnq4fAQIggz+d6mZA5cunlUzOpfbsHqwHPTOS6YMbfC65GEHBm
37Ov/NUidSwg4FHDydCwMNpZthb8av+yrHgXnAX+CdClgTJj4+BqRAfgPO+CjgXM
pjzDtPJ6Lo5TIFhDOzPGD9Vj3n+fBpdsEV6g8gg/IX48qX0+l9C6z8pSvdZXGqMV
lwrd4WkZ0Z/9Nr7jNAt7BauNMfZp+TTU6uK4EJC9CtypaLYBzQTYU+IJ7YjrhHDI
K/EJKhN6eCQ8/ua4ms/rNpHouI7LmxUpQ87VIpF1seLIbwc31UcYZb86KgeaMyUP
8u3TSCe2y9tuYvTHL/I6R1aaqBm9RJ1e1n5in+ziuaf9KFH/qFL6pgyYROpsqiCY
/h7ITMmwa9LDGF8dY8qQq7qpAOrfrb502f+QTx3JU1T+tZzuwfyA8KNKgwUl8957
d6YUD/FD+6A82y0siXFI4WileUtYD1ifF0EiV4ee5L4FoMbE8mip3QKG+ynK+SOs
DQk0LdRXYZhq9l2AmT2TPuDCIDcBfamo3LUWvE9UBUusgHNG8SHmTye4tm51RrkS
l+9cGXpiQjP9C9fwuTND1FA78J1mXFd0quvw66dc3wvLmrMZY0nFcHj7rcdYYoaY
KijCIszo8BVsOaG7K/5zACAHuW6fwoSoYolvJOTsZg/ZdQXjWlfuEv5TVO33eaQL
IyukWQOfUHXB9OBOeALOr0pXyMxnNUCC6DXeKhYcTpkB6LcRl0quRiwTOxSCkYvM
1Vl/KLyImEMaurgukY0GEb/EaO9CmQVLg1A5iawEI6K+I+g/0+11b647v0YLqEjT
4CXGysjTnaEhA3LnsspiQYy3kljov5b1Ce4pUPCfAHUGNIu6lzHrPjQWYxMi1/lc
lfzLurvxF0dgJBP79XsL6NleenJ9SUwX8Yh8REmi/MOag7M7+M7NvO5h0pEolTN3
bOD1vbC1rOGhDtzHouuKA+dXFkT8ryRui+RGHeuSrzLEYD2KHKUB4e/MEEx4GC+O
zAeEXmfU3JD1WjqSQ8J7g1RMZ8MXcl2iue7o/G34X9Ki8UJzdUUH8GM7sbrtxPHo
RH3D8sAJF7H+PwYx8asKwNsqpvaWYJTbrWJ7bRAniUBkEinFBWaxnnXWl3TEqNs+
xa2N7Cxu5HRQtFnNAc/O8U/bLnJEc6GScGmKAyftUJ4oVEqlcpEh1hY1zC8E9RVa
W+PCEv4o4eyx9o5vMfADZsNiun3cA7Nt6mSb+9sOIgcc9w/YUqe2hX9OLzbY7lTd
ikxiMdrAmejTM2Hv96fXLs6Q8/A839AJGbQU+tfXzyglTX8e3787JVzI2Y+/ImZi
KSAjKN7j+Prv3EGytA8DA80nwXhOIPgO5NrFwyn6CGS0i6fNM7BM7d8dCBV+/4oI
LltlC2lk/l5OETaNardWXlv3pH5lEddirs3MwJPlI5ZeeBETTZJZlTZIzdDve2fF
1UO2ICqDi4yTuvDxGzMmIYR154P8mI+2RYZWhpq6SYLIJox0bhdktIwPQ+8h4W+G
bpozmo3IRV6vQVy5TWpY9xa8JrprV/AqvRZC5uIQIJboiGRue3pHPALBLj8H3lPW
IJnetRGzWs2ZcrHeTELuzt60pEqrFKHZ4iAdcyPRtdtV7/oRizn3B9/rkX3qy4rW
zz9p0w0hTEvndxpkJuheolzx2IvRQJHC6SibCA4ZoJfDmmeR9ITpghpoZu8K74fN
gtOFzJYqPag+0qd5vpDSOWP0tJnPWi+faQlyZ0clkbPFJjzsjCrYxgbdv6ykfU+0
p+qc/ANWGSkNEWQKIpjac3Jk9188tjIsZnMhg62Qfdn+tHKN/KpWUPv1r05xUXo7
OUfafnY2s1ZWtx8qOYuAGGvOif8Jqq2VuRwNEoYTn0sZwY/O/9xERSxDWV89S8yj
wSGNr/VTYaVy3mGx59ZQxKGNUjVWBDbrcJMPjtnAF+MXDawDGa/FiI8AR+f0j0gE
tx0yB9pg0OT5Q5ci1mHpc0fOzhQBNsGIZ+9Tirk7DkOZJ1rg53+zVarNtBVqHivT
S+LCy2c/sIGu3OSy1Pn43tGQ4ws55v3TBKI1dWy1zY2Cxf6Eoai7inApv/1mvh+n
X4W1Wp73gdJ8d4gJ1H0KSxy+wxb4iOI9i5e5wkMmZ3E6vVFr2UkyVx9kPM5mqEZ9
7OmFym1ffp2X1zymKQaX2lrDxgCAbPpmYTNP7JiDcEDzDh/P0lDH9pYvZJ3gihJC
nRFGpGKojW0hJnQNLNz7UEIwRsxjWNPbHWHTB6/MAO3TllNy0115F2gx9bbqpnuZ
2WuUdqFlTPz8z4FdQrdMTuj+EX8JG71tIX0U6vdkH9VghV67fFAB5Yy1NlVcCga6
GsoVCfbFtpV+ZXVKRcoPLrmtDrUDK8iiB/LX2z3kvo9tGwtMxUldYXescbWEPZgh
CqeGHFP9ZOC12pIXflUmppc9HDeXogT+HdXKOO93Q4HFncaqN10ErIl29IK9iEvF
lVQc7AlQ112eUvIf7+6wG6UWB8LsBaii2QU8vgKo/W/Akfo1a20GF+lB7alPv0WU
rdiDZ+mToARdbIVuulXvHJbpE7fPumLchDPa87AdZ7g0AOUcWKMPxUA563nXoqzl
Asks6iHJIoWFeISN6tQxuOR1HYPo/mKl880aDbXwUJHCPx9Y1vMb65gFvkLJcD+m
wJyutDrbOV3Tm5YyNTwm9Rowgu71245IgrISc5FnBcFnbqdSGf6CMfkpgrrtPIbN
9b5DANCUv0kfi2uOPEt259MGLHXyqK90k62ggQd5pGw3Df1a6jhJuL79ZZ6O838m
zZK7BIKeZHanOyZvKq0UBoy4eEzQGvcIKBpniG6YySUKu+UPDIkwulTksZP5jmY9
Wx+EQgAL9sl0E6Yp/Y8NhEr2a5cP6cNQOeFBJ+FIiGnCZCvW4ZkggqQbrCWoDgqG
nptejNah+d3UaJcYIwMncE3gPFp2+sYZGHhZeGoc3Hv2vaX2eLqmyKHmXtKw8/Sl
weCMCeyQdSGC5N3+ZDnTE4ha48IAvQPYsT8uxrd6n8NhAS+rowsCp4ASwbK4oA3P
zP0NGrGAJqWwJbss6aaR1avhJALWbVeQUGlFB8AAb/4W21xtVuZ91jephBDr302M
gFzOw7WsQtPMg9niQI6oMst4vzuCMxIG4s+vxibeB2Kfj0M5CRtb/h2oHstxtPU3
ySPdfvRQDnuYz2NXUHe5uL/4CHKZ7bkVrDuZLOTIgPiRBZ7LfNwnLosNNgGyCnHS
+LO6LN267x3p+3srztaP7xW2GG7TFXNx/0CdTPlOHgQFb+Boa+60H4K8/cNi6B7s
olJ4RrATxuvvpy6AGvbkiZN3CbYxszS1Befacslms9THJUj0Mv3cayf6LgOECQUG
nDcXOpNnMJumdL9vaPQNWUMh13hduVMQ7YacVdmg7Fr7IurL4MGdrKh3OPKJ4aw5
KcBeBZi/muz03yMmcQKfb9VHw1ihQifYny6k2rVQSGgrk6/FRDTgy7zdbRJe6m3N
86DJYyN9p66yOtDNZkYOq/Ybjve9XQ1kSHH/X3oMiX3Fm1FzzYEriSAgZUKsOZKa
wc+zSnqKPsbDumsyaXo0pG8CWoSYQCwn2gDuhPOee+HGK+jyPbmSULRxQmBSqRfr
8A0/ApIue2Z+mC5rQiwyLEF2dE89zXey9JfTQwqn9VkNqwmY6LnZ53JzJ93qEwAp
D/FbvkgNQEvHYH5jhBkhdVE9UUx+CuMDQjIxjURz159lIFAF08sGGxD3ib4jXfhR
3pUbY+8t0mBm67WCSF8O6RAgWpKgN0uQofizEZ64Gtp/HaityjDZji6p3vNb5W6W
zMmgLMPf7/eTNpJPpvD4dqeW1Ks0h+Xr73G8amXQ7yENzk59avZf1ohj5ejv7Ent
ON9b/WudWZAtscwZCmLlvTrHwobANn5efcn8fui+0SMatRv0yv0OzBEqdo2NVgwN
98OWo/YGMUj0rmoFz8u2/1v5OOVRvvrwQ8QHwPczf0vf5lEb39fVQBuAGLfKhlNp
Fpl3aqYvXXUy6QgF/3aKjr6CYIcdQSeHONYUHQ4E7e3/eOtcJvKqCkXu3kwGKLxr
1h4sWMGQb4aZcPJZGDnp5N2HoNKrpkjtwVIJsFS8yTUGpbxLI6JQtKLUSMsw/5hg
siBd0FfFi9hJ1uwEW8yTndXS86KP6NNSykV52PkgmXonP9OrvkjwKae3iQQnA+tD
bvRgml5Hj2IHAFxeMSzWYQZq3iq02zEsSalDGLXl5UE0u3xnbhEDMeaUGzOdxhAQ
nmi3N+hA1+4JWcjeIe3AIqIom0Mlnam6VsFpcb43DOjkNaR+hX221a5MDw7u5leO
HwVZwKpekiZotBqG1TXX3nIudzqfRgmkUzV1TIGRzcCnBX3zGBG0uvDP4LHMbmOw
T6zfwGFvIfi5dQRGK/u58r49nQnrCfEmbnl9aw/CtF16YaYK8Wsmww0ZKHD1ilaO
iRCuOmswY6ZqSinluiPqP+DU5AUQcdKuYnpYQuVZeEdyGmcMfF5PLXHacCtMJVga
F19977CBM7pC2qo5AgiYRWBSuOg6X0aJuTH797hr+RFvSNJERzGeJh3rlOv83CpR
P63Uap3vE+oPzTatDZcvgHkZR/UiLdLFw6yLACuWQs+GqgszLWfTBug0+99ikjdx
Nb4laCHcG0lxPP4dJpPorDucidpOdFCZonx7W7EDahbvmPr97xvLR9+rZHniOgBe
RzqeUizqW3v7DmTirDr5QXtp8iTI8WWOjHUdUBEy6ypxvM3NwyB1nw0r6PCSzIa2
CB0bmjx7euurImGMIzT1f1ZQOeTmTRePNnEGp9+XPlVRNMKxQGNbZ0RbJX/t+1jT
Kr44JNtM5Xk3iIXRTmjIAoVN0EaEk0lVL/JVD4zrNhZhexj+cXVUPhqf8ACLZiHy
PmeEkigvwIRnLWozSCPFhjhZeaYBXnd+95/jNs+rNzqC3D+KuA4RMgVJOc74DXMB
/ZMREAPo5YFmGLG/p1B99mY9Ox8sOaMER6UpB7LOveU8NP5UKXgnGhPMqswz4lPx
V08BZUCn0ZGa+IpEgp2Xydnrcn10ssXeeFGyhmOao9fC+TISmuILYAYgU8DEs3nq
jkJ55LcI2FlRN9xwizv2zN8/6sSYFW28V1JdmxLRegFfLMyN5sV9yPCJ9Amr2hyl
7XtDNA/C2/xq/ITbjmBOBM8JD3wXBf2+sfpZU5VTU1cKU+IqbpGKbbu+L8/epE4g
H4l/DUnuE/izVbO2qC1E/BZdAeFqA8uu01kHQLEtHKbrs3iWzHhVjd4MjCe/hx0b
IUk9n1oczB0MY3PYVlJuQGWAUKYQg18lYkALqLPxN+bfcmen0GCDe2geWj+z/tDR
4NMXQkbuLwChWADsnbS2HgS7Ng3Ol21OAv2d9E+WrnPcJwkeho9Pw3tklrNVH7W/
z9fY7CDyPnc7oXqvCeBQDXJkNlXG5mf83hI8vPuDwOFF0x6wVMFXCkMrelJeWfOu
09nI2sDC7bn1ebA53VaRSdhepW8zQ7OvP9YaI2c5yxCoxkNIapViLiW/Zmm4XeQP
AV3ffu18/5F98ip7QKgZtuOzgkfhrtRWeqlqqg7fMDiCt13tHchUD+Iyrk+rwmRz
lUJd85VKc7+hsfztUHBToUvYbKhNOmOMKvAbMZe9SPGlTrXQqRm9QMj/qU/yfzAC
i3EJzR/pVtYvlr2hEe9CzMYdvYyAn8cLt2/m0sGGrHTe4eWywzXcy3fM8ZlPIbiV
xrcw+ebaNGJPE6UgpV/G/AI7tijJcn1eWhNlOivxzxkVebfHXd5Wr3/i5CI7GXML
QspVy/o/i6cGq5DTLXErvE+iN8JW821y1CAFH3s+JSxvRXhH1CEhMteCV9aKDbnT
5oz1O77/VV9Q1fWXbOlVuYEeW1wvbhERgF57LfOLhAuxNY8rlu41EbmgyPsuQKg9
+gnex2VMsofUv+nB2UcQn052rg+r7kH+VTEuRNZJJ2VRhN5JUQUodOB43vKhkFL/
yJkwiZYEfChjMYkbGT49ZEojQDPf6w8NckMO2tLKBiCtTuXn8/MNB7aK1Y5+1+if
RAWZgWk9uIVa8sB11N83+uoVZOhbDaIQ/OwhoGhPrkQCb/Oqi6J1QGGd65K/Iq4A
eBEPywyThKoNF/U5GCDK3X03/a1Mt6pC+oEoJtMfndp+YSFT1m8VdKHCmEeR5ERP
iMpL42F6VjKUXfh7GpeXFu6QPVV+mrL6zFcu9oUDB6jI4k3YtvTCuAeETBr3MioU
mSfGuy+A06NWv4xUC+f9QDG///skN37HUP4+f7Ew5SajAeLh1QYCvxSlMHzsbngl
A1nJcAcxwd4Zhn2lJsNm4dQTiPlxp4RvUrRnaD6GYosjIoq9OepRpiN9Q4nuPA8f
8+TJ6mYT65kEc9PnJq7rRFGxwbrxmB6vzN//iwEoPIo6N4OzK0Y1A4U0H6l7T3iX
JN2/gXA4+rVmkDdXL2ywPsZuOGD8lrdAmv7AFqkGsHNbPnRFIh8Cq/Wr1JhcU/Z/
JxADHUxegeG9Sx+8b7cpg9liGVBJFHNMZaTkBaGTn8WcnBx4SFKfHUfj3DlBJRsW
5es+F3I/yAmLhE+YU/nhfsuhUa1wdZ+Bhn0h2Yf2faD2I/me9ztJqtnuZS/7m1Ti
CTLpkeC17tBQ77L9fUSZHgweHFhK+BN62UvfbcYPTWf32bR2wiYGpifvdZ6Eu4OB
/kMQdnydlJjpcmiw/iZkR0p+MVW6TaqXzW+sEOkHQkjGG8Gsrd8G1PsTAdwqRIwv
7qSMfbBFvawgVnxMhGrawMHXGJnPlDFaj0ySpXfpUZYv/LGtmCFvc/bYFegn9P8U
ObClwFpWFmOMZx7Porcvncckz5j6OT1nJYb1rrBhWIbAx5rAA44wgEyAGlJy+u4G
XeH5rq28uhCAfWOdLE7jM4S8Vjj3kCmI8XnhP9pNEseIhVpLIwe44CBXKTmpwVpt
D4KcH5A77fhys97bfXTFUrB8Wqfm5nj6kTfckjXgQLt2XymNXXjUfaG9glScvWen
BDXRI27G8MxOxsrCA87NiMWo6ju2eXuRY9i5HPsdFLUj8pNjQbMsfa7DP5T98Y50
cjbAFk4+tUJtw3hqd4HJdHxXPY4pDmoGNcqlgJgbQ23gEIf/TxptWN2UFCBQC324
3EbZWPo/SMx4JoFVtbqmIEFqCT29OVkPA6+ZT3Ho6Q2MNNZ57ADSbh5wD5FJeFji
R3MqH1v+0ovtyOI9/Wp2Q4Sp0V5yGndkJQq1cct9b1iuTFw+4/omO/0IwAsd8oS/
OevMTz69KQb98BbYxA/vdtMobuZ8TmgpNcl13GKucbzwmv3yTZLJI0GnZkQfmzMm
tRD6Mzd84pESiDmgGKCayJiEPEyAPRV+DgKIQBNhZk9ifj+FCiHDT953s1MNc528
lWkpByfvm8PAoaDRlRirE5l7UJN3/FZYyExE4SPxEZBzTSZa/X3xD++BVBVkiIvP
NzLqnbQc4nFoEdrDj0tlArQ/+OWfL+0cbM5z/7IC3oC5Scu12bqTo0EuMbgQMTme
1yXZfFHOa2W3Ui3ic8nXZb2UqUyQmJOBGxOi6SWeoBS7t9Vvjvbp+9jxS8JB1pg6
ERmsDEhTrS9zLPIvOJ196nnKraIB26FkuojKagzbUCWUa6c5/vl8yxaF0WxGZtcW
vXCoJPIq6hBuQw7hldVIJXLMZ2DG2swOh4OSX/TznJ1HIUvmr4qc487sm94UkGGB
dzP73YkcC90EU9k7c6MhNM8kfKgn1HKLmsJ4CwnP7ZVgYrPMMV+R0O91st3IXAVW
PJfWs0VHQu9TtweC9fFWsb3WbcEAIz2kHBgHUjWIalDhBZL2RFANqcidiEWKrhSm
TUcnQpPSgv/rwc9fDLgByqH6xpY7V8STYWqi3rellZA2DUMV6yZKM7C9ZFG8L17V
nWfhji7cMVEur/ojxCzxt/RgUkNpofmhfZBSB8Zcw7sSydZCX6UFKu82+TomtTzP
T1bkxSW0sgBQXT4RJhk22RmzsPnL7X48/7YZhjoXUxDgNnq7nH0KxtWp10eHsFd2
yXbYdkQsA6MWHfR2iD3X/7ISSxgS8Sr/SuIuxBvvvf3R+/iT1hT2jJDCZYDjdMw6
L8mvFh+e35RMn91FD3NNlsQWqT/X5m81dJn9Lo+BwpQYD5EVLY0h/XdAGjt00pUw
90MDrs3iq/T9RJDMMR01oCCN94tDlAWywK8B5BAo5WBbrubx/GM/JpIhXbwUVng+
q8lsxTXTSdKA3/Hmg2K3HqOe4WXM+jmwqKRU17NRaw38jJhPswuSVoDbiedVtGCW
8tVKI5sSdMRtv9mU/FryM20CXoL28Ae60vtjcHaE8SowRcxIXkjjyQ1eNv3VaZKl
+FvmXVUKF4KcQj87RftDu5bYviWV0+3qngii3dcdPAg2vmL5D6ON0D0aKglmzTtQ
KuLJ/TzE6NlzOzUihvYvfdTCKC10Nqw6w994TlD2dygwshgZEfSwrkAx1wui3DI0
aHZ1oJyvpH1MHoRsv8guX+GT5DPNan0iSVHBlllw85y3ZkZzfvfdSCgvCqSl03Ls
KRvdK1x9CbO/6MORMcfKWMrt4BQKVjHhBYi5rLU1IUPxqtifMgfngmureS5ho9Z6
h590y4VjPIZkXV86eRknZNV1MHTwnQRLIkBEpGvRWnMRJlVKeyHBsLa/e1a1N/NI
KviVuoZldMNxw9Dipb9g3j1gy7H5UFTggCHS/zqhaBnHGphnw9X4D8hU2moe1NUN
6pC0z/PZNZmlj1NrjTuLpi65grclbZ7No30n9EpQpr/sSpyox3q2REtSltcBS/NS
kONod52u+JpAZi85aI2AFav1fB5NkQMAE/AabIyE0hkIhJjV0uNZdeDXzFwEDDBG
316dbkgMlzDvmbB0HPx/ca5GU6gwL+LOV7BC1BwXOF5BBz/otxcPtSg0MbKJe0WF
aswsFOD74kppNfk4PgdZPxHzeHF5AHCZzamQVJJ7Qa0u4j7dQqK/lnFuhoMzVOIU
a/FgnWKQUPO3wrUAXGcfL8DFITXgaqVtd1PNPIiFKyPjCtanzjyR3pLMcc0ngE2X
ap9XRYkkAUH6KTzYg9EC5h/pvAxEFcWa2jVuDkRxpk3tE3w5oi5t1OK9R5UUHxUX
QeHLS8/TASSuaXUTz3QTZeZujinUBoFqph2/AMCnEpS2qFEEc6Pa9vxOpTg7xYOo
Iyp1D6Axs4nOS6nXUnL8mbEppH56oGZOZisvWhEXKELmERTHVRlvWTWH51cF+Vqv
LkrxzgVZCo9/RdbhAWcii5M9U0rswsD0folfzmiPx3ZgUoiZw7zh+4LgPHE6FEG5
y8sTKrhOcQndzuIDzQKlXbPfR/Dge3Dv7qfdeU2AcA2yGLRA3iu4M8HzgL+aMGVg
sBYr74d+qVImlb475TtLCr81Puqj1mnG1PLg/GMt8qP4Wsolkqf3AqU48l9roceF
fKuddoFDAvs8ta8cFo12xEnvJKe5uBMp10QW+/S7ntRFRnY0HTIuIPC4piM2j6hG
4sUh48ZDuSTJu9/HEyAkz133Qj3yyHKh5ZJ6p0IX9KAiKlETOHgdTmJo0CI6gIox
a+meaV1LOs+KWKyRNvnaYbjsOxcLr/RjxXoNn8BDxQRPZFxAYRcee2taISPHD341
GVvwsd00drRUdqAu0Y25RTclIqd1Ds1PitWJ9BVdIv75tEWtS3/wHD0YEM7L00Dy
BMjqKMKjG/kVbWMeGxPSQzGbu3b27fUFcx/qpD3fz+SqnYCsPZZQAyUjqXXpQw0u
AhuEuga1g1iToam6Jeqs+SwPS0vxeX0rkp/f0fzHno9Jie5PWXrLPkXlsEHD3Kw8
JYX0X0CM/WkUarGf4CWwRIoLQKN6XQamld5nySczgBHRz+vCjXGg1XXp699jsi/w
gRZ5gl97ySjmRqpWs64iijQoJaQjNsx3kYe44OWwGx+i229AEuvGiMEbpL4DDNtf
jaVDP/BMLZDap4clHW/UZm11eY5UlT+AcZE2ezLb1E0C9KdvrDnZejesHRNrQzMd
JXIr1DQaZj9+H8KYyiNHDEn/zlqbY6NQAfV+VNcqnSDM/1N3wP8yzgLkrBn2TBRl
BByMREElSSj3jfFEOQs0RfIJa7De3WlvkUOkEqk1dy/xwHZrK3DkKlg3anKiLSQo
dZoKpu8NjvA4CPn4hPiG7AZwKYs4DN786iiZue+IHo+/8iVXg7Oeb4LpXWVhWwqf
vrDAuqPmSnEV3MC2EdVHEtFak039GWChGWlLzcl5+YwEhM+rNM0sO+WFclCHdA/q
ODzE5C5v8BeWmhvr/TSBf0pWJxMyPgMHtJ70UWTVqZYE7Jg1kuNndJFpUjPmRaL6
Y5KYQXa+afQhSeWiyexg8Li3VYW8PVZaedqvtypAsSEJXKCzYt6WgXiXfs+2xWwg
F8YgTlNrzHsDwo6TyRA7CLFVR3fg5EjGXqLBwK6yEcHsD+qp32Psa0TR5i69jWVp
i+KvFmy103FvpjdIPrfsGEha2zMIvdDHMlm9NmYX4wF4VFP/9fmbgi0CNwAUX4MX
FRJSPg++kScPDZMbIuGEXggpugZjehxKQVb7CNzRcjzDKNrYQQIAxAR7iiiAR0Wk
tN2KcKdbSvPyBH4MBzfEYO4UgSapM/764hKppx30nZcBvwp2BOz6AJyJUohez/hV
QGVqGhUPnPk/Y0QRyKFUSTaW41WNXqPgpDBOKi4RehyHWbCc+GICgsDHsxukvXMb
bka+iN7asSmuVv7b1tz+CM81ceiwqGXN5vyDwFeFJ9jDqfVWLCXCiOpLhXTEt2g7
fRQ0M7y2pV5iAbhRRlwjZ4OJX6tRFWvuzAl5R2xpcuzsjmOkC1R06aF0ao+mJvPu
SviN1fwn7WzqDy0htzOUur2k9Rn/JPiL4mXtUGC1GGY0txGPoutm93qanJSDZt/M
LpODcVXmJjJunsF/DDaa2vfn4aaaBDW1KafMeSDieuDQfnR/hv5lwj+O6EWsDhMm
DagZ7krVkxWiN2Dfoea4jbSRNJU/JcTp3UzILs68eV6ZQ2oTzGU7RD//WjnRqDnG
t1MJOF0N1WY+D/LC/czaFYOwNKBKMRIfv6FZHrCCEe3YuKRs1BFW6JzfF6q13g+l
WyKCaSwNuBfDhVggOerVuTHiF4yFiJBKS8Y7loD8fRCFAaqQA7hdWCWE+l/i3azt
KGWFuN01NY4wISgit2gaqM3UShRL0LtnaVQDjhLc3AauqfoKhcMiVVss15M3oSft
jcXSmxl0y2ePhd5OvnqVIHrlz/3/PmU3PLXVbkKMI/V3K8Sw6Qjhu73mWiiL+HwC
F1L10MVR0QgLRe7hj9PNJjritu1NqETNuKSInr3gntn1A8YlA/8nxVapqdf1GtJ1
QUk2tuqafYSRShWwBXCucqOXefh0y+PHofCj6oA8NZ4kvwUAAEWDYAnG6P4v/kYO
YfHIrUnH2rDR8oqgbyD91ecUOUojSkf2eaqyd3h1B5D2Lhbrb3QNZFGLH6M5O61j
hC9tk/Z+aOdu/+Y+ipG/xYpGu4WmoSuxfdS7Ht5TSSXM4gCV/1G4amCjmHfwaN7e
nTdlNlUb+vdeSx3eHiytGZyw7kCXh4UyC+x79wvHr1YzA2YVsqlbNktWKZ/QnAKL
fZ29N/FR3xlxPHkeuVR5+7VepZluNbm+Bn/Do4QUTbPAF7X93hIfTp+T65p1fBXT
Cco9E7g8pC9qMr8j7X57f02g883zB+SfH2Z1PyRAwSbcEYPv/V0FIZWr/78ruHjJ
XhSKjQ2TEfs9Gf+Yb9ufz9iSR58XDFcYsRDgrjGr+fBR9aK73L6p7/AVKos/kLad
etKi4EAGMc9qZaHHt2Si9VtIZ7HeQorqS86VElxzpJyzXMWe0jvvIJF753YoCKSE
n0AsEh70gIQacUOJfDGjmzw2lUj2JmsqS3B1D2/dL5mvvz70vOrlFrSwTNOEi2fL
cJe7azZ84Iyuqx6+tv2qjNgbAwpw+ksfgG6ooXCtzqNkhBOW1qbPrpGOmhmJZBJM
W19vrM2o+KSA3orsE8HrUrWkdQ32Vq3/2eeEyvvjOgDhrATqarcPXTuZpJ5S5dfk
UjkthKjjP/ft8E8NHXIRWWjN9tUM5Leef1ySIg3SSpvCeTrkA1bWSR0ZrJrbqXuz
XR+/P+h4HWM6Q3GB3TjZMWONmDxHxIYoRQ9DC2XreR7cVEGBBKla+QI8u3EIuYHq
uyEBh9O3PmOGEqnv8+HazAxGwyjpMkZkWSP7st3mIwFGBH1LnSuImYroN7oV0+yn
LraD+eVTnVOygYfMPYtFGzA55PWao26kb72tOceLQg4uNoTt3/JnECfWApeD5aQV
vQcrxNGdx1sSpYe99z1XJeyHl+jSOkbpZDgwoGMYeRUUJNn/E08AFACvUa8YOusd
t0Wj5ZSGX5xUHDYHYtg1XRubAYkgHOj9+8Ys8Z0ZpEZpqGtMfD1usD+YwZYcZwBf
Dv5GSM0D2n2zmc0Xctv1DpDVKQVb9E/e9sVU4oFtyZtP+dv2GpAWLZ77hqV3Dq2+
hmXiyENzORM7rRfwZioduTZy1ACAKAkUsow0kMSFBxRjBpBtGj4cmghX4dxDBPlL
WEcs9sVZOF3EOoNJuYECeJHfyXN/IhX1DuNJW5LuonXLyh0hwt85adH8Uq4pcWh3
8nHpKZ3N0mXveT9B6hk77NWB2eogljIt9cGkzcz0LF2csD4GuXX0qRjpNoh10Ttw
pQp6ZmQqXsmS6oq7q2FeZuZK9nuDXsFLVWXeBpCu/+vMq8pl/kGBL/ntrWkJxtic
4NAZa6KyZxgrmJ44GJSJMJsBO86on2BV2DQBxwKMsYsFZZYQ3/gTLAYfEl4/SDN8
sp3g9f7m6CpRLHP5bFEJrfFdx23Rh+VOFnXOEltAijTELDIQT6VjZPqqMm1eh30Z
CX9QSyhTanvltz6aJTEy0ld8DzwBaM2iKTwjS7yvuBJcSVAha9vN/oCZ20hFTf8X
5dN8kTPJpVx1XBeUH4RMEYajfcfv2aWtOX+DlxTIHlRu/OzA32iQzSD2YuuGq+br
2OBS82dPbp9lWT2cwP93aLqaEGw2RdqYNAl+kjNQ+HHmmRSGZlIZy0/vPFeA94Ql
RZTQWisNUjeqmVxx3VNeMiw4dkioXS/hOE0Eq5ZytSYpeTsWIBdi9EOmiBfmVQsU
NJu06t6sR6j8Y3eq5TrHN4hgJuQ+Dya/AKt1hDdci5nwFO//hyy1xv42qfW/M8dc
ykgRsgMpbUR2imoJnWhkvkj9fRG56CXQDH+C8/KKjNB/6/Ui/hK6G/v5tgG85zSG
t/6j9ur4D6nciK68n4JDEsblU00fGE+o78kYmvxBFKDXdw1b5xWWgzz3ZbDklcJE
LamzGVVLqt81uNk93RSF6Mw++oRd7Pc0AKIK/Q0eMFv1agKsxReyo8aLwZB2uvGs
iHvi9JdAozWy07QqhJjB4G9gOwPYYWFMBhP8a3sQsvD9IP3gTSnODCVjSKMejciu
gV2epHMENXGM45tJL3Xxgwf7d4mAGiTt0FepyBkYV1bXblLP3QXUsLNDQSE7L0KP
Xy7ZGKCohfsHnuIzFD6+JeckE6QEWHYWzqp7t9zeUvuklVhpj+r461ix/LcqHbcF
BgqlaabILzJJAFiqyWb94111cu7fotHYTMmaGzqEdG27l/qhPCDG8Qujo7t2GmdM
anE8J/oQpdqEd6oSHmkDhShFczKVacBadnJl17R51f28cEYU/y5RgzrL+jXepdY/
Sxu5HyUOHCd30NUrG/7dV38qq0eIzQPqaEjcPuRsChp7ybRezk6MnK1YWXwO5Zmk
SXnCUExw/eTb43HakvZJYsN1I8M0U8bNL55AsOdCmV3jiddzHiLeGV2YQVTjjZ4S
087CHlXa17e9sa/h77WrLhVmtkZRSvQmJQcOpp24wk2JlcYrC8LD2KuIk3VynPyr
8XH08aDycY+Iw+BUURcINzOUFNB5pIY4X9iukL/olP+Fke7bZPZktVtCaPuGPyW6
Y0pHYcHQ4SZ96V33Sp+35rlmliIQ0n7WGvzX/mQLs6J/x2PvrI9IkmDKk7TBHuvX
ldCRhQiQDcTVV+clHRAjT1h5FgjrN/w8j2tZNeWSolaScBMPwRv3kokt0lJ+ST7I
hWZD40SFCyThngTx9pwaW3VMR1oq453bQR6H2hzls4/r4pApTLIFs90QpavdolJo
oeaCgi5ifYF/ELBc+XTnbLrYDaBV4L4442vrswk0yPdASwhBeok2KIb56FHAHp7/
kz9o4w+OwySlcAx7Xm+wKIySftiKsWUf7zdg108AXIr9QW8FdtmK+TiNMkPHOK6h
mmT/0u4dOL97XBCTIMkvbp69Jly6Fx3VHrUeUffn2k6cH4qYH62yHHmyWJTdIsw3
Yo0EyfuC8XmLmScHLynuNLHohpN4NgGIB6p4aqZKleIX4eOTo/m1hfUFBF7Fpbzo
lTO1olt/Bvo/vItIpdsW3KmiLnPE0yA9aPs7eRbCGy+mvCMAbsH30ZE0Yp8zba0S
sqIhclE/abfg8Z3hNZEeQVrG0P/lxP5caMDWiSZ4lvKQsPCKNFg4hyvZJdWiXNq9
/6Q1+JWfXp5Swtyr6PMgIDou4DyZmWXj/UvOQpn4wyarZr5NEdoq9JeDlVv5Oys2
kGOQ9ZdcdUcVtCL75bsaWySifjEIaX2rptYm0WlpqALRKyBiIVTHK4DN3uOISOCj
xuREqlIwMPx3+32Dbu1pYJLIlZmyqvYxD3VzOIhvJhYA1FIHJrkBPTPLu3RKZZax
26vWK/GUz38CzqfifqvTsTxVdVVuWJlnpShxZHsypZPAKH5I6pQ76HCibdIkxul7
Pt0ZCSSZX0pfas8Emjs44Wn5//8KZJdcdqxqFQFtZpbunqNEAY1PE+Zq+2Fi8FEC
TIFDF6iPSKjnUeuNB3ZWYJhBRoN0zEF/bBsFDNYdmarSa8/5JNENxKyKdR/6KZbz
s7xC61H/8Mi1eYN23nsycAvhKD6YF1TMmskTaX1DTdsh9wzOT64wlViLvEhaeFtd
oKWUWNETi/xuNWo1O7XEbgN4kB5vttKdcsPZZ236w/xxDFkq1TeYRDX1cMDXLlFE
+l6UjvsSGvmhG+qH7VcdrOcywDbwVhCdLGeWnMPm0MCKP6hm3km4NHecUDc4m5VN
MY3LaVMOgKzp4T85fcmDzRGbtH+nW72rM5n/pVhduteC0x4xfQGY6zwjF1m60GBU
qLBCkMwiZqV8g0zFGXTiKq0owB9ZM9UY/VpE+Ltpz4XcLk6pcB2WS2FPRRpnkkgA
+F6uVAd9lcSGGXWteAfA2DBjJKeLLwMmaV287WgXpBtGMDMX03cPRdHdlmI9iR5j
L5/XucnO0RczFC7r+N1WrADfbZDswe1fpK0hrBZv+7KfqQmjSG1GwX+M0cb8wbZg
oOUDyNWefW3ZoZrCe+vsip/BsSKdAbv4ZDbQLOiEt9TNkb+1YV2W+9NCRbAFCaZQ
d2gMlKoDbF2oeJv6Z+qx0PmFYdnOLqxzk/trbXaXbkZcZ10LX9wh87r0AtWsIk1L
5d6rALo8fkJZP9ahgM/OTCfokP7RQ5plYYpU1W9AD02Bi7ELowox7F0ihj7yDaE+
NC8XZYWFnc4kK2Xz6RCG4bf2jiTlEUkL/O136cNhvRiUn7ANJBpIdCQKeFPXzSGJ
sNfm1Chf5T8woVRAzZGUK9sm7d4KxS/uDCGEqmf1wWR6WpbZiyFZJ65N/bNbfRLh
o2SgSaGEUr1/uUzJ7ov1f+E3K+FrPluYQdGEYFcQHE6/fZ9hbg7dE7awJlqhEg/E
fDtYXJjaATstGhewR65jyMAxe05KVhMVRTucxGrzojhvMBeKD9GWLght7MbJUz60
cUXCfXu604TLUKJqIYdU62izTsWFRBmtFh8U3g+QtXESMoMCMp++g8KFBjGz3o42
hIq4HlmL4fvQ1o3fYjsu5Qy6BEDFql/qVzLNK/3rZswTpeNqFG0TFKs9jGzUgoXY
b+H6eMLe8H+HJ1vGOUQzi+gtVJ6W3ickD7H7dZvZsPTxSMZ0j1YI1dbvg1FVVqZj
T0DoIClPOgUKVQHGe0jXgO7jVKAMrHQH7FetzMJ9/vnkVmqUJaz5hPSwU6DZ8X7Q
bfhetfuvv5U1cRz4HW8rynHf5WRB6GjT21QMm8eLN3HbPw9zD3LXTdjFXaFxAwBo
0X3Pm2zxZn2o3pK15bMfgMADEaGzSxY/PSzEeqoOr3xxTSyXSZQlavi9MQ4v2mjw
k/3c6KcqQTAjoD5CYznp1lGFLPRNCpR4UouJUy9IRXRsO/4A3E8i5Of1XaJTzvWC
Adb8ndZ7GxO2/+DvurL8kvpSo3znNrzOoBlPsfMpG60JXvLNQ6uccaO77FszF7r9
CAFam1k+wMZZQHxB7dlM9QuUVxJ8CcVQC9koKsiQpAliqZ/fYZwztQKEYLZgtjxo
BF/U1jhy2OSqHqOVpA92niaT5BxKvHtUOYLSmuQopuU9NlpNZzaTZVCxeFKQxFdU
CY2d3DkA4F1As1y8vDLaGXomH/jDy3FH6z/df6dTufZtD4a9vxzRSLYwc9Z33qsL
JkZN4mnIst47YG83Lsa+QLCnxvjAE/3dDOBWjmX596jQAWLKA6/fJHdhBIe/X43w
Uz1ASgnSA4ZMG3ylVxUT9vdTr3QkoPqGeVxEKpqx9ZOSxOKS+SkoBm200nfzPEQR
TCapWWiJk5gWCR4vr+TTH0MsfLy9sqUDKg/Gnsh0C0RjZ3nSo4v1ASK3bRimwoWq
65moNySryPJz/g+qRkkqUpjcaP9S5IOUtHwDMbcHRtFe0VG+oAdSWCmUzLfdBKkG
CQvLn6QhBG9NDyqV/S4ZkG081koi3y2Ze1tK4Zcw0lglU5K6ovrvMKdDcOtd7HG0
r1PEq9ZeVKcAbKxdsoKlbQnRsNY85XzlwqgmiHZcDfdm0ZdEs8PVRBeZPHSI09mZ
9J4felyJEdW0a9vJBzQD3sfHG6J/MmlvDCLrxuP5IkpZ8Tt9Ms/zyfk8PcnxMNaK
QkgKLXV3Zu0iDfi5AX9JxWtqb9f6Htm5xiSBwwaA8Zs6bTRttmG2OuYPSpvdq2FY
8adiNQg3b772cq6ZCLwiTa7x2D8olg6688eGJnoNY3UcgRG6zg9UL/dP8eItMQnl
mdiydOQmQkKXEeY73omBFH9bGFEg8pCf5c6vF5Nl6zEmgfKa5VNcTpavoHuUaRTg
MQGL4Eayh0bgBInSgIK3a4uYB1JMbFDTqtBBUbVKVUTn2t9vbe3bt5zDb7o2xhgT
wDcw2Vu2VCE9d/80IrHEeSFf5WFDvpdFnY8t0x2C15RbDI0EcxM9iueQNhyyp6/N
1ug2HL7QlI9JHu6OkRyje2CqeS6t4L1U1okZ5gYcJh+jvG3n7JazyLXLtH52WkbS
hk1Nw7nwavEmqKfWvRmDi1IvA13uBfdMFUJ3odJUQj4SxBE3tH0d62mNrH4nEpHI
ILjBzmBaAdB0LMsHMA+focG+XOqi+7Ql3z+H/DbtR57e9ErrShVTgvLtKvdmOrC/
1Ux8B/malFKAiLMyhuqQWmMOqsW4dEhYM51sGE22q8WtS4GtBXbwNUqxo62dcZ3n
tsDJGAWIYRarepHj387rD/QGUx3VsGlQwfU9SlO/r9EnErrJvFfJs3G8wqip5wjY
mRLLqOqTDagXWMNL3GRYC+jxZBazj3tPyYiM8SMC0vy8mAAjJBjZ6u/TiXWWjZJJ
Mvk9mw6Is/Ek6hRjKwbRkPG2jMsdCLQSEuw9G0XDNmwpiFESRybzdXycB9VmRQPt
xfimSDTo/8xtwAAZhyzngj+dsWntZ4fb33aMCCuUn0Y3L1kSpgAhLZWyx/PbZrUp
ApR5wDhEHKA6EZcwEayxvK7HmHwUNBHNcEFuFHwk+Zn0bs4mxY7igF+eR8WXiYS/
qxw8zusI5HG020zkbtWdwAO3M33ema6/jxYFXzqWasfIZh7/ckrXKqIqIXSEoOy7
J3he3dooCauVpJ3LBwLd0bjRa9rYRybjOYw+ms94fpqzBsr/5Mf3xquvzPH33IVw
sRJQJqd6emWs4lcHGx3yUGbK2Z8QgNndkrUNPf4fRHYVXkk3PHFHV61WByYNLu2+
E1AKdjFvfFCnziySbAUbGVcIWuH/k6y4wHY0+3VV2VvPBAgB/DrfDWi6VtBDb+0P
HwzurtrZ4zZCAIDlgDHo/gzph7rYb9LMD/ZtgekZ48xh3gugsSsOd8mmdOr/sY0w
5FhE4OCDcUBkpsFmCrEVIaOw91O2h/bOYipDYmSmGlMjNAEcMSJy9Y4pjsfFBJ0s
9ookmFgD/oRGHSaMVAh+uR6lqIYClc2InZ1v/e2+71+W4ADaS/v4C9rX7AqYmQCS
fHKtbnwp9O63iRSkq2z0njQqaO1RGB/Wi0HLJspTv8s9ppOO7CPeidpNnwCaFLNF
HnXDNtYa+WizzyAzqsqKZ+Bx8HA1cZDUxl6dohPAfA1tnECdJwIrtT3Ph5YgRBgW
TpAmtUQm4IcDrg6fBz1il6oyqa7RszBf9NfThBD19X/wJy3EUv2DA0mSpEAveT5Y
KbGOXzabd952SCwgYrZsg7Azc1FzmRRg1NAu5QXJhrsmFeZ8IEdvuHi2nCUAKCYL
2EVf9Nf+i8CAluShrV+08SS8a8e/HG9RIYw+9UmPmTnPyDvr4Gw1HGN3ngZuYSF4
LiveT8U83cMfjoXgurW2+2flX//a8IlyipEsm6tvtbd37K0Bum9JjQFmdheX6FoW
uk3D1CvDHFGK41lmw34EK6e2yHHtjOnnFizjkOST9xc9ujVHrJ51kpgATyQXXyrU
gOLOXbBYP9tBAJCzSDQMaQCZpJBrtyWd7zhv+xUfkC+W6MBKF3NPOK2T8RepZ0tt
NMf5iHGolD0CR35GwaJYfFARf6uv9OinX6Lv0GWFji21XTOhzS0HDbpp1hhqCc/4
zBxEaLI4yhnVb0L797dyKM3R4UOFllmyJhd3AtjMzLwSJVoYLN13WV+vGnaj/JFE
+GGmp5XdJITGsV7hD+Qie1A2HLSxpQ5eng8H9zmBd/J9MmKLoWNy1BYOn/hXWNwr
KT/QEgdlZOT+xS8y4W9FQjLTZZ/zx1TwECuvx/y/VeA2DBemKyPC+dUVq348/fkf
jZvBFr4/H88R5HdIxzRGhrpZ/ZpcTaSf+vofIGK1/lTgcHZRaqfkd6VouyeQYvJU
8V0Kb07M73xEHOAYj3RQeWM7XxkuJTYwkknWjUo3fn3CvS7Srf2wlhfC3Em1ORSu
Yz5UK3HTkctyS0BAbDX4PcCm/No2uGb+P6Ji4s3Hpf4BBBGvxV8lAbaGuQd7wGPW
Ww6+wdAthRkcfg65XU9pxmya6zP9MKNdrEhRiV1A3lE000721cwfEH1qecv+KtqJ
12onHslhsIhZPBE+9fZeBdTF9+JDZVtwAZwExP29DHN7k3GM30m3nwUqY2Azdl9Z
hEkKe+x5p5SD802IRg8vCIZSmdNL9J5y+rFdgpYAG4iQXe6eLRCaTMXaItqgmqOO
CqyFhCgLvALkAhJrUOpm2XoblgpPOJjQRktnh396yn/d1ko26jKQj3hQCHC/3bgi
pWsfEUrCuRQYDIAv7SJaEkZn8nYmV/K+XEbu6QMADB9uj+7/jYcsSx1vwOhXTH62
acSVEKHpVNYT8/sPLZNhr84Czfmn/FJD9GthQr57T/+KTKM/9oSUi+8TougYgKsb
h7Za4eV+3xAGn2vWOFsCiZxs8WiGVg2P63JwZNtlmGAd2AI5Gw2TqkGSa3zbbx4F
Qx7HpRt/YD2pngz22o19pQDoLeEWFz4KlbPnZi8mRCA1nAqM0LRY6uXDktp3KrvH
psB8Uz0YOpJiNUnTUsJd4bg6xdDVmTgA3dZjwj1ddyxyX0Vp4SZB9/WGnnbVAvHn
drN5fAYL5M87JbUPrV3ZjCMUx/R8nCPQC0ltqIwp/lhdvFth5Bchs+iVtmU/Sl3S
7UHgUJShKe3jSHBRJPDW1qs2gJfoEJIfbuhYmgp8ko1ArhWOry7LazSdaQ2qdU4M
WtzcfKC4Nmsydn1m87KWqcfS9rJF6MjoAvMTz88BY6HTuQFpRSYCZXf4k4O9vEB1
tkQKarlj5Ck/pENjtldtIUgP6Ollet1uH4ul3kRAsGE+QQN0TsTljKZvLGRr+SGd
3VHQXCTav81ummLzgwFmN6ke+37z5zpHcpe/LEEMXLO0Nd8RjCNOSFZbr30pc6AJ
xbsAYtNDqwwBtnXCYTvj27QwAGIybC1nGwxZqfKdn3SoGa/KBoWiNs0aD83LbTxv
/8MJHz4xbpuO2aiMBuGVp76oGpWuR/w5KvRf0VrVp+Lc/YH/vKDGY9wYrSp6MkCB
Tns905B/X7TnnybDSI5PGexvL5N11DnxLJzFk7m5t6TUbA1eCXdftIoFYBgrL1cE
tAERPIqj0Nu7SVTbLVjphq9O5+/nKH62Qm2nZ00f6BpkjXZOWr8UlSkgbA4oeZyb
vxqIxcYCMmB+cQ3YKqoUG8WC6WGw6gnnwMwfIsXjWu1Q81Q8CjoHNQzKoDU46DpI
5DykQAiiekqRMxuVmKURe341cRzPUPqPGdpzpLoLOu5ADp90Uo7Odst+taUghlvb
Hp2tenw4gFBBhxqZn6il4ocYTrfAX7qElIIv6mkJ2CrBRXJS28v7uEUa1mjS0clD
ZgsjdBiMYoWwalX+zS9xhOnpD+vcR2+RP4FBl7uS+dUI5rxjotbGnfjdYPzvcEcX
y5k2TPZKzu1p6Y5coh0m2jgpY0isnraRnu3jNjhDaGYCyETfu4/EqC9jJO8Ngjmv
58sKzf+UUOKMODs3ENlhzUQO5LlLeQ7s+X1Syjb0BUfYEWGINVHsdnI6XSGj0WTc
jyS28bkAWCWJshYFZqKhWGLgUVgFko+9AKFZzdUwgtlxK6X055M+Kw98BikxibeH
MXEnp0/x1RCqhOxsuGstB/DwTF3/Uww+PHPGcgyFJ6qkHd8g741MqXNOKNXwQhWb
y/OpODfOCpti08H1zR0QIU0tAttYYTo9HgVwgmvSsZLJ505cacHPwOYh+Y7KrK2V
ac7xMCVAgXWioMJpVX1fihZrlOWYAooQdjMEG7P/34LBfDx1lGFVzv49DJWsX8+o
4+08yQ0bEyqhg/L3oNC729EHo+3XZQdg1jFl+hghjQEKAU9/HyO9Z/Bby5IdI/tu
XfmsJEPbqVyoBHoOseNPLRmRzTvAe2psLwpSfQXqOky5s4FdSy7UzpoQSuTG0mp4
38MS2aK6RzIYAAUgymtQUT6AwwzE8v5WoAhbcVuhcDYs36R94ghRA2YoGisXSCmk
8M1T4TBTkN/Um0bW5dyqNL9va7OGVainpcIrhllASAUIAc92YgFobba5v6Nu0jN6
EcH8hvqCqja9TPEbmM7wCwAw0GAf5azERJb0UDGTA1k/Fa8OZrOxqvz/6ouPLs69
uoFUgLrTx9hgA+LQXHBTzBxqRCYB/8lZuizn4vvvNHvEYnXuyQAaRAMIjhYjfw8A
OIx4C8bGwUt8GVpMMJMdaa04WiQ6dNWa6wEvZva7OP0c1eHYl0rvT+9PEL+AOGBu
Ezk7zmGO9H+Em+ZuQyBxsK08NeKk/EELtLWckh6HGeC1CU7wu9Dy5y+Gf1Wey82L
iWYBJk+BY6JLqxA+iUz9oLqrsbQdBurzMnSobpPiJk5wAb0Hna/vzr9kWxZzJmTi
prilg2cjWaj0D5oR3VXzw0vZwUgVHda6nF7OYiO3pgOHh4KfQg3EquAUNYoTa+mX
o48rMfwyMbC5PXlCme1t/mbXbz/PX0ygCY+3sFgWM5x9nS+pLa/d1VgxeX1DzNSj
iNa42TxWpeX0jvQw3KTr+r0Foj5D3OE4Tr6asU77JnkaDKzKXmgOkU5P6G2jlSkZ
BV0DDK0Cp+Sp8WG/qaHh8sCJDi9AvmCrpdJEdgARYIiqKq9IYLGC6Zq/mQsz+x7c
IBOmkhvLOsYvxQVOiMtjPEmT3huDEvB+NJctigl1lOnA+Db6rMivObkGP5tM9On8
EdKhHxH5IWTn1RsQNqJLSA4hCbVIQ9SyrcoPWp3cX39sfsmREWvNcJJ9ZhJ6DsTZ
jIAYys42kKzUxBDQhsKXg4MqYC5/CyqFOYGTb+DTnbkrV/bJKizKPQK3czRCSFca
kkRa9tMcryZY26OLhTjfSE7LWpRHAA/ZsV+0zKw1qhZiX4qKEbO0rQv5OwLcrY1V
6+kpTHwpthGXWEzDKIgHwarqpT9QalKcCKvK0194UputYS3i7Z7VTvU41HBOXzUl
wLIx/261B+IAX3MQJcKlsa9ex2T/SVNCfJ6iZX+87i07vyU72bHLwe6Qzw70Xz5v
CiFrCMDmp7wrU+bJiCpPIkoGkbwfiKVo1KYZxrhJSulGb4XxpgrDFrFmdT1paYNH
pic1Q+JBMkgbgXl1qYuMENWpkR01jtGA3a8Q0PY8IdZetlGN/NLoMqOvcUWb+RVq
9WYgER4pcSuycXmrQ0bvCCJC9Z1zAlLmsLVWuWcUZsUEUO2wRt/GD0G7zVLq8Jrb
lDfmnHF8eppVKFQLhrj70hzsuDVc12q+gsHj8Qsmdd6bGCHFq/eg+AiR4LlCLaqC
ZCH+fj4hW0ix2YMmE+wWdUPz3eWl3f5OY0cmTGNL7g6snX518brJQMpHBg0MGcV/
kuEqyerU2eGUMjQB6mLpsy2jbO/0IZab9MSefmfrKMNydDI6sMXlojbAYh1HZO/c
xbPDuc8xQRCuQH6PxiyH7ZhDGYODERynmjcUUGNNgLgqlMcAI/CQz80xG+vxpVhQ
l3Q8sdZUE6/u5qXZ7k6D16VqKxi/c4A/z3IWwKTylbPMXb0erhrzurnNxBkTxoI0
Dmu7IuFqNVnSrYHr1ssbZYk2Eg4lKzznUQTerC0SQ0WZ3tcJtmWPbgOShzI43aL4
k0BBzFiFIjkTyBuD+0F1KpOZT8M22876WHPmFgCq+gMyblL/L9zCo+sGcMHquPfB
JahXEcBSdjFY1OkDjVhaOBeEllZq2SDfOU2dsnzplsYIbiF8AqTc+bGVgITcV9z5
mvTrOnZEFoZUtBA5SmmUS4M6T+Vj6db2I5A9RGSV8oWqxXe+QQ0ql0XtQ5MFoIZz
Y/2gsQ+FXN/GYeeGoQ+oxugRfuyZ6nlB0pfOeORsZkrRw9pxzqnNDePK7+HVjGQ1
XvvmfzvOJXQLMxMiOgIzfO4Ngle4CtBDkUrKHPoleT2kUty8x+95ucM2IvOyf94q
KjeE+noxjP0p5iyNVRJCc+rgwVSe2/QpmpAxgvewqe4qREl+u0c1nN4YADqCoUIS
M5iljmYpCpapRS2494lwhv50VQaKolBUiEXWpowfRLRztUbep1F7SGlFiJX67vha
IHkL96KMR55/EZkyskXv3WOVgSH0TEFlAAZA7LKw67ImwPzigBQ8N3J65ej/j6EN
bC0nyC3Dv/JSDVl3AE+2YNPyCXJaBJNHMW1PTp6wMOVGxsesoPm5DMYFA2qC0L4G
QU6gZ7CfGajsnsdjBNsjT4FvJlXuSILbMbWL/vBfpcTbbWfDUFye0RHp36H/9Yq7
13ZCWvzYGY+8VOIF8tWECZ9PAvvnjkFC3n1gRISMl7Zo4b1cAJqgZUpQhmTwKGs6
l/ZDS0BOt9wwsZWJU0m3hQlRVB1nC12C6C5OEV7hpy9n2aNgTkmTFRqaLaaeEcvw
CJTeOePv8ZlxyxQmnRQBI8kukBtNVtivkFQPslQkfn0rVWyLctYWrNJfFFPFcn5g
FSBST93MTHNC2gd8UH4Wdokl6Cr8gvu0Qc3i0jsg36e5CGGbdwzqxeIuajln3ZNC
OWJtXsvSHw9CTnchHTLv5cXKpAZIOLpXyqp5oiywlabrZd69U6yiGDFZEkjNElGT
BekpAdQdL+VXLSS80yh6d31LYG9LN8CimhLQFb4Fg1AkL1UmVV1FvvNI8VNK6l2X
J+0OrUePIqTOvQPaQFa/G/K68ozidgmxZH/Md388PO5L5MknRW0VON64thYn24b4
IEOFS5v02Soz496LyBaxd/HMGFavq1YEYjmqAcCbqkjLlYZiO9IWBxJgnUJ5iBQX
M6U2Y2m1lbXF56MTd8VNiaekK+Or5PpCSjmFSym/Dpf+YLhyQCKPaphGj+YBKjSp
i5F4XtYsFTYRNBi8Yx4KDxr/G2wn4uN7Gm/bwezi92X5Kj3c6sB4ekbHHIq8Z/xC
81ZeE7m7cHR3U61jpfw3CGlUcVtMWR3C+pMQGt53/KV0waqUh6buRS+E9x7kGMJL
vbGh5e8DRJhVpA1gvcOcHQYjJ/PmVH4MYwSbO1dmCNPtUU8K93cHQv3T0aP7TFXh
T9Fa2miVtwVCE9dkVZu9KNENDhYDrMUEB3xnPHs8tY3387qPF9GRxy6iiE+6oP2o
MBL0bCQG3wC0b4ZQPjYjOQtxiWa3hwIQdPYhZx30cjJzTiEXquzKBCT4S43cgqZn
/uNWmmL6leS0xstT/fuIwJyk77kcrbzFeh8gQuN1Ef6GRq89RqCPZZDTaaTAX3kB
EMDmnMZkM1acvm6/EEJn7fSH5gCLgRLyROfU4mKN/+zAbUZbr+iALK8V+S7THysA
lCuAOQGOCECQ2jx++xYFMIc94yWaWZm7E/qzzUKowDunjq0hhwQ1EX6ssZ2hgOAf
5pQHuS43dIAUO4K+7JVEq8gQgXYOC2F9ls28oyu6KvkW3uXVurMIPsgXaIXcZ7d+
YKPXt8pQ1emV7EyfxFiy/bYpUd+sXXey6F5E8AhpAUHLCRLJL/zpRk7bGd+r0BYC
MIF23xTjqJfGplpexV2OxCp9F6xtIcv8QWuqEzbZdB696McyyhNxg1dDVVVUJeTP
niig1VyRVhKrvZnFmMlTr1CJjwfTKSTxyMX+9c4/9SlQ+l48IL8c4gC3TmDGH5uW
rxfI/v6QHC0tMscmsn60GvJeQeevbWBd/SPIKIkusio6tlwl47Li9geKBYg+Riem
thOIdDaOdCcx2FJ9b9P3uIfnYzQzRenrSf6hJrQJ5d3aUufA80a1rPDTbgv+kMvA
phMl2nufFOmCOq2FgqwXmjhiaewkj7A0AcbE0YualqtVRBu6vlpbYAVw4xz4QP94
NTUkKLB9y1aphJwMhu40D6I2lFc52Y0Sn9U3doQNvk7YE22kpomQkgUbdqjbK6XC
rjwO8t1UtKIdNZMFmkEGD49FGlBep3OzlH76VeQ5Y0d7SJa3eGflmy6AluiUHBLw
yEKJIdDwxDfE56Db+x3vI740i+PI6X+Tq4e+N3jh74EFljR7rVRKUR3KoeMAhvoY
ffC/nkD83bwPBeqO4f+2+Zp2/N54EuzkV4o6J85fS63ywwpIyqmeoiEJarrfLOPM
+XY+d6q14P5BnGDPT+hdUSEi9wSjhppL/hjzPTYI4nPHKovNyUnP43LSJcgdGE/v
zg09oWtQdEFlcx3N+RebqOAYG66hTNsdRqWVGZ1ORhDEd0dnO6WnLsWN9mxK1Ae+
ofRWDFTP3RkQfMzH7y8IOEPgZnfp7A83upxTXzLW1j+rD2TL5D0aiEtERm5SBaFK
4X+SUB46+7RqhJQRdsQ4+wdzIE4aJkKjDP5H5vFMS4apCc4uvXQRPlk1pDGMwP8A
8XNGUaY9zl+D8OH0IuCkD+5Spjan2p84XM1FOqpIyVc38ZLfeCgU2rXHoxDo6b9H
5/TuQuBurZBuHP5rnli0uY+eplsw6UMIgAhtxLkMHocScMcBytG+evLUatDUf5g1
uZkLjk/DgKpqhiRbcYegcKx7tIuK3cR1dYT4INs1vCBqMOFoObjnBQHIeWtuaZZI
HA9AnuRbwiP6P9s/OnBWHWHXHtcFpdfXRxeuPLBW5WiohCjaREUFBqj+msuE1yxF
6zPriag/VL8SFkWNqMiU02z869yUAW3C0OUsXOIXYCGjKwiOknxS885I2GoAZBGi
scD/wqhCA0obMtqYjyvWMIrZtAlfpOB0rEUgBsYwu3jWujPNTaQq9vI3gZjeYEB7
Gwi8hT+RYUgANxbHFmmVykjOxrJFeNuPezU+G4mSvDcXaQ4t6A1eaSY1DZQel2O6
Lb3He1IrEKhrTOyVoQHstRK+YKzlX+dPwQis7E6Pq5z1XM6Ov4G8qQNIlf3sopw8
+72vC1fJokoauZsIQbU+aCk8e5IQuZ++zCQHqpvwh6gUb4t207AxBl6pycnkYAfS
R71PdNG3nYZpDP7v1ymdsvqnZUYVGFu9XlRPW61OEtrKIO8ns3QH67nYHRFmDBsf
Nwu+PzgmBvwcBqCnWjIhRM2OLFs0Jfv5GBVUzBcM86zKIim6Rohm6IuESu8L++om
VwvJM3BAyF1fODDxIo4wLWMknj/56rkZnXWXF8EkaRBCRPKOQqQbCNN1Ux9eWxLM
oxIJ9XzXQBL8aLNoLQOVuEAamNNbE0epWJGVBA4WJ6ysFjBJYowt8lc5Ke2VJrqS
NouGH+62Cdq1UIKqxAJvNPVSfT73aDywuEY4mCAVSSGBiGyW2P/82n25vH6Bayoz
LKLwyyVbNVdQDR3tsGNRCpA+TouRIdHwQpIOHKsSjrA+AzEwGru3Z40VDgO9iTek
fmHPVocxuxFApCaBvH1qOaFmwLNDgwCbrZcf0l7utEOCNxCC/3wUNliyDjGa8x5k
i9xwns6y1mYS3RH2owlvTWfz36twh/muweLTzFWINspQlWvtSEcfu+VRQQxd4Juz
Z9Z1hw7cMi5l8c8vGnlH1x3hESQkcD8WiVPzm6y8fiCfMgbyhHBJMW1/2DQZ5pcZ
Aaf4nBfsbKg53zy9VmJNRUQgwLN/gL2RJkVJQTxD+GFxUSeMIwVtsXGIYA15FIeT
YBKBFi3Fz3tqmIM0QfmVopXKpgssY9/FcFDEGKXnQXs9sCgYBJK+xXfsJSnXxPRk
db8YxW/FNffM6RblZLx87RPPkkdlQR8X54fvJ8z8BhMPo/b8lcism4LfFngnWJq7
eJVHWrnfC1Uulp2JPf0QMcz0Vfc8CtqTkPYU8TiMKpok8FK19n9k/vMtNaw7dk9F
cm6XwCtanu7R6fehY8cPGnIZI94eBGGjJB56V6q3QUhLlh7oiilyQLXr8qx6oI3P
hPLl8x4B/PFi70ltKb+uy5Y1D//cxKo4MVI85uo5z5lBibOKNSDtW20fkap8+lFb
h76zVF6uEPs8RQ+aewA8EAX8WItM6NL5tWSCe4doTt9Ea2OsEFQ5iJ54WRBkyx2r
3tbqXkrv7nxB0yi7L7W2lu0tZnVA6RxMYKAnV6Nu1FeUezxcUKT1RUFfO07kZiTA
TJmapQ+6GvQuQegHWXwoY1UHcdkllplbgfSbn+BQtssXoIEAlIfeaP2MxfWnymAT
dlq+9v2N4lc2+e86d5PhmAu6vnNks/ZLkqR+mUE8KYrWaQXshf6F0z6xPjYrrHYr
DK6bcBboHW0eX/aF+rfIceWWxowGhHH+nhd3juIjAVktOd/VszXMqrLKcMbKDSgw
PT5RS8nmKTrBqQgAiXtJoq3oMYBu/w0FCy8aT+4ooXvLC+W2hwixr4Cm43dM3jWR
huBGACu9om2aaR3k9BLMHGq7RqdVIca/Ul7Nur3msB6ZHiKu3EF4ckak+JPVU3NZ
bnL/N47j9TQwjdAqgW3m9tLzMVEmGCYoBtY+ulNN9Y7EbBfzCpCABFPN9bgqtwda
jYbb4YZ6HE/1V6gTfprw0A4jwHCMGq3ntCnSRnpIMtVL6y2UBhIWjZpl1A7SmIrr
iiFuTuMNXtQ9gWDuvsXHAeW0BNGpdnpsCkECX7O7L/1Lz6PG0cFe1BN3FkmoNOcQ
CZxqztOIhCsnj6dOUcnIrwXzzfOeYCnpO9T6l/6mF8WAoE+YkOnp6a5nuFNOORQY
z72cboQKrTcCvZ/gj08QjT/x0CVbnsUiWgK0UDAqEYPisf2egS8PbpBQoX9IZnvz
vkc6S/xYiKw7rgp1or9ezh0/vxH0qJFOyhhNC0DN+F+KjTxdfZePvSP97/aOJd2V
p9yqsSNX3+pPpcj4U+sBhrrZeunywdyxe1IgAw9avCijdLYxLHlun6H5e8KLqFJP
Vn8WrL/T9VtjiPoPFcZEwU8TzHhb/O52QCDwQgWB+SSZG4J7Q3X84tRHhxgKEDt5
+p8vS6bVP05X3/iymwn9r8lPL3tDN4coIK75FQmNMVsAUznzEhxDxUZD6UnybzCN
Ooa0mtVk7pLTmJ42r+vyknp2rKotRbztdbSAcmw9v2jp7UdW6iLuONN8h3EbqT6E
j1L1dVV0/45cpVAzeah27drBjSVanFgG+Wxr9wN3DLhibDALDE5xlYjIxpYqwYPC
5QCZDJQQy5P/d2jtHR1JuNmGwtt7ffohqdG/Lh+m7s3WjqAWfCF1st8ZrkRSbRp5
rD1JbOZAzxEUX9/3BxOMcDsuCTTPHvlgDlIMRt3D3SMbRduPmhYpGzLP7v4gh/bh
qMDV0STnEEZsSKhMIVYnM2lsAXNrnlTMtLlv1yRE+z+pngMxCkOIShrZEwvdvZ95
IEadWfyK0YevvhXfWktL2cFlo/lCzi/9DGTCy3fco59KUOfCjxCH27ES0ZmS9M1m
HXCP9kgBuxma7wjlv7PGEskyYtP9fBJIHJsCoS9Jgz9a16YGX8CvNE/zFp0PqYzH
fuGQ5p1fnqkZxlPbOibvw7jzxVlXi/5TlwCuC2K9VtyrTvkF/ITNSOfiFxKax9sF
8QOZouqNd5NUMrIqX0h8CGRVn0vQPz8eeTm02KB0M7I/AjurF4ZY/yMV1CnVdpFz
Fgds4qe1+h0u7Y665fN7ImJvG0Vs2YmQTyHPIohUHEkXH3vQmxo4VepltX/lwrrJ
hAfhnzeOKdaN4riNYjW5WDfrDOzGvX7o7WDLAfDPfo698JaZk1P6MIewZB/Cl4aH
xshJ7p8oFkni1SjC4kdoeqto05a7UKlKE6AXYaAKBGMf8oOZ4Oz58raldYqOKgWc
UImG5Wx/cQ5gUXVG6rzcJXNKVle51zoEV8Ki6fJ1IfQs9t9FUaeNYQjgHp4g34YL
gsSsT9xYGXA9JqsI4uODv1naBWUZ4mXStSyPsjIm/ayYnM0G0+deHrTyPE1F9Eet
HOd/6R/ISJknUXypZYNJlM7xHSR5gqyKXQbL92rGw7h274DN408dftkpARgN0eUW
dS4NoWOTBAX9za7jGp/z5JLs4AnyeZwYQgDagHkkYQoRA2+RJnKnBj9i5hNT0RtL
YjbDXWCvjGuHTcBWQfiePWZ+sQFh96f9QpvnxxyHlp4ymVHjFCJnFMO4LlFe4Q2i
vR8bdCCk1q44VdqtkhMHNVJOjz5U++Tb/hgfM3w3Mhob9ZzM4xt7jTHv8qJ8ITOE
Ge30VECsll1MRdjuHojLlhnK7DTRJIgIqWpSFzGHoIF912rrnKcCrLgejI8nzva4
JnbxzNZmJx+YWXMhrCwNLZ7kzrvkBDEHL93zPxkUzsimJ+J8GNwH8AZU1Vx466NY
d7MqczvlZVyPAwUpdmJ9ajzOyAZL9g5TwJHmXVUFkHuNykd56ZXrzhtYb6FsOdji
iYGagGLEZ5laCldD8czMA7zrUX0XfLf0mkyfEVtin/+uH5UMfviH5MQa7bL8/kfm
dxTCezIoHHst/BFG8oQCJ8U6jrFmXpjnPa0hC/r5NfOBMQMo04cpfh7Q8pvs3YEl
LDFXpsu9PZsJQZePTFGp9G3dr1O2bqWqWFQnQG5zHqVmK1fJ/djcm3V5g3tcMjaz
lfGudkMNI5EiBuv+dCKpFdMJh4/h4fSl1sFIUDYbXuqBdAgtfSIkndwd36UBr924
vRf6XXb0Hj/8Z5DNtWa3cpXZJx+E0wk3AUrB+abJbMaZep/g5kVnD0L/Kn4iFEJW
oWHuPAaoDkNwW+ladM+g4t++0Ybv5RPgCjvX3INw7E20R5qjGLctsWRgSyilk6Tb
d9ZBNSxZhEG3aNkzcdRRcMsa5dQTFvJBXwyd6vge0rpe9pdL4Qr89T44UuylaEds
SDGCOBk2QDSYyYvQtYkfRktxsruY64bR0mlbdQ4nzNb+Zw/dKJon3OdglCJbP5uI
Q6Zs+659+Hw0zWnBTGsyUrW2B3Z/bgqGHVKmW5DuBVU5Otyc4lk8JUWDsaGiXvGZ
ggkiMeG1fS+aZ8RpTvvlMcIbwGzcQUG9d9iQpPzcc+U8addxEwBW0zwFbjXwsbuv
Djh1XZwztD3wppdoGBfmXwC7zfMJjxihLbLRJ34PLQvfQ4O5WYIutRveS+nwtcLS
sDaiRFbeO+aY1BuJudRs9+YOaYU7OFlfp4G0hT2qtfCS+eAkaB2jnu6LCTnDdV75
QkwkpumLNnJqI6+HzvID6khFn3RiKZ8Frv/oTLzYyzE3E3dTfRXguIaooT+VVUtC
cWWrxoaeG8hC7mXwNaWL3qZaR7p3EospoQmmDx49vt6FIQWIPpy0Ekl4lYpl/gBo
3gbRr79as7r+Xu6s8mA796ou4J64xWJHxYENuEjZ7E3LuwkKT2SWuNiG4khbiUOJ
JhtTR8HQCBctmbGc8XOVbygsc+fQxlb72FNt6XxLHG3CiqqGKPY/KoQnfEn343LM
ajMIKnHS6/pUr7zxzLvPaH6EL80yUVpuT//h11LFFPS6dssooTfZA71T3SbBEx0s
unidfkQxBY+oMEhcb8fChMM+up6ZHgkkUnUWqcFnmHDpJkjfrGThx8lqzZInPfBY
JS6hfV1vP8CFjnrHhYT7TKnJ/rl1VyBxS6h9pnIeK13nt/L53z7E91OjKq9y8Oom
y6MjaDnCeDYzGGqHFkUOiKTHdEk/72MJmEapYNliR6dnNIBLHLjXdwVLYY9IOLpO
OSKr4MOnl+Ne4XyH/M8qGesER9Xrb1PVlFfdKNd6QUOGUnLEJ/pfED8qswlDq4ff
ovLJ+7TfAJKHICqw2ePZr+g+rJrjb+7JPXqHOtv6sWSTTZlMxpGHxQbZvb8i/jqH
HXWOPMk2ltWLLItd8kGYM2GwSAtfUQDusYHArQ3Pl3tCts3fccwa+6tczQQINUVT
mkaQ7bd01OP0Jub+wvYpKyXPJuvM7frqB545JKAnWzCNJHroTPagTbn3X2kAYoMN
BU6pgbeRjyjzTT5xzhfhoFDeEzZPsZ2DtZULHOfs6/B7w6umiIzGuQWt/sd33PM+
qtXXcymNf4bInojrqBGCfmHlF0qYwwNIEn5Yk/fULZexTR8AJ3fLVnjvhhmNbI11
6a2ZRvzIeH5YT5SkV+auQVpJ1ZWPZU9tIUv8wY9awXC2GoQFcmiGGDp3xZuC0VJx
hbisjEUTf3ttOYCv69u8ikUD2894PF7gAXkj01X/omjniWRHtjNIE8Kx9VkmZdR9
mbctc2e1JpLXvqxhFS907+YqeQZfUXpHRukkJhu5CqkC+CZKg/NATKgbguAzQFIR
j6E60yasKwvQhiSmKJmoTWC8btzWpbKyvegEVgAYwB58H2CC2XwHk4cADWPd6Rfa
/406H+aWcczCGf0tR4s6V/tVPV3kvlgXmRMkb9M6kbLTJbsd8+OAkQKYvoHPsQPD
NRPLAfFQC4quZpBxf5yLExVmazyNl2F5hc3qJm5yDYASvA6d6k8d2WIquqgC3vde
RFoH2Hu8qOqXxXvC+vEHVmtJsilTYRSSYUYBPevLix98WM+YTmTNjKDdoFxPtwZQ
fPFK7XpvBnohkXyJB1nbWPtxF19cKlwl9dPz1GNeuU0hWmMUTFrbq5GtUUcxNOTP
Gmyoj65Xsbrj08UVQRe424tRgM6RnjSZTVJ96DPaswhch+j2mKJ1cPNujC5xg0w5
/Hhoxl8q7M/y6YAqBW8lPrylSRcEoK+DLTjsmNf98nP5RUFtx7JfWjURDGm1Ubwl
Oe0FQBrg11OdrBG8UvzcgkurWrYtLRmex8iADQD79nhYAK29YZAWUYTnQOzQovdj
h1hCnD7o7TfR+7Q4DCEiN5Uk4YPbsfq4q+SH/nHj6hwdE7klTel3DDa5uqUYbkZy
mF72FgCUA1yuK+QQBmZpGLfC7xrIGljOEC28mgX069al2p7Idr3/rwtiZw8PAg3B
q3SRt755RapTRaKu7T5YFlsBG/5cEUSnF1v5LavoawjvaFLBIlDWg9ZoIsJwh0kd
bxT4IBzrbk39S4eCjdAUFErUDcmcHleY1m+lyqZDdIWmf+av6n7r32bw5fnktfOF
1iQi10VFu4v8usQnPnml6oXOLftT4zkBvV75+LCkFsbidZctmWEwh2eWq6RQucxu
fi4PA2uzIvKe2RAohUHGiwN3qhJk65Lpb3GK6Pk7cy+QGDYyn/1217VnwX6g8CSg
hU6fcHgtcy0XVz938ZGmtWr3f/HO8ajAxLPu/fL1lKfB84VgxUvSsNlXW6nnBYDi
TX1Lc6y9FQzXFshEDX+HafnVy6RNGO6i37hUnuY0aPZxrR/a0iZfp06skDEo8tiS
xm7+XQSNySO0JptvkN6LqAWuE1wZqnJx+QNtjwhmzGXL2BbNNuDW4gnVEO8Nyl+N
knBn5JcxAFIoZKcddwsd0KhgTztAhc1TgNFouwY8HnEiV7Nay8X7wTuCB8Rtj8dB
W6fXKn5mfXhBdC6PCb1Knt9HvOY3WhBvJihk5BtSySw7SOS1lFW6pSgf1/9zbHmr
wY6c5e9k18pJdZQcAc3ak4CC64VpC5KemWiGD982w4uX+7yaFRPDUJ/jRsJvl9AO
jX0g9OQbd0hMNp1R858i4CWg586dvxfbdlx/jT2KUqlA16G3/cL3IUIb/Yp/EOCJ
vZHQ/UIx5KH3y/a1d6UAdWEv1iX1Qwhr/5riNlCI//jBIV4OfqNvZHktG5YLjeaa
osYXoDbqZiKBP/vIFDc6PmsAcO6zy1muyxKUwTpEQAcSInaZuMCo7XId9o0bnWV9
KXxMtYH00XngxKuzSPbJb9fiDBUm9Fi0mPi8Xi/cXttlw5/uMsyBnGP4d7epl15z
TkTyMs12TmeYf+sAqSxrNrooWcctNAcYZIkpkWp9k2fhikqtUYp+0XFsWEIigdqj
x+MSlyWv6TSAN0VVoq25CsPev+UliFK/3ckfHXU6PcTICB2CJyhRxHgfpIQoTc56
ueHRU61IPi+fTA/IN/hTG/BiaDdFPAkZc9nSThdW8ViVHPlaYuN/t3CxW7DH4K51
JviZ1co5PuWJLBnbleI7fr1hm8ioLy6t41tATkJ7YGXPPWh2tTDUPVQgC3W3ik0n
mncIPFCT1rrPgGZSvS5SdUhkYCR2KBFZdVQ991NtVuMwA7quxq3zFrtMjmnNQCQi
gxVYxRu0GnokCIPKYCNJPBHlS8ixx/k8rHnhiyd1GefSm/vXJ1BKDFpDvYSECAI0
BvD0MubIST887oISDVZWN8TMQ+w9bSfVaxRCkUaRVI5SciyYCsN2yiIo9YAyltKu
KI+4GXh4HE3Bqit5jvM+Br/bifYcYsMs1CIonq/mEnOkfHhvVOqPpeGQEWqRY4Vy
WAJW5WZzI+p2uB98t7zcyJiN2xcxNMarHC3eyPMs3Yp9jwM33u4WzlGaqZpiautw
ijiX70ys3E0iNs+z7zj2FMM23Rg3/Lau8MyeVDu3W/7TSUIStmysVlOUqkOCTKnD
uq+WFhymEDrE663dZGIOezPhb5FhQy1DdK1xYK+KF5NVPunKo030r69gjvlRaWr9
ItQntuCtZ/0qf+9Gf7L+RMrdcwaGbhCEXMN7Bd66ZwUoFqWsqeGhE+OSbXhJFS7S
i3jJrJc4v2wCTc4QEGEoPzbtgknw3wZ39dh734Kr4eulEGlibsiujb66BYGL1AaC
QrxfPTv2putyhbJd+702aZuduPQPKMbf2PSsRL/dm15Wu/1ChKz1a00iD9xgMtN8
vxXrjEC/fIRn7hz2nIn98GsLNk6lnW0msG6ST3Kwykt3Ue7aOB9x/cyt3y7QvMQC
hrknaOcEcDJPeL9LhMQVC2L9T2/yW2aMOW0CuEl8VzcQca4G08A9euUUtNZKYKmw
0keYWAIejZ63i3EIWodkTTSs98zyUFA+fz3Ee5yw1eXc8v9nAdc7PtkWVixkblVx
nUtdpft1FhKeRmRlvbuY0rq909JWQ/8GE/pkIw/NEeiMyf1DnPi6zl3GNWL5IeDh
+ZfGXwfTGNReEgyPVJP35smuYIljypl/VExo277j8jUecUQkhwLShekKsc4gdLJU
7nACLIA5+s2gX3Y+OoIpJF7Q+g+MNJ3WHd7/mQZa1SepY+sMNYRoT9lBVF/jexqG
ofIJueyuzaGMBDWq51E/+LO4jBUtdbWaHepnCJUEuP1TpehW3PzHtGtPjQIISY7n
dHl4ObWErqxx281fPdopX+aiKSK1v8hMNVqUoyrKTfyP449ZgxozUZ58S9VjQn9d
K/BOnUnI167+87uBNi2BQdC3I4mtQmVnmCY9qlTOXRzcgf6ddVeaApnDpEU4QWEv
xlb6WHFesirrq0etRs/NlzGeeMQIhjKh3BeBLOr8CDXsrVB6DBIHAocSBeXIHUUg
bJ0wl56J/w0E3mxQTl/ggcgIqfuPOwxtzoltxu5SePu7Mz8FFW5oQgBswpQlMzQr
kx+ScLe+X5rjyqgzuKlo8sDpRLFK1/j323rejKbXoAzqvp/eQ3Wt2KEVEi38ZelK
6uRvst1imBtjjbt5KCTpqKOqjrdUwxm9+Uhef9+bNYPjSARtgL/6PwGV2J+EZM16
f2jLwah5gEpdejGe3HiL34ZRKYrU0Ys5OV63VX0mQw4FH6+7stx4llcnEM8mHAmY
VyqjXHRCc9vqcQIcmOmaaRtiJVfE4987aQI5OZxDDOI5w8w6nWjd0dzb/WoZmwDj
kBrYi/M2li7SxtnBPueH148UYom6ndj0v54oRDFhPkyzBvigTeppT2Dg5U8hTDVA
GFFU+Bw6s3WfJKqXxNqG9tTIIRm4/0FkAv8paB5ZpHDzXwLsNDcRGuyXr7V2ijfu
Eu4s6ddlCQ/GcCzHsevFD8yrJua6IVx0yTUB1cNCPWg95B/CB5F+DKDvx51HLmXQ
r+zt4jBJtL8TNgGlALsdLSd7OrIWZ/fuRIjsQWCx003R6w72j4KEu3AILZjmtaR8
vzOsX8XFjh149TUFPryz3cVFBOjvMlupBj71E67qn3TXnGZKd5EKGqyzXn5YkVME
FlRpVlyiRT5VoIBneiCS1psvZL/kQ6Wr9k/iFgydzOgL+U/RQxGC8oXniTLp7dbk
XACISukkwJXJ0LdbFSrl8K+9WSs0pFjlnyhvRUuf5JIZoy6EG8/+mjxMl4dm7cHZ
FQZoieBDW7CEZ6zmYzZkOukrg0WbVFunVbxLzlsFwiOFmKf2yneXqLfeW+iExNcQ
E5lZpmDqLGHnu3FZPSBPms26eYFjzBbyOezQusHtE0fOFiAyttxqv+ehrMUKLSVd
FjNI6rhKN6P2Z+zH4QDuG8RU3FnYi247WIjAOfg6a2Iik9yTeTYEbN1ZvUokIOqY
HlvnlOxkPyXgNX8i0VuEkk7rNJQ+Gij0egqzTv8U4abc4kN30kCb5uQ2iuRDyZRj
+yAqqmNXxLM9UcMDLSukZGHSd4fPM6/yk7Yjh8x2WxyRNzGA1HXxDvMEjweFAxlb
Cpe8lI/h+1Nyi7HPmQpMNMe4+/8lqyxa9Wrxq6zKVkFl/OgoizBElMvblNoV/R1m
6F8NcnqkNzIxxoOPwOanrp4JZS0DXvFu6Loy63QhbsYHvolzZNItXELStGk12OzX
ecPmN6haPPI5d4/RZNmB8sPoCSm8REqa1VBEORWBcqo6IXV3B581rlzcznrUU5+H
Gc/GHJubv/KE5ZpJHzZF9yY2dP8ICU3FApWLY0jD72HkqYM6NlUSP7VXqUlvPqtM
ecl1RnAm/JSOLa7hQHWGmap9KudbHp0oOTWf8oAVYtQ0Hx8zG0zxinS/To7WV6vn
oQZsfN90T62NfsPTzjwIKx1ndu7lYWT8Y+3uu7wYIArS28ZgE427yxMrUgrtOZNM
Q/iaDebunSPai5KlpoU2IZPSOEIeMvHErIGUwam5pkgl6UXASmzcWAFCR1l+sZnx
Bvn7eMgU0nuFbbJMb5KVaDVUQIKLw5ozRrvJfTMCx19gmjKzXyVV7qt45lsl3NXl
szeY+rlUlZfVq0CJqImdC/eAz9M0+yCd3xcuxKSyElp2VA8wWV7GX2mrke4Oi9x6
Kc8zUk6moOXud4fe20cbihouWiCYbuhkEPQE6XdQWav9Leg3RkOcgSSKvGZEgoOv
8xwklItwnaLJam3Ou/mOD7dXCelo2JzulWF4e3533vYssXYgU+gqbS+fJi6aqhB5
1hzm+5c7Tk8cMmotFKFJbu8jBDrr95tIZu3ixs8yoc4DIlE7BbUHQzYXRaWKQz1x
lBz5qIv10PlS8HDY19s2GqZUzqFhUoLItusUTEV5ZZfofcQlwRjoLroLSKUhwUo4
d6RmwseVj6Vu/55vKkPhXBQC+KPqrQGgiL8hPV123aL5AipJvdXpNpy3AfDPZDbI
wwFEfIQBsfJUcsAe08iOnQB5LkNviEfv2JZwIaWW7Pzmx5b00WFMp42AwGvG19ko
YWAWr5TEAfLGS1WjqZ/aWd0TMrZXibkTm2GALipl5/G/DRDg5PzWblzjuHucpSUo
i4TaSyLFYxP5WqjwP4Hu7Kh/tQmMbqbY0Jom7z6Ky3qC1j1oVd2GRdUHnXJLhya7
NDDHDeRNOGtYr/O5bTOHYsFyqmkskYShe8Z4Q9Zy1euLD50Y1QMtfi8Pv+S/1ybI
kNrWmcD1HQ7dkIuz5HV4VmlfsxpYflekum4aeAW69/BCPcfkz2dZTVQkrZ1B3VId
ujNYbep9xGqEMt0x6cG1Cync7DsN6YTx2A3LQloN3qFwUa+92Cpaj/tvMDv6cdq/
Zc+lerKgv6ncHbRvsqFTlPyyNnwqjw9NIGXkSOmH19AajGawPbbgsmzhYKMxa3Uw
lyXJwDj5qvnXmZ0dqp/LlFvXXxcFN8hC+1ryDrd7pEUpWJIH85iIOdWSDEfN68uP
TbJ2Ms5ABk8gyahIF5KGytQXqpu3RlmQK/7VxtXPVhXUqcIg1QMJIlO+Vl5t3ryw
wVoY7/w1tKN/7jUcW7gRKHNPzgqrm/v8j3Ji6TvbNflo+P1qOpywRGEAUrU99E+M
iwhpq2NZ4FVaB7zQuHymOGuhgbbnc0mcAMTpNfnyYIld/3FRrFCmAr4AhyofOPyG
ueV1hR7gtYO5ppCaQPq8jj//dHyDjssJfUBIfPrsDv7fDM6MBQ4xuREeVOwWCTyZ
P3/nqLqrgt7fI+DRYFCUSb/fMgdmFM48O6DKHvy2tZ471OFx6T4zo3Jur1/eaAdw
2gh6r1Q1BHb8VH4WKnU8KQIQNl8H8joHeJMa/E5AqoeDT7/vkELbQdoABsQdkV+1
K/E5xHXmyKCKCGWyn1gj1jHvIqCUN06Q99LIGOyCKUvEVU0/JNU+HDllVFb6NoyB
jGBDnGz/1kB8HkWf3FfBI6Gd5f96aXaQrbnjm7ZX5PnD2f0nu38STGDGgW3ebit0
nE+WQjNYJ0s5oukX9Pt7L95+F3oZo9vPB4i1dB6lOzTxYkhqHlD/v1bN009E7OjE
QgSjlZeQkSe5peecTSFpn1tQ3LPss+4f9ZwJIyNKhZZ0Rv1RjdQk3diJsYJWCg6n
PwheiQEf4dx5InMbwvPpb7UIIWadEtGzoCLB3dMJ/3qxkxcYiIb9n1832f3ZHEaS
4fwRfw5Cu1DccRnm2QrhD53H48lMXl4R05i3BqpGkIsuBbH4xyWWePULNM/Lgxwu
4Q/5UVzXG5lw9gL2B7nu43d7pyp/quBXwbctIGiY5tUFOX14KmpvR+7gaCXvSde5
OyipUZ7bT+Syvst4a2q/SsYCQbAWysJdyYJXeTEkfGUG3ar3C84LSnJIbv2GTGns
mym0oZ1XNoZBCdY8Q6a9n5U9b68B15l2hgGBkF8Rn3q8WH+137wHwHGLT4m3oSrD
08WmYOjN1w/KOsoyxZ/eABnT97+cii1X/QPKZNsiYNxmOnYJJlOL/XPbNdPlMcSh
aQ71OS2O016R8CD4QN6VFpz72ZHf577DyG7TE2etzu+w71r3XqYzFufZxZL0VTyO
FNbBkc2HigulzgdZdDGT6iawqeZUl16AMJhKEUlQwG6U5pN7Pv5a2Tokh15mWtkH
C4nF4iS5VHEZkyX0kIOEWg+l8KEHlXGiW1Sk2GywOnqBaxXHP0pA5nQYfXKibyIR
7hyZyXcB1F6s0OcP0QWusl/uKxnmeMoweRCrqqt22Ir/iogl4dA67/oQcvKWMI12
AqaTaV9jST0PKE26g098gG5ainwO+BY6xMR2gIhbvumcV0ptLkCp9iMfWZvkOCtW
a2W1TqUeBY50xGzi9rKgvaucQ8JQXgRYauEwf1CdaCoqeKeN6gaGRIDxLLT8S6w0
SGcCws9Tp7840pb2oBsuqkZNCpROhClI6IKH/O1PNSMdM5OJnMQTXxbp0FaYYlHE
zcTYJCo2HqwLvts6FA/nxr7t1a+ERuTTpoyN8k+m0GtgUoySf1C0S51a44J5sr2s
u11m+JSeo9WItoGA44DhzG1eyIx419aNLtdDkcV5iZc4VPjUS3zmpemppYn0fx9B
9D/dJl3H8LuIe/MI8VXxfUcuwBKQGop6rIulzl4OXEGpg2BnKO4iF0Oc7npxdFMO
thGZgrvLApzyn46QIFS7UxN7NkM0rGYXmG1z65UvZ5G9XO+Et+G/XN9Hbb8X7qwt
FzAufxyLV6UVaoBZkrRlqIyNoVynhuw52h/MFXbauNHuCRdIeniHTMG3cKCvXC6N
rMXqvPAKJWEgK2v2h8l2OV/w+/NMGGZD5PlYB6nv+BlNVTpqln0DX8qA1ALF4J0+
QO+GXJDFz151Z6u60n0kJ16JnJgvn9LOorcIr+gQjtZ8uOBVYSfACEbCHKj1GG/z
jF6fNQPjRv8dn0bGGeZZ/h+hCskrGaFw3L4WnNWKE+UXRzSWL2e4VeWKzQsrJ8QN
mqZwlZT4DuwdWjhIKWc9cACmGxfRIFxYgCUAZu1JvLaN7RkKNc6Lo5ueGR2Tnk8q
KfOK30i/oots12XlyMLvOdQ6a5FVETJYhiJaMy8N5ocFI3Va2pVXxpEvk5pQI21Z
qPmuE7yFjT6gJaPBWfhj862H8+vHZFlxrq0ms71IX5qWwc1H8D6K/RrjuUUzrquR
irLWN8IhunygsnUlR+h4EQMCxg4f8CLLqHppHTWGrOXzAOKwHXsNqC4f3u5Dneo9
/QSRM+e8UcUJCxoLbdpU7jsqTyjjoaYs5mAXrKX01oC7Q6qXxZb/xHOFEkkglyfp
DhJux2hdGACmaUN3fpLefDFg1pKiSUdoPLKHf4U1ZinM2NCVt/0gbfSCmqOIYFJV
ZeCCK1rqLza/0Tps3O9UCgYe41UXa7W7WzGAhw+0UbryAc87ccPDfLVeALaR6xNA
+88vtm9kzwcrUyeJ6BQODdcEVw8lhzpVr4ftCSG6bzSYqK2YnDI3n9XH0cBqNHhd
WS0nFBBcvjGjQnAEjqzzQthhGkdEW9RZ2D2opY2yOaKxfjO2KjchRd28cjoy/SNB
OiVsgEEdYL/4qWRZthiIWkDtPuPBVCT5fxdDwqIIbaMYYK4Q/gd1EWIA/lOaMtKw
jeZWwXTX+CHrNML0Pcly19FzT9f96D+TO4CWHT1jT2yP4HiP2nVxkqkJe4P2QfIl
JIcF2melc9cZLkpaxOzEc2BFX0X/BqNDOQyyyrpcFuxmCO64dhJbvQ1yjMWByzYF
9dPXJIYQW+uz3yAb8hDFAeZyGLCnuevbPpUMRrYvbKsmkmOH/a9VDrrS7dbSKCwx
lEowntBvdXYr+rz6sdwIBkDzKQTZzXBQZSIdYgkPOdPTidZyVaOJaUeETuzYCEjX
M0iuf1+WzQaGYv24wwKcSzFXRaxRDTVLrI/luvNH31l571bde8HPJdq5F+0+tvYN
hLzfU/AKlH2OI8ahicpQDoGa4Y9Z49ga7G3Lfhs6DpuGZO+G0vOUswdfhg8YEfJo
vOLWezKCG7DS7EWQYx+/hkYEGq+YfKhhBve6nyNLWxHSC3FgK/I9AP0ln4kSljjc
hwG4rbMkx4CIfaGjwl0FmNCb9WD0q4U7sev634G4ON9Qv18xuwrzZjHhihv9xJ5I
lfQUXungtuko/joQUjsy+H5FZ2PGD6neAvLsA1rQ5UeNq9lvWkSgOLt2sUHplmAC
YCydUykAkrxRJG9JKAyaSRJiGMRiPLa0dHAzbbZ+zHc25Q4qky8D2e7oaBk42FyG
xO0cwcu3zhGC3N1nK5OOin9kAjVaWL1zaGQ/zjHJwEKdh23tw1D89taV+ggQwLmQ
pO+r4YaGYXXtT/JSXQWmVMZ8zEKpNBnVWDCkTb373hixMO8KEp7thPm6MYsWCogt
vyT4AmQalo8kPFkTlwsW8mOJxo0XKfVjEPR0tdjmNh0Dc0+afKY/Ldwd0FsNTisv
VPNMiM8fPllkKAavkkK9eIvTy7tuAacOaJ0YKVk6+SXlnhoOPoCwitodGUG/G0XT
uUm6iFVFiq1rnXUR8vbvkyCSZaQrFlIJdrBM4eYQdXaWqmLE0c/deYcZnVWovFCv
fvdTBz8pIqWpKXdDqhqvj/CULAaw0iGiBZVctBFO5rkhV00ksI6xhZ1hItC4WW+3
TrFDjUBP07gI9f4fwoWIheE5P4yVinN96dOqOCmMIFRp2v8jBPpY4Ktk2u5Bft2w
LZEJzY0X2ldLXkxAWjRMpvLxuGSQTrNYxqqNM+LREdJKGcZgOWy4puYkPMjQfMii
fusYO6/JqoFBz21WXx5RBv/UBiwIKQJOp2IswCVRzEaYKDaZCu7vPqc6eKO0Xitc
ZUZpJsRdliH/Oh66V1EvHbHyBvQxRYc62egzs4MT2u6hicEwcv6WFz4NsipaYpHS
8PwK0bHHRrW6aUvkOXrxfD6V4eaerTuxOV0H/2rLUCiMAhraPkRHqrKAES4ZzDYq
RGuoQxiG7oeDR4j15XwzlCJ32GdfHhEdfgI60noCvN/82S3kGvQXa5+2JpfBXTF4
N/KfEu4pqhIb2pBgTOmBo44d9G41va6PPla3qBf5Tly3LYYgGhmhOmucEuMBKMMq
lFzfLHmSnj3q6YMYFoqyu1Dru0KVqaakkmoGwUR89nXVs1s3H3F78Ca6OoZRUKmM
bZtacMpMPKUxHYTASwWO3cYskZkTqmm0bd7N04ad87SOiN/cZDkfkvU0ZGRXTVDb
8ZxTn20SZ8o35VoX+fPdKWjw/lCGygIXYyCoN2LROCdZUfz7zvl+PTSrqLecG7sV
mkraN0KdtMC9pvdlEj6xevg53PV99yMrENcUYp9u7pKxlNyeVEJZ3doBEw/NvjS1
50IgsHEVaN30f0MvZWFw0vQkrTzqP+P0JkcOIbrsKXh9kW1Cn765Cyuf3EWvYQxg
rXZYT5a/GSb0+GkK3Qoj9oCVWTEB5vyiXQkMWw+gIGLxJamfXgx/+powPcV2PV6t
h7NucVEU/9CUTyftiPo7ZfrmWfBdpKWa8alIf9OHqUY1Zp33qY3DMrc3KJXSqSVq
mtH00S4dWmJ5R9mH6Z0rV6rakSf1m5dwz+BOIygVKyjoizhcfVLvU0tHvlL3Eth7
4szWLnvLkQAKRBy21x5Jv8o60gI2iHFvt6UGFB9Fu/gc4qICkFFCJe0gbkRoEbIO
2eacgKV/f8y6dqyZsBKw+nOzuttUos7qgzS3cEzh1ExR1TghjbdsR/yQBqLJf9Nu
DjJbbilANksxKhwuL9DymJt6/m8qTOQKMvF15uV9TuBnuIfLm+sqJX5rRIHtfAGI
8jGYKa+0CY8gHIAwk5CJxbouxkNvO7Xzw+yOQGwDxWYbqlq3LAE+s9VVXCW0+iWJ
YVN45aGWZ9kq7NMN2u/NoDhyXxM1c+/Q0zch+vP5Abp0D43CYGnH4bYWP1bg5QFD
6fFxtSMmE1aoi3QONjuZLRpE5wh+rywmDHGh9/8ol71oSroJjC9hmpeJxzpVaPxe
FbtqkkvYZ+CEP2AooEYGLiCHII4GqGSx0E5CRpCcBoA9JpGitw9S7YuKz9wYlxch
94IH8vX79lS0qVlnMFYl58JMKsFKq0+7u2344CXztRsxSMeWWqorYUxoRxeHnj7u
tCiFMUNc7utDpWoZnVgLhQv5+3HNgnq14IDnZsHo+WmvbYfoTIwhjNvZa/LDAiB/
d/FOkNjyCoRhD8fs5836oV1HFUiSVT7xHqL5PRFKA/N8/glBIbhLkyKZpjHpn9E7
zOzZ2yVr08ZZvF+QE6mnOH7YaVdZs2BCOKHioNSiW9Jto8YY6eYmqXXo5iW6B5Ox
+RXh5o9Y7gFLXpqLDJnm9xghNEFrvGuacbSNxM4ICbhTLqH2de4KTHCksbmSgCcZ
6edZlL0Hd3Cm6HmKdIBJn/JqfriyfPIAoKWv7Di+ozMPKY8d8JYFfGYXU9JPR1R5
cC/XWa+tP7pZ2FR+yG5RF/akzo24YcTv67w3VF1T4bg+jPNaWohrv8t5TfX9o3V+
+FaxR3qLdYz7TsT+sEBuLggoEkWbx5T6snvxnbXLyatArm3DX+OM6IMzmuVcTR8b
tyFXa3ybt7UV9aupQADwo/d5YWOi+pj0/eAJeMvG6rDTxqWX4x1JXsfbyy6gIFxC
S0wh2/T9Q/d5ZuCBlXsHJwMVZaZk8Ybn8MFxYssuRhiqgzJEv33hzzWHTqvRylkP
zFkUomUv/SHAcgbzGrsnD0H6OCNnhpmtYYbRc/sRANubR1BCQYg8yBs0z2tLTKGX
z98qpl+LZuVRKbycuA7kHn0jMY4njY6U8wqTBcvVP4Dfcm9xGNSR/UkZL4q1fYgn
VVApI4rd7JvJw1zrNiz9JjQYTtSium7MkjmNBMsEva9P3gHHelp/5p4mncuna4tW
lJS3mbsp1D39YmjZcC3JhV0tGQxr04adC256bcheZC77RVYSN86QrPpcCWYeR+WK
JgLml/8M47owCGn+8kb4vuO5isl70Rm6JkuyGIliRp9+C10M0iSb1DnBJyQKFTp8
dOkaxPNPNcgVbiG14M8+yMCwX0XuydXgEg12zN5o6hi1pdu3hIkS8JpmqSnavK4K
vep8GmPUsPvr/lPd60mEP/NZIcoDtEQ2CjN6ETL7HkyCnjhQgxSJhOeOJr1bdxo2
TBkFMWy1lHqBcamZCE3YEvUrk0I+BBxnpgx3A6AjQnIksYIbecL0JZv5Z/ck5wRk
UFTZCy9O1xipQNeCMGjTHBLG0RD8qUlfqYhDkTOZ0nkj8LgSrgdjkC9ZLAqDpX4h
ZhvZJQkcsnufwrnL2hE3YffRUwbrH183RaVDSfv/PxKBFHin3gXBcpqTOl+xOFpT
RkIYWHSBrVAPDkeRgcblkwvzoErLIt6d9Hp1jbMVEsMkky2Ui8UdgZfUj78Mz+xF
n8bB4DNZK7KTCvstypNe07Rzu5HzyOasjG0Lk2j8eFOYbicWfuokE15SKMztWryJ
xadDqRjt7NQi9nFwpleTs/nGgcAx9i0kPjVHwkjWxLTx6zZ/92DhgDFuYSg/vOki
qBapsAdQirqOgbrX4Lv2nmQLZJDXElfIinIW2EbLNpdAMqEY1WAHniQT/zUQNyzb
0hKUfOSgp2yqSKkL4kvSkaKjGUM8CzedCvi2spwRoBkYtpYqkdChceWNbVTuzQt/
Gv0jII7plOL4oTxyyPS8sQfIDT02c5qgOI3YLams41kvAGUmypo3SwM8lEaRkvAz
vDR/b/JjqAjhUEiEQt3HpQM2klM0tfZWNvUGmWsEJMEyQWhPbPYieTidvrooV/iv
dikx4Pxfr5CyJ2Qkla6W2t7mEDQgcfmyPBrFboOUYxfeWbOurwGhdtGgoJIEs1n7
pXwZSGaRJlK9aZF+wL/tmAUoVt60XjorfBkllebYBMiH/Oz6hNnOhTt6yPzfp1kk
hZdhIfA5lfiUslNEMNGrFTg2XQG/q7DShbkdl82TxUWmDFFVxrzHoFAOk9rSwyFn
A9GTheAy2LIi83X/JxNkEde1FJXMzJTEgvO3/X3tlbpQKXDSeGzOnV7j1j3MP6Nt
ydxXcch293RYrzl1sRz7ta9rtin/msuOTi6zRlFoT8eMCCP2eVwG7eY+DQYecpOG
LeYxgIVVJx9sZ9BfYzcF/znRaRwfPjwswQ9Rzuct6r9UjwD9M9V1SB+cP906nnLb
FHPNpgrNukqjWX0tF49BWv/rHYvsOS0cQ+r4L++tTW0qIZZvyWkLQS4vZsZolwcv
uFNa3OyVNWFmlc2JBVelY/Q+UGn3YW92B4Guqfv9JnsG9vB3tcWkVLc0gXp34VoW
5S0KvaNUmtYvrcq8uAni8n2Ums2iMe+gyV4lEcOEtDdPsWQfg7L2dQnSIqDpLylO
DCRVb0wUyjMV8V/JE7Zi3HMMU0E8iK+ijSrEN8dX2v71NxU0nEGQNXgyTEq8/R9G
QxtGUq8cw8HDGizxDdr0mDGpmFbmvq2HOfSiQYbbgKxJizfx319Fui5upnbEIILS
j82hxkUkf7lOcdWjNnoayS2BS7HeyDa1Dpt3XnrhXYQj9dQPeJ2ATPPUsRkxSMn7
ASEh2FmHf81qubq27GKBbDfmQWl0CVu2eqmMOlv9Gs7QXLSV9uEKdsUF9achpqFR
kIsE6RO1hoDmG3MlfWgmzDMCDn+BXpviv8cUzOXgC85l744ndO5jnNls2qXp0aJB
oiNfDenSvFuhjAdB7aF9H9pK/2FV5YkY/HXVcxIWZt7eHXDUnBYV5ct4Aptrl41y
bkUd/8xAI5UmmPx0I5jUwtgd/yvaFA/Hqok2ATdhXluQEvzL3N957YuQEeb3SDdu
zR/JxkHg/CZIohJEwgjhMaqFJsNPSZnHSFnw0hbGWKRW38FMdB0lc8qVvrnoQ2mM
SaCcY/z9SxriysgbnNaLbI/RDxs53FY5rG7bruJv+sQd4xhr3zfgVSRtKktes4c9
PLaLbAIQe1VECnKu/44YStHK5A53ykOe8cuE8N55ciePtSvcG6PMGhVP6WuVi0Ib
Kn+R+5jH+ERRyGajZRJ+MveUDBtP6MB1cOIk12ScmdXiGwHQP5HfGdtEBLpNf2uC
IFfWIwVlbdTkHPXdcD0qEFcWdIPXIGccTPNmz1AQrIuai3BbI0qKuoIex0o8B+fZ
S3y5UIS2dwnqSr/buJJrZ7UJeDJ8mYf3SAMBT3An70AGZWAjxNPaVUdpiJKDaJIu
Memw0g2B5sZJ0CSWDbqkqed3JEiEDSGVRXlZdkM9Ns3LcjqPCyjt/lAWM5CsXC6y
0k7WS9aE9TGHeQq2a3+GnoA0mNEvBozbFF1fxbBp9VVqdJA2oK1YaT2xcGsseoaw
i9l2Xyjjy6/ynXooeEpVrbS6pDrw1FdnYG1zu8cgmrMfqP/ngxR4qHkfLgn2gEMO
zaTQ/hfxiq74JsZ9WQ+0Ur84PpHOY+lteDOI+omxKSKcyv7k0pImaQPvmQAVIuZB
6cqoIKvnO53H1nmzh+JXG3VzIQNjwwBK0KQ5dMiVzRjlIXP+52WckoODYrdwnqaA
nG9xpaZ+vgCdWoPcaPHvQU/981scHZu4xDy5cPTU2D8MayGmHYkoOIovQ74B+08B
Z7x2S57SONy/NB6tfhYcA4ycyAHvW8AHElOWUIJ124MHFk5aqpZxtYMYU3ZXPD0S
rND3qFCUoBKW0YyOGJqOyddVnJkws/m0d9vVqc+DLydd6noBc+uOueLjCiDAidm3
95coai7P2yRGxjGYX4d5mTapwYczUIND90DuD7nlhS2YlGQMDz0+WId1gaL34dHO
vEdf/YAv9xp+90gK7tb6vRqY/e8PVLO3otw1dt6B2HXWHr1qBGXRyZnEVHF3JWUE
RiU75JAZC19AS0LjlGf52OrZziAGDRUFRM5RQPRaij76rPyjo3tFIjUO++G7UFJq
ODhZ3I1FKhs38DgROAahuPzcH4RifO6krCEDjHzAbEBBJGV1FPoBSR8vCkDfrrZf
30hiC0y7KmzTR1ahc5sJYY7mJNn8ynoQrB3yL+Swc1Xyfezu2C4TJTUfgqUGiJGZ
PnKKvJXKX4o30fb86ZVmf2GW4yUd/my0DPO5qXpzuwgI35whRS1vJXgZ2N8qZdpj
PBU208OGCDIz53kWtNkx8Vz6m8i+YTivaqk3leJ4a+ojqohwACaDvBY/0VFhBWsQ
aRxXEcadvLaMn1h378+7p5DnU4NSExZmOHJDwTNMhd+8s/ShyQ6/MM7CnbIr4SFz
Y048lNSfsmldom69/w/F++ZBVE8u/IhLMcX/kK1OHbFL2uZu2CVHDaRK++JSvTJv
LcRvpVwVY3WL5HYJ13Vmthde7I48g46R7OgL/K9B54GhnHqN04goOjanK/Bw7NPT
U+r0AAo+gdx2ZvkdiV94l38rhz6qDgVvQ+j4U3m00r5+scF2Eesx2jLodiHanOC5
EoEw2S7BwBflKBeE4JFH1sfj8+a/QD5E2aLzc/7fq5ogDJpG0y1vSevN/vN+JeUH
IGZhTx0enJrfJvWwZHTZVFBv5VWUvUoqBklkW6YXv4kU/CbKHHiugHpGZB8U33Go
8pZAsfbcOf6ggzIeO/W8CU0ZoUF8P05SKUYLCgnmoxyQfvAFeyK84zA+gMk3/2v8
66p/kbz+dQoIYjFFcj5WVlOMkhrOyfWpEJSdZHZUUTF+RayJn7CdIGXPlZHEZKv5
aTQvv1NCOI2mXdC//O7s4aBNNSVn/4DqejbuLtTrbizlaffczE9KS1SSizCcIFSU
9KQR90LiR5xG13YnVCuVYb1gB0TKXqmTHzOEFId+nvZd9o+nujMe2IFxeXwmW4xy
+1wqH9rjaIwOCaC8r9HvbcSPVbqm2Vdrcnz0ACxUHQv81A1Lgyauoi+iHOxUPvXT
dqWIYILaIzMDg4l/Yq8Om8AVWvX4kA5hcywgnuAy1N5lG8zyJhxdimIacGqpRZPN
AB7I8X2DIuU1MLRWFjRVWpiAnvfZ6r+4JlBcqaau2KMx6/MHvH8a4Lp6TAc5sdr/
Rv2IYatMxPJMn/swMr4VG6af7A0YgjEpDOynCFBHI+RMImMj3dBFHww9M9SueCOf
7M1AnKyG5TyWI9/YLALIjBwovl2imNqIsNu7S1T6jGBVUs5Ix2gf8WkEaI57A0P2
qsA21270Vgfaztqb73tGE0J/oRZ8b9qSnCi65RwcO1yy3OaEBfvxmIoJvRSjzFrP
eeXEtOv9uYu3h/XnskBKYgiGfy5n9Mn3JZOuQS4lrV+GNnAY3XkFbQUSyZfdJW7u
NBmqzN55oKtmR8HqAInqfxlfnRCrqxAsLFJU+ANNUwgrXi6ON0BQ1TYlrj9QJg/S
4oI1E6K+p930LhlWoJz4QMNnU2k0MWgEe4h6f0vtKFFxZmv9KDdCgM+k3CYx8mrE
lOGiEOviz+rfxpLJ+fLRIhW+4c1OAMZkFXNq2KKhAdMoyNMASZpHUgdNUaLP4qjB
n8+TLAM0PeRM2YdupQIX4vBgJdWOWmUmtD87PCEaBSZZOCgt8YcWARvv4MunMQcQ
S3X3wHoGwAeeh0bq5uTuD5sudAWoikmRRDXIuPawiGwkcb7hTpWmm/o/aLgOuyAK
AAG3MHp5BSTD54XPwPVIm2pxf0mjBkk2tayJHgc5zaSIj9S5Lipr2rBykIBWT2Ce
tq+bnVNTz3E7lSaWE3BdKwxXlWDz5fsIiRvJZCJ/fE37/gDxiyr9sgsWzsVoERYJ
jmOQ5MrnksYRBWJfrEKDDUfm9fIeWiotxfzDOMtAkWRcGGP5wrRJ6kgWRY5i9rD6
6j84vIgdiA4I6E7CzssYkvE7nntj7m4Fan2bo/gxHyRKYGWG52kLSyNsbLUb8iaD
C4HwHYK4QIsG5GNds2FxJtLSXb7JMBBah922PXihw+Kdhag69kvkIGcXJv+csh8l
2cxkhItbOlwCweIxXgMZmqyrB4N4uFEVEzN7aC+LKjTlEkQE/hqguPPkMppvWh/J
qnBc8HxFOV9ZJMSwjxtO9fdDlIWXT/vCSFn/guUJrT7OtpTKsA48bTjVZt4AM5NZ
bCa9y57jpq/xC/R/aSwH1WmF3mGim0Wfta40mXg8nbxXC0aS7mRJDcSdjPX04UA6
T5ZsDhz9afByKboNsVWBkiYgml/geGwxg5XqKIIuJHexMwOX1m6SzB3dksIakckr
Z7ZJpiUZ4WkeWSr1xVF3dUVCmLc6QnZ7C6rMP90PM+ev2Y6DoeT0wITykv4S/lxq
0yX8QgdFQyqZwsARaZ3yKvfDm5lV6isLBUAGQ6UmMvluCgXm2vW35UL0RBoWjKu4
JTg3SacbQTFZdrH+boDVVLPRoDehXdexrIt0j7n7Jott/975jOViiU7uBG2aW8Ej
gdoh4ppkqPo2bDm/hkhBVdByPKjKd0Db0KHm/iaL6uA5SRVjBiF6vcs3VnywbYIV
S9CgAZVTFkS2rbVIlKL0KmFqyFneFU+jER2Sdh+YzXhHxRlV+kr0VbTnHvm+HZcS
tnI9JkMumjSQF/qUMaSpoDeVgHcY5HUh28+f38fjKvZ0/14tW28mkownIy2ApgdP
Y1NEJ7UsS6N+deUibeo+mBZEVAvxhymIGv50+GGeuDKUVUVZEeqtJVZl37aMIVRb
NLNV11cXsufbKWWH3mkdvvQU4l2IpHWrpMVsFOLAD+ur5APRHH2U9Smx9RkkuiLL
yQn9k0y0DT47WGoJWyW1DxL/Pp9f/uat13at39jvwBDOgXCemUD9BrVj1NK/+3ua
8VC5PGHKjZG0PK9nRS8CP3GNw1eshxHDhZqyQWdW3cDSo7zJwML1xABsgkRZOvED
V8/Xe7hQRSZaiPXA0L2WHf5zH/EpkTo8dzvaVcuqUbhJtSX1NY3PLSr2nvxNDBOy
IFvPF1amNt+3mU6L/ypA6u2TuL+7lm4lWxgk0N4LrxCfGiZ9jlRt9jmqoy61YwcU
P4j9k2qnpmVsqyZxC+EXvYLWe0tBM6di8EiOEHL8jv2khzNwdKzZUNn5rsDpXeHS
whBWWtu5hmI/DIZmmEVF6/hZ8Ooj3y8lUByvifzWX2lPcU1JeFPmgRnr2ut1bmDC
bHB3Yt7RfDMku7MJLjOSfEJLmOGIaH5Vysi+IrPQcKC6TM4n24SQstBQGS29To/H
ubuQAcizrVTspQPZLyERLAmwzSme9kd2ddEjpjHNnnclvJ+2SsFmnutG1BrGpIlk
+n/blvryoPesWD107Zn3CSjuvdP7Vetsv+Cu0WbnlxOCPB1/wntorinX5E2orUHI
pvmf8LY7UaSgeQdnaBZDAgRYDFApsykMAApKmLiAba7MH6ejsWHyXEvIUtVYPdaN
TlhAp0IDf+c82gvufbh013dlhcOGXhBBpPQi8fnuYGk4CGPLS12gvoTJB292wIRM
nZhgfMVkHh+Lmr5VKZeW5IjW4O68n6RXu8VdGox4OmdSupPDDS8SHZZNrIbWLcsq
GR1gbRHqGJ2a5GJLFiTfVMzMWBzflX7Vn5st1hzYU8Xnpx9Fkfk187wfuHgPl+oW
FGTzWOaF0lZWbsHa8Eo1g/Ee6Xd60HEPFoQQ9BuqIiL0aIl4+o4CIhEbMdQ8XLsV
Dy1iIXcgZB2yuJ+6HQS2xTj25jA2I1hPksQV/KFTSHSDBuA1mI6C+eg9pVSvsUK2
+QV3IK7LBc7hdA0Ps+2kd8VSbhW+a7cMofPHXKgeqgv49YZ+xjJwuFs/DBzcocMR
cfDF7F1VdSz09V5jTeVImHLbx+PEl5q15rGgml0BdZUveTIDqrEenX2ft0nAfaKn
0gBq1VwYod6/RCfAjCIlPgyB7LR2SAYgw7p/bw1nasTLVdRmyF/zU8IRipU2ptYP
gxM01FwFMQvw+AWcZf+Uh2aw75xkv4dYgxquIs8p8wLHHcuhJzHXkFgZlBkWAAXP
yjfT1lmGnl1SKQy8l4qKR16KHnB6HaucUJQiawIKUafNwUpTMYBpIq4bGrYDK7ce
37db7GG1cfiUTdQ8wCXVvB2lpeRuRT0hgG2Uin23cE1ZtDXiMNvFlmneH79mEdJ3
14iQyuf/dLtiNnJB3EAuFuyTdKFnfIN7ViwU7oUmwp6M9viz8BQ1BdJshrSO5woR
o529PLWlVI9fPaCmWJWdaVmDnJBpcIFN17Hn+wHTKG3xjKY6YuexkysIsK2Y1LhI
d+4OQdAwg/RwEdxeF0ZOAakyLrf7mF8R+6GGpYc9lDpadW/jTNcLD+aRpmIXeAJY
3J5CK85uSQjRFn0awG2W68F4PcsQ4oS/ypHBPbsDYhsrdJnW5SbRHzJ927HqJxLM
dx3d4ODTE5cXBPRggI5IRqx2kI3LRwU/rhPFSjPlaoGB+S0Rw5ynQIjUPKNS1Jd7
jgKiJILRvd2+2SmgPJXmOGhHhIn17TxASaU6yt1x3/aXaR93iodj//mX1l91khy6
P8+uAQPosbescEJWoW33AB8/1mDUz+xlSYtM95GgWiOLUGw2KHg8k+r2tPb+PK9z
io6c2Ti7PjVDMjeG/MYsFNjQ8TkYeu6dg4IbVLnMPkJZL6yd0AWAVyL/4LBzQQzK
s6U19nfQlun6NzFsMixbJt0w4WWJsVRrbpQTfYUS+n5/efnnJUaupyi2ODuuKdVO
3wUQNeIqu/S5brFX1JWA/u/8Mzz/ZZ0vCYZ/rGRxql7fdEUZct71kwP8fyZ4wVfp
rbzblcdrhYXty9fdiihLFwpWzOqCYyDQEe5V3mbzI+1DVGEbvJfale76QMstWajC
bdp31hd9Apu62OKZ4QwmKh2/en7x30IXqc8PJTQxS67MKr/QsIKfWSWosEkyxtN6
W1CVH6xiqobAIiQ8O9Q21TkPJ6CPByeh4DUNJqlXt0fK4yFXKrt0sDMP3hhtp66U
WRn163CifATU8BgAXPki+k8McsB1z+OyGCsGMMNoGLISHsp6f4D9sAT0uRQFEtcT
RF5OtLQDqHp/2PRIraIl1emWss/PuxG7LTYsCYY4I20kYBCW5XjS4sqaRFMmUu8o
MDxeo/g3N22TcXoIQTnKTWz+xqdOku1axsns9yzUSrbY0igaNZJM9hU8xnl/p4wH
zIvTnh3NJn5/9kF1XnE3YLqOlHWo3pV4RZkEnjjPFUBPMop66aKIMv7MmUCGwZ+y
5lkPnRJpfdeQfcRaTLT4alk448gLf7NX2z+6oaI18rEnE1Lk74WyZgCfMGjBVZWh
LGVotOECCv+TFVa442nJIRUG2AxRVdhkOIupWFjv3w0n/jBabyNoPBE2tFHXBPI7
mFeu8vk9KTBgNfa7xYM+yuCQsazpoTZ4stFo60kD1vFtXXFI9cIzkUBwEMEN7gFW
WChoxRmiUtk/RUooGa0HEAy7PfGjzr1RGjlJFKYgPHhqaMkK1lnj7rtj8uiveuN+
3VG1hmqgV5lsr5N+O8q8rEi6vwxLH+FpcJNSYKM99laPmfsJfljvPjSmuEEMDSBK
0IDYx9G8M1coELQD7k8L+qsDUsIL/XV1jEfx/r+gt878KvR10CV/juPYxx6lKgL4
eBgK02kWiWwfrJOk+Fp/oxmejus0eJyid5EBFNerz93gjmICiNyDglBhrzHaEx8G
l1dTj+i01j493UC3xzetA7+kIAB2libg0deuteyKqRqLJNYd/wty9GBlX0DbVxaR
A05iPo3bmOiOjC7y7vuhIIuf4FV/7QavgM8PaZlOJwy2q6dxe6jnKwyJlk9hQMc/
OxEqvdaNGd1NJ7Wmtf9yZQosPDPgvLAiu2bxzhmyPiOrFq/6x2QYXowSsd/Q43h1
Bhpvs2/KNlWIzAeH4WSRuOjjWjU21zFN2AtttIo5kjGduAuaFey4+5xV9xN2ph5H
F7opWLNY1awB51uP3tbGwT64lhaoi8XSi5Bsf1bWcO1++Pn89laTO0hghQkgEtNJ
AfUgsCSbymmryTHsNItuIuJL0qwuWscD7hZNXcmGATIJXhSIR93IGQrC40gPkABB
15Low2saqYQ39d88G5SBlYn/vvzCOvsTr1M+IL5b1RAzTGBXQdRbrEf8D5Meb9sZ
NnNTFaUGDaZWrz8FN/cA+K2L71wPMoqbse9CwVpODTghEMdKp6swqlA/wXFk3lWT
g0XkW5JeA84J5KCRG7/fH771aYID0RsRDZK09SYkX/hBkLYLAy0Mby1eOpC+qG8t
zCiNCPY2PcdWVEoHhbuB1M7TTL3jdoGkJQ3nSVLC1BrOX7O0Yke4eAPoe5E+lvWj
lNYJCxe+WE08k2IaCyB9eNxOA3BMbXB8XyJGE8IQbN+b+/RjTrQC3oso3nzcNZJr
nBOS02VuFbM8BF/B6HnP2sVL/N6oF0ehwlhiv3Ow+DQ2RZKM9RuIio8yyuRSeIy1
es4OH+Zgle1Wwt0VKiQN35Med2SCaf1hT94vbkclHDZTiHp0MhMitRC1rm7mFOSH
SOnQmKKeZs0jiSnYEhfKu/LhLI+mnT5lj3bwzrtH8SjeUheqbz7n4fVbh+AqZkgb
LNg7nnvH0tnycZdwgt5aCd+dwIdhDDwvmftcbbh5x5EJq3s9CrUeuTwHARRXdYow
CyufUlKlg85TxhlAZ5LA+7Rg69q3QidAMO7668VUxbZKlTnaB9xJ3R2CAeZzAbaW
TE1UqvbUxlV5DYQL0jC56fibOWJ0AwuA4BktJ/JP38m/2k7QXvbnDDdEjTYHrngx
+uel4oaEcNHOu5HohgBRlpaJhq9iwhTgEi2SS/1Kry+hh4IgSYK6Mx3OCFfx1F63
o7TRlnR+rYJJoMNETsn3B3vuJ9waWuutzAS/oqWLiEqN2KvikD+vIkXF8ReKDAMk
Y5dQ0xnDWw8jPlnREGTcMH2evRMe52kZik88WuKO5fD7xRspHNsCyGed9Al2OS3h
2YqG3zY1eGzQ9CjTUQMJBCNvOnHTovkrdc0N6pL7id3lxkUD+0xxHOUQfJ3qs9g0
HqdUlFx+jJcXXNH1ZVBTaDvhxU5Doz0hWohhOK+B1t59ag3kbD1oVNRL3Ov66MVz
cWLBWE/5M8+En6PvMWZAnxG0zvov4T3SSF/oVW9A6JoJSwPahhNElXZrcHBefkJd
TtypT/HV3S97fQ7CbuCJNTX8YVROP1aIFUgviRjNCfH6/GLNHOh3L7AcYWCK61o7
A6FyhQG2GOO33sYjnjJ29xHnKTpRjrdDEtzHrR4rIbORrF/OpLlNCMX9v+DwlTNc
lKbDM01Tti/PfY8I6EZ+Fly4ZipoCCKtt79mEgJ1GNWkoY4/xqFLMgt0ByFAlw09
6Q4b89+SVOYieqzgXWNeHlDD8fdp1PjnhIPsDqEHbCSCZNNWNzyfqGnZEYVVsX9+
jBsY9vBjKq0uXZLCrDP3T11ePdtca37YDSKcWPydPDRl9UcZneRuRUGJcvYSFcaC
IdPU2N5FxfSTJEBTw8KAO2INraWOvI9gIu6CSKfpR2gZRgVovCSsEj91rGW9hDZf
tuq7+a7J/xiw1oItjk0Hrmo1o0C8B3ycCX/eRXSquNR186k1o08z7bjB5jWo769g
+SweAkSc206YrFccsvylTsC5mq2oRLbZuE4FcLNcyTo3pt/K24GSbL9MdLqOZ36s
ckq/IwN8nYShRh0XibBx6P24CdNk48rm8+F9QK2MvnkvDyVOyc+Kt9HBpXeflNQ4
+A6Xvy0DuwMjXKf+anTy09Xgq9651CJqdfbASL0M9n4dQnfjb2v0v9OKly/5VsOl
/MuTe2pjxLI4GGsMq26JSrFJzjHLJBT54FNRfl5lSYo1WzNPHNiFwvi/Z1m3V6cp
NyGjGv4f7eFXl9uSUx+cdCsVN+AP0R6wV5o9XgrQWpWQKqPTrBJPjfg0jt0fwDw6
F2OomjytG4ShA5wA7IReZSqEukc0MZMGtglBXvtYEj+x//SrWm85FwaV3X1jOJ5j
7Sb/Cj90qWWC01l8ZCBl0/9zo3SzZLPDCE32zKJlc2xm4LK49DjHUdqeds/dCOhO
KKZMIqKE8Kh3zZ+FI8CRtUJ2XyQtGAgoeawpmTa353nz1b3Jg8jQjJnvIekMmhhN
st01B2SHoj1YZB0xbrkoj8bvfAGJCL9Ys9hZQp5wwkgNe+WbSyQn4RwrYhmW4DLj
TOz9coO2l/jxBRvANNsHoV4rNdYgjFbN0S802LiPqi+RskVNn/zcQze30h8Xkd3Q
osBvc//XneG87SwcaNAXSe7RlYegmKgv1wAN8VD/FLU+bZ/6zUfyg2MSKOOySNsh
XxG8CaoDQrT1T+i32Xp+E9a6exHZf6aWNvfXwvMuxk3kTxZByvncbtX6zctO0B47
8XGa+0NMQ9vtPATXrkX5VSoCW7f8gsAeFIUBWMvmjt8FvjLT/EtSAMij0AhGXVYK
4LECLeZq79hJdPNw5S4SNCibK7h4bzQ77unMLQUNR2w7z+PDi8B/GZPEPESNvHJJ
l1fEDgF35xskqgFBEYBr/HEY8/Wep+l/xCXDU2fq6/ALPvvq4WbyaOiMDBOj3ZiL
S5+s4Ovr056+hmondVaxa3qSiJp+mgIAtZgsAL28lGQuRZv/M304SftSMcuzgl/0
ZSdPawPrF/put3+xMEqyJXtZ4OYuXR1K4/jWyx5FTY845F10gIDYuxSh7R1ALjFd
9QH2JKNDPa5ttB3WYFlrDTcaLnKW1eri2P5Xua/NneZzkl3ezKkKtjaW0ybSGnoI
kwiYmNgkO4qOY1OB8o67Rh6+nLBnyzhmVCe/zatT5Onwq62jnaQ1uwCmjJgnPXL3
Vxyvhrfn80f45BFFiI7Xzw7jeP+Y1ah6dMl5vZlNxUjvmngDchdYR4jRqaPlL7ck
Wl6B5nwMF9o7GE2hq3RtIqPk64XQiuXM4MwbwT2BCeL7FGR7Hz496WOFtZRDYZsg
IqMc4slKETFC8nf3VM4rJWgn8GpuBDShOBXycV+lrxOv2xfcZ8LFDKSZr4t7idp8
x7Z7zGKEfT+s9hFGM5/Bj349yI2HTQ+n1ceDB5/684DY4CPbpIhq9eZ/7zF7M3xO
NQ4dRYgHEjG+K2hS+pd/9ujl6WX2aqaGpvn8E00j0gd0RS2tZf8oZzRCtED31HfY
V6XcxZhe+f41iDhNL93as5mRSkTk9iRBOLQyBwc0TEpvC6HC3FP+PhxzP5YqZaMp
EnhIvdq/mS8se/MoQ+4OJJ4/yh847KQtSRbfnDBbFFkrm/HrKyHUe4IdF7i1+1YZ
WfQYmncketJSDUDodUiSoMwYP8SNiYQe7I5Pc7xu7RdaXvwFYMmhpYSZuYaO7wcj
UPvmls19VSq1XnSPNmx9sT50RmkFa+F3dsdGx0qW2AkqmAg0ZuxoFi4OaFDhWVOQ
Ns2Pr1lnZP2l+y9ouEv/5ME4bkeKhC7DTAtwHF8cbwmKXM2n07sj0DySYEK42CM2
w6tx5k9WfMa8BKEkBgMzhItobZSrBcRicVoeECPO2VpL3zx2//mPpQGMSyzjwzAl
DX7UXIPLmpq/Afq9LH9OrW4R58txb+dEQQSIMfHwMK+oOI5i3XyrNkPjJV1ePpm+
YihObdO3eX9K8bMTbDdH/mb1/74rGK/OidI3KqhMIx370qbYybARky68EgsGC4zj
D566URCK6P0ygTFrjqCAlTGR2XuNh8nL4rVIa1531oOk14PmnwyKqt01sl/nJqbz
6u6Dve7KZNP4unBQR+7+hDWTuDtT5ZgmmJBDJlYwJETrr3F8OBYHibxPzWeeVBI4
8DzWLDQJdCpGctAC18ukJ26M3WUn14IViLdslosHHbKESjlhfwwGg3eQZznLx5FU
Bk2XEsSO/+GhE4Ent/dk9G+0jXUpBoGR6SPJ/FucbmaYWhnTjxQXtRdiwAyl3JZX
Jqfrrk840VI2GOzipqzdlgULE2E++RyVavhXAbIOtV0jRAa9HtNb3jvC9ZOVifx0
JZTsm9+RI/XNALgZC3iYoC0opj57JFlXFWZzfiFisDRfFxTRvF4+SfrAGU93i8jU
zcfBlW1TBcmPiphP4F/pklohElAzbnGjyamWrjsOhVc58KMKJ8kDJTmSZdFh26k3
9A9XQU0OW4PKwACpXsdWP2WkIbxNccAeTMD1Pea34o968oVcMogQCFSZRnVF7PcY
gSOIp7gxDetSJZnrfKbCfufuuQ40Vh3xBISTJJGXlKjg2zNXbnVEKTJjBAiCRtaE
BRZbJNSxuZWMCxLggLCZGwHnY2oe6sPE+rVWO46GoWdV2+T8/wx2HSFHZVMzE9Kf
YHW8hO2ujhHKQZDohkMTR/fWnR/pq8/tAhwhqNTguRj7RE/PMQS0gVFbha/ei4+L
wWvo+JWnHjIp6OCp5yspzkeZQ1YrkG35e6xy8sWEdFtE3M4873NYx2HP+o4hKO9x
Z1jbDRA4OOY0QnLjnATIr2+uUZFTVi8tGO47h+cuSl3imVTN4u9fXaHGrdjfVSug
3mARL0GdC/8Z/wplj01tEh67iKpb4p1FhhfVEbo4WR9SUpyPrY45B3E1uPBxTGVK
Pv0WogL0OhHS6f0HI0WEuvr37vF9KzRQWzoatZvhqxhqUwYkGVV9HcqbZUQj0cuP
2fBThiXBMp21a1cYR8KqefGUaSx3KLK2U5dSX2wQqeluROOSwOLeo//e1pvDUGOV
wbca/GV/9DRvexLKr35mPx4DGj6m2yVypzD8H/Mef7Km2i66woU7XmzS7PWpf6hY
oGru8lZRpneJ6iNlZ3Co10oLP5PqPK6K8E+zG8A5ucVzj1U/9HgYOBAgfcNbQdC9
aRvMKKneWD6HSpoNkiwYHcWwmsrMUcNU5dnh/EpCItia8Ia/qqnkRbBK6afUVP3c
88rvC82Pa/lNcVTkkHK1OCfA4gynZJOT3sCz6M5d/7pm0oDk184u+ibEPDkqBHWF
VWQDNpAIflaYZmfC1LssS7HSayJXJOtQZaE23mE532SZylCuR352pNv+v4oMA33x
h5sz1ez9z64aqXu+cuzTeGybxPCZxVtxOgNXG971L10mUlmUi2SXX1FtFvRenbZC
6mVkzVBde/kYRZ5psW7NAodQ8KW47Kj0zCpQvE/XkhHh7dPhvljM68sR7Oqrg652
QBsWuVdYXNWSCgYWgWu1+Uy6Ap+SJSCpCoBTwsItIiQ0mUrCkvnrcxDz9VI64P+W
CzRctVKvMI77KKskPK14V9+X5x/UP+C77rR0DKu8/7+0CfXnimT6U7XnnUh8nj/u
uhAPoP2JEnBNXd8zuR0KGmWre1GA8N5bzMp45+DaP/mwu2s9RpY86jyEVRg3cmrO
PWgGQ5OQu58hbddQIibSjJ9Cq99doOauOWR5GZRvSLaeyVs9U3UlJA90REBzg32q
uQ+djdcbh49ji1Jj59v6UdguNLzBNId5nAMiTv9Jsuw/1r8DevcGa6zv7YhiJ1AR
gK56ZZ1sBVvI8uSygY+6MiP3xFqUS4nHXHOc+RPBWWd0kUZTLtgDQpmIpLJRNVp7
OHRWhUb22rumKKrXkKUroGdiDQRLuHvRg1Me29cE5Ib/ZfwaWvVtHi/MWq2omzBV
143q4tZCQplLNDTwtZbmRCSO2/fijCtgnwyyiWo+afGagFagZU9wdMYPNZUROkDF
gsLVt3Zk8i7Zv3xo5dizugeL/MYgyiirkxuAQwqEfYWzmvkVonUAo8Ggv9BFcvzE
oHEe6DpIWoeM0dRRQZa0lYlAcNlD+uTL12w7SKHJeK564AlgBXxC2TR20YdJ4K5K
B/HvL0EH2Hbe0U9KPcSEhjhmPtIIX1YWqnn6NRw7SO2TAowOpx7Dxf0ViIFFBTPe
/UNhDjb9afB9P81TrrYWYgCsFMxughN3OugkUX2XCtp7Zx1X7euzTEuyS3vlV4OT
+D4HH9ZnQ1ArzWII522Sn4ugHNRxIrxUnO0xCV/Ymi6Dd2bIlzL7tX/aU8MAInnQ
8+y9MBMuMjOpfsHtMkPWGII+yedpw4ov2dtsl9kRtuQBLVaNISQcfG08kpDlpmKb
Dp93AiosywIqk6ED8xhRTFJ7bLofmEXBft+5daKkzV40ZEiHsh1h9WptdA9unH5S
EnRDvlhuId8it6hjs0JS44jMWmSKLJh64zj/RnCW3w9MZdc5Xvx9gRzVr2W41TrH
C1mV/LGdLvDs8dg3VVRAxOW10pgI9Jf0tdEHYpNnV7kNkaSkIocKF7k5sjyEg1lv
F3RmqBp9Xz4KGlRBRl7EpY7In2ISDK2GYFO/371FpgOekvozjftKb2QSyqCD4ZwJ
Ik2kSzhF+XNumg+xPM8A4ZzwY4M/9foiNbZQM1YplY/6De5onuUmF/1KiptCohzA
i1OyFr5V1KXVO29jmOfXHKg/Ed3wHUW06AfViWtzXCTHfTupBb2GtmkXEhHKo0bR
VRTec7cE8K0Y+6lV4Z+9iyomfiCJ4vioywfQKO/ZbkOevXJITQ8S+StDULbaIXeh
+CqbqAZPe3wUgdAotWZ3nXiG1FjOdVohqwcx6LemGsC8BtT1COex6rUA4xOPjJqD
u3/vl4svsg4BKJx/5qqHewEhvGGooVaP1hbV4vQD6zeSnFxGSBm/zLL1fb+9G9yT
YHlL4zeH/tf1pORujF7YNvVxGyii8b9cg7F6MsGCtMvL/8K5yKe9uD5PxysdFa1b
0R4NXZnWgqj/p0YE4erEZ5oIE/234jc+gWzHTuH899+y99nRvjaCZiJZwRJN1EWS
yXde7Bal7i/BjN7sOl/VrHLQ2HbmMmyu3whLqD/1jxQrzwN7cf4JR9+iodjkJ7Gv
DvEevmSl7lt8qY0Z27Djox1Ntjfk2Serdesf97XrfQY3XDEx++/NCBLNPL/QYXHJ
X/0JDKt+6JLnADh3TKlWEdGXZruXrWeXnVVJAI8ILwAgAqnRuJqXEkB7YAnC270q
asbd3Rqg2qVS3O7Z7ILHhWTaKfg2FehHVou5IrFPJz4Ddmv/r+i/dVEGhawJHboV
CUfQID6X3cPn6mHAnhs7yVNOZypUk1TEBhR/6ZLK/FJKhwMq9oEy34uU+YBZ+PNd
PYfofb1BdDQqQgEbSn0mXU8AdPwX/U7o2LmsPfPW4PPlnPeNIld1RkcLWo9hAaet
bvyuH6YhcLFR0JaQDecb9yf9Q2qQruiAUOvd3yfeRjaZLFWeQVWHQGzeA/YrGPDa
aqJOKHx9nNRnwWmPPUASCYulXcGG0pNd6zBEDZtYtgJoUHcdytI0aGtv1JvVFckp
QBpTNtQNadkaxQLPJc0FlSq4+REkithBXeHM0vzJf0U8vwUZjspXrOB1GRZFZMl7
jNkfh2/2YYr6yW9gYKPi1bRo9R81P/fX6QZxosocdh7cPh0hxSLLGFfRM5tkj4aE
/f1lEokUNuH69spU2LoTXkFX+q+LlTjZVsGwOAgNrS9sZGIIacCgZicShYkXujG0
HuGjYPNpGqUUIlR3B1AmV57nQe7xUICG4h2RZmU9i/Ey67Z6/SRk+4KMnkrVk/FD
5lsQ4nAe7wD0eb3/h5qt4AJ7cTAH34R+43VvL6zTer4dLHndB3Lbyn/nbQngExIK
1WSr1IPc+Uw8XnNScyKnGls2Itc6Bd8n6PgYf1uxoFdJebEqRI/gxGBA1XULOOAi
b7KKSGB9uudRYgNoHzXDs8Nj4g9Ufdl90j3JTxEkZdohT+EH5ypTFpzG93dkSda5
O8FrK5/UHiKO2mylC0CJhmzK5Y2090cTQPJa3ZP8G3WQC5vwa/hCpIKDbBTe773z
ItutyYPPZOx0vafHHCw68MVtCQueZypNOvlpwHiLrWlYjd816jSokrm4XiCM9FWh
6X6c9a9/3OAxY29k0nuQA6fjvnWipWe8YzySoXM4A3ptUJLLu/pw914MtIXeKwCw
6CuTNTt4FgtyqSK5sPOcslNe4Cv76oSULEh5sibp4NeFYOmAxqN8OUGWLiAAh2+j
TfMmDjzRYsefcIquzK8N4f6zgQtgIRucS37sAgi4hkakxomPcjsL5oaigrzc2+Nk
CQi9Mj73lxaCKXr+sj0QgXgbhgKQvW9RMu11fGJitkT1E0oB3RtStQbWvzPqdxUV
gat3J64qgUoCPtP8BGAgEcnOGNRw+kIQDZX/NiY5xf7SqKVBuFaL8DgiJ5pIqZS3
PlFjt6yFvcgCWPH7VP8dfr4o3tPIKMA0ldMtMyXG+tZik4boQ/zsudDQZDSsswkY
Q5V5RLHEmL99udLcWMufnqMn54e7E9HQlCgc+UjfW33HXvF4K3QV1jWALRaAhaYV
/yKgWR6biXgFEcw2no8JqjYhKc8fX7YYrqOGGBDIYctXR6ydtC4JT8hGbq8f/CvV
rUfYx0DVgPjMJF4Ig9SzFiADx/tzD9sathODk5OXRVJ752AyNteOGEPjSlq2vozu
ZP4O6mnuTCLK/gtBggVfvEn9Z8SuZMnBZGy3U1dnECPB6F4AxqlHPt1J8YOmF6pl
VVGmVbHCWNegIrMKsrrYlqQVCoHcCvKP1XJ85pUj0dSuUPe5E3BV5yh+8Viav/+o
qXoVXRyR9CWRVNwqMhqPBT1v5QKViWDmu0BAf7N0h/fmeFkteT2I2DIHfLcoLM07
QMe8lHM4tDmEB6UCYfj9Ai7QA0shb02st3A1/7MhkfB7aUCloSJOWb1o5xD78frQ
XF2w0uA37V9VQECmFzr47rIFCNVCY+EvoCZku5LHsxBAbHx50OsRuwB6ZDPqur28
CZTdYJOJMySMB+A8RxctvfSsYuu7HRITWPHqc2xhmNp+2eC+2RXaW8DHR1UpVIgJ
mp9BGebXggsVPkq+PI8+dnhljr9gCE7JEOZ4t9BjSZfKD8Gp8F1Ce9Epg9sofHks
ZMxb2xu61i/6X1NilSSv9osR4O0HLPnud/96I51o7Sxr0EFV4zAwQKxsUv0+oers
/gqXqyfrJIS8b8CYORKgb8+dNuNWD620zM7LNRueZUKWOkiTdTXamat0OL/kNJmQ
2HBJE8rB9JgGZtyxf5SjlQcPoiRIx2Zd7iGpi/oSayA9npHKKqZijOIZ7wRwoRjy
SivRcNc1u1ELoukjrlVUIHzTZxsKyu/V39cdiEZma/kQdDfyog4wJdrTwmZtvpkL
yGAL04vdekwW/vgLXXuezWZUzc5TCQFvhq+IN0GtliVEv6oKaPuCMj5C3o9Fey/H
OEGD2sKFS5bvkUiio8n9NfSr0S4XQGS9Ot6yAuDGcU+Tnd0onBjXTVKRnZQ0Pby5
zLf2E+zqyxZFLQrfDHnYjUm+5jmn4F7Ocv3MZ7rnJPzplv6PMSUm1jUC5+R1KZ6N
Uxt7CmG+v22vmgINrnCVib0Hkvw9zIx+1o4XF3yKSghZDOga7xuaDK1eaKkos7NW
kW21M6fWbpW3kNXGecdRLBFffD4ldmdwaD/ds2ulp01HLQ6eOVKoHLG3hcBJ7Xo1
rCHwyuzo9Lfsd5FO3inBsy/4IPn5jwvsfqHYlIdIeYayQ4XConRr/sVMDk8/DvcN
b/pYhBZFZ6kS8yeupM8D5F+LAtH54DpnO1YsVSTHLQPL80yrmrhmZy2CG3z0YOkR
GQ1tD44kPDgcLt/vEScYMaLtBCmmTxinNoh1lBiorIgOGs1yv86NCS6pTamrfE2j
BSgFKrufEmdsp2T1FLqe9CtB2tDKLO1zolFEt8F3iUWE4ffResbKjfWXPdRNmlBs
WlFZd7NXtNgRm4jMvlrb+cf4vXu9rgSMVA1PofqSiiNTcW9e2Y8lrSlQi/rQJmOy
crYQowJvghu+hB0uYfoQb2YQcTDx1guQlgHvi66QH3VilYdp4oqc7JVRQt7LWi28
bpNDxTuJq59x83GFZGQbx2RRuexr+ldh/Vq8qNmge67XxL/lqZCDHTrNoiGiF9KB
BQge6s52DO9GBPVAN9YlNY8/BY/xl7mEuVGTdEHIeVFIjoz2JnGeW5Z6EUfb5jnE
TwQJxI2Y3dKBn7rPOe9vfcPcNvHF9sz74Aerw6wRfyDI4RopEs3O+8ZEo9k0sJ3p
Zg+KrsEEkYq1IwF5xewU9Rmwh5wBMPdhW+fOfJw3EJ9qWa4O6lgGOlgAIrAoRrsz
wqDI4p7cMXmFkStux99Ky/jUh/Kut8hqM5PrUyO8lEfyXIvDfG8bmupbYrl5BF3F
eZTe/8XBIvenPkF44IAwYXIKG0xbt7jyfz6JIShC2PTFO0TCMf92WylMC/gUc8Uq
KgaK55KJPrSKia8PHelr5BK4vw+FYKpey0xpq8HU5lYb/v+99xzq0qCY4mk3qnZS
4RkqKJYrB4emV0qTkxognWarFQeDzRu25om9HkVXgXTNcZ2nQt1Jp/hUpqDyZ4BO
N/GnrY8vrvPubtd9ODXzleZDcjW+IwEJIbRIP06M5xrmXU90byLPd9k6pUBKvoWi
SzefJsxqFPnL2ZvCkbZykC9lGns1iIsZ3LsmtGT63vX6jcwEddjlJkIy8KV47pEE
uc4JospAjGFugp8amWyKVJXM5VVsyx5F97m50YiFxdacz912Fc1okmb9EZvyYaHV
r49eSvhFhzfscO1fZhzqaPygyDO60Xiapn/vM9Afd15GjL8sWK1B8ann1m73A2kB
u2mW45PHnXUjl+7ED2QBIJC0AhAlT2/j3dIS0MXOm9kMO7fVemt+dNM7IaDBCKtr
cWDEtAyHoy/GQ43Vyvfluo4xVm/qG7nzWHYvn4uZ5HIi8NXYk9eplpLwRprqYLUr
dZt9YHISw2O2pn+ITbF1FPnoInUM5tWE5Ya4TpAOFEHiNq5JW7Jq7xFJ/tlvJGgd
/O9ZLHfLiYIbgJUcwc7vGUxsWZCHy07WqiXs2v5J7fJT1Qpb7m3n5MyJ/VlKBtiR
K3k5vYZtCCQDIwB3FNeBDEbrs78KLndij5n39JpHXfUrBpbfpsRsHCsnXTfGXPqc
gpaHF8EeJBpCjqLTWfM8tw2AVquWDqHFW8ss3oKKq9QS6JK+FHV1IIVzo+gllLsV
rgFWlHUZLZk/Ohq4KmUTdE44GxILgdiRHJuaop0j+fCDYZHoccLpyOX7jZBPeakp
Hjuunvz11S2WqKqef3II7YY4IT6/wdFcRuZIpp+WeGuPxfaLkn9xl6vWAKBdQqFg
wHX9/aYgX7PP4ApaPU0qA/Es5SXOdzr3U82g8CqupEKRWb6wkqRKvl7bxgC3umrp
DdJy/XeIr2FIaNrLMjzGox5M7rYXA1AFLsdlKY9w5SRjsBZexpnF4JM6uoNPsI63
/nIyBqLzbzvXQGjX+Z1A8GWesnrAfc/zNFcd60NvZ8cx/AsDoSqP7N7QBNh/Z6YZ
jpjRZNNxdjdSEB03eQNs9mPnq6J+ZthcCfS7aRaRQUr/rW2dg8JD5+CA0GROWuBP
MY4uVvl1v7Unob5zojjslpZBdNI0nwWz0lfRgh7LfaUWEwn3YnkkPWw9mDuTa5A+
7w3PgAja8P/nkIw1X23oHx21Ynt5rMd1cGpRt/swQTAKAtr7F0qz8co2u9Ma9PS/
PZwcr+qZGZCYw1P8THEK/Z0ObW3YjfsCgcGXd+N0Y2qKxobVkdnxC5RSZaDj3HbQ
C3F2Gt8OoAWEmg994Rx+CmRXLKhMLLWW6VAuqWEGjT7gKi59HRw+WnWuOjf1WO/k
ZH+WjOzdLzbx41nHgNajf/xGkh6XfnwDVkejTLZBRtpLz8E3VNhs47fpUOyqAq+H
XiIzIgNegyG/RJWEPpeevLaQSwibtJqZouWzf25UeBS9qk3sLtdqFrXD1fauPozT
HyrMn1/Cbr4ixBRA/IetXAKrlcaA4oRmJP/YtdwKJUrZuamON/fHznbQOLiVZdJA
zP2NopHIFvh6+OnJJ6Wa1WUC5czVDIL4Q6V+wz7cRvABZ/+Ekk8D4obpruXachJO
R/uoh89z1lnBlPz0mP4vD6ABipKMi+JFU8o1drT69A3ZMpTVpI+h9SFV/amww5wd
73D4IW19mCaI/2r8200C6pdgTUs2B7PpDg/oG97yDiIloUT+wrYNecJyCdQqBK47
pdayO6wS7+XwZg8O5vnnSzrxfZOkrBLUBSB15VNcZjT6r8spkZlcqycGKwfpG4R/
Eib7lBLJFqsgnFZrBjclvQ48uuN2Ebo9f7vk+X1ckaUgxBy8Is8/5KUow5bEt5uy
jaV1Fl1uhlJBuQUVld2Dq+Zxe1Jw9J0rZP+fxshrvldrZdccXqQhGtTSbugViiWu
Tm/T4bILxyKRTkWUcrawwLsiI2wSxBL32zNXeQVCRXK+CueSwP3Pg29y3PmIwM/V
EV29MSDLTpXalsR3/Yoq1jk+6g4UMFJO5zLOVmMsp9YJ4sdaCFJhuyhDLKsmnaEC
HLlerNzdkiz/mi4jFyVAsXaNp4VBZHj/HiJtCFMvV7PzpuvNKkSoVrEX+ao2l3bH
eQ6wEbK6gLbsC/011yRzjf5f4IFB5PglsLn63zGCte3gOIJ1S9kByU39eNnfAErJ
qi5GVdVvKlAN4BILd1X+eWt8w4Wm6+aWkRLD1uCFx2SuRboIRc2DwDR9Jc1EwB5e
h30rL8TmySa+OsU6O8wiZn9oq8tGCptZLRV2pCLUfc02L5cx7E5KDn++gTmSn1GU
AJezXO3tyMNaf+XniXbI0WglfsctnfvvFZUSlVYNcauMunwBdhGIlvV6O9hiAnUW
zTIXxth5IPuR3DZjIcY5O5Uc4er6W9IKGSVLDCBg5n6HtrcGhggLNp7qf0Ho9FLa
jJSPci3vCo9FcFElBFyR7PGbUDp0R0hX1h9Mci4f6eV16kXHOlAI5zjJx/hhtG7i
4Z0ZYYzOhf2vchYvsTo7Whv3EbnaZ2zssX+/s8/QZ0wnX7fYSNF7RRBFK5OHH/3O
lIym9M0jJ9rsCSkLrKLK2q/uHCVhK9qXCJmeLzXQucHFFO2k8xuShp1VJJtqIOOH
F0zEWU+8pulTinNZrlPkf7YOMGB3vjCiyv9+dSvI+ZtNCbryB5gCqtlp5eUkQLSv
xBIWS3hR83wbQOQQOC9ci8cr5zR+LOBtzjJNDvS1qZM3BvGGVBtH6VXBeP2ulk7M
/SaKAw9RCX3W2faHul6dQpluEdWLRbTmtvaFNDO5c6GUs2l/T2TXicn6/e64xZzS
cnZnga5TFlCOQm12d1Im5TKEXrOvqWOH/sHbeP1eb2uPKsrP2cn8J31YIDO+JO4O
0vsjKZOr0Pz15TOEVQ5PkOFFFKuYDihVgSlgtFhbKNWl0YjvkWLLD5eAa0sO+jBB
c37DG/VSctHPVKgZpgRiisZpCzycTNZUggv4OwA/Age7KHqY26JKX22KGi08l73i
cV9IyFGvjMQB8eIB32I5bo2mQ3LeNN3hpEDD0wz+ovXzEOtZu/CQ1wJdVYz0DGih
zjwW/M+VtAs6y1EK+xzhlHAdffRrccmyRDn4Gz/aW90X/V+SMshYnSX6v7nQJqSM
OIbq1sEgjhhWYU5vneXXf/FDLrR5OFDp5u8j3h5sS6gSkoxTipUAEMMEa8+QUDs8
vIVikMe7iZXftEzldrFIUfY7vw24Y9Ujiha09qG2dYdpkeiGqrPOD7OnwV5vmWux
mtaK0yOUzyqBtpLfHk73qMebwsWhc2tD1oLScUIIQUKvNODWLIkQ15qdd3EWBvIi
inlwyrqUIem20AeungejDFf+cvNJnnLMRPk72bJG2NS71a5gTeZzs3ld+ttp96hw
YtPRCYQoaSj/lero7FHQNr1YUYxYfU5o9nVYR1Cq7OGp4ft+2RuRjRi1l/Ncg77G
W+Y5tAGmSEJo3vRdTBtw+WnfsKaJl37Ng6D0WUpsHToa+MNP3uDvQlP4y3jAhPvH
chxwIAs09sKErZRWaoAjOxarVEfVyBPbwHuv7oC1Xz9QCWI8qnYi/OHd5nF3sC8U
LTi3TEijvvhpVSE5Rf6kLA2jnMKVDKAAojFCyJ7V7o4KM/SWC+FAb/gTeQAk0bT4
NShsQAf/xrjsLWoH5fLpMj+/5ocHAiCtrFFDCYtJ+HJ7rEsyfA59hm5iOUrHrLjl
u9AUuTq5kwjYrX9CL0K2Qh32u0s70pvDheK2bVXRLTizn7goRWYHNc6A5H4GJdC8
94I4RRVE4jBtORoEPxSs1wXw4CqtKEXilVVhrCDSJEg8J4XWkJCGDarUkliQHzgd
2FLezkuKjMhcW/J0dB7+vmFuCqNK347yEXBRi5ZyChPk2Lm0ARJbSYE7BmWA+kVO
vGL56svcUXhr7B+IVkVP9h8/jUTrkQ51Pns+v7tv8BpnYpA6pNzgfOSoE9n4pEUM
+qkPEZZy6LHAhpiJCt0pYJMS+OXLo8GY7pn+X+H8nGCgdjEpllBVwpWR+avgPbdY
miaprKelzHO1hLxjRDJJl7RA2vchGBtB+AxNL4wSYBK4XqaGDpRL9TITMx3AUdY4
Wm2eB04Da1VILiCsIOakZpSTL/tV5m8E9Ic2uSkJY4/LoTqpJVWn8j+wFUnK44Zr
ZcPwwDy+i8trjeNDB1kVBkuphwMldMFR+ZBnH4XHi0LF7o57aFZ1JE+lz5e78Ti5
y/CPTYw9xoGZcSDO5MXExPGhJrjzi5dwPJMuh7m7BK9F++xmoULlpv2fz7PU6cqT
yoDHYkmZ0nMolxZ8vem56PT5fg4eEWM92Tdy05jZ6BcDPdnM0VhA7gN1CvpW6qHf
AAYCMkFcjFBHlUT7ma3eFK/dXTXuZyN+BDa2hXhdzzg4NOzVs+j4X3aXT1PSkCEp
liEF+d+tpwy74xbe+FsT9Pm3DFNnlcF0k045cSejgKtKnohR7Y1YY/Vf/+DBhGNl
owy1PMnzJ9FkmXFJ1xdqe7t2yofrGz+de5L9Xw7fQepLroofd4OG4d8QyLhaglXk
5B6jP7iIDF0BBMSVtPTnwBiMGelNrk2YmHh4iOIo+cNyI07N/TOvQ4AuJtKVYy1G
Q7bZE/+6DfGJug7z7ban3Ekqz3UFLnzQ5HRdAjsasz3pTX2cUANjdZPrA9QgFDE7
5EJf+RyblJj+2f6KUmnO51Bz0Cr0aZJBFksmls8yR/uuRqmfzCI0NiN2kIAiLVAE
ImgAs8U3RhfA8T/xrzFUBa2hJ6de3SEFn7TsyHDHWODqQCFmjBoir/KO5qDDQVuw
f/bBjRB9gaJnfvQLqoNSEVP/W3dciYHm7CzyaydAlOBu52UcJTMlZ3td8YJIlirC
rDaY2UNIBY36kyczMXHw5/sZXSQsqqiKRo58ZknmKIMyzBgDeB8ZyOkn/l8zKijV
21jzr1qD5oM99MBZOEqwgm4Mc9ABK4aXi/vzoPluNjW/FWTosTQAjobtuojBTIYY
cGgG93QlZo5phKsvUBtdtNM0AX6MU3GKXo/5UPfS9wIxoUcIWUhsWVI6E21k7OHS
prsy8K7JSRKsOeTPRYVmR3c0NueWaDJonjVQGEuB4Y7tL+SGXnfhTKcSdpSb4/6+
J+d8VajJ2+zVZmHbGNkpb2vveJk0KvhEpg4r1e7i2q7ipTkceTKeh/jQXeIZ8ZCu
b+ao09Wt9hXddezAPB4VJpq1XEuxqOtYuKtGEEM+A4uc1+gW2BoYNus/KFuQXRq2
c5FVUW/MmrH6elYnhT02hwUZr15MWdLqOgrMcfN/UJDIcqsPmcDaf1jURKKQoQva
vI9DJ/aHbcQdDRWHSOJs2At2koL0R+Hx6S20YjWcrmR4AfSbfggEu/1QJr/g/zVI
3aatB+m5PvpyC7G6ihL+ElE1TP1zuqhIl1zqOCNb4XYyR4b73pT6k9aBcBkI/lGE
UyIoMPVZIZR11qQu4KvYiZWFLjTP+bnbmsuO2c84fAebxDtYMloWIVRlaQsRzWAd
5VOQUbviRzqr26Xoxv678n7V2OjvtZtNsvzuyi/okkZqalG0k8uQm1qVC1Gju0RX
aoKygkP1LPlDneRTNkoRSNLaw50XTOeCJ/IrZ7nLGpf43gXJeV5dcIFJbm2t/lYW
QLKBoYZeXwGyaGIYMGAFnknTQcieKQLgYlrBBkV13/FK+sscTZEqQqu6F7qfP2kt
hMmFTxyxeisPmQ5ZoHE8q2ozvhXuSiOU6fZ46aNmDRCH8Sz68zs/cClmYHQMr4w7
PMqXPQWI8eIXV3v+loyuDHv9/gPHgXAxBnW5ulVB3kzm1M/kYWb/nGjJiqjr2jpa
mzZLcAq45uHhR+w9z9zMAQFtNJuayKscDEEaYmc0IvR5XGAfMZawctI6oyPbyIl2
8Z0o1c6V5Cc1pbvVPcK8pNdTawUKOhn5EEg06XEhrTKYqsyoE6bFwfWt2gcasTU/
i/rwiDQuz+ApEK+PGJRFDNlsM2IyDUnEGjzLT5CLzhiJGFOn7SRmcyDQ2Jo2nWRA
eTb0vo+61hh60UJ91T0yk17kD6Tan3McuY5uvnjkYHXe1/tdCuXWcWQ6KedaV5RP
cS5vjbVO3PCceasgwj4tDKQpo/T98bgmrRkj1zNs7Q6WM6EybzQl2mLP/PpwHX91
lAe3sRoXt1nrak942uyx3AsPfXKwjO/gZpItpN+3XdHkHuB/Sjj2tc0q4Mhzo+Z/
zwZgWK4bUTY+QYrpdwimOLfMVGS/A9c6Nz/8BXQZPUsXqN7fpsFz1evHazNv2EVT
mS977qefLgxeiAmPpdD5uaTkH0bW8aJOZhpiA+Jh/W0PUaQWEkiUBUM9iaWt3hnA
h33ux32aK6KXPsf/wKn3uMGpOVjA+tMfoVtG9+zAtqQ0reIisDhA6qLpIsUJM0Yl
H2BvPC4ZP31Yn3s8euU81DJfs4KcokfxXO0XVQ5rbspRCqAnh1J1rS1D41VK05D0
ZqhG7xM8UZPa/mm2xLBCoPjOKFY54VwDRjNxPVRLxiq9uRatF874Z4HhclvVE1j0
b92+SBjPMn1BDe7B1R919FjQ+ed2CuSkIaIYuaMUoHxcbrTr7TXzIXu9w32joWTq
rtSN4bd+opEyo8hoIAhRc498x8uxBk6l525J0vxzebOzD5cpyoYl5ZDGkuIgAfk7
0HbiZvclO+G43+ppxwQTxLArJycxnUGWo8B1IkYu2urkT1r0vTLpdNXUfglkNgKf
EFaBVw3PQfj+3feLE+3QaAapJqcCfQY2y5SX5VbLFzXfokHNkYT/12YbdlzS7QZE
UCl9FrjYg1wvmnUuPe+6oVlsH4ao7H4XrMVfKbQXJueFMT+Bs6TdjwugN0ez0/NN
ysneJDXyuvbzM0lk2vuNAlI8qC0zcTm4SNov+Trv+I91iunhHLvWoxSRziNn2Ay6
U+Y2VPr0uVQrxW6H/LFwXH6+DlzATIFWRR10GFrCv7CfgpNgXXw2cau3ipToFKOs
yT0x9rHGaAfmOG+3bVGWoAkb2V1MJol5fIe7sEbBV4G2dfJaEO4P/BgoH+iX0bzT
rpLVDGLKXOWzlPaOsgL0PUHkJgl9MJsv5uGXaA7LO7j9Gr2+U/eOWW+BF22F20Eo
sXZFtv7wfipGz9Ah08XMrj3qQ3qIWxRGG3nOiUrh9S7z6qQVAUu0l4GE2Y0T1F+l
/jIy8fInS2hUVqZNOO1LkAEEBHDI0MuGBuH0n5gp5y2YaJZN5nUUOOKECkhcryXs
clyLG/xhGjtLcSUYRqi8OpbbasMlV2BMZo5irfEz7dO0jQonscGE4Unur09HXUES
BMvjYZoFaEon42mnSml+IeuzPdTsEiILA4MIxJVdHEOGFjgVkb9XlLjC/3madXVS
8m1ggZugM913BP+xu9h8dwUZyrMU72re25mgVLYoqU9//4nnf+E8fgVVRi2/U+Ey
rkccILUvRc/V1WiLZU82KdRHQ9Bt2KD6FFsMpDCXhFFJ6MTaFlKOoISMZregIrR+
rF9n6MMRa60IJCjwoJBdQjLb2dl5Kz2Qr2iNzdVZg9nsqBdYYndCboJK9F7L+MCP
5s1Ll3scgH3DQSNlvBbSrAJiNU5o6N4s1ZMHsBh9ffN91t4VgOEIE2oCA6md03kx
j5ZQ9db0Vq26vRa/Ku/0YgQ6Sifz+Oni5zWtMNzhUs1qScM1qXaEcbyQHA0DaWE8
/E29goiTCfPFcq/RQHeWmiETxgDk731d7q9u//Mi8hT3r4xaCUJa7pmWEQC2PniV
4Y/ABr6Tb36jAi1LkhMhp0EE9Shjs8UtIVSvDghmSYMVrmZXag7Zhgknp1/2CG2T
yRM/F3W3NnBCV0fYDReCHwR2cWsgG88LCMqb7nmCvpLiKJ3r04uBShpOO0XZYWuT
bl17/G81+NuQfT3shkVkPD2JbSpMxwPrRJTb+ZWYGVBzO0LreVPMDV+86kZrJ6xT
KOqjan18TCr9AufyFAB0HbxKKito8JrmrYpjjbShzVCJFzjfb1QYI8SNv/qRJWuN
VKNnCHGpHUjhD3YEkwmVibQw0k+TGjtevOZi13bdu5vzsCVX5mzS0ALCdSXKrGiH
gm5lKKxNZFjMUEBpuwwLPFCoEZe88XdWvNXgmVtODXxQ3QsnnwuulODVNw5qX/d/
DBwYQZ49dx5+g6DxlfwiSNyanP3A3fgCjz9vk2C5SVKglG/nl5kF0I4CKdSskTSv
Ir7tHyAl/knnxCAe3CFao7DHCQUTws9VR0CJvePRR5PdFkOePooBOYPeeOyTrSdq
6jJEP/UlTBGl3BEcu8UevP2eItQ6cent26nnHf2CKXWQntVjEs+8HvLPliep/xDv
FbCXUH0ZMX1wLp2pOjWkxiYzobfnOvF96UC22sCkIZDIwfKwHpMWz6ve3OHnuS8A
XCKCfSIRBf+YiLTZ39h+g7QzTF/gct88l97fD4Y+911dP9px7qeIZDZQ423kR1pg
15ysY5KVZiZVB7w6SroULGo7kLRkuiHlnt52ax00nZpsgV1kuVp2LstGujKBrS2J
k3pHuezRL7Ys8Icm18qb+6erSsv+pst2abw2OFiJJDARm6M3kDH4msEszNAzr8T3
qcqACwer5OFfVmMrDboaxpOLsKSixaerzx5kp/c+QmhCw0ejpxxn7CZhuT7o8ei5
Prze4MZqkXB3/D6SA05YTwmY5lipwCAO251j79EE3h41644+b919TF9TAj+xFyuq
uPxrP/1UT/AJ0uzrSgdegAjvVDoWJYV23u8fFvUWbaqBcRUersAysmK5VlP0K6dJ
lSTtqYCS1+INnViZ32BKdygt3g4AWF027rxJQYGJHownXtUcrha1ctZ8ewrgzo5Z
sdSjJ68e2JSOScJ8RTjBa6NAtemix0EoyvoLX5ZWZsEIEE+XxEFp8XDU6a796rQN
tlABkJx2U5d9zrgsq0ancHmC9GaAPH9L8OpGaF0t4/xTRYtKs6LrFVA+bK5vTr25
0U8g5+rV9P7k/nkq3/qMdjdirVKGYWrOqPKGoYmfJ+tI/1B/NTJ8UaDsBg32YML0
VtfBM0EvEINv9TGomMN/frtDCx4vWwozEVyNYAjHKu9ycQGoc0CQGVjFLqF6coWn
wZ67BZ2Tll12eua3/FFybeRM0Sddli3/lTdgXA1Gh0VvCpBr7wi68anfmhTNGV81
JuRLsOI0RIH94ugwW49QPhxQouwfge5J1pfZC4IbGcHLd2NGN5fhX14zUzfAfbHJ
EPAupI5lrcC49NGpM8KwG+xlFcdzv6+UnJBk521TaXiyIgWmaC/L2ZWY9EWU4sgp
iFSCr4GsVpXYvZEIDCl636/9uaIhL/At6nNLXXKsN9dArRCai/91i80ObTMMFPle
UOnES2W57L7zWNEnbAn1GMetpLvdVD2XxYqzRXBBnLIft6k6m1C84OARIjUXAX7B
D4H64ixwKdTfpBVr0IkgdHIpR8V1Eicd2/NhN0XPRFfb4XdA6pkVC0J/gUYVo142
EV5SC0A1MWYx0v4H14gsSMNPDFycWRo1OfwBJ7ROkibvbR5p5vKbr4sC9IqIO2Ll
5XioWKgaba7HxeW/0XGpCCLb+5GHFpFagR5ao5csnH/iOdCdun7doo9Q+tfcgvVJ
tg7DM6PZG8+mG1YNdhmmNBhndsQVP8kdsSCvoNyYOMAzoxEiBjFVN3ESi/in99ax
Bx5FPitgt+XtBzM3i8Xj377o9mFA51h2IBuPbY3uQni5eZjHyO/AjJ0TbBZ4YiJd
Ech5kR2MMAgeI1gyD1AA9ubf7DKwfeUUw3JgTeCMwsRka3a5ANY1XmsNzKNVQjce
nprHyzw/rl4gMFeSvsIHmh49/cvUjrV/3KdGi3933cxO6F3nVJeJHwoO4a2XSKpl
sHF23Yu0HnDRNgL9GJ4p78JLOuF4PYcxCguCG2Z5ZqdHfwhp2Lzle+vIABMMEsc/
1zvEhbDFVYpeCiYrNA9PyeZzUj82+nCZf0G9CrCLV8uF2QbWSaW+K8PB9LlA56+O
x/XAm/w9YDHOEIMX5lm4tCEKX+RNtQj0P7KJ9d7nEBROmDX968x9DLBwrM+4YjnI
PTDxfpNfQG+txpFufKOfo3PYS6ZObA8InLwOljlMTx4falFPPzc41SelXAEfvyBp
8wG59FynHtRF++pS5XS4un2OgULPREeSkEQ7TKt8HQg9Tw7aEeYxN9x7XApSWOYh
vvwRvlwmaQ202F0ezThZOY6SVM0zlPzE2pvQOWNqeznglYFEahqefSx22aN3TSjz
yqbBFRQhdt1pLOYeTIw+v8vn12PS/lpfuo0AGancC0x+Ks7oIqb4WENSUJGY5Sb5
VeLK5mfoa4F9HOROh0oFj6H+CzcV7s8HTV+1YRDH4mhuxMiPAnlbZ/eLeSjune5N
i9TXRY6tNFfahemyKOQUQPUpWvEymn1/ZstJrYcAtjgC2P1De5Qiq4NZdM6e7wZ9
qR/lfdSPPb82HgnpAmcLhu4bkIhieJqohzsQ9uU98sOauimQMpvgQ9hMJraxhaoo
k+9+ZVys1LEGd82q3iMGB2YBBs2ZWJoWO8wBfVh39e4R1/rEWjLd5YtdbTn9vVBs
8h24wSHVpQ/lcoY/XT043wx380IeFEWdQOxtjCSi0580LiHw1IiEoEeDFfTx1x2x
R2vv/Vt9RWo1obARd65/Wif4igy/7G5Pq86hfd1+/+aiWlK6f2+gIdq8tpPyJ6w6
qhrb8hHPasWFSWvJMBHUq7zP0MfUOU0rwiI0QD37Q+l27FMBUZ7MfxPM2wlCsvT5
2OfeoEwqEql1Ogz0jYJhx8IfFDxdd4NaNWz4rneeWIlxMGI6e6ZXYM7C23p1cDkP
3MJrh1yWgGFKh0mGhINroGGJ3SQuirz7FvrpDOTmwHYzm8+YqDpiRk8RJwQ7cmtM
PRLgdxFsEOzwLRF60DYsqWPub8VMW+EHr04AhkRCSmcvqG8GkIimLb3rGwGqBDAP
GPwXi/gLRtFWJuwHOGFVNyFSupuv/z+moXqbx7yQFKINlSwexDyVM5AXbPi7rKmI
BMym+QbL1FeBxtZxLfSQjcOzFTE7GfTqjSwTeEfdP7/F0yfuHStGxBTHQejuZpRE
vk03uzSlz0bBgQtVIDqKXv4929S1rQU0qPmr3x+kr+E1GK8MdnfMzV4CG1IKiHBP
rArzo6ZVQMgh04sw1KvWg01qrVBNlPX2tEzQQLr523/ZijcRuYroeKB3wHffHI7j
c1HH8+jsEB+qxA6K89G4rnp8pxurh34cIqXz6Hu0In/u6Yk25yIrtcKsDODQmxb7
K8GqyrSdL6urQhe3SdiqC3lNEAtAk7ruzS6TTad95hGBRt740z5SGqYOKRB1C6iJ
DPmflgsnQecWjFoA+9+Wtw85FV2RFQAEiVF+swv2wSKchW0gBrIMFoOdbR++FOdU
22y8mrZyJvu09U2HTlxueDb8MIMploRQnG0bYXJC8vA8ICSKSHqsAKd9f2dgz+np
2NgOAaXYDgrv8i8vLvckMNrIHz9PAIhmFwEpVkqpwvQlo8MQ0OUz7yrjQeedSlxU
ePE5yo4I17ZKFu8FZK/3D0t4iR2CQIcINfu53U5aDtvxLPiAhirPf/q9iadBvkS+
ynl7PSL3RsLEbz08tdr1K++DJQRz4pnSLdfUMxYf6DFEFOI2YwQyVmPZslyEq/cP
5+0UOAk+7zIwl3gQZWtxdUfmBsCk2dtpzgbO2LTHY/kO1CYX3cqZs0yG/oAdx71Z
54nbJs4kBi8E6NqAA2Lxx33bXf6cOCAheyCLUrYlXfE3OryxDiALClfEQ1DOusjz
cD430l5DNrzQUL1Pg2/9+g4on6jRn5zW0WsANHhQ63qb3e4iNdJNTT2RybTGEpf1
f78QHOESrMDfjTu7CDGfCp7GSVaYVi5bAJztWsJmz+GJHY0IWr0ptFCunr00i80L
30JD8iRydfG30BD+Bm6Un1y0S0OwJzB2Sh70UyWvnyGJBlrDzIuSia/tfXBjvQWW
9gN9PRdIsNoqVbjev3h+dyyz9+3/GFWnbG2UO1cpV5YZUNHBQrqCjI5e3GFNHa8g
uLgARvEf/InQQt2ceiWE9Yvkfv74uHnWH6KRfvatFkaDF/2FKm1m9s/QBTB7EmRm
rIePkEpJ8BSDny4DRM/f03LGHNxpgf1bxkGZO0rVhJQT5eqzUOdGHgGf6E0PH4Ut
mOEn1m5ksOmTyBBwKouIvdolchjnvApdDAliDbsWVnED0ZID8YgOB7cvsiHM1fc6
/XHorvwnKC7UpOPmdpz4j3xD2D51BEqfdSmbgX46291yHm0f6D78L5OcgNw9BL5D
oIzN/BM1ri2LayT2HREb7PObKmFSUrsptSZlQpmJdME7kVfA7NNgzSeHRxlE0tXu
+XJX9RSdzPIxw19utnGH/ecC1RMa0jRj9KMc3zb27v/MjPFW9FMJzRO9/9HEP7HQ
jTe6h+zvA1+2O1q6mx3GFGFChXBgHvovVgzssWNljbZyguV+b1Ozaut1vtjf+Olt
rfjYYbxgJPJNqotJdKNRRsEnNuaiEQh5CKxn1WykZ9jkWxdrivQCMPSILSGi5gRS
u3vK/Vu1T/pd58LMQtaiTI4rmkaRtxSod0ysDNmvaJtoUIxpggziyXVPMbCWBtsY
5W7VpWdYvTU3SdASiigX4TLdnoF31cwdEHsKdU2gMPWx6U2/WnzVWA8h2ZGSkor9
eOEwq06Cn+PoZtHglh5q8YJofy5NGEdpuQ3FNHt178hrioW5bS/V80+0WkQqXNzu
fMdwYgb4DVfhDFvUil9W0B8Z+rgpcn6TnjdkieqJr/ot8WI+f/yt0lWNl1ffHZAX
QU2p1PluAIWtCZDTzJ1SqjKaTkl3GkkyUAfRrTPUXISrZeOkjz3F8pIy63m0pJjZ
njUJ8OiQIGtV36i05hCgJr6xAwYvP5S0yEhKZP+j+j50aZVvjjtU6hZOKDTfDwqY
KnH34nKT+9i3cVmX5lejzUVIwQ3gvV+B13aZuRXIlmDnjyQ+kvQkzbZ42StdQfWw
dhtwktwYeOYA4j86LVpSmok/dW113eWeS8bW9ACkPjH1v6RTCKvMYWGvhSLLNUsV
OOoLvM4GkF5B8mqF4+uzfMAij7sq57EWoEIpQrL5B0AF3oiEgc+ywdC0CfVVOaTN
5ELxW2nhu6OMnQouBh+lZCXxvZW17NrTSopinO0jBH879hKkDlI0mu0L2Dh0BSjq
yD4Il1Yobkg0JKb5T1TTPTvtPcJR1olpu0jveIRWZHHwwhM/aB7YCUZ4XTDlrmD0
ZNnveMq5VDazxDcZUD19shzA4gzHa1xaOD7cO1Jr1KoDL+u5ZrCtl6PkvspHb0Jt
DShfLXMRL33+yywtmFmUuAVK9bX4JoEMEk6sOqyEASDe7eDCIQxpNbOS8Lwj2o+H
NcIgjufA20X/dJtbNKUp87NLHNqUvoCJ0kxI5sd0+evHVzHRRr4Y9fvIqnHF/C/f
kax8CvMNUXRQR0PZdLdbzbkwBAFzOrHAMuJ+zVi5exk2uCAKpIqi3p3SCsAgTqcZ
NuKIv/yocu74mOWm9xmTtfRCCKmk6hsimV5+/Z+AfLaIAMno0pUvhi71iUVANXIZ
8RjC8DhUvxJ9BHp9drKrKwNiApWl4wb+0ndCbIshw6hJQGoZ3HfRJDvGJh0s/zMb
zVitdYy8bNjxGcP/hQGw/FnX7xx3Tc4PIt47kBhKtgfFan60b9cBfhYliqSBnVt8
HyYmAZj/NyLbZXRwBgpOlFSaxtaczsPj08ux/9VdQYACDpKOU6mqZVuaD4BOTpWT
L2nYKTB4xtniwDisKjC8hxxcVa12rXPjxhLO95ai+1DSm/Olb/h54Y/o+nJt/f5N
1qC/IKJYlw59u45PExMm+QmDixAny03TwAgWaOxLH5LbMTiWjgXeQtt8FDmzXTBs
KWVtLTv9r7i8VnOFeiPOR5uiXeEoNrXkWhk5gfAdsifCzrY9iNfwLRvVPUIFtIvz
Y47ndQzNtlc/AGp0uy5WXRpCwUYHtHvsTSs2mupBEZo2I6zZqkkqq9JYon+8iTdA
e39B2lUwbMZfu/IKVRQm/4JxLCPfrw73sJpNVhz4uAOGUG0/wb441qg+zC+d+h3p
lLKgBznz8wTslhYxJmGHot5KsRzKYl5DK66bcdrX71PdfkcToK+jOqQEOpms8aH5
WglsKktnFc14W299+tu7teGqSQCOUpOZYBF8argg5OByA5hxcaRwWE9i9qPwYwCg
fCescGjQblBVScDPL7pjySno+pvNfTxBv/+d0fCDzgcxsWXHINC4jCqCGQ0YK0Ge
odA62EtlUo5DZE/jdGVNSRurkSNFIretcjRi4tqk6LRs+VUr95tWixOhT/fIJXSW
9MhAkqCYstgwU84N7TKhr5YVyJsVWr0hctRFIkakNt+fWISb35wRV8laQLOiIEtG
0RzSi7ltW8GyybmF9TqRQawjMoOvCN4L6HedEmveg0qh9zMY89FDK/2cEQUSwDId
0/LjWT4LUYYLhMhL+yZrcrjrxfHGCa0Rv7aHUVhmmPfBkkDRxUUKMLAuWon32cs4
8FWThdT19vG87qpnP5RCOgDfmsApWW8CBSb7Gm6c0CJfe+DLvHyhl2PP6BUU8XfT
v/WOn99ufTNFY1Hy7xWZZ837lhgvNwJWrsCwIc7N3QS8rHt3u85Fud+clbONNCxE
OFYrWpqRTBS4sXSK5SqjUUAXMpbKoPXM7Yso9fP/CUaauO5UZjFltHe9K8MAnBm7
hL6qL5ch5JLX2Rw8p00DYsvyndzsC8tXt14sBnVxaN8qrdI750rsAVvv1IYq4pDZ
7XJkPqjvyoBHHF3TUttwQuELqC2yZIuPMhXnK8dMtkGrLx0fEElfcOI0v9T1eSgv
JmqLoRx3hJG6bkecHXvYn3vYMIvb9E0OUoZfRfTPomGEmo6s5V8vJb5IscABlT+m
5q/OzweRcjF9uW6mLGZBD66RR709FtVeU1X4XpaOJXxy44GXlTp+cB3GWPvMMWVW
7KXQAEHFPt4g+ZVvpAd7MFzICu6WmF00/H1u8rcdjugNlgNUOCYjXW4wyt+1eYde
Snn+R6nVWg29TIqa2UB8LdwSZfPOIqsDVgK31S8KzJa/t7sGCvqEMRuJ7NaPDIKZ
QQPEyR2fotYme2KYwwYYkalzV9nfP/jb3z2MD+483IgGMCHtxXYmi9a09F98Gn2h
AMl/b+vkE+tUC6XOQrRk4JW3z0QetttmYUwVtt81m3z3/ZwyJ46UeBvOqeHaWUyx
9n4JFelgcg1okhOsT/h/MS7hSjLZr4YRHVTiCRjK0uuHDK5aTHF3GeSMdKzb6RU0
Owp1908EIrNk23jXMdDBw9qzVrUwGWNt+dZN3g/Jxm0K6kUFKNxqCwa6aNAjbIiE
S2qcmMuX4awSSsGLv38fb2XB5KhAJXvqmyR8rVTpxslDf3iTO6eo+spjJ/r3sBNg
26Cr+eKSWCDBM11rjbqV1Y3eKsVYWTcaCGZUOZijcXKffZqIFGjqWKQeGRvXMaXS
cAMUexJLunoOpp2CoVtYPTUZsaH8JYVrDlx3NFDs4yi1WD126g7KZ+vx5ct1Vuh0
nCvRHHC5Rhrf/wqZfsN/0LRrB80qqUjuOmJNTsmeTNYvjWuRNW7wi7nVHfxlPBso
V1tV6tG+RioRI5QkGhKDTb1zVuipRCIXdMyvqMfthglobYC3Xnz1LIHqiIYHHpTP
CVXmhZuBsZ75BHdps282HCKgQcRifNxaf/TEuJipV8iQ4pV4YxytnmWM9+AhsQZG
FqJ9WCkfExMKxDQWOaK0gG11Hnwa5OowqydXiN04kW8HVa2dbLnZJCcQkT3nsQWu
+VIDMWt2ToMN265322scDJprtDm0mbCDLQ2nqMKGAekaI6ZeRRdNYw1+iewVJFB0
xtHTt3LvjLxlc0IOa4WQ6ZsbRis6r8+b8ytNmBLAcuYLOgw+/KQPqxM4WSwNT4ru
/VpL6+yvFPFSuZ5x5CIB6q4nn0NE6+9ft2PpDOLsemvyIXJxrm2B8dTkGjmEWOmI
dqcwvomqigsT1h24nWBNavmccdz0+S9qULBbvx99tSnu2Vef0wAh1BfJo/mMeXrK
fXU/BjBKW2YIFWIcoOTpeEqesw/NyvFHGi86yEk1tQobXsvgl2aZyQtYlIM6g/cy
ErUm+Bw7LoIY21tw3yK2JgfoAKo00/kBv9semC67ylS9jOZWGW3/DZsjpaZF4N+2
pxHX5iGV+wJUePyCICDjVPI1TGAtYZGLG05EQHYEveqjjadUrXJPNoeq9dnl0wtg
MuupLWdWZYEwBU+zzhL/PzVhCrTM9xu2e9KgMR4wsmqk9n3s78bmMFFpl1N8ZMbK
PIyqZSBnBr+6vw/XaJwgVKITQB2VpdZDcr1JQWSOj7Bbxi54hFpK0aCIW7ViE9r6
Yon7uQhtpoc2yfXYcsHPBqqZn35jb4YcvaP5KKqf5TO76xH+XwMlN4VJATItX+fB
BYgF/vMqVvDo8fmjcRUaUFbKRcSpCFy5HYPnO2EwuYeaSL9RUG9AttgTAL7o8VQh
oDhg39D0smBOmioOJ6QWedGit8qccWzLA60C577x48ImgwITI9Gd2IKKa4LCAwxv
eEYtFzM2aiQhXJA1uNkQTw11pdvpE+/GVReoHltHP8JUI0b1dWKRnSv1X+bV2pWb
9atLHlPFLkxZlgu4y5nrObAgnFe1x+GbSefTbI/ZTDZjaxdBjO0QoU+KXqr6a/D2
9bgU0iBXURRLjGRggJH23ifc5AQ79XH0RrXEEHsHWgAx0N23cvMd/tAdRBl7FxQv
OPClaMVdBqoR4L8WpVBA1kN86nNpZFWHqTkUPe5TWjilUHq3/TwHsp0id+7PRu4+
ydO/Pa+o0qa/ITsJ2iRUJYcBJVb6hacug332HtYIcnRgBX7UmC2K2+ck7+urvNyF
cfO0Tg4DtMsgg2subG5+vzCgQTz31KeNla9SaPSMGkkhbnV1JnJu/OhonmPx0vkh
h2VoDgG0DyMLrPcN2WHhVnpNvkKg2S4WG/Ve5VZkJVA+lVtLZi2FDi5vzu1MkFBk
IiG03Tgd3iMjHseC8REWKxD4JTNhJen/pl3PzNqCPUGuOOaAm27BrYytMmzKtOBA
HlA65NKSv+v/c8GJ8yoJ99nPv0JGUJ9TSeNZqcN0+bh+3KEy77lyHiuc+UwkCSQx
qOYSmNHlEjg2bbVKIsfCwbw8GhNpz1/AJLWgwJ8ERC1g5yTOWq2sJANVtELx/QKI
5KOaVQpIEfMHSaXeDSudLkqHkmVoh0Io8RmEr1LZ246KckE3rVDGvgsTPnqbLrJW
Un3FCqEAFfXtT/BNCvKwu8z+etgPnmQt8xIP266hnbd0QqnPTsqdfvRx+u/xWuKw
f8N8+9d7wGkhPIo5wmRi7k0nXTLXSAEgTn3XVx9tVHigQP7daSLReSjQdfI39Nk0
jXmcLdCaS5BCJflJKbM5d1VP9sfEpJKtzFwaEpaaSrtC7Ym3rO8W52WqCKQypHO0
Q1jNqosu0EjdmFzvJCqEx7EfNYEgEL97ob1N+hyld3k41DYAcn97+27giAflQhZN
Z9aAZ3P1KpesWpqunfOuDhVwwOtx9hP32GFtGwKmSD5WPv5y78gTJm7ukrgeUUAd
BpauZ39wxJQ6dQZpAabUqHANIjU7jZcgOczIn+tzgZj/t4ChTvg268+t2vSIhxo/
FTURNlabFW6DcsyFo+YPLCxRkuLT3eVFDtRl1n951csj44TzqpoD4CwcjzwcsXuC
1nynnGkluOUV9ipyMJ3Dz3D9C6m02uTyWvxuqWLQMMUXR+iBRMV57rB1j9VFwN3x
8hAnuu/ksOeZtz9bCGerDnB1TvIMkdmdHpyDEf5+ZjNjKK3999avH4WNm9Hev3AD
1LocPrlkEngSYBFcPxd4/qcS3TQV7blhEagmwjmfruJUL520k6+VDS1y3XdQWpkg
yrmte+iOZmmC3HXe1kGIhJsqJ3NM35yrIGo7YaiViu6DxqzB1V87c0e7zmNYUag9
tq3KvycSnbAw4RELw3Npr+D3VWhvi58HApn3t2PeBBA98nStKeQmEKlqDr3QohLe
9TT7wwbchdviXg7d4jS5O4P15T84c8IpU/kvW+PblFtdgDKdKMBSY5/T65exV7mQ
AEHUeA7S48P45dcORR6Uvcq16fkOglrpE3htB6LuOBEVEaSBVqr0UKl/i7mvxgiK
u1bdg3tb1DowrhSWcCV5hYgvWppsORxc//xizZxazKEj15x5toB20f9hBjf99dNh
fDOHxWIijNhMCdFcx4bNleHprvIgRN4Id0DztzYX3pBJOAmeyhVG7nHX7/3/fIHQ
eYWh0RznxU2aFao2DvrUJoiOZWvu/WjSpVu3jWRTbqmVzbnWxTaotUSoGjmIGGK1
RvlYkgPwDq0MqipKKsZ/q7bwQ0c7dWCslRfEDgubk9fs7Gu3IQV6/13zLqqj8+Xu
bpoKrV2cGegdD/SN6uzE1YDSh5fLm1nY8jPyzTx5IQ/MoMK08/4FqFLd+QxKAb+O
xiXwyWyw1/M+K9ELJPWBlKkoFPninhYZBLw66pIVsgIiWE3OFAtWPHZV0d1Jdv81
SY8QO4GAH0Bf/T0ltVnU5Q8ORcckq8My8BMVrwIXBIFRYJrpsduhFnoMcQm6TS8m
ulMOgIIHXPipMdilN3FyT4qHvBI8Mb357MQOFUYQlDVp1B6cSJKk3v/XcNq7SxCH
4RSEWjEt+ziaxmiXgXVAnICOGMGdCmDIiON8x5vhwsaZ77CdJn9xFLKTwPVu/mWs
V+kABYoaUGJMFUEjY2/NuB9y3hLeqtYQ55Svi7IuxWlsrc6tZ6auMryOuCfG56zE
aioBYXEJe14T9jbTJbsH9wgRI9mXYdHhBVGlEgUEqTvcmQ5CAo6555GkQf+KgEet
HVHTsrmx7PT701/nsUZPNJDAKc2J8ZfifDPmetnhHEOBHXLER0OSazFWx7TnbQG/
/3uep1ah0HRzHrJE/ViCkQDHMpAy/LrG8sPxNZlQ+1uUZTSAxqIrd7fB2fX88vf6
QJ+s6R3Vqnl37wtxKA2Jq7ccVOQsen5/ysafORrRQDGfSCjktUkUVjwat+xaqhrP
5MbgOGAb9iYi2FS8J4oRw+SAyhLcTAMYdFEA+o4lxxFbsRIGyjbt+O5qIHXPstzB
QYDGN8l+hPbdS4Wk1A6umnXG1p0g5YwWmxmD4SxPdIsaJgvqfkXgr9hLg7GQkEcn
iN3r1WTRLA7HKFVRN81ZOoyjxsptt0Le4DCmu2uOvZrYpk76HHGx/Crp8xWVxtk0
YSTGYmWtuqi2SsaJeZK4ZcWyBd5NRuT7lVtDxoj46WNpMLGyn2+ksr/wUEkNnLkm
G+FBUntPatmcZogT1AfME+Pt+SnvTWS8AYJgeqgR8QlpI3FpgSN5DGloTXu2secU
XZpOxv+aof7rimBQdbKom2nUSIMwHCY1mLlbxP7nS5X634zC6xDwM8symjOBe1l9
3m+WqSoT1RK9aOYnppa4i7C3Hm+9+SipJpgFApddMiMl0Jyj6R1si3IX/zcA42cd
UzjuWwY2/sBMKhI1WpH77vv7Q/TKGB3VJZtdLL/1OzctwyYG96Ewu5XOghTUJZhY
4sTf/WS7/8Z7R8abzWFqAqUCuHLGkSE2mNzbQ15waIyPyPMsKiIs9tshYVQih5/6
qvENseHv+m5nnmUGovy08IAt2cbOMf2g+SvZEa4GcY/PdHhD6uxN2CgB9QikZ0tv
K9MPrY16II7Sa9J/3lW2+thGJnTgm5kYnqqi0Qk1x4fAKd4Nzdz3rB4DbAL+v69b
js5SXnR6SnrslvgU5NUU3yhrVw62dw8DQT7fC6mFYzVdshP4PqBlGtKQ5si/ETjM
ZsobI/3h3vz1DDwFOovsUrMXyOyH3TZYAGFfsODqnSnnT3fwsV8W04mzHAQLvQl2
NRODo4L5vNu24SuZP+NfyqUvImKDEFut9R/vaSbG4ID8hlGact7WPjWpWKWY8Uyx
X6lfzhNKduIp4deJahCxU+fHisTPxOFByIkJ8rA0VbY3nmxfFDR5PLcPV2e2QvqJ
0hGFr9IjKYn9Ysl9orTtLVyl7lp26jLQuVgeskr24lq8yeKqfASwZ2Aee+w/MObF
XxvZoaXTt6G+ySXizyK3VDlYBHQSEPz/UQZLzFVlbFerMrsuoIzR8V3P75GOJJnG
emGH3ghDhRKXq50Lc1G/vVVXNqEw9AqOtR3W0j80xFzYaNAIb6RFDxbRJfkUTC3i
IK8/qV9yrZ6CX7gA8UutADfiXeNDE2qUri4iIAbEHFJ5nm8zVGwl4XkgX0P0nhAn
cpT2PZGAYNjYqQlO536FTh6hqtoqZLZpUv33rlWY35Fobv0Tk4d5NAe4hFkMFoMk
ZxGhquUYrKqb8THPbtPcaxXMucK09RXDeJUwCzZuLYT1r9RA7u6IOECWAwaD3gJv
rRbrTAebgxxmuH6/LHJ91HmzMOe0RWMfLW8fy2CDK6g7xKk+nexSI5vaTpHFMnLt
Ms58oAkJNzYZWVPnAoc1JFYEXSJpnElXS5f9oA7vfO9v/wf+SSTaTEZ3f6rbRG42
UDM/vFweUfOulkOl/6eWMf4STRHsryT6VsEczrJjTqdr6/go0ZWYuBVz4rjTpE9y
xJqL2l10ZWYXu2+hJgDS1qu2/A1iJ3VXzz5qrnwf2OPsNP3mPFaxC8dWCpBHZLL5
iqfDEb4gROodH5MjiuZUgqG+FuqfBGuD0utfo3mMz1wzyE5L549oAu3CNK7WPvLH
FA/Kcn9B35g0hrHBQwkB2nn/pYQZC/0Hyv+UC46F3AkuQ1nWRGit6glrWsq9X1Fi
31VhMskQsDls+8xnQcINo7bHaLXmyunxBfjWUT+dGjpG55TZvhdb5TQCpM7F9IDK
bQhDGxNkfLNwNi/cmLYXRQomKmYITHGqUeuj9e0zkcKEng76JEmZvw6F8jadYamh
Rwmh4TFR6nn/FSOMWiOK0nbskBSrgONAu79caxjwecNky6JscdMI5eNdMKVW8rD6
HZq/7FTsCuplJqBl3Wc65TP1q12aBvIc07mhX096oh0V2v8El/g9zBASq5HhDEyA
0yr46dZRSIP9LvR2+fgbBe5TfUI2nXmWrrEqfIR50XvflUQadlO+JXJuxqimS/AA
tWnCxUHEPVjxaLtQv3m40aAjY8IRp71MUmriAvm42hE+xnymBVtSANuNHoU7c5lT
Y975YLb0ZY68mDm+fw1TL4MUoNm+QNZMhho6j6SLTdx1+F2/Duo2DhKAobBUcAaR
DkgMT1UJ8H4KK6ipY7JJx923v5ecPEPPZD/7zmqzZuB5fNnGjNLpIB/0AfOiRNwu
hJd0vdBUo4VqTT0ER4n44i+BhJApX/kGzGY/XfZk4NeBxzPLmvpqAz6j2ua56hAc
UzdetMhJu3JsSx79gM4hJSq061q6f5T4ZDodZYikx2G5ilRggtcfUFFVZpu6XE7G
YcuNaWjmxv1eYCMP75Xqbp/ghqTh6CvMX5rgmAmZEm4epJChFZ4O5x29ZCr18lrn
2mNwKifp5DxPmrpTAtdxyYjfyEzsTC9y6Cyz694KF8F947WPjczNyi93ykCuAq9v
VV8truMRhGdKRI+7JBJyHkMLW1myJKu/9SUFFhHKVyZGW1VbO55CkloXcYhs0FAm
4npDBYZlfO0wikaRKtyh/leH2gyn+qVG+DRfmbPxnTrvp80hiiusWIZEPPswpCWz
LSnRqnw247GKd4CowtjCgzrue/noApyq3MGW63gDtM+epEcfLZII2tansF8szSBV
Q0zivP2IkfcGt7BKcifBvJaS0LIfnhR/JwC9bO6BDdsZ/c/JhsvCQVXGLGnw37XX
qHALB+lQxdl386ZHHyAjJcz4l3cun18Ilrbv2QlQ9n9+ZQ5UsN8VNupcT4FClG3O
m80vJR+NnMtaSPvXY/zdmbCfRPmYQQAy3j7XfxM9xZuVOSYyB8RmI2Z7OLpvWp7T
311EfFGtxC7H/2xxuOqtRXLPM/06pNhtW0UKC2UurSVZvYh8vvMLeAH9UzlGjUvl
l9pYixspRMm5yAYJopMpXkJMvJV6fd4IzuF9v3Dqhtd/HSlHWTH5JmqyHdAqP1gr
y7li3WEUvnJXwqNEcAvNejwoM1sByeYR+9HQNL6//zb90/y96L3gykd92k5AWNnS
NY26H6AMGHrED+rgGE+oLSdaWYMJ18sMPlGXwbywsmnLPCSI2cKoIeMi4ibvT9uR
chuaJabHk5hLGE4W4WdzwVvuvGxdXjelycZ12jijo+Z47c5oMKGDlr4f+GTkdmvA
wFYFwAlPvll8hSEyhqOE/lbnsnT3EBd+FWkAtgnRRoviX57pqAczJlszkuX1Gip3
BxEsP1srQkjdgBHr7wSV3nAhdNyRHJGvQMaGxkizWAwpoukRSEornO/wxbvqdTZQ
RJvrevqYAE76PQ5w3gtejYrEIAX8WGxJZZyAwRj+bvy/ZP25luwBOnn8LeqdPLn1
dRQ8FKG57Nft6wuQrd7CjoxRoEKUk5WbLbHLqYtIMa6Wqd/MO8Leu52MI+posy0F
SIXI68GtYINtr94A8Em5vqTO8rjal7UrQ/YNEG6oEOKQTNPF0pWl6mkukKRxXy8/
q+qSCRIMZYmRHD3tckRGuFPfMOpJJmFJlOo6xMkRKhzGCcVN59/kef30E5MyA2Hc
yfla20pfa/Nxpfc++9ZpXfgcfp72NGNTi2woFDfvfGsEyPh/IFydyz3XM7Th10Wl
wQ4K6xMKUwc7jRYUg6K3PeZjrU0W+lslZU+7zApJOM+S6pfk686K+L8I8chBD/vX
D0eCD49V/C7mKFLuqL+EgmrxloPog+jdhcPbk4nIyik5CMxO2wWylNfxXNufht2o
PyYfsJzCIFmauYFuT1LWuUufHOad7FZdux6Bjdw0PkqwMnrSvUWbacRO5TDEGrGT
bP3Ykjhv+EtRjeRajt4aPtCv6S1QkmNqp1fC/fGemX9bkbScq+g8/AGTTha57U87
rRbq3W4/NHoL8a/M54h/yimOcRsuz3H64tG/htz5s+DCrCnEn6X2AXUsh35EYmOH
waD/s6X3MEnmpcbqVRljplNepV8GXXtRuzdzA98vedQz5JYGar1OZFFlIehJWuC4
mkCV4VBa2vx1RdAMunKPhKo/c4M/wHXDeWRiRapvR/MxZFHES+gFNN9upH9qoBpK
qZpTIqi7UyKOUW5uHFs69E9tzHKswhn3AJr4P1CQnSi9yauS7mQ3bkh3Umz85NfH
FF8j5lBOjQIZurzlfU15sJS0lQK+IUMCrM6t9NGigsyzUld5VsAjOMd6bLT/TPTM
Hu/oNEKh2KiyO5lkC7Qx+3P4vEwN1PRsPX688CpAbhCHy2BVR//afnIUEzoTopdK
zwu09GgIOwxXFJQd+a8oGZngOF6Xw1C+9mEN94P1JrbALi+uRm5+vbAodb6RkGNW
2Z9cZRMZWJhtLGSnjBtdqvO+TwLJ7lZX1a+DnsI2dD9Ah9MptDh5YmqvhQJn1TX9
1MT7RC7tPQLw74QyZZIZ+y1mbaG6SxVFlk/noPBvCKeZoUd5OAz1xxCIoEaUlEr1
WOsXn5rY20kqJ76723EYvj/wD7/R0vC4Fw13+IY9VqHe5ADmBIZNFGbW0n+t3Bil
JpJ9YF7YPAIqUFVROLLE9zO1bQUWAo8EJRkp0/rlUymy9kFHUdKBk4zh3qtXlVTv
JpX4qV6MIUpSYCTgivn8vXNn/ditHjcGDCZYW3MrdUF6JumRp9cpxQrVPuDmXKIJ
OzETLCXvUIIrHcQ98Mvngm4xVK2GSeCI679p4V9nxjtd3nQYXVIv/onbcWf9eLVH
cIcJWS8kq6e4F6ovdRvQcKin6MpGNaYYIcdhVNLhRkVQ7vMf/yEOoTks2iFkXkOF
g+DIBjZGQNMekbqmcsdE7vPgltgGpfXGuk9KVrELYunsnvsQofECO6pPfOTmZKg7
0QZoJQRfbLs8m94qSo3ukvUrgxDyqFz2BSik9Xs8Kq2nzmTpIRPBhjVue2korY7g
JCLb1CBu1qgDsopcoMAdwUjk9FZGrDAU/0/pEYJYflWU4WxZU8/OTtVlXZMeMOg2
NLyVTRnVEBcnJmfjbE7+Of/Woj7k3sq88Emq5vDOaH02axnTanNqyXWSjCcW5zhN
OQeUV/GP4NIQ3/v3YHeCCNTeLUTsaa+J5s/KtrbhdpROYNuAUjkZZz55ZDd9B1Ul
9TEKkuqAf9o4Tg6FyhPnP1FqMgOjjqdg2qvqFpPWc9PRqPXRUQfFnxZXGLKx1eF8
WpxsdQ3OzIQ3zsiHDwiZM35MHKLBB3N6eHMl77hDdDoLG/CKxNSqJl9p6XFjJ4f2
7i6WzCOEjE8TFidmNdYDYi3AJSHBeIYrQjhQMs3hULkFUgC/Tx2d8i4MEcn/4D5k
7TRlfXT5Y7lAiE8bGMSlmcUYKyvAboXYkmlF8hStSlhJLDRJjw8Jc7Mv8+ro/UF0
LvnsQA+U7/4JlpeL1kVCLzOTYcZa4F1Z5ssSYXlT0svTIAMno5z+jmkirNcOH7/c
/o+65jqi0PhEl+a5ay75+iyH3poELD35MRDEakFMaa33WZIqvIAL0FiglpG2L5mN
Jqu++W2omL0oIY+SBGUL4HlYfYCx3qrLjG0kZDxDs2umAGlAHyz9b+spGpMjJzaW
6NmOXgbwV7vJt/nD5B8Sraviyr4momEjd+UvoqxvRjWxzwnDbMXQvXCVHKTKmFir
dD5AU576Y/+VENM9Ueatuk1JHCbrZRgdmp9SdANrznr2BckujX7aTNfQvSvxEPrQ
rBh5grsW5LD1WPHPgyzzsuLJ2L6iTxzJDeN5aOApEbp5HmS5REFMLiw7p1sqrcsP
3SQslWRF6KU1l07ykV+VHQVhNnZjs8y10DJSYGIeFh8RGySUxhsn6/+3EUnwBoko
7YdeIQ+ZBpVV0Jj9wtp1fE5l7RT6E5UW1hSe1jSGxxDgbbgTS+lHNEgPLqeWB3/A
SZr5Y2vqlDZMrXTTGgGnX6NzEiuvP8FbfVVkBxPuc8au+1hUo+PpCltwL24JIGWg
2h9diM4FWajR+Xmdfa3klVwl78uuiowq2LpjSpjj4uqg7k7Kx/Z2JyuSzpBcUp65
Rmj9vg6fzZQaJH+d5A5fJEY70/5KebSMBDeeyY+GcrRdNXfEV7eEmji5hj/nzD5n
gE1bCUu6xj2hzh6wLAWmE+dkGSHAEozbYzCXxo+OttiDMPsrjcL0YNDu1ITxb6T6
4cO+/aIVR1ZnDexT10ywt69dPPF+k5PjpIw0ER2PDMfhoLjflAKJrgJNztrHF0XM
zNWXcHBIvzrEVJoAHuI7EmDr+Dzng7XXSRxeBwsjLHrFQ5LO7CR5MzONKMyldzrk
87lFpx+9tyuxas01lVnNji7PEuI6N42KPwSCZ/IFtXdoRK4j160rcUdzxDZdWZsI
xHOrqiQNGyh4OVFcPSu6bFUvNvVcKZV4L7eQDF6RjQTWrANEzmtUDS/qsVp/jein
lTDT2Je0kPLI1Ysz5bYGGN4HSf6A+d0ENlBwj3yZl8aRLT0SVDNiWVPdmJl9rjiX
8blqAIwbuWjYM6rkmg25zntLMmzJiLjDSVwX/RTIU8zTtf/OHJTlacrDeJYnu+yu
QOzOUq313VP1qVrwgnqXHollJYyZ6oQ5khm2ty3JtdKBYmAzfhvvynUOgyWeZPjj
4kuphTRbKiMp+KWya8mhQLnO83BHOcL0CRJ0ErEKd6XuKP72+zV7GycTT7IvTy9s
8bCC3DOmp+9vAMwOnI5WulRgphD58I9XIdT4PzWvgGcxk3fU3P8WD899Jihl1idR
+c/bQkieWGoj5+7ehDGWOtwHwzPiE/n+jb1IeegaOSnJa3y9AutN0nR8S2PCFflh
R8SgrB8a6H8cI5mMa/TGZIsvk7Ak35d5L45Q4p3zuZrRungdPF8ybHYWqGhZw3Fa
YiyhcgjrvyubpaqHgmPIsE46VavQSTL48mptTu4gaf8Vk1s5V8K/rCxL2OQmRCJ7
zXFAT+LLPYwvn8o6rdNGD3wT1Az7+h0PLjREWlWe3BBykrwxL2sGkTHzQ+wDhzbq
1Cqzw37FAOJBizOKImtyqUQ+/W4BfkMQXd6PKFZnOsZuEtwusH5klPBiaxxBpZBR
FXAVQRMFRR0DKzvQn2zQHI9ncgB8AJnf6Bh0VtP0s0ZCXJmwmbx0oixi9wfFwKBw
OcQBmslQcbmSRvG295uC9Q2zQfw2Z1nAu9aXOpLDYf6zJMrBBr35twCHuRzEbQ4u
YfFpmIcovlMntCa+KgkbqapuaGLpUoK6cT6F66bj16DwYpLtYtHKcgd3qnVJPWbh
jSX0qRZl4n4twHcN8jB3KbunxNI02D5mXzQNUY1JcUrfKNMf2cFB09vbRLQb286B
mzTQ8QVALQbh85zw+buZ2kI6c7aMhjfhSenpSpzLMXI5A2F2rXceFrfSlIkPSqQ/
UtFrwvS65Cy68aJ0aTVNnNX/YGKbMyCyhvpjKuLkC2UrpVCNPQcM9WoBgaTA9OOt
qIHfjmkEeohyLPWhHEh/qdKjIDGreKEeCIribOCuw9UtUb5JPWMzP6zqJ6bXPep2
u4AEKX0tCY//ob8Oj1272N2uz/F5UDsmS1hVCZ09Qdgue8NnQVh4i1kOIU+APVnY
TegXS/zlITBanRmWieoyYoIndXMhMDqWHcVD+MbCp/ubpX/A85/nU76NegZX58/8
oK+kJx7kBT5lHJt5cxQ9pMe1BTXZxCwp5g44EpjUCVqJmyDFAo3bencCWFExA6+B
K0SkYznqxXrBnGRg5dlqGICbGAgN8VeM6uGiHgfCLzR3iYgfVvt6bki3ZoKg265r
luwNAohwCYwHfU95DVmBaZ3BmvN6F23CFGPmH6SouoUs7fpcizZ0p/A531fi3drs
/dsOF7wcX8LwwpLK3xSbDBkkLdA/Wp3yzmuxz3L8wa50HbUvVufrdk+2I1nhUPos
/XjIVPLUo+chI16/NTIsr4b8i6y+LPuB7MrsBtx1vsN5XG1MiADFPuxxLRsonnjL
Wpw/Q/mj3e67sEWAt5LkMObLAvoQ7uiZzBIvCmD4PMi3QD6uOIEQW/cY5koaB/uf
HmcLE9lznHeQA9RU1+nBs14DT7xkLg87iWsym9rO/34m37F5nQ8LDSwuN+Tu6Nb2
O/w8Uhb2L28uvSli32ZwDhLFnNuO5b7KX0c8qNPoxC5rOYHP0KY8wID7YiBNOnmW
oJbMGaRp//uEGPflYtaVnsDOhsflShKMhfQx3cZvVd03r60sqZcxra7HuOsbc1Vg
UmjW+fZ/CikScGcc2fZKGn3axhMPZzxnWTnwDBCB48pO28/8/IkYJDHhPv7sg1kg
nuvC2KbqBEI4eSJA5IqCxBR4RLw6UdUwTmSHmUMuX4qUyELeUYPg2bTfjhp317Qb
H6J6tYUxq8DFEYGzoOx5eHQviZfKCezhIDMugWp7oOxe404jnSCps22HamXPwLtm
JQLBUOAeOU9C1FbDxiMAnDBwI20R883wpHQxZS3jL3flqlCgdtZ5ShjGVLHVjSlt
7qZB/BpOBKGTU8wMaYO/PCrDa87GPnsma+mQr4txqizy488r1+pcf+TCjcOkKcsQ
6GmGGTRizt/06sawzSBnvSedn4sglQpnBdj+hTd5I+YKToiMm3JojwuN3VeduNr3
p3DIyZHH8IKPZrPUSF+3y49EzdQouBNvq4CxZeLyhpRtdSlyK4mFhXJb8xlxIplv
y8GlFLTatwQapMRSqaJr+nroHAU9hmBR6EB+4z+HR8hLn600w1+/J9pRQd6XixZp
vFtEmmn48oafqkORij6O3gAtG+PDOJReB9w5gLZbJoIPfRCJAWDUqYAcCv6fz2xw
7LBGWPuJvS3BgOmrt7c5EVDU0Vngaz+eZ5aOB1Z1s6VeV4mcPciv2DQEpvkvTxWe
A70oARqbjswe8NR1KKcC/t0x5/LhXMOPe7XhhQvlzlUdIQXv6m3ajtwby4v0G06d
H65n3wshlxvloKvWN2yB2upq5m5YV/6w6Q0IZwRJdiwrljHfQ8VyTuTWFKptieyw
v6TB9rv14SfCsxi/EAWsB1f1J1pls/0HwVf3PTPysbnHcuqvFDU6TOM7IrJYWb84
cPlhkt5sMIc4zcFIUbJ42K1VBWre4T7PwIHDy2M9RqDzyuiey5/ExzsEL1B5RJnq
0nB4XnTFCviK9tXZ2PsCJC+dZ4AgEO096LQklhd4Lwukgh8osKN4RZ1E5eNxzSLQ
zWSLtO35rj0Ve0+6dAV2wtDmwKywmeWp5muS6aWL16CkcY0SEQcXHj4YK19kxm81
7gTp5mEXlLJEuuWLyj/yqo6EKio2A5WsxBWJC/Y6nGFQzrxl/qLz5HqIZrtWIlaW
G5oIfXdKCBpAoP9AO85FBKM/Q2w3c0hvDtL2TvpvzakUT2yJFGrC2hnPfGiQWZoj
uJq3BMia4USSwlGomG5lNLzHHFj3pzhsUhFTG/+YE1xxYBQ9qCV0zZ6nOZ7yopHx
ZRUqC7MmnEFSFbvmvHlp8DXdR2I1rcdQa5DF2kLYmiq+ftAq0tmWDy8ylUvnv55E
SAajgl2EKXejMIfDjozSq/2w92zoco9+kjY4+GmgqEKfoYiEv+eyJhr+pZXH24Oh
gOVPqbgb+ebOy8082KbN/9eL2stknRr0IsLaccjNRO7W2jznneXymdoxQ+WovXZ8
sVKReFeA2A5hvazXjZ8N++HfdUpZ0D2yx/Gy5N4ZkUYYxRN6Jn3FIPRnCXakBEkG
gMdxh76+aYR2C4qu7L3zQpYdCAWCAjZ/FSKmRCxlroc3JnOrh1vhbwv17YRP1t65
6DZi77CCc0Dazxu5QaBRmZuu5/pMLCAVUcMobaP74Nk3H+9VOd/UKxEbNPQqyvPY
cK8eaTNbXy7sDQyXSxAu1GYzdwy2ZBvK7QAncW9AJPiNQ8UZOnoBqhMxlXcrnJW9
bzEkBDjAovt0zmEzTKhEaPhdvheqvrjehoz2tWffvjGi7PuSUzuSUr1WqjpBNXK9
xxtw189ken016OuTK08zZgz+f6caT91ey+DG47p/45rLsFbkpCSSEFJ4i5tsFSDG
CJqdfrwxfxgPYtDLjLBnUTauIWYvhItwBsJqKb9IVUHtaytWolCTj3AOnDU4zVm9
DVhBXMZsfmwOZp9rsWf+2PUeX4DpzSur4Rv7iJgAIiKhKBWbdYe3401UmcsMMehx
bflvkNQm5zLFaBSzZoDo3HpdAAAoDjMX7z9d/BFCJeTjmz1V2GJmU07nEX5Dwex2
zUxSXJGG37U/ddQPigIwQJReAcqv7tdYNKSgYK5/c+RQ7bXW7IJAW3PPb7K6Akdh
Uw5C6yf/Fo/ozYx8czXA/x8/ae2qMymiWCNJuZqzOeO5BpXLj7Eb3XW5Nx46Wwzx
xtRgWxfxiYJE6rPZpj6rAmXvNbEd7TzafTAEAqar2q91C1LeU1BtZf8JVdyn8psj
SAfa2hIu2WVsLzr7CHTwgt0DO7qLXAUJWPyk3hJ30KfQTdeYSTqcZHPDo+Rt4WEr
pvBH3dFx2LwRl+B24tiEUpXYSomsmZq/7VHAE+r8OQ10ON42wz8wKUz6e5YOEdnJ
fUEak+rdc6AcslVLUcIeFJkMBOUsm5q3EZ2p/Dsm/2EikA8ZfQBBBLY9MjNLdpBf
UW2vYSkXHYMK9HswixFuLoYXYpSRcapCgG53aJGUiZEGQ6GtGzGPv4s2TjHrQ8XT
KUdJAeNz4ldTXLTOl+aIWJ+OeLJ08JuFaCLnbjs1lPN2O7+aprbwCinLv0sV3YPP
8H2UiSUFssBWweWC8Y8Rp9YBNOs0F73n0sUYbf2vK5V0+1zFqrwroJqHBrIt3TU1
gZjsVpEH4MggNRbqnSSgqEcuUm1ErklaRj8zo63VvvlKU1FhILPpWa54dh+P+rI7
w7g4Xbdg7pceyEZpZVr49WST5B8ljexIZrNdkdj6hILEZ2jNie+fElr2mAmRrPsM
qPtonTJ8FnnMEK8/1xKwlagdMh8crHyuCOY4BTMMcKDLewtK8M3GRh+JZMKgpw2M
cLG52bFYFytpcocw7GqhUm3G+/cam8baWBpJeBTJAojXCKiEm0fEMze7eOdlcrqb
bGFR26HqVBnwFzej3md///zCmlE8gu7djyCm2ldJAyexRC5kmOqTyCQF5HDIv02z
8dGvmqbrRXm8cBx6wzpmujr4ebeCp9z2jep8dCtMsqFM/Ho9A7oyHW8HN16K93P5
zxrCPuha4qDHGIcQuq2lpx6vMnvje/bfyFSdCfLgZ9eoIqMlDq29RI1QnFK/40F3
4nfQwWJPwyk/VwGQMKMXC3ul0yhjeLoyZY65+itcO7+CtN7qfEGrXdZ/q6Ekb/8u
uuivluTaVC6WkASPofL8eFhcM6/IKC1oPU6jYnaN5HQqaeBKLJsN4r+tEtOYmCJS
NGgpRazoEEkkk84xGiiJEXay5rtqoemlfoB7KMnCQDPsSD0R3nD9GYcdI1P7Eahu
X332LyKnA8+SabElNNraIRzjgac1R0NQPs0NIOaodUpm7TIU1Vq/fKMNBN/BwYg1
2mjQfJ3RpjKtSvp8oXWH6N+scirTJpY4RkrzwFY0jmwt5NOVSoMrI+SHYskM9n6e
9zE9jIu/R9r0RnEb2jEBtsENN3brx74ewE7wDxForneTidIGgSctBbCMf55+J1Lk
J3OmGVrXg68V+f+fGXCs9Rnzzly6voxa7VxzV+QFDvqxuhnPRk64wi5uDNsvRAp4
F+3HRyxWvSDpSFDE2gjQxRWk0ydfjlGvGOSsiL6bbl773O/Xu9pKAOulwQUn10Qh
wWUmR9AFgGoIWBHXrV1wxa75HNOE/9GsYnxy+p+abZ6UHgEG+rNaygHotPQXnZKM
WoFxWfdNvUimycWf2vIHza9xucmXTKPKreXSkCzf824Iq1WPnVgWuPfQte/e/sW5
bkHuL0J86gYsorH011c9MJBFCepXkxbOqXtT/N40TN5/pDgpTSGh4UqiCUCFM8ss
KwNyAsVTgQ5z6aX66prLa2Ck38Uyh5cohwPIVYxdYQhPSmuWh37j/oBBGj2wcuX5
xJtLEpPsQdqHHIe6jk9F55qPARW7eWSrZCJN6GCGhdAb6QkGEJqNx3OggdLVu3Pj
tdLPp4mLdVM5Z3+oLJ6P1DWdnb1j73Y2vqACyPxq1uQx64zVAaiJrK86xtrXkCLw
arbOI5km6sx5+RnLOQVfH6hOF1H7Wk9VgqycTfX4DteV1KorCRRp1lq7DeJIfwIn
d5NKgUUMLCngUjtQluaibNqoKsWmSqL6y1K/bOFbmRHJyv+qRAHNIt0l0hUwLs7L
57S024okD3NsMTmwCED5j+pAanU0E9F6qZkNCVasL57KonV/H6RyLbcxl4kDK1/S
mDLzCNBBGEsNdi2ZGe+ImiY2GTT9VXlaLwkhoCkPmNIFlQcs/8C+p/TeZm3t5n8w
qFQ6DxACTwmRVcuUwwpeAzy6lbgNG8Vt1apCQiiqUlWr23ReBthPDmcWMwQn1DMw
ZTJV9odiBeJ/3Fd+aftpyGELBMpPw5kAqY00+TjG4M0NIpdtaeFkVZsOdmzkawbp
k2LmF0ojupg2nUMzGTXJVxjsQUI4MKowX4TD6vYlsImMJkVlsHSYAd3gF0Lx76Cp
DRXwBPVcPLT6RmBK8cJeY4QPnnktMpWSnI2X1tuudWl63H6lOz4b7bVkaEXe9uha
W/RvFfxFBb3BIz5I0NpiylBvrD0FYVL3JNKwTs3VbeF1z9hsRnV5uOX30FZETcWy
7wKEww3R1tet1zvBJ1iH7QyuYrUgU6qxTGVf/Cdo7E9OZHyKvoyn+uYfzMi2PSGw
0ZuUXI3svEO9vrTEWgcQaJ/9kfO/3NnxeU2ikfTd4rWLdY+QO9NQVTx06KZbHtx+
8XNsLXAVS/HxEEMXPwwgAjF1osdGhO8Bx2PZ1oJtXyFI8POKzUiucrihcFbzma/Q
vnSuaKFvLDc/rLcGdpKRIWXT3idlfJAeDu1ysxmIrr4fLmRJqZm9gyxkmTu5JBqg
XPeqtXfXXsljaoZI2jpb5Xz0uqmbXs0Y4fNEDreYfVf+aahVua7pDYRRvKQStqMH
OOAyni0kw2PjZe8ufit/GTCBW4hels0yl/Acz3gU/eXuDHqlmtYtFKZx4ne5rCTp
XFzAc1fu5wFg32qEpA9sGkWj8YHD8t40oLZSAuASYY0W39lv98GGV5lBh6SOgYUx
R1niRKAgWJ7jAedPJHo5abNdPHFt1XeOpNn8Gejdiwzqx/fAtXBjicPveEgX5ncN
EFzkp7c0627eZpQmZLbcw3bB4i/k0xVU0OmJJU1rqukfRkb3ehzJ3f8SMWs2dHV9
FhLz7LRrmm9o42Z96voF/CJGWuh9aceMZsP4IB+V0rvnOtOvDwHEYnPwpKC2LHtv
clWJlEk2Qeap2T6eEyr4Uq6wiyabczo4hLlE0EQjTxXcwyQA6OKToyMClNvce+yr
HeYFahUQC6QIqfrICx/fyjbmY5JE//Pf194IW1eWXN8eKHpbH/h3QIj3C5TSmN5h
ij37iJR6XRKs4hpBy+sLBkBtKYYRm0WBXxEZGaEswGMlBPta5I2x0fd95yc5uZTa
XwyageCRxmISOdS9w1CIGOO+L1Tlq03/qxreVPO0zI9bVtDttwsJdtuLO5t4224L
zM1dThWXrCZZcGD8EtoqJBoWRkaasfGiMxvC+9ofuH4yU1FAy0hbN1HjvXvrEDVS
P4KQKdxR7zSlJKIeXeMr2N9A4LIbDOOJgTj/FTkAHXY5WpWd+4+r6afwZmenFcjE
njIADeRMEUH42cawnGRIuekcEZLD4ckjHEYvEcOAAmihdXLKsMVyUpFP96rOKlr9
CUlQe+WEpRDB4vK8Ag4SAwwVhdC7XVMwlsPndUWITmn26GAkY98Qcly1E9rd3W6b
wtXgESn4gWgf2FaGGxf2Jm+9z0rDI0D3KGeaHKJOXllvTiPq5rDv05t4uzp0zb/n
8Rh4UPZDXyMdOq5g1Z40au3G8oR+p/y0y0vWcA0Wzocp6Na0fDprjCzeAG2j5hN6
tz0murdo66a8ZlszyJUCKeyJRXetamYl3FKOdqXb9HdDP8YyNPEiz2ZE6TLWPfXU
k8p/wrevn9zXFrcgpiMjQSawXUTz7FeHKHBTqY8fsPdvkSpy0fMZJ5lM9YRXvkIB
7kmfM+TEMXPdc1+B7TyXGiRco/eYaDnk+3K8G6nuu678rlF1wXp4/qIObaQg5UK0
7pCA6UPagUAhtmF1RuO3ux9z4wGPQC6RbDkke7pBg1Y97tK/Ha2HTUN1YRw+zMHh
1yx2FQew8x4EBRuFe1wKfUQGD6MT1WhBNUZesEqWtkCFjTxK27d027b3B0W69wW1
794JG+WG6FYN2bGDuazX871VNAKd+UiS0Rfq260kzP8rSGKYr5H3EQt49ArVZTiS
2SG2fjvao7kzizEqr1rTffyfx2jPv04xMyuF2oO6kLZQOwjaMoHcMQIHg7OoKMxD
/9Hj6o5GPbVkdbU50pnXkRqZ4vN7EjpduczRWi1W499Ev9DiVrXRcuVEcYrUorJL
Do3IBg6WrrwEf2KlY3sNWMulTNtAP/LBr525Y8S8DY0motNHel19sbm7AHhfZH9d
Ps8UeDm7giviydPNPiFCjintfWgCiLeyZpSZswItyxphL1eAOe4uYt3gKKamcH3w
mF+bVWy7/2zxmSEwPXznLzkHpW8U+/c7vp/qQIU0+Ub4dC+dfiT/BVTSkn4QYc9c
ZZL0X6MCbzLWkNwYMBP7pL3+eumANmv97oQD2NIKDS2zIZr0QBs8V2dgHrx8e8BY
oGxFw+k57ZSgkAI5iHPmga2M8/5tyaY/hhKX2aoMJA4D+WLJz5zhofzpLGiEn9z9
6LL9uThzzIrTX2ZyONoLGoqq2MPB4DCKf1lVITC5vDcakQkgD27sVCxmL1MbZe+0
fGUQMvwla9sWOH5gRi6E9LeKBqrsRU4B9jkXrgKb2YcRUZgDC8Gz3/JsyaqwPITF
U9ABu6I5E1/pavqDWQmPzcZDoevi7i0yDV7J3Cl1ZuB1KlYBBNgysgJ8Cb2ksrSE
cdupty3jfTu3ouSP0hUDS4orusB7JzUWnnXATfB+L6fXajTFa6E8+lAkJ38QRwV9
xpwVy0ytIBjAPTJD/2u3qkYwfmL965sgXEIaK7ectfTCri/vU2jC9SX4ayau8vZ7
QKxWi+j36j5CQrHRbS+lhUgYyOo5prvrTrTchCWnfTMdRQd35FMUOXVXTUhUkT/L
/ltVKpanK0LZqyMGB6K3giQlrQaEayYjdVaKNsUMkInCZeKwas8VxGzx21C3tPaV
RbUoko7Tp0hU8VRzI2wTeu9/gZZ2Boy2+bxGgyAqXNp7o6QSVKJMgVv9lCQVBEGF
DefcKXoYXRVwaojXowOWtv6+OPvk1g7RIOOhIT+Ruczh5VHYS3YsxJyuOhN4SN68
lIZkyut3dUC9pgSfEEWHuO7vH6wWGDEy7AiSnYAfZ8y/ByvrrT4uENSII2NxfGEt
K2GefLVJmA6esIp+ylSONoFww9bwMOHbmt0oRbU0G4ASZRRww5knWP1pBAJ2uHrA
jLyZuyB1hvGnbjAuaJO1pOycrUakb/vFX+5oo/KPS5QDcSXO37Bi6Urp5PqxzPl7
PMba7PmKMJt9PAkUX+zRcs+W/cw0VofCW/qsXuLYbfXf8q4TuJBYeGt5HwG+uBPs
LaksEAXMCRiRf1U0iM6OghzkoETLKNhzlAMIazXevSM4wWl/Pntzxe37oy++8ouM
hHQC3wpI6GxEuRNXFv3wb1RdKDOv/ATJ2FMd2yuiqJz9KZKoFiXawTykRLOVumzI
fxEyUxe6encGisoqyjbxxGdUDRG0KPJ+UD/r/+EikxDevZ2oAImVjuyVKhPW1mvv
EJG0Eed0Q17xIkLgdGg4lZeZvlKQBppHgS7hT6vze/d7tfpfEBOzquj6qXhcodOe
xG3l84jHQvDB1ljk1lFUmrHp7H/9/GKnoLD+1Qqow0M4JAVbqzjQf+li0Epg7M/x
lgtaDmmeH5DQWkSzkbKMUdciHMFWR8VPquexsDza42vCwsxhLIpfrGXp+itaYDuM
u3T/0jdghr8ukm5eCaObiZ3HpMpPJNDbB0BntPWkApkBOqLX3l3wrJWIfrDqvFid
e/8ETgLuUO2EYoNJ2GvAD5JMxfWa+T9S/p7L5jiEApK9BJYBpd7gzhiEkJ66hDhS
Vyc56wQBTdsxOdhFe3ZPtSSU/hqRP8tlt5mO/GEfdrSUZKGHl6ix7vw/ZPtmBRd1
42Q1UlTWQpyEvV5eBp3T/egcRWVHYiHsh7XDvhzU4ohb0NhyklXOSAhwER4GPemI
0yeUrtEmvonxPqbDnz7IwcjM5D3HmpwF3F/sNQHTVp9AubS+R8CMKWCHq8fyfVJU
3avjKMXJ0o2K3B17QdPiRyFFUwlkMpEOZkcpUFEr5Hsk6QaN9KKh+JKR0M2D7rR6
LBdyGqGDvZ8I39uWUhY2qYy1ZJfLkUKqcJUOQ6kWdvR3gMgBeWj6dat7Q6qHkp5f
StFj5+SkvDBYlqHpdHSJoHE/yhsqiHC+8iPGTN9qLge25aNH0vp16L//XeuPQ4Ff
P4I9Q1qix9VvB1me18U0tN8+kGd4CyeXU1Uo4Kn1vlwJ5etUP+LPRmLpBhOuVQsD
hOYAoHDzyPBcTvBFWP/RpqBCy+cD4fBbk0fQmjomLN6Z2PjB6trxJsFO46+b3RrL
MkTvTTETTSGwgqUjZqlyp4NRIxqzCG13T1uWqPj10zDL3Eac0s0YCQZxG/c9LYnE
T7WYPJstXAxWuMDj9FBL33RxX8MA+cmFDNjE7GImNcOCJ/SGN2zypSven0pDjb1y
Pf4p1cRAT4qs3MnKzUxPKxF8/E8/W7ohh0mtcrH5EejFqAtJ2JChM0G8+WPS+Zrd
0R5pGX6IJ0btWHknTmmuwkpII9rT+aEuHs+5OW61eUtw1sgCDB6yKvS9Ns5b4uXm
u+C2eZa7hw5/TrZxdFdalQlD9AgDyv5Lgf0j75vhfAjqcpZXJdb4aQxwfqIWMrIH
cOq57JtBnsNpjDgwmn8JqWT135iC7pH+EjKUm93D5TiP9dwQklnPgJ3ZyvV/NoV3
l2wfYhsCbAEAujGSGRkCu0e4h/i57Xuq49iL2ElX9SMsadbJdOKRMSTfYmzefOCf
Ay/51ucfaprc1m5Tcvv2EYAHONxOQHvHkWpiot3zkEN0UMSUa3anVX5Ro+M1FzdU
CEYOEe/CVelcVNc/hx7SiFk/SEW6ZPhPCvZrOsORNSuH00P+8ecwFQ+EBXKONwXn
i+QTK0rAI9MP9VAF9HJfxmHsYxCbfkApxXC6aHHP7fwRk4bu9tWX1lZAdFMAHMvy
G7b9dU29qZi2bHtMBVSHEmnUwGlxL1FW9ciiwS3W6R4+HfevDXNxOXxUt6lvnPr8
29iNAfOSsc1JgUcmrlW8JblTsbamNS8UkpGqeCXErGcoiY88DVq8qPK2yZPq7n+k
AMLytYGkWPGmOOnMounoMyLgYxzUywI27UZ6AAiqbQpwZYEEX468RWCL6hyXTsX/
8cbpRQkIMZYhNGfqW7WB9oyGbtq5QAf0oZgKEX/A6+tFGcKeyvDizZf8MUr1t9Y1
sqSGK+r1aYly+xlY6sTu4mx5Mij92bg2+NyTOEtuh8E5IMGhND73VLKFcSSweDIJ
++a0MltzTwPMyD9itw0Ik5KjFDNFCy4OXAXD7afHZDtabgpqvNF37BFT5rh8HrOq
wE/ScUgXEiiSmpxPS9BErVPCJWW04AbsUh26tesXpw8rUPZC6Q0Ab6LHQYvStBrP
xOvg7E7Ch5K1VlcsSdMLW4+sVs63iQgQ3Cx1TKYpG+0BV2sUG6sR7PmnLF67bBGd
b6Kuq7C3ZoCPOTaCqIs6XH92+/RTnX+2luj9aOf20qbOXzbyIPThwrgQt88pn5cc
INERZazglwKB8NO82TEH5JL0tAj6NaufDdVlYD5Fx15teHxUOfiwnjtDhV/I+q4F
U7aAy7HamvgfBpnIukjl95aynUQenHNQBv55Phu3LusRsDo/fk8/mUk6tqK6jrub
EpnW1DQm3hjqluUP6NNK1q7up89wl8N6mQJN4lN6Ig4G2u6zo1r/GiNegz6BkDAb
HtUYwQDAtQtpv79wR8LpfqtjJbpwQSRdeXxx+A0/HejKAcY7uA7WQHP/UtvcLXQB
5KFygYMsSB9Y+2C7Lez401QaPIUgAmcXEVI4ZMjQ8gEmuG9BU5dY4JCtNAGSssmJ
MrAYZ69EzYEa4PEz2CudxocuLguvaT+dSIyv1draeEgXk9tlNrO3730y2wvb89Gs
Mnktiaz9l3XYrzz0m46J2EsbTNHX9/mz6cbxDu4UxpFdhtCjXqpNItEOb0DSU6H7
bzpru37T9hJywW6RebD+VerLP6xv7zGoDxaa8aRDPKQtAqle4oP3AcNBil2qaTOa
beCXUb/NY3sXlN/xiD9WAsUPEG3vC7nwdcaZOik2fZxP6tzhJK3TWJjn5+wM76Bp
M2juYmM4pYO9L1UT5vROrQcvGimSyvyOCnqNvIY0Ws7UuTU7IisXA66JVxjx5SNN
iMXiDilsIAK7Wzh+RMalCbrrrm/mFUADJwrWyYArsR4haNXdCtz4IH/3OUoHwOGq
YV1lHxH8vgmT+fvnXmWgS/wyi902tJ4lyVB8ddllbFO5C7ya5Fekh/JwXd43Sfhr
vIbBG9Z3LrnSSQpEa0hlwPY91ikqqIcBnU4+6qTrRHVPVNR8KYgUzEr4xVBhevxf
ZeCiheZBwLs3nrnVyA6i5tzHvXLym6IcqyiX9rOa+71cz7QvAAtL95s61cBtAn3G
EjG6GEBuB/6Hy2O4PJr6qm1ieGLSCzPb+L0GX3RcG+6HF9FsogJoYp0ihUAMEdch
cTvUNpw5qq8Zk7uS/eCtnxNLbcR3I1pfeQlTEetCpN3mR00T0p2ANA4xdj8J1qMU
oL3FZQBVN+VuJSptB54XwnSPcbfMImTKJvvkHUyatr5dQOtdKcL1ddj3q9PPB3vs
A++N+VUR4bj941vxi3yicMapRobp+ZA0M73lWooJrbUCWzWbZboz9Us15mpvq//x
hyjAhdnFe+nZ73hhGyXshLQYUgydMjnDkr50zCoRCLTN5dH3c9YkLzlXc/k9BDRo
JhRhcburhfZs0X29f7v1Faa39mxGsX8Km7Q2d7TX3beRkChsJI9W0qIzvdYPdzvg
LKKiOUZm0R13Gatle9Dkf+17NotsjD9plsV9mv3dcMMkdH0FhKIOb7Tn8ArWbQt8
9xifrxPgzMf4DSg505g+KR902LqfYSEmInzMnKRQEIrohOOgc4ncfxwrVERIm4bT
VLPWgnLoVWC+Jgb83ywDTzHIMd8NfM5rjJUPkfI0piSWLVcf37Tdg6p0iwfPqXvx
zKMko2otOM6WEivr/Jm4hF88eLqO9AojrtlI6sZQqbcxC5yMtAreXhzpXPi3WOiY
m6kboobLoD7n8ZS5oiGMbtL+X3gxLAy5yFXyPJ0gC5vqYU7l+pb1OguC63VXQjmN
lymW03pjoprEFoT27z/lku2IMgUdHN+dZOiEHSbyhVZepQaHJBPsR+UOmFKEQWNG
1frRbTfUFv8WOiSya4xtQ0j6biv7vOYJYjK4dO8trQzRDA0hObeUokB1Ic2kzVIm
2ln8/JGxWBkJS0bOzDoSHW6vIDV4w2hDheYlZAelEhAnTMH275UjGRz4++syXWCE
qSc9Dqhj5/5K6yHLfT1HwLgrO6mxSRXa//xSNSC+SjXracGekXfYqSnW8klNRS/o
0ACezgRdp6eNq34xbJbPqe5V2qmkpGdNDX5v/Jt6N3aoj12OOWjMRjt1AXoSssf0
IDnZNhokQ0WkMO00FnF4IcDuRxG5zTmMJ3vw1rm0YGmjNSwcpCDIdioYzMojBLcE
LXSzjiweptiCz1sivBXMpUahz/szFaWZTctsK6xkfoHU3VtBrEunCbDI/VtG74F+
hq/wE3gWRrBAL4d8W1zKnTmBJpO8oaIJQGM1YcN6j7Fny+yPGjR2Who8MHAkJdK8
mQPJB4ttrI+nhbV74wf/rIm3x4ZqAXT86wWbpYLQX1KRTMG9q/qGGewcBG0oc3hc
4PNoYnGTcGskJsq3GldfUNOancUkr1OUWxMGs7c4P4gATISFDqfCebp9dR1GW+S6
eg1diq3NqYaCkTs6xSXw+5Slwm+sNIdiFRdoHaY/AFWyjK2WJb7wopGrXpRcSd9d
TzdJUjt6YQ3syQY4AUVz2VUytNJpo5Ebxmeqn5JYjgt0cVHpUVy7t7E6DSC/E8SH
5BZZGcRk6N3gSOeehEwg0gFOeYwN6laO63x8Op4Qf3/Wf0HR55rAN1BuLDkMYfxH
se7CiJwyMVMEiBJkaVcUmwgBIhD0umEOv3VSXQdOjUQqv2HUeOM+VBlJDa+XIihm
ugSdH9fFjsxn9qToQ/tloxYIrOxwBJR7foJ4HFsuH8J0yPHyebU7RsOyJ0Bbw8TC
IOY6MbGxUnd9x4zED3yTDX9XzYowxPw39IkojQ7/ajTwFsxow3IONHhCZuWPFqED
96/CdPcMRYFFOeW6lzEmtyd7mkPuYptmuu6rwByuweGqQKS9lpTdDa3sxzwzD8GG
i027mPZgbxU5/EmvWqF1+q1bHnV9kark57Tb3vdxXeJzOzZSk0TQfvZv2SMStKsj
1+yyanbDXjJ0JESJATrvb5PRroSLrI6TC4TKUjMu/P9z5x4csS6ZCGhW5FqvVBTh
9sMe5WoJ+qxGUc+TuGtv5pvovwSdZKlSKpfoK/vb7on7Z47d75AohCNh/OD/XOAd
Uwji8M0rW3CFxrvfo5JrksA/LHdizcGBwcYlTUz15sigmbH9PUzMXmfRPRswRRKu
MCc7t35waK6myASA2I01LOOK0ahOoztjIEkWWs6lshlZUwDrsVwzFfEH6ttc0dxn
Ay4RVxhLu9FLPabUBfc87iNSbPIdGxC4EErmGWu/IEpRst/Fh9kS/eH1V6y2eaUE
DcuV8WGHCyA8XCKEwKsmf+QUgOop9uuSxD2oyieWdWjkMJvoFrux0rpGmkNDLsHv
WGokSnaJ9cBIuYyCzkviIynbDTHFkwPfzSJKdAf7hGsTWD+yLNCzqP4/7QK/0rMC
MzSkqnq1wU/zZ3rcI8OhY7uFrQs63W/wT8X3m8a1J9voppYzSlz1MFO0abfUzdhk
F+gjl3gvPjc2bsYnQCJFMpP/XU1Ml1q1YIan+3OlQ0zd8NAKMvcXyFRYgG75FOyT
acuYsyKKiTSMHat+hxHHd7rGMHxDqm80N72zPq4gtOFjV2iPqrL/ugLTlEb+k0Sh
RFRCdx8B7Bt+eiONeo5apVMTdJqRtnWOvI2LlwQ15xixiYnosUy584b/wtEonFwN
yc6lZOZXElzlgY0nGEncTU3KScaHS6yNBcGj30ZR7iXjA52dZFYSU9cGiIsv2GJQ
ntXtzTkv5cyEPXiMwl7WjUG3SHvQ87kiZaVSmPq4HKoT1/r9/mlqTIbsNjjyhWLE
SIsl43jy2hGNQJrp9XwKVfKw8S9X8nt8y9p7qeOmXey6mpU0us968KFnqmhseK0A
bbuX/R34nge4VBOpGotfXtJt82a0hbq+UCAeIvxk/gGPxj3u9ZI/Vy2PhswuZqem
EyHTV7u7BJeWXVKNvYNz+0riiFgizx8MUOZn/pfma33oHhuqVPxj2MX0/9OeQd5w
fsmpH9c9goDEqfITYl6xvQtOAhx7C8aozH7U8tAAH1w0nSI9ieUv9xjZmYBrBiAC
y8iHopMV8Tlt0geWxbO1Pk7wCC+joCUUIrSyDCeuxqt/V5bYzHCLeyKqN6Pg2z8L
vADGzRJKURgNrf4hA0bvhmRI/vcczkmPuOdWsAy6Tm3Z6lYFqANdVgTthRFqR3ez
LGq2Hsh7td8OvAmpg5IMmaiA18pOc2JL5aHPGihv/GqP9L+DKoLZH2atqGJr+0sw
rJA+b+znuISQaHJ9/VAOn0YiwLHG+ZfNNKnRpenDNTHVKe5NBINR4jmCgsb1d8p6
D6gVLSGcyRrCIdnzdPcBJw/lGQlJt/brDA9Ko4fBCTkBYOvFPrpXeB8SnEWmyZ9I
rxuMgdUwQODC7r04XWV7Ry3eIQYdFRjHQb29AuIV93S3yyNlvQcr6l/yrFQbZCm2
YNymuXXlhZY4ev0WajVfk8BsZR7/6DH3aWcDR+pEJycF98dpYVPpDRS6x6QzExvT
vphz2Wzt/q+mjRlN2+hAiR8uTiB1fvYxiYGpSBJ5FoFlnjLnqwvnXHoUy4PGhsSx
Ju64z7CdZ6zB9g2FVavzltyse2Bem7hxUdhxAMkEGLRzOCFO4fTyeZlnEmjWBJTK
XXrFSMyiz9BmeKFVipGuu73cSym20fNxUMUhe1v4uBHpGnhrHpYfN2dWQrcCQl5a
l+pzkpd6dx77cneZytpm5fIGvnFfTrjoj7rQZmyxtdPWkS7Z6LIkXXgAKMT1kLcP
0ADnCrws/aMJYFNa63jHuYESzy/cU0LlYP0jb66y16u918J3sbKPv3Koh6ox6pB9
9qJUDbXHaygU7+GFVBt+mN1W4e25J8/tAcCmcAnuHfhEZfNR4YdxpqjJggnf9wQ8
fpdlvIZTnB0bCGvf6U5Xqzu0K1jnSKqif5WfgpUt3abc8WoCTqN7npxpv+Xx4D9i
mcJaNhFuVOYBjznvgeMzc5puVW1a3G2VKilkGmbEOzvVeqLdwOLzNghsmvDQde4d
K63Zk3Fn91UASOeSaTmlNUG6HQJWIVswQ6g6O+orhBQSr0HZoo8QkxwE2CJSamKG
Lh0PWfmJRn1xSCsbDHHe3KqHcakySk/BNmMOnp6l2r0P51in5pSngdyOuNZY4xdH
mKGg4DccpvaSHQ0Pwv5+HD9I/JXoVXfAA1CBOk6kvrhYktYuWFryEPn7Dbl4Pz54
iFiq7el7xBbGsMytHOeXuyT1IJ0MkB6NNhnDtW7ofAhyC0wQf71R4oo6bAjiyzDw
gZhqEx50tgcIC5Jcv98Kf0PQzO1UyhpbTqYG6Mx/YzosCZsMs0MGJOKUSAFWvYbU
0mEmhX67Rk4NaEu7795t1MS8/o/juEUQ+G3Ry7guqSHS7qbN3CTtKLYFS8+T6iXi
Eg38QWjdbFl81O2xGLPV1sC+Fay266FsjFMy1Ok3nWmSCgXdnlfwp5BOx5pdoE9d
aNp+Sv0ovxIKQjg/M70sQB0II7jMiZWBFrbvF1/mMgdaSWB0F8EjaJ1gVUp92xcD
NiRf8zwRjC4JV+ULRZcatkFrV1a6BDadlIaYaWNLp/tyhftYuQNzaaivCc3Dz/PS
IAFOeClA5ow83QyMImlLQ7y8wBxAbsSJs9o13mqZk+E3nL13Ngs37vErX6rEd6Ak
mOQO1hGJZo6+b2A9lSoXZxgP2AyQVGpTEJkp+uRFKiBqq27g1o14BVEyiIz2QN3s
ywhbzeiWck3IXuKUyC2rYM3bVwQHjeP35ZiGmCftufezR8DlvuzJwfLd7yUKGhIX
62xo9ixVbyClKPY1amf2ac9SEpdnyw9hLAnqFglDWtGv0kVmNSsgc2UoFbsUSd8I
wjqVkN60J2YT/fCrqNMpgNw5TL2JXnWoMq6X20BmO6NGN5SkKHniexILdKEMgFh4
pbu2c8d2ljk92TBEPHzwrUHhctnKeOh5MGffvB5NhBk665kT+h7YeZbqAq9eFALn
D4caRFgOIO4QLC7bPafo1s6zPwtjWFm0vFKygyEoBUYgG+ZQ5avGSg3y4xcAsMmc
3rYe8G8c9Agr0tear6LC+/s1/45WveGAX340VmvugloH46xJM4xbQz6nJa7lOOuG
PtbtKPySLe4/lvtCcXIiEMdzxwn4c15TXLCRqknc7X0Ck7xwzz/phPi8rwKymp5e
CjhNzxZMoVFpa1USp3cBHcWraCnQuknJ5Dc7/J5vpS4wCs+41nCaiygSrIU+QTBm
IbaD+7/oaCIi9ZL59yQvfSZ4i6SxSQw8v+6c+h4EerLc3bxmsOzTtoMosYORgxe/
LEsJb8IiToh3uXZDhsANYm0Y1zZqyqzWbBHa7PU0WWL0RfEcOQCepHLdFlH45jo9
LzczYrvQwR0BVYnqXccniIE16rrNBz2VOjL+N1UWGLgCBg8qOCC0QpHpdDYIBLAm
9U+kQ4QnYGctHij/vsADXaqS5mGLFEdJul+hDh6SbxCvqNsTfhfqtPy6cOZTontd
bZaRJqebCQL3D/gMdEtEUaZLi/O+EvuIwvVnQMGdzaAfsSSlu1zrBqu9u9iVD14a
VFZDNhVfTxRQI2qaY0OiSd0YWdy7OmYtHK02PwyEZ02dzLRFws6TONJxpy/4dexl
N4AyOuQ/haeml/0IdnkU0wrX8a0ScdeadQhpsJxnUQtIxedNpM1a5iaZk9AAJkDq
NkSccH4u0kIaVdSFJ995wnUoNGuxgnk+5xrREB6C7eK7838oIYzEClYtehMVGAgh
wIrkhq/QenL7jqN9hLMAx8LwG2NHQrHW9JKdBU+JG7eeANOhIr6YO0TqDIHWcFEm
S4rEXaf4RThkB9c+Z8GbHEvaG4Wp1MgGF/zj8CZdZiYFFD4YkyatAjmG0odOV/EX
LzzgA0PUWUit/eLDOmZU22s1Eng4hEn9Pmy9E1zeqCeKKsoMINUzKCmkHD6VAkAP
/u3L2WpuOzXmWMetlyFDgGJ3U3ppHGwwMgnaE/zKteMrZOB0g0f2PxweIYjIKafj
LWuDu1CP04V2WPaTvi1d93aONrtZzlD4LfiMLUHzOCtyRYp3K0UfwCXdCAt5urbt
vWL5ME12h4S4zKBdoTZwD9Z/lLGSyE/Fwoocf705/iKvaNf8M+xEe29IEaTrrELr
xKY4BhDItn/AtYL/djmOuyJCA1OvxXBNxqD2+p8tjUt6vQWkwcupQ9fgouxRq0XN
kCxMGI4Naf5WPCZrnVyCi9p/cfKHjWiLkwzNkC71RYVPAiVrhxfGSYCLeUEmMvze
ewmJOMpwB4Nmvg3q1AQ3yNapdpVYm77wRQqkkxLeXtzU7H61NIb/J1016ZSUncWs
r1VfqY53D3u3A5/AaGrpHI3+DD7e1PndAACA/UvQuUppmbr7wbQzDem80vOKHORz
MlyWkTZFXTMMOkFEY39JbzD+iDh0C4P7guSkYVBEqmA03LRvfzkkjD/9ss1kFaVA
weEGSFSI+PcaYRVrCRIhM0UGi8rfu/T317c/h5Ch+wPlL7B45jeX1GMMe2ujTk8S
31o9zHt+Zt5HB3OCn1WStpSWzyBwLP2XEJ342SaupOB6XxB+HlK+ZaMI0CtPIEq/
VKK5ODtoPAfMXQ7ZjudDpNoNn0fxLbeBufIPOo5RFWRHfcoXyH8a4uUt4E67Laey
JfXIo8ltC3k2McDA1bCAcUac8K2zTpFQZU2w+FzMIpZsKUibbzQlBb1mqDQ6daV7
SZx0yx9u2LJ9PQFEy5cyd2z60F+jI3wBxg0ki+o2LTB0T6GKfOpT+XTl0yJya6fg
ezgb1JEzkwzZQ5slsCDyYDv1VpPc4sSmrYn8xFXr7/wvKoRT4ZyKumwLYMblXLt6
YoYHYETJx2rpLJHkbwyhdwZqJjt8OZBLDz41R8J5f2CdP47xHLlocPrh0YSJCmme
IQJb01LoqXE+2CMHPgVa7oq446UBHwo9J64tLPccPQFZCvBI+IZhla0eLwdcJKUh
w3JMVFvdALdnKlAaYWjxn4BABfTfKoK+zOJeTme1N4UfS+aI+T5adWZWPmhe+fVN
UEcyjpZ66HVmLm9DA6m2bjB5dFYFFLl04XhJ7v8RShTVt71KiAtkTdk9OrEaFhlc
4dqWTjTIn9UFi7/aFVEtd1A23ArN35+E9DXg3fBKn20i1136xiXueJ+mgC1WUQte
Wsvew5Vurl1ZjUzE4S1XG3z+1HYyefvIEYAYTh9AbPu8Gbv9Nr7ErlpJHzeyPUUG
ygtsvYxUkahGIQDX2Ni8mkE5DbFOOh2f6NUp2PV96cffzx4WX69KaO/ekKrUXYUf
zNr1LqbgPIgp3C3TMCILBAyj3YZE4txMaHLe20Vptp5wXJN7P8/Fiq7ZlrsKmcYp
E6bXPWdvwuCX+NqpCCBv6DZ7nNoU/c+WKQ64W9JTcr5apdzrsf4J4BW/Byyej481
OQnG5wCxvTDHjW3o7nNG8RXUn86xn8VfVVgUS6cYkLQ2ZfxnnaRCT2BlYKHPBsYd
yUx/dT3PFdhla/rcrEGFz+1hR5cd8p64xTu3yg48iCQ862B5jzfrjHpLSR1AuRYC
elhgRWgLRD8Yu5WgF+WFYmhYpHPq42t4VfJLdsksUE7lH+QomMLM+XKEdlxt7NM4
FJVRkR7M8ohEBgThrSA03644R1MYUMc4yTREgVuz6ctG/PPs+5LYfQk/5W91Ul2A
y0aDcFM4kq5fmGXNFciRmITstX/3+xemxiNmDg3pOEc4toON9ike6I0ceI9yAMXp
P8juxhplc1WIClnR57G+g04kKpADaxBijy5JUPtx8vjeXPM3Wfw+IlUTxXPt77n8
L/Kj44kfotPuN9gydI4baJ2YvwV5eWdpLkTIn6UWXU23rV/3Gysoc/Dk/3YbJ4hZ
THBFcs/t2JLxr7LynobCjUN7lLhSlsKAG35EaysHK+C1tIOqmFoW1gViOJQGUeTD
PJJWXR4BexuGnGsbjcRerc/7uSIPN2A/ZjTM5fIXnUG7rHsgFk0CGsRs7g8rLtC/
8pLoKLRlbcyF7KlN4Y/CoFFyeYWwNIWJsOaZ5RaIdnHsXcDfb1M/azne4orzIWfp
QaKpehfoa8eRvh3l9kDHqrss1dSG5dy5cjQKeohxgY3a1sqFqKvJ3VkObW9rSnSU
G0/G4aDLhbNu3RaBomOi1zgurZMzeTT+SmgdzLhWz+QGai4wKkZ9CIbEK+YoLv4F
xK7PsKhPnDiHVLfvXPgZMPiquc9Mub8mHH3n7v6/EJZnctf9sBnlPmNORK0bDXV6
MBRrNfnEhbtE68LyXluUEGhHMvnEFIKpPpwb/eA1KbhUwwr0wZgtQxplEr+6Iw63
kFx00IMS1+scyhBG+mId+AQ7LK2Mf+B9a9lG808s/MbXlptgMxonGdgT7PYAYjHT
QpvcOxKullJ+pqvsaaVgg9jeIl+IcJi8PboPpAFQX4+Nq24JQz28/i5KBRtXeNps
KggC6YoqNYnXa8+Y2CcT7yzG5QGbC7etfW0uTHlLIW/wCT3sT0afFkZfHMiYR6Db
FfGBhzb4OsDF+MFAlmF1fmBNXnNknQ+tUx/1Af2A30tbsM7dDQM7JMim3OLwazct
GV1KmIDJUelrrSa3oTv9Qbgb+MZ7yNNIW7fQCmlkMbwQJud2/71qFbh7JOOu7dGB
NJ+DetXhi1de0zd/FsC1oY8GNHBGAg96yn9sfOgkYiT03eJ4MDejuAzz0N2Kia4T
s1jsqWcBZrjrh+f0mAOmdUcoGo9ui9hIVzrAjbQoK1HAFrCQULAUmUYUCJkqIenC
0ikpLIqJwxJahtzwrlV9GR3iNt60f2Vf8E33fP2panqpz0dWqWhQJrCFUiAuAian
qwMzxprCtdJZ+DQ9WLlSLqP+cweSWYoU4Pt4y/72HNeLwc/BzKYvKKAKZkP16BuA
k2F8GRnp4H6T9Vv0TMOPjHLfLxHZ3RappLaOVeZolVCG3MuUMV6v00/a/6HXFmCJ
pd2eIb6ts/ntfl131gmC6W28iw6k+ZGCOsQzVCXSO66pT4Rijqr3QPseOpdyWwNJ
eDMH2egfnXEEzvaq02vIMfObCG8I0qK+CFkhDMP/FLjO9IAujlonpWJ3F/mMr0vd
vLVPQpPRJVHktbPFe9FmLazQu+F3S806TBDh86tcrT9JWIVKY1DRbNRJjXKVpRb6
rCeyofL0a26Wl4SXA0WTYLe5cSEMxNSDnBJrprCzBpQe+Zb8BZ83zgB/RtV5a4DP
Iba6mzgcyGU9mGlcxm4/RM3G4OSO5g4B6L6fEXRFbaVbXZUMvbFkfudA4vGRschN
E8/LeKfqcbC/Yf9ovsDpBXhjgqD5GVLa3IHYzyIRQhjWbn/24qqdAE2aF+kYzTVY
6kfQoZzeiUL2fX5err9fIbBYaiz4lNsbmgDwFRtwOJu1EtN9klSrdpfGwl+8H1TP
5hWp0ONwxAHEIGiZCDHLL7ExRXLgEv1tcH67832m07D2516F2uiLB+JDYSXwbPQu
+FQp78zNPssoDijudjDkJU7x2hI3wdXectkcPkKdzGYob0KutINHP/mNN9aOIMpo
UU0aqCb4aAoQ6drMbkEj6IZ5BS6/BsJub/oYSlOPe33xYbA8Tgv+uR7ZDZOJrLBH
VYcnIdggLlU3XC53Rhy9Cn9pczHl94BSp9EXteydDH9d6Z7cb8XWE58wyHf6yrtV
meh83V3nx6djzAX+46uKnjpv8BDdXJnREre/WTwAHV2iUxXjs7zbxAfBcwncmN/v
/8JY4s/kq4/B786HPrzH7GUL5sib1n507i9cCSkcGK0pCjl35r7Vdhhtp7fJpfsD
RSsM06rxRwbdWm+ey+XsNEcNZlLaVV6+rQpn9498SUBe1njvaPC603jf+nrXzC84
WkKDNZH6ytFXWy+shy3+XJGfq+zsI7GOHHtw2ATpvMkuzHMIJBOEJTW/sKO4b/CG
ps5AFlwAbieO8q5iFF5MCadgxcmsNfrCoTVFeOfQUyou+2BxAC0lPUKFrZf+NZ0L
7wGWS8+ikoT+5aBswL9TqwL8fhNqj8z9LFPuVG/2UVMGazd/JqfkVZi0fKvtpgJ3
9ZlP8rBPyUTeCX7keIqBvWij1W5y5Mz1lhty3JHV+70N5fdEhQJyDLAdehXZkfxE
wEzIrzAUp7/v0C6iIjMzqyLtUTZCbkEqrEitkThZ+JgWUi0p+fCszXwU/DxuckCC
fMm0LjusvKOk2qmUUcDRK869CChNT1wNpNZ8Tur/ziFBGRDLTA4QtEwPFeEgknqb
4+nCKNbaHjS8w8DS4yL0FbjLsDu1YKgkUMgOVPp26ePYL/1L9mufOIOWsHNeumy1
0NoROYdmfJWKjbpmT/w2g1ccslew9Iiwn21kSpeKxpoc3T9r0uA2wI0+GoiukCHD
38q/GRnS5Q6AsvqBziSgoK6GMmPTRcddmXqeO8Lzn+O7dH0WOOkCeDTAID/XgROh
onDRV6dihjQL+PmaODPG0f1U8zzi0W2UivdvmXanE6R3boQqiP4Ryr+vuUUYXtdp
toK6pwOVLZEb0VM//g5n4VA4WVOssALpS9dpRH0xax+NH8KoYxHyl9nezk8vaBlq
jjZLJMycifd7wzOCX4PtiOArktIdwZJPJKbosubUrvSCFBCZ0lQ7cjD6kKlNhL6D
0eg+Fx+KFuWo1p7pn0ZJWMd1vIgJtdrUB22CYYSG6lHDfsfHs9dJ2Zx9p46NyP0t
KDaued0ov+TZumXWggVlOHnrat4/u8aZ14m6OvO57m3ZjE9IpJbbM1OwmYk5Ivpl
/4p5nvFxsW4l2SCO2Nwvgc1QUNMXWljwlTYCu21JRla2JwynSgjv515gR2PtJU5z
SbG5BqY5Z7FhwaFn6t7/8NMBNGZOPpWrPkSrTzEmjTMD3vrv5P5Ez2/TKJmD5YKm
HjJRwxmOBYW13rNOipwRxIE9zxWtu8FV0UFSV1S4iBMF4XFkXsWNmces20Zejg7X
1frCA32Pt1/FplaYYzGB5gUBCaFIWM6pFEE8X2y/8+E9dF0WMT9RPD5J0UZrUeGF
HuUDYJX9oZ1E4y0xop4GSkOjfetTft3mAijqUIMXrA0yBCjo2eiNDRbkg2YMP/bo
/A2omvDrzR0pAV06jD5nWPNpoidVIytqNvky2C+Xv6UmOh4Ygq4CwGiQPIW8lUsJ
bhuP4M7yByyaa4bqlMk2hm1ZyMXLXgHE4bou30Z079w/pK5hygbG77w6uazBmZEl
jll9pJtHYdIYIk62nSM4N0LPHo3q1AFf5SiM3jXXUrN7JUNNQN8IjLxNWYMoCect
rPtxgI6CaqRpRnTg28K2FjOKneUQ9eiAlFynbb7hVrb2mVTUVvIch5JbGe9VZhYm
kkGMo6wFupWEQ4uoUPppQW63opcPecphUGv5WiXANsxn1whLXFLsZHBR/CMEwGF3
kzOg37ckHvR4a8Ca1ysDjcanzbKcK4nRYub3Ifm7hQ/3gXrjiv9mEKnsNHMy6jRD
cg1x2L2uPufjdw7B6o47k3c/vnM6qYCPAr8AabisIPzn08JwADidpT65Klj7Igy6
EmbySI2+OrqHzca+hVd26mhyuKSvSNzYKe467SQY998mjOzotMPNkjWM/SvR4m7L
PkLv2WKpzyu1jqfJeZodNUXtUY9VFXgkhSigHFTWoM/luY5ZKei2tlAE6j3p61b/
zc5OTZ2knli58y3MtEqEqxDV1N4rDV+c4K+7/1t+ajmL5lykX37z17dc6XKTN+AB
+/vnlAt53sk383rbPZGPIJhOVXaFNfM/RnLz2kAj03yeqB1/ugG4zkQg6wyOnwv/
CRnXUKtjPaZbSWIIkzb3DnO2a2eL1VS6h3OEKHLrpvMkZ8NBcc9zDgO0S4qHpsen
x/1nWuLTOPAN805+ZvmBeZl4UFJZ8+raDfiDCAtRQoCCSHQTk270GpxTt76+Fqsf
i9INSdnhFJvMuIqGTmgrWlQ7BCjrHKhcgM26HgtqLm4TJFWTlVF7GOU6ZBRFjW0n
A7vTIEVXE69qMj3r7w0J7NI2QlJNmWsqbPpbKGSH1YZhkO+J5HeO/Lux20HNf0hS
XEXEp1f3kM4SLR6HCgVsyeXuMXeZVtCeO7X8fa/pxrxPxAqhlzMPQwAS98rChesD
r5h/lwQ4ei/IhNNt/0Twv1Nmx6dl1D9EpOIGAD6+WREBfxRFl8AgdE4vIaxwq9mZ
CLjKUzbtWCJQzitGZYgHmUE3FmSWfoqpP0OBqrfFDkqanO4/W1KnKe0PVHXANbJo
Ys6CCk2cir8Nk+6ibLj5rTubc4W8x4ps0rQbYU2C6wOGPcF8et6mjur/ITlNzqa5
0NQe1JLHW94clbOin/YW0cKp7gdA9Ren5iIpMXwaalwddRHot67031dlevt11Lga
z8zf8MB4bLhZuWUb0Z6IRoz/ehJRZ1OeXZMo/3cgEbldsSUQYTvUtxVgiyafOF15
DdDbkFXy5GsiKL5nfnlIdAJnmG4kaYwMU9/9N7wNyk9+ugCCooQrU+NAxiE1EdKs
0EPjJ5cO1R/qKwagPQW23S3kZ6HHz2UTZgYdr4rJpSBw452NItS8P4607wgr/AqK
X2dWJ1nFHPe9F6byQ1z4PbgRZLq0zsaTv4XXbHT+dasRouhcSpMUADehj2F3g2Lk
nwohrOL1ay1qqvVXkEHIkCPzPpxuPW9+tv7kFeIecjjwnf2xHJjPFsj+hxHpQf+z
detccDCjNuve4XcDf/ohzfLjHMA/hbuD0KHUdzrLmVnI+vLgelW6y7TQ+J9Micz3
p+GsBU+VMpRBW+CsY7wR8PmEitPJTbNiFZKAmGqivZHnpz2cT3kwyAOskdR3fOrR
DlYZULl6myKInsoqwMtJVjW9MaA7llLnGosfwKuaSF8wycNYfnlYXgDu7ie95hJh
Q6h1sPNSzU96F4lqQTZRZDE18Hhkv0NGn/EKnLCK8UmWjJtE5qPTM1myEXwAdU0L
M4m79wK8E1J1/FSGnDMnr31+JBr6+fMuKarBP5jLhd5UAcgQcbxNjwQsPtC8DJbl
BhZDsTzuLvX5Yv+x7SS/avTSaTxFZ806noAiFiQQQyLtyY6+UQgUi8PgX15xwR14
HGu5WBt18eXSvKDm6CdE1mvvAh3HSMV3b/T+Hty7lyGFiiHkW2pvw1awIWTOH4lu
/Hxld8RX0u/CZ8W9J8OS9SeLjs00BXid9sw4FS/FeJU294R2lr3+uoGGvLcDl/9Y
a+D5sriCojnbhBnIOga3mbbLgJMRRLlybyaWxD3+5W7aT9361eyPcp+tN51L0wfh
2p5T7m+dmyG4EChlqT/ED4yDJtsCfwPpwGGtg//cB+pVRwZQQcm3W52SHnweAQv3
k/48UcqG4eixalnga+bEkM1xVyItwdoKsiYSi+4Qpimx0tR204hBF/miW1rDhjfe
Rg6fXXRCeFA57K6XLrRqwYAdGTZG4U8YukksUsjCPPbLY2NgCwBuEVH3vtyGMwr1
ntmTpAc2G2v4lnmnLIlHsmyA2dZfPbfl8i1D2JEJpe/S4MYy+lWGvP+QCAPTKORF
+yqoLwQ4bX0AQbKCHijtfrlYfhFLugvowfGxWXtZj2w/FEmkI0hsO89vJ40yylgY
HXsO1kIfCK8p4qBnnO9sOksUgiGpGDdsLVNvgzNLBoM+zoitA6s14UpUQQ5TAAaY
o1bB4EAbadEYLqrZfKKQneIJf5CyqWRYMctuENPfZ3tDrMKB79ydF85epBSn5Z7U
AHK2CrQGhlZU5SQd87FkZFhoAceymn//PZpGzjhcDVApDkuKabeoCDMU742pccDc
X8N3q+LZ5UNnxoZ5txVBSBBK6Zw2ntsk/dA5FMRnYdaeNacEd8TG0OuwTDgocLXT
N51dMRU/N9Vz3fT43qRzh7SWJhnqOECHL3b1krlWRrequBGvHCYaQqNFfkAp1wMn
gIbXGa493PNaTjULBM59zjuKBNT3rb5l5+H0oSQSXITp3uBJpPafVdk0tWgE8F4f
TnO5y8U688zJZML2uKXjTZ2aUKAtJXE4mH7vw9stnTP09x+glnGWZBhlbOrY42Qi
DWxqakjWx7hGRO8ENlV3gFzbizzZB1aH3Ssf3Lw/6+Zm+nYZjaQLkIB1hVth8rD7
7cmJVccTIfUGN6Mg3m5C9vGkOFbk3okQp7oIShwnODLY3ZqIayvcJRem7Sh0WinA
UZMFBrKW46bERBJXM3P40PvHQblNHjuhi6+qWExFdYVIB2yyyv8f5MdxkcBPba3C
G7JOL5+SuWqQw7q7jDDxyzRZLLp9pDbnh7pA/RYG6dQktOxGzRnjUbOdgU/JDdml
HB66BSZYyvsds0qWMDjgPdsPiNuzE8FzcpVM/XcT7PGLf/A2sk21usiXHvCKBl3B
D4jCtU7avDfpCAgRWDl3HfcBUJe90/BY5/nPca6QgkZDIzMzSXmbAR5e7S/2xbOk
SWg4w5fPnUcXf2WVqVrNTV/V0m/oW+uVAdGBF1xlWw5Zxcd220obuu6sDTL5yIpx
3a+AeECTpkGtruLgB48riIX/UOPzwXrrQdIoPQu/5zQ0iI99rX01l4KOfCD0r5Et
wCEbKYqccBHYmxV7MSME+iw5s3VotDry9QkjNOpxmXI5r+VkY8vfQ8AeYF9oW/4R
ztXKTr7IhzrB+LUTK04zwVR6rg/EsNvCOLFcpvfg7tq539SNrCbEofl4nhjBNDYU
k0C6RtXck1/baEXKp/zk4cF4Gm5pUPcd+kQeyvA+Eims4B0jjsAb9y6wtaSLvryA
rmZSpAxdCdWi4IP6FdWZViKmVTmZP+54G+dRnrnZFN3G3sOjIoMbJ8XLe1Gny8kf
2hQYx8jWLzhEtqFNcaftEQ1lzKWSiSMaD6XvFpH3DOTCj3/TjoJe/DRQt3agUjcU
nG83Sfi9DYTWMdbaEhh+/u3wiQ38yBU8219pzrxwbapUnRTAcpjT/nd8rG7hSw3G
V0FFpOmE6uKxKG/0zVloh4u56V4e6FpkLitT+33NxIh1yFYD+QvUeONm6BUvbggU
8bdZTgYGatgc6LQ0ee27CNwHQcrjBepaQHqYRPeYONHjEEh7dUv8+cWb4g1FcZ/v
4XC12usEZm7cV5HczmVeUulTVV+CYxy2fP+uhuKzHXzkxIWWSAPp6alK3JGU4k4w
4CGI/FevyEB+X3sqkwixHik6tLMpwKxAGn4HeggwkxcQxXSzqEIfcncvC94x158F
1wOvlPHeGTCbTCVplKxkX9nin2xSmucg9O6G9ktLoUzi6Os/EZTRYqba9Or5jeze
3IXhGkcvOKpOCFK1SpDu35Gtx2B/LFATq62QsLv/5U4ExRirvIStif213wf529B0
avWkuZm7X1UX+wmWVBZFH++JaIs84e+S0gDABzDdtefcSdgi9vg1Hg13H4NaELW4
O/DIg7GGsu6MC6d/a5/UL7bNq+YRV6/1hYChmFu89t4OHhAPbxnT1H96lFo9uEj9
LlR3ZqWx7PgqH11NVRemu4uwXq3fie2FlqzWadlGiF/jO84vTk/h764WqOoSO7x3
YK8Efyzq0ymqMo4uhaMvhTx2v0+M9X4D7/I4e8Ys+aU81bWy7LemQaOngrYMEMEW
RmecWPbTQJRYd6bvmbjf/FkTUpeXzh5ktFXucBR3ziyk5ky6WAPInIf2udKQoxLR
6vT/tnLwjC0gl44sSN5oydjanZGNojyG7WMEOKCSQF4T3828UCPIomhgLhf8BXOk
Hqx0w//aOszkqCkcPYodNzgvOfcVBQXVdKwpitCPt1Gkkbi60d5FM7WDMgezqA7T
hceoUNs/cJ4e0roih4Ln6fuSUsxdQTCIMgOsrIpPomUDkTHNC1+DgbNxiAr7UWFL
TuucFC9twJgFBKn5tG8bQFHoh3if/s5tWmtz/SN+wfPc1nQKCznA3CXOLhm2gPvc
qhZEpOIJ8mG35hHvmka/iR9Dm1xzQwFV4wEGUcMP4lS06HHLXOm6NdkKk9SC1+6o
rXGH4QCtWjCBAa0jUD2nb3XZEs2q9AgXJkDH7R/zhd882xT8v5ADwy1wiPjunqX8
GUyO1HPzsiheltloU1cXa5a3Vg4cFGggs5yxgho9PqhywTycSdL2QmnXXrA9Tuwe
MbR/sGYyNLYuMmdjf8ZF8rIe9BrCiAdmgXoj8pnw+w6LXAffnTFVVZzW4TKicdQm
+aMRtlncn403YGo6JXY3CCMdNfDPSX6BTPodToNZWhyd86Jorm5x6GSsGWMWmhQj
gT3nxBYMkgj0CVTJjSBYtlU2Bjs67etHHANKiq1I2hU5au3Q6KSuE46BuNrfzINn
jA6gT/APuLwJdjBKyw75mwq3+yBFADchSctF4AUIWDYiQ0T0iqp41NP5cnzbwDoq
XLyh3DXEZN59MKhx73/A8imV7B4ZT/xm5ljJmKzjegc1wUiD79CSWBlsnbxgeizV
fPM0SUYGfc7Yq4ipmXnQGjKXQHhUdgXN+tq2rLmMZkJAB0WkJgOjUmFJuhHN3q8E
MReitsTjWKtLMSDG8z0He4XJvSQ1lZZftcfvQP8uyHKmNszsNg0C5Gvpctw4gR2U
F33TdMCZFT7ke6BlQd6UFicoaHCththhDUiGl7cJwOj8JWFaLc5k/n68XpjMMLUe
6VR7XUoeyaoY6/YHhljuM5tf3jp+2Ov3sKUfWcgN6scPbhKZMYXf47NlRiQNpol4
EVCCOkHIAhf9Vry6dbJIE5IHZnawnf/3V6uGcs9jtxPm1bibmEFeYUwwF04UeS+w
rxy8wL+0TPx9z7/TsuuMkETFuroRlw5teX+vdHzoa04cByI4RiNhGI/GCOKJAnYo
q6JGSwoqqhcuQMtYr5QPGovnjBl5JvuskXif+rMEkyiK6o+S8EGCLT38gWcR4JPy
/Z+ohVbiJ5a0tgr1wBzNBmUGX2x8qKRUjL7ymnWo/RCn20ZmcYbsKacc13ffP1np
0RmINOy9ESe1dEWiV14Ge+uJYmN1KW+clFnbZ8oZieFcucgGXY0BPe038zGjAxyX
HMMF5+o49MJnc9eGorFIhMH/54Mtc5fIZOtl/r1EJJPp3YiJVl1emb9sd2L6e9Jy
xOpATgAvTPPjXk3zHFceybNiVcZnCiLPP2NIa5/JzvUV8VZZjwTClTl4Ctfsl0iN
H3hgvS9E3Wg+pm0zKiu43UNnnQho81mbsAhnNUN+8OXromat2THSl7bKNsJ2d+iq
IbkxXEOClHlcv9pAv5rozlj6qo2y5jhrmQRmmZPVK2a6+fLIe5YK3J/OBLJrKGrd
Jw3SbkHRykptauICbCrktAsmFF/RpFUnlkhkGwehtGSxobFmfk2KX9T97i+C+wnY
qXV1Zdwv2AZYU99teiUdtIHhyPwVNKmXndu12AHZUtu4BStMTqJvCA+xauY2dPUH
1dRQmH98gkay7L34ItEu2V5+NSfYEFb8/F8UCvsAj4WYiUHMjGefCuCC93Nw08G0
ATzbWhipVWgXZPUR63bMiLcyRF5bm9+1Rt9dm4ifmBgg+kaasW1pMucI/PyuVDy6
R1ib6WkhHu0AO8Vk/tZL+3TnAW0dM8f9CGbF02VZeTj+JEmHtCKSMnCTJG+vIvkl
Yf5nS16QNHfkwV9c38ZMtqtPqo0WisxotKX5Ckd7lxYArZAJ9RfneGnBnNqXO+/X
3hiiE68V9y2rlDCacCkJtjwT24ca4woEGeU0sNaKZSkrBqLbW+rPjRyk+Eii6a7t
/OPfYPSnSlCyMDG2U5rz8F75IiULU/UrkrWOuqCilXk1ec9kO588Ipj3bY5txzg+
nEIFIUacunlFzTk/pLIpvazFGe0fplw21ca7YLsj/7uSaSMCY/s+/uNFrNYT4imP
ps+Cua7CoJYzrjRtpGqtCyKsFxy1CLISdmrHyVnKrdxH5jGpa6M1Jfv1nYUxAkWV
qyCemO5vEsQ0CqVFj+uIELX5y5kGiQRReBlaiYJriyUlAa6TKMGUOoh6I/RwHNtu
q3Vt+P/iA+nQfedlLn0soKzDTL/IUc1Fr3pSo7lZrFXa1y0kHC4XAMTEesIiMLFc
BzD6nRIBgRocdm1bZdnS8sz+KEdIlxp/YcX9rJau2547Pwk+vQ5Ker+E19Duzf09
d2CAU/Oh6KA0Ou9OhXMFTpzwJ3FYZDkvd4Dfh0tsUWpyT8nuiF1R94V+zSrJ5xCR
/1OPeeHP2IpPWMq45Ih7y1CxvsPpvxRlDq1Iy4anh+bOY6loKC0uqse18b9EceOG
upUGg3CmXreacXjda+b0B8g+OmJ8g3SbF/X8spInA/hoZ5NqfyNccAW7YgPejcUW
GIZRUXgZ/cprqFFrPzuaWLAunlWsAm7tKAhfUjxTFHvZM+5TYviP5qarfPcd7Ivs
zhksSCllee3Qu+njKkf+LdBOF+eIw6i61Vf1xMuyUt3Id3B/F7hfSRQ1jrDYG40e
KoXGPKSrBKaYJFlC2oA3D7s7Dr8SuP8SkW/dWzUav5gumUkcbTeH3ooSn4z8XM/w
AdWGXRutHi1KTwkwzivkB2dHoJzCwR3UuDN1PaNT2Mvom2YsB0ZTRpTG7VK8HHNo
DL3eB63L6mqWMHDml31eloU1uISvrG4cei1SU8vAruRVrjWMXzIEamVVi8aV9f2/
TKbZqyVPjoOI+2HEVApjRBsemzC+r+OSfr/LKsoKSwds6nXDsdwkEZBudOY/cv4o
R+BAXCABPzvgLI1IcgbLxndbHQ/b2gVg8T4SYS/2+r+utRtRDRHHBcz8e3ENWGCo
C4cqoFZ5mHXC2bR75mfJh4lLk9MkdTXBBP1P6+8BO5O0isw70FkaiSR6dZ/D4l5J
7wVV03qjxIk/VIl1AKZ2l0h2WMss7EziyyJd3seImkW3pg2v8sPwWEQXqEqWr/gN
x/Af8BShpNUsGE7onBYGM8Gdb1ViY2nYcfuJN41PXpagLPYfoyIg0E6qax5XT0WO
1k8eA7WXOZshZ4oiwqWp63ppSz8/RjJ1pvZGPmx0sb9MrQ1udJfn+TWiYMVot6qT
7IVYAD9LAIFl4t8CS0pGaoMZnjFP4l9hqI7kfHHECIlaxtHVQNYT7TKbKaJTrR8L
nEgry5cy1ENGQ4h5s3hYOs54IyDyKIRNWL67X+SH7FymOBErMyi0FcxMKII0pHYo
lhps2An1Q2VyNIEY++CbkJEo5eDEGf6PHW+n05B7APh2RIvNtMw1tDbj7NTBQm7U
7MZnuo8wXACsgndDNFg5obeVT6jCForH1Kx5JwguEo/vtFtSsom5pSpNtb+5LJ1w
pvWMhdmDOjusevFOjo0RtPZxrXbpRrCYulRhV+ljgTzX5aqEs0Ebq2uyBk8R/mbM
BsdTTosVFnaD2Aa/K6XUC8VvJ48mIOKJ34L0k6f2nUruRGH7ZvX6qDHRWZqry11u
IV7Ery6Tan6eYYQi3vqIc7lDI7Cb4VKYcJXZRZxi1DloVX8KQrEJeT/Sg6pzELR+
Acc/DT+TrplhqFGgN0aU+6ZRKvqOSga7remTGcFYIhjIHRRbXbjYMsyW1+ZUahhb
r0LlnlEOCTNz/Epmwrbrsa/3YQYUc9NJXe6X28ben7HCGMdkt3wQNz3LHJegzBqU
wUPS5OKe5Nah+PClWYkxdH7C3p6+6DyPv3R+4LjsTeNIJ3/IPhBASMBD/HGyzn+T
FJT9/UZA8AM0UqBt365B8unY+ibKDHFCPcNWfw7ebvL7BD3EBWtxOnba44jBJA2x
MdybewiosSZ6bXwO1pdUIIdmFyiEWXNF/L8g/XIPji0vXoS6tv1+7qiOhlX+BIgI
S8qnOt681x9wrg22HjcSGraoI3dOB/4KWVAJ5ICiiC//hDP8m1yfc/WI4TF8XjOM
OaGgfpR0faEW7Zbu4sjl5tR0eNa9gTOblNT5GxQJre/ixVZIzr1HrpNaDAtZhuF6
xM5ufwk33j0lnyTAQuSU4X3KtmJuhUy9K6bu81AVqIEYyXFyvLej4HUxSoFxhTSF
gLY9KyyfIoO5JQsBNW4Cj6whKy4rBriYqqz5go/tGxXwn/3WdeodQQCgEokVj74X
N9HasA4iDrq7S8d5X7APJtH8xpPxxj3QmumS+ucKTwDgBQ56vBBOFALPV10d90mX
D5P6mOvbVTfgVywGyFuiNuX3F5S56iZVO7yPH6OztLt2zmZSDI4t3/wCoiNPnIio
5Q298Rf2C1nJHBr5GtrTxFKrQbgrL3nKNRcMPNxMqomAQZ1Lhx9tQGlUgcCBt97F
Fa69CiTNvWNc66Vjvi3XMwg2BEfIPH0U3wkhzHdjVT1o+97kB5mOg+ZTKo362Qtg
1pNn4BbhoRSQfUGCKzFcFaMZmKZs/FzAHDtJLXlT1pGkKj5lBdA6Hq1vjzS1lVHY
qkR7V0CFtI9lLVsjh/NghqkTDaUBjgShoFgYFng68qXhocT2HB51bEWDx4oCq/LK
x3Qz3Ug+WspK6XLDo+i16vZvBnNFlIsZ+q+EisNJChj7GT2XGfBKQoNyytyPZJrO
yt67gKZuv/VgrqcvOzMEpSH5h+WcZQNBYQLHy3TZBhuunX4OMJHdbiYfDVYhNOdQ
TnxyIte6a+0hVIH2rizR4oZVzTxcAi/T3uZPykiNvjHq0+Is5YFLT7T4aoOJgi5l
IXb00rUWpNe1lzOdfgfGPm0gHyoQISAtLYr2b9Z6HrsQOliZlYTOvZIP8qIxtLVc
l4j8OScBvYRX1hMtIYC8MlvmF2qiG6JOlnpqU/Gb+47Rx1eF0p8Ax4Y0n9mx1f2I
/2/eIkWLe8Kh5JKmnk4oAWfiTP50mFTojiDZEzwPCyH1B5YglyWbVEr52RFEhKEt
aHT8DC3vnm8XdDv0aOUwxzhA92JDPIMMDmPhE7Mbr9khH5sXcWx2eoVUBK2zs9EX
WGKiQ6h5yXMZfskSY7JTlegWV1x2ATx/KARSX4SdZuBvII6Of0lh0UXCenY48cCk
9vULEwwOuDRf2Iz6/c8aMjTsCvkhAdJoRb5URND56kEFhCKowBfJ0ClTk2mSRfD4
BwLAR3C3P6t60btINXqDKX86/VQbM5CJHB3YIMXuv7455C8cCV/7RYif7l87mLLj
N7KwKZeAoTwXOCjUEU1IkR7Tq9UuuabuMnyVSfWQSkt9boONMgFhCf6QRPuTUTAo
3oBoVx9UhM7ScohOnlDw0L7SYVWmR5puqXIkX9psGyzWFIv+Auywoo+vadLC2Y3r
5FOOmtHSSHN2fVQwvSZJfDltNZJQKWFy2/zR4COx8r/zlYTCXaR95Vx2gbq+d9C1
/MweOTKVK5oElZfPsVFmTQcA1vFKX4tFzMmfRcXPRwhwW7vlrYB3t9+jjZu4OHfz
UKHzI1zPlX4SLlmAQdWBLI34sr9GTCOzDlR/ITXz0dYWXuNEalvemBmxGqNcE0iP
FaK6pUASS1ntEjWAgGoAAjo+6+ywV1F9ge2kiYwyFMUxtb+pWjWxraYpufwWdlUw
cmNo5c5JnNDLLtSPxrlK9zpwGO0P/3Zg4TTQJu+wOnUeLkH0gtnncXhd8G6uWwOa
DHX3XM8u2dcjL6X+0GN+TZqumPlLPA6Wvyv3ORGGNkREThY9fTPPN/yQQOODsYxB
mX9aCOw4T1BWjhGgt6UfDlOr97y+7Etc+3OvBJ8ZjOq6c0f3eJmrRgtkcoAGI9YX
4EC2XfcO+eWQIfHsHPNaHS7CANFinlanW9GPTnJ0uXWioUoTMBBEHfuqiCedwnd5
xld2HQWrDMTChG9gnSezCZJHBm3M9YnTk9x2MbikVk3YiUuEChwiLiKL+U02Z73t
rXvmgnUiYER+OUyOWl/tBN3BaEW2TIGdP1MFwWtB+5S5ekDpR2cFaWCrU4QqRCfy
jZKhaMnUf5k4XXuHqPAxQWFFS7kkdfMNk4P6ODINsl4x+XSgBDNy+8rt+stO6ouN
B8UO9LXvTYYIm0VRvnkcq96A3ruMY5NwrEsgXglMES6x5OLfk4HUKMfyQLaOGiZf
JN7usDCLK1iiUcGIcSyWus5HtnpfA1yRL+wEOGwRdYGWL9K9yAtXtpYNSkNRIt54
SmukehLfbrkX8yJl1SPpzL2fd6ZpLhP1La26H+DvhyxV1B6k45VSyKGDwur98iul
mJdwV2Gu5+uyau8OOEE5CDMl+0MVd7AcaabwgYNCBJQDVjvgog3YN/fU/5kcXL00
I+dhvzrnFEjmaoYj9KGbeEJwDpdv4YySHlN6hpvgYOlbRNthG4mJCJsEF0YuyEYZ
+3s5CNNRbTrRjZYa7VG0cNMPtSX63CPSmajGh6q4PcfBlMtD9CU6GKUR8r8HyHJ4
L8/yZV/hp0eyyCmNqbN1kAtxoQQrMX6KuzKptIffNDrtqSv5T7GerkMs92fip1Ja
bJiB15rIbKrVWLnyxa3/rBEQ8aIm5tauFmhsgXy3MKY5/yjy7Gvt4BoZc9f+O8ME
rq5LeD5J3euo8B38jeLAgYu8Y+QeKUMgW/ZqY5iRTouSXgXOG4G7o4NWZeeVHUKh
g4fjUQ+pydzSfq4AmxBl4HF6CH3QHbgunxPP2b8oJ8555yk/+Wz8xk+W3hPydM0I
LXyujWXxlIDSrANYUj9WhtnvgKUJB9pbtzUaeu6R5pxhBnVHjV5CLfaI7suhk9WK
U3d3hRlU82rfVWfiVWn5FW6YSsE48q9D0jT6iqf4gC+dtFtZOSKKRFmvhQDrByZc
wxc8dYUvI3tGnVyxKEV7UCa0/bCAH49nvJtnAgRf4mdUf9Wd/Ad7v4S88OBHQAtC
2qlv/wfsIrXSkS1aiUvcPB1fR8AzEwcVOmpZmIad5DT9tfdUFAWmo9gJX068wKa1
tTeKKe4JDCX9d8y3ym722V+eEOUe2aHGAgxqJBgsGhPGNm6U2/CFPCcc/p7yPyAg
azBA7TnNHWEvUEakV2sTSxo28IpRtrgsiRpyLsgftmZplhTtOe2KYxMY79JnK/NX
L7aw8t8EV7GJ8Kvb2cYqSEhsA0ecU7WjrvOB21nbaMy0PLZD8yP/RB+rDQQuKObj
zwYJv1QHq03s6uCHyQ/23MJqX8MTclXcjuQYag7mTw6+/o8CSykbUpjZF3k7ZvHz
Ygp2o37iRpEou0RgCEdoGymX8TapIcqvtTWqgaYQ2aMsFIiFxr4evpi214biQ+Lv
G9FFYGx5efWhyaLsKW1Tmou2Ysu3DWDGmVyuU2K9WwEtvT/odCVIiA+w9Yuv+iRO
LMfHkJJsduefGMWxeEItNWfhMR4JS2VxxCPb75L/4L/Frpp134uB+ItHhKE5aFL7
rspegKIQuUfZAhvU9bv8JCGgoAfALL72nHpNcQpte81x2zhc694C9SPJmfPR36A5
+r7vYchniDwuRsp3atP2w1EtZXd5u1DfHWPTf1+kUx6AHq/ElAFnJa2kJ1tXvBCC
CxPw3P9VXkY7ME9nO3No+KCXS/4HjkZAYktY+tByrzkqEe9VX8YXfhXsGBDWEmo1
yAtUEMdfdV+Fmg7exAkPL6ivobVE9JLHnx79mP7WYb6mpb6fhbrMEQiNMqJzBEAh
N7Sl4racEqqQEwM/8seJS02xKGuKanAUmxmQnD6N3YVv8a1swRL1rKViYoz5TkzB
kl++yCzF7H/dWyu3Pk4gUZO8ulVFostfnEP/aWpqqx8gBKordgNGs42YYvfkRrIF
+TnWSA2ytjlp76tpwnHGuzeJh765qSIoM3zi+qaVveJwt1CulJXeehhoA65NOBXb
ha2w04IkqV85afFFJSDnk9/dTT4HAtBtz5KJ6DJ2dV4tVOfGnwGzvEq1gqPk0pWH
ZWwnSgamIcs1q0p6SzSecf3BvMC8iC1NgoQ2RuBw1HwLl2Wv965bUIpLO7XAbjHJ
B/7aJd+IAEBKb6PPKhVNCrwe3REBHwVNHhn4k8bglTJjLIMZGLgziw+t4Omoucrr
xBgTafALjx+vZCvi8pwVGpOeY8ogsyO5JaurKII1myO14Zs9EPd3XWr66N5L/KWl
6FtUlOtUl1Teif6aqroKcmWGu0k1yHv+K+uJD707lCgEFy5wCZLjo/cNafeLDz11
5oIgkeVjbtBjpdnnjMTmptyHyQa381HSZqG4opuobLoR6Yrv6nPpDsGvemcsEUfT
+5N9/X4CwjvGfeLn2WZNBPbc5WIN/pLhgPARrpYfamKcfa3m01gkKZbOscKolzfK
YlVWlva+1QMIXTOV0sx/Ton0EeKM0Ju7kx3qy+V35sucXqCQ5pJIVuqvpUnSF0ia
opC5vIfX/lGgf+8B+e35/twfzog9s6QFNkt13Js5ryIVEGAp7UD0NvAop3UA5LRN
BPc+YNQklUFXcWQ0KY1eJAcMShxyb5uJOLVwTzDnl0ke8nKXFfCYu1UWPzT+1F9b
2LVcX2ukkbty4bzi74aSiqujUeVCYbRAH2MknMkHc5P/YAMGT6xUucbUSTeczv2p
evPS2MVEFoTwh6gRMA4Sal8a0j8SyFwQCrKFKhxUZKZaJ5u2Qc58oJQe5nGr+SVH
n3/jz0bIWTHCEDXo8EHuK54V1df8jZGhoxO38pzGQRZwWJ3M52Ymu4bPPMz26dTY
Z2ossNc7Jk/TkY5P0JXTGMlki2ByGOlBRMgwCTfbfzyvulwj9ugVw7XsxALPZCDU
90J8EsL44JgKvueBmgh8v9lNqkDd63EblXXXsqPoQEuSvgYCOTItcNQS5IChtyUA
GC5eYJZFrFqFCTWwG9QPewhscIIzaEN7CI1HnffcV5Sdp/mYo2b6s4rLTr+bW3yH
REhRsW6D5dNXroztsTev8IwkUR2ysAwlOufk6JD+Z1FkU6laweb1LumGxkk7/uOh
UWqfYM7tWExL7lyxYAPUF2AUUR/kf0jWe/YRrvdW3FgeeBtaCaWt1Ev7dwcAJNf1
5yLpkie9lMqUGQRbqtMPROB20KpLqjtKyntBfz2OzQ56eOK/mgoULok/9qVvGUpy
+4bCdC6q5NUSx9+cREAcgtElZVbb90VZuEtwzfdttno9tnRkwtQQe9XTFcNCnRkx
qBHV0rrc/IAJSqbwkMuOJcBvVczQfZWOVHuXI9CKspJDL3ojh6VE9YS/1x6jDA6U
jjXSMpj4XpSmmyk/Z36P5G8v1T+dVBoIGye/JDgJEE+TeQMACTEBP6/VINtamryT
a3pbYj4nSVtHnz0A1O9Emz+Q2JmVN406eJq/5unDWkMmWdCyewYOBR23htOgajov
g4BCxxJfd5xZdYB0QUKc4G8Xg09SeBSiuxBnf02aj+6raiwUveTkqHZJtBdRrTad
SxauMa1zOVIkOAfKNyOur2oQUeEz6YbFtPPhnu6EE/Nb3wctMFqCGYmc19Az0EUM
hoW8frBv7xVrIdDJNzMdp60mezq6n+vpOdb0+iDQ8R+j1f2D2408YqZtxBHimWEt
LqXgR+pdb98/xg6c8jjdh/ICnfayUCbt3q86V9yvuE9GWSMTM7OGYL/eDKOZwXv3
h8YX1WoYTcSJPRLyZwRzrHydP+eKvZ0JvWlb8ubLrEJSpwqn90vZxgyXp3CR3diQ
nVrUliyCXus34rNbfLX1I4zJKXe0usCjER+HJ8Da5wZTzDTUzlMlDeselZKBNZub
wkBIndoUfHgxnQ9wyDQe2U2SkYvGgxaOwRVsj5c6LqQkk+zu365bpTU4nP5WUhrN
rDd87WLo91S2fMyR9TsgELP89yaEHAT1peQ24MD/99qn4SlZVaS2Ut/XNyJsM926
imZ6Ec3UqB3ODNyIopmkL62s4J1qaIQBiETdZndEA6OA9rQVsadM84XU7AvR0+F6
f9ssfWJsBH0qsjAiHY5DRaYpYjV1qNLU7v1nrbWzc1a7epZMOUzcOqWiI9B0vKiG
bumWT38fV7yUVw606ANriaPOgKQX7wGiOZbXQEdMpzeiFEpP8dcMxfifID0dP2f0
Z/wRnlB/Vkew9UBzT3OoxXWvSiaG7nQb7zbfIDGFTYFprvxvfZ8otNAeVGkH9tPw
akmJ7xSnKUXO55L7XIl+yDz+p4BoDANwTfCg4I8WBuaNKi/cXcMlNEnk24wnpMBb
q+1Wy+Nv8PBxZdTVCA8LnVxCG+cgLUTVoQiAIEX65Q3/pyMoFJF+E7lgvAgPdge1
x1Fw7YKQq5AenpG9WZQp1CSWl+QE3Vh2r4fco0Q0E8QIQC6ytMdFIlWXHa7T9VGQ
IPw5Z/2F9bFQno3i/79Fa7vXV2mf0vlRh9lVE/W6nR4rRBWJYAsi+TiC/4OWtk7q
Wgw2SWL2IXMWcbbwDq3IWh/AE+w6ulfLgUWuG6jRCkfNidEqH0Bdvsttdfp03fnD
AcHQDNjZN7ezOuFn3t+2UJP2Bk8WjPYkjTrmvTxD9lbuw4By7ANbPzkMi3BwcDrA
5VXwQ4l7kegtaSh6fjGRvs2JQAT+XZA620iXWQWGty4MupwVi9QSN8yAo39Y5kam
qMILpkbH80tj0VqE5kqDePZFEp5vevhIaCfNvdZqwHPFWZQ/JiGECG4dMyWss9Th
uqoiZMKlcJH/dDL4drZDd+92pr+GqZHD7r0PCQFNsWvqGs4YGyEr5vJS/RmZpuJg
fQo+5i092n7K0DoSkKXrylEiBiyP45/62rm39/FZm5lFw8Eoayz8FGhJ0Mw8Yc8O
faPy262j2LGG+EYP8ZAr4DGEOCfkHEe1tc/VSh/hdXn1UnDDKZpyLodlXYmXt9J9
ovhQW8QBy028oVgqip+N2d+7qC8blZiVUEzu7oSBmalII8rA/tcytqPm4B+8l1CN
kTWSFJiSWmI8iZJjUzDUrVlsnCTerVZCgNzpcthS7789cQDpKVBwVRY4gUdLCncb
MCQIiRSEp5VDgloTiJPsMFgzXmCRzH7FQgI5yIIsEXejTz/UxSxa4p1JI/zxU2o1
nBnMvY1/8znqnQOtCljBbclaZl3GJx6MLIsvvoA5wCtSQuwyZVUoLx6VOI8VK5Kv
iR9qiQ7IDmKS8REo5I0BLRYHnGYoar3lbwL5aRXeNDaifeBHdJkA7Yulk8U3pZVe
4TsRRtxdY5mR/PRdMWEbAUhwXXWDQ9QiUgS2SBTc7WVRSTWgxN5j+t0t+apdagM3
MJhVdI5O2dB87fOwJxitBu4RAeBxk54VwSUIq/yeLayMa5O4PVJn1m/sUPaofOFj
ME8AWnm/gVLNKB84TXYUN5RRn9Glq/iBP1eYDE8Y82FyWiVpLeVCkhGE8zKDIR+A
mXZA7ozfo9wONS/48weIvg+MsZQ3U3TVydZfvjXpKDiLYbbDyl3QEQfdy+M64tNs
b0l/se3FhY3WMVST0/IS2MgOImym71+7IJArmNKw+IldbTXv2oPY1AJJGfem0dSp
2wZ6LMQJLwgRX3s0TOah9b0UMlUVUA9FCEkBk91di8/pH0tHnHmHUl5ZAGIZxD0B
EW5qquiZHAqJVCU0HpiC7IeQC2fvPCqHl4CO1AGMDd6sm8BBVEgPh1olC/SZg+CW
YxkSqsyfjWRc5x3vrkZpKu2De51seft+aIOEJgVypXwLVI6i731pjmhA4AYotFO6
DlRH7sKyvG2IeCKpkvJSCYsrUITRhGoq/a8T+ItrQtcOy0Ngg2yIxs55JbsVqqRc
k/F1WqEclj0vjehNinI73wp+WC/aeP1r8+ybnSla+ZqOpLufLH8vPWvrNfueiArM
GXmXVF6+SFu/b9rnc9Pg/wuQmU3nYP4EStFHylQse77SEIdMbdyglyI6GkcOXtFE
xXdJS4JDoL4R8HmSgbw3o+AJwTRP3Lllifq2mrmVatDVw4Rtdx8p4GnaDvi8j0p6
vExu598HOe//OC7/+g1qmuCFswotU9YriMJsI4Qb+b3R1I4riKUHeDjmbBtoSKtP
XnCurKcmmNG7N40blRSETCy5aVeaKDw0f9JVBLgHXPVhvKa237v9PxV/NZAkXzvy
igBB5PyjUtI40mStwfTQPvXln4mQAaAGpFWZQptyMUYGH0xVjXwJI4F03UO6t91G
WkU/ebS6HWzfjXGldSv/wWdVptROvkvAZwpOYpKeRWMNKngzzaVlzIXaQQfiaigd
+D7MPduQaZUmjTl3pbhOdUTmfKTWokE4HbU9PCbw/qxzA0TvTy1F8PsxFyvVEJZI
6m/A+mK/ocij1viUkJ+w0VZxmPpZrs7lymmKbPr7nxDpWFJ3/FHLTa+EYEXTxGhS
T3fo2FqSHEdOpy5QXF0R8pOdSd8OontNnjs+q0bRlyXxp34eneTyMj8fVKuqrmmr
dSw0OUDqfBqrBOdLTA43TwsFfVQyTgprAH0ZJExtgW4MrLFaHJ5GsU8H1yRNbgPl
njM0dW03AHW1mRRxIesZ/8sr227AM+SFRQNNBXF9md0XV+Xt9BYZJfCU4uFrB3Kr
+9QcKGMpKX2O+HjAI0cI5Z/MnkyKc2kK5E5Eux7Qjt4gd8JqMrgAY9s9KVj+J/e2
JsIDJiWt5glGbwIaAgFdnWq/bQEpovcPnfKOcIRzLvNGgElRPiiGI/9MU2GwEy0g
0CL6vt/tmNgsJgjaKuHtIJ2ZiyyD+Lf54KgbZBXZKwUJTHygxWkx9Fxv7GTdt0JE
aZE7KujIzjxiczlFvBJqrqeUbk4FguJR3LiXeLB4asuX2hzQTrKs/BWawBSp8dH0
nllvFDEn51IIJacrTvcWO4LSCuhwfbOskprP9ahU6vquvsGAtQkB1Nv3/0twjakY
2gJGKx4lbcJSp9aHebK2S2LMaFu3cYM/ROIKyF51QWZNxbrEmLgijGZUeiDvbDN+
9TF9h7WyoyhezkDeAOGwI28kXXZGQKBay4raP+rLQpNML+v34+94N5WmCBUulB/2
76/15myl3jOkUpsDGlZtUjJM9lA3n0SIbFEcVHngCsOiNhD70qrDqMThf6nfBRKr
wumhp70MJDwj4s6KS5Vm8v67FwGTsdrliF8mRtUks4TOYF0XgTPfAnt9A1G3FRid
JR/bwUP1KhyqZ355pULoyyqWyRd8YRGR76HBOaqPa2BHRKi5DmjbPpV/dOB3AZbg
lEwqcF9eXmcIhDrFFE8WZYzY1OpfKwl4LUoK1erj/zs8qxaFYo5VonLvOGkywZK4
niAKFm/1epZpDzy7nJxYqogVF5XSzGi34Fip1kH6ogdAmx3S9es+F9tX+xWAk+DR
BHyPwuq9DYVLTE5rhsJ4yohl5zxscdLC+0g0EHiYlK+Zpk1V9mX6JRIBdVna+ebq
Ho5xDJ944nP4E/aYdxdP4I7URqnyACIRcfvkGw9AKprJhYB9aDaFIdQ8u6fFw7yq
d59cAlSNnXO9LwNqygrHpvexQni6M4oeds9mN3bLjfVsdWuOuNMqypDgrmwCLsma
t9hs1eYDlawMqBrwKrxXNlZjVtUg6MBgxuZDoSMBBNK+xIFeWFYuAjK4jFJ/bwRr
8+UbFrI0eJWQMvitmvKBMJnJQDSwDP9vO/HNjzjw7RD9G56pUx7dLjOgzWPQhhoP
sjM0KYuu6iMIbH7V72Uu2jyeSvMCxq8BiRk+T9h8TC0HYjHRa5rpPd2rCgmz/Urw
21afOQQnUUGRmSsJqcdrS9nbFKD8i7gZSQtBvTKsGytcT6b8Kb4PnRxPioAQgS3t
Wg1hCbdnOQl1ts0b/25K2hgVNAmnKJOin8KF1Wb62FHcIBJu73tHAEefwgfE3Lmr
a7b/krfg4sc3ceCIcEVvnpGObTtPqgSW0r9UMnwp0F4Zdmh2Wfd5wFFsbfJhDYKE
CItVwr8BS8AEFln8nGyIzPmJkn68khqsOgZksL+OOhhDqv2rml0Bo8IUyxIxMWHZ
IH0Lr4OH3G7TeL9Sv5yWAOHpREXC62Vx4NX686ZQzs6JeYgfN4mMoTmdw/dNMkvY
z74EJra4k/jGLg8jzsOZvEz3xULFXnjsQj1tYbsHWok+tXYCGLHymk0ebmYtIk4i
9rCDW0QNDHsst26MZJnAgFFGtKMjxx7TONRT+hsgF7Eq7eSTTCyOAqwM5v1dUQOK
GaYGcvYD/ku4pfs0m80FVv/mBowhW6XW2Aid2+E/uxNbi+3ZEezYPtoQOrVclIML
b+6B+d+9jt4WR+yoHpclDTTzYZeL/VsZgz6K2DyPmzl2tD6ZkhrPcoy/8HouRVj2
BeJtAE8brIaeB8ezuFsO0cc7LqHQzPhEc00dJsFERIq0CDN8VT3WJK6SIJXD6GLP
7EImJNAcevocFmtt9R07YibpkxlgoLz5zFAbOscFvisQlD9z0ROlEeQB9wJId303
XmhQeqBnmOy+4Mw+sKcsNO2pzRkh47+s7qrR3ra38d7Nvdg42nEbprmtx41FklY9
bKSQ4OSkkLZ4HYY8kLJCx/Mb8QD954WKPRfrEMS02+dufIilxdYnJ1acOSCGX85q
HCUbrnj8AKS2gvVEPm3kGD+HSRB0aEOcX04yxtNvI8D+zhwC/6uF2ZAHjwfNtdoB
/Wa8Cb9r97RW4R8YDRSgKZROCuMAcu32HQHhD5Q0PjT5BCpcHf7qI0UxHxdthLTt
aaUX/jpxignt20LEyML7dvQOEnmfq79Chc1g2akt11OYfL+zIB5LMh8UZfH6z5K2
lvcG1cLp+mQUPBO5BskkKRS1Jz4nQL02Afxt3DRCMxpamwt4RqIra52MbAPV7a2G
gWD+g/1korDzAejDBTCDcn7ur4kWZyAcO3tgKV/M7Urnic7xOkqPgifkHEDAjkKd
b+b9ne3RGx5dti4iqTamXAjUeUPjozRpi+0lu9GcxZhlGTmlq56enXd/nzA9DhEZ
q+UA6k+FNvEh8Ix/sXYnLP2Dk+kY608u27VB11oToQsI3wSJksId3xQqtkRZ/K/s
N4HEpmvx1q/GCGVBbu97mNNupL89/0vARb7pvI2jwCQKiEAW5PNEAezZHY2qjxMc
OyACaEChxpdnH8efHT9xZE9F03zzhbyEEl7bJu2JiNlSAsi/dPMUJZalvtKNuyNc
bIJTuK8XhIvLXLgn9EE3XIyhufXIIlsXmhTJLT7vL4nf1FsONkkoRZbo2BRqhasw
+nq5vZ6BDDx5zl7fSTnKQejGTLSXY+9YUyfZt7JrdosFBKypaeVmdDjQD4BVNFx7
gLvgXPl5tZnP6nzon01UEyJ9d7VyuVnlkDTRMNZoCfYCw5NZKfxTwHHmjWA766Xf
ZriSlB0qyx3JfBSAusNcRNbdeGWvFSJsVWCTx7qt9mKji5ro3b40AX47exZFj5Cf
PFw5SOj+tRGxbpbLcylNrn2kHm9HQa/CriXMdZmh8pQtVo2tejXUIvSnczbW+jzg
Qys2SJcL/EAmGpvqLTKbBm+4uB6y7Hw+vncytkhqMC8p1T5FupENIsj/b/FXA8mi
dUv5gOELdb7Chchwp/ijJLrvONa7IxIPlFOw//rXcf18nwyDQkYZ8ei4TRgOtsEO
Vyo66TpejNp6siMfI3lGh85B5pBqqWnyV8vxUyt+OzvpxkE0VbkQPUZknwcnZA07
Sh0VQ1KjOEtvBsE6uhwTNhJ43vIWBxA3EFqMyuCkyCAttTaSK3TJVn/UMnk1NbdG
Ksy5sPusApJszSf5EhiVa3O8b6hDE74DMlSfpsqiovjkN4A1f1M9LIH6rYzZZDJt
l8UHo/17G5m1SKRxzbkupN4SGuGsmqZ4yiNsBm/h5pVJLIIBHV/9SwG/gBCMP1cB
YPT8wAdkIX2yateH3rlIaCZJlqNXqTGrE5/M4fkRD9hZHSOOhfkKxlNJMNUh0XP4
ZK3pLzY6hfn0VdI5OXG5w7MCzWpsl8/O31wITnY/N01T/wJLD4eBfBWTfNZx/KUu
eu4xIF075C4TyVlpMdIBB6w2OLPqsv6MAMpmbrkS9Tz09ueXCGJ3XAlJcC3unCX6
aEV+jxb1pBMpxjQS8MUa33mIPvz/XHZcWrNW2CKR13GS6CqP1dTFv57Lao4k/zMA
rVJ5AUR4GUJrG0QgDkdm4vuFnJ3zdAoJ3x7WQCMpGghPmkkEvQNY3iGJ0jy7ESju
j4/Wr/oThqSALdIz87sW/aHnkVm4ofOSwkq23OSrarIwqbWULeyQGVA12Fjd5EwZ
qx+91LhSw1ajQYbP5yT9p1WRVTISFWwl6PANYme0MVz+YW3HIMkAvD/2MGSiHo8S
1CyLjg3FVRmQYDTrDopdy9R++Bj4iqEY4dHFVTMc6A3R40AUyNUpH7oXSik4yzUm
tzp0QvUnKBZmJq0mHgDRV01W/EDiBs43DsrJ/wpWDe9XUPhQs3T5Zk3nXFP0D3Dn
urVwwmixZpxiAdSiH7YzES9saoA3ATjy8lptJ4a2+bMbb+BOua7JedutgOA8o+U3
buXEIxxOqM3+BpgZZ02UyvgDYOTTT+FXE6h3hKI2hCSVz9+TZLIIPB4bfAlmrIVL
w3+TfAaUeMY6/C06HHY/5Xp8Y++QcoIZLinF2br577YvNxXCbHXcIJEtuu76X9ha
s6zIqUeEWnk/Y9d1wXs8TNYryGvNrJKOjhzEd+R9HjRbuTo1lLwCciz1bsXHkO3v
5cJqzfFRDdcmfaLIWZMzB7gMthCuIucCVEqv5DiqB7RFjErDDCOE6R4naR5igrsy
jCMAXUJ0wR6GyS5sIqnDweqN3e+FevpC54Gzz7NFpm/yHi73EJSHvk8SJkWGcSuV
Tneuof6jkz01d7D1iq9MciaOLllva/5hevgXOc2NvD6nZz8zdp2p8KNY9KYwo6LV
7nX+28ntYzxsJCmd9jLGiXHSFE6BWHOBhgwVaZ6+CWMF03CQc0TZFnSo8khERj2o
ja5FBtOc7WpJmkQlftanuyB/fvL1ttq8YJ/FkVOpnz6fO4R3ymaeBM53kjYQFfn8
H7otBUr0+wlxX0heBejb+EN1DfknDTzFC0hbdH/TJxbOZQJTtyJgxat7z5xiwSfr
ideQF1FOAZU0G4qcwvwaOvq2g60bjxzW1AtXTEuJ4WJcpPOFeO3A8UgAG9KMIHhf
+VvCpIwW7UhyBUACu2f2fdb+3PbtYXEOc7simG1OCurSSWNrkwaJXcV+4lHlth0v
oJkjj2rOnKqFhOmm/vDgKpMzxZoy2JxhTd2muD+7ngBeRFTstYR4szraTLxB9zzk
ZKSgNR4bw+lF3t44gXtjtrNW2EhJvtgCuHZZPBtGp+NrtR4twA3LF094B/FMPYfe
3Wpl/7ue/iIi0VXCVA2Hupu8Iyv54DQihsMlDNtW4NplvMBjR+jdCjsKFywfqmzP
jFbp6sN2xxXlmrM72sLRq8kC/pXgYme6aZb3BskJcfiIYLtponArrOm3I9fyUVEt
XPyrPAedQ6+UV27vpMw7TMrQAa1qyia0dx9cD3y4SFevjNdCPwNZCdjF/e3oI7kF
OlY0hTKpdb+xpAL91Wq/XFYLc9/Q2ovQNKkJkkuomheYePvk9NvzkJvkpdOTRu3b
sy31RwH9xE9YzHWYcxrtjEYL3W+k3EKwtGQ1rM+7E40LGtq1O7eqT2nBAuzPdhn2
7bCefo7QJPt41xo8jcn1SwI01OKS/cs3e9NQRHXjZLcEqTPNSxNqpDXi/pNFcqJY
79JlHxLkIUMSoa9KZhl7EoVZsY0XoHQP17BbwidcT4+zJBphaLP8/rVoZyqEYcba
TU0dccMl1rGlqd/GiP3AhmOPLUADUA8SQ6VFPgl1rlW+UjxP9BYxEdKcDcdUE1CT
GoBvJs3wzX1WNWcG+ZRAL09Ur+jRve0lUBfUFbznHLS3hf+8epQgEjJRKde1etf/
k6vSzbzr6UNPk3LJOqIQntDeip2OHlJjPfrw6wrZCgg1lG2Ry9Tzo/evdCSHLKGk
KjR8/8/ICqLdK2ermdF4lDxIDPtZWygwnhqifiFohYTg/LDBixZZPvzRRl/8CvXZ
WfozZJ/TXWoztWev3PXutz6yGjATHZcaWHt250+8aTFPnCtfdpmlh5k1wI+2kt5Q
1jFPoI2NCq4Gx7UmsRahjabe/6eQh1chcKUrDuOHtGZosU5q4EqMHfvUfOFkvSP8
1V1i+ckyIN+zGzgJKlJxIkam7rQTLAZXmRDinM5N1WN7T3abGDEm+J6wgvcCKHby
K0ZhGJ0410Ie9bNkYGDa6KKVN09U+Jqbrqs/u2mvykxx7sul2trvk6J+BIuTQ4xZ
EQbVIk/NoEMoAjZh1MJDTW7UZNPPt+DpJJYmgcZjB7PnVBqftRiienPA262VITah
Jj04ZrPik1iKqGzCldaDx/5BFbPSgMHRC+4DmEaO9l3fyQjUyVD/vzOFpAz/T+bl
prgFlnPi6ChxSVyFTXteQ2OhLxrwWj4n8zECmbHFFK9Ztn7hNjbKCiU03qjogGBR
WFiz5lOu6HgoXWf11LQJC/SVoadgkU6n1H55Ieo6jFd4Bl/ZFkN1qMJz5q7wjx9l
0HPJYI4OLCLyTLi+GCvTy70c7QwLiNRHnNK4k3vIG0jRAlisknH9zVViCDO52kEQ
tZb4nDHu3+JdBwEKAn0Nbv3WwpjPDqk3Mt8pLmgS9vnTGrCZhResmgTJet89wEKx
Jd7cYYLSe3qGZsTr2Y9VpgmfZc7TahKbw7gjWQ/DyqzzJf+Llgv/hHTTbWa5qZSD
n7auD9YCEsy36eWF/QgqHODUEVLK1ev0n8zL+RSezyotlePoOpmQ4+iW5p2B3KZi
kGjAjedeYljJQAFd8PjtS9rYpnH6kmlVIgxJNv9/7LQBAJ3jpV2WH993Ohs1nqKR
Os9xhRaokBzcv/xacDeeQVAD/tuhCFFkpfI2bJXtTOexEdlX+m14qrezhvcmV23n
YVYXeH0Ka9zzW7QjfAIT4CXzbvgHgnp8ohPuYEWmtRTLdauzuVJR6zRiJoqelY+l
jDYX0vo5fu+48ZuYsR4su7Py2c+q8A+qUTKeMCR2TTRWTDb+48LlXklWdDozSMoN
YNKh8rI8FOSOcYV0JAEMaPPtCtfgvOrDEZKPwJWbWApsUa0vz5xk4m0deynlFRYo
PW97CRumZn+54xkrwTw2NCHfJBCD1v3i0GnBPNXNtMRs/sJC79DceamaTzXtonoB
2AqW1D1aKeWg8m5cplmMtPs8TTm48mP1tEdrv6+DEXTvYbAuO4QQMYQWQhT1OE4i
DJxS+nsSxEeiQsDsq2Cbe6dldfEy6Q/L/4VYgTzamr4zvNhqz5L8cfTiZatHPqHQ
mDqe1ZD2zVBAxPppRULEysTEzYWPKYv0Lh9E3Eg0MSxFv1GH/SEWN4XYp5Tf9Bza
Vt6VP/PhfmxxFgmIq+GAggoKVDo7SBNqvmTjJDHzmlKQu0k9nqWRSiSWb+XbybQl
ssQxNvrxv5W4kH6CK/lNC9gH2NE6zgJHcOuGh9nN4JDjQJ6nPrr16wAluYSKP8kJ
3DYBobRkpRW7ouYMlCjHTsl97QER+zDNIEAO7Yn9HeJNF6j3oSMoeCzjIxeTOPpp
nH0tcvW+SsgKlfQRgqGhpLqYG4CAA22omfld0LxaVFndQHCB00NzWAFA3Ac+Hmq1
8/0H7aybka4fsYgVKAjTP5uM1sIKmN0xtcUMcUJXy3tSbgZxv3cK8o/hMZgYaAoY
n/3F2DCYy5Uu4XjX0sScdJ2mRN9RdFhP25e4X7/D6fWYmivx0d4r3rnq4hL1owBj
q4BVivO8QjJz5ZFgLiOsEynWwL8IQFeI3+dV2DIJw2cZtOm0nHDJZuTtt8tUYa0s
ycWCIqojGvsABteXzgXOXcdXHpGDLXm8yb4omhFhxjl2HlGy6IZS34ad1N70gNTZ
jPsaMfqjSsXLQZZkgcGesscenDNq3Zdf0t0dj2g2iOB7yUnYOh57yebPp84kcBOU
GL/v6btTbfuE9xNcsHg4HAT2UCzIAD1Hpf2QTYBBCDqgUUFgceOK2ZHx0OZPzpQv
zajI5w9wZDVaCt2lzbiHRi6gCuBJqlzNuO+V41azvIGRseQG/m6e8Eh+5uCW+efI
SZbPBLGJakvqpcoNgwgor5Y9e1OL4M0AtWdDO5gJcSxegQFWMe6wYMneSHTwEcLx
bCuWjOvMvAj8xevEWRL3uj1+stzPLsjXU2WWYkS9XUa23NACx75+POiOptExmRFY
rNt16pBB4ebjizYTOfQwmChIZ2vMDYk9QfV+GXV8z3ewFzvp8WKzu1FOu9NxbO2a
7U/mQGyo9mkCLV4RJfBlXY4ABYXb99e3vGywpq4hjFUq8TficrlLojhIe8EpUxt7
eWOWJf1ck3H9791sPsXv4vfARyx9pxnr2k4VHS5ZKKV80iYwgWwqSNeRH4Vieqzp
tZFRPCrnJiZAc2OYaE7iQudQKGT7omncZ2rfIz31Adig6nbDVyvyD1iO8SJu4esm
Y75Grqyr/MFyZHxclCtB15fQ5l0SjJmzXap2rQHhSLAap3iijStmpYCiwofD9hBO
soVeQHsRA4MGNFTJyvKgIS6a8A5PyhIpXUKvODfZ3q7cKAWoA94xK+hC1CN+/B3Q
9bxWDEZ+2A5LcinKb4UzCmFixdVBTa6tliOXf0+yYCSjoiXQoY46H49eK5asGnmm
CJZmF+VD1nlEAgbo/JvIFthyt1wG0zZnuajNMaGtBgpdvD1AlWyL1ZwbmErLRUp2
EzLrwqgVPibuycsCM7I0kUuztdF4syRT/NlCD1E2O8jGd2BHPJSLRA1dyzgrXLh8
45VidCeWHpf2vvIIf/3/3MixuJ4VcrCuzIVYjhR2qeZxAOTUtKeMZxlvgy+Z5OsJ
ZliYUxFLBqvse+vFTnhMsOsNKyIhaBujIoB+IeDRZF5truy8fYfD+kMgbJnKlU70
SMR1WJ1VT4/NOje5zmsouPvkP6Iw/nSwXSBRNMcVTgfi0LSV0hknM7VIW8KLIPVb
Vj1r66OJP5aJz6q5UEHBr4XtvbAEi5bAjcfbjd6MFqy/CgJJf+hTSW40/TKERFqO
DkaRMibHZBL+T1OQfyfXuDOqU4QCrK+spiDgi8JjZ49TpnyohrL+63fAxIOn14BF
V1FnXN+D/iC2urZOjwnuiv5TH/QVd2VV0znXWNlFkcxltguJjaPfOogUXufAhThU
nXokjWXierhzb0fcEE7Byb3vGYC6m540TiSfKfbwOZnHCb2Bw3l7gATIfoQAJe3J
FULExRZGkTWVv3OoYOg5bnN6PyW4a4IAKLQiX/DqQEUxIXmUvoxSaDxJd7Uquhh3
ppOuofZvhilXaJAwPiVXtoQUoqkfqX0tpB8BA9EBltX60F7ojYTjtt3qdZB0eWod
hZ5ZGIdlrRLawa2NdmSzjEMMoCv/sWqjb5qgNcew5GS/5Z/zAFrLQEnJz0Wo9KrO
6rxujTUjTUnJfbtA5zyf53JlGzCU+GrppBcsuvLHDjp+kcXrLguB9UVyO4i/In/9
7bzei5TUX4kirTGLnJlxjQkRDVUMPR+OXxjzZps+IokCDNE1kMQqWS08Z0i7oqN8
QyuCuhdTaM2u8pH0mIQKSisiMcZb+hs/imEE2O6GwCpU64PAAaeImVUOsv2xgETM
gma5NbH//JesAMb1M8h7RmQBLrHN74nYaKWme47Rpair8T0FCreh9zgo+Fh9EM08
sSiQu2sKWl3Qof94pGfofPAGUMBSjan2Gqbh0CpUvClRxZshY9q4HuI41HOe5jmJ
i2ncOjgAMPk35EpCPpf+ns8Tf2tYrp5GXzk8CJRTKtDMmtfDT6ms/f/ro5CzO/PF
7SU/S5waKXD7zNGbEaceYTEhQUW61kiXcb7gMmsEsCEuAQ8jOCZYfdwZET2GhHED
GwZX2g1oxxwX2tmboRVWibyEYK0hsSchlL31R33G6ZcsOg73Vn3OiMuxtoPt9jMF
QnZGpF2MxUpcIsNdnpYQmGteVZbM7TRRpRZMUgqEhvPbzs6ZqZhESO4sgYt7z4GU
FG2nwcoLqyKX0K//bFCzpa6+CJIYHBoRBklITAnNIuiWhLozupBZfJx5zoJCQvlp
7KnLsnv2Cr2X43HJFFe/YcpYUWb+ZSmrtIp9B8r9WSCSWYc6D2UnVZYPiNSFj2zf
t9XnDOtwJquZ5xz3Ugi4Cj2xKH4qhrMU+sovKNATSURhFHW7E/hBne3WSFa2moM/
PHxkLOzk8EAaJ/kGHl7rRnpXDmpe2K6P0Wtw9kmKTDcfPhN8ZU16CQ4TD1Nb1SeN
RUrGGQy3WWxsE6vEAFSdAZMuCWFTLmbHp/Q7vjK7uE0AR/W5bxz6wFXyzXIPUdeX
81erdjGP/vUoR2LbAebiTBJtN8SC8MjAC32cxv+VqS7Bv3hurSOk/CcF6vRVMT7e
N//MGww4FOXf2sfSBCD+do9fKmu3inx8vHsDvxHbvCLaCKlKPjQbsyzuXAI7r6fO
RZdNwPtYSaz1kqBXptCuqBytwa5vKXajasVb+da/+yNSLWoHdZ0ZMlsBqxjmGk0/
JicpfizEkp+dYysmT2Oxs25wgB3mYFoeaFkl83idm+gzbaP97rhJo/yMsemWNM7D
iXYxBTHu4ABkAE4A7TpnIiN4xP6d9ZeIlrNPi8ROEXeVovKjWdhsoFJtNJZGjyI/
+I4nSJ7PY0aQi5PWMa76MBuA0EwtiBuKDJ+jgPSEPPYc1TPF5iT2Z3Gg08YbX9PZ
JFvRFdlb7HyOD4EXHNfYs+xAAu1UOx1vHC0g6IjlSI5RKda5LWFTQorA35vSQuC7
AC6Mh5iQ/l8KXKZeZOkKl/KXV5opDUTcl8n9zXvb3GoeQKcOh/XH9YrR1ReK5i/u
Pz2vObigqx6QHyDkL7C87NG/dt3kL2Pp01nKeGOgIGOREp4yi0ZvNgjBs64aZ2o4
ZQAV9I9zuxo4CGMdqVuu/qRNMLSIyFIkq8AM1JNgRLAVV5pCqegAgXdq2dfi+P7Z
HBttq9xqGzcpEHfnq4TJaJrCsq7ipKtx6MsxC5u/xPSh/GUlXs7P1xVRxi3LNu5N
rVW+jPzaiY7NG7x7ipmliaAJDHD1FDoQHCOfJb3Laet8vban8uAPyP54rZDsiZUs
bY7vFwjCFGTeblUd/nKKUdbTIcz9jVftpD/XYi+sitkmyOtDnYTXrxnIFU3rfFIS
+0YEPbOFQYYFla4+eZ++aWT8Zx+td1M5CisM181MitOgbDmb8SEZa9su4rkrss1+
zySdCLqWMWyyqMVTTm/xDTLnhC7CUgWketHScr7+3RWmd6feHlhpC4y3KEn1X19B
eNmoU5Vd/24hyTGV8piec3XlEm+StT5t+3I5gRhybZzOixHEgWyZPNe7XR0Gpbre
xEu5ICQa/YFaKqF8MF2q5iclgcb6AxK1I51XvcW+c7BQyGphmrzsldCSeU5MfZCl
dpnl+PI3A7tvM+SxUkJvvb0W292PGQ0nCm0r0OHj2tH2fHcHRlADRbixgkg8uSVj
OSc6qf6UMgRCkdJ6xrwlmRrVinfxA5Qzs7SSJip63WVkHO1RWNGH6BvksgaTAviB
f5w0S09todGkkBKpr8XwnvfqMgw7bAeD931wJnu/Bkab2jM0KYOMqSIONcyGRcao
q8u/Yh+ZqhoH5YEAFg1FuxJpCM8jpZloGTjfZ2931Efhj0QuPBleMIMiLPYkTq3W
HWhZ/BDjqxfRVqWBvV+HP6ooO8jj687fsnFpjweRZqVjEgCS2/MgT8SzmGbDjhRM
ei8smCIc8/bRSBR1UejJvVvSMQITZHCDN3/AcR+45wGSMwUQ8HwKhMhQ7Vw8Kuni
Yg1LcnbdLgSGvdkTK36olzwjvOVA4TSrsFWixyWibvBOgbIUfZDEoqGyzUjohqAs
0ikZLtRwdYxc8WnA9FmV+5hW7WMUqchoJuUpue4GJ37zJKjuF5SgPEi6yTvv2u1+
8ORbzPXvzKbXQca9yiyygyHU/vm89fkAI8sCRarK80u/zNikmIanbEBXUGb0Ansd
OAcV/xcrFeqMjrFDfjA/tvUnYWDk4TbKgRqC8yRaZBFSxRaUznAQdDJfQg0gLK8G
IHyQGTM75sgrEAkN7UcwbFgYyI2dOFlfBwrZAeL6tH41q9zyHrmlXYOTWr7FwFpD
dEaey6kjGz6jVcfqsd8lZsKTdvXFkqYpaNaNeSUvxyaGlk2FT/7dKNvDk2xLWjui
hn7pXxPMGXYo0ZyCxWI37Sr6f8f6nUN+VTW8sdSv534BmC7dAPxcA6P/zZk0cU+q
X0d4uvtweerpYcO6f64bJS48+fH24mtRYgphBQY9oLa/PU4rw3xD1UkUv+6PJe9F
8g8NfPiKk5+fSga4I7g9PSKyPFG2i4+CH915BZce4dEOOHxHcRLfAXphkMdBfyEI
mTghHtSCm9EFI922za6Z6G6BMT+06MVQ6K/xq+sGpTWVWDRYZGBWM4FOSwsQKbxZ
ZEZ98sMJmJZm9I+AzTJH3+dVRZuc15FIpqB+k3wmmrE7IfqjWOUoY5bXTzjk0RxK
cOxCaouEuSk3liK4cQnx0cJMRXaOLuNPW5y+Zq4xvWWmMyQ/nBWyELrSfzGGn+kD
x1fQQde9VELmM0D4uoXMP30W2PyWAodJKLZpJgt7tcNyBOsd/Qg1WqaMJmeU8ES4
bwEtNxVv6rtiWMFvIr0bLvEp0AG8UjpN/jljUnh31bikOLo4069EaIDEVwK+5fFs
kQm0vdqEppBabWduQjKXMNNRe3TO9nnfqmQm4oj3ouuC7SLy3kyUm3MhYnC8RuTC
j4QrGIMhBPtBrtCKEC86P34GLdFd/gEb2j4UVfWS/3jjx3GWqSFERygSGHlHUNEr
kPNMdwQ8BP01N0/VY4KpJMoAkVcPAqnTTcvddyno1H7jnhhXFxZ1nm6P3GzZXV8t
ZzOK4kkse/QZ1K2mxxq89e/LBwDmwdkxSiEudvmAW6/+MqvL6Ef8+c76tnfM1HcU
6wCYngabzYuaYOq1/3y0stdKwmQv4+jf4uUrwkEAN6SPeSWsodgAhNdNB7ROAII5
VTzzchMoQs6agmkxvcXY6/iRCLG2hm0Jg6sl9/t+7fKnE4nNnmjG2HxFsyjjcPs4
Bj+yUWdJs168+S4VbgQfwmS0Lz8GBRs0xuaYeuK2WjPPbmNML05H7lBNqOjuzrM8
+U22rpBOHu4SfEMC5wVHk41ZHDEJZQF6AcgGkZuIRElD9rKH6jgagY0QTx0zemSU
fAl9HHzrbNsFVETK8Q55pHpYoLjqcKhqzZgPcMWkH/Jh1nNolGRpkvLg+lWUaXQ1
dmki4QLCUFnXkPEGTjWyrBs2vDVj3Ib+8IdjfOQ4dh4SQsAe19zJkiispscGq+xk
HY6v8kwa0NyMo2odomSXs/QTg/1RSwq9go+Wz+8+d6dzVlq9mWmQu81ieyxksjl9
/oBsiBX+DxbiqHDyKBYska6zXSsOjdl027LypOiPEkZaNb4mKdpN226VqQywSUY+
zbo/5Nn/IOZh1BX1QLLTMKMoWk84c30QsQu0U5AN4QLIdqWcrUfFuX6jmxihL6he
R7Jpn5RU8aRyn0h4SwMhEH8iHCjW5Z0Cjbn/cQyd3xAKV6hqHr1wzVc+wxDhrd6n
XQ1j1TXw4CcquXPfyPcxoLadobiM34JgrG8Oqsydn+hG+z5ywHxD2PA4rIr3mvlh
3ivBuQUM0/orZ9hDTRwD+WzuWorUDafpmbhoENV+SIf/W/zyQhbRqnPQle62y0cV
e7t2E6LZNG1jhwkInoR4NQKkMCKO4Pyy6JdzD97zWMCQ4RShQsauWbp68rdRedHG
xJoLXmrXXarxMgKxx5q7eRYVXzqSwqa2tuR5R5shrrJX5B1CusDLopXnptVOPN6i
KuooOffKV8NJHN1y4hEG6iT8GiiTjQo1JDWTmHKzLIS3JofoQfkiqlZfsx216egj
k3S7B40VyY40uAeTCQ7iSAUYEnSiclsiSvBEcZJOURLION4G6oz96lIRI54dwyse
HkkdeCFZxDMpSTvX8sOhKPV8POEam9VkO3G2Uj2nLhZLCTGGtwO9jrWTAcpE7ZNo
i6HB680KKJcEsjNoIEjlE6MvH9c6iIM16xzGN5lDwHXOENCR7AE9NWEpt9z9roN6
xQbv8nHVovc65lg472sjjHBkBg07znDJYtTnvTau1EGCzkBuQxbCnK+HnF8tout2
kc5tflSmr4pVnUBpdqZChylREm8qHq3Ol+gbBoEucc6s4kQZMSaQZS1zCw84JeP6
hUOCzKwAazedv4Y2ANf8/fSLGp3gIhJsoFLSZ5rflTvxVk6BfE5ed9a587zRn7aY
uyF/yGdo8vgc4JFzF0L/N3ZBd1Dbez/zzB4BwDzqmtG1r6yW1Z8saEKJ3Aow355p
sZ+I9J23YztRfWq0+zJ9bZLQ+syWaIvO+GpeK4YRE+JP8LiQ7gNcBcMtG41n9Zxa
hXbcay62PhGXJSRjXBAAqmeIFM4Tjz6wAQ9K9mush22CtINu4tudup+Y+sCmnX6X
tfB52Gfyd31N0DgdbQkyyW2iJ+4Fv01z9AtGuyXom6fipgkg0kpPlWwYGWKzAJhk
1pd8gZ3yIaz92hQPU7mynvfVDpe4/N/MN11UsXEpsD2yxe/NsIa+i4ed7v1GZf/n
vT2gGdyDKxehocbIoBw/ICDh8alFcZQaSxIXf2oK1SxvD8c2ppgSj4EfX0c+rJB2
3HO8oVN2irSRaTFjFhF6AhPAyVC2XKzFxyZb02JPN1JFBfZaVnnSYmMSxeObjoeI
Er9Vjl4/c0MTPWWUAM9GKenFGcAFaWB00zVFLSAusyD8v0X+JJyfpzlKGD+7nxTh
mBsx/44rV6kZvefeCA4KzqB/xWLwRqlaN+jf8DxTk/ACYXzF1WWEKoSpHamnVr7O
GDAzDcKopSOrAar7cwstV/SLYDA++2aJarHrkZMGVtzLimFxmtTLaIycvjB5bVXR
wZ1JQ5nty47tbb0Yghzc4g+M2Hkr57CFITiVvDHiHTnAS+8GScEplU9xWw8J/v+7
ujVrx2XB+NTUMiogi2+S5Yrq+lkmBmlViu2rbGD89/yJsCb/DWDfI3qsL7/GI6yY
zKlmScZMJ3shfDEXzkZfc1pctZQa2i0/NZ/OjaZtWllCFnm9vdvoEZEb9POPb1xK
RGyYVa2V+13omWKVwYf9+DP2VLRR3Uw+JxPge0GbK8NBk5sM1xuLxa/H8nRFYuJK
j4gcMR/oLRilsHzXamT7nIzeVD6ONLBX/y/t0msg0A2lpbgGva/xm8n503NVXHSh
CcltwCp7JRWYUfjYoeHRtPj/lDReMBe5wgpXQwGGpdbV6Q9lH2/BkvSYe+agwTap
px1ElD+sj9xHgGAH4O7zEyrhQt8GFJ4FUYhOSvQsV43NtSim2mbFlglsnKSC+XxL
b8oqP+fc82J9WsiSyY00KXdBIKex2stM3Abimd6wUvVL/vLWDWAyri4m45rmVeqV
c81QWcxEJRBwc5uAM5oGYE+UlFX5h4/gHqHkdxf8fs7xIBuDpMdjcKZfOK3OnyVT
iutNHIPKSv1TVrJRf5QutaWuX3HNUNh/MMp706BepmVUnceeY7oCsJYRYHAZ0fM+
y45CDztX0gubu7RhArtYD32xDNiY8+mSGrnx2KwLkGXjEqOYagmifAsxcUgObZms
Edl4o/CZp4kZqyky4gEbSYN82Zk6CGgDMyQNIP/rQdw6mPUcEvG91GY5seIi7X4p
atsM6UOTmQrh4lqixbfDVzPxMxv7XwUF6iJEVgRuoYEbLe7JCVELsPTujxMf+Ijm
ZPZNfUp6wWdz2sUcmIS0Bi0Qo3IZ8/RJAzpL8mMNT5++Z6EgoKbiAjPB5Izxsarf
8HXXpIpVMutbQGU16pu1sFLQOjM7BpImqN+l28o29FLFwf5BxMhecFom7X+7jyKT
4fhQdHGDvC2tTWGOw2C4AKpzCEC2pmfUUj7U+fn0M7/tINxgxBAhI7Lbkc1r/7sx
MmB347Zd9zrf54n/ZfSZsJiFrG+z9hKDi2WHS2K1tDSyKaqupku2bwYv0Gq7SJ7x
rXPc0qQpuZajTYVX5cz72KxM9hy3v7opZTC+HF+1bO4IwZlNewonUzwRFo6QExZ7
d6hXzMaMxQNuMGowlQJH529EVHtjlfvyNASnVTZuo2yrc1zL0yU+yF0rb1nko+Fn
TocahGFYcA6aYr6PLgI9nzQuCbGZEnS8IQanWW2rehk0AI+zsWunUbV7t3D+0jC4
fA+HHFBp4rf5oMj+w8CtJXlKuyJqyN5y8GnWCEp6aKeed6jh2wAB85JDsdcJdhdr
1KWgAOaH28WWJX8iX92GQZc5UgXwhF+EtDrFteGsIc8G8fE6VreIn+tQY1xnzT1E
cNoxeILMBhlHWO7ezwK7LvT9llyq/k8NBYBKPw+H1qTAqK/mTre9OHocMwv0BpyL
YzJFFVpWPhZbitd5aVdAS4g0tNYGDKs9FvB25AocxR3uV9i+Gue/5IQBtZhR53S1
ENU4enrfinI9kGIGwuwK70LR2+Y72dSrY9Da0txTbBqePlr/EtUdUA2z9YYq1rfD
rWOfyRtlXTCBy938By5fLqmjYZ6qud59p3kEIyVAbc7U7Mr4l4RgXpKqGmpm40e3
+5eBiuleg6sT/5c4d645omi3yS2mc+TmI/CV2Rf4RV7SJDRHz3H7bNV1VmP1pKlj
vcc5RiwuR8rbr9A6kyQNkmQoe2TmtXyUXNUPJClC2/wZBpscH9dXL/z7X5w+o0+f
a/31UG35oIlm6cibAXM4D/BebFLPRVN2++il7XVaJrpTsH9qECtCT2F+AIZlYkLd
wnWR87P3wcoTCiWawWDft35We1PEMr/9Jgs/C20nZjZtECwdSrHIz84/fiLYXzNr
U4nevrFKTKM5zRRsM449CrvHFhUoHhjek8J8U/SRzyqDL/7AWNnKPUDFMhYi5kn/
/4QBLwwBGm7YPzV9Cy7W+mZTKXJTO/hBtt9ePwr34ZQf1fIHlfuJG23K372VGLVZ
wiOaoY9hJnAFdSQ9P6Ncrr2oZel/mso7VGG+WmZqvmIjVx1uIx/86x1Ki/QKNYXI
Ugw0rO/dUL7bi1o83u9zzu9ndd899Ekj2Uo1LYs16Bm3XAo6Jl2gc0QdiskEQxoE
96CO9ZTpvGfDroH53X3Cd4hsw2RhDpzc5JH1W7GeSCfMan7Q2ZUsWMlES6pvc5S9
V+Eq7i4TxMjKBKghbflicfKor0YxiMUTPj9nsqm+uC/ddpSL6UtmCIMLHECGftq1
J4Jq3i3giN7uJQm0gHFUX3tnoqknSN1+AwO8RgeIcwK2EA/hfUZ7TmxozeEHhJdx
6WkKKJrG+7dq1J/dgtChF8uge7Qo3D6SFmFpShSxJfB903n4FuWl1+1lYJgzU684
1ea1cn37Q0W2Eva2gBXjsL6WQXHpkQDvE8S0B/LfBBhYf5fuYUl/CaIwuw4p6yqc
uffq1sSkxWZ6P8H7wYaIDILR6rXGiTA0rybcYaWjjqILAYKQbvTRDoRhwgJqxubQ
KAgqHiuQ3higugxNQGyyhAj5ez7J0dyrTa9n6ly7z6SOmQBwvkB1uTDW62GErd4/
ZS+Udeazr52t9HvqzyeF2SlW16NAKdSPqJHlG6WMUZnEy2/49Da5DOHlSh3GyfFM
WGgGhzUOBBIekxVoaDomTZQl76+uYfQc3I/YghW1Ss6/0GBHVLJm16qR8VhI0f3j
RW5Pdzwud4Ii+sNUhVwbENCiTs78/i/8S+JH9xFQsxDvYJEF6HSjny61lFqm8cAL
GPNoAt28aFvG80SW1tLbjkWfV+Gj7Dr04uJSkm+D7w6wMX2ADi7f9UiMzqO+WpLU
nF+jJr/XEB2ckuiQBzZjLdgMDdmXWwTEzXU2jd+TzSitypVZr6EOZ1PmbP0PJ/pp
yxP2p09qTIFYgaa66TrhHX3ff1q95GDLukzGnzc3jqi2Q6MV9gO+9U4MAojuh1gq
x2K4LCnE2YcAUnJ7qw2N+icb1YUlC2OqSd96h+Ril7Jk1F/hVUenh+MXPK67G3ki
dDHXd8F2Ey8Vc5EdzhqFCxxOUyvSd+788iopGjjCm2+NPVU3lVKASNUDEljGWL3R
YyBpmoqyjZcgsiGaatCQ6wqbFOgyL8wxiO2TyjwmInu/0FMdvHeOsO10NbcTXt/Z
lqb/+v/VYf4/K7ZpxfqF34glB0Jmc3XafJk78u5iR0yzvqZraPxxc1hVfTqEaV/N
G7HCkbA08FtRvWyekIxAvSJcO7pKus+zoIEyPJnev+IpMZ5/17jKawYlDKgSi0Y5
bAdZRmqX17a/e8JhVCPm3sYQVU2nuSqsDqzns0K5bp/upQHEyeDjoqfK+8f+CRYN
wWHMSJGZHw525hUx3uu65uOCvO+P+0tEzYdtiO0CTc1R0QNrX8ywkk/wqn7jn4TZ
blKS/AQra0zG37FXiwuKrA15GC1KsGtK8/rhGM1ncSxtS+dSFDQopKbDgdQ86skY
925DhjKQ79TbZwMiVwk8x6xemHM4AJ4afDoEFNyGzC3mKXzA9zeyKlFMhgqK0TD0
KFAGSotUZtdYRwKxxt0XmiixbauDFWCihOtOlARu9F3dhe23rjdBtvf5BlTV1Rkf
aCpa2IhroJUdxJSHkJvWvemuTuw1WOlqSkN9LjBCMmv7lxFfKF+9dwJda5zj1Nqe
FKy8pzGCQhE0wzFofr5WQ4yX3lhG//zd+jaNoHkeOrdHNsRVO3rk2+t4v2Yzl5aC
QjAPskVTPDMcb96SbJcMV3IRRVf0HJpZuMq1fmjszcJKsz0+hBaz7sO+mF23QTFw
YCId2wJ9zXyO02ZcxOHXBL6CQcnuueYugFZPNydAEiUzc6wt6oFka0YS6QTJOWjr
8yecnHdJw01NkPB9xWBjX1QWdEPPhZStTYsiB5Xlci/oBmHtCw3AbXqI+aN3LR3R
Kq4LZcEmfRlHV1IywZNmr9I+ol+hASPWThimqehVRE8xUKu5qAOC09OipbhQNSbH
k/M+47CwLrk8tMG4St2E1W+uIO/XJV7jc3dSn3SA7MGVT1+uDMqLsdbTb4TpTjev
9ySICxSMP+aBsDeLdZrEpsG9s1uM4uniOgqwMN7IfRaqm9tSSiLG3hp9JLtksZ/H
mxWpOibeWLafSLwn8/ipDV6MY3FlcCGzs8H7vxLX5qi7olqGvaSkk2SYGQSUZHca
3LwksbTmCKrYWruUI4LpVK1K169zaIuXApxcXR16Yobxqa6bfBkL6sLsekdxsdKR
wiEpD8sK/fI3zXYNTYv7kSW4yFPGwyD66j8/E1E67H1v9agcHPP9YlR3N7yjLPMI
gtkgEUSx836wQbob9xbjBVsrqwjw0hdYO5HHlPqZVRoy4gWrpfr+BudzVn/bJTUh
EdzMXGAvHHGXT/EuiK8G98/BPFWmVQuR5X9drT5aMR9FGzPfAp8F0KkhQESnxqAH
A9yL4sfSfDc6BeghcYSXBuc1zSKExLyev0cxPSW5RuyIjBVX5niHpQ0k8iztGVMU
JGk+ZIU+obd9xOh/jDuLXz97aePQRXUmW/tU8Y7BdgcDf5d8gvBQDgVSBBittZxe
SgP7Ame0U+H++OUDTU28uwDFG5RY3Zn6OYGbVcqZX6jhg46mZPlNGvNMjQdeE7W4
OmIa9SlE3uEbU/+GIMAr3vKeSRtp3ARrf+2Kwy1GYFxC7oQhUyeLYYXuFAdn+ayw
LSk6ktiDoM28D2LTRosD1CYnn18+M8tOFWNtZ2JPfNlKARsuvyXRZkdo9knEfAU/
BQbxz5P/lIMre9pcpsI7eKp1aEQHADNWdzdcnzp9P82od9MfTe8hIyEts/jkckJS
o3cxjsp1py2vgtadlDtwCh2eahkajbQ/jqD37bZdUxKu/8p9ZzHuqF8AmDJnL58r
iPrx+TObGwq1NUgf1Bhz/RDfuS+qlZEIWqkcLW69Jp2s5nl6g3OW43CvTP2LeYed
AWkVOu2rFecUA6ILoDjPMUfi5UZA++/RMOJJxGrfFz7QfcVkxTV746OgPLQGp197
v3nNoI/ZY49OD2uP85fJBi8pf3I77bftjme/x9M/i7DCXNMcAI5NTNEx5A1gKcIP
UAxwiW4HLog/OWtri5AiLuqcVX+t1utjo93/hbeiQ5uOIN69WVttRCu5gOIARXN7
KgqM8q36GhtQEcToIepeAvHC1DxvHg93vA7PcQcCCTFr89q9aCCZw9VhGk1vdPFv
kYUKxbjTO94Zr3TYuDlxsGR+dqaPYpW/B0picFiMewYE1q6mapaUL8o2nAk/4Xwn
iZVbq+xBDV0rpKI2UKJqaw22nZV4d1HJO7gdx5FqnH1mSI9Hb+9BQ0ZZi3vR1zCl
vgpHqWKyl2c672CxMtqoX6eAkuiM4xJTT8K43QnC/tFulvwmxxpv7WoD2w1CxdqY
gAXyyQbSULSiVi9seXZo94PgeZEulzJu0uGO830ULQLgakVWaRS1rFLzDNHM2F/C
CqquBnE0t8DhgshMW1vUm6+Mv40iBUjCmykWhxcX5nR8aYaygwOTvAzD5RzGm+xH
ixI9W04dsz9KUIWZsWrBvhoe4W8L5iLVggcKssZccRAl1XSp6C8m5aIvbAqpHmCe
4tSVZ3/ED7KKGG9/YuwX8ChHcwkF4t4i1pQNSjPBMRRXqHSyhT5dtg9LCj4ylaD+
lpi6yrUok+p8sWrtyc5OLOwL4Yh7pCU1zxqmIOGpt1x1Brv1dRWG/x6Rx/nCqpI9
pM7GkbYHUb1VkTgpvVWchyHTrXkTejJFhZ+jcY1YutzysvEAWP8uYI9eXad/7C1n
U7XA2TAysJtN5Qhq3zS8NfzvbhqBuSC+8PcjzTxPmIUF9EVC7BRI0drfwFJSFHTJ
V5Ahwh5fQMITjJ4cc5flPFaEB67cmzn7x5AMdtNJFG0CeuqD+TW20nfHEoQmMxBZ
nJ/VzjnNPKhAWfQ6BsJ5xlZPJCk3Y8SjK0QldN1nRw8sI4IID7Eg/w4/5ZPfz91y
bp9Q4L/STLBCwtYtWqsGRrUcMMtTI8qPXHGdUCx/VzT2tr9GGrz8LEOqfnCTzx68
fT6iHyjZvZLMJbAePvmXYItGrEslDcMavL+EsCrK3BYwSIwkjHkpdseCvL/qKYNq
6pp8qFRhFnxVvQUsyvjNUrdszR1tgkXXKM7eUKFs6TPlkOq1Ch6yBOmChXbaT6gq
y6yx5MWYXoUWDWA/ienq2ErqxH4xfRHG1FyOI6s+igrQ3B2jXXEFQnPAEFfiDt8b
AlRcfF0QigyM3Pi2CoznYPB4OZGRp4sTsDseQvwwpKC1nhdpP1sXmtcQ6K3Px2HR
hEx/MYKD6b8CTMcT1fSoI0qPUmA0nnFvsSs2/V7bI5iP6BMpGwTsGJDpB5/niU76
Mfhm5TPqi593eRQ8OWluayr33/QA82/gHMVyk/Ea9Xjbidpg+f/EZVKZP+lYp2XO
cn75kXOiPZMxiH+InbiQzI90d8bUTWemqByH+UVVgV4ziJ+vHuSMxT3X3hExFr5j
CNLsQq9QVRxSSkwkP2z9pU0Kt2GVyWmT+dfl7+2yqbT6qcFzMA70Qxk28CWjKIrB
cvNqwPx9zm/uxofKuPu4KbDsKpwD68/PsN8InPNwVJrtef60xt1+O5bs7XqqR3BS
or9+2B694PE4HvwsnhbXcY+4Nm4gu2zqKer8lkAn7L9Vn0LFRPo4/1WGpraYQljv
dy7j4g9GsDQVGMBaanOS/mBmqZJIWgA7vg0hJ38PDxLGKzDuJ/ugeF0zHcyim97V
qBEJ+cDI+I+MqQtNkAaPf4bZNPlMw/eEg4szp2fuebUP8CcRE1Y10AiFUJeTlOLd
miDKPAhte1zqAqnAZmnTfPZ9ABWseDuiZGgOdU0HKavO1GZyrU8HCec/37GMLRzQ
YfqWwvQTz4NT2DzhhYdwDLrhGJ/BXm9eZefZwujW45i4kF9QJMEkASIyJIf0IEKo
HO1/ioo767rGA3vhpc4Vz1NcI4aR4UyPKT3daANEx3IPrtMr3R5cJ/PwUXnAIci8
EXe0fm5FUHptp5tbfyVPGjqePavOG9JcH4htMuZtQ1q5+Gn+FmmsM4Cp+xDYHOQr
XvNY7+P8m66jP8m9NnRygIF7ACRkDmQZOF6Fm0/uZD0jsmE8QRHUk74n+8cztwlJ
VztvgcolrKNXeqZBbD56zaYieYxcIbMQN9cM5ZDyO0Fo1X+kOF50AISZ4gveEuYS
cQsxg8t7d7ySdIcorVPmAsM/eVj8rgFzH4xyPxTcQhON2Zlm+7Lk5HiIU77AZJE2
mkfS9HwuleOwYka4mYaJiKkTSFeWlVtMv5g/GQAni2nv1NQ+yQSvRBAn8CNgeac1
i0VP61gAgIuAOkJrXDjtJ/Fh7evopEccpqHcg4cj/w2hY9vDoSqH4x3KP3mYSR+7
TKgzWPJEtu/DgEeTgcOT7gteJEfnEYDyoCSjpQbf0om6ICTjV4NLh8fNOsf4jpoU
B4ZXjjTwoLyhoefrYBk8GvXpZjYrF4feA20MjYyR5+B1M6Vo+1omFZSmm2W9Vfzw
uUPTEI7j5IMQqyG7fsOR3YIlzG9vpalO+09iPrDG708NNTZBsI9gXdT4tSMX+G5/
wtOzO1tkxN7WbUrnOh3JL4UDWIxYmNXHxpaTzq223a7FhfMRjV35+vhRRlmvROyJ
hiZAVp1MdTd/rr+JnEGp4GoDVMqvNYe1FL469qsA1hz6H0ar/mcJptkv1VW3ieLC
Elh/ZywS39XpDRF8qFxy9P7GSpf3bGLr4qCMDwmEveKM+y4nPSNEfMfXaS62p++s
ZKozNVbO7SQfULCIRe1JVId9vyygrK3SRa5tBPqfKMLgJ6PZFkWagGBmbvWDQaIO
0IX4sB94X8NwotubS8qz+ei7tPJTiL35GJxvej5p9lS9UVmyuTJj2MBC7ogLKBkN
10nYWeR81xsvumGbcDSXSVqTUIjvy65u8tkrGk1pQIyZnl2nD/j7XjZJT2st36+Z
40wPMG4MW4RQ08srUrD4jD9hNzQJiPiy7xVbO/IjeHjU/p1TOUvvKXxd3TLTHkGC
wLuXxCFlDURSxIw3X8L+IuHkV35kiwZsfuAoqhSBvvDiYtrwNeEx03l3Pr9sUJMQ
9hIAq1WpkzMs8WuEWtEi3Va8zruJe/vP3vENvPgTBCrwYhbP2SVmFeMhaOphE5em
SNZP9ktlu2dFnZWFC76c5ETdu0wyRJiq3etTVDrYc8zwYbXo33Wxn8I2PHIEkDen
fB8KJESqZMuoJusmRlSxxmQlLjxQ8zp5dMai+obpooxMykDPM+ZcegeQxBdfUSFp
wnqvuFCLGSaO7MgQXL/xZPIzp745Xlc2B4Wwuz/2fDpCjYe05CzmozrPFiaA9VJJ
0i0/3qzS8XZKDaU0tYP8NkEEZyjdwP/RVLwoQuKK7RzbiGmWWpw5eSlu6yvfVuf+
nPpoiO3n9duNxjNs+AGQ4W0Z58eczks+F20ag3mtk38FPNPbUNlAPm3Rjbtv2z6q
zPXo4PQ3+0TvMdVEQciZax948R+76L6MdOdG9+FslR5nNtkZPuPAdxYTokDB9mwa
bPxjQG5P82dm+grIROktDHMmUX3/vvjq1OVH/b6Pgv9UTn8Xw145X0M//ljLLs+R
jswA/THDESBPCHaldD0wB2OAYxlMQP/OsTnHqx6MyisS7q4dR/w4HGI7CAro6UP7
zTnUz1shX1K3476yHeJa3Mc+wnOUb48lc5yf3xBimL6mVl3TwvXBVMpegM0RBPSs
kmD+f7y0cpRdG6IaU0yrl/aAMHGUoU+a2Ahs6GNrU3CuvBiX5rKbBRuoH+ktt08S
rXSJRSVagVTDKOE9sJzhQ7bvlwF/5CzPEYCe9bwqkFuBbKGl++KqfTb2J3jCLW6a
MumY90YPTiRQvWB55V5ionrLd4/ruOqZBCmDlobD2BiSyA4qMQafah3oPOgwzhvI
goLufRM42NpfvU38rrVjQ/xXvpSWWiNzgGEKfCnV1FlEsqL/mi1gHZSlcn5KMu1X
CeMoI0uf9i8S6HQNK0c1yIdLjz2fGFZb2xMuuJsi1F4qJD5+gffCkIjU6zOeBjUY
0ViIbTuprSNAK59zfGNAgP2Rub3f40icrSBKas2rANyy6E/c4US772ZQiugqiRt8
KtYQS2bECX8ZaWjhpAu3sYgGzmO1lM5Ngeh8/fPSBP4Ym9mmr1vs+WUqTQFnYeYA
gVf4x2vtNuyRMoBTw+k++fFH2KU/notZc7Xq1lWbn1u35OSw7Sehd+7w7fdl+HfJ
6BJlMXLep0U0yO2RbAghcKXOyPukEJuDqWInShmFol6JDxyfgHSSJoW0kOKcfaXi
r38l9QBUxQu80/sAHNjiPKYCKsGH6l/NxhgfzrTp2UsgAw4HbnkM6cMl+bG9hHOC
KUj3AtHqQfAuILtJ0nSqbWfrM8I820w9LegZqg5nIWlE6i76RDAYDLA9L0IDUj6D
LJB53Whv+Jh6yur9rbk33v16Ejnyb8Yh1Ki1l6KThnL2lhl+Bkxh3yZdpn8A4aIv
gLLFRRPxO40Lq8ipPx3HZM7jb+F2ltsbek00RMNA8HX7a98/Jrh5YZ3aPEktmRcn
xcnNqQFiVN6LYIxd/MsBwoWv/Vc2+xEnyvEMeKiV2sGi/hl8EeXBZAVOBcA/Youa
8sGKa62kqBGK5eCZsil6ditZ5VAK9jT/MlGaqDKGkd6q9PGuIRpcEcH9r16k3VYe
Vt1jybNXx+N1yF+lugvBCJw7ILKBn2wVtq5jxJ2EOGdPtslQvllvlxWcXo70c3ph
F1+D8XJr3rnuGH/aXa7xjFYrnclCXVlzFxsA9oCeAsTYwJzdm61aWRU6RWN/FE2h
qpaYcVv2aioHY5vsltOGNnnJ9Guo2hcrsOpm3mqNEeqo/oieEcX0s0LawYAaFBpm
4hHFJFumRtND+frBotI3ix+RHfOtYlJxc4cYdSHqHUh20g59YNWxwtXNNlStcWAI
K2oDPXr5yXbWmq62IVbUiCaZdbD3h5baF9nPWvnbXqIsLrENxor+uykauma1dE4J
2euxgDyp+RI+RoE3MH+Wg5qVNrSLiKTWo9aBS45QcR7cAJmWnYqNW7nl76TezjSY
4NTE0+ecJtwSXK9xP1R88RIUzIHpnk2fc5rBIV1HTOu/aSUiEQPLPKg1mfy4x6mr
22qXor7TSSMBVHX9HaS8SL2qp8OcMmxGtSa7BbiEwu2wXztKf1UQfqghs0WnuxuF
0tOEEJke9i9Wz3fBQVwvy40vFQS4WRsbogLdj5h+cdWdCFaH1Kebo8K+O4kJ/fUq
11BfA1B3W6ZrDrP9sIG/AW6v+rUNnAth+aIwfgJf9jBtUm3cqgrUBVpNxHnebNQU
JXwlBpDbxwj3xL6JucznVVCDYWWFqLSA0nUtvouODEFSdKoJwPDAmUyHxLLTbKZ1
GZiZ+QacZlDdVDUv+dJKGif7AzzTh9Ayt2hkqAHsPrbSQFHqzbU6nbszBKmp+3pz
P/jmVfwwLSWOuNKGk5Y8O0jGMEmKUNzrLa9nDMCaPS2YHGFDJidJXaIs+qY73nUd
n3u2R9Kl51pGrNHDypZJubGp2+8pQAoiKzO9HTx7EaXlNbu6ovqFYJ51D+agT6Dy
iriSJidCX4g+9FtZVwSR2qtZzxudmuZfbY6e4TII81NCDqsHVFvu9EcUl2LtRH6P
6KnnMe1UDgTXyGdkZt6rxNs7hSb7U0lq/f88MRDu++ukE+ni6I/WllBFF+03dyKb
Qrfx9+JreEsCbznheJHq1gWtdUwXbi0vkMdCq6mSnbV0S+61cauMCosEgrSGb5td
cONnb6lGGQMXnOF7+GMwjeGU77buQdHMMwtTq6A8bHgyP1KMoCRPefKUSoBBYJoi
CtFuR1jx3Cwc+8UVYmtLnsMmZLiAB0ZHkLvb7cSqDySdVkI4DzpTnGDUKSyvEmAo
j1UNZk/XHoenVvX6bNCy8RPQ2fKqIz1vn18QdzqJyRqSkTDO00fGHo7/TP99eLax
iH9RZSdYh//4nVAsy1jA4IztG2HOBQXtbWIS4Xf1MB9JuhS4jq5cIRbpT8K1UT1r
HYNPGycwprRAI21ZMWQ1lu2Z4/DVDZYephOuoq5nEIZEXAxh3NCiof0yUZepHxsI
gFtLyqxYc+SskViMiX4PZ/EDMaZHQDkTR86SAc16zTHtqqSRwLTY1yHuqo1pOWQL
ryFPmts9vsmCWxg8orwNkcHzXoIj9bo4ZX9wTleV/Uyl/3XIaYz/HcN1TDv2LOuT
6sjfB60sQM87oQQVT6cgKk7ztsil0YC4FgIR4Pv8oJdDwOar3DuIZa3loHB0qoR8
lOP1VX7pv/DKbqB0tPqZo7M/4x0Fbj8SENGh1rpJlQPLwW9oGahnNk7GM2RFj4pP
DFc2yTsRHglVhxuauT8bArpQhXmCm7eib0IVoQnvq4Z4E5M+nmUXEWH/pOsywT5J
IWQfl4gh9FBDn5aD8YjrUfDf1XWcdkIug+ynZh5vq82kdltyV9TwgE4QkiaLUWYq
IlbG5vf+82Hi6R3VUpPwARimb8+U0bk+10SqhBU4iPlzezAx97wk6arh+H2VA08A
lQFXzdho3OX1P5HQ30TSJESzqFdPOXLNfrfOeXlf2pEH4rIxu1KHBKKbOuubDViP
Rns5MGGSNdhdwlod4/9sM5u6WuaKBHBFO8IAFvFg8U+IOAontIFAWRdfMoAfHX4B
+tFDhcNvQ/ubz/0wz3jNvmEy9rnthPn9vPuFK6dJL+y4IJnnJ2b722x49BF6JidT
0w/QkQ0TCsaXQewOEbM3/Wauv8S2PMy8KeToMebPa83/jfb26dBgdpyV0s+uHbH6
ptPcDJmgUlchSWg+KCNS4tVkdx1Tol+cmpIraoCJFCSYoYP/GRxYdpkuHV2cYfha
1kYtuVqngGodMCkhrGf4cGEHYouo2bv/q1GexnGORiBhoFjf4r8MdbRlhQ2qwo6Y
/j0oj1Iwml06w9NhSCXXgrYlSmOGspKc7UbPg1QwBQqaW0IMPQBZZ75qS2+nRlxX
yfiRD7WTdXELMhSMV9V2tEKlk4uUjI0KtfsgM38nr5ExZIZ5vHh08xIwdS8a8Pm8
WsLTmeExMetZbbTlrsm4ewS4msA+VoWxauR6aSj/JQ+z+HZ4b8zRwFicSJHVelPF
V3i5veA7Tn0sf1UuGK/1wQ4BjlL+PqmgV/XK/0XMfPE1W8XcrXiUTFUvaLlf+hTA
VY/u6Gnj3S2fQM5NOMknd7a1g5PnTz4FIz/EOo3GXFu3XBV7iCHo81YixuypNi18
0iild0davroh0+ekZwWnRcU0/Rq4gV0vewZxmuNJeojHwJZ9KoJzS+QEBfiVEah7
xVwjvgK/mAE/0x9PQoc8RzXnAzesF/Ms5XdB2nULz/i5RmNiR1sABcpPRGiiYxmP
qDRTzKpF+Lj8+p5crDGCMzk2Q0b/H3T90+7l1SPj8DpCj6HtDbCW/o6zESpxFhyr
0Weha/l8TMYmTvVk9wuhgiKEgN9xPzsPa+3ttAi7MQKrdiFiFxYMvOGQzCDKh97J
CJXzy6q1qylcPn0OVn2Uwaz0M9u4u9jJfQ1EKd13x/vUqTSENGeji4S4DvPup0e1
pDMupsFKIpV1tNAQ9jUQtVksBR/ICEU0EouQ2OPEeXmlrbl6hiGCfupplQHlPywW
vBK/YtgIcmchGnKW0v7SGCBxdOwKTMXUGuyLKJJrPIko5p6fvdEoh0rVuhzpY+vY
oMkBf9+si9ni+LrCb+3WIgKpVoZ6M/HqVGyu+aFv01FnwrQmquOhaBnIQb8OtvMk
LzrEwWnOM4ZC77jT3ILhySj1gIaeW36qIDjOSyOFCTkoLxBtJDxoHDJEhHQ6z2zo
nPgwIWI1dFfCwhjK1v4JhsHcC0UXNUQ44q8kEPxo2GDF4Flm7U03OXl876UD3kHq
5sxsA09x5MRAZJk5N3nGfbducjRDr0RXyN7tYE9UG9UGBWAnWeCEM3Fl9Ux77drM
YE6TZg4wq8wRuE030UFyrsDcU5oiwQds+E3GBBO35ahqMksHxdnDMND0xyEE4fqb
5r8ASB+xulNmEP21F1pwFbqMGKoUgheiF0C9utGiifN3tkaWp0pl+bsCZfN0MBwu
NO+sJIayRSfQ7W/9T/PWirv0zjI6w4qeM5m+TS/Gx6npwS5toy0uP+SOyAoeqgcg
OTK36pH/Mw6Wc1uPpJCRhNXhRqdBBBUcpcbNWK5wqIqTu6UluUUtFEP3CiSt1ZgN
EtQrf2xuSF7PF2k05HojJZPR7fcjM20kf853PzmIH4RixbTvJBq0ZqbHxR4tLsWR
96apmC4qInczgAi3mreWz3+mRY/ytZQqkgJMIcWh0lfSFcsO+sylAoXCyHuKM8Oc
viGJkhhe+PO2wUfEf0HeqoJJF/gP07hU0Ehd+up2Mh2xgvU1o/nLMy3dRriiZb8s
FHNlXrbSPZB2rcBjFnpGiHU+o5NlQ8rYXoqwwluxQveGcfq+AwgAlDhSufqbDW7w
18aQEDkz//KBWHIiVwxM0sIL0E9XQGjzzFPvDSIBPYzPBv1UwGTM2jfnO/LiBmDu
x4+QjxpQaGmaGKpmeAQsB/mJns3zUgqRg4HwRklchm2LFy2rnz4mV6TjySkqiR8i
OXM6M/Gaoc7ilEB1o+jKwNrsbmeKsbyRnoz61hG73Zk+WWhUtAYYCovU3JbkmmnL
bHPFwYEIIlEtIjvX9PH0chZFPeKzZ1Clkzaa5pf8rcFvSd4NX5DL+K5S0abhSMVg
qCpE6SJUGdMHyPqEZErA1HP6R9ihMvM1Fspy960//TqtX2JSJ2Wx75+x6ZEtTJPf
ETT9dVBuoLRwaSjyM1B5JN+3NlvOs/9FiVCfrjXbq68kZ3RGQlOtRED64PgCXuL/
HdkcozQw99rkA5rwxB34jnQUbWW7jClxNzrRzfJjQJp2sAVPohldiekwzx8CqOME
H1BeydDZmaCwDs8yFzWPQDfH7sY180EH6pph1DoTeWGLU/LHVydNM8GFaANzkQVw
JSGzaRAMeNzKbdKu1Vwo4F4ahqTUR3bp4ObGNwqFwNZYVqisBNqNbiIK5kvgYQtx
YG5St6mKduJ2RcRRQWtiqPbsGvbaJJTvZULUl02q5xK2hnjGE75miM0Qmlr5Fiwa
hWHUb7PXMYzo39UlW+szIhHzImrPD2/zgRhxxfkBIwyrro64fgat2uryTuDW3JOF
1dkKwCssN1PKOuousekUKYkIZm+NXrYxTB9Q20hwfm8B7uIAfsLyUeJ5xrUkLByZ
lsfpAIPfYojafMFrJ0Q5zCV1EYLG14cvRuUFMXWUqFRFLLdv1q4NMAMgF0+oWwVj
eN5XohSsY7KGJG0ZDRDawHn8BjeXCG7b/th5qCSL4FUORw0KXH3dhJJOobWrD9Ts
KJOKpbex5j3lRCcoLvQm8aOlXP17x+7kur2zPxPd5v0CtpEyBODuBgC/E9nFerfi
36GHUF3Tn2KXfCAHcw9prNvCweZMll2cboQrhynN3JVUvFdBjzVvkPaw1Sm1m95Z
CIgaG+YfOEalk9tlnn54NAXpZUcc4yDruUCggb3fUocqDBUpX4I8z0wLsSW4DQ4t
0d72BSH14+ct2IoZEblvPme5Q4SMcDdd/VA2Co4EuijjnyzOjh0lYXrngL1S8hS4
97y0lZRTHIfEfG6gqBVURyyWBMvTKUU4DL6W5AnkgWzjiWDN4EfzZsjaXON7peBZ
RtybuxkEL5/5gCNc8DrIrAnFthqU1gozBdEa2gxFhmbYCIDt7giykLcjmfTh74U8
OYJVLdaXzbH/Gd3SUFfFy5lbT6XQ+csQV0Gwr/+DpIZaupfyhx23PyJjeDxsRlD+
sHsLcvFEXFwwUvH8ipUiZzh0ZlIS9mPVXayDw17IAgcsvhDp5Ug+aLM1op1r+3Ih
A7+RBzyvhZD9ScMYL6eIVxgJuHRYNjjmv0NvXmDTy5KxEClFFPUpjaaYRbU7T8/+
rFQ/PpJZkFoRluWQDlIwSqHWRundTxLokbOBSmOyAbCtIEIuCd8TcgPiAn7wEYVZ
Iap8s0nP7TxLrnJnnw3LqEQaQWVJ57NmoqfPDMBfIKWSHcn7C/UcKLf4tXn5i/bc
O3HRAtjekU3OESLzy2iBinSfkpvfouxuwvKdU5+38xMo2TNYj9KM7gti18x4AARm
jOCiWCzoKf4JH0xWJswh8BaSRnBdGDXCpS9oTNyMNc4mVfycRhss1pwMYPmTNMQH
bquRDWowIhh7G7Yqn2um4D/HFQiPdCPwFMfwrOd0v1JsaO80ynNumEHXLgr5b3M6
eZcVfsWm/uXMTMn7xgGOle4V8ojEPXVGNBKBZ9FluAL5zRHJKnfJ9oeL67g/MQYM
rvqpEsbE1GRSvEU/lWEg4HWKN7HfkdKOQjjlOSW4lUX4yTeB2GF/+UOarM+tohyB
hfaaY+CxvGs5u20LpEXxNGT3c2h0XFmEOQp7ACm+V445AuYifpkkhp9zuJUwZDbi
sI4aC7LyCFCLqUMrXwCyVor0kpzHj5jUadmfigcr1RfwO88Va+UGDjUZzSawzLOa
udoHdAk2fh7xb+3yRLlMsBhjklQZh6M4MoRFHOSei49s5s199B0U/V30secI5YkU
Yl9UXS060JimFndsKv/M1y31DG7w79tptJRq3QU5BPDxOawCFQ8S/GRGxs6aKxsI
1QPFJwhiDCyhK6P1uLb81mn2cDMSbU/Xm0+LefDI2TjqdNIUk6q8WWEIZd+7sHyh
aAA3mLY7fhFTdd5nlXmNuZx5mJE5FnNMRCfZJEntPAI4J014TgOq5NeISRQHMg2T
T963LhhfphQrfThL9/m6wmDYb7b0rrqQDlRLFQBBcooEtZzN5mmn4zgb9ke4Ta1k
2NPazOI4mrl4ZFPnyhhGwUx41L1v/1oikhUL67rO1uvSvFdv9P2jsbnP+5H+SCZl
YmHucmZaNhJ1SE7WLkqOhyYxSFQkou5Ae8pNhz+k9i7F5xCeEib0YMLDXJ5vF0eN
wqs/2EeCsYBc6XRt5XdMVYavQmc3Bjao8ATYqxrhG78qjnmM/oY7OM+f4d12er8A
tcJlcszhbCT0seTaS8UpQVSN7kx+oFRbB4kJJwjuq2O956DURYOPuCtyOfA0zI4M
WANKeIxkMwNJnLfOCzn16rScE7RM5l5UEuu0vmuIcoeXnXA+vNkurqbjCpOZ3kEp
J/UFtVTeJq3wrtqheQWNSya+MseMNNAWOo7/ZbKoVZvdZtWRrXY0K5FGfiYILnwF
J/ys30c7YnoRjWm6DB3QtTd81FKJg05z3EBjjtnEbBf9hCrhN7vXrDFhlOsWZtNp
/YB7Wq1LkxxMd3nizQO6ZjtR7ZVazLnFn3yTchxBkz/fqC8Jv2iZ9R5mYqp+aRgK
MK8Ywas2dsA0aCKoUpqs8GAP3RQKvkhDnvFw92SZd/kdmGG6044MHJvLzdy0r9ZO
+CIFvLT++pXbxYOXkChpWF7JNZ/P85QmGXRrEOG7I0+MBhO+GazcDQzguWDVtT1k
9Bzz2SzJUBEH0D9IGt4g1D9YC/lZN6UOmpdp7tAuLZc4gWwAtBUJWhymrVUDQ6we
wudPYQ+oZKmYR0IWn8c/WzoJ4VEJeNhAgN2eFSbNdNA0+2tNKQqMzUqKAIBSv2ji
eSSe8ITnGn1nYttd2k7PCuMYxkrO4NsjgWKF7l7n3Aqle2SEEJM1GcRL7caqHllG
dxhSZqYQTlDnaFztGQ6qoieyfs/Re2+mqLiCK4TUA7tD7ZLuydOKu79HdR4tWP5q
0Dv3R4FmyYaoFP8h8i+EvgsWKuik4YWTKaY5ZjqdPIhDqJOgGDmoR2siZmC160BN
z0BQAHtAxDk1LONKatXD4r5FSRcTnKDHtq01eh2Nr64xMCJaWn3tPhdz5IKLYaI+
pHZiM0UdI4fwXhkhjn0OzV28rtHlDK5u/mrAdxTHp0rNjfPrE709b5ax9a+S/XxD
2sYHbkw9v4gREq9mV5akO7Md6+TtPumGMPaUYXZ1r2HDOHJ4CzaZbB9ACcF+L2zD
+1oiLT+eozKiEQx1Gyw94deaTw4a9nRD5ezlb2Wtl5BKISkypPRQBLmpzYleLHfb
88q9rCZ+Vuh8SQwtlccyEVtnyO4znTu2tQr7CyUKpWJPDbkJyb3IFHR+o37QncHy
TDC3v68Cskwzf6boZT4onzatzzOI94kl43VIWOIMeOaG6j7LRxix0s5+N5AvDVct
0KvkPuG7bBdPeEs2iXZEDq/m55uJ8jc93xUuF7L+GiJGGTtRz8nFfncAEQQgKoLh
9s9+cHCc3tC9t/ZXTeNERDaCdpzTXNQt68ufI7FAv12h4DoLLHMPN1+ztzDh+Mel
h9ocFPDebq419e/ZAj6w984Y/kpSALGhaeOGzjaZ6q/wHJ/ITDPviND4JiTFChKf
yZSBm/bx5x+M6e8Vk9bf/gX86Ai9QrsEIxemlExWqb87ZW+ezHffc2G2sgWRbyNa
HFOJShwXU65xVlYJ68iTxxUTTi5/ZQJiPffwDudhFKnqnM9IsYXFXrGDjKmBohhO
9at6aToCIQUmKS8EdiyF7YZX0gm3RN0pI0NRMXk1/QUoQfyG9XYQIpBxWYi0MquK
/WZFMcFdOIIitxY8QcekLsPgxI/mzyXqDe65chTDyuPJSmyYp7ZiJZ+HB2rG6U6q
GOrrzrFNjZnH8P/6ecii+jMzPjFDgsLAPCF8y5s660Jy1IBXgTRwodHnNty00c3a
QQqvBsLVPF4IMWdvF1yNd+44esptPyeWmgTHMrigbK5U78mX82H62Ebe1abZM/za
Jk50WareYM/1rSY0XNLeK4rZLMMG1NgpziL4H3TaDl3MaZI19HQxhSLJT+qg8QnP
+VKc+xxajuivizqGWBrCztzdujv0Lunk64jd3kX9H5N9cFWEGq4JuL7grEMv8h1d
PpvnMYVU8tVXWENU209AOkqQshz5XJHE8uhQPHUHwUpu1HlFjnJYpzrbB05avzOJ
H7cuo/dlkwEp2PRmS3d6uOZ3ktKzkiWfetLPygn03KKiUxfks/o2y1+hITWpAFKw
6mJZj2n6lfgjbGprJPV+x70KAA1esccKF21tN5Dmchjt/qSPk1bbggp7BsTjz6Me
xaPIaXI5jcTLMbAffsR4HU1Fadk12Tgb38QOL/dQwRtAsD2g+3Cm+05slUtPeqGc
k5sv3K/PPY1jU9hjcs8kTRxxR9PXes1dzM/7juySB5raR8lfNOKWhAQpA9n/e1tV
4zrusirIWZXS8lc/N+zLPFFy4e+STqHgUOugtCygldcajP8/xk3e7mOiR+s0LLce
y/bTrWkHBJ4YggLPK8W/M7U2QtwOs6CKYoxhS2430/pRq4JaagofoyB1JuA0KWEK
d6VBGgInf7p1Px1bpTh4TeXS672hxtTkRn0lIUYUnB2N9UPdLX+JXaF1hq6nmTJg
i7uBvHq58u0PvUHp2DuPOE8sbQ4dzaX74VE38s9A0AtczLh2oykR2/GYd5bMcugd
ImTPtgUd3EPmk0ReyeroG17R/OZ0XhMniNEGMSJEWUy72j5iEdBvVWASH8j4dMHj
I5zXxAAOGsiq9zDaIt9hBsYaZep4/Rvo8A064jclV0UG2Q0hfCCeUllpUqj74C+H
6c9veOdMCyFMNCskWsRjdtNFR+HyBmLR/mOLV3dFvrvck3GxnpwYEjav6i2aWxkR
qDJjZHTb3y7zK2MovaWuA2ZHCOmNAFteqmfqxIbqGVC5LANQWR/Ls9pdsVFgiw0I
ehAbGuBN/pkQAAgvwBQwkGmX1HKK9tXTRnPmeI5RX7pdfYK5iAeD2Zgk3IZtnWAu
xMOYqrOxURn2lsSmb9GCgQlPmmmWYExAXS+Pskf9QxZm/kOq0X26/gPVC00mGFBv
IZVbTscuylStPQAseBzGDbPZZan6EfiDCs7/PbhCiEPOdx9tnLlMnE4rTB8j+RhB
2PT1UlOz+nobT7rMtNyYo5981eRndxJiZiq1LKsRc65RoUAQkY9BPzcRWBHyZlG+
TUsH74F7n7ZkvRMDkXyumuDoDmKh46resPCCd8WkeH1NeaKwRD4jfHtReECsti2z
yj1jk7MNB1muPdZNxeYoQrwLv6B/HogXYkoW1TsvvwN/jX6JyqBKhgeRAsxZ7IlD
7Qas6HJ41Nerb/evTtu5Aef3gCLvTYHrgMCLOOkzkoTwUjLWE9ywj47SX4r26BJ2
mzzo2pkkyg0et9lOl3aAB1rUhbzcJd7oFq5yjD3tbXxANY76z2SJ+sPATmToy/yI
bAtLJ4/yRftktlfRKNyZNCCo/u4sCVM5A/L8drVvenP6TDHpJGg9SplGRe7czdLb
IwP70zaDeXlWQEdJz2js1TbveNA4vGhKIJpjpctu5aWy3ShwdDSfoTmajMhtlddr
FURI0Z5Z3JgjYvSAehVGaxTCTcwYtsntuvNQ6YNSkaUopTybv9XzDi+BTJgPrPs9
1IZTySSYiyaKW0+G7VcQYm+EGUpk40DXo963T7iQnCCfUREKchojocK0Rb7FSEeH
bJVlkddC1XACCxGA6nRDNAJ2c7F2YqctDHuzL00aswW9KpEjh+W0Jco8NUraGD5D
Im0iudTrr0wHZ9ZlkBp7gNYAksJZMPwsUkJQiVzEz8Bpipn1HP6WoLtZd9Mb2bCJ
FXYvB0Yg2e1XJJl3g4uemdIQqYE+fGSB01bUZR6tgxFvV+6I3WJzMBrpPxhaqQ6+
P6fnsJiXkFrBiG3dxWLIPw3VaA83B0mjNx5POd8asJwmUtp3xB5N12Q/FajLmPOL
JSOTueLhUuGk5RanG8zPJ/vT9rGwFWoKK8zGWafbGb140AEtw+Lok6TleEbjJpwR
wOI9KdXxHxqvaQWJfIktA+0xx7zlOaLPxLxdZ2awFl6sK3FTQ5/xddZvKi5gD/54
KVv1qOjaev6dbxNZ4XUq3m5qvm+1CjHgaV1GGKiRXWqHuzs/DVlIbOznQnO4HQv/
jyO+bhb0kMGot+R2tyuIPB2vnXr6XI+zCIx8yMOJUNTn8+J5N3Ui7FVvkOGxMf0c
VsJleG6ZF/gRitqCoN4nEgeuCPMWfRRL9jX+Ukb2Zr46OmH5+lOULT6jHi71627L
CwQx3VuIdJ7b1XUq4QS0rSIiAN+nXoALQFBtrYAS3h5d61HlOsM45VQI2w9vCs2J
fpmTIZfRkur59A3Jx9PbZ2At58yHi7bkfOOjEv+wC2SpBnxk03dsvNeJSPAx+od0
19nZCG+XS/k8FOnX1Y3zv24KTojtIYrX9+2Ot67DSABbEwGQMDhtRdXsOXbI+UP+
/xkGL8QtBUIWzy7FQfyeAD5zep4XQtItJSxho+TugzekRE2t5LbEi6+XXdB7QBz3
vauqmq0mp1mIYoXUpMligQxl6B3KKOkCCuYR+/DvDrhyZPhUCWPLBwGxw78bU2T2
aYFyNS8mFqsZVSO/bVoVzwBpCxLlQo7mNKbepvhvTIRrp65xzAJa0rd6Do6Ebs+J
WgWKyXe7xM7/cUrhGPpuLdci/cZ/cOIisGnOgvNQblQQ8Fjya79dk9P4g+B6tFD7
m6S3+UjybQQgYh+NMyVsj3KfRA8ZwlfZwFzHuB/VM+jTDuu3ymrVauMX5V8xRkri
xaQt9Mm3BZrIbfO1/vDhBCW/qeq11sPOL7+25jfdn3sa91UNTLMi16bYYNPw3yrR
AHnZhJeUvCdhAjLjfNibn7RWdUyuTkT0F/ixYxdCvUFH0rp7SYil77+fBsZ0N1eb
rygbYpQOJbxqLcUeXCgq+OXCgyS9rKv4O0ZcRj43OAoijfgd+cJQN1gf7C+3Y7vb
TPhmgbcbELT+XOPQhgavJQydp4wRzcBj9bPykroaLvGiPppnUCeMiS3kHMyOYP7W
Z4e7G6EMh3xRp7wd4TGFZQSntpJmTAzxTcVXRYz49lWy0encFQWlU+4PLVFqX4rA
BtXY4UFUc/Hs1CQiEpyceaznjf4M0vR5W2Vn4vRfKgSEhBbJiUlFRP8l7q2vrmc/
MQ4q7UyZjEbNTh8rqSHP4x4seOGWTDR2OmEiklW49rltVeijCjmoHMZwUgeqXKfX
yEk08+3g51i1ZiqEv50EmmE2Z9GFM6khLCUyOT3bHMNtMK+3dn0pGWvAES0Ejeme
aL7eNpGYUOqhHB51Zydikpnrod3Zu4p/sM0bRBa71+rF3chAZN1GAZ61udsNWT+6
CVFphwJcUZZw4qcIFjUDJZFYZbTK78VQpx6I/kF6k46vnow74HHXL3nVeeUDH5Ss
z1uphK6L2CKCeZU3FCwjmX2V/PlcRHYoC3ZjCB3ErKDBtoZMUggOLRhWjmKUf6n8
o7nFLiR//pCXn/1DeMbYukGYfkv/Zho3u3lBU4cckgj8T+8+XsNtTG9qF0WAkyWk
D1FodnGREOott/lRDmKLgQqCOyzAvqZWroj5vLY3GlYT3csqutL+EGVHDpP+9Xy/
Y+FKLPbGfElm65DvlAdHvZ1Bn1lu+gqCS/bsf51bXFr0M991hWveGJ6Mnm0s5yQf
wALppT4cEa4vlvsHjOBWnK7ZT/8CUUgZZo1UZ+cfEjRsJ2G9ogAu9wWLpTlDHp8x
ctexa3mL0IyvdoHUqrrY4AtCElw+rToGwPscbvulD4jPcATPxoMV1qmJaXv0JfiZ
ULXERNU3GjGmd+u+R7bzQGOX1dZFVSHIRzIa0mNnCXlR4Gr65sCsiR7XY9DBOGxi
NAceAbJ3MQHAgCMRCconwSFBH3EdJi31wYOoZ6XS4HeKwPIjKTtbCZuI29ISym3k
rIA5HcteGD3xy1xdbo42A43OoBfV9JVbDs4jU/UxVx0LglWQD6IcFAjp/4baOhIc
ABTgtEwSfZbVrg+aAl8vBQ0y65s/2c689JVOUWKsAZw107d8v8HMv15J2863bduv
vlXawWcDvfONU4FgFU7b/fANuND4mVZkHmcwrlqeKJD5W6NkyK6n5nUUTMfhLbmY
ekveHJ+vQTjEoYSMA4KWVKns1PP8ycVAsrNifV92MmpnSTLo5ZoqLoqqnoP2Gtkc
eYAdFPR+YWx1QxBhPidsy3lY+iESRO4jDnSjWtjbEbDpjY/ZSVWZLkawCgotl0pB
npLXxeX6gaeaik38GihNx4do5yAvos1Lzr6pEXZBTP2L1FMWzhmHiH9Zi55HpsBm
QOL+1pfcMy1VL52gFQEABNjUV76ZrhNgkUxf+xp6+TxCAPJ34nllk9TC/LIihwaR
/8XzS010gKajtLKQHgDmA2MQ5vTGHwy1ddICVHsZLtOIaktzqxuDw8FNy8OU82xB
OWGR90jTjwMx9uc4HEMcZQOc/Ui7C3p3avAyMYSnOzW3FTBdl4WkC78e6lnOaepb
mt4SimHBwaEKgsJczhTuowG0RCgguXXm6edASc01aDaJEFuDp15CXy8+TrZ6htSp
ueOur7Odx6XRRC3DvpDkEgfWdPYhsfSQ+jGGU6MjgvR/Mq+zRhiSVr0ima7eRMkR
CIOZTZi85bbSyC71LkNg/HkGf7Fj/oCV/AFBrNd90lW1O60nXvnmPrPlFlVz9JQm
lsE5K1l8z7V0d3m/ojciMQI6NjMCY96wJ468lE6yBOWEGVRE8Xkzw7Ar80UFHKi2
NPRbSxzr1L3KbW8mWPiRiHI8EDD4SJ0VfPMAXkCIcawErE+xdWx/48F3JixkqKlI
SCM6mHqvN+sCBQ5mkuyjnKM32c3K4oibIj/yACt/DE8tupp/OBtG5iMHSz5Xu6WA
tTRiONdtyuarKHe5MNG/JcoTGoHnhUOXRrEbP7wbgU0N6uU66/7nmjTNw68BJpcR
9OjD5nCJBjzcLYd34178u0s9e5b9N3YtIvOzlRySaI2I+0Ecgurf63EQhDGP0lAx
7uaFtb5YM8EtpRcHrg5o7xvtXHUJHAcGYFsy+BMbIT+fuSrPjpQ7VUDlNmLgyB8p
9h6ViLrHRN3SeE8gKr7QospC6ctOVNaegujht62cpKx+6VZwV4sy8jNlV/EBCZIm
YUgiiZkoTw23PvYZatwmktr8SOcEDib3Ys4/23wrfa2xMyQyk43XXYRHkYsxoZi7
wBR2yhmoxxNfw/hW9vHt5yUWlMGEEm7adCg0cZTs6aTaDv+Ob3VZtWUL7TzSQQH8
VyTaDOen1k9Jqp4ch2HUlCPrWrNYGZ+akpsf/3xveKmJyAzGAA5K3q3cx94DdcWQ
qFPvokfEbJ2SZ9CScgV7U9LvuejO6LNr4wKMUsokzUHB5iOD+w3CTmk47FZ6hiyR
K11xligvMRjd/ZipuY3dMXegIhqXXtFdI6jdfTtvYqw32Tdlli0h3KfQm53YNsOs
U1L0Bq+vSUgzQNM8WRqXjiJcJzkHuZMhfyHYPmY/lLB0iWH38X2QFyBQjpXyQjIm
3o/1FFKuwn4hS7dJXmvMd50OGpYQNvHl5+ybIpkYdgCiHBCLVFizLN0FtToiZiRh
+2nnDnkcYtAaTIvfuCb+35y/3miOVsMkVWwkziSZI45v+iQZUz2/+90c9K6VuKlM
zJTFiUtC4UnKWtQJn8Scq7pbaoQgWl6nvFUjLrd3h59OO4K1qs6ipDL4GodSxXkF
Gu1IEiOyL9iRfI/USYFSieT1xyViaf7ljM9FZvIO9/mC7is3GWL9P17Scyx1XhEz
6P00pZb6ZkRAHyyKKrwJih5bxsgk1tLdPH58rXJ8unY/t9/0jtOC+EaJzLfOv7A5
fBHxYaFYfs/ZADj82wjIWiJDNlZHmNsXqpK1dYCr5VNeovmTKJe7Y14jytF6qe+H
wbpw3ibYVB62QV51L2ZnmOpQ5OABFVEF/t6nZYWvRZsKrMYo3nDZX/HTJglg2KkU
T8e+mitumIEawZBr9IB3DbDahknjqKMcLBeXI005QfKAH/iHmCLFTeXIEGWAx0Ys
MO1MnS/3DvlrtbZARn6PjTnsP5cx6oiB2jh5/J7rTf8QQAYSdrtQFnEswhHBiqkN
6aKuzmLf2V5ImdOwGL0tzDxcLbveWs/1SHRlrX15aId4DY51DvNtv5B+nZkvchPR
09OlOXlCZ+tsu2yI1b3W1A6MBtmVziCKBZR5rjlAJS99NK9wof4xaBz0TifdtPJt
s7cv5vLrOefeLTXaU7zMsQrS6N9vZf210464IhawQGqnAiXDuDg5Kx75vEc3aLMo
HejqKLTLQ+Sv1oQw5MJdMICKj688EpgvPkdyrivnAhW8cnsK8WUzfScWZxlGYMsv
fjevHR+Yo5iIIWkPps2q2nCkSMSYq57fqpvtbX4xmBjpIZcQpnB25Od+3nbx9b1n
tqLrJz0ME47qRVoZpgSbAlPe3uTwg6M0H1LTs3wrh8Ds+4L7XDSKrwDlpbGBaESw
UjJ01Vk9fYK8pl8vqp4m1tMdO2liKVrKVlz+nhmjG9mJlpojtrKYoHfeTE59PlHN
cHm6GnS1eNhkEmvXpzkkev6y7Hl2QJeJ1IfGUW63gZFMRP+4x3f0O6hfUroKPxbp
2CswFPzcenxrjj1l8x5YtRIAH9blPqTkODWPBCZydSgccnMF9MwBSjCXxcxchKEZ
zqdlyVADOr/2mSD1CtCFYJxfWo5KK+I9nJM/aONKjtGx2HIRGmCgnYqloAsdY59P
lO0awUba8ZAQRfQKS8EFFRpcYS7DapAVZmHCf2PGkises2UVvYnZO4NvYvOUL7NB
L7eaniee0nMrAOx5iHtQSL2Jm4NNvS31Ff3DdijFS9qsN+GIExzw5t5C53qIJZca
CtjqK3Y4HxGh5UA5NP5VttWfgFX0QPFc3ZqDn7k+kfvjdNQA4xWKrQ+nNx7FPeNc
sHKXhRY+Vq43+preJb2u5BAhvDZTyK9Z+hEWStvd7cEJz3TlttCb2EgtxNF+Lyoq
bpOOYfqY0S9Qe3yJhRBojEq9I3WUwRNlYdsVrFKsO6jbcVbzo2MtfA72NT+oWbV7
0+xtGXe02UioXCtDgF+yoZxnEaNhCIgPL+XVlotdiO3gnGmpMMydb3peYAoPtLTi
mGlSsQsg0BeNMF6u91/V+a3/e0ZcacjomEcaOsCZUgFfvcoNEEleVI1f1P0Gwx6q
4uxyDZcTHYVSuW+KvbFV0AkGZEa/SJmGNcLl2cOhoA7YrWwE/KfaVnWs7lnd6hju
b8/ptYYlJDUutjR2io0ur6f2FTE5VLBKfKN6TJQVo5ZsHhlv43584WB3zPZp2ul5
4hN61zgfkGTs8ktaF+pqfCgw1Te6ewcN25vYCa7aRuv+DQUoWss6p4IB4u6gpAt1
HIjI4XH+wNMQQ2h9ySTL2+MNw5xoONYm0QV6GNlFrblOipBrVaCFO6tAEcyaXmO2
EUrTN6gjOSU7tKd3fpzseN9m4zZ/sqNk5XSxbWLIaLEjVhsRuPq6xgxjLlEnylN3
5v8heYJO6ieFXn3QwY1xzn/t1JigAUnOTqBY3m8T0+P4Dr8EWMSp1mTT7aSqiIVg
x8aYWSRD9a1HV2Wn056KOCa2o1naI9DqM8vb8ALr635a/v5nLbeUtm8j2nXs/cok
AWdMtXND3by0CJQNi+jT35SuTsgvS4QVZC92Y6tywRqGDzbLAsUOakmHIp0mGnja
1RDyb/K7pp7dE1aVOYSaqg0Lscwn7l1H4sWLZDMtzxcKVZ36mGBV8nbm/ENdA3hr
rXAEDZzh4XenPuHLdMSTbIqSyYU7Hj6gUt47mmuytWlz8W3Iz083KujEX69sbLmb
VgqB0AWwmQIsHDQVcgEBqzM0mJBA6DIr1oLciLhZMAyZQ+0NbzoapCDz4TZDhDKi
LbDJi48MFfOQeRlEHX+WWZhsXuPQ8+Cq9j90HF5hapxb7iA3W7MZPbw5vEmAMkgJ
vIYrRAJAjgkj437dbkQ0LAG2HJJgrVqQpnpv3nb/XzvlkVYjQ4/m0397eczHSMDY
AKIpof8Bf/7nFX5vNJ32L8hPHSwXlTPjh40XJrT9bE8ze8jHEPik1mkDS7ZQYBIi
CFa+VCq7mE/28juhgshTAnu7Ogq5WRArouBTpl5LaEcNfwxfyE5q1lrWOprrUXFh
zrmz0MvqjlarF1o+xKyB1NcS8KL/yEH+/cMdJXBZl8W78W4o8zkFCzTgSNrOkeHT
dEqHrZlh4gj3VbSFl2Eo8JV0EkcqkeqDQqSgmM9h9kwZdb17VksqGWlFzHCnFlJO
+IPnZfFncoOe1a5rpxdggkZDqc7xbnI4gko8PyoPiOhuzb4h44Qy9QPKG2ZJPbm4
94TUmC/hFPuNCd5VCsYc1YmcPXva8HD8NagM2OcTfxpg/G/RmI1J26uMjgpa9PW/
Tm6SLA1lrsOmdf+ZU0BxApcQ6z2pw+Ye9DxzN5QFp39VD9dFdmBTTZW0ssKSz1Nv
nulIpRbvxB8nCRUtHUNDlzaBpXHGvzUhZk9huS51n3fSE6IqBT66bUuPTMBDOOfC
fLHwbL/nCeF6lSS4PNz+BBYhjZoPZYkY86PYJ0IMaCa+tXSFwcoxXpnLEzAaj4hY
3T0RBFPPaD6kLqIW20rOsNt8t+EKuJF/97gWeLM3BmTsJ+Ux/hs+/RAlfVpOwWG5
YFUYh5K9mnGDNDAifBmp6jyV/oeSmctqnSoSqfhMJp51GwcWAWo132J38uG0lmqU
PEiKbOo0tVsLdFGCGYxybyNbKrhHju47BFJgatFa2Ack2KJOJOjHWDnJ+lvbbxr5
/oj5WDnbtsxCF/Dc/qNVUnPMyx1BSF1fXkp6zsowrFdoSunjZPBDnF7nawChBiJR
PHk9D7INj+o8Ji9jdLR4fV8PNd4KZbu2RN3sNQoxNA4vFey4o5wMavSJyJfLdmjc
GGaMlzoM/66WQZ7hlLHP+57wsmnB8wZSx0Hd5bVGA57p5yuw2/17awNf/0+7S3bq
w0JqBgblp0XHl8Q0prVROZOV/LK/tI5Qf4h0PWfTVeNDPD2JRID0sPBSaQx2zrI0
ONNo1IyFnhwyrr1qbEx6/VEJlouM9o18d9STp2AWx+hao5aVN4s/Q+34/K40c8CV
rHOW5L3c29stXSLyGaaW6/VQS8BbUzBOc6B0kvp3p3y7gqTKl8QF1L13BHbNe/mC
Zm4Dn9RJ0zKo7xiuV6ZwR1aIaghWu0h5BdohayScs0PEcMuaFhy/9XSxgmHWskT5
THswmfcupvetvWs9JmcoWyZCFbyfT+JV7vI6gQua3g69XuKYnoXN14CbXTio6KFT
gf6mcy2lAYuURRTKRWj8r3Z7ogYxynDBzPHN3orEKu0IYUByiP8H0Els8i2nkTQh
kBrzVI4GKG8KewxtevAQD0qpsrjSTBnanPgeEDkhXhFOZ3teMpstpdd5d1k7rqCT
h6tCyeVrKytZQxNd6jJEla13EfZlxCDtuRYE5TsSdifx6YtsWk7EOqQ2CCAbCDkJ
p4Af+E4cquoGYCEJIWmuCrwNGTHn6JbYZOSfx204B+QWHVb8b7/kCPb77TcFw4r1
lnY/mAtXhQ5dqV+J35tCfY1XDsXAFL77wE8zyP42T52oOTmqX2Dl6sbihe0TG4lL
6UCfMAmZ5xz+N86DP9QeUMSaVdOdayezTHKnycR8mWHop640r6pqcHOI165S38+M
tWDjay+zOxE7PJdlmWZ33RNlu2r0Evp75gO1Kq0uTF5k9Jvuk2YCUlMjIu3Dv/nu
ZHUyg0WrTM7tIVerBkC6un8arbNiNMDHnop7nCFXqmQLvMQjf0wwFbvhlooeWMgX
u0fGMU7FfHOYCtvSd8o6lDKA92uyEc4K83QrwCZB6bP0tvqnHJJtGpCJ2f/cNsfC
IHA8G1rpJrq6EhnoBNR/E/tlL5ovsKSKFury5TmbwBCbkMdIuymE1vSYe6xwpHlI
uPRGQZEgYnfzq5kYMHcIce1kW/SnV9jiVc3trzCL0b+DbZHh31zV44w2IjTdOHvd
eQgdWEAJxtfe27btYlaSv5gQtDKKpIn63nNdIZtErXjaV+swqxdu3u/IHK44Nfxu
cxUboqDCAHtME2T/z/qpQqk6qG7as+397L0EEmXYnwIm6iMXqWkqVJwgXR/uARpI
Kt7bnOk42+B6PA0gMtP2ohITUNBOuK+WF1PWjKugSE7BjLImSyZCnEF5Xz+wc/+q
lq4qHExJUBhV2a7osLlbY+ebTzoOePou1zqHapSWQMYseANnufctvx42vzNTO72g
spIzj7fHrp9nIo0HJ++B0sebnD5MEV9b4LE00148v2jxReMmiw45XHDSmVU12912
jNpt8yT4rgGg5xnnq3McFNF5xyx6rwscPz8WC/N743mMDhqb8JdzxoxP+SVKrBDW
PKF9Ps4YekmKhFgtHfmhqtgDhgQDIlu5TOXiBsUO0I7vIscfInRAaoDGk0pu1EY1
+CrIxF/eMNPj/nzdsbcUDCh/ZDakb3pv3Ynr6doi1UhuXUQMX9cD8JQDMIeBKaJU
2LQ1rdLTU19C+l1fNBPZ2b8iX23+/y82G+/nq71MpwEC3Er4L7p0LQEsx4yzyEHg
AUn0J1cbTKLxsytrj4COBdsBHOb27VaisLEY+C6vMivg96HyHWq7Ph2SWJ2D02nf
ieU22WZNfllqQbEU73h2xOwk59t0oZEi5hOAC+gA4MkZeJ0ylo8zkwmn4B5oq8Xi
3EQ4e4PDYpWkPhp7Ju1PSTegP4jJY/OU/ejsiU507KJuAR2kxXWUFb0i89KPUiAM
UCvgxgdF4XJ64FOVSzsXuF4MX1hmKdH2sLYdTEGHP0wxqNpupELWrSCH5RhIPL+w
j4P4Fkh3gS3wysSbOI55B2XrECO+xrTu2ttQG30tlyQFmyx3zOwvihjlrtiCwi8v
JCIX1FmWTgAxu+F8er2SUnwua6w/C9N/xpEyQ9RsShnplr3T93+sJJslOwr1jcjW
XrsoynusW4cnZHl/LOMC9ByNp/JD5RF8OeTJ5Hi9+2FJpD/c1Udl/s8+BfkD8I/0
91VcUJtmmF88oDLulQqHcnXsAibZj5VrK/9BtL4c3B+OLDdP1vlpSgnUPqsRJMYJ
tREOPYPVwBvFtMr3QdRnD2SAHk6mIANXDIqxwRBl/5MG9Whr7bI2WY6hUuAGqFTj
FdIhRIMD0NrVeDzM4MYbRJYwqjJOQvowP5HWa2IA+Vo89OH7PKx/c3oxaWGcsp9O
Fb8KogCYqC/KAWNaFFNws7bBI52y3XLqgcPiT2yazr3BXIgaF3BOf2pain22mUXr
Y22BOV79D3e3SXSOiwCPHUbdkv7be9cFWGS38QJCUKsD3THScMzVpo0Sf3+T4SV+
ze0Dfbqmb4Ripg3EVPhs2S1WA/sU6xwsV2hArjvhYN8YbE0GUv39FZOLQhDOJ9A1
aZoHFnZN6TXZqBSoqtd+LbcXdRh+pi3uE/xcmj8Znh+IXaoY+dTpyJhK27tpvakg
p3jKP+SQHI7V9xLu5XrbhXcuxs2g1XN8jMY97JUi1GPzGm01F3/cooNCyrOdJTUp
P3hW0p5mQxsoaHV8QcOD/q3pajmgFST/pshctgeVxYVBrcHmsrkbT9+lvfCuzm/s
PdENa56iI2eHZWhS6v404OS3GfJ+ud8Gao1icgByVT9+GZOnDBYI157aiZ3/ookq
HC2vtOfr4InVCjieFhrv6k+Lc3i244Kojr9nrRHRCcgx6v6Ibo/1RM6PBPrwGsLz
tBdWjsURyhRFlV9IvneVL9rSFG2i7O9QbGuYfxTnD56kEnpKSa4M2xWJxG3Hue4M
10KpGds1SBSZ072dLD5r3j3RS7ctxHaX/OCELvJ9otZiixeq7P47HsS5iLfsDa4Q
V5VvKI1iziFtdDPIzL2+FcGzutb68B0kl+LCGt+HVifPm1d8eDa4Zg6L6QWHASDL
nRocbEY1bEUtHuSPV1HPGMySxW4mEp/T4PHcU+qQvxWhFsdLStajO8evGsJ+9MoC
9R8P4f/cHJ5OI8AYk8uiy2mKiU/lC1DR+8Iiztbb7w8RWXaBTWM7MEP0XpQL/sfd
10iN9AmxBLQypMH18EsRxyPSc0exDhPr0O0USoZuFggBeBWY7F0Tp/YbadSOxY03
njJAvx1lkEFhNDtReB4/KmD0iuqFUdjgXyfNVP+CLjW0NrJWPsKSs4pN4NogdO1c
avujE3gisgWtMzAfLc8bDVMYtnlEi4CVKF6RFKC991Bg/xuennUXaG+SnpPkigY1
rg5L+QnKsYDvtEBwVGsgSibmHq6nh8XNZJcsmz0t8XJV+q7iflqSIbwshBks+2+C
gF/iN1VYmxpLi0q+E7Rg4bPI8/mhB4mY7peH9WuPQ9Y3Cke03Ci6AT2l4nY9s0Kl
8AvFWf7fvakiC3Fcc3RaQFIaCgiI8zwU1LcxlSCFl6yCvjvv8bmVKsSExIRH7DGo
6PC9ElT7zp/HdsXEDRjgR1X0sJycRDeGLclcHl5KbfNJqyua1I1pp5XiJvBFOuXX
i8K06dJSnkCRZiPEnU8fn8UEBDWkH+oVvKwTtaS8zfPYZVgG4lAiP/bas3GPAsig
FiA8WuN4CCZ46hhRs2g7ne4OJMHDJlVnv1CppHMfITVA0ZqRX5jb2fBYDTeNUaJu
rbI9buxnLv8zQDUULUPAFsi0uOIJjZocAH71qApjr+3UbpZkEgYzSuVpQVsdWItG
G75pseC9RoWZ26/7qqcVm+bS73w0aP0o0IAs0jvSzvO+SwZ+KS8VBFOHRAwCLj56
ywhjafgnMZ9Dni1xrGn5kvkXU68UicSmixgba6WibhbYTql2TULMMBu+VKXznSaX
pzDmppCpmv/t8fgyoUFFAOTX6D2WqtSadotzyCzQcv4Q4DpOtm5unvR5UVlGp6l8
xhL0UzoR1xMrc4c5OZZzziKH2rQ5JrufVUENPHhAgZUy2LKCUZiUmlGhsecUfkCy
A32kgvHjnm0mcdV7k2OlTgp0QGJkrO04tfel3AuVBCzdX9nADYEw6ghhbXEpRM0i
zA4SvmVuBJxyCaeNyhVqRlqDlqWBM8trRyAts1/GPrxJSUOdPsHjGsClypwaDC/v
UiwZbVxORBcw37QFfi7kOQ1vxFUEes914nm4VLDcWKn5rvYBLUGnq9D63fCi9122
6XxQg6mNHcjraZENqB/G/rkfYw91FxFwWHVV82ftC8G4+lLDsEedHMxnUftzNo2i
ZKm7GBnicuhXpS87XduJ4V7oB2qB1tbt/Iysyqfe5UoKTqSi41PJ0dMxgYazFE/r
OgEVHd5qoPe6tZ8oAb8SPXtWyHjrloGRo2cYXPRelg881tVqi8toJbs2tWqnOuja
cruhqjqfcLo1k3b90pztnJblBp61cI4P5ZQwLgrcekbJIGj/E1w7XMwYfM5D4zfK
7haMBlpPbOw/797H+qttb9AKC90jl9tf2uX3tHBjDsPbqW+kw9nrAAdcHChGu2IM
c9/aGLpld7grPAoj4ikS+j6u9q6FRCClerZjamtXWJwd+65JpPN+1XjY0d4w9Gr1
RbkC/j4TBrFxB9ieOPPCwBSBQNv2p4VXsl1PeyaLTCJGgaGkA4FgCn2qNhPAK4hn
qV1pyNjtisNykKA8jy8w8D9iru4oh5KWm/x8bosj6TXbblWyXGV4MEBuIay88Mn4
xqemoZrhsZVndj6hsmVE6YUyKhnW2BFuRUG3bqRNTZ2/ncd3o/UXaWir1n5E0IFS
vlvcUiiweYwq9exkKPtwJ5+t91AJsePg/LdXHtJ9UebJLFIUjTsWjwWPQBCt2ZJm
UOwi1H0PW1/FXsdyVduoXI8jc4tM6Ud/4Pqe91lD4yo+fmw/Z2O4JOnb1N/laZYp
eI1xST49DwS3Obxs3avozj6X3+cqsqRbOmqDpMeaRJStZJ0nHpbq7r+JLyIWz9Nx
62RyZp74G+EgrgaeDWnE/8t+rINL9hHLcxbi+kPHh5KW0OfG9i+DkX+sgwDr6H+O
A2KLm2wG8JDE7lllT/OdYfH5teyAxi9YHuP8ZY+7x1q1lp8VAefWWSrNtUs9Gedq
HAZzlyi/SuNaHGRnJYD3KKvCqQnsZc5HhdrMULja2hvyAtvIRvKwjcWVRVNJoPcA
pfGITvD068h1YZwmAMpc5fBgSo0KEN9uMZQWz1NsoEQx6zkYC4A7BrPxFAz4SqwT
7GVCy/v5HGPclBwSNxfXKw2i/DoG4zSsGOq3u7xmyJ/4J0GxeJ5RO59mcYYN8QlZ
fzd4NWQxUgm5KV4NYiALqR1e47xNzBtiAvqzczIOmv9QSBFlO7LkR7PBGixl34EP
bR68UVQUqmUmB0gqzMHE+RjtK88V/i7ltp4pl7JdZGmJqT0HjZm0bNw+cUBpfXPK
xHZvfCrZsmwq3gZxNwlEgTfVa9FES/ylRU39MVddsAGJaLuRaPRdlFoigw0CQ6nz
Tr6PR7b+ozhaofSCrAbNsR2tN1fRvQ7cCobpaNYwZSX/blwV39IFeh2JXQsMYYCH
/X6GsSppQLexAWm8J8GPKMW1rU/DrnXBBwMIF9vWoNP9ykuzi2ujpr9w9M0GonfA
1OfIk4meH1QwhX2Kne/Toe+xQe+ySb7UHBgiwVk0Zq6T7Q5vkXs4VT8NTds9DM3q
Eu2leDwKzAaVPVxK1wxpUPvitb4PRw2zeDZKXP5ituvE4Fi0+x5f03/82zAsTWB9
7RqTNTdBB+STutItW2kE/zr2f+yKUxZ/GtmXteTwRNHK1PEPI8PPYc2Z7J2c+BVL
uNt8w9sQteJZEAob/51tktxlgLViEBIASeWZi8bwnqRfvMdC9AwST1OYXHON8uHE
EfnLWXaYzitvZ3kPuJxq2/cwbv8GR0/CqV74dKjZB49Fan++B9bMZoCqhnNQspPw
wR8mBFNScuhGct4WbxmFgV0+uiCxHIVcLY7avqd/xeExvAVefb5JolfD0Sz/XuOZ
Gb1NSt+0voPGWnJdVUIfuJ2wbtIRdulP5kpceba492NVC09wc3bB5ZJlz2o5/1hb
Xi3F25xfY3JbMTdhMW5igwdc8z4OlfHVnQHEqWZCIIbpKWmeS99xQhQAsEkgBCt1
eC1H1WZzq2PltQ45zJ2URIdmNoQV6hu0oivBta09wOg3jwsLp2JmJnt/n1rTLafO
nVpYHyh1Vk0FiD9Hx94WwY6wVLNuKDMCa6hk/+Owge835jji2xax0m/IFmXAjAj4
xSZHZt6du08lkgzDqEZ+aBqhfyMCtW+zFv1aDLo151VWrd7aaaQnsKsuS81conWk
AS9U9/Dyv7jmBvATGulR5yjU5npiqjK1wEmgfZjs1hwaHXj/ufdZRYNiSZxR3U1f
sI8HBET/XUA1pZweLitNYx2uvVznNpT/3DRKWtrL54ohHuLq3QBo+X1lg+RlOPfC
YaY8lly6HlmBJbdp4XH0VlDNN+fuZ2aGIIYsvxyHu9kwu9uiVXvYWEUamwhme3E2
4dW2UeoCXqs1/irKWLrl9f57RPFm9TugMAvvRt6aujQwbj42xIEFtGBuhgS4Danm
WnW6eyiszTcB/HRaj9jSjZmVblvbufFMVEufolveo/rpfFtiD5fuNqBaXuLDpsSq
PmNsqUm3znoLU6txHGM1LlIcrOg85CmpeQDeNqa7Hj1Hz0ZgnMoYQ+NWAAIK8B4I
RXd0mTPkNVkJk+zlpFDd0qt8rx2pRacnS4LKFJj5WYSeL7Ts/vmNu8ddEoJ4qQMK
dshG6luRwJQKtM+Sjvo0hzGNmIqVFt94mCgYN7QwdCUU6k1PB/NOqcoKkfCzlkXc
iaBJ6WaZzeb+AIiPN4si3Z5entfSELTno48r3TNIJ2FC7Zugz1L+fkfWYHh8Tk1H
/wRNzb/WARxPFnQwDeMxniN3ZNv1w0X90eNfbMke1X8pvIhaBJ8/heISL+zMp+8V
Qupm6fnkGPBit8DOPwoOjJLXGQYNBudBeYdn0JzXf/eC48zdZcUsnSpoPbwxs6aB
yY6kMB1AhQdPgkbqemQYooKAwGAL7yl48fLiz5JGy3Rk+2ZSseK78KwMJ5jd07v6
om+/7NBzGwVuXSXwaQDxTkmhSzqj6J8hrbjd6t68fIvak6F5SShxIy0wNTAuFJ5H
2Q4B5364621BwcFacL6jr4UMK9vXH86n4IOTF6vBnOggKTktll0WsDa1lgbLfKH2
rW/r7ZgZ5eMQnjzMkgtpYrnOQ14ZLoofokamWD1MzhrKjN1jHotBZwtVNuuNIu1W
bvGccy3tCWrkHJDwzcydJqTeQODGoFJib4qP1ul1v+ZGBzErBXB6VM5OaGH+TjTC
imez1rozjkrGDriMB69YMqOWhR07YgFOeFt/l8E1qHprR0VqD3+EhSE8gWyroUbr
QhzWuzR4fJYXdZwnZjtDT9s1JBJHPcAgDK0yQgPFO1P2+yXA/QHwfQcT9KddNxvf
DbTqkC814FMI1UdeHA1RJGU0oO1MNgyFReP1wkb7P0Mb/k2qdORjF1+sX+JTD4lF
NxfQ/S8l2bu9aQhLLN7/+WTGQ0gMDlwrwCmNfRrm5eiYJXBjVZBrOPTkTjy4uOly
F7W9+0N44N1JtZaQoTLUPMT5CVgJQV56Ef0RVPfM028DOaRARyc+eVMD9/u98rFT
q093QtyRfZ0eXUNZpipVeY12UwXSQXhpyPLfnA6oixpoAo2u2O3HsGtU+98jrctM
eQRYwKQNe6c521D+1ffRiwpL7nWzAEhsFafgDjkkrIZE5TGiCyPmO7Y+sE5RJbur
RUHeg/wpN3LWVz5KeKRGmekTOGyUWxpOOE2xg9P7PaghksmWMLaTzXHa12NlZs/H
uSCBk3811DXoE6QZAvFdHhf/zTyeJm6FzvPvmrZ/o9K1BYJAcyYOqpxz6uKLHS0U
L6jo2uQZCfnzvvyqtRb1mBIT3z+5YjegGCoxq/pjGmJ5rovpiRivcEMov6Onjcrv
Pg4ErgXMHn2dv7GSjxXNo37c6HDMX/xs/szfLE9tDhOpL/inq/b/4p+ABMy1cWN/
6CWh4yNrVtZbdjyI5xB9mm4tLAg/LKcavcteMpi0dSZZPQaewNZMIO5TKfMOnXvp
HQS/I9dv4Zw9YQPKAWRAjnrm3DOHl3E/KAMMYMeqNaZ0WBTCJgF5jUhKjUo5v1CQ
bWZPYlRr0Kzxz4sgykVPUAZH+PS7WxOEz+GMeLmZ6B8N6CEjuQ28tXF8pfRJtOMZ
IFOjOSWXMpDrr5jrXkEyJp+McJh9/uCXh7rPm7WW3QCZNJtSHxL9+qxldrEsXx5l
eAL3L/xn1xi8VAUgfHLqJvcDMyjUnn7rXAJITtFsW4wyDy76aulEdbJvxNMrp68Z
MpjXYtkAzyqD9SlgiXXwzMp/DW/6KALkYF8R/t6nrrA5bWMZ/1D/bdlkMB1HyZeU
TFOat/CICpGVThKvYFQdSzjNc+QZ0ZakmtK5zK0QIqBhhML2ICOk1DBrijzdtT5s
ofCjDuSeKmyxg9T1wwTzK5bxDJaFGWhrM+Q4Yl4ziIteK3Cng1US02cQg29YL/49
LITlTC5LEcKwNhKo7Ki4Jud9iCvFx2JqwS/ye4gkpUceDm4tO2cppHA1g9jxL0kB
sFgie4d3p5qBjcaCZ41x78FFu0xMtaoVymntyUnwNqXyRvBqqyi0CyyVvIykE1lR
wjJLdNM56Scrtx7NZp6qN7QhLHgdMvRq+ig8Gzm145DpC1VJOKnwXOKlFjzFWgI4
IjKxXsYGnP1JjBJF5fleBHMP02lkiqoxKG1V4ZIax2fnO6s35TwQ54nU9gcGRyVn
GyARclt4mHuYVfB2Eo6YjymY1hT3vb//nibZfqD3+3/OwlEm4gYDtFzeQO1nVphJ
IKyHm2r2NvjML3QA2aWELYTRSg1ouyj4GxnNNdTBB06i/TRqjYkEHInlPp16vy+F
7qsEM6kRdRnSJHA83aR2FpGoFKGbU6K12e/IvA2n/kDvrwD0ebT4EK3Kb84LF8jk
N7N1TaJtbCjwEXDZE/e4Dg3SH66NgM2Khnk8JKM3SCtqU55ly2tG7inGe7PhQZJs
f0f6RuSsBGumJghHRy317VLEtceAlZSJO6gVsYWj5YyriDuELc4yKbY7S9tFC020
Osfy0dRo5tuxnRrgp3Ezf7W/qKxb0reG5GzOpPdIXDzT36qfNobMJ7JsXD5SuG6l
dRmeSxobiZqop8MVu1cIZ4OEXiXHcxmY2AJr0ozcuDxW7Vq5aKjNK0fyM73jDjVk
dJeKSqNIGfNhuivmpi/ht87M4NFrotrTzpGLtPnyT1sao1uTZxjmvmxzKet7HBQb
1JByeySm+MMT2iMWwGMCFY189nyfY+RtHnNibF+fGHLMMRIDK/zHpJLQJz+M26vG
Y4UsZ38aoXSe2xRREfqZGE8aIcsEX52ZVi8Rp2TFpAUOXdo6/J1gfjft4pluTiPz
0EWTGf8zTah1dxsU/c4UUigRh0h9YtAMURVFUxIJjBYWrnJs/bk/+4UJ7HwMzjLP
+22e93Eb+8aXkhXr+pKzTNxi/WXY+OhuJe7ee08sgT56XJ9UOZmsnjkiyO+hZT40
qZTWVs4FgaGIJgqBKwTXy+U0Tpr+wuUPRVjAfTudpAyPtE/zxQbU6mqu67pjerO8
u0mWWSR9h3oOM8NSrHCcnJkBTbk8AY87YWFWA6loQLijiOeWpO5ZOMvN87Sw8Eop
B+2Z5j7z848um216cCASspSPyxDeXbMFhAPTo5yKePrEpDz4jAQxHAdcdkmsHUAX
c9upIN8Th4Q0U+pLBaVP35w08xD/Dhz1k3in9NQTVlnv9rPQQKU6ChRrhWtbSU/G
FRPJZDpGcyp35vjkz+97Gs9RVPUCwxYIctkjsAupnKKghlIlpAKiSWOjK6zw61pr
6l816nfHL9t7ouEwI+A/osiRh1rjDOLuLV/wNOLcimwU1aNE6w8xdDHeUr1fR0I/
q7zl0cOg1StB1G4NQBZCiGXn8wbausk9JBxXbd9PhfTjVTNfY+ffs6N/IE+t/0B1
iND4OLf3u6lt7cXgv2Ifn7cAXXj4FJM51/ZgL23jpRKcT1vg4xqcx09S2fQzJ8aH
3H/1rlxjXKwRAj/vjLOkeVnveplt3FvYIdP6zbqnoMuDOJhQUC1tqXi13O4sfqza
3di9SvELOPWg+tjvdpp0zOhR9eX6Qr+hLWLd46bMeWlqMgCyHipvqxTBEZXgtc1H
Qgni3fkmHe15j3O5/I+z3LrlFqXAADjF5YEyu5F2ZFh5hfrMILIk2glGQ4lxLnKi
OfT8lIWXCuSgr+HjhqF69k2UsYkDq0s78XVTD6L+Es8epfI8pe2DYsaSiyRNQYVa
3CrYRWdc+zgykiktUPJeoajPIcrdXeRcL8TakjKs7Q5k23wk1psxc3E/wSMw5Vsm
BMA5iFEbfbJgZKM8kkpwRU3eUCXoxGJYeeLjQqm3ZMhlDfwflcDsBZi5EVuchT4P
ttVkgDWLYTeQV1KlxCBPfuXM4t6L9a3Z4f1EoFEgRYkzdFZ30iegYyHMkV4YpOLh
mLzestrGQ/KOeMO++PuDz+J/fxEzJX/KCSKtb4vI7FcpYnTJJU/54SPoupXG3pXu
iC8RdaNR4bxG3FSIll0z8JFTR4VsXd2x/FBZoV7JKph+ZwfIu70OaioULP+8ydCR
juGamz/MPNxRjeedWBFHnFy5VJrkt78ItjTS3zrXiiBgMfsh6aUHn7oDrz3hAlXw
LjHFlj4Z4vLtJUoFyb8JclpKeCAFDyMQ2FrFT9X2mXp8FSDG4TaCrHwK+fA8HZxX
HEo9uHQgVW5Nseu/xHtIyJvb3Wq+T+j6lcW6oYYezpOMRwWXLnHIWnjeXy+T0XSa
LldKau539dlAkhtiUqp2uz6/qE6m2KhMfjqfDim+p3krQ+0+RhAqmV+vTRJvSee7
Kwh9pVBDf+mQjo2tkrk74c0H/0BhSiIdty29Nd+XM07s9ej/1z2Fej2qlDezZ/TK
v1UOzJK2qKfsrxMuDXPV+SCQnbzxIwudD9XtrKwnSVn6h3vs7zlGXJYHNGiXmj+Q
d5x/Fw9r04Ty1VHJe26VKerwCNVeImbaVycF2CFQfQN0rR4zlOqKTJgBepfv0H61
cGBhi7iymKch/y45bhVBLuJ+P3xxnMRH4Xwa9icqIgOtm5n8B4Q2HFPfxyeEEjnA
mVIqUE9ehTRn94+P4tvt/mivK7q2/fa3evEX0hzEidxjNBR1dmDfuMcMb06HzUFn
nnVHaucZdg48oagr5PzpoC06L/t5gDO5xtqRT0Pl2HC13sy47uvUw9gbSoxHWx5M
UHBiTIwO8bAJEqSZX5Ypa/NU2OiKr2oONJo/5pf+fefp0ItA3v9FIJ0VCvtY2dMv
1UL+u9x+dLsXLRjn+5XLd5fLMDYFjv2lYSl18iSI1hMueDHEkTF7CeIMAlDcGOuQ
9HwHiQOqHobFUjLVNu/TSn2M469OJvqJks3VkuRiYkKG+R9TW7GREnfa6c7HaLfX
Hz+U1sm55E7578K4ineYPdd5xzb5SUnTqIFCUfOiD6I2tYOa6fG+XJu0AFkvdTeL
KzaG/UOsMMxMKFvmCNHxK/jhTICDrRzoPzq1NJNIpbXSps4LTjkBmstRpUvX+ocV
MlulQ7Xar2L8QgaJ6GcoAhOJ43BAyowQhFWNp7B7E1CHn0rtfke0ep1B6bFoBT+2
NWZsyVUHwPDRa9Qh2FSoDkdlFN94QKpuXaEapEOvt/WR1rHWvJZpcLfcSDrAB+ge
xZr3D6fQvk0Dhmmys2SfFBAtTUBGwQkGdchhxsanWHK0jL+wENcE1fjCqvZqgxG+
tg/ZiV/ydGBlC1AGYCbPFUb5z3ltBUQN2PYfXwBQFuaORHETedcXGpXllGYlbSLj
qYElc1Hv0TwuFGqHHIPKuK6sdQoSi3xbGW8I+4ec8xyiWv3VAusqG/8FNcvFfIOG
iAljTlwPCxbiCQp3/RXNwv0OqpNflsclgUnvemlXChUqXTFpanD1OqdocvyPDChj
QipXaWfgyE7vucfsZhiAyY8tB9m+4I0PtHQXSnozL/FFI6jPOwPfuo6G701QsQPw
qoYu4YohlknUKTqHTRDL1DAH2mPGWP451kuppFG0zvK+9OZ4gABSZUVKF+ku7D9h
6bxeGrpikWwV45H0rB5b8kFiCn1vlxQom5RkUEtR6g7n7V8F8v/QCNjmg9KqOydd
KYw+fNgEkue7CYVCEe/xjeaqHQlMvwErHVosQpRTwyHGFPqAznZFNO1lf1n9rhU+
PhrQ5Js2ShXBy1RA5QeKypN9emJQT905SBWcDVaMOTNP6Q1CE0V9Uw6tybJuJHfq
2rW4bBH4qwvA7ytXxqyY1XifTpHodfG4bP+SWVZC0ebtlYrZTzosmNaLgKhkbMUi
2z9km53XYtxSHlYzxPOrFNHb1uuaFs3oPH/QIlP8drtHW0nAvloPBrBxwGNcY7Ey
Ascw0bXDYbI0oEWAfX8/9DN1vzOSh4iIoJpFB178QKYu8c3NZUoaZT7t5F96tzTg
6IpDgqnNlzWuiD9TOdGhyCz6181KitwXOLxp88zvskl70oPuL2iEV3vNCHmLsAeY
+I1seJI7BuwLMK4GsnPKsIzssxnAJGPErQ5acENrd8sVpxdAugIk13TRwIaj8C3e
SaxCxvd1t+riqXLxcCOQhmo4gCTyjqYgkpj4XemJ+n86Ke7u2hfLdSh65xHq6VcT
raaGXfq48/4adFzBEkUQbo9kHbOaqzw5wQ8P1kJ0ELdoE1K4kn4drPYBghcMj1lP
i2XZ7w+2Uw/7hbYGVWwyvqINz8k86Nhj23dmF9v3e9SY0cLstUWTRYetWRJmts04
Hwur7NOQnTNCNjFApmlZeA/3vQqytuq3NcWWmKHFGdot+OAIyewpQ9jz5BW5Mp6E
1KD47w7J6qQvraktVuKe7FaHNnst16fSYD0xybrrUmc1V6Q48eJPRFpF/Q0e8Mk8
3yy8CjCqrAoW+K41jW0QYAyNkCs433Ni34B78ykpZDljEjaIk4mUbMGbsbfTJPvQ
//VUOTA5pjxnDeZ3bWpRyD8Su3VERSM2SIrzH9gqv7KwDaVpMZeMAugPp9Ay8GN4
4ItVGmj3duHbEc/j9bi4PODJBwYBBYJtlvXzq44C+lMmur5A6vitej1QFO4lPilm
f2Q6TQN1Omj/fU7jsjOCgkzcyiDlIv4/i2pgseQExerT9fYjU/T+I2KtqTmw4NMn
QW9jL+HL350vOYyGVcY5HTmShEJHFfbFRsNB/P6LQn+fJVmD0lz+2l3SNTAy0Peh
r1tmavlTp+3eYerz1Q43CRs4KqFB3sDIVroRzg4nFEvZJDS9HOmwYP06AcOV3YTc
l00rdxPqi/S2eb2HxfRDbun+l5VyTdfAjNVSxxpwah3GWQzKpLbhrXWi5Mbw1CVT
i/FmyD1OxLXw/ADHphJpnDxbGFlrZMFIPcg494GJOQamEnBuwH1dshRe4sUBi9oN
Qv+aKHyRT2rDnj4ZRdO5PG2NA90h/l4MxPzZfrQvnxnMkw51GMY0aFzZZ9SGbk/g
mQthizNq7fMMavivX7U02XYBaQ4yoD/JopPqCPwzowF+mQe2j/akAEN7ZwLSfyXD
BONCCsf74FA4vmPkMFfHgGXlL6gQbZroepY4WrNXWEuJPNTj+gou49aHXrOp41vn
v6sr7IatFwvMzNA5hPeMf2Tk4pNOGqgvYYHKVObiks9C1O8iZ3n8utLRpJcHyc7e
ZrNgaNxrfL2Sw38ZnUjSOakUjNE/kt19QL8Stq8vVV35lbXOCR6yJ0OZWfWquRZK
44bd0AGP5qDmeDyZ9xV6b8Yan11di6cEUabyqnGl/p4hfTtTdp2zus8MB4+6SCtL
T+c5SDDgnIUwQdzOz25gG8fd16zoVlsrLUuKDHdTvkn9N3o4ZSuBLV+/Uy38Ehgp
MrGBwVo00paxelxHUf6HpkRzBjZWASOP7McqZ5UxwYwpiEQxMcCRHYQbRV4OPHa5
IXXhnLtslOcXQX2CX2ORWPE+ZangIWq7+J5vBA+8FKuwiCee05MMgDenutpaODqX
O/dipXfF4HovNpCNjZVJJ1CKJfdgmCrD6s2g7H54IkiwdBXKbaE4a2ZwQzE0MLdP
pNWVGtND9BDvaifkRQYL6EQAkoNr8oH4f8AjdNYVZOzrWosyykPfQrJQ7EBBcDtH
9/sktInnqyHGvriYO3YkQsOjuhrQJLHPUMr/ePtactHCDbFWPKSYUPEsVzbKVFWU
g4Le5o/VttG9msyAZ2CEmehJrGqol4ISA1iTp4nQ3hJZz8OgSJpFZ90DU32uWrWz
9kqofziPe9rH9u2//hHrtKIKKez1z3H4hLBmIkbvee4FBjvDDbq7sHv/x5xX3kU2
Lh3sZoL6eicWH6AuHOvDvhzL/6dE0zOm8jcifUx3uQ+YigTLcCZihxu5Q32i/joW
zHave3i3GeOVFX2pxKi0Ivl6G49+qNfx3Qy+KO/MkzQQRse92y8d1zz1AEv1MMLC
qyigCoyEFLrAd1SoS5s+uFM87Xzsc+zGOEL5uj+Vqsnw/nlk+zg3WO/FyYebUgJA
FeXqVqal//lncbvtN6W31fvQJDq29U07y29YKIeZWqAyqh01P/sJbAQgSjV1l0cY
sFXfEEvyo9zLLFnewoHOF4WJO1vXSgASgRd371aqp/saE8N6BZeFG8sdgL2gpLpi
m80iULRG///T7t6e6oxExvNogh/j22+LnlVknSey0vvJBgLY2aad+T0U7dOwLoRj
4CYRr6P8iZbTrcRLgJMf+swGgBaveABfiEdnApk+eOYG3GU8yt90ElDgT6fwd+Nj
zopylAmUKrtqKP/3c1iGLkIbu5cWF/l9OBeWv18LWkMPrvOG97E9iMsTmUcuahLZ
+22Bhj2WPE5Dp3/Abk9k+Mg+uWVRvHNPwZAQFGBT8Z8IV1BOkQhCjSfTeZG8vXP+
3FP2d0/CgA62bYpU1XTZEQyeGlT6nIhtlH+oHaokbtGTH03tDom/3g7jwP8F2BkA
noxMFNbpC+FKAM0Yn4uihNMkmzNiyFSbhoOpfz/KtbkkSmahzwtURQLI8Mydo1lN
EHTGlYNu+wEuWCVNQutHNpvDuYi+YOLwAo2YwicRjAgb57sBlcusaFhWW4XiosSo
zCgfGcmfgGT8TfflGeEs5yFfRj43lluxqGrBfdtwtN5KD51uigV+lUFsX+t6rCKh
PO5dgwt7PBNzqo4Zbx8DSldyEfVZdb3WcFK9Jg5i/2v6ACyOXJdEV7p8SzAqR5M4
LTR0SDdko0FIdav7txixmTGyXt7GxJ5snmfr/7xPo2CP78EcqLtOjeShqBauBqu+
oekLR2SjGO9alpv6Z4VAONZRA5S7lzz811y03QXiBNsbL0Q6hyV4KlfuOMdeigTB
k8H2j5pU7CGy25XqzFwn4so98HxSbMj3N7X0Yrg+I1Qzs7YyCjxQFWc9ITrcbvcq
6Hnnv+65j0RfNAoM6diOSYr4IL45mEJcOqBvJhF55dAejXV4hc6F3BLyX5iV9KNQ
BcZz/nFLRcsUfH3Ut7jJr8i/828l+0YerDCMRFvuv+1VqmWhq4O3Yb21g64cRAiN
v8ObG8P+A7rsa4mIz/CA1QjPAmQ4fg7SVPCZdyeVPBXBd54Kty17vQqfQ2jkg+OE
c+PvzcoZY1Id0I15vgT8rIl18kglrnK+mf/Yc1RAtkTugz1pPNSNTavc+81DWdDC
TewNHY6veKTafHoEeW4DSPYr98u7XbAc22kVppleXTybdl3npKLgwlaeutDlLV9y
tTJOPKHU+vYVIopvFHM3dGUOdAxsf8KSjL/vEodb4GOzuSs8IWnerDwe9q72IJYV
ZuuxRf2k+LzmNIOZP6zR63fkfh+CtEgNHHnZD5DXSJ7TMvfQFGwlCVN0M9jDbXah
tYrwGMyH+8TLX9XdnPYk1Hi6G+ex0/DEv7/D84dPGNV1m7UBiJQXbludW24fTMEB
xdjS+wdzf+vQti2XoXFWEg1lll7dBN8RgoiF71YeiWgvUmSRFWBui6C5zth1PRqp
hlNy+pPJruhGpuxgJGSgH7ivaLauSi6Ts5RtthfH1nlOEO85fctzGxWu0zYff6U8
ZfRPyKjk7HV00W3qrFq6AcRz7+InKnp7UVpj3tl7jCrgjfTH1spd9tzUz04K3V9a
ZNm5IRFef2SzktS3+mUDU7P5tVol/Eni/Yeuk8EGzMXp56tYdRrAIwTFVnw2GOpp
09odkHVXy1Hrve8Y0TyveI+EFm5K1QO4nD/oB4kL4XHo9cTyOQgMw0Vc8PtNuLhF
bc2iBn0Us1hCA8GXAu/wOj10VUVQm0BmUm8w03jfMkiUbNfGv3J+5I0yMdxehXcN
K0GEedMRb7rXE+s6IiE2tp/tPOzl+XxUjRQRBidyQXMpi6DywVMK4U75aoAms+p8
Tyf98RQZQYDWHAY9zF8kc61rHMNoG1ooFmwC6uZqR6njIIUJRRsDp0z8IzxbI8Bo
Fdsf0jRn+vGhMbmST3iUtRPvQTQIJKPhuN3cQU0TbYhazFVfU3Z5VlCV0KN377M5
4EES7LYdTBbQa4X0Rd5Np72Y53ws1VBTevC3FMB0Y8EDGSqlFIW3TnfevqO0zEV7
pa8MnucLa6Mgy5zp91yJq/IVQ+WcMmBeqCw2Gqmw8JW4w4ZaS3xVxSH0rgv9RGws
hoTAPtT/kCzOta94PX5vl4t5Nnd/uUzkJ5/bwsFXPcWdzC1dzl5VPpoy88ucjVJN
nhLveiYsSRebOe+dbeizwu56AwHSQmVspfu1jpMJ/AxYbywl5vvaTP6gILzPUe7V
N9nyKn9BT6IwxQ90WIaiXEdv1zc2CjrLxoTxcqyizFZn0PRUelEMJ5dWPL6wTkz3
oQB3fR40iJs7VCfLPbYNZKiLSoW8EzcGr172t7Kszz0U0p5//I6IQOx6nAHXCpOM
KrbAodvYNFmciWJQtd5J58xOXdtdRP+I4MlP6Sz+tZZjRB5PJWcXJ+7L36ONHreq
SH5vj472s0WKwbF4qceHAo/QarKglhbATwaJlJ/xZooLP5D/FCI8U++TzUaEU4z0
oIuZ+m/RcCSwAITj47wreZqua54XUOQYMEMGYYH1KCPFXHXXf1xn8Y+v3wO1nQiT
R/FdAkPhyqv2ku40UoAtx8+ddbK8DTQHNqi06E4NEnZhFouGJns0TXuT6n9n+yqF
QOaqcTQNtsWk6h7WWEU3lgdB5gDnDoFdZs/tTjU5aEo4HbQLxZUVfNcjIo+v5t+r
Hh7cwN1aIg/rgrhRX81iOONmQJZU8ZJgZId+vWaVcPK7LiaxCVaEPg4osXGgt+hR
wAHxwWFSAo84TSKq2TTMseymJEo3xrI+GpwixIZk3JVpwyEZusvPdticZMVdZLlb
6awKgYywMZgVkF+t3Ka1FsO+w6CwUsdooje9ueucCkqELBAPb1I7O7FsdUpKuloH
QnVY0GhNdCvNvkLqBFJ/Vg1qOtrhg1xdibjHMffmaM4ew+YFE9e9UyEoXtcldlHZ
eNMi6U6ZgK1xyZLHk45DPDABZhyFGbqeIK8WKthn7QzgTIj7L8DGayxEcTzAbkGp
auH7oHhk5t880ienQ7dcHappqnGzlvzBwMca9gTVLJvmhtPpUX2t1/yFmjrkhjMV
TFqge6L3pJ0Rx8o1BQOZpaFzTxoXON4blKrDxVINdmBbL0BGq9OJqjZ46OIs340v
N8Z2c3GIn+VAxnGNgUq/z7JOQR1aMlkAE+KfG2kC7svp6NwBo+axwiQ+Ux4aKH1k
7I7tyRJqDRjhSlednK0z5oeAXyTrm3Y75VML0w/TXihOh0jqs41NgutYRioeePOE
kpoQijiIE6JdxYIeIkNNxSNQXoE6A6q8/6QUr29pDsJt5VKZ2KXJMBAp6yO5sL0+
xIm1AiG7Xnz4oMu42EstZkT7ldvw3xktvTewGRBaui+a7aCeV50diN3xpUovUCrc
zB9/T36Ufa8RrTarXL/ni6a7S4FG28BR9FG/F0t0R9bTUJDBkihIfs9eH14nbjB9
V+p7LdPgviHRZGPWyzUQNGS68l7p8Zljp4O7nc6JXM+kpZRQzIhPKendymdCtNpv
H3TiY3JzQfG+0khiH2qOiiIiUtgse49eRoVODtQ6pfMyLw47Px8TfMi2DyULoG1P
Bn3NS7qf8QzJIhtjZ1ny5MNNomR9k+lkxAcxAHWNsiQAcbNh5tIFB/DpSHPxVzPV
3Bq6rZogwujSNwBXCQzfGGkqxp+X1gf6E5TrOb5B/lGxilyW21ZHS4BDoExyST5z
kppVTzU6zHNCggG7lXVpe+c9IPMIxfiSDvpiyopdRc4vmfqCpOeyjPTM553dKKQm
hbV2Q3rPxPkwppVYP4a0Sd/ym57R6qNJoc2FbaM4qhtteG97bH5OMDLTIrYRVGPu
8HgdJqqQfXjfPcjyecOh4N50xJBOCc2ANm0mwuUtSUHz5utMWVVovoUj4F4Psqxu
5ERhsVLZhueGwsCw6Kp6dlVc4LX7kfzJfc6xCHrXPIm3/k3OjE/shubcqSu/gx/7
k8l2xQXBLr/jttPpFenKdh57YUZ/eVZUn4yix0QlygbomDYNyDZ2Vak4Z9+MfDWZ
z3M1g3xubL9gWO536rX867ZxwIKgQdwY7yy5kkoaMn/eGlA6zSh2FvDYbTnIk2yQ
ttvivvNoFAmaSrlsMuXmKnkDtqxeytlRl9JIADPKbSh4tFipBv/IV71oKpfjIqHM
dtzBOQ9oCzxSDIBC/zt5RGuj+V8Dg/0kYBGSrAPymIVCAwIywaGqJoIQ6ujr69Tb
hFvW2kWBabchZ0dGCdPkVmGeYT+4P7qvMrx4sMdNjgzfPw8diLUVK5Jcr3dR4Fcl
4X9OKPXviChRkUvLCgcvXmHD6oTUDNpAZppV+mSoI/sxqMeDFW4i0uOHjzC69OTH
Wqb2V2CXnyVlQkwgemqx+P8xNMJSOBxmsxC1zeJpJcQOlYdT1EuXA9eqV8guXwGz
qdV4FrXRHxd3L9pagKxDYfE7pLM9bHY689soLomkjp1LolcsCe2pByMmRDe2F/4n
tfTzRUru+RqtkQblSLQuqyKHA6rLJqN7cCNSoOn4MhDBEL5E9QoRV89WXAgcowiO
FzRz0Git7PvE5V+u0B+SNtmSp2pJ24kL0awFKTgR7bi34h2Uqx3/jmjr/to4CZ0U
8CJE8TPzEDDq/Qd7ieTUs2K2q14qw/mKDISj/BYbvATapQJkPxfZp+dsrfnfGQqw
LI9+kGamXDFxAfSIkz05J1sHzBY7OjqRX3AQgCWCobyRuxVuhihdpi3ClURxyYhs
89y+t0rT3Hh26A67/hQ2Y0cnqQ6KP83WKeIZY0nJ718z/F2gxokf1hZhhXefndlu
sDBOz+F6VDJop56fJsC1CmjQr6jimj9m9mZwUyHc6JFeewIDQAZuGKEWJAmdJIdo
4/Vz3b4cTESv+1W4lsdiaFAvEXmiM6zBpokx5ihmxtsit/DrbO81k/qVgPjZl+V8
pqoKTCGhgnwqcGyUDS5VbQjWpQkOPkFTLRA0vNTReaWyojfG4bvLYYk8Obm67VXw
YN4ivCT6U2GtUPxutGccM9zeiVF1s0SjY63mpUAUTDtYlRYiqLh4kuWBvOFOCknQ
Alt8kdgNK2S9NOqVketP3/5nNrHVznvfhV5qSzbPiqvARJK1EPgTb5rOK2RtCTsH
jb9O7dAL0g0jw5cxsjF0r7rDhh/ysCDXcF51gDNI35RknCFvnSnIDWv6yXZF3G+Y
2tP33ZLlFID09on4YvoztEty9emK5uQJVgMe/DqXGxJdrz2PjcKdHZ/zezuBK/SP
4zDUc7KaEIj2bfYsfe4H7yiosWQmxYwSMVZBJD7k9i2u1LNz1U/HljPYiJjhhWVT
mLGZpiJWrJCxV8uc/IoTbaloWi4T7ZCdiCDhpEp6kEx0cnKKhmuDRBA3oY9RLjU6
WjMVUVdJndkXZLlkeMNMUhbrNjjqhSSc9fSn4pgaLFNoZ24HWYgw4SGBebCgS91O
2QyXA0q5Cs9h40GvixB7uuPvF37Ygek4cOMRxXBFeqV+eamU3d3Fr+OzsRo27Qbt
dGI/Z5MKdnTbMNdKafMEmCQldOF2IGmEEDIfLL+m/xu3an9QWSpdfXFnb4KnLdE9
SeUObaRpXJFrsBbphr7lFNMjqII0GOU4lpjMPC2TQYK/XWGnW8+4HDGWkeN4rQfJ
b+TnqYE8MExcJU5t6cwIabSWj5kq0856OWijTl+1pXpe9xBpxx9OTzP6K/2EZfrQ
tnKyca/h0yaj1cHqKWDYfgHYvfVcnvy8KrLT8RTxjdG/fS+JMo5lF9oXq+muQz/J
idcY+cIUmK21mmPZl/B55o3XUqwKWNcmBAL/E9F9fanVYEjQj05VjwEbimkcdNdE
GZ/OQCtb4SImISdM1WIzaK5RBWBE+c8LJTByC85SwBOl9Fa55XvwuKRegXg0OL/l
BXw3qumN8LfvvB6Txu8nX3e5nrozJ1IRz3wHxwlsA9qK5xVbrk4OHY8TwWVe6Uzw
XC8wGPzjjDRyTJHM5cVY+A1FG+on53BiTa/xOG4x19EAdJGpeRKT3ylG2kb+g7B0
sdUVIOBJDLCu2yRY4Wy00m+qbPjayDzauX0qkNg9h5Y5sxjWuzhj0fFUAtN0abiu
fqatooPhbgN6nHidkyErc6dijfm4llTraU5C8PpWDGIOlMmFU8W4Yvk6dAMnco1x
t/4y94hohgScTpiUmT/ADvBtUGukncbMGsMdSdh3uWgGkn8/2p+MxfqygL+GbogW
zQGFxRk+2ZwIPFVVhyqWneyRTKPMz7D02rKFAqELZ+lb1lWKMLN+s9hIe9uBIq5i
IQZ0hpypNhtivmMwKJG6WIgRNOF447pRs3FIj4FvO19hKhVUq1C7zCr9yVhoqjSV
AiV16FtO/uy98pfsHyE28OxzJsUU6qAZpBFF1P6NTZdyGkb3+m5tP3rQQ/pyx5Je
gQ71Mc68bYtuRd0K97sB2vgCtDmtyA1+VkdmRDxdnFTRmY21Ho1jtBzaPeQFkVj0
ZjrgsTpLuoYqG+eCN4QAAsXALjre97CFxdxRCFvzmo3/iw8AoAoD+6kybC3KBPec
oGW8m26e087o8iPGmdRyHrDdoNN2O9q5IkfJHSjLVld7r+9JLBeip9whWHI2HJ9/
HVsnCMT5rom+xmePbHzYNgZ0XvRuoM0zKUtmBEU/vV6pC5UmHZKxBa4onUAuKGQ8
hTEqCYLy4ILBokHxu4197lEu+0ANJsSwMAWmfBRXnHeHZRH2BGOQAPhJ/Zt8RP7C
LitUbgPRdQ7956AD4v0gCibYtB1y4fsUFq3RZSb/fuVBQ8V0SZ26A+OZpOpg8/IR
l7ntdfIsYx5sKeTEVTvyMGZmLSZ1ttEE+g3DCNVzlC4xlZaXBW7BYLyBxfGv8bxd
/9i2lqoBCj8z9ftwjEZJE9lgwwKP2Imz1peY7u8bLx40AWNVri60YQhmxEMBvbdJ
lehn6/81xXQFCyAsbkld1vvji00JyQ/+04oirdd8Nkm36fshfCxOZMfmHME4oepK
ttmB8+xaLXiVoHqO+qc4Vw5eeeWSe13xu9owLyXpa+jdpPgpkO9kW+1kH1hzEPbY
Hja9Hn1WDnImMM5WILfQmlK35Go4RB4KxlLf1wWwKxN0G8xd/zBgdKuZbpPvvJzO
3msRVO6kPKPIOjW+xapV6aD1NWEp/CJp/9z/gpCL8oSBO7GfxHnq8kyBKZKgB1Y5
Tbtaa/HqvU4K5yMZp+CE1TiaW++uMpgs96P18410l9BI5aSeiiSYAxlcTcXgVgO1
Uha0qJmca6wErsd3+EKU20u9eE1nS6NklkFLKYKqu94OjKm0Ws2N23v/zBUiaWDz
hFAd4+U7gsY38Rk6bxWCHk7nM6TpxkZGuvMRAl0QHjQeJL3JqRDDaY8eQ9t4FVKE
uV8LFqJPQkBZ5w9Hcq1jQDcUsa9ygK/buMY85hs8HTz0omwtFZTrvN6I2oB+3DuB
Li7FH1B+w6lfVwRIXw1ays4mN4K7NOwqlOHcUp/do7J6DqRnJe6p8+vxGlXPqM8Z
Gpg2mH0GcS83ME+pc/E1JeFU91Jkn18kjnTHpXXyIsG4nPCL4OnfjtuvPieeohUj
UdpUP1ZtPfPTAbgFoCciFOjkDkdKnbdTp2N+jO0ZPCzq8Ai8g669ROxqIXgneLm5
dNXcDGfc3T6Nnckpg8SxNrih5v8PThg19RapcCuE+W8SDeAPrk6Nqoi7YjQjsKmO
pJcOjPALL6umUdHyjniYguq1bsNARLk5EYh0EmfCl/WubEHXpD8GqW+hBaRemn3U
paemgITLazR5Vn7WA0c7YlFD50Jh2M92XZ98u4qzsztogQKQBlkPEeZMdfeb35Wp
+t+kaphN8iR0KrIf/yDhBX/dRVDmeREaCmP33dTUk8XBAlbv0fBAM+qNNVjYLlao
h6FSvYE7/e4h3Prj57tQAWszM7wWvaO7Az+2RoTO2HKe9gNC4im5dHyawKJymNLA
5JPPPWk5lcRW+9vMZuTAc7ZInLtreMzOXqU0yb5OsKTP61fJ/Uy4RJBFwOWD/8ZB
0CSCMiXr76ejUPyzdaP5Roy8WBGMmA1CI7qR8ygk47KwnSSmNf2zTgU+dlyTt24H
6FaoxlTSm8xy1nHLCuOMJYD1xdJfnnBYgPAgcgkOlCshMDJjEZgwBbFUgANey6gX
liLGnZHrD4q1QhYok2wLOXERXDHM0CsMpZN59nqwNA3g7m9KKSzY3Nzq851BezP/
t2USPDBTjgRwOXWifNHODPy6JjoIC21UJtVseJnWvg3kfNQvI166qC/VUs0xFbzN
kXYTxaBaHRmh0iZ8xsshybBfCyRbXRA4mYOiKPDjHc+rVlAoZld7jM+zYpXJEyBE
xHMkNI2u4GPSsHGxSMVyKKj0AIkvXP6qFMWvkI5HEnkjHh26WjRDwFrw0pj8QSOs
dVxDeWFN9XLbWkFooDJS5IEVshZpPfzYRxsL/Z3opiYjMT+Anp9VO/e91QbZwOLr
qSOTIijXVTmk2wh0kBfYzo+T2BTBOlSBHIBE4yaGPK/B056CjiuBbim60oKap99B
wK3Mgr5zLJLaLrMeq8SfVlnx6++FVS+6vVM1vppNdznVlKJLGOxZkn+NBU9SiNdx
JbJJYhqunWeb+UNEmINe//+/V4hwIMfByJDIPw2zF3Jqo6Qboqy2T+8ozGjAcxhC
CXNXC/G5eTw6b3tqQZEJR73+oTIOjTtZb6Lqjpr2nu17M+pa1YJ5MFbUru7lWpqo
6kWokJ7janx6Qv2pIBPHvHRiWikY/Ky8Sm/1S1X7bAIyE5CbQbj5c72n8fPdbuXJ
FtCk40qp7DhrPk071CjqnHIrv9fmAar5RvS5Tw9Q99j2atjabg9qvkKUM2zYBaIb
1K57uT1hKyTnBPlfw/n23+fwYQ6xtJnRVYOyZ43YFMtKUquRMTfWybPShwDLeGEC
tPaPCqRkr7j/z0Fct6NdBsPtoMfHWOee9V+9fkHdrwMxfhePDYDUBeuB/lL7WPhM
8A/yWhFxVB5XZrUnmERlxz4kSILEF7y3hvrr87BAkK9qaLULjNsE8oeAcXvG/MiV
DUsLdYwHGz2ajEEj7HtG3/pJg6m+9jfWHGAa+6K2O1+GW2c1nXYAegcXvMfd1OAo
V7S9XuPufGDlkAk8kDpsnYRnsM9mlsZKG+s8I+/FA+zXI+OdLHdj7v9cJlks56mx
Mcz3D9jrDTBwh2z1oNqHUF3Ki3vHPscRaVGQ0den3Clw365gMffgaYvABGIkb4XM
Cv5ADlxJNYQBa8WHrDKgVc+P9TpFhFFJNpz6LbAj6sYwvw+BzdxVOUjfThZduku0
7FoPjAWFpB3jxmElUO0iA8PgWkGIPQ2D9zWuuenKllon+H5JbI9TCJE/f5smVuZB
e2SXwxvir3ZI1WdsQCV92ERJx8UHY5lmFSkmDI1PqeAlq04/1DWnQR29Ln3wYJOT
VxuWyewFrLnSGN5BkCnlI1pZCrlVOKjMz1YuYhclSyagw5D2bKhO2gA25U/nNSiR
5FIo1ZFFheM174xLXd6uKkLYZwF95CEyO+0GYItPjJqL8hPHRpAK6gB5qWhk1eBQ
ncmIaTtj99ejmCDBEsDGI30kVeehJgB/lk4MQTqJ0Vmal/+whtjI7bB6OYF+cZn8
qldGBSYua4j7NNBc6HZlVSY7tyKtcsKtNnh4jQJ1jDN4E+HjeShXaLCDWPlevynh
afXC/nNLXcEq+JmIUvU+19z++cJzagDDhnD9kSilPS+U9R8CDE6JQzaBMly5swoJ
0Ec7CjHQl5GIHEiHq/eJgVHKHoV/fZIDCGyKXOyPozjEd9u7nl+gGy3vy4SzPBlL
k5zCQ27RWONF8fKccqcLFuJGdelKGRUlRhHtsbdHe45W8Vn1S6OsKKinoqULZcWE
pomx6O1pRX6PSmYJe0XwMxgLVZ5vYUIrCgni37lJIBzk9CVukiJthDKn5dwgy6Fz
w3HCd/Yf/Lw1a9qNbKIwHA+uY/gi+mTlZHFfo5dlPVsyoRfeaPYiReEGSI+Gk1pW
aahLN9lt8Bk8o5scPCOoqrJb2yNZKQs4I2YY8rG/9wHTQUNEMEv0J0m9k39madYy
kRYwGEyUVSC2DOcDx25wnwtL/INaK5BR2JAhH9aZx8AjqomjLj5f3lOQyGV5o5Ep
yewk2+OW/Ab/u2jNKQirNnt8Qq/XVkdjv5l/ytjthGExuRV1k13+8sD61YrrCabk
atk/nU/XaCp6TxhFlxqRztRJtIGPn0e4pBmQpl9o7KKqg2LJ4lIbKQNEg20Hezs+
j5duAJ1tRQ5hKqtIMj0A0VM6vHbZYUM8msjDEq+E5PTKkEZNc9n/lliII+0QfGyZ
UnNPXgM7Erj5XeebU6qzi2O4YTalOKOn8IfpTYcO1VdzU/oZTrsDEChG2+Z4sVkG
YTOO61thnLz/QU29zmFmYt077jcLVe/1YZNhvDAfnG8ftuoxXACKtxZauPJYD8Ih
825X/cwrWugiCVpmh3xPgcdYsYg1pXz5qAUGdfxSu8RZs7cdJZd4seFrSQQyoCZu
WkPuWN0U/nV1YXgaGfasVdsAwHecyIHAuovMBGi86Ulpqh1bAWo3dzqHcRA81R6C
x7Mm8kraQaWxRoPCzS4sD0jOXzoosyrj00MZksJ1+YvCmMcs4WARARGMT7TEW2gO
EtIa25wbEEVQYuKKpDScV6NS6c7kKa3iFTZDcsZ05jnJY/dv2bckgE9o9G+0Oa7G
qeG/mekvHx7ofOe+XRqQfCi4Jgdc4chsfyO64+JJPUN7/HnpU0VnWy6uR85gEc/O
QwQBRmxLnLFvQ1MjWtHCunVFqHkdztCOAnJB11MmhLXN8rUB6k2FC0PoZfVCpCum
BP35xDWNhnvqFvV3kREjLapnxP2LKtHRI4RXpca/nN2hZcBsgG2mtxeBVFzoUq/e
Wfk5cuSoWm1ieFuqxbsVe1lYAOwQFNuQZ+7oJVpodbXDE01TjE5R/Bcs75JD0FEe
5kOegx8bp5wrk6VvqIUEsHJoeR9T7QT4X+QV9Y4bTf3q1BySNjeLAZDqZO7m3IkG
MvT7lRi9bvMSytMq8Xkx36RsCkESfZ+aVkQ9aqVjyFKop6DoIyW5yQDo2DeLHw1X
wTw5d0W9Ema/u8/ZNDEtTSnORfBQ9tKnqZZ/9IN7+pih/rl7UXok3EAbB2eJlUoJ
zMZ2VcTTUJzRJ4c0cKpusSkTBFJRUKR/igFgrmKu0Y6OVO9tjyfXQWGz1ZnSJoys
GyrpZdJ6YHRb3W0lD8BA11Ev0zmcJLebgt+EGIl/qcwNyhuzsBsPfWTQYzhJ0Q46
9eRqyq4wZr/jZ96KHDxreLeaHWhgj8fUcfu+n+vA608a5zbfkp8XYSjSy0YQjC0o
i12D4w1XXWOVMOTjpTMFFYi91VMplnyAyjUtxOi+taClQwdNnYrt2tY+wD4FTNve
o3lY5GxH3SpN1M8ZskIocZO3pA/kevCs/EiOdz/Gmz+hdyMbK1lVVjSelMQoZwRi
RLCb870e53wzaMD5EodZUOydnS0/a05pMSrWrr5at5fkvxcRVOblwoDV5nryy1bo
HwE9K310v3Q4YXBigGp9TMjmxzxArzVaYqTwfcz0uebzwGaZLmknNv8j4i02mUXZ
QQD3KXpM4tjy9twmcRb02i1mLBw2/Ffe4aShxxU2z9oH1a1NZnaRfCmHuBL4ju1r
+CkDH1cuYiJIXKvyOnnZkO7BBRyoikJpMXJkMHmBTVId8nUJiW1SOwBDCOmO2jT/
qQ5GY1h9FHNKd9f8n+mBltHg8ifK2QBEWJQjHYGI3fazJXMMQkXYi33gaQOexCUh
3EjAh0r4iRKx/H5k75b5CRbRfJHwW0NSNK+StsZyl/TaSOlspjHPkNtrkQiBVtFT
6aOlMPidtql9oIIUYyCqD/5cSPftOlayk8pbHn/5UFjQTBBtfcQp2OAEG+gb3Ype
dopQZPsigmdOiPVFan3HTrGo7oSc4YUQJm/B0jMqWzGIbsuioe9s0lj0o0n2Ei9m
4jJyE4gHARo3NmiuSbr782iAQbFV5ec8gqIsZGDOfE2naixDMCc7V2ajBJZWp+jz
nk8jiKnFEvCXBRi6Gq/EqL0g/kn5XGHwcTaCGFPdAm/TZIkptDOlU9jZY4mVyLwj
vtXOG5eEY2lTPYInOWqGNA68EOj/Vr3W2JvcG73p3TVha6sFJitNv0ibd182DAXY
Fe/AITEwMZ7xQwgF8slHpvPB9N2RZ5FK//50gGTmNnLj+Kmwl6g+9Y46zaQ5S+bH
NXDVVjL2z1m/3TLrroP6DF8ZNs40mVYuZeDm9pYJH1YH8rxa1bBQKnlSVl3qP7uT
vz0Pn7S0D62EE9ihemBGvxRfEM7BEWd9dpek0fs6Xmcjo8vBiNPiz86JVGeJ9dlU
iBVcUVL/opYkWwyRp9MK6SIoqZ9S9Z1Fnb4INCjNP8qY45RJ6RU/ZdtwHTGz11HD
tFFtsGMLrZvcITEq2FixJKGfud/7nrqetmt0LXxdz4/HcJ3GHkZGOBJuGPDaxDZv
Gzio8MFrLm7uJh2d4QXTbx0HllmwtHCu/usVdV+qb6gZwlZzhmJBUsHF3WRGnyYl
0PmnUEKAAVtd3CxGzmkaGFlqaI/QfWBHTK9hffFyjSbJhXQM51wWhdWMhXUTk0I9
+0kP051iBZXIERIOtWM/+s/FCQ4JH8ZoMuabVJ0ydkCDK9E5eun2XZ+07288vkWf
iSNf82Vzggh6JUcfKIWMrFDfsH6qJBZkEQs3SX0R+DfJF1UGNxJWeeqqDm8gjj9A
4anEENNExHy01GXefak2qhyzRLmDM5w8MjtNbNVLC/3GVw+eLD1S7JvT+TZvE+md
2Hi1S8lHve+gMTBIrLPK7c6jGoZR/76CiItx1RK4uTeQeRUEJAkyybQ9xA0AbRb8
na+7sIOe7D9CDZP0H/cR9AUrAb5rRybwbM6iuKtSoedTFtR4GPWCB9YNV23w6kPT
HjvlJcjaUsJmWYvSFMzpSlYk1bMLs0z0cVZHZTiRNH80BQR33gwH3bCNZMdAP2Kk
YiS3gQ0XOkA0FTLfvD8Neoh+TSTHsk9LvjeIOIqNnuXN4JigJn5DfsSdgpJ6JZbx
yGBCATQr50QbaqKsOHvg7DE6oqoPA3a0W7wiACvs+Q2NjHSF6cuCX2O5g8KixCAE
79aIiQz7x8oyJ1Yl/O12I9tXs4Bc/fWdqacEnVh9+uJkdePZ+Ey2F+yOAQwYyxXR
rI6PrLO1SP281n9iawuXeNCXfm7FezILNETFHgm4qBIR981vyWomso5iHIPM00CW
/M/41qj+9eWuGBYMDsQejRLbUznVqa6l1Is1noew4f6ecZXlmHCweil4iKZjunWh
WPRdpey1YGVAyB+AYN63/sJXnf1MYg8oVLu5gDMWcrzxOS1OtvYVam+1sSKkm2Jt
c5suCuyXO/N8NOiHlbJ1Lh5pIZygSDKxYi4QuO3Ra63bt3p+HqmwrPp79l0lrJzn
OUU3UvVvBMs1FF5pEM7MsobQ0T0s213z7IbQ5nU9OBBWdcnHOQEhysGR/X+FZ7r4
sY63AE1AqQb01K7IYlE6XqVUSBwq2SRvkRJibnyTnhqjJM9mxnZsvo/Yedf06QTp
Fr9SKPPMCAYKtH8hTdHfWS2EZRsE8c6AG4qxYRck4slCHd+eIQ8sSk/RWp2tP5WN
EhKBvdc3NlQfeQX/ZXXPFHWzwcirWWKmVKj0NsqYxdMJuo1ewmpZu5IaXQ68Q6N5
3SfzRvuE5MY0nhfKwPqtvNN7Cso+WVILpmSxpQ0h6JiO3miSlACoxxRcZ/Es+YRt
vO04KOVCSidDN+D4pIEdjLK0RgTlOtmzVzypJTGLDkB2gL4E2d/8FwOGG2IZqr/Y
YE0lL9xmTQmOiKZl/3oLqW10wr4TAjcyli29nDzIod145KTcLafVKMUo63BhM14F
YJyQ76dnTsBylnRd3gCVGqI+GP8waZwKGlp6Aa79WqQfxPBEv4eT1hgWCts3ZMJl
m28kgnj3AyP9iZXOXEObBwGaNHTjXz3LnFLhPIS1KLIMsUSKg0iOmQrQ0KrPsRcd
O9yKeWqBpjt9cvIM9Edl2P9Gh+Gcqllw5PlR/MHGRfkUL2q5Db5VFdszhjUj9IvX
shitd5cTTanOWJ2EUQcTGJg/ttcdR0yaNzzJ8/e/nRXUuZk3hoooqkiMIRtfnlZd
Waubqk8Xym1JLimt+8V2bpwIlPQDbFINVR+dJlFYQdlUyuuPwFUyDxkMjO1NAqkf
kuC4JLcKN7vj9xN+D16eQPARHQslo+f8k4YNiAWgtQoEc6nyYWkQOP5GY60+7Ckx
GRkTXycXjfvwCZOimlijklL4tuoWwGHgKC9iTu9L+2GKwlBNqfAqoDIFxeq6ALbT
0IwIqB+SodLDCHI3yv8CnUi+s6dK2cbIu9hj6mCJCjt2KRrPFjWHY04m428jh4OF
wodA2nt8nafTrWU9Qsjxe9OQ8AlcLnrEowv7cdmKpUe8DYUj5yRJrSSMlxflOpas
cSfMTJ6HaJyU8Un+sZeACB0wbi/cbfn0S534+JDlz4alXa2G8LxKZtCna8hNF8To
kgwU5JUITkai2r6SqcynfP7BGGKr55jEDmUE4tcXJaMARIlFkXy7YrxjFqQ2fG7Q
f6q3ktYEj5bATWbZsrTNcb6Cv0PUrYeTFGe7aFfsczmNw8Wctv3QbmAFM39TmW4N
roWX4EE5lIrHp2EMIr11c599PsQy5dKIBCOrk4l+kB8bkFCutDQSxIhlxxvtKRLP
SBPFxVV7IuNQ6jelRbEGYLGIUP6Wv+pT+Yc/hobxeeaJG4550SEHgx+vrDch7GBR
MBAKa9kf//uS2DZWRJpYB4fVRoXfIv0x4lZc+L3Q+AKFZsPbInNR2mac6S79DNhG
9+QUpOduEVGe3xMbJh447A1dGetTf9/muiZop9g1JseBee6lie/Ktud/SpkGcHGm
WF7imXmEegwIWWpFTTaxR3IwHqol8HoxpCrhzKu8GVrO1wXZNxXilRlefD3i+PK8
W2K1kOyGPxTj0LQFuaXDXvAjR36mNnk9JXcZftGxy6P169F1Zgn08vl6u9eDj8Uc
KsibX9iWWWodc+x3d+hLkACfjMmkDmbRdJoKo/QzsIT9ooEuWrRoXWRnCfwmscG+
f2Uq9bkoOzMcJELplt6nBhPUX5MmGZmGg1EzK2JVzZUVSnJuR8fqP95eetUGsfCt
onCcFzHhDOg19CdGErglsEvIsCzV1VA8HMncK8VQLEBeLr6gs5zN8HGgqAvfIJdU
A7M78Ppvbos8VMXrv5KJgE+tuA/HofhYlmX9gn/vhS3L9rhWyMYNCod2G81Trxax
wztPYrVAFmHGfDImLXfAUhDWUBjewScuH4DDXTcZc+iRU8vcAwMATWgUl7Ey4olM
KF1Lbto0WNOlM6QVDG5wpuBwfkG71TWppelSIcGTs64cbX1+amRwufcjR3MQdFiO
zlA/KqUXojhmTuQh41RgzPC3NO17gKnTr5ASX1gorBy2LdQn6lG5+Tbdm27BIsrh
8wOL/g6A8O+Bli6/HYdWBZsoy8cTtXsFxqwosb+zzXZOL5mSxEWcfDubILOc8Vb5
s4R6Ejs/yNuy8O3uxGfxpLA2x8sHZOoDNdrQN/4r3cL6rzZ2bsjlIw8xpK93YWV+
KQXVVRIFfVlDOKN8MgPt5+3YrkFb/sl1CR8Xn7TPen5TsDfsMfbjDJdzPAcqlwAc
1JhzRGD+P5gWpNnNurl1dIME+lpXVL3gW8qnm0u2QQvGkC9Qla0/NUOp174xbs6X
wknfo7a1WmkUBZSGmBNnh6OhC9VKDkNKmEK/lGi5aG5hPS+2aXfn5OAvfpgLqnP2
TDi23+0cfT/hS3bLpBi8lKn0Gdv5ezrVI5zej1az3SQTUcf2P/oEHebcXsexdYAu
PyorCWdkwEIOyYletmhr/abPaVGUGFLhZu90lv1+Qvj3XC/ftmwcR8gMymYR/Two
l07rCoOFpyaEOACCGQn8lHH4yBkiEdGP2djl6xk+ly9Pe51ItpFbz1JBRxW7t2Gw
yNNydWkU3M3v92IpPOc2UoHQbJu4QZnSmteUlxdYuO4Ogd7a1w165LZOGfGoQaYJ
xR3mLUFqP6ELBz47LEPNBx0hnszJxIHHwcgvrHLTZjZh85lHlrVIBAYMuE/GeTh9
AaLs2WXo8HAHGhEEIdo3xflRnlOSfqdiJVtOUMfgYsU+g4efCJ/5Q8A0XkHFw83v
YaChzJXEh/JnF6eSwM6co41VWm6jBRlVSUu0C4egQcc3J9xeYLzC4dnciYmPwR0f
qws2mNTIfLEXN8S4XXr7RE9JpnWBqQbYgatufeVKlTkclXKFzBEDq2w8nFua/9iD
ckplOq6BNJ+FTI3eS9dKWrW6P4Fl+UaOWkmZxv58/ERVzGkrXAfhR+SoMt2BP9ST
6JP11S1dTxf0ffDfAvE9axvCUch4m0Zzr5/pXyPdpvZodXMi6A9f5fnzVVjY3Gpr
lDNs43U8vqCj/TgH8DqdM9fu4oj05VMXsMrs8OdvxEV+nm2CVKUbx3DX/PO3zGN1
+kyOFne0MuVgEdj/fewTZUVRAPMhI+vzz6MDYVcXgms8p8ZyzxdjVzWWWXita3EV
9W1Xgn9kImP4wA0bbUH3Qhabg5YlJO0T5Mbq1JRI0BKnU5eTPgWGvKJ9/CQTHa9e
bSldFXm/c8wxB5LAMt+mu+eoW4qarqGWHsAYTYINyzSiglbFRHteWC+xPNzqfbk8
LypuFi2vf1W6Q0HXeVDLAVcYS0VyW26Ij1tpFQkHn6jznsJBum6J92aX2nlFM71g
5FVvGGigx2ohLdhRipX8uOS6okmCxiOfJAXKb8HpFH+K69gve68IKPOHhKQE0VEp
lfPANJm19CdLvAI3+3CgbkRZzYqwgfiTpePhF9zfa35zObQ7y2hnZscGvC/BPzYl
kOcjbpkPgjIUWgZZLLwOOwzAqK3ktN392CSz95NOWQjZZu7NOf7GP8IkQDLiHSGw
64NBZ2DFlcy2YDZ0iAWpzhf1fUdBFxmZckOgb7RN9ZzBF6K9VIa0trL/s2+LEcHA
xntdkgsQnNMF3yOI6jwlsAzArM1Ong4GNAtxQjFEJEB06c13rpCcnmS/7zAoOq6q
RKAq2G0QafHrNmRt53iNhQ5qVXSgay8BjkMKmgkyIT2zBFIGb9eUOewYunHjVEN1
NDlvQjOLongublWYRWkM9vMRAmdvo7dOlhb6ZlsQa0JAdwlfxeL9mTerte4dE6FN
h+7rRuL5l9DR4y9WoT7YTcUu4SxkMv6z+1rGeFP3Bxa47jKHm5BN8gkPA3DtSs6+
ue1ynKDrp+l105ugN/NJxGEsnq/hpstgOuybD5qQI9fMl6eDZvavx9suGlC59Iwo
rgVZKA8jr8EyElnkQCIiJHAvAzA6o/2cfVVcbDd3BRB7fZ+iPSSiWwE9AUWTwnYD
hOMVSOYoqbXHBNjWOCTLNmwStmH4cy7btUsVGSbNu83Qx71LlktdUiDCj3MelVvX
6KKcZOOAvGMRvRfoxb9K42YWQgjkOLo+/MMSS84HglB7pGr8ibRulVZWrkq/al0K
PyOX2pBD+v257RlLwTRo4xXUD8+y3fubc/QlGvFlOhf1mwiRb9XYObXV6Gmr+dUf
M53RaJO44dUVqLTNXAG7RxLR6XNwn/Y5fvoZwowWkm0ItlY3nvPAEqDZT69YQq7R
gDX/V2ticJbsFrmY4rbUHzwuYETrtk8dYjDUCMjgQPSn6wv1HVBMZj1qrReRrRU7
5xa6JxfSvoo5FBBD8NkQzkYyywH1Ssuow3JRG7xhtA6xN+Rxg5pTZ/E/KrIoULLm
q/7uJ1ZOwbiVNS1Lq6F8JEieFDXd7+nniNVERdSuPvTAQJ0vCXOEes0Qw4bCAlsZ
HW9lYACM/9M6kmGR1WAK4zEXIa/f36tIiGnFgkLf9UhyAHicXIll45l2v5y4CVVo
CJS6g+rRSbVYs/OLI73jk3joAI6LFIZVqn/pwtivNZnd/24Pi+2oLTkgzNQP5JIW
90ULUVAPWAHhUNYCmNm9ScCCoo77weBO7W9YTNsmcl/YwHz2S7IFFU1+oYBQ+4eb
5Hh/xUWHYZtjp8DbxL9kWo1xQUzrSgVsMW5yKW608LjFvV6t/+IfcJ3bXKyqSK9P
FwfTEfb0OWCNf3VylbvneFg9BrapWCh1fa6yBlXdBPRXj9NAyRaOHM5N4/ZNe5P6
dIZQ1UDss8H68HXzFLExQTm+bLUB4Jm/z/eExKbQmKHHE3z8v3FobiexVfgey2Lg
/zDTTGZscHS3fCio8H4L5nQNU037goWyDfnPFqdRI6fejounlIl9kstu6AN8AHLb
MAaIHrfqfX9g2bMnM1TH2Ptd3nmRyGgplBHcUx2mGPeANkNaqM2KwAvxCjDhhB81
DYmPW82JW4MX8fI6g0hYSfxwfZanSQRoI/sRP85/2b+7VTZmD0v84dPxUPfAf9vO
7JexdcNHs+9Y7UCbkyew5nK/OH9JlBa1IwDsMf/Euo35BW2CeaT/qFUcmDUJztRt
eJqDfLKM2RxriZCKJYo6mtvYJT4BPS8bUsJameNcqyaV+N5v3rfeQhn5mAvVDS3p
2s9MpYE9W18wb90E1aAsT6E3KcwB2rJM8D+I4iQYM3a+2cD1CPsUQ2aYieRjY44t
sDOAGOV6yq03a1jIKdjYEv5Y7MOPADdgCatU9tfdtep0rva2xslj4WXJYb2k0QH0
VqemS3ej7wi8BYVRv+kaieW+vKSFghC/M24pYbwKrb5pVUQ7b4NNFEMFJebMXUKe
cCZYgh81Ih5Bl39o7jymhsip35SLLVD0m83YM1XDahhkR6dhFR/ajbUqRpFTjd0U
iiHyb/Pg2baD7OP675+8dtwfSf1HQTWMJPoL45H1aL1/xPTZL18A+fkaSK6gEPnJ
xigYWuqfnKr6M9iGzAX/MiOc0S+duqurPKOuEm+UXqvyo+gJmAae/77HX5PcX76A
O9SaNvz1FklNs7d74RUnGVJKqXnwwlpm8Irlv9uhxIwMPiGA+eTyXcg4JYxbw8q8
wEd3oRFqKfrc3kGjWu4WprKt3OIHtLSjyP0l1DCLyxGA2yr0u/5sNMhto7V64ShG
xhgeVLRLePYrG9V/vwjaPxwGNCjv7ZiryHfvTgXMLyVfYgLFsSGYx5zJdPpFL42T
qZ+Qt0S912TBfO40RkOTbr3/g+vKz/bZM1KoFOB9LiwpPzFMfB8Nw1sYFmUCx9Ec
37F1tlt+dUmmIEVYdbRAWq0gsRBO2HEDpQGA2DRGCP/2xVTmpyRwKuKL2JLyICnD
z6hmhOjEg6sJ6a2BgmIMP9xwEM6MXOHzRX8g9W4UKReZHfs4WCqHcy4J84axFILg
usP2P9y4kjkdqFTQMdI3p76YLiV3x5QrsFOLYrFG2qKgPxz3Py0Z1z7hWQCKIuj4
trj45eF7ecAUR1+NWJ3dEWC3sgD0HAzd61P+djzVirTae0sYZd0EuA24rIMAM296
diuE+Ya6aIYbXVb1/aKBFANOChXdTxMB9fv54dycwJ9naMCcULTnZFwAA2CcGCsp
+8peQkg1tZk0ZFUtV1iCIqoYLUt9/lHoYPgH5Q1Irdxaxcm+MeO+9YOxizFdCT40
ehG7dBaRT/RvNgKH0jZmRvRuzW+lc2tteyUq4HfhzekAh73NnPfnX5X94N5mJWHH
Sp5gSsi2KvmzJE1b/Yt3ff7coE0rydc5AXr9kuFoJs4bM9HcdZegSlvlRYojhtDJ
Ce1rWfiYHlmaz+QED5nYeDx2pj8AYTrZ5O0doB6eB0uR4kkmd9w6jxfj8TSiItwN
DRJWoqmWejRNQ6RdLVOTsYhkNMQ665W0DWkBmfAZ1QR6l3BFGj8cw9pXp5g/7JQO
xduFZUCP4q1ysapVvhPV8S8WIeUetQE3S+6OYqQn7+KOaRyj2k4QzaCnf+KBn8Ht
Bg191QNelRcQ0nabnrLSdIFrOe1DUnHvyE+czeYIlRjS9gaifWzytzgb2Ic4Tt1G
4Khl8570Po/SBaFcyd+NBWfpmOpner66JwZHQXBpfIKeGFJYtkiMlaAttk2hY+Wi
DTKBTW+qcx9czwIRfE+GsGpbP1ZrbGOnoKNXgGWHjyF9Ab2iQtvpbUHMcEJlNpLC
z3/ztwwelEpRKCyGBdIks1owb+nwpCy5amKc/HlCbng2TfWjTurj7NZ/WJZ5J8Ii
K0U1c1mN+ZmjEbgxFIdRV9viSToCh/7RTYzXjRhC43vPrrvVtxUgEHzD36e1fInU
d0JSSiDxahPOjo5rzPlx8FopPRTUhCVPRcd4dMGTVWp5zof2ZqESghIZXM/sI4pB
or4RRbGmS2vTE8HME2IzH4IlZJNfB6R4p3OWh5+uSqilHdtOlpB8HtBomOjiPgRj
Ei8spLqUuQQYKQRLplpCt0on1vy6mupam647ZTxLy+l6JzhV38XblRdJxGpUwPMT
TS9d0eFmgQp8D9etO82pAtnk3saWoRVh4x6vscRfBX8sE602YjpqnP2+iB0vJEYX
oX5bNoshX5+rlcwOCgD8EvIFmLHef9EyviX8nyE0iRptYd4HnWZXqGqr9ErA2isK
6MsSqWmTbUMAAiZ+5ojBUya1nm+hMYND+3Os+HL5bA49CObLfjnyFV0DnjeJTh2B
e385BLwS7nMdaynWcjKg4rCre2xBc08dbvycvPGNx3OabyG/zPKGyQDLE6+48Pqs
CEaTaqnFuoWvQ7aSHIqBVUCYOi9oHqFl+ruKp/FKRoEFLuwzelL0ItXfBQpgurY7
skc3Z+18I3xM3+jtJEz7VtCPvS3XdxkWcDauK4IiEY6OSYAKAbFPieag1aCj4rke
HuxYsolrTeOOmF+/X57nW+aD6cFZkvsg6w4OFBrpfD4hzjczprBh3kTTSLCSHUXH
sh4wXOOCKTuUwb2JYB+a1CmGYNy+nl+BeTMhf94xeZwnPh3L+Bxv5HbWVe8mwgH8
CDqo50hEhNtSRZNnpLsAT3axm+K2AbRYk4Aj4G8ng/IlqkL/PvySvUQ2F53riOOn
jcBcBBiCE1jX5TvcO+C76bzYWodtT5BdpIu3wzYWjPg6N8zRVtTlLiFCS3HGFJYJ
BlA8RvZ6x5h0ubPBPQwIWCcAmmvWbxFkbk7VWkk+VuhFZMbmYgq96c3niNtX1zCe
u5WRxkmqYf5LRvbeLWZbjQitIhUSbpEDawyHbBOZiFe+d0shaFTk5URH+V73RHTq
pDLbqJ/bQFY+0AF7ojue+m4v/M3ZbDJ2IZraE+dMYtWRmiqZoZCIZWiP47ypVsc4
WV3UF0ShN4jEsRQm6OEXxoq1ScbSwOZItqkSyMXkXjgOHjXBI26cZonmuQlWOaxf
EwlzSoUObZwCuwhGODoJlTzDy+ELid2ms+RzQf9UMXCTZuXzF0vhhNMT6vahR0xT
sKof6rPw3dszbwru9U2BXN9cB/KlybCR6HGjSWq+cn/82wN52Y+quJNOTbZwaPya
wD/cOhz0KemKJ+WbvhP6OSdhE5EkO1sY83RGzsEUdZc4TFKcKkmb9uKfIOW067WU
x+5rSQjYKiHvwp4DqpbsHmiNcCnIHboBXyOn/QwMGWeCvtY3cgRgqZVZZGcBGOgj
ILJ/I9Ish0CnAxSqyhn57nuaWttbFWYt8Zgww6g97ToKk3Od5GxHjUU7I6gsuBvS
3SXZf+UOshDvabsKa+ffzPO4NShlxOXDlnxIuVXC4gRUzXSeDhRiZn4g/bFojhY0
/g9svQ79p+0ThYFKQ1Mf50++voa6xQYleuW1gpJKJYVyk3dFs+xrfypESNkx+ko2
rj1ULndNph808ozS//IzQ/xQwZ6bI4+sC97d0/sR8HRXsiJMtfUKSNCL0J1aWpUe
1er21zPzqVijFxPpknXFxW4PkpzG69kBBG6nB1+je8GfuRBe7e6z+mq25lM1pxo4
El7doNTaFBLw7nDrAlbJ9qiaHFJHkupfo8znBYAOz5CyI6PcOTgSiypGBDTrChB3
DM+efl4vJ7Kjq4pYEuBvCQusNBF+PvHiB3k9I3ZK3zr9iyiF6diW+0jb/SVUXcpc
TGE7FprcH4fE5j4RtoGUurIbhkMGI5ynXXqXeL/BxANU8hXFATrAb5UlJR1QduXo
/hiBqv1hgWzDQ44jVvI9pNRwbVdVL4K6lf5g4ysnIlWHRfYhUigj6I+MkYG8YYyA
tCkUj9BTd06j6Sb5cvRZqEv+6RBfOniob3e9OOmagHA3BL/f4BXcjLmt82D4bIZ8
lS/DDfIG2Gs6BV1Idi5n4aQxb2XvK3FfgPRLf7Tp8RnPTbYU+qxfBmg9uJSt4KoO
Bpgasb3k3bcRJ8bjdFXPgKGh4HYpmzzF2xwdvT9CG18Otq34+YNNmtwXmSaNbRiW
RKgQFsBeFpY2R80ZAF/iA1tbMnkKml11esI5CaqLuJvhzymrcXI0JDMi2AfV/Urs
KKlnjuG6wIkLu0Y8/S9YeFG7ApAdBu9W5yN/EDs9419gj5erURWJAdTPXQJkgfT1
uycthZql+eDffqFotgAPJdgLPEZr3ge4CzgaomHWR5ukPhL00qu0qd61ebPENZl/
e0MXYSnE3qBS84OPKfb/rjVU6m/CYdRtS2TgmjX58cnbRPQeQfGHtqvDB9Yydxld
FsqBWhwZWrDiJZo+vHzf+C2EXk+DaXsWyF2GG+bjaz2xMvHjZbsCxNHIdd05Uh8+
gF/yPFdJddkWm76WQbl+fQO3JlD0NNX9ZkF36wPWPCsVmPqvtrSwMGsB5ovWfrgv
zGFOuapmQWIuuIZg8D/ch/zH4nbKR60F2UeBBY2LkQaUtPq22qkXFwXm4ZDv6t0h
QqutERZT7sQJ4dG1v3D/I9rzVTrt55Nb8sS+lvYsaofU9RuBUxeRR46k1jdv57L3
B9XN/V7KKuz0diF9pZ6xGN41RUc92hAqQB/CINoU2ub+F2nC1pzBzI3viO6waowa
AiDFlSo4S3xcMIAZuh0tENov0LSJMR5EN8JZIvJM0zBlKtrBFTJeLOAVdmybfTYZ
ddZ9mPU5w0YIxHXwRpch+I/apTYsABsClwbGAS2SIbZUNvjxJEj99AzdKyDE9u6Q
V/3a6e8gXYfhYHbDzenk30EbrDijYJmvRXdrLJkmXfGG8QhhZoJDe3xmiyTW+kgT
enWWtljb5kOWJGKBf3lNDbF9IAjhcAd6tGlhpnAm2PH1jybvQ5/rJUphRV/Zl/ph
76OTm/qZrcs3hxsSS3FAA0lXNiatfqp/bNO3i3r4R2k6Zej72VJfrLShgKETxL2d
ij04Zl2EaVzt+vv9fPtX8/WrO8XqRPFfjiXCViMtAhwGfQ0MyHwPOmJSLlvW9LEB
xp98fh+ZgQEDl25DiwOHmhUrzZjt8jW20qLkFroBVGkJ67GYNGd81J6t/7HGOshk
HnFOedJdYgq7GJvJ9U03QJ4SxTLyWuJQeCE//n7kbTsMtTnlvH4WtK7slyz/SCeb
ocwEQ7ooZ4mAWE/1uY1ezLSWfXfMEtcPnUFSPUuu8sh1VZpuUsRRE0iXEzIWd3pW
QQ7EC+7XLPUDv2/nWLLbCzhxkza9z85OT1fuan8WMTJ8KWHVwk+1te1Exa6v9Xb8
NS0IGZaPJkIJZvsJwG85vkKMj6aT/ZZy38kxNmvnYRkUvEhqEuz/3M8zZCk235lZ
CuF+U9NRCVaP91/RNt91sPIYPyY2n1hBH2NZ97gwcX0aDFJ7RpQBabDTT2eeSVqK
JMVuoewXGf7KtkMW7cc7nEFrXwO6JaaaPs/F5waWqKkEzTkoHv19CpPDE27CHIsp
Tf2m1+E8RKZwIDOIx5hMlvio9GHb/9eJSxTT3EB+X+opLazlnSBXapvSxIoliOe8
n67I6XeWy7V7Y7jm6hDsASbBpQfnGFknKfGTfW/WqSWIp9l7BN/Xt4puCjIi8lYj
NTOt2vDP6Ket2rbmmguUZtaJH8MaGZYJ8us662glnTADWIvWezVUHxP0pe3MDdje
HVbHH8FmglNw07+DCaihxxc/GCLrmYYqCj69mG7M2h2gnxt5J4ZMr3ebEsy5N1HW
nMiNJuCHxZeH+R5ZJI7DjCFdm7OJaRzPXfeAJKxSNXSicLm3exK7sty4iwBOjq0Z
4Akn1F658t45GGbszl7XineILkstUYRHLWevBqdvb6C2FtC8B8IxuPT+i2jlU9P/
+rl9n8y2IcNHOERStfO/TM6ARtv7KvkQPRExEoDoASB79ljBI2FwkHgUkvqwiy4S
8oRKf5drtrtlz0ohGZlXEdGUEc6YKz086SOxySrScnKDbf0bu/LCLw7FU/8B3gnq
1aiGG8D4Z8zkTQ/Tz3l43Y9j37QI0poNhohO+fwERHOFiBjaU1ADrAJKtBhg0ntR
uVSHn4NsNAyPDSJXI8Goz6786Cg3Q5wts9QpzD9Ju8GofHGIavtorzua75fK/Y+3
uowWKFB4h0FF0bDX8Cg/7LeFt8YCV5p+jPWZPTokjT1DQbaKgadGW9rAWs2jPCnW
o6HIuTJ2ju/qr+cBJ3RQqUQAnCiDKia94DiFC1Ldk6uPX5vrUMHKx56C7Bq6tyfV
ZR9vxgRYRm4n2Ahta/i7uGxCEXMzFsEQOhY/0o54SkZhpk72wmvE/0mGbiFaiC8e
wS8yGIIfs+w8QifSGwX639Irsr4wmlEviJuncOwtctYmi+MI8f/ccS1hLeDrC7GB
us6CNGngLjhIPjJ5yJayQ2I9QwGODSoc7y+5kGThOYB4lZmLl5LT0Z2jFt5waouk
zAZ0hn1VfqV6GKJXIKJwNQq9xVtm9q/3lv/vWi9Qv8SVtSRe+DmYPtJ/sx1+ZYEA
mNcbOeVsh1ZQmrLbeNc8unOJ61em98/JU0pSo6AbO+HuaBl19h4O2WczvFbFj/Ig
mRvSy1W27sANld5eaKtJFO59liMgyanP1H06TnDNhQw03w6uq2bld/rIuYOO0pxm
0iPkeXmRc/UA/93JDFeilVN5re0F1sjPrxAUloVBeReGOrpJUQGvHYdofmoY1gSv
EnK9rvWQJyaMUFj7HaoA2GZfhRaK1ArkvpqdI9xjdWAKIO7hD5sf3PlYd8FTLx6p
Y66PXTKUuFi/HlN6G0Fs6JBvhxI6p2rjmxtq+I5ZpIwnKJ9mD14PFm7ZEUiDlR6P
1JodJIk3VyODVhHmi5ITuJ71LR9hXpCPniD9GWxNPILdK1KmqT6uyL8nhcHrs4wt
sktjX2jiEdC+D1mqNpO+XrdqQIbPxxrN0n0eDKBFUQ/DqvlxVyIjD46pivZdcvcf
bsySGqyhWjKgvqEmeuZWAk0BR/SqeXje7jhuMs3Bu577iEnRP7kEEvD3GNNLk614
Jqfu6he4jjOeCdT7yF7n8ZqllttmUqDcAG3gk89vZSUF8PWhrgfRIU+ASDaNOsMA
IB9yc5Qo6xSkf3KTeyBDjT/2mKGXyXUkVMoyuY8jr/240QzJQ6BcsY9+b5QWNNep
djdCBVuOREX1ZymQJxQNlPjif2iz4eRI+Xm9WfhCb/H+4/59ldt/sTJgudGx7rIf
PjzsHTo9GE3DGRcqr7q5P7G42o7QKjAkn191zjoeUAgF9rmKcYw9zqZE20NiDPO/
u7OfGOu8UOga7e4O6uOLeWwqulDCwIowaqTL46NAPWorRi1mdPDT5Tw5bJhImhnb
JEawpT8iUsyAoMtvJV9C06zvCKVzHLJ90gaRl3tRMtwEJmMIUHo8P6Zo3suvL1tb
fMNKEKkhKvEC9PpUUpOAAhWjPUcWVGq5ZWSVDn3Tj2wOEylkb9ICwgqCDPFAxG9S
AX31vJghhfSdAVLu6k3PfNfgqanKRsus1Gkw1kMv9xVJc5UwpxVfbOeX4sTMKmIj
5TQiZMr6DE9lAviXSIe7974kUR1Okg7W0g4Av4hAotaBpmnJsQXRUdIuef0CPPGu
uMqxEjCPrNDpF/LsWWrUNfgdkOMFeooP7cINQJbXVKEA6i+UOGJP/WhReQYPrRau
RYdrvuaCaCaSQjvH7+l7SMz3CHnrT4P0Z46iXlItodnm5e6Pz2P/XcY29Uwu9/jx
XfIpsfGOlgikcWDyF2RpyZFr6PXuwvfmUjDDLfoxz80SyD/7/RATYFbGfdmv5a0i
1joPpHinCqjyY4NiSizz1Rx3wvuMvfWsV+lqwJDHEd/tDjLhwpHmzxHd8gtz7JP5
a140ztkYKHgmbskArHulp7J79PLrRgiUWad5ymM5k3N0YIxPanUvUSyB1BFpisSo
VSTqrlPCG/ibkJNflRB//08psnpFMFtr2p0Hx3wRpgsen0DJmc8OBUrmpJIwttH1
eBAammqPbRFIEyNGoLE0zjBEIcRV5QDB3jaHVyZxdGR61e165wFh93Sp/TBUXLAU
BZjnUpJUnF/mNnDv5ubBrvsArg37PC9H2iNxR1Wc2H9LXH+moYrzsSTPTinSXyL3
RPRndBWo5LRR4eFXP9cRvOLkGM6UXq9I4p4EEWnf65jzcxqkE3HB7k7mt8dJBmE9
uQHrDv1aqxUVSseQCR5/g5C5vCR5Yhshv7qky+RxsuL+uP7tvZPFpzD02d3rRGEs
BYa5cJo+Bzz7U6SCEW8jDWj/21E3ZIIz0hi6hB9embyAHer6P26aJvl1tA6MczfS
vm/H1B+q0x9bnDPSkea8K7PBGhqZgDIIoTbERtnSldEgoqIcZ3r+m6v51n+jJ2lV
ZMj+VSCcq7Gk4tXzbTwWRfPYvud78ZU5iTz+8/wpgTo7ev0VYgGokj/+L8SoyAWa
kGRX7rIMICuit3yNEt99BmwM/aVeiQkGT6/ry767Bpez1ule6j6thdU7PgyvPmqn
9Iv2Gc/hPZISwDr6ZR4sHvXbjIQ4ML1fF3k3bB9lS8GwshDfOl/dXwDZqjAHqZAp
Q50oHO2tgsbHUNg6XyvpqSckCUYHR7g3rH2Lv83v9W8V/Mvt2ZI3vD9cmEkSbKNs
ejVag1LTVgz6nCm/1PKhSFMNjureJ/9nx0yOV5kMaZnF1RB+aUG+BU0do0pDNR07
wpIJhW0fbylqFsYgFBNBiGUFyjZe2cyGAUo1co6mqBNZdkvqLLwI579MPzJWG0xI
EAqxt7icCmWaepyX2r9zrDg6zPmEM6zrvKXn87irMSVkKeoXIanOGYNy4qa07CPn
Nv3dF1YsADZWXEoZrh0p4IANfQQuliKMLIYzlcxgki18lrAm6qSFS0lsea67j2EL
fbVXPlpAk3byol4a9x3fIydRuTVohu8TAZZslTvgvr5Zh8m97+QG7CPL0RKA0tGO
OEtFhk8MRQCf4By3aAevRiUDZeB1igr7cwWXyFPiCRNDnChFJmUpHUCtWZ74T9mN
KTzqQ2sfapDHRxVmhp/Qm9G+5zGtGGHUigUDHP0zbozf597CyEijNhxtWbh2/2v5
ZB24SDVTJkwqy/CmnEvmeyncapZE0sKE4qKJhGnPE9TSjhTbmpwt/TPthx4X6y5s
Gjzy7NUAezYpeRhZgDybU31eUdjupVrKIYukf91EA3ilYFVTQXxw3IDOvdJJ7qvN
913Ir/pKqN68ikfU7fszOyCf/TsUzE79nQojX4S+We+335nU8fqlkM708P4GcDh4
sS7KkFGjpOmy+nf08HZqGpxbfNA1M1AkKfiQWSQQFih/Iha6nzMfqwCz8JwuSCd2
NwaWkcZJNCyd3NaFqdMh145yR3mpxvAuxKwcbbc88BmeNpR5Q/GGh97QyCGht4dg
l8krO4QGsCsJR1+OP+Q7l0nxSGOMh1+iKWKj9LWVP70m35WTQjQfSX5DA87GOaGS
hJbi7bwFyyYkiaiXZrqV4uxQo4es1GbA58X1kvRf4djrGInlZULZGnAvybRdsour
b04rqjyPU9f+AbzUSBJy9v6crygR7MZm8wbPDRx9uzcKWc6tsmhJ9YRLQm5i9BL4
ih+f0CNqf0dDJdzOSzJeIYNmy0pTrha32tnq29AnABLyK5/soyC81DtH/LiqXS8b
YVfUnI79xd9gYR1zKhCQDdEGENc2d/ozKp6dZoK5Jwgn2f4KWVxXAyuyJbsn+yrL
BT0qBqTrFoIJdWMYElNdGtVKd8Xb8iVuSFo8n90JjmoNVITF9I8+mR2tqZbml2qQ
AjYdSxjPf9I2Eezmx9y9i+UsJ/q1lUq/TGY4Lp0yH4O6PQuE74Iw8Vf+B5y2uNxu
iLsknlilcDNr8JmCxoLUg1Q1Jfnv+e5R3eveyQ+ckR1V+jdgHhYked8HmNByJZK8
uevgI6qM5LJCcwzoY9svKJWHBy6Q8rqjOlPY3saChbtrkqwtjY8+Iy/y7XLNvlVJ
221cwy8vdoBQsxRdUeUwO4NKIdT/iACUc0I1uTffRhMPokU/dCifl3FvSRJ4jbte
+z5XHp09c5T6JYmsfvq2yHTUIw50m1ahFIXVBp4s+r2bO/vG2OlzyZJM88w2ozUb
mX9jgj3eP57uK31VKOmk853g9JZa4gGxUUXMa/7PiUedzKfI2u4QOe7urPZs6Kkf
6Cz/B0rDtpzRk9HY8P/2wWgGoxgA+yaAvI/m7wvX6Zqu9EoT/Egq9KhkWKyVpXDG
Tmhqy005nRjBr8PSWlEEgukahuwRjfK0lL3btFwMrURdrpDTMHHG8QcuPwxx03JZ
/ILcf+TDSQRuULJ+R4wrbY6sKw2KD9Rh9LlCtwRZm18ogQA7ByXNc9pCDExBU0VN
IhJRGWEZ7U6wnVMPJNiSoVNLL98lb6diT6W21I3MZKAu8l6072TbsbSWfFJyKo8x
+M7JsdjKsCennCHBHzbOKC3tSvK0zpLEeoPgy76iuTKO1viKDFoWTPs4DYMIkINZ
OJpBVUtB57CNlRmckZMZhdeHvLL3eUB7lSAphnQaiCY5Z5Fypmmz1UZYgLWLXjzm
L8c8qvUp1JjT6mJvAUEam4DR2xcf8ado2aWCupR6XQjbrmMxA9tS3C4+dX9UpgSY
2R/IzUfH39MYKc4fYDep5aOiGImGLcjvORqwXQc9h65V/JtfwmPs9h8v0vs1QOyh
vYXt+b5A6hzae4O5b5z1Rrf3cIzwpUd3mRA8Wx2angNkvL9BElt6hmpB3KIeU+de
ZniTLX7HqkL/HpdfOg+iaB26OzLodgI6Vu1DBUBQn/aMHh/a9gE4ATBtL9ZqxZ4T
CE6DMq5x3fgvCRQZ5M9TouGOTqNmMCRsvitc3Jjrd7WN9BMKXPkz3zhWO5i4fGdS
XMx5pvQXT0Uo35KWAAj/406pA4DCsopFiFlr8j5BZpdiUxEAIs/oSzfMyZvi+UzM
WR0v6n3Iu7+OfFfOA3ZhG31hceAwrdwEqejiTOVjCWEn3uLrXxniEJpz5dRLoYtM
Tky/Qz9ItTyyYS+e34v9qpWL6stcStuOPKOYe4fvefunUJdBy6WSGm4+HSYSCdtQ
Pd6m1WRUAOL6OLFG8yhsSu7bYtVyzFPtQ2lPbcrptEFIfP14G+SYTJQwPJpNGt9a
QG2TOfKWZHVepphoxDWiFr5Ie+d+Tsfrnt7yONQX5/yq5zMZdhk7gHXhYd8FEPU9
UmYK8rbAwUi+esJpyVbY4GXIqu0+zm0zOk4E9vy2rovTDEQ22mesrrxK3dVtU3Hv
TkZEwdYPxSZm0YguM4GPREVHfVmHbwEHjQ11zNQb8Yard77+xjWDd8Au8NFBTikE
kL0lzzhvIgnQEf2LdR50fotcMjVd4TLjhNWSwrzn94VhclHSSte/RZXBAbMAVgV1
I71xzzO7eWfuaB22sr9c+zisb+NvUGZdtS3TEpoWlY1ikRzJHCZm+rJAYw9ByK7Z
cKJc+IyLFUF+So8W1WGak7IOf4fmX5IEMQegC1ltkCM9edh+Asv9OIwFEPSOhrAM
BHjdS0lwwMl6vdIAs3s6zGEdkfhvkMLn9PFlSzHV8JRudEL3UQnn5lcMxw9cnqRP
A9u0LeO0Z5qQwKb8JSWwkjcIUDL4hmARF4bxXsmNIByE6oimvAyjp5x+e8e9rGKr
3CPXuwOvB+w0oAKAAmFA8Xdk91hOmiOQMIiqxdiqueNDlPfjjnm6mmJz/iFWWLqB
yzuYW+z2+tF1fLf5V/Ef50Pl7gv15MWLQRGFItSC6IcfDCfVo6HD1qrQjeyShEyS
DS3JKBc918cgCqseygAjVLh99SPjROeqg8c53N1pDsGqKSd7i1Z25S36iPKGT5W/
D0J8u8qMXLVVhfW4g7x0cMZtw3y4GiTLFjZuhaKBxHie3jkUhCPZdAMvP8ExRMBi
sNu+ozpQb8+J5vyt2VG8u7+9uoMms5WI45sg1YdUBhxg3ncz4ndGHTE9S78AH+GM
435laRyiRXrhriILc18C7IF1Q0UXkCh8akfH6uUbLAHSSqdFneLJ+4LCeshLPhTC
xBri/UvHhw1/c8fKjjKyC6qlymSVD/HVQYu3lBpKHAqkPpoY3otqITIuXY/bqkaN
odPCOX+J/djXLCdWY4vY/QwlTf8hio1KG48qru0Sv6M5Uhi6PGgEXgxWWe3uJlAJ
IJokUzZCJ4qpKUMmmffMAtBK7xT4KTN+4VPAAjGFGRJdNjc4o6AiJyke6pmqYr2A
syhg3mR+07PWg5PCjNsLZNrvdaoNlEwBjzg3Nk+lOPgFxoGMXcLceDFkxcxVPNoA
Xa9PiZ/6K8/WQDLxR2zxnMIjmPArdxsMyv5Ds3PiPmiBIRfRGgiGUucQp5+f0m0h
/Ybw7vAurRpgxmwOpgFTpeb2ifkz2budPiDqr9DEGaIoZUQMhxBZcJ8h4yMmv5l7
ndWgt5+PL2DbvoPPvKaJX/ccmhQr1bkhvzXAw5xyxW7Ol3Jh7dxYhysdSU1lSb+8
fHrCKIlcKcizszEstp6jyWKZTimREe8wE1mb2/RwKIVK0gKg1o28tKyKY5uRZoXn
Ii52ZTUN4ABbJEPDZtIQ6zwcrCt47CASutR81qeaFrXUuM7BEgSwhKxHrbfGqDrz
oGjPH9W+ZQI/pNfpY1ntWvrtrPu+ZadMpb1SbL/4PXsHDkY45wnBy4NYAoeoDkOg
eVsllonrJ5A81gDIJEnHEutFxGGpB2MR3pDWa2B4gy3OrvSkULwK4EumL7ZghjMX
yjd8szbgDRrv4zgKJOSp7+olIHOigmvauNfKbvwjN3gHgG/mGVnA4qmY2W8io4a9
0SNIPXnukL+OQi+hjsKJH70/ljfG2cB/m1QDYkkyXJ+AD7CTD6ok2BghFPOPY6kd
IsOV5wguoYEzdZEmJEoYVwz5Hnz8tLKTpAR4H6xOfX5ohwG2zDVw4wDpa4pDvRl+
3cKAYSqXDn9mR+XTjf5mGbhkmw9YKx7SvZWIIDuujjoM95mtZF8Al0IEZSxeQUwU
+3ZnaXaGueUCMeF7Z4XfooyKki697uqmTWhZHXzBMfu4fSAVzsxTS353cCZVrcg2
E23S/Xwishf5vKqaAbOvPdal5pUbuF+P8ax4sy+JwNGMmFJTBwPegARBXXUlzRxB
H0FfpYbhc6CDIDuG8n2P/YKoo91pBHPbojmIwnDhbLU64HrVwx9q7hANGq9jD49L
Q9n7PYi/QLcjyoby7jgFtySqNipnz1XiYdZZsrRSxX1zm/V9vGNrEv+6sNjKsCG7
5NxnQGShedtuozcsB4u2Loa036cxY2qKJ1KtD6ZGKpiAmD/3TqtQSRS6KwvLmTmO
gtz5dv8zM+G5pziXdLU5UES70TafTH4gHytPpF/mxCdFBYvhYtm+JwhDhS6RGFw+
/XBm+ZacKxRbP34ZTx0nl4WUhAk+32h8Hr/WRUjX2960aSBA+W5jqZB5ICKQ3zRQ
67M8DIXwtdmivzwSL/2AJ7m2wQWqsyVQ32hedDcaLWhTfNa4RS99GuDNpDR3HcJy
Oy0Pcy3lwKVZbbrRi8yxU5S460bzMSbay8r12ZL4mrqztsY/tXKN5O3m0WRRgZAG
x8mK97soItl71cKXOvwv2nP0h+N6AWa1jpb4W9ddADqINuVH/u6l18+SXv0akUjX
NLRA6Mw8WmNOPZCGYkaIT+e1HV3GkOACzF+pNJrF8TzywC3XESPqPnlaMJDOYfBd
Ei0XJ+ywhwFeKdJsSum/we3E9S5McHdiAyQAJbXrtTX+vlWG29LLOHXO2N8StgNZ
8KJE1op12mf4OxjHq2bdLI3mgYdRQ3usV6nQAgMVwSDmQDXriaGB2lf2zOezQCf7
76lmd/R92szRoXWBoCtI7KNmrNXLS+AD6yjQmE8alShaqCFAjt58UuDX7VQbbQms
jh8VTO3jwCIGrP4+xac9YaoZOw6jDlhSr3TX05ohTanVV7FNbco+RCinGkSfWG6S
idPwxmXnAGn+kpb4YmKs1CfBk1rQngoKsm6yG3hxMY/tw1R+jfkpMN2mymQrqdUQ
vJCGhAKC8wGep3sKsMUPkSyfrL9es+r6YEOgafMxzKfY3qbYDO3oWWDZpXpiSWiK
2f7ahlIzP3CH1UZv1z27mbggOB47eOGrv419E5ypLweUlVfme1++OSxmqC73AOcU
W7B8kvADy4SPCHiHkNaGLSYfYwfE8Yw+g24b5SFb4nCLk2xTjzHJ+yiKdXrKLNs1
yv7TIx2JHuZjnRVTakk43tu1QjoO+320Wf3qzLZ1CE6M1KvpspUGagHfFLrkTjsZ
Cwil6Xk4gjfTDyE0EjYByGFzoBJLQAyGs+HzRsDwF3J6sCwcB2/jYh09Z+53F0ye
85Tyy+ztWo0JVNGL6M0cFBCprjJHdtyoksnO2whqCk+pbh92EHhXojoERhAltBpM
9rBOf2Dh40w+jGruIeZiRbuMEsKnwRxkeQMok3TzaVMp18SgiVlislELUF+qt9Qk
XWxZbJ5jFGBxzBMrDKwvwrbIcgfRiu8rnbJZqVukoegp/sN7K3frtu8Z+11N251S
4OEkHPkuV2hVT3eWirAgn42gfpkwb/yPuGRnFM6RCr3b0Q7v+AY7z3NZ+Gz9bKxX
1cVdWoS4cYOV3ypBeyL31ZIQf4U1r/VTFhwXXNHyYEqq36ouHNiQIeNm5dUe0gI0
Nb/IYVooKUqJ1a6pN9Qd4XmSQtSUGIcrsGdkmXL1OwR02OkE4uxmhgrI8TCqgjzf
aN5/knOcd/FQhGdl/QKznj/UjdFE8Dbm9cEZiEw3n0artmI9Rtw7m8xVawtFpq32
fd4+tgfP8PXfbQcy4wZEoVUOsb/1/hlIAOjtLPFSoELg2YkQCuxKvvNG4pDz6c6P
PgMeJkvCBVfKWXMBI5cuzCg5L2HTClEQcteCKXsB0Fc0E8yEwxlEBdn43hypxDKM
dkbnp6FSMCTQ3XJldyWp8CDZtwkMTHxNlZDWfv7utkyVQ1ToLvHeKZz5KuWWnc2+
C50RG37aEkPRKD4pYgS0lwDtTvBlN0b+pq9KCBLor+hZ2BZRLwgLtk0oGppRK4Gp
1o3yiqXuCcfgZ6gKrwhd3ZSxdLnmSmzINNmiyl6rNBFrUhnhP2rdJI0WKp5HnvdI
+cDVsFpSHVEqMUciY6xDdpBdaJfCsP32WvHTewp5fdkAsKnktNxujEHA3j40Um/T
MJfLEkxq6gDGOxGSluO/iBNIQfthNExUJgbBBuxVIN3eErfzfDOKVFwdj89SJgXn
nUEFFKFNqIHsg4hw/U79PQncVUqzVyHTYYQ5P4FnyaVzhS92123rKoBAS0e/cJ0H
ja6bVevevjW4d8srZW7dlgX3N3jAkfXnMm17db648GoXK/lg8aD9YIBloy0LrTZk
9irNEmAk3l4vP7XkKKKlCfqB3E7Y2L7MqLameh1DzI9tcOIJbmX7chp4S42tT1IY
b3UWWA4jSG7kwKqnXsmIo67Hm7Jf4TfDYU8ukiGfBlXmgIiaHoTNLgPQLKOypnl0
TcbEYeGFG2S+LKgStI9S55uThmqRgo0+N3UEzpyiZmun0js3w8iTVute2QOoQrQR
VVO9ubW5NsueSGV/knS4MFAx8OlQLl3YsoGK+PVYoIwLiU4+cBh71aRybBQfQrQm
mRDyyNkEHuqm1iOvTXaulQn4T5tjRaE98hfzfHOP7tizlPq+rnSoGC23IuQ3kQlh
cw3WzgSzuWjbSb1Ry02H8EW5JseNB9UTM/F7BMKutbVqR892cXAr0iIcGCmiUBoE
1JkakzTgNaGRkgBQps+/eZ2DbojXvAVJzwyowqeDh8R7VFGztkzlK58sdQS2/cxE
vecZH+kCKOU8NLiEkAA6zEZIhKEjrLAAx3+vcb7x1ioyR4Bk1D0VGJv3vrI6DBbm
17PCKCwu8qAP18bxnlYmG98F3rtfgu0eKM8RTRnbZoEcwONrZRt08qzCsJFGRSRm
Ad7Blh97jcLBaCyAoFSUKQmIHtxgKiLLRgTc/JAPx181QQOADWYSxQxIooBgQdA4
5Qtt7z+9ObBjXobxGAGcGWPL5DUG4w3v4c+Q4kSH3hKZ/Ke0bIBx6srSsaPd4vfK
yVzhJTqgT/MVsIxOKFIomfuZIXIbj/sOHzOq5DEtTMGtG18BC4sYLbAaqxELd835
o/ObA7T3fpQ3XFHh8+8RjErSJVDuNptpR/6tJQuliZOZhO6GB8ksl+35zV+OfYvI
k/clSK4TVn4cMhhshSOZ5wHMBW5fFcn8ZozANvI0QU5+OFof/ljcZZp2uBajwHDd
UH5XwGunYVTA80rvYmTRyy4mpc/wyr5ZE12sUWmTpUloBFz3HIORJjU5MS3sGdoE
SHzYtlkumqAZZ5YOIT2S0kmBUedi+Z7W/40NqclhZtSJgZgGsh1aChvJ+3as/OYy
lDhIAh7frPnMMXDjkgZvkh89ccSwxfAzaZ7Hp9siNRnXoSZ0UxM/Cbwab77PSXkN
p8InZx2f+l5CVXfQu59CMCW94Qe0I+QcHx49f3BRyzcu94YxeOl5/LMaNz/AJ3yn
w7zzvLqEQHwQQQHTWXB2A44pBosOt56CtaQ1EJeExGrNsiC7ykd+rH2JoHJlWLQf
X7/DdXFB0zFbQU53CMaqY7ljlerlZs+lG00/V2qG3xL8y2c2Na8vJTM9g5QtROsA
xjgAdsVx0euqDD7BbirCw9mG/mVTo1KcUlHhuna1YW+rRhXFh/oYe1rE+noT5qWE
AutufUySRIW/8fb47JIFI3w/+UF4jOTPm1da4R7Ln2Q5BC4XE6KU3AvtJzdn9+nc
em5TL49igFUF3CsjHyIX3JmDZojPU5m7VDeLaFExlGghszdfCp0dnMiKqPwB9RSt
ECBA/zPH8dX5ZEnPD1qxFHMhSENdFbdx0/nNunDiQkjoiO1M/SJN2DrtfJpNimQu
6z2BrVpZqzSA/JWrOFlgFGPfWeWx7GKFB6FRnnUZFLCMIhWHRfL0N3eRLinO8hWL
9ePVI4kJwn92+V7UfcdyjHbRPNQZ8zA3ytuIQyM6QjYuXcEktpa9dIrnwIHwvgca
sNKvsuWdCJWpBYltU3mCueI+HPuj5tuLs3+ZkeQDg4/z+Q0gHH4Hk+Q9oGe+S9BY
m38FSXw7jey/cartWztsclnFO3Knw6coig5XAcpQ2T8HI0Y+jsZ52lhxiwvaNYqo
+rq5l2f9Dr6Ke8mp/9t+QQMEAurWeuLJ08Dd1Idl2s0ilBJ7JLMYN1zrbqj3rYMe
hP23TpGaP5cPoIF8Ej+DxE4O/3NlG+IMaC9PVDIgGAKLMTQ+8HWuSji/J6o5qRqD
pQMb+sBeXucSjD5AwT8maPfww+1kqWsV2+pSrx1GSj4RlQzABzkSYny4wnJKMSeR
Fkgdp9UE0TqfAhuwHeYKygtSh9cKjxvGMYPtVw+7vGiM/7ZupRb26Ug1ecUuJNzj
PaIpIEXQM1GfLIgOZy8Mb5uVe6zFAIqe6/zYQ+M5QfymaVEwRQcY4u4W46QLuD2x
UOfkN/YgsWWziu81POpa1w6fuHUhyrTZdwbmCR6AdsnkGhq4td1H01cH5MZ1St6S
zS0XzuKAJUzHC1S41VuW7ExwM7ko5Dv/uiUj+zfmQUNfA9htFkPpQacimEx6M626
KbkQgrQtBAD/bxYSkkozXea00hRry1iSVSd2QDYhe5VNuXiaoGF8lqW75bJezLPQ
cLQj6cqUvt+MBV5dAxw8F0XnENNlsJOWYAt9FfkMfbDvAcCe2X9io6LPWAKbO0iZ
7T27l0KFNM7TlgU6+ORx53c2t2P1quvGaGhuexXvWcFcvmKd08EFx9oFMtbUZDqj
kcpwJYbeDN38TAWNf5hDVN0FlItBXAb2W6p2CZXwSJaDmYqL5xsU5D2jTJGvqiZu
zZzgoN5+6gXZ8uofHqtlViQewD8K8x7QyQKHUJTYvfjMStMY/Ielt2vcl0IjfkgW
t6qthHGs5Ngs+CyxKuwwA9fXSpSXg8vakzRQTIBlbVWso2kHwgJQdYP83KwjQEWP
BYkn8abj+lYFROGcuokBPfQIrMfbbILsfs1bM+z4ttAqPVCKTYKSeEnHaUFPnlBU
6hDABHJSU8stXry716Cc7XLBUQhQoqVw1yGrpXqxXHXrUwPfKSCRQRhYpJ/qCyUD
D6LeNUBZgK2zkDtaR736Na3dA5McEkTobAhtPu89dMH4/xR1G/XIY4ZraQBIYTLR
6uh0GNGTCf5xrYgsKf1hCXFY9JJA8l8zuZXwAyN/cixDCLGWYp8NM4NUb7twCocR
jM/kpAPE+fifOi5jqb0jtlrzPQZKsB80BiNc/p++TIwAd/Q5D3ktKAmINOjFC+SF
8HTxCPhvI2KRVnfNbyEflojhnwSOGoVEbWb6aPjFjEF5r6geh58K+so/STPmzlVZ
MnjdJDdn53KFXlH4x9EXsM1wRYq34CMuceCVrMUQ4M6ayRAnuuj9AKOsQEwN9SYG
svR5C/qQK3q8M3RXWR1JYynjvr16dC8EJrHWo4Ps22fLJED75NUNVKSi/AhEE0cL
9WSdy1Kt8BiziYPqT6nizw/noKaaiNqS28UFEQADLa1Gy84uWUazbmNX5n6QHA29
m/e0Z9TQJLYFpriCqonwz7m5sbD2NcECkYUlF6VeIpPa4Mkto1wZjLFL5yWb5Plz
lweWSrzoYlVTfYFdSt9SrpYywsj8PWCpXnScHo4ElLJlYUt8XeA1k3H4Xw5Go1Zx
l7Dxy/WfEwIAGOl4kKSDFGTUNcpgtTX2LAgJMRRb1/2v9viG/U+kOjNf2d7GYuCu
r7yB7MULpoepP75wZpN+kru21N1avuBBW2KoFjfsDm0igV/dwlAECpIVoV3++apL
5LkXcodVMn7dTLE/6Z14pXALbQDSzsAYmFifiYFx0Ke9SBaIsgxyq4FTVhSktdiw
B2KkMLLYgCw3FGvujtnWi5C894LsOa0ViLV0N7TUqrMSEl1PawOZ3OrXZVQGXBVh
QZ1nf2H69AEPXtdxv+mAMXbzPal6xUPjbkMoLk/cNDT6jdbHN/4ZQE+2Lk/xWzSP
16gsDunMsSXulNV/vGpJ+Sv/8wKLt6DI8rMAJG+0SV3EBkjJk86wsABuydr20i3Y
lqop54ygZo7WGdDr/et7E9zTjBmUv1fM27dDwlkcpL8kNg//VjMSYppyDGyh8MYS
F8SyF4DZQWJteuSYpJg7CJjpa8i762NO/hLeEV4X1LStVBWo16jmeQigifBw1HFH
dqsD5E8o6GOhTkavmQ9/rJOdCpU77SiUe8ED47ro8WKEbzWkaspkh8NTiXP7IhKX
T2W3NysOFYqUmPxsHisNNhQaqpjTGIMrbHQ2jUpNw0cEufsZ905pze4yIQ1eaT1B
r1CHnkCFlFNo7Y/H/S4qVsUfQ9m+f1GrwMvRkUqtOY9rqk9KX5w92LHPrcTBQ2WA
RzSe2PYEKW4k/e4DhLoKFueHV1zhXX3wGyHAZHwTSo8v/BlSohxJQ5DvwUqehx3s
lylV6tTz2JEIuO+Ku5WoxBqMCzGnUk+hB65jc+9XNaMx7DhC/DyMwBtxxHaK5KW5
cb0cn+WF4x81tad5L/1rbWEgxyrDBcnSJFiTTtjbZk6XuzwW8GP3fZ64UgDgq7Ug
psw12NNxtHGpMy97gXr4NALvV1nRaWzuNUg0oAkqokqfj1vl925lhj7/ddys9o93
whAARzYvTa5krkFEVvDkwtY48/SQblSaFfhYFePd8tNIZxaHKk8km9WcasZadZER
3bnzZqspXThntx1MqG1yhmhhkEyXsdzDkexeaXTvQHsYvga9xtUeeLwGjEsgSdcC
H7hRp2+nI8mAU/SPuxLVmF9mUWVFRfBjQuJSXr8W+sLSFFwD4doBJOerYO8lSRvM
XqRn6778T61c71QdSAaSOKJA1Dby3LW1sTyJGqRyIeN7NuAHB8WXMKKLknJd3bEJ
JWkUI2V5+eDTy0wzFaFniSl4NYQbzXDbfIklXWVoAxn08SH/A3W1fJWiFf6keZCR
fEQhmEx6An80lRpHZ5PDYb9If8wDdMCnIjxBoCgQnrUcF2GYJqyPacikILPN4N4v
NN/KOpX+niRGxR5OpE5VgfjJadgDjO+/iVXe5Ianv/Tu099GdYiNIfPR5eH3roOQ
fGolfXygJ8pyWIRQdXFgoeFkV/a82/ogf2iKW3SeQPdFfvlnEdDFJum2iiGaJU+3
AXJ416+JC8m39D9YkkTLn8GkZiI+MLE1FpVS9DtjinoZlzfQsP/vnVWutnxz9FVV
4bozErvR8K/zmFwcChgj91Tfmlbvm+zwu6VpArFgjt972D23rjEsedMdZMZRTdgb
i2O4l5CD1F8w40JKhlU7hRAoUp4OY+KdNREGnzrh4gHxzej7CEC2leoalp0a0rEO
ZoE/zJTEMTYE2nAWl/N5aiNb2decFlFA+TqchOZdBG6Gvkd1OC6BvjXrWfVb5a7J
D9A7NsfWVW6Wfjxun1EZQYc558R+LmUvvqHvqUGwWadV0kdiRnqNrn8hUtbXyn6q
NIn/NI8TZVAjdd3QdMYJjV6RFJs5HDa6BkvdmUd/XIa6juKV4ZarV92qx+CSQyRM
UslFyHiFhJVQwNmCRg8cJ4xokEzeZggEzuv7PFfRtyaUihZ+O1hCd6pC1HIaxXkc
awBAkkQUnXCpl3fGnwiYgNFKHT9UkdTsyMkgez1vIYXjSBPo3R8Gp61Uv7Bbm3v7
8pWXt4sNXX9pCPgWqURx3gsb51rC/2yDNrvuXtuOsZjPmh3IPKIgEfNKSjilgkCK
A4tczvRJXUaKLbaPWzMMA/hQQ8pKBPnmMm1+n5+a9qnwtPNw0BOL7h8xREj1iqU0
oaCQHzDxE7CfLoEE8hakzI0gLOUDz+5/PtP+Lxe8ZXnXqgNYbsPyUWvpodtPvi/k
WHOB3znyWUcw//RZmfKHHYRPeNboImNPsR3QpyHwgyFFWuMKaVsZhZuseineEdHH
MpoOy+jSCK1I9mo+YeRQzrFRo3rZARw9iyZLp1C2W14cY6KzweuE5r2gly1eW9cR
cj9UKT+XcQRMrbfikN3kpFdbAmRUcl9huMz88/LNrUhHKXo/mWOzfWuFK3J2DewV
crktmAmvWtv5vHnklCTCfYesMtpwOs5pXzKfdkcpx74PO4jw/5hXpxxmXwVJqqpA
+feqpQxTFM1QZtL2KI5P1GPsZAh/2AjVqRTwmzSQ79J61h6YrE1qTtxkTTvkwJtS
huj7t49i3oTNQzWNoaO9+inrLdnYcmIdq5lgMzh0AwGDv8oHIgDT61EKZjKG5le+
G6A8OfpNQ/UaIRp12Z232vMrkWRhpcaSIR2bxFICuGOYaC7/K7XKrM2Y6dXxmKDo
4hPewQTP9+GTCjlPd2HTU42VTe28M9bnmHYGeo/OL8XWMPAS105KO8nDsHykSFid
jMb5Lu3kaA7l2i46JnA/Tyma/5dJXF+npxYCpSRzCiULE6AIOKUfccQZNYPwFUXi
5H+vffHdrhTJzc1aZipM2hu3UZfDTqJErSpF/w44/ThvGw2MeJRK7kz4UnEiLsCH
LTlekYkhpx2pvEiiRCirA1Uz35Zuoe8ghqNaXWtUMy5q6ztuLY/YmC5bPBP/qEnv
2n8arTOCF+VewmpO1cEXFsNR1OFE8lvbrgRG1GZPmCsqwpanXo6ya9inyowbT/tB
2L+MsSHwjztC9SkbqAtrhwP5UxniOStdj0uzToR98d6moIu1hNOqcNpUXOP/AG2e
VmFR4mRq9hRB6yfSDFvIPLWN/IDWzFEekegH1zS0sTroOiIYg2V2W6kYcWfVm415
8LeG3QFNd8je9uF0Me68uNlRWINP/wQoAnDXbmVBdpY5zWEOIeVv25g4k3om8rb6
b2DuFi/Zj71Tmfr4Sc3pKsPcz8mNu5JttTKy4Olc5y/PrcsFD2ZQLJ/x9aNbUnch
0s2lABgvDPCV7n2vKQjC/R12qWn+luG1qAqQXAywwerHAkkciY3SItpAsID1y4bV
n+Hng8n9YjykfinJ26Ko0i0dQEABP2hp/4CtDqrbBMsNtcnfTDZlQ0KYjCuHcxDn
5E4mlbx7eG2lZ3fxnbqc4vXmM7u9JijhVqAyFgJgO0Fk/RPuZc1fwZlwa2ZvPC73
LpSBaH5sO680moAzTflcOeJXVQ3YHbupG9spF4HKhEfEL9POYH8/pVjD3Szqqk1D
M3sFymTh/MFDAwJXfnB7a6cV293L+Fh9gyjKwNkLnz8KA0o1v1fj05nJvGHlfHO6
x4FwCXWeWcfw/l+WsAOgVycm6s+52uoirhD6JBZS5+7u+h7M86Pf3pScSiyGTBpX
ovZMdFmCpoY62WXYRz/gBFLYGrWt2RlVwTj8Pc4Nbs1tddgYl6VU7cuXsMAqWgvG
418Ij8pZl8Qi9UheU26eV7CZaLwNAZMxNwAhTwIoNwa+qc2qoklPVDwLNJATHT2f
nLYvdfU1cpw9EoT7zc+qRLc3aeutLJeo96dWqZCz7nuRtYCd0lJvcdB9OIBshsdG
uLtLAyW4tajIbCjO4xSG7Adbs/WOkJLdp69lvkKo2+T+CxHdbsH3dyguVpr5oGrR
7j9dSERod2FtpGh0rBjlTI4g/SfgXOOCKKczSEWDAdw2YPHhF4QWN3aY3uYz8GN1
8h5SuBbLQFTiT/DtVQTZERSG9QmcbOu1KQRdzhCJY6GhZHHHWL8kwTYPHrWUbnPP
JEu7S+jiZZa2epzY3ZD6Pr7JXyqaFxREkll9a1TU2bixdFK3GMnd6G9XnDuJSjQJ
IsduYov3vRZspIiGvuyFtPVice2qvJclhIT/zNhTWB677cvRDH+EZRV2+yl+9IV+
HeKDFK1US0ybky9QbFJqoHYZIpaztFOBDTF0mNVGT22lOraMvHEPjOFLQ3KPafWJ
ujWsnbMjUZBJfr2eSxJdobrVvPrJ0suFB4V3vogPtrq7oqx84wOSzLJ31oGWznre
4JLAfH2VAWl82gOjKmkoyBAiaaosU7+TmEKVT0q7Iu+WdNX4J/B53kAccTkJZ8GQ
wQ2LiWfR92BWHb3C+t+bauSauHlUYNoQGvofMOd48KcZuo4MDBHnOkxvs/e0usua
UyJC16EYURZ5PEdeTbIYOw4JgKGBuTHOTGfirjz7PG/5NocnIxXjyFvN3MBULCbm
OzKWM3H0Go3ZN5hXy77Iubmf7GDEqwu1vH4C4PDDygbbAQqfrz9kwEqm+vvP0IPG
k/xGugCKGzT9+ggrrbCcod17hmRxec8BDmhhbrMPjKGBobCBRfUGEaLfXpXwy4ER
MuFlr0wiTPem7lTscVHV3TqMyxolsP7TumEtIngjCU4BCauRwYfEjJ5erolQMVKh
2fjd6QYlgRA852w8uRps7RgNzrynrIMzzn3n7kyMEssMqjvFmWQ+JNz/i0EMA8rm
tspXU/HCj9tguVkyoHLKMp6GYKCCng/EhQPcw2JUvMJwNgq2hmLv4V18Zhlbl8gB
vKhW8dSbpOOwODiYSGOPYpiIYLBinPHUstL+6OCJYUqWQPt2gg9GywFrVr9yPY43
ltZ8fNZv33B+8IEe7SGjJ9Wmgi1f+pYhWQh7m0lx5s/OwP99O8v4B8h0pOfSfEVf
CjjyJuMYIBDi8OkjRl8RtePns+ezslZOTEkwafgBVppjGYADL1yVW80spMsN6XPY
nxyEGN46amszdjmmJrJfEywupO7jq0EED4yzeN6t9Fkazl+IkGn2hpc8373ajdS4
wqiIZpnUcRyW+MOOstQO/PSnV/B3g5dp1AnMWkfiscwxx9EBwE1Z4FeBjYmF8Dg8
ioYkRbQXoA7UQHHt3ZCd+T01yg8v4B/O73yMSMgepMKiea15FJp45UM0BkObN5r9
xbn16ZaMPbqSIdLpYAMmdrpqswrKsG0/tlbXP6v2FNzMPet9l92C3/PAWHX/Unqf
xGKkXTeWv/F4RJSADGFGPTEy7AUV6+LCE5Rz+75hPFOOS7mnVut9nNOB8/Teeuga
roTHpufJ4Ok3p0Ih2DjVsE+fX37FO0Vq20USZtquhdcl6P49zIvv76Wlz08Jlzvv
ldo6jyA9+Yws4deyexPH83n13hYO+pc4FTB3Kq4tInzN+uXTYT0V1D9ov5BZtEQs
3jdX8veSSWIWfUglLtR+4HFRn3xeuz+0DVF0rsJoi2iPKjPR6Wsn8FtLjD0j4X3o
fKbCm+jEGAPkRiiJu70+MTr5MDdmda3cYPWvF6CDQjplxzz6sTTT+QM8EQzFhofM
NWMWUD0jtFo5G0YHWs+5UO3UWhCtV78LkXEXQVHWE4VtUscBXvbaZGeaoRHFA8b3
IKNKJjs00ShBuwTHRT9XKTyhXk9KyDTiduAEB/FpryOV1FDs6VCEiej2QR/4yoJd
Njpat51udHss7Mq/0AjRH3pGGGbli53o6G9kH/KCvXnCu0JVicO3YbIh1odNzprc
rugvThTE1ysUm9YaSLIhn8PdB8jyGkd3ReBpmdjrtr/j/D5A57XJImFMtNzOR3Wi
lKxx2ZGnCX5CYSbYnpURo9bLgf2wQkX0pbIVGmRNH13OxanytMp/bcJ/hlvSP7mw
MW7ePalIq+qG2Mdj+1vPP1mR7fGROzizaIpPB2HmHayxNUvyXz3FhIdFJ5bHlpjA
yu2osfpN1X2COFYhjX67HdDve6CV9N3cF/moEmfr9uW4W1Od7hoJfOkEWczV6KUu
wuOCeD1wjj5A9KRNDvfbfzMW3GeeP6F0c8XkpUdyDcBdk0tlIkKKAMQCL0tfrrHw
YzEAmqAhUOo7a1tn3mPuPRClXbrvlzboOTaoaYhCCYHgySSdPSEFEwigCugQfvil
EiJk19+9g6AuM42ICQjSwyXV0aN2qonb3eZhBTFbIrTS1mRVRVl3G4mi68DlkSnY
ptf8A/5gx9hUCZP+WI1ceA0qnKSyKRk2m1YdOU8eGpLz6QpDrNO0OkszjkNrDZ9Z
ioW2ymiDF6n8nXKeWLblX0ZL1hSO0e+qkYM5re8s4fUaxjRGZNyfOeT6fETxsvTY
ZI0XqJZp7qddWO73IxC2G7hJcekPWFPzpB5tssUezEfdPXiMAv9wgu5FpyqI6XJz
T4Em9rsQm9yMd7mb4yCilVPiuDGITRhaocTY+qAxZ+ySQfOs7b9L6QtZ8Z5WTO6Q
eNbmOP8vsHjCC4pyOMm0xH3Wne2NIgV1iFq7yjsXqCOg27qSe0sw6HpXZQODQwdf
ccOR5j/tUGCQ8yArLkvY2A6IlHX98a51XmMAa1OQJEMxnrO2m8VNe5C6/6LBivA3
CAsbp51jZfs2pSEtf2sfx5eAx/PyX+LO5159KSY8ej7YuKWoyoXsnfC1PRW0Sn5k
2VqwlDcN8z4lk1eU98f+eljGPKlXWo29vGVFTSw3yyOUMoAUIOugfNNsJvFaqq1/
6c0W8NtdRsXyKTi9l5FD33Sg0XwNOxS4fHHnJDGg/KDQPcuTjNVC6UrWAuICBEW/
kSszHDhpTgOEFyKowOIp1s4srgpyxm/dqjUxkhIdqJca0wPprZfHOoywKQcZ5V91
GnSUdQR8pDSx6c6IMPa8yXF2QCIgZkdwRwqIf1mMbjQoolGiHSbwCW0UEnuu3lra
7/0es0dIr06UJvtDLt2Uq9tX9/fG2zG4D+oci7FNeQ9MCfzzWsmYLGKQEM++IAJ2
T/85xsuResodnM5LmdPEWNmuvGU2y0DA/PZ9QOtFobRvQ+QiOzbBxFbLlJBHM69n
TZ0zjf+/79rh5WL5Vc2rzT5sCINHIxN6nPMkCFRnYFAKP3Gl4mxEt9sJ4W8FYgh6
V5C7blT/2fYbypQ0kl9GAHTVOfD/t6BzT1hdymn1EHhjuzkQ9WF131eMaieDrRpt
t+3s1VEmN/AHs5m4jJ7E0egDMYlcM8+DpUMVYoK8jL2YUB8c9GD4sx0cbXmFjMIx
UTgb0KNfbMes1YVBJ3Hn6umArlKi/x6IBOeOSon2Vs0t2SJMPJh1c6oflsjVf8u1
ycEC8h70QacRMOekdhtXuVClXDhor6/AOSVGuYFCZ0JVCg7CRPgS+YzCAO4ffF1r
5sSAQRCx0+1TGpvLF0FQPTjLMBkgbiQ0zi3c0GtggYkrYTjRBZpfEuq7Vu3cbFRF
KEGmeAL/5GjTivLeR2oOALlyR4iWblSy9aw/6tbZbuafFBA+Jajngn0UyYUE7DcN
V9kJWQh5vDbnN65CMEHuoFsTStmT8J9dIO/ijcGGiIb6mkq9l/sgrAtqhy7zT7Zm
APANVUG6G3TGYdtgJ5VBqoXKLqwTZS9Md8aNfMcWq3nSIaMj6499sMWnwFWQXaje
38RKibq+ZWzp94K48y+er53N00EnHzgrDmG1Fmwdj3yaumHGJ1/xnMUIR4Ctrejb
k8viT/cZ5hdtQEHBNSE0gbkfYOsMmY5elhLyadC3eLWiyqr1ILT02Dmv9l8Lk+vK
Qwa73L1H87pN5DLhpqCey/JVzv5Tk1Wuk2OYLldU3qo0DEHgpeE+fiGKqadHr0Ud
W2+fqDRiPCHSoCeK2U3jQOvAVej57iZHmiYZC/sOYjR9AxiGZSuoqI1gH/C7+cpa
XZP8Y5GECgD4J4QFWuKqOnV1IsJdMZ3lDjz82XIz2nPRFuWud+alx7XcqZ8mli4w
7FSjoOO8PQv2u0T4K2WFZ6clp23KuBqgLzvzJkrp2/RzgfWlYXnHOhqgdcfyfEEb
DM3o6+Y9HxjoevXFkYnIyZfLU3thvXcAarAAPC0hhid8ZqFgh8FX0THL3gBdhItX
K5+yq2kipDH42NiLzxmC4YgM63keYnw+H93gCSP607wAoDdXkecI9kEgoSxS47Rr
/JRMwpk3jfpcy0YdjMzLjukPrZYfPW06x/1VhR8JfpEw85bMrJKN3Vy0deIQi9zc
eyTpYmIVmxBocPKXPQQZWWL16VucQmpL4WSa4B95ksXHbue0K/k1Abf4nsTxKzbU
lWKlGBzbjQQoDIwZbS54sSiZY1XD9z9WDESCSz636GNeyiTBOHgMGEwAQZR6XW1d
hIkdilMq5qhEwQ1veLu6ejhnyrp0CvacLBMZ3DlNjbIWzBmoKtX7TYLA2Yu92ctr
dCVhZ4rfAVNADhKXC4Hb5J14w5BMg2+W7KCIVW11maH8xWfajKN52FgCojtORklS
9fp+JZjDhd1+NQz61TQwIRKCV8TCgEvDZI5cDwrzJcWsdPOJN0TNbhXm43tiPiRa
0CzzC0W7xqB5zLcLAo3gPX5+/oKUO4idBFWJlDfWau88IONed9xbCFV1gZauJgGl
AoidhPQtsU6t+jf1gLE84n21m6UehiwI59MK02ejbDsUUddKO29RorhFT5Plog1G
i4XB2EEZWLJzsD8n+fpvrruTlhhBaGP3AwTZ9qNdDIHhBCAVbpPn434fEzgkq8zv
P5btYNYdTpC4jxmBbPpgQS3T6kVWPXDP+YJ74CeOfVbQmDeVWb2zBlH1zN+VMSY8
Y4u3Xu4SxVt356vBuOFNTwcpGnX5FG4Ju33HAi+NUPbqae6+w20G35LDwFWL42L2
0jF0COV+rCC64kp0Qj6sP6G+PkVxhT35u0O0F1yglKGF88NWTdDGfGNzfYJ1Xif1
W4aNGiu5Zn1rzfev0d8bx7z0Rz59OTMSHGLQNulPlXeRMQGEfQk8oZ51gcYkRmem
OGwcn93/6nwAvPqUCPqlLgEBUjM1cQY1GiuOtrKl/D9pgmkNcNgl3fTkzzGKF3iT
Vqayqid7bB3V315BBes7+yzaemowLy8uonSzB5nBr2qFa5GMEqL19f1FI0cuMoYd
cHsn5YLDGaw4saocdu2SuR6k3Y29fSwEsw84oPBcwBUBah+1oUqiOSWDgztgSQwB
I4hLtumYYc/q2mghSyo9fMlboEBmHkQnuzQ96EkfGARy4dT17EnMiSIVwfumh/1E
u/4yh+AKQSWSJeQQNfbbg40QPtTBgReFB4O1QJJOcyWMlCu726uByQ9h6f+SnPA+
6mVizWEOU/C3TvL7J3gY1AqwAHN/Dm3yA7QYA3CVtKiUxLGT61bIpl8pSab5kdDQ
68B9LNPqqBw7+EsuxI98GRBqqTfWCH+m5LF/8E0HJtrGAFnGUZ1bdSsjXxiyXRwZ
SUGDNMFH7QAs9K1ixzdTtccI5iO0yFUcv4zh94BywYxmh/SLcQJt5Kd4KxZrXBpr
utLY/EiRtP5E9/LNubXdnQZ5UiPITCY+r8BxU/2GWB3+/MtLwE6Xcus5ZIzehejN
vVJO8a2l2leFqbiSSA3kdBC6xVb69JqsY3Gf16LU8eLmrwfsWhXPpT5sngzZ7iZ9
QHl5De3I/Vds/kYqUHCdmD4K0mabF06r6GJ58nNR7+Mu43pcaST1lRl3YMOh9fGa
9qkNyZEUa75qyjPDHyT32jEKgjtVB5Q4As2bkJbIIpi3jtHIc4W4sb6wWuWpgwz+
s0vpaph4PaeRRjH4dQWD2M0J97o+LBNzYjz9VeZcwRNWjJr7xfHQnfKiFbrwSGU+
l01h+rwcU6JlQNboXDbkhbteXDDIYPoK3yTNtH9k1zANZ7thoIUn0mpjFe1gxkcl
Vy4fJMH6ZhEhJqDsWR/bYcN/a+7Cip3lpCJyG0PtpcZtExRa56bt2Z35+nSR7CqE
FPfTkMQHXhrhKFF2Zm3C3fP/7suW+N0PsDgmptLsQ5pPI2a/UQUKleTnUcIlqz4j
z4HfeTmco0ddLes9DqLy6WWOYl8YMc98XzD8fCF/S646++MLrUXEPViOF5iLfLYG
poYudwXhmrGTh9oeLF0eTS+k6jpryYGbfSm+S7PpacN/4aLeYvk51D7UFBswzUQn
bxatrRojCyxG7hza4bfDMvluHICj0JurWi5dV9dgXB2RSayeE5VM4vfGTkuSEP0u
fho/1nfAscci9n7hRqltTlWAXX3NFMZfpyCjF8LESNPyzJIi/ylNn8XDn4WGUoXo
vVDUb9iisIUttYBTQGr6yd69yO/RR61QGtWlMkPntbG0Hx/Ybl9HWavNYxLRew9b
PaMXc1YVDGAX6txVNZJktdobCVOspocrXGgDhgNzyQ0lTAfuCI2Fxbc5Xx6yvhgD
QzrnJ+colApbMl2N7l8660oz4cugPu/M9mR0oyNeCZFZUGG31lQay5B0McdiLv3Z
w8gWlh9CRBX1NW+uuY/QRyAb7zOFCD9rpIsnBE3Yoq/CsNtE+tF6eJYegaKwms/K
zd4ERzqnp2QwC5tBRJjRs4YMMvgUAy9guAiwmox871PNQ8uAXT/SGBedhhNIMfHh
LweB82Pw82eLO9By0o5iff7rCUELLQlu+XELXFR6Rp0fEbid+iNSRch/p31vTAeL
JsP1T5qb//t9NrYH7df0dVlnvJGBqbE6ys9mNqPv8/rLZ/tfUwEgJ5D7UfnROUbD
gistQcTBjCwslCAheYAAeVc1EYkKFX8BJ+dEiqNBrt/d7l1OMyyA6BX4gqItn94l
x5WWmCzRUioixqfNqg7CHlwfUhDO/oSYF/HEHlka83i6h3WcXwngOeYxCduswEtD
JgKmEO/DoRT+6dgcK5LorIbZZNdAYWiGqOzc32ShlauZ7rRqwKz8vJ+QDJ0MGlZo
P2g8CZOi7opkG+rEqWoDpUblD/3yYdJoJxEx75E5aHY9COU1wP+xwkjZwE/4i7wK
4cmDub7PGkbIsO7U42FCmwB+OL6H7CE8Cl03D3jnEjov5QpDlW+mORanUaz8nBUK
/JSOlJ15SsDTeM3+KyDU3Mn59Rt8a+2xlK+K4MkKFwIY5VuhUxbV8q10sqt0geAY
g+oLyFRLNwXUFHWhzW7ITHnBeu3Ms0TvBPLTOFn6SW5pE0+6f7OSdJn1QsKXLrEg
Kg0tNhZo+dm7c8ADaAbiWe/SvNoFOWxpflroIInSi/VY6Ms9wxWX0b35c3xFN3cI
7SAQvNMIHvqRaG/xIbjBvBMb+LotT2CXr4RtGZoLWranCfXCZPZWTDfrWgsolfLq
tb9c4R3eMs960Rjubq6WiqlVPDWs+nFl/GSZioxUSa1wsoz7ssQeOc+EufMJccuG
5PITTlIQKDHqvvwC8H7MQq1NO5G7ZQQFhGwmAoOzlYQRiavVymlYZQoeQoIh5iBL
6L+fJkslSbn7nBdomJprLaOYtJ8Rw6M9RtZ4/JckXJOcUPFekCtOP5INafx+Lber
1GbbLEfKUv4RO+B4pb244Xq44lZyVDWDFEjoqJRDAAkM9T547+rZaz8aZyLV2d0n
kHzxuyWFUaCkZK/80mdOnuAeIr+bpUwNUNTIRQ8dqpHdMWQtpI1puV8HQ9PUZXi2
Clu2M2904ryoRS1O9ERhCZmJm/rBF4/wkEkmx9x/2eEuiO+y4G+QIZN4xoUDOF0l
aEFwQFLf/v/2TRuvxcnW5262eLjsWAKkvAqhm2uNiCT9Q9RjNJ6uaz2GFeJLoSB6
8KxBQYU+rXWx03NTGDCIE8FhzUWhZOWB+88dNu+7YufjPpwWCivVAP59XiNX7RK4
jRT+K3az5a/JLH3bRFQoSZ7OhZGsJxzg8aeR06epWOjQ0DzJyZbpFNWuqVdUKfUT
+E3ztEcr6I5Z5FKqz5rHVBZMj+7aeUQd/LKKK8Q+RTfEY5YnaJE/waueEbHmTpeP
wH5ZEMVMtmUkvtw6PhaBkXtOlSCZZQP3IOKiN7GGmERrNPi0S/AidVRJAYXu+WCe
WC8ezV6hhuakEY/rj8Rq6muwqQm01Ap50RNkv482pEHTOdKTXRG/Km6qItgJAhuo
7QBHnXzUlIKcamhbfm2jaaLKb5M8ZDuD1O4ouIulAOBxMWy6ahBA62f8Cd2xTZV9
EzRbWUer+T7nzPBypo0qVyoUmtG983HxXLFlkz6Vz16EW+Hrc19Ap127Tnsl4Vo4
PZahEcqMNHAtoTiqHqFUDgUnXZSndocW8hgf5qoRmXYPrgKJ0YnAhFHnMlKUb7LV
ZzRStg0yHggdLq5t706EQsk4oeq2F20k4X2TxsZcTY99n1lhc97fasx6udLOtzUs
vcY3DuNXisPuXGt7DaY2EtSUKL+FW84i0a3EDZvazsV53P6nvbfPYMLzPRfRLUBG
75flie2k52MB1BrJkOKEkG16yrMBZnnC+3mKQvygURBlc+B9ocglqzbjENS8J99H
AeFlLIzWnTA6dtazyAvd/i2cLPkyQRZGpF/mAVV/uOvVtI1ZgofqMSDRbFe16mAh
Ue/0OEpnHJHIeMGTGjuvHV7cvj5j4XrUo6LeVD4VkWfTKXaJoWImuFNzAjjdIcnp
Whsax4tzjiQBpyk3grG5bcUzqPMcLyyLpwRTGgNezM6xzO0o9ehNQJX+HpDeJ4xX
zvN5USjJIvz91Hm1W3leZ4x3MISKx8iEgQZVjfT06masutN7esSHsi8R/FB46YO4
Adec9qGnf/y/xHpTseZKLTEUrYPDE7XIHso/1+y+BqXEOQGKKvlTV7tsTva1uOTh
NQ5ShWElU6SHDY9VoALNi1VBKibcck3pJTHVgmljlO7MlTP0xescT7ygNZnOnv4G
ko99VGfxKB0iLRB22j24uVNRmq4DTS6WS4u0cKzx64xLEr4lLym1srqU5KsR/QzF
pXglUFM2POWnIhKW9QapP1kwzv6n7gt5XXoKCXQyI8cbHt5h77om4r/x1GZxrmFq
jgvTOaVlae35FSkI67uEXJt8OGExYVHcfLkavcqSov47klXBc3ihI5o/C6RKw/3A
bija4igeJvaDV3lxa1xc6VAcxhxrZyvlxrZBaBz6eRs6mAWrpdh7DdB4VI9Unkjb
2dWIFVNdZh9imju6QxXCB9IPxJRGqD09USImKc/kDBvqhtib0XGD+9SbZJtWSj6I
SFde38tCEXCk2CuhVcpIQSHuIuv5sYhAtLGyT3hBzpc8iMvEnluGN4G2SC3Xyzif
X3O0OKqJ970qCxYR1qeXiZs+XLBwXWNODnrgfF2jeW8wMPZ6F3xGkK/PrWi/w8fj
ZYp6YokvDb4FRIF4sXZ4TNo8OIe7FaPZlByDGv6njVS3Q7M0Gfd5bn4DRzi7g+YZ
HjIP4FSgbFiZ9zc+Sx1VTaZGVlkdOt72qC6CMlSms+1TlJtv9j0yiXYhqQK68Ycu
5Iuxt1GaY2rFVTSu+IuYLHhRRcCmoBB2gDljx4HZeDzrvDQ5/1ElRFr4vZ0rut6X
IyIJgNKvZn85cf1QktMLya9SDG4EJeUQmv/Ie8YcFczOX4T73S1UHnyTGGHtSNAA
uc06O+PMb7dLAb3apRU3Spjb2zuLkbnq3UWDNIInsXYO36PYAJYERRTfxWid/wM8
Dqt/tCG8wWTP19noD/IZ3BmLYZS7ICORGDOKVimUE93M65rPXak7y8j2IDJEdfK7
++iMziHKOQzltwn5cVlTrcal0yBGEx93YOyjco0EJwJzu/Tb/QiUxbYC2n1j+RIz
eBstyIz/OFK+IfrCcRG06bz0WqgdPx8UTDZCzcW5SfpQrw9Fj6Qrcl/YF7TwczCg
02x4iWBcqyW4xbRO6iy3jATU3Bou3dvJk1mmjaYjtITyMqSjCwVciIjILcA9y1Wi
kn5fI8IirhE3iL9E96oHFuNZFUdint/Hutfc9rutSR5PrLn/08teZmXpFqLxwaSF
KP4N0Yx8FiT28frMm0jjHEYK498H09hGcy9eOr7+qegAFebz8eJn+L8upPUMqgMS
td8DLlO0seIgJ47ZScEaK7/LTAMiiuz9tN8Ijc9TTgs8B9U1W+V2VLjmg3pJ49Ya
T3OtAMwYdQ19VF8yerA3avycDOgqd2GcydvY5ucrgQAUylVhWQk9gIuyU/eO+vMB
6vQB9BbpcyUZPhQM7dmU74LZofJJ1RrLLILL+PAVwYSTsXVB3aOOVBqov4U9+MS1
wKHl1VcVSoyDwsfAWbyBZZTt9tv2yohSzD2jwj01uc+Oi7TUBsG2DEsqfVEaFcP5
eJ+5X10R0jVly/DKcZ+WS/ZNCxOYm+ZUYvcdPUjxVUqkt8cKWOC+O9Xn4bUyqL5f
ZeYa5ZDs8yX8bSTN2G40mmM7ozP2lzh9n2DVRihiqa0d3Avry9bZVnJvCRLZxk1x
QPQ3Mu2mMLJoF4CH6v8owea0+HMQ+KwNM9gvKg7VW1CkyN8fkLdsSHsNfcPOJVIN
MkNObyqzN9M+FZPsfbuP7PeFcnxOFetr7+K0ecRFWD3sRL7GhFZxUPdfD0HcBLbH
6QcwQbKUThg/vryc9Sx1UfN+wuKIDjNeReutoEDvzL2SVt4xM60iX+cMthkJa6oI
Ado9/xmQMdTcE+FPKlcPOM0qFWFQreWeXzb7cDoxZvv/rASk1Dc+xCmy/N2C6HUt
0KKAEdMIMF33P/D0Rj5glzqma5dog75lsDGRFV/nVV4VYohAbn685mrCx2227t1X
+64FB2eDihDi69JovCNjFosRrFG5DI56VyK4vZUZFmBw+n8QdYBaziGJpP9OAse5
zEPT4CRNjD7Etf064vbyVsz1l1216ZywAahTRk3iOg6kZ0r2b3UmRB9nghPnV7Ma
4bzgReZlMaM76MnZ0+DzlJMD/76kEx3MrwbWEg+imcf0miU6U5XlDWjJPbFTpBRu
CKrYLdqdXKKemkd2j03pXJM4a7fkIJzVmYeR5muVIZEWUkrZLi4OJWDzPTTvYgkG
mJhFiFYNMqlVw7enlqqr0NGZYDmpG6nIgiJ+821JHX/jiupOwCxBp+n16kGS62Jf
Z4RH+C7oDcKyiJZGAM4tOjQn3F/1J75W3yCWxjpsvxek7+uWBHFY9PDZJRD8iJTR
VppI2v9mxPogqSzr8fVb8xwyjkRqGq1ec/YYOA88f4WfgXJElUW2hfI+ZcSSWfS3
1dsam0PwI+gYvdFAS5dRuDZRWTaDOzGGBsLn2K1g0e+WMw+b6xkMBKqa0e40Ersd
d8Z2ng4JKhXL1lz7agn6valrpD2qja/O0GMUK61IVc+2ORO4UZ1qt9SN0c0MMQEi
txMEv5DVkaKes9Ovcw6nXRvrNLsMEPMlzmKo0cMzwUP0ddrCqa810XACGfNucSy9
nUPMG8w+xO2EHdX0zF8dNrjFQE7bqrKLjEany/crtUbkavH7Aq+QqRfYaSEh0YRz
S/c28nPvrtc+mCcBUGgMaqJ/zjhKfFI2AX0o0LH+Tjyaen59J9jGgSxhTfSRgv31
xoINGKRA3dKc6CfP4gCRSga0kf+qS35KchyhK7Yx1wcmBO/PwwWw0rxdi329bI27
1TIG+ZWv6sk2q5GtrJIFwBsDJmL3enqClSp4or/rWcvD/VM/tWQHasClR2Y0nkPS
slrhVCaSosAnMnfHKLnfts3/85/UFNgPRS0tpdZjOvZoOBVolw/Xvl57FZjWljXR
FQupiEA9wtE79S2Pf011d4iDR5Oi82j1ybRJr1QX1/2Z6E8V3iRNdjSO3vCbVdcJ
HJb/NCVduCk+vWDUAX/3W6BpSSkfKM4ZHWboki5lWmVC0Z7VP+Ul4KIc6Knq2Zht
jMJTu2vvJwAyN2ol4Wf9tyQzcOB/6Ho3SxUBXvOisOo+vsPR5aWxFU71a+/qwmf/
8h8T5gqycSSXhLUkJebRFca9wxoUfVnA73t0YKR5vfdxIrRubR9THp43WzFoe+1A
F9OQDP54HM+1/80GnNe1PvZaB4m8bdzG0GQBSNLoXNQWAgOEhOqooX0nO6vAysBk
Qlfu3aWJBQDgUIZcy5vNyBVJ1E+5/YTYgW8MZW4sSB0H6t1/l+ZSixjreRmzHU4N
NUwtOA7sQ+GC57zVd8IJxxnRT8cpYIWCRLvvbhaCKFdy8pmcD8a0drcuPYrGuue9
uGUF/ZWpCsMsvMhQ8IVSWv1vdjkbaC6eepIK6KnSajY3XRXvDC1q8U8Igu9zh38X
1kxIjsNHITPPahTnmVKSmjIZUlLL8ivSaSEy2W+PtYwmvgWivU2pAWodc245ylCl
6/tr4CtYmY7r+4jm85UV8dCj7nPWKZDCfDGoadmjwoULwUxRB4ctM0qMHhwRWUY5
7H0GPCkAxLfaBgv1Ou5rcHDXW+59+QSwyovfs1kGHkMi0Am35FR0THwbrGNJZgxX
ww5uNRhj7WieYzk9zf6aOH2y4vzYVanue9X9O5Crb9rg1zuyuiUPVvvC5hKsuEsH
GHi6SPCvzpwCphVOzpgFPo0SUxAnHTJPeq+OosjiHNOPmztPAfRc8fZopxzWWEHw
S/BqDpUFyZt6Evu0kngxITRZoxIWKCAuzNBcyKTjXBkLMsM8GlGKkLw/O5Bim6CP
YYsRMpfPRMUy+7lYQ5K6jPTM9ZjeDokubX5EUXpsTTUHHXL1wlxS5HGdmkRbU4bI
gY5AFDR3X9HWnBYhglvBG3gEoTUNlXPV0e0aOSmIznMbSINEijx3wiPfe5Nq8xN5
bv/m/C4kEaPVjAWYRKGZS9NzMdrJHb3fX8V7i+le8HTmTScOp4s1G/ofwp5ifJuG
UDQ3yDvblXsNoMZ4c4NOvOGIoAGpRaPDM6W2zeEYlkHs0Cgehy7CrTTjgUT4pZIs
CJRUOZpNG72mHLvtDBt+ojp+eLcDYhdiHDybU7jClf9DRcSbB6gjP9z/K6TqdAGj
7IriTZ4U1ZN0yAMoqKouLEswpx2yA8udJIXJNGWJcuFOldXFikSiGn1pG3gpBsrL
4f8E/e1wPJ+2j3bsjb5cGqom2zx9Xxe1XYzbW64JohHaWAgE19W7S+pTeB3xCIgP
K1jXOhERtBcywTdst05eF7nSbxCkrpk3bu6nAbXtg6h2vBvVccZUMx5ZiKsPumah
p/W1dPvOQC8llv03R2WFC0xb8sbcbbWA+7t4AN/SqXCOCW31IX9+/92JzxXq/50a
RuUf8RoXIjcImHVKr/qdyhLjyW+r7nEbeSD7PxnPSZlDw3Ou8DBMVBWszEeUTPO4
yGXtBm/FvBUExIeX8niQ/66n/YKJSKbRI0nAbmaszys2tB1OjGhlYw+HcXZPoNSp
WB1u3a3CVDxXGjchFacFEYGVxgyCqPic1jFIy5aDN0HC12hnCNOLaT9ABOtF4gjf
+7YEGuVLD0JELGb3PO5ZJdLqZfNMgFszkqKLFHEM5QmVxiVkPXSMlHgoias+Ls8v
7F1gUXX2YRfoQU/m4vz6CwNp+uUo/V+qir8kybvUyYxsdTH7UytY6ILeK4JtDF2d
AakqhuDK98dA1MdSqAttB1xuJaI7BqEWbT5hH0Q0DNJZ4OQ/Y6PX/DPXz2tjLS1A
omC+LQqBwEwu8YOeNvWJ9QnJjDsPa95o4e+h8SEDHZyn24rtqlQzVmOOatoQGAKD
OHUgS4W5SRF2XGj06dVz7IC6cw4w3RFmzIfOc8H9iBNBVWRBBlR30zh+CvOHM5Ly
ukueOFDWeR/7lYP3EjasAcl7+cFauCdxM3oPjBgXq4v7ncaWX92195U89VIgg4rr
RaHg8IyyDIhVPRWIJT6RqWY8jQlIZD0ZuYzJzAdNoQH7Kxq6RsxBHK2SgoKa7JqY
bTsGn/+JCHn66kaQNNCKYl/vOUZ8As+1fRClDs5xSG9ux8rLw6DENG670hajJ9jr
zS1FbtCb1KzjhdkCZ6daqV3uHS8+sojQZppZzi5FU3DyJgTjeKgsLenNqUCXPCMv
kOEcoG0+Ks8GfwTthFLCEZdoAuE5CWth+3TTdABbB9YA5CDpIB9euDSOdUVjYcNq
FFxVfChuAvx1AcbFMRaKel5Nh0ykU01yRhpdo18F1FuKDpfEUhDYiwAljW26DGxu
bT+UDrXvsTJUtpcD3eBOH1dIqexVf8ZhJ0aoyBX7CLiaeXIzEZdH/q5zYYkN0sYa
lE64jRFchvS0wSoG/IvVVKKk/cLtfdiY+JvnCIzbttuedpHiYw6YP2zJ5QC453Lu
Kdo8lfBgysptIlDuaYWVoV7RJswUoggpqc4vXiKuGT3nD5wFVnFH/wxC0GNGJMJT
Jx74ZUNBkfN43pTyQSdN+S2kWWwM6Ne/6SQyhFOsEN9N+Vm72lYyeWmg6du8K7fP
cJLq5jw6Z2OnQOSTSAgEwgOYv2K1OraChlor5Emq1oJw9gZhsGTy0wbbVJ5zrwdl
cWnF1wZaxeiQCI6GQTkJeWmIZqUB9+J7vvKX4udfCx7KztDyA4bKGPrxRvtKCMl7
zEyK53jFk128JDHNGSGREeoHPvXWXT//IctFEEl++Q+4ZiRRWbsr31Br5ulyH/bV
ITIUuyc2Nw41W66tApSVQ77uOwXc9pOvj3CNS9joTLlDgN7I3BHokWUDknVImh/E
usy7otV0MufzVV2MQIlwInFFupd2C+DvSJh7gieVdxicmM7y2QEqKZZUSZbzMVGg
2p3eFcaQ0MfAOMFvrC4XxrwOEq9fo4zofWZSQfGlh+C1EVDlFDR6mSyg4L+abZ43
whZ27uSJkm1tO+LFY8hArcz3KCxqA8yyFasmPMd4sk8jSlCwEnJAxQzHZGzXQGx9
2RCLZOlo+q8m7U6WoW4p2/mZwW7nm8rjKt+/2pn9SdJ2qv+sQWgXfgi+o8swU1Qi
VG94o+S8HhyuXhr2+gNeyumG4cdZIDcZoDDxl3T1GQPIcsb4FvHazzK1q1Kdpn8q
S83/Nbgw45HcN8737IlXKTTHgmaCF9A78DOxIw/Gzax7Bx5YZrZlPNrPpSdLQhCe
u84MsfGr9VIwxjixEZOjsA2G1HeHBEl+jQErbHFLcdcI4d8RZomVFHsE1rA3lhre
41THPk7JSRpDsLRRYtdJeeHWZ3GagPlk5grrksqEJHC4Pq/9jqt+bcp3lHfIY84r
kpV5vfsiU0cFabRf0+hubvhkW1sm9+NaUAEvLsuSW0aMs1C/YreISplOHaoHZiFX
nnlNfxdQOqRwfg1gut71iuNSzi0BfdHltyweRr0U8txrefF0dgIZwCkYzZoaBMLf
DLI8R4bDgcWsjkjd8+kdZ6ZDxDrQvuVGhZTNUEQe4kuaf2uQ/ADiAGHQonOgMQ3d
mxcQ28zcB1oIYnBXL2wVxcbY946GgHKtekfSBwnWhuNNqunspowjTrPuZILFfHuS
IP0PLzqx/7GUa4jyQ78grojsuX+cf8OF9iJj6oHwjIl6iLSjlpfW5thw7DqqHyDY
XrQb3bHhwx86QqKq/Gay8tvqkBeyHq+4OhfJuzQ8sJWa8wKoY08LH5X6J0OLUyby
Axugyl70cp0+hA4ypCiQrPZUsWDzjmL2ZAw3Lx878FyoHiBJdjw4NsvPVfsKTd63
SEGexthIDbUvGcXTcUHYwqtXCxSDLoWsYeOlJ9zg+rBUJjWp4POKtF8Hs0yvMGHt
4gs6yt/zwx7tJHzyiYhMQhqmP/ZyCZAHkcnuYs6AnxPYLBFAty/IaDTZYcfGaRSh
eQlWnJcCs9om1sVp+aJ85KXy176BXvtrlKVTHCBwJOK5Li2NWe9anyAlQ+DmlB9G
PHGn4KgelS9fNKQbcn6k1Ic7Wx35SquVaUKStG7zFl1KzsK1Fl+0YsmP+5+TbTb0
wur7zXfDuGPcoMVkjO9+eSSzfDnc5zy4rCLKgyPkfmDRwVrFJD34HtNBCo6Xt/2e
3dHRB0ab+rBbpJC84Hoa9G+4G6dzmWMm7tQmlfKM62Hqsa03A+EOpffsHzZU7umF
TO1weIMaYqKyn/WsUTxi4cUR9vE7CRn8gsvpK6A44ZXI9sDyoOXKnE4J31sKUQ6j
Rox9s0Klpo+JBzdOZM2ruXF+ChRIY6eQteZ2rebX8dHQ319Ft8rZ3AujCBRFMHYW
qy7LEYj1omVuFRBb41N830kfQ7+4mjNwl/BArcRwivLPoEvPqBQw2bWoEzd7Oq1S
VlRwmSXo1UFk3l+nfYAnC+FQ5ng+Xjd+YW30VbpdyPMAq6ZUMMb+sMqRnV+yDqZl
tltxk52NxNEtgvp9Rn+9pg5GioqFy7Wi74BDRyf5bX9fWm6X+KLauQR1ReiXh+zy
5I3w8oJHDt8/+/YLG6DgTL1FRiK7K+YQxUe2naJjbL4wQiA9MQDccCwXTK6NviI0
qsjILOSZErw68klwMVL87Ri8Vhjwu5qwm2E0tGiSTeU4ZvPeFDO9KoHd8JsH2eX9
7pDK+2QEXRZLpxHNA4ArFRg7u9+2Y9AAu0rPWdfx4HfYPZ2llSuzJaYCC8XN2/zK
N4mZPs1fiDSFpi6z5q/o2GNT5zgL6QQzZ8Bc8FSW4uzM5E4bHbRR06gEx+rbpHhm
fqcp2ik+PSA5IWJG+kgky7bSuFvyXi2puEeT/t6R0iqFoXTKwRNuUwdSJ/djE+wb
WvHOfjDIoE3Q7IjG8Jjh3ADqyw3hFjrc/NeBTkxeblR1u6BZm6MF51PSAxc3aX79
30G/0yJ8gaDKDUOEGu+FHX3dtjymvT52mATygbYr9HTyt8PCuXMbv11NrAnVh2I0
d5ThFvp9kvV0i4eEFMsK8f1gmbD8vWAJNu6ssTlKO/priqP1hP/pT+cRxrA7CyZH
EFneoj9LGwn+4JKB1Iuh98B9dmmAgAE8r+muvVrZfjjodp15kjvUI840XOuTeJRV
WP9Mn3wAGvpNVn3pDxpYly8BWrP7VtBrE8QNWD6g3vz+MmlW8/uPxvpxpToGe2bd
cv21OlJS9BKRdK1oASqpvEjhLh5kyknvgI/dWZLFzkkNg7p3o+o9UF9oRyj6aNGB
LFFtzYZn6Z7Uj/jOEOajECNpHkIe7aK/3UyR622zbEZD+uB5tZsYz6IcwuuHc3r7
tDn6LMp/hcitLXHOdzm2ol3PNdCDwyoNcuhWzmZBYboio3MVa+HhqU9+ZOfBTtFh
6idDBHzyNd974BL+lI57tcTZEgALy7PPvSfZLXPkMKM+TjNaoA6TvaosKWGzrNfP
TSAr4mWUfDTukF7GdApbfbadrk3kBlyCuTlgShBm0X+z3jOkf3AddcyLM/PbNvgG
SKqP8MDS/ejmDMV1jJlQOEAptMMTX5Xnbz1mpHjutfq5NPNOw5kRLuQuZaDXw7tK
0qCwbUIL7pQxypInYD5nCttcdIh/ZSQ4cFc7N82GANXR+oH9d6t3IfOLiIgO31y0
l1IcmoqXsOnAlkf1hvrxRg5RORlaXeyDvROm/YkcAlytz1HFtO9z8599cX5U3zdg
xLIK7kn3nQ0IKEuMN5N7ZAiJAnqYs3bJNbJ8XHjCC0+RRancx8zjZvyIjeMOR0HY
dqhDTeYssCp+91Mejb/c38pUMByFf8JxI+lfUsClNdUiy5GOMlhKBUj+WBKuSKti
xlg4GqpvnlSZIHQIANL8uD7P8CyMZ89Nr0kKNtr3ZeeRt3Ps4VNgxdNWrLmv/xxy
aGzPT2rSg3MW0k2ddPVbY2ujOFvioNU5Cn4m+IeKsFV6ImrZhA3ynQJ/ghVg94Y5
pnESOlKvpREpj3sGL/HyJd2dOyBmu8Ao9pxjfHZisy8gcKDbc34sgfgoBPCY737y
uNR+Re59JSBOPlU3vynRTEjKR75l/inYH+1iI8Xvzfa2ZLdfVkWKH1QqNX9NAe80
JiorsXfOvOp+l9RpaQerON8bWbqPb/buFjetZO9B0hdnmbCkZ6nWHsWOh/DOYZx1
3X83fs8dwfHUTsb1SvzhyRPhIpoYcqSsReJNaI3fNek9PMRHMXQIKu8bA7FTNQDw
JZXE+t7lRak9/HzDzfvJZta59ajFrD26kK6gvHjH4WNIux/VBa/lVfQUhfdb5ga2
qyMJDyKKkJsN2T5ldhoQA17gGHZjN8LHvaCYKJXFTIGf+M120pEkwahePUlF9qHt
rLeNKqHuwLanhNttw1TJnbd/F4XPzOKTTzrt2y5d5sl5y9FRnQS75lHkNGDGI4P6
JeDeWcxKe6V1CiazjNm94mbBeJ9nPe/ohm7OnHVk5kooC4ZN3jk/cFf6c++41HhV
KCvdMZAzLQsYeoVrZXsJOTG4ZgOrDcIhMjqsKrgPF5TUkfFjYQRM7uBft+0GdCTY
8QagdWTZfOiGD9hKAh+bG3vwWMouz90W25zGJrddl+D2wTsgfJ8i9emId4IeIfJO
m1QytBORaJcejVkjm3hgNhQvwFy5FTe3CcR1hOrgwftUfic+l0+eXgpJkuUk++U4
yh/GxXE5k6G8vWIGQEWOFOJmO7yvlz6EsS0RclsqBQqiVTyk1IWcnhFAz4blGNFe
WBt7QJOEgNDmuySlCeTWPs4oHBPbNIgFydpz7Xo7FIKh5a9U2uEU0jKoB8JDUFNv
ktEaTd8rlzeoGLGEQkTzycFgaaDEXhBrOj9WVrUnn1FiWpdjb9u5egavQ2QnkWLq
jj0DXlbEDaqECBUKLI1shTdNg8Qs7D/Cr8qGbwl83N2+Ji1JpBfxu67E6xbgvccQ
/A5LVayNpL4yQhqBw2/XCLVLFfJyHYOHbIn1PpQs5KuTfYl4/gaCEzNluWG//uTW
HO3DCG2BRzuOe0VWOJ4Thh6O5k60VYseZT0ae3BdgxrM45qjLQ2NDCpSJnkjfLxE
xTGF4KfDmksk9zxFjcgZ//m+M7xRjCXP7M82P9+cxtUVl0QdwC7fBd3aQSuV5ShT
DAbmf+VxqvqkRhRL+O32TW/2OY/065nndhLz2Z7ib7qHr6EPnKVYBLRHAbBeY/Of
b8f9ciRv14+2W/7QcpLomcPSoelIudEuttgEeDFm75a3PtvfXn5LfFYxi9fQgxi5
enKa/G1wOXAiyspQSSmv6I3RQVsroT+8OiJJ8820ij4FcLW5b5FGFLSrtCCpgCj7
PoMg8YmCxw+KS1XnraSvD22dL0mjFisK3sHKh2F1IdocstzV17m3c9ThMLxjAHh7
UxbG4hsU8EOrCbSgzIemjr9faeqHbB5QF5yMgMAZHOSC8tFpwKQhBWyaNfUTl5xd
kwCgtUEMp2qIAdWEjoHrKjqXAnqDupJ20ZRH41vuN24G4w8rQNwrFZg5cQdvivgl
28RMcSNHFCLNokA+gcBViE63ODOuOHLlwj6BCjHR+aa+FjSE91nzb09fHaKW3KW2
n1lU2ZymInf0NHhlehdyaE/8YZjWtNY8djW7FEMacflD/B0iU8RRS5uypCE1VBZw
ktPofBU2rb1PDTCEA/ccQZi4R2kSI+aKXuXCsi3kKKWuJM11mutaKI9YnTkXFJdW
oTKV2RUnCKPiTC1VeGLVH0QtoquqBEmuSqyMo1CEg40MqviiYuO7T/2rnk1HOGg0
/uWXs1iOakN8HyrEbGi/eX91g/j1Pvm6CmOS9mgUHES6/IF/zPt73r+NpkJ2iJjj
TVU5w9ZCP4w3B0+3vWl3VJa2bX/cWM5lwwh4D2Y6LsszioVQcpJx0EXQ+/s3/bFf
lShrR+dk2beA7HTlp18j7HWYZnra1jpNuxBqUqhmzMzRUtB4brXJxFlkjellszsn
Jjyc3fANonwTdtmgq+ZRJ4aiC+Cvf0q/9I7jppMx+g2VRhHRO40jSmbZyvfIjoRx
bXpW+Sq4BvUca9Ev+uXxUXRt+/bz1SpEIWJ5EvEad3aujt24eBwfTp8OMF1tTfyT
LryVpcv/cwore4HQBN4LveZzSk5ltpAEvc7GBKRJPdbZ9FRH6cVLTwqKJv3OdKIB
bIKKz05uFKWaqKYgmOjyyukIZ5Tv96Ge0dzmTJJ8f0PjppRIlmozGIdJtRPO8iv9
Uu9ALjpjsffylPb2WlQXWn4r/T48JjkkkUTmI+AfxJ2zWY2TXAntyNsy2fi3C7e2
bfB2MwsCxcYxUzTHsl6ov9WEr3I6X5Eq+HhaZqsIWx25KsKGle8F6VCOy217mU7l
VwPGVM1W4bB2xVsrrouNLv4T2Tc0WsvxD5Zf4UaHnW85qsywtMVhdcFUhC8wghtG
7EeM6sPep15R0luOkb1oWvb4AlEs/1XivHNl7BNFa6M7oZEgnHHHYnq7STzxp/WH
Qvl16M9xUL7VAjfF7dXYHwSAV9eEF9gtDfnqc+02wF3ycIunnCaCXwGZYMtxg2Jz
HQS9Cs0wHJbdyMsRF/i4mrN32Bor1BpCGjl2LMiI093Be4VvIl3fBpCKQH15E0B3
WoByXjT+/S+ER9xFzpP5qEQT6NOlhjQSwyHCrzgUxTptUT1xEwYyWWPUDFn1yoho
V/5bvkX9eobMVL5j4zZSd9lQ1yjJKYdEDF8QGXBcF+Hc8J+nMVjb4lUDvVeSwQsE
JmqlaQos6fWr6dTSmEbiXUEL3pEb5U9ZzxCCz9BLEMHsnYDZr8SxLLYQxsaR9hcz
/Yan+uh+NA0wiyMco0A1oODJ5TfvE+5ApFhBdeIsmDMMZuyX/AzWvRdJ+iMFzsoV
gr8pJu7kZi1YjBGOH4INKqDdSnw/jG2UtiLdkkARpwoclA2m6xElcdnT9PpNOBNq
JfLvuC6Qg5dLwMTPeYysJ4ZmRYVP8rC1IPDbjeCedFuhJ8jkTH303cJFxheJOQSe
mAKpa+Q21edu22I9RRMdabSCPsMyAvlT++6GlA/raQN8sffB4fFON7Ya9FcJA8Kk
IDImWbCmY4MuacWcU6znRXgHJzteMHXBytPV5B1UkxcnkTYRvn7mRqA+DFSpLKz4
+SCZdXshdSoHU8gH0POqi8dmXrw5DRPUEPy40Zurb4RXzYKS8VlaTP9W//mNb+3U
O4/C3Z2qXxGNtQtAEbW8d6znnNesdMA4Kree/8yluLxWxk5arbaLELUvb11INIJl
98iCC7Kdh3qTFOxjxKVqyxAEhwjNzxy7prKj4+Oc+uDXZclBHR2YRuuQevc34fd7
DF5wzRrJhTt64yeGZ9UzHdBD9zd+0elvQVDgZzfkHo5Kj+X9481PLdLzuf2KKrbJ
dcDo+eXwvThyRZa/Vzoeh6g7ALWJx5BpE7x70xK/g2pO6yBDcsV7XeVbKWttxNAU
38gFY0PXYliz9e5i4d4meZIRlOWWbeeZzFlCXhnYCiOw7RvQFjh7gdRGRLSUfu+X
k5+u+OKaiay2/bcM6a53tXd6TYAMgeR/4Ue71s+ygGBRGH4XKi5rWQJNaqK7GOoz
Ynwwe1ImEwFUEjRDkK6MOHhNDca8AnGwirz/71b2lAEpofchpFQPllrvMfO1DGmz
JbuM7frFH8ijIBLeXJNVh/4gvFLsq5gDoNcZWCgsVDqG4vzaRnu6DSnix5bGQ5Sq
O/rw7gbty0XDbdpnyp3gdjXKt40bkJoODpRvhW1Pql18Slo3L60v2tMpum/xiGbz
BVZPMk4yHClsCnF157qUh1gRR7KX5JT5sTPfn/1+4n3FW/AxqEWQ9D0B/qI0VYQI
XA45paoLTrCgRxQku0CUUibAogC4gRPTUo4PNkxP+NbeocxTYTw6jGoOFTCpN5fr
vLQnhTHWihG0aBfuGAVFYreUMtaJ6lYgXIGkLEG1rR5YX6Sd2MH8/c4BvHuRmeV7
yUO0nEPjl8Fv6BKm1vh/aNDlWrzdQa8559MgX/aNJgCUu/VnP3XSn5v/0DYZaueJ
tgouUAC9WEALeIVDrupULcwDwZ1HOO2DSEBwQ9A5iyKtyIA7C2/iFoaoHuhZRYs1
msRjNAtj524rourHeudD3SlKK+7VIJ0UIK4vlg2vY1gz4h9kr2MI47W5BNFz0v+G
ljp83fwaQX9CjvHW7OIfMD+XkdQvFq0Uo9C1mTZHruIrYWxnSutuXhNXfB6mq6D6
/bucV797sdm4xizw1T6Lg0boWoGJ4p1/vpni96k1oeSr1w98JOVos6fcm8cw9GRP
uGvsgEgMCh1XMiMnMDEPlqV/MyY47vIi2+UZJQzzCeoKe2SKjBvRwWKOieJmLxYp
vzsPXZPWqLHU7aWBqkIy4Z8H6d48ZwO3/DoXsyOTR6rFpVYsHexFMJLcFE+Mkpvl
s9d+Tv1xAGV4YSpg/WEqHWLGRWjZnipW/ZV2qNg9JdfGxZejFh7ERmQqullfxzkx
sFLMD2W2fYx4irtibsbAEtb/R8vWU0Dp+LBkPvK44on6dTXShmNPun0Y7LalUTA0
u4asFvTAkmZKk3sLXVFjp16cTH1PuN3yW8JeGs7KcD7CcA4eqc7xmHzrQvI+llo2
lhlzV5FWNdsURGaCr2VYb8c38lgrXWCmrXolX7hhFLD9HdNQz8UpJAzIDbSMGcxz
lPRwn3F6Wue8+4Bd50BH6QRgohbigs7bCJMgy2UU7eAVeanmZ6LnkIKUuAk6iBe3
cJagjqrqyrKU2mPQ0jKMacplXx7RKbOpSfj9F4sdOLeG/BA470DmdVMJttRWiT+9
XZx43Qy3r0q5Ct3IWsiR46ITT6o6P2MuyTVoCPwtb7cxSngf1mB+7JfusDBUFr9t
QDAjkYUsPFaQ7SqNEc1yv/GAmCSlOMtvUz2ILKLJXs7pIo4tS96UiKNwk5riqCtW
k8jAXxmhVX0oLKb3xVaBB7wMyBA6IPsU3UeAshXzGlu9t5DmUQ5tdQTue3x839WR
bK+rM7fTJe92ZMWqfwMHwTFNK/tUwJHUpDIEQGwf03JPazVSmiQD7o+FGFaWsF80
zu9oSn+WTnJgcm92UogKuT+MWQv1vy0uFqDSXEw73ktoIDj6P2TiL7Y7SIuaLAxS
i+4fGqtX4Tlwt+DMhzrqcFzi79dZpWuy+wRa6vRE85SPbMknJIMdioM8BB1n9IV1
p6YW70pQW2Uatl8yrKMDW1zhve7Z05b6EababMj3GLfwNqnHIP7N959Yqtbtr2ZA
dT0cb6/Epi8H1zYU/zEdy1KA0ppnhvMa5YNAU7WVE6vEOU+vlQAiaM66f8To+TWb
dsqJmxvOfSd9TgGohRxtooqULd/GVe6hxO1s2QGmx2x7KF6whY9jYL5pGvbvS9hk
+p3ZXXTKz7DdytiykP3HiIP4RFgLky348eAI/4z84CYNowka6JMpyHXU9bVX507t
pJ+reWxE7kuO6Fvt2EpkWL1cOfIRN2O4GyHGxVCpjrbrpkDCWQwT+VYK3xIe3swS
59WhQfUVxWyOsw9lskr3bE+wj+7C3h3rYknSF7yR7O2VpPA64KG4XWFpqGjDpiQB
4Z6JMeRTXkU8JrxV5/D8TZv1DO+4yXzeklFOB25u/12F2X3irZP91dRoTWApj7o5
PziazWNAfUNMdp83QBpLpmR2VDz+hIYMLlmHGYEEn/Kbw3JCrM2P7IEpfmPJeFgn
6Cym/T8tN9KCq7abD//YFpZnVjjyOwEmoI+0sdUN6gMLziwCBXoyOgcdkg/sORDE
K82S9zvGG9oIha2Gw4WMrRnMVu1cgn0i3OcoEO3U2B0bAZQqIS1UCthYxZDkXrE/
SrRaDietXRPl2ws+5mCOmjnpr/vkwIEQKntaUUJFtYxT6+wcvy24+yDaTHhZC0Qk
q+D8gpNzXX/7unMNjqjswxMQNabro9kr7wVag0Tcr/2OZ8KSPQqQt+yd4YdpxPV4
NUmc5Vf2rrV6YlCxIokiYQxtDeab8sUtOQjs9ZGMahfShC4tXWUP0YeyoN8vtoD/
MbMRzo1YP0ugW2CZLOXhq7wUP6hiwtkEzF5dDCLxjx78a6dqMGCdNuNoU8JfjhTE
YstcWk/mEfNvMV4e3JBNcfnPzZVLVs0DxphixkZAcH1ySoByCPoSidtXPDrZzims
F+fvLBOnTqoP27I+k0LLwEhawo57HB5rKfZTSsg/sYrkYBfZgUVYMxMELEWxFEyX
0/7u+eKKQFTOE0uqc6oPLD/rLqrCR1/UpGp3zgDgG2Bsxkp9ETtcziznq6J5NPSi
n/SnHQ0mz4gIPHngZMMkaZgyYKk8WqLUeD2+w68nMTsDtUbNDb/GSI1okuGy1v5l
kBDvX5cmdKfH8cthAROpAfFzOnICRR1dzoaWY/wY9VO6DJmg4rzoVXR4o9KlYybI
d1byNdVnK1AZeZi9k66Y4dCkIDbktwwLKjq1wHvG3wBhraVpzvxYFvNVwpkVYePh
2Pt+fF6Dso1o3s9bzkfQjjL629vB7KptQ+gv0wYFRXJ/u7zxzhNZmOSPq4KqIYo6
1xO3Xt9nTxDefP6xbRmErTZpae4KV/yz5jvq41Dj0NYFiAeGhLeVWRh7FkZs9gHy
R1uNHiTttwxzSrdaXdwGzXHHkdJHbbYPqpkJIljljmksNgnWQqr/0QV5qRR+guJ/
YKJggEUlA9l/MXMIrVL+k4KXPYCpMoFPcF3FeDHSHpm6CgtqfjV2Gd4PiBPucvgT
bb8b8RtZCgFb4MvzoLp/To4Gvfqa9rg1PLGOXMFhAayEPlcISs9JMqCCTV3TqTAP
0Ibn4xzkaIaOYFzBKfu3EaEdNTJmc5a2kBTfdCHTp09gMdR/RIO7MLFmGEVfodx7
PsXZNlfal+/0H2YVznDN+hwLMEntU0nHYtAGmIxLBrLxRzLMeXks+dRAtSej/naX
K/d3wV/R37J4zRKFOW47SaPZ0rXyxG35z0lMsUdYugM50oRj0c28NtYlUePkPuVI
VxJ+QQQXIpgfSt0b2ek/QehXFn5ndS0MURqH4f+oMXitALmUJFZ30UyzJFiidAw/
mlJibttrst1bWji7UgknEuHXfB9bcyP0D7WybCLFwFrQlwHUCq0WJJHgKYDSDAI6
jsX9ibDJs6pcKY0I1KC8Gx9INaH+tOtIzEgj9PAf7LRZAilIzMbghUw/OyOi1aks
L//hzGPZceRKhDS5iuHeBZaYrnC3rZArlMX5hrjgHNh3AVXoIl0p/lFTNW08Bjpf
hdu2KKwBdUZI/oPbdZwS6FIrI1KQ1lSXQ0OkBxglnCb2as32tR9gZvWOlTbC1iEC
N1YK4cySjWes+ZGLQUmgMZzjIDE3ds2CNo6k7dANu7y065wYDxZRCQMqqbaOP+23
IiSqjr0+C23kamR9rBovgf5Tq32NgvMCiY3Km/5sidGg9XI7+jKGuU6NO05omVP3
5j+dCfvzNl8t/CU8qJuaYiOWDzhI1zyp+nEN3/brEkkMB72gRbuDNF9YvFwqnyne
9Jid6vie4rRmEiNg1mGwDvwLabG1j9KaRT6UK7off3MXzjMAFgvGEBPxwYiwPqox
QeYlKGOqM8HlTedp+T1XpUwBFMnzr+kYNZY813aIppz9KE44tB1jLnkjmzbP6CAN
gimyPZx0FTlIBG3t0SLJxvmjIAGEMuuPOemOhaZtzTf9QbdmoydyrfasBAefsp4p
mZNp60A5TGQSwrMhUqmmZHG/kP6UqObMNTX8MSieLYiVm8KcK80T4OkLjx0FU/oc
41M58dyquNhoP2QH1+4fq+hMtdkeeIUkFnpJ1qtIrA+zjmi5mJp1sZBckYbv19yB
uNo/agLsPTQPQOQi+Iv4kTuGPk3OP2lX4ssiIkvtlSTM3GXK1nEkkjA0tsPztH1h
xYqdBbbLLa8iESlUmFn/GuqhoSc7mdBLVHZiZMJl7ODjXqcvs/VqbGVOYK3x6N9C
JtDE3CyhaqvhZ1PtsLTjPBUgtClwjqERIcoD7qa2mupB1yIqIrQVPjkSBzSmkHJd
Fsw6XDO0afAm/8B9sThKFBGq4HqIL3pE3y7nR1Xg4j2YOiiV+HBTeFxiV2KD9nfN
BI3ilHEISYgCNQy+ys+BeOpVDXiVCLxMSfzx+KxPos0xUVPflLSZTiZ0lUx7TTO5
0VZ+tzrHMqYhGMOfNZ6iQMKR4QTLeS+hxpG4pWJCN7A0KSVNbEet6ftbLSMSJS71
48MzV73tBD2xEKar+E0bxUE1kJfFPd4qVVMIJFMtATZk6a2rMxhSF4v3bx8p+FeW
MMi1g27fwhhhCJU0y5kMnKAZf9UnhhNdtTJ1fdeb3f1znYkZt6/lxXPDzM54V5nO
Uh3kjiOJTUBFDes0YHs63lurNwsxKbwqDOsIY4sNB8jHml64OgaPaW/t6lqNjXS4
olZt79K3Tcw65zQfBFxzzuHubKz1sXeC/J4PIt8fYzqhql5jIKgdPvNNImXGMjyo
l1i9CDUe+3TIhArqZfj/bAQmPKyknjP5AgPA9iVV831mWx39IS1YnrGnHwwePGax
vzpFFxUKWNW5hETD89+WxHCsQz7+O3QhL7OKRb2CaEig8qp0uxjrR2VTsY9bh9Qr
BYBjGHGS15DXlyduqgdDuacARkwweZxH3Tz/xv+gX4quyN4IGaD2VrGERoOrYm5n
ZfSiG40ojgTklt4vn32Xtg3c1PBBiBh/rKmDmJlQGyGazFyEjGBze98pL6oqivqF
zls49JaAYWY2UPWJtULbNeKEjeTB/88tV5U6wIMRbzQ32nBsqI4u3TmUNFOE5+N3
FB4gTwsPjIPKB7/e3AWcT/qUWMDCbbCnKzQgMJVrwRPBo7dAQ4ZRWeDTxKePhcVj
IlMiwRZlxPFqSHsfpaJGaafjltNawjZ/qA1xOPD5InctjYQgaTpnAvr3SDnteHnS
zpMzpsw2DdhsEfq86co+jmN4NOE+bzpSfo89NAmxjeJK6o1cbeSocnYhqVy8RJKx
vOPs58ZE0RFyn9yy43B+6yqGvasKboOx0Tq0okVdUFHo3Ae8Fv+wF2GWTea6O/6o
eeiJaU8AVt51mq0qpGC9f6JpUolDmqnv3osewAqXlOz8B+TG6KSajbiPhpo3lLCa
J4VAFng9mwuT0DSX/QIYM/4w5RNbNYdYwlysjmmOACAsswUHGCMQ/XGBkQOSXtAT
unDVqO15sB1qxU1Wq57WOg48tIPasSxzzANQlJRjGXlM30eYiStwPPdHZhlfXnmc
58ows1gxRFnOBGsUEWd2gCJxxOOhbGukqlI0HGyJCE46+1EL9phaYfAS+EOMt2pq
FpdLlqp882jfmulm7YA/DfEUQFx1/OUumjdKAvTPRdbwtWyw4ZZp3TZr08L1tAoQ
UFF3tZWWRxoyc8Q2tUB2WFaUtb7OPC5RSJL651ZvKyvsBUFp7fuECCpLcCt3+CQ+
6yLkevWWOG3oTCIkgF7B5h4cdW1EdZEtflIFkfBQ9a33qBArDhob9nFN28R/iFcc
Lvszgeo0ZdCeXlZCWNidFZkUpJTEo37gVnxI0OSF/y0UKvoVidJ5JHwl6LIrBdIm
aG5daQJ3jV2QkU6acnJePonT9AnrAzro06w7HDYkT5lqVqq3QGhqV0spfGuSJ8WG
S4P6fqkUiYSuFTh/xPrFbVhaJr7XyEcw+/HEcU+gGlrHKtvdXXAfJZVPUrGDRPM4
fvrCeAVKhyrIfJfkl9qBrbNLMgWPiqKGFUiCk/oQVqnQl8pBrhWajeGOU1z9orTa
UMNegJ9x5gCJwnZr0TBFMkzTigEx8Xu2efn4TPBvFw9Zk+5HPHB834zhfF6e+lHY
Jv3+cEsAp+2jq6QbkfjSJVYyOU4HWN9Vgy9MlhYIGyxStDUjn6rHoDzkMRMgYCwn
9Ag2bjV5FAjGmCdb/XirqIEiF5+baQZ9YMXLgh9QYL5cvOkCSSd59tO2GecQdpWh
cXHUu6KDG7wmW2nTYoCE54uto476UgR/lR1MUVvx7uIYLSxgbB+nQGGDUD+EwJkI
5iSTzlIpvv6hI38dBUESSN1KIj3dTnN//rPRY/HuIAKstN8954tqH7OGqhymdVYl
73Kv8S+hbbqrP2hdByNdE+15DCTZ5Qv9SgcphMu7dX3oIAAwcaMf256rCjMh6j7p
KWeRGkiCHboI7Cge7r8NcVKA4Qa+G8h8gq+Kgm6toPi3TS+ZYiNKpEI71baS5jN3
DQoMhDJ8vsaYsLT3X39qvFMk02AR7BOUwQzEUJqO1Rst/EfiRgtqwqmFVmUvHSWa
IFdXt8WCAmZfBH+rB+tiAEe/7eh2yKqIGv7yWMz6vGTEh8Jv6O2sA6nruRybpufL
XJZSXjImSqYUOL6WXVR0Z302Oj5qY3tBK2I4N3IqlF5XXDLSq42B/Ym+9jFc6Z8P
9GQUftkeGvi/L3dTgHvjWOGEZ8QpQRJ7m10JK1LTrupJhPAURghT788qCdaucFp+
Zo08ViOh9rXzoTJIpqJTm+N/SzRv7VMY+XLnC3lAxHdUEHsHcadM+kaFTVGMAw+s
wCw2iOZfHb2vSWxbIU7aJxazHtXgh03d/AXXoR3LeTWiGLC99n4h2tpKcwqACfZ5
gMLraZAsIRRofNfCLq4jQ8W20rAbuJtDFmnZtVaW5/DwmlufarZV/+wl1AvkyTD0
/HAigyGS9LBKITXgIaQM3+zZVTz7A4Dy9OBkn877ZhiPGCof1ETu4txJFlP2kFc1
ZIgaI4bDhiZbgfwLUL6Gj1qef0qbEQwhC8+yfNIK8zkjSiQ+hJ8R/b4WKw5UQAmN
nHXqFvc4cjkFmyBqEqDv01VMnIG935oWji//2UDNoz8qiB5UI3oKuDD5mhKjSTUZ
g4YeBekecAunBuoZNZq5a/UjNlVjkl+yhRKVPC84v35JjDotZtgSdNBwXukLA0G1
awFNfiuDnmRuDC4bBYP6EV7e8TnYvJBSRkAGNvNVTgQsL/i2KldiBzGXCoziLPNh
OtObMFRf/ZQ64MFA8XZRgFE1hbaS34OKrMjnWmqGFOzErKm2wj06CmkGT0+8dtKs
nbPO/35cSHvz3r7wQu2A+kgNR7ehBm/BWHQxUOrcSKn4C7z5BDlv76sW+bhPijI3
FePCZHhj7TpGoDVbJoIKykBAwUCno9hBnCGG2T7470OalzUbLbKT0KZaZ7cVMQ8m
KlA5el10psBTq34TjKmk3dn/yyUlUBVuHkQrEDLjrAcGArTBEZUWBw7LAvAG2s+Z
uFl8/3ARMNL3E5CoL0+hYOHY+HKMMna31dfZiIvXcMekrPOvxdvb6ad8Ru9bAdQp
Vo4z8xHOREJ/NF4VU02vaG81Ex74SFQXyC6u/4kKyouwtwmBArVqtx+ozpEHCEET
gZD22z2JwEPfROdS1osuZ0yiyEGFXQwwbE8NJQvsVwfSc4a8eqgBRTOae5dBAU6Q
pT19mSlvN/l27RkBoH3ZlQmoNx0Ake8vOLJj31+FP/J7uApEuS9MnVRqKxvdqO7u
37G0MQSCdv+xv7/Zn3K1jnmLrAVzbnKoznnawsxefvATLS7YgEJ3xPGcE93+Dy6K
q8SZavQCItap037GuBLsnnHnm3n8aMZ8sm6JKj2XS6YwzrY4kq03uhA83HkpkrdO
qbSycncLshEJWXJBO/E2/SvAuFDurrs9r42xRwi1XotCbtgQ2D6m63pZe9JoVgqI
y/q1DPhld/NtUhmg0E0kR1c4jtVFwefvOqxQsC2xjPhNPbIuRECd1xfJDq4t6uBS
9z1Z/bv1SNy4CUCUpyuz07/AlpTQbeJzbJUfovwOqfQzuZquinE1ggFDxylcdjeW
SZcuNUeBu9wkU376navriHS0x285X/fmGvSI82UzpVsUF04pYE2gjDZpVGawiwjx
TVe8mmoXKdwp5PT79PF0yMMskGqVSSk8B9H2Z4ubAMqux0Ds82lt7LZSX/vUHHVa
HlZebldInVXJi6IH8BaUwWeBoN/NeMYW8QA4DSrcDzSiMi5aXti6hHtozF0XW2qL
3WDIFR9dglhN5mKrWjZNyXzqk4ra7ERy5XEiOi7+vG14rFGCQQUoFRLD3AasMpRh
6puKXpO/f/iIXAK+LnZ1McE6JrwNltZXuoeVcV/Sa0kV1x7+94DBjsFfWsqSYAb6
19PkHFDS3wvxVFoeqDKUhpwWHOG/2uNNhboTCo1kGJ1lxiMxPvcXfq/x2x9JXDHK
82cTErNpDnKH+PT7g2Wyi3Ubn3TaftjDEffrR4/aLZfykPVqHTC4NCnkEz5pMLFA
4h75qObqqf5ZadE1vtuq8u6Sr8H3HfrOgBaIDfuAmUuyhS2W9H3rplStrXxyLstk
pxGXdWHQXsLI4dcPRTRizew1BXkj1WiYGNbNXAYSZjX8Ra4As9Lj1fenGBEMg+Py
nUDoy67zwSizTniRbCyfH3zyvcNDvAPnQI2IZ6fqU/C/yrBH96xqOFpMEhVOWY9a
YIDmAKzhYr+c/578WtTfMxL6bKJPikuXH+fVQxazfOGOyYBnkjSGiC2LkpFsqReF
3YccVQmK8aJex6LkZicW2c1zS+Ky6B08v1vKANjzDDCm8e6hsMdQQBTvJMHEaps+
6ShgAnD0y+NqZlH0fXuGitt2AjRo3F1JOTtI4o9wm1w/4lo4qXVA5WcuVaFt+U9E
UdJMpUafs/9pmTNetl6MbrLxdqPpz3EAeTY8DE1GnSmkEj16+6FYLKyN045iSEVH
mBhqsGlZlmbw1x7q24Pz6QjSEEYLf62jF2xl1f60pL51n/8hqJTQXRoWBVbBR7Qy
VvxcjYVeyT6XjkHkssWZ09Xzmea3a6KRfKjNGqwsrGWdPfAiSKZ5G8QFUNXTKUOk
CGOz4pJyx1JWXuSQ68aLUuTbQl54xfVhraMYf/LG99Zzh5/iza/heAgoBAJLMCM2
r4HXA8j7xCM3qcVecs5iFb0GDqlrsDThTGCcf8Lyyt9gHnb+/ulJE2c10wy4Fi2K
wlKOffCKyVAwjSukNTryURp/8Tb0OVSCI+6sOCo1wldVk3tb9cOSQXw8VmSv1TJg
KwQdGj8nGuB0krHFkLmkTV/gfKWbupsddI6hiPOCD/fyKx7+/OkX7CIM9e1RH95c
mAqKcOx1D8QiJ10K8nzXK+/WbxTez56w8ad9ungm1WHCo95Z7K3r+8qPNpXgIkhm
hR/Wh4hmjJuUSN3hXHk38UlkpRBtdhPU3HMc9JvijyQXxoUmtC4rPXwxlRE9Doyx
c15Z+46zWjrI68lAT1E7UcuOqokLIryA0z3UzqB07+FBNnN1+X4fzfCIRai2d9Y3
1+3kslVjjcpOG+D8bHk2uAXt6qtnUnnkRCCSeoRK35zbdXchDY/IqzSC2Em5napX
O3sJg9UOB64O4WHaQ9pUcbdXa4GILHz9CXpAYJxicNi6Dt0+4XkDYefGkgfTcBlH
BmvmmG9wRwcgrYbhOxdX1CbwxXoecEn4tfDBcRH2/WUgbYqKDnb0ifwdMyge5fvZ
MjWiI368X6qb9NDKIN4XK51tJWV/8OlFR5jvPFL3cQsfB4yGKXNGrmUQHhbCREPT
kF9twMCBpOPXR7m9bbg2Dw+lapiHR9rlW8pQgA0d0Ri6YfP5S3bEH0AA8ppP1XEH
0UcoJReZSWUM3bjwuiYvAyZPuT1EasVShkNodnuniUyj2z9DYQHuE/ZfxQ1gszN2
GNQmrDyyLP2oV+KzoiwRxyCwSxxC0A7P5JejSPTg5KaIBWMhBmMyYIICilOc/9f0
gTh79oKBdgSRWRKkOzJIwlItuGX7Eu9Q+0c3GpyeABE6Bo9yXYbim0DNmSE3e9TZ
FcAG1xKqQIHVNHUQJdgRsXiUVA/gTPGls7sUNwNzqyxgyx65Qooz2pIXKQyiFTt0
+hCpt6imvAZRribkkrrR9K0ZwiRbqigcyiHp2OAiTk5UqWnLuH88avCAj+Gm8IML
gbHc37GYtoTm+yk39ZKE0t4fqU27zmwLDVlnqRFpmwD+ypl+CeNOvepM4p+OtHL+
26VrgCgPpt1p7Nn5CUNSEdcsY+a0UKSxHHtWvhDYnCrADY6E9K5w8QT7SIvSQC37
sE5mxsUJr1QTaYbQRxvavAaMbz+zFvEOdl9iSPDSa0hwGr/3HmF4IVE3k4m50N5Z
AGO2IJBufCZMOBmoXg9MsUI+SRrPk3h8hfDg/hNFALAT+aFdvTCwIdatqjSP74bD
dcIFcrEAqi2O4NpIjdqCpNmeU8QRxPtv8B8NRDgnmkzLIR/NkhS7/NhpM3RqqoLH
6W1o/eh2BzJgokm8fBh2T3hKGiVHQ6VcHjUxJWRyezto263m7jXy5hfjMT4MZJYO
QWoiayNwW0X+fPAuNiMAt5keByDmv/+FS/6LfNfeDPhlZrnhTvCxIGou/NVKaUI1
4fZzQBOPhJYQcxLyu7EWETUNq+2X/QMm01Mojddq1u16bRT06giwdSTqFVjjjdZv
xoQQje0Jq0/v5G3jLPJV0No8lmY9KDkcgYMGnJ05xGTsbxk8VJRKhMkm+Og5cGQC
GvXRBjpS5h2B3t5s2+TTyq1HS0xxHpPWZzzKYkeF1tVDCYoyCZuGSnvKp2CM3H4Z
416/Nqxj5sPMo3fQEATFDWaEvsTlq9z9hYb8o+AwghutSXUwHuuL4W/v2aXRiVFI
lmdAaf6Om67vOVOFe6LZ0ty2KhCPACqeU4HgB+oG3gDi+U/B0/l04Qv3SgH2xOla
LHOATlhu5/gCTh/rOduoOqiMkHCk6KVRKmZzdqUjHkdw9kGI8xl4qs3dA777gY1+
cTbM8yrCgePiGTUpSlZxkaGAa0FgdTK5rvAVN0agXa/QlMRdAaolESxCz0/PDaaB
5ZPSMEDW/q4B78S+hFI41mQpjLHvcg+Jai1BlQvQnDYeOshpqT+580EdHGoJO70B
wl2UtAgzDNGFJELi6fPbmVSL08dYKXQr/19g7PNOIdZ+LlLj3Q7pE56lUmHXi2lt
DcJ+JkQsFvZRvzpinWYRkE2kTHL83/X7L+v409oFsbxCyy4JnrKBRKOaMemRZsl5
64ujhdb7iyXDg6zqbBdPxwhdcIpN/eHvCHbhXGpD/Zxf63Cu8Tv9YbtuDkv45GX7
NnThvAQUuV+Yr2HpTmX/19RbVTXfXuzWYsVUla0Lk13L6iq1WVga/UAxnSrCvyCA
jyBhTPmeDiAldCKFG/pbPf65TZrxqxZ1vYZJURzBP52gaSQiDDiuvZ3h9TY8YWeq
sb0zT73zGWvx0hOz5VQhv66Qd8q6nw2A129Af6KSLxWJQ+OvNo7f9o5tLos6j2CY
5WxyJ9cB6aSu7gmWUfB5yDBDDaT4bUF4C2L7YxpXGXRWCxu9gmd1M2CeY7ARln+e
3ouA9ffJJYMRFtt73Jj9I6jWNsJ699i9gYvhOlYHpu8zmMj5bG2idxy40LacD3N0
RLNB7qHzjGv6WhKM05GfpdByY7ke81XShZwSahMcyVIfP2Cr/Gv1QKukrVTmlADj
MQWHtVU4xHbKmkNoHedihfg0G06VpjTvKPoobOyh07XRCtv2DKQF7DcN8162hFtw
+yhDhZl2za9KQYvjp8rVfpF2eurtgCKe3d9s2V2u5wQvvyfmPYul2YA137PDuBvL
Z3IQPB8Dc88cPG2OQ+dfryQcL4sE3LV/zNr5tMjf1KSnm9UzdZLckJlI40W73XRa
cXuEkQzDAfxLtIlE55oxkytFFC9qhqL5wbIrKYaMLqnM7SE4DT2NqWft2jnXa0wp
Ww1+gXx7GqcmLNg3nSbTkbG88hmkyi+ikcVpEnlglWP8rN3SXrErFHYvMTV5yMpm
AEzeWivufkTzLpevsQweZWAHbADiL/fJacErHzvyBDFdHmQRXM4gxZ5/kHdHA9uG
NSaJfcB+LiO78DkVFgld7bnUoN1l6anJMr0r356fab6v9QChQa36HFnUNMnAT82f
DwuHxUxaSmTW36K0nRZ1nDUTgms3nfaEXMKGLtMFwYDVlR7Jr9nnjkSwgbJvBRG7
j1yhgkWfEE466ULV5vy5Ssd3PHn74VC2q7XmRiC/4DH81Z4ICq1Q0nWOMeMQFIRK
R4aDfMTpnY3WJzxLtVEJzUi4zGhp8HZWSFOVvqbEil6gfAkAQZfYfHFkgs32n4Uv
XSmL2eSRhRtNStsqQU8xhfmk8hO6Zzsd1kw9iOCA1Jn0i/lCDYYx/dbnv2TktpJq
ToahthYYvGL3tFVdAfPnKC5KiM80kFQWEYZyTNiwEYUkXKSR8cnLaCcvXC3r5jsU
CbOFjxvfWxvI1aKCZv9gL+w6qMESjCxcV+QGkhvAgj8TmJT4uYeXRAdlufZrvV3k
aPEkn4JP0iRhihb/EBfSffA4+QhVRNrIMnq/xGYOO7nY3k9KD8Vocul/nVNMh0jU
chCrPv9EiGsgLhC0cMUsWjgupkTyhmBmT6E5fNi0JojsT+FGI94QSfAs99PFYkrW
KcHNdXsXDtK2y5TzYOWDrfwMXSLHpkXksBh8hUGjTjQa49c5pjqRZBdK2s12YyT9
e4YkHtEHTgcTsKSlSFsrOZnHO2eJfiuekZYXdnWxEH+CgpD+trdnlq33qn8ONH8p
VDP87XvbJ3FH8RXtvQ3kNVkFjaKYTBil387z7FW04SV/KLG2F8DQxZZ84pRVdTY5
dK0PxFguxcsVodmDKkeh0LHXCpJvtEPZi4jLBUUni97FzLiW5F+m/slHXFLpatlM
ln9mM6sHFmuG6J6FTrm4bkJy/PVc084N3RTVzLurX1FcPek2eb8sbuwgdwhDA3rc
rm3D6XUzEN6OnrO4GWIHGMFC1OaPiBra1a3ykhNCPrFVqxKsSMOQSdwNGZLs4yMI
BR/F/yb+Ylw6/Zwhv7UAY/kql9ewCkcSF3eNOqslc88RXRINDlAjqD0jxYlXTIHx
hZvGW+n9MhYrtMM741KOkuOJvnwwnKBKUh2fjboqrpn2BPTGn3NoUU04MXmDGcRb
uKTHWdjYs3g/Z9D/79MM6eKbivcOXECAj6ry939Igg5n9lkPs4cHTU9vFUq8cdGr
y69Bg2eTkyN43C5buwiI4UMzJV15szFZS4SpqQSQuJoi1Mov4eZ7dW/NB+VlGtFY
1WHogtGb9vGAXeGsAxOlc0Dt8GQOSWVBsA6+wVuITrDyCkbUT7zx1t3KwTMQ8YL7
D7wn01Wep1lZDeTx48C3PhSFuuH+kj4CA2KpxVT5SsDz2UEL2SB+FN9xbzffSx3M
cWxjn8lw/wYreZz/87gWyPXTWRZ8EO9t5DVYP+c+OfxWCDe7Ul0fphXfJhgXgZHU
srcMY1HitIj6LzPr/2zYebBtbujelHah+kyCuaNLowUCkAI8VxA6BVfm+jpaWRI3
ZHnu6yqOSDy+sbbIw04YFzD4f+Px4ZCmztVOqwmLxI9gY84F7MeD5fZy4oul4GQX
Neqyr/ioqcRe69jEwjovjm+5og4buh7G3XQMeCcmrtzP4JRqITPfhv/+1OIuWNYs
aOXFcQ42PzdhomdlQSBPMKqjs8jx/C4hu3t954SolrXweVB7ccTYL8Mkd01R0c9U
YW+hbD84fTGWVyxb9n/deMJhGsboiOE+e6FepXYB4e8tAIp/ppjctx7mVKKN/NTW
qMJnsU3k7M+0KZItu5FlvXh4lIsMzQkoc0CvOfMOZBCIgbgdoVie1uqzmGc7NIOv
rs9gP7TcC6Wc38knSW67oxbxbcFeyBA4JVqWyPPD5FZr4qYhFjz9lgevKJVC4csI
CWxYh5KL40VDgg6vPDEJ56gN/ukC3mxCgvpeeWG2Fu/OgMbsYCWOJuClgVb8jOis
etE1cHiqvIOK1Cq7HSjTxyKZgPAyDr1BUR4tAngahGFlQk1NwIIStgfJkiH+E/uT
pS0Ju0u08E9UU5jeZaAOKXmJcd70OyB0ZjAnK4m9JZ9txFHi2FKGu1tp3qx0y8gg
qluspR8jJIxmZFmoRmIL4x5Ewd47PCwwM9h03cOuGHmTDS9qyyk6lkGfiEs+AzJT
tYJxjHauvaV1u+beJeFlPX4ROlMEEYvDyxprQJWXEgEBd41NTMkQyjZfn5lIxifl
nbyFMlU7FrqGrFfy1gnYKb5Qow69VsSiQgNsVNB46dwBer+6nC1VGKonHkhfGh2B
bTfbVSC6ccgE5pRpjJQPru2mwamwDS1ce/ApxPf7ULii8GN7pwhph/UK04VMsdTX
TvoMblQXIl/9ah50Y0t5IE/IaTgmi0mf8lFeFM2mLQcf7RyYXf15rPzu/rzBdU2u
KWpVQMJyPSXBVP5IUtgiI9H1Hn0i77DtH31p8p53Lz4UWMx7cpY2ethK4N4WG9xU
/c1Ymbaxi4etcxYbvc6wi9XDRB37qd3C9ncIxyauTA/1b+jGAhba82qUUyqBjhZl
AHPwFxTIibP9g3Kz5PrZOlsKD0HYZ4Ed2Y1Jn8wShgcu6A44ZRv00N7VFD1uMV65
FCvV6GLDzbqQr6KBPtD+BmhVr47//eu0BfDhM+Uc2i7NVmfelx4WBi3xt8dB1UX2
dVP26ktnhwDchOu2Ogde3UVRQIj9Gpiw9FUkLY9pheFPEoVGE0Ld2s61ov/bFzC1
CM7ymF3Lp0dtFmv3Er6i7YkPKBy2ffV8iWJlK39htV0jTVYDHamF6GOjt2RS7h6D
O6y62PKiGHcdCzY6dXymmleLzmCwLG3EvLFwdBJ3dZIYrItdn5DUthWXyWol2UPn
4ohJzB1sC3lAB35UgN6IVppSWp/raUxN2gEAB+9SdUN4XDECCdYr7ofDXVZzDBJs
wsAS9mgwTouF8nm6aFf7UM6kxWIhS2qHd01gdgulZujF7OptRulvIr7WdNqiYYIG
IAjv+mMamcyKlDPTFXyDcHDA/36Q0Br1YO7DZjce0MR2pQplY908mu5rUU+NLCuh
4zc/spHX+e+i8toIGAvQjfQCAAky9bqv6fwlQ7qFJo9sPRrYvl16FHcNIcANqbw1
cmuGcnqCi8CMaeY2nuDOWuh6PN/Li2q3siwelg8mfO8/LnCDOyuz8u3z6y6e/NPe
LzJ/5+QzxoX3/LTiP0vFbRDQmi9KFR6fA65DJBHoiYawtdbkywTXIEVtUZVBX4XJ
WjTgvBFqjVMtFzwVvYxZn2TGZvk/HFZb2KfSrTQTMyjGoMKh8zdVbEXHGmZXb8B4
zdFvpgDOdRO7GGH1kdodS0RzJisRRJhKhpZrIHioHoaQGd3IChyKjfALmyYppRhQ
tX6Ol0X5el+14ouKI4yn3prXUWPRVGbCKXsHkgJERi7Sk4stmITkPBA+20+GLIH/
N/4hzBbvCDoHM8JHbfLm2h4qj/k9g9iEad7BAXfVoYHJBLhoxul5x+DoJ7Jxa7wE
QEHVZMkOLCvn24mcSudPNJb+lJFyp36mIgJ3zyzjZ0CDxhWPB8HgQ7gjD9Itkr5v
i3YymaSm97IuKFT5VgS1KLPj77b0QfzL699sbcGNFYHf0g2atlA0JgWDsgUq7jpJ
wVC/qdJ33YOBxwehWOQDpuehAacezgZbjxF83xz0omS3dMvo4i3hNm8V9pr5F4h4
S6bnRK4ggzpz9qYXGF3REFXLbx/Ygf4fJ9vQjAMrf0HJGG+G7NgSo62VME9P2Lgx
0P5FTM+aauj3POiwZ6lRoVo2MGAewseH1KGtCec7gx5XizssTWb4aPj7eko6ey5H
/lEu/cqGG69bRef7AQ8lVEV6TjuTRT4UV9xppl9ZXdYfyvkgTw6zCTOpcVy7/KAc
wUmy8KtwW1bT4v+6+AQiQDEsJlesLoFjLOXXUCuls8gPRn04UHch62lG1H4TBFxC
NklVf95RHPvmXAQs32LFxm2zztd/QqlArI8asV7m1xzAQrXpg2N6tvKneHTaW3dZ
xyOX65VlLJVw2y5NRVDPeIYsd/gXSMcy3zDdPlhNt6woKzcRk9oXKan9pD9Iynz2
k3wRvQAIoUSdU/R8vSsxK7+zzM88ty5dQ8TJRAOpf1lzPsjcqRwiSUscfph26Zeb
xktk7NzEVkjzD+F+D33qvrONZrtYVqFuI2Y6iHJBGP4jz1BwMgwMpqehJei8YD/n
0Ls+kFswtJbryFCqKwuXPDWGGTwdMJEORt9P9Wm433qO/ZaoXm3/LBbYJ58/FDQR
6h/R8nwnOhvAflx/+QosJWcsO7wr+eHZRPNbm1eB144Dlk5kZmXeFOBmUF0lmOCG
fhmxrVcDgkbc+axLLFppS05ePBbk5khPpXUTSa70BafL6XLZWmRsQL32K7yr9egv
bTn0YWotiqPZ0XxsOoLtPGgTU6BQMT5QCF9CxmPF3NF0xt7d7uTTqT4FNnElN8lC
l3t/lLcp19CB+LaMVZWJg2at98ueUwlFitv2iytD376bJeD+F4vo+HYwOv/SPrW+
SkW36vp8MBFRFl21EdiNnmrP7prH9/rx8aAsMPs/CN0uUfsD80ZVjfmwgyCNK1rq
Y+yIfVw4lLbhFg2bdu5b8YIiy0WbEoSILutoYCaxMrWPWfoJDW8x4rn7Tc8n49ub
A7Eui0v8Fa4So25Qe8qBRugc5kuf87hF7Lo5NNdQC6xLlNgoj1wNhLrWzoDGp7xj
XFHwMukAs2zoTosyXFMI5CptB/OU1SmevFzjFzzMQ8+lBh4XJUWT6jUULHQ0LXpV
WP1tIhC1fcHhLXegMZNZ6X1x4835ttRagBeoxIbcfb2jgLzUXemSFQhcXoRpXPsF
vUN/G3KT6WN8Le/jpc7TS+iw1NTx8Uk2497Fb52wUWZDf6VH78CdZYVcRHFISjW/
0LexFMYZGXEgY07aJC5FXjDd0CsexUArkvWlpiwezf4ftJSbx/Y6tvzSjVdwWzgb
rEGDHw2Jy4Dr5UnYwiJVv6c5Y0Gx1ju7fqpq95kY5nTWtLoDq8j+K3I3vSUc7KQc
P+2pAVukNbE0DBFI0KY/XPUTqaqtv+PY6nCm3hFOjUs4hmxk6fWepAHt8jqlsSk1
YCDL78jeJkaD2e4Nk5LdR4tZ/10ZALBup1LvIkMviun1DnQxaZzDI0PljqlVsELE
0ZpL0kWm7xJQE/VZUq7MnkcG20mfsF1QqK/s+1SrTcErbyjrSDzZUI5NGVYWXs+j
9WL0GkalRDR5+ym892nVUoJIXiIbJIDmdgCKko3OJ7+RGKbCq9Uovm/LeopUMmGp
Q7/kfABB3Iw4EAnE8IGFDgaLMJsVuGVUbl8u3hChlQeLVjKvhdxQ1sc2WIpLOgvb
LxVwP3Z6hnQlwR2rWskDPwPKfRmuGC9bisRhdB+J9JwXMaku8POyXIQK0CnUdHRF
37S0K3KTiloxHs5C2LDOuc3E3YrwjiJwl0Ur0lWJqN1W9Mea12iwGL7MPZ5a6sQD
BlG0eg5fv77jrnBOxL2N7HBwNuKqYBL32H9hf3ITBGRBrzQVP16ZVmD1uibffFLJ
aY9pBre8UoEctvAAQ5X/l0wG173J9l2LZseSKCSuc2PnCMbA8HjIf1wwtfzfbDJc
W7nSNELSyNLkx/2oJisnvI/bDDSDGOZRaNmmR5Q6qD8mVB91YRThYqOY463Inzbs
sWyeMX44B9XOKSzkYpB6EsBnoFKgoG15LGCKOZELY5fqNe+QUl28CXwcTggIXozS
CRCIj76E9yMTohAFKetMPkflWeSSaz+Mpoq3uIbQ9g2npGO6KSJq4srkN9wT3WmX
NLz1o6kCQNGWaiQ3VkObHJNRRzZQUq5NJuWFEiQILOZAn1eu15vB/o87+/9DwUUe
XKjNeC+PDPo59WZlqAd4176Qh7mhdp9D/hqaqBQBhfOea+F+6yy1ZvYwuy0NNJ1Q
4805esMuNMLqyxLg/nk6CU9134QRQ9Hr9bt7OPOvq0K+2591LsY/n8R730gGlIew
bAgCBxLl/OMzH1cer2Y3Pd/xEcKmoe30cDA9vQu53KxOLWcZsioYTlgSH/Gf/TJG
NpIIyefi6wjNJPZTO1u/TP7UG55Riv6/LBfLFvdkJ1Vp7AcdTMencBflw0bkeTW7
zEpzUPRRRpW1s1F3VcDqWL1yHl7TP69XmVf98T6ksUa7raxHLU4ncBO02JxO8Qrt
aSn8mtD/rvkvgIjO9MmMVEJfBPdPMFeGJimbtW3elMceaJM4XWPNp9aojHVfHofX
D33vcUsvS4hBxEG6i+Z6alX05ucF2F+w2Nf12m6U8wLQVwiRXWsCTEK4UFcS1Ccz
3S05UJtTOWuy1QmbwsINokjsjp61EZDyPBof5VMHKpitSF/iSPEgVZs/+Fr7z3ds
MBlQJITwjzpHVqRrsiBs6BM/gjaCODSdD+zDnXKE7CtvSWzbEM9TxNS2qjpY6zls
5IoojbYb0WmXZjY8JZUezjcXpCWKOD1CxDq5Sjr9I6axpDUvwhZ8j3z+QtNmZuMg
oX5A8gD5a5icujZ8si7xSfMTnUjhy9ijQUVHfqUWCBApI2S6aClDuynCqDklPwEo
eIvv/OwpYHZ9mSE9PHgUqyZuhtMxDtwXy8k1ML6iQQMEs+ylVvKrr73r4lXc5NQQ
Z5XgQgIZnPUNsKFsIigueHhWkcLFd4Fnzr+AqA1C+cLgesC2jKeeF3VoirYF279W
Her0TA0PZgx/GMu5wUXXQqv/Y+ifBm2g8gI4AUlaHBbIv80MoJiUpry+AMuZ9fo9
PbUTpZnjAPwq1X6Z3HDKmOBFaXM1sFmPTdD9QEhOJcYMXtjTt2a1kLcmzeUJf1ZM
JX8ZVSbFJKiEdto+XJed7+QWEkr1FQ3PPZljft7hfI8REKgiKHNTJFe0+izxAEKb
7tsgCTe5DJHMKCalnqOR42hYh/qeQibEp7W8OX+2e8waWnqH9xUaU11s/PLRRxJD
QvKbxr5uYArNfIhNHQSEh9wpT0+4EmrnJL8WBkBn1WAKuLBbCQbulDt9fDFVdvg+
ECrBVtf1ZYelS2wFL3RpCtzbPY5y7aLfqquA9ITNcND/qt46TrAvKQAHMmEMPdvE
MBOIg7x/LxQ+Lx5T1eUYxIzfd++fNkmcg3Ds+WvBu7g7IMci6MWWZiYN+Plm+CHN
34YRxt5Mn98tIl/OKSXDQOjI+1uGVNZZtOgKeNF/iqRmIwGYDGW1XrnQnUuvwioM
+6NKZ6ESPenkt3pSmDw1tZyl5fS4sApNc4rO9ku3jPKPfbm8TzHE7fgHBKhSVd2k
f5YZdSwbrq208BA/sIixkU4LWDzSUW227vsAoED3PjtFA844T8UhK4pJyG9QoCjj
/H+F0HsbDjxdeBOMd8qvk7LVCk0DOL+ns4LpctWwi6aQXCOp9fDi9F4f7V3bKhWn
hyNUVhfvvhNJxrQpxtEP4sLW96x9p/sP/60YVCpm9bDj9jt5HZ9VY/hJKF+XQnUG
tB5JJmXr5BKdv3UnLsFvCqvOTMZX9sL0gaQUSTR54y3Vs4iS1BdIiu31pMSNOlpX
0XHoM3g5wcV9VnqqCQakvb8KV1gasIsBT2fmYJgdb/ZilA8GEma9/N6CJmWnNuvb
HRDzw819/uV3Nu7WPBEcjNGd79YhPQL/+LZVuV0adJSnFG7gxRSArUDj2jHx2ECF
kbILaiEU+XB5iGe1CS3q8YnPCeQbl+2Q9WYknPFZiggFOUlFoUoOl1Te84lrK9qJ
S+zMLRGiNH1Hs1xa+Me00AO9trkkmEYrLQbe1yd6YWa0qnJPNZB6vm+HO3012dUn
pcxftnZxw47LB52GkEJ5Y9BlOKxK62tYuHXC/bQrPM/GlM68M1AqbLLconxf9rzc
JetIOvfRKHvoBFBseETV9xcxSwLmQEv8cxqDNFCNclRhDFhd0Z4L3cSEGLWCtaQ3
SCbFVgGSDGNGT5dNvDyP5dd/LV+8hyNWzLhxKfNNzp9Wk7KqtZ3ePTRT5DDdYg7m
EJ5j5hR+RyRS9GTeSz76BzEnx34cWmCsaRfx9IsSziYSRMHeAQLUu77Q5LAmPFSG
Kkyp/rgYVbcKkvtUf5xQnl1uP7whWgV2h7FhjQdCz2ftRaqejhKlg3rnenz8Jta/
DqZojaudIrYhlWUqqV8TUtYHBUovhm79zokAqq2Ls0IITjycZ5O3KqLkLmSyORew
QRDl7M3lN9ucAqB00vDoqXboPwK8h48SQ1TzWuzQwX5QlkPrZTjXfaUduyOA1QND
2KBrFQQRruIN8jPFMmukRQ4e/5zEz+7pXNWg7f2hgEx9aullRWxlJEsajorUKpoz
np+jt4t+jxbZLsXNPnhf/kXWmUfqX/Eo/xNCgNEQm10PzzsQ3g97Z7u+8U0pATG6
2nkYc6/KZ9HjD7izeK6Cl+g+vFp3BVnAVcdnFDNab29b7fRE9lX/3Wzr+PNZLwWz
DdrktvVyFT7ImeKh1HS+qW/miQU8CUyPVhdN2qd9NfN6TRo7CWXBi8np2efhMGEW
AyHp6daxdRxejFqCeeImVOwMAXogJpuZmPcR1T7K/bf2n3KTC3XOyhuubVD5cN22
4AsEM2+odhDxblilOq+w6f+CdNCKuMW92bbHgoxQYi5Rh4ig6VL42BLIUPjk5Wgx
juKEhn7KDoa5B1n0FIIuYXl6+V//Ajdhvj0iRnfzIYgr5/HigDKyDsZAeQeOByXq
XZIWF7Pb8MHIUDapb6FgOQa+1tbLZjbH65CYUu5ciA9RF6AxthYoWbsEQY5HVP5z
c5IOjLWq98mXdpEnmGy1+yV1W9RFVY5qTttb0+W1M8p9Uhqffnb/xEv0lPMY6iSc
FOkg1wnu/gONTDA1yfDKWEa+nckwyzAQwruswBYoGBFciH/pmmHQR2AqH/hNfSUg
IKAlBqtOFAqEDTLa8mjd3eP4RUXjqQNxI8HNidGiC163lBzYHGYevG3bpPj1nJj8
c0r96qrMVl1E+KbedaTfkdQYEVOorl+06btG64kPGTiB+E4KYycZ0k00FLk4y3OW
GTatBbWKevAeW4ppaZWSyqMhAde7okjNPBJRhC7ofMrE3OsUF36JFJgHJ7DVcmn/
KvqBCOkt88ANURGMlGVuucHJ12bXW7v97jtAUgjL2BU6UHkudg40oW8tkIvmg636
8VSVocr5n116TB2I5yHzOt/eshbCinFQGfCqAeVYuhQhKt0DOLCBKZgQln2zME+X
kg9c0CqHllqn8xmAgab4rmzPMEeyznZvMuPMSYGKciHs5gBmmOGoSttwnA9TBejV
KxngDigPIT2h4O9LcjwsQCws5mbYdYLdeeAFNZdJWyzaJ9VmHU2YvQskEVZ4Q1kf
u+RTqvHjgYb12z+/lJSOhNOQQGD2Zvv3bxlZIdYIN/yZ6cOqQFqIhg4iYWk97k6m
Dq2p2IkkykbyfblvIiLlqaDu2wwrltQIY0tQj4xss2U6pQHOPM0qXKlndpDQQADb
zWybiEs5AwX+lzqO6kFC+iFHAWptYYYtNodMVFpOxl1cOkYZ6sPhiXAp7WeUeAHO
DLrYX5G6K3e26NI758ggNFr3mNPwR6mQo+qNqBoxy//sNPis5syBhRKybgSktXZD
HGhkhmzP7QJXLpKMREe6fS657JO7XtlD02HLbQMSeCBo+k7+dHq8rab/iCSpqw7d
hCqAjTOGCnr/JIKWkwJgMpunV3QC7F4a4/3Fo0+TKUzkHUMcS59ycTh07rUDyhck
H8LZ/oKo9vfwfmoXYTmq8DxExd6bjstrr3xe/CmxEm8cdGk7eAQDbz4/f+Tnyn2V
cjABJeS9X0LQRbpPpnOyUwSSGNGpLJ2KPCctLi3gbf8ZrtgGMGs+IzCjohyiC1x9
ipUqk9Vx2wvper/n8sdfuNqLKI2ByOanV1LiLTPhyoLsAvR2ONe3aMq/NQR8HE6e
cxoRHgn4Ae18yY6peXuwzexLe4glCUqI4Yh4C+u+zn3YGyPIkdj98X/oVwT0uwvF
7SHU7225g2/BMmX65TI5PS1L7jMpqgMPFZrViZ+rMseoXmzQKtTgCDcuwXMnOSfV
TVZJWDOAU/NGyY/ijI0xuhO3ZYuqJbRwR7InUuXS5fxgn9a2Tmj9/wK5fatOPJf6
jBOV1hEjMpOt90X+kpX1PSRgLb0QiC4YhKbX05kCZLmsUWqF0aXv2pamQ2L5SMMu
7IfNBQT6BJI31FxthcQVMjKApvQrThujkXlyauJGlkzqsG9p+EUAnxsm5p+yhuS7
p9z0pkN+Io/RfgCnAkRj9EI/d3IomVK7LOPE/KiwhKqeZsnlRGiLn+lsQGFt8/Dg
7fJGZYbBENqlyZMc3BSqMB3ebMN4Tkt+rHV8IFVPZ6gy2WYq+YKhQfCsCOtoZcE2
BxKeQjESODP7Ani18+wT1O1Lb56ROda+lB7y1WbfHvAs6l6qnzcrVd+t6exu9dz8
/LQMDUNJCSvUwJWubbP9LZ9+OA0Gd/UG6JPVDXYDVTkEuyLtzY/ebK//4ZwN5Az2
753sX6T61Vmvwi98bsveW6Eo/dAmcSqEgG/nt9NDjTjT42YK9OhGFydvBF0vlhJ9
EjbmHJKAuLtsBF42HowZFLIDdxl8XRxfIxr7pm3PI2YdXpHMgDOBXPoFeePWlSlN
xxjFH9KSQRSJPmLpwIaDGqXslKSsa4QFmuWnA24dRrVmpLYPyfOBPQAunkgpMeu2
yUkqcIs6j8RMC4Re/E24rSlx/hxsHp9qQqGiOS0ZZ1hjSlu5n6290bMc0Pn4uGzg
ERJ8K8rmzFyMt4RAE5Z2KRG5dBQNUPRZGQlV/Bbjo5CgRykxBeUR6ti1SB2ZAcsk
+beJRPvceBORU+B6ORD9aG5zgJKc95qgoJ/TN3tJ7LcyISb6OHgEnU7JBwrNquy4
odfInOFqR+sfPg1ZmlN/+/Gv4obpAyn+ZMSZE50zAojq2lFOvqPcwYznmVS67Nk1
FHbUUVj1wT6znpcPwZ4s6Q6yV/KM2j7BscAPNRFIwO9NJ09weMAsF+Ekmnn8K5QV
S3LiGSerw1xneF4Dd916q0q6WuV9rVExB6I8Lg9aE2lL0KdFE/4bE/6wOHFmvZKS
QwKRjlAAPfmi2OivN/4Sj8CaPSpDcHcQ/+2oaf4y1nZ5JMyaeJ8vlFimc9DQQ+Dg
brgArkP0DLCdRcwQvWp8ljXG2bXmoUow0i6Dwt7MU6EFB7TmtVe+zPGWmg58ZaRb
6J4rLPrPffuf5BaYleiKin4MrwEt5jN5j7TI73XOx900mpijiB9J6aqTtc56vh3F
YyKffQ6II/P3hTwI7fmwL6aIKMgmJAtnOBx+hMDUuRKRR8BC+3wAR6AGxnss2Hei
HNi0w+02b8iAn/l47dO2QmPlym08ye6VWDjlM1/kgCr2OHfZ5rSDQfePeypFe79K
YET/hbGUVbgTCEb3ZW5mapRK/Yh+CzoDYgWERhKVoXsqg7Spvt89Enbyp/eu3ykn
nImqd1aK3SJrnZWy0AgOTUg5hT5Xmk+PY//+9SSekH9Llrs5S+Mc5wHrAbwJkPiS
IGyjB7NLMLaH2NLFodGN7ab+iaExLKwACstE20atsV4vhWx9YM78ypL6ODZaxMZU
kUPnFCzdlKx2IU+lMfM7RVGIOncXACdeHOCZG5D2p/rZGPnD1Pa27c/FHhRPlqdv
hSDc+Xm5+DLZxbMYhdDypzNqZ62a2OM4GCnz2VQMXWAwGOwahhWWae4SkDZ9/LHF
4OV4dMGk2fYObHTEQC0xNq4+AWNx7d32zxb1QcpBfWA7798LUmIYMZV1srjZY/dO
vyMrhx4WtgLRetOHFIkARMyY23UQi0HpHHv+PtoNgop5WybiZPOxj0Yf/WRTVMN8
1QPQBm2LXWCPxyuqaBICQd//0AYwPKgyJI62VTeRhUJ73/+v2JcyDxdwHX6vwl5j
NiMjPABrFkvDn/92pYgQlI5T9TAqBxftRJpuQ05NZxT5A5+3VJ4XzUiN640cdl+G
L6hMmPjmZuHblcofhMBBSG0UzJXptBHrYGxEMeDtbCDDNcv1EecTyiJr+5fsYjfn
RtXf8/E05+CDUJOchIC10XRDo5xeuyMy0imk3+LMr1i5Q9vXnG4eF2WEMoPAaDri
/UdRm9IqmmN0S/2RzzIGfeQGEdlcDY6kryIh1jwqIJwnY8WGzzvkEG5sHPo2h7+7
vSwdTTLrHVOLI0FA1wV6GIQkG7+rZkwZHpi0AWocjHUqS71pQfvbL2XnSH5sr9RQ
s3XCPUz7YTxSgNe1LtCYrveNORiRfesmV0qvXXzXhJ7hQk7drAstfSz2Ry7xvpZq
RMNkzl88b8lcm9MPRe76XvFA8hnoLvAIwAkkmYKpD1YrS0bln8BpxJGBX7IH6vgR
X3zXT0DZAWiSjSEDflA3uA908w3qpJamjSF/pnFf19G9pxLZ1UOcfXVBPbVhOewJ
G1eI09fM3ARItJrvCcfTbseip9ivt6HCxyGGYh+AddRKVsYX1QXob1jBhArT9F+R
i8uwiAnd25oNIBH9Z0nGdVNd5HQ5Xs7m/YGaAj8mG+DMgJmee//1EL0DHfQRtehH
Cy/dpII7gaTg9xZmbUGgMdsZkMaaXmCk94/DbBd7MEGkwmZkDQdz+ZmMvNfvCEfP
ZH6d6GV7QtQ6PayvLyyCMUR7dCrgaiZga/giuCFv+gR9Lrw40kRr7AxgBfW5yxpn
wZEhU75rd8vVciBu3nxubKwOcXSg+uDkHNUAqp50f7POilWCWa8PTmfZBZgusD7S
wVFNGhwIY8z81ZJbgru0vB4QaXkde+n9CyRHqsJbPBuHGjF9B2DxjfZL+TTh53ZK
QkaSfCOpQYvaTRuv90WA8AeQbrt4UuF5uRj9YSEvWNDmo6PHfrXCVt/OxcLMn1u5
s0VMaFwzYALiq4rOUWIhNRhJOnrNr2RmdfsPIUr1J8JxqwUFdSrnh1xI0I/s3j/j
XuLHnUuBXEbYfN4vkeCBuY5BCpNnm/XG8nEpWNTWHiLhOweE3bRQisQwsMFfvgxD
zXXWrvITCZDAL4H7MvjMfMvyuK8BQhuaLSFiLsbg6hb1gBz5qkErVQ+MGWAuTCr9
Q+7ag+l/gOh0xruAu0NQAsQasqSznMppcFkA+wkVCgssySelUxjpC4Wm0LZxNx7X
RjOrHgo7QUCpDPF1lcPT9uKVX4ZH5YDax2eHN3wgrw0Bvsie2EK7sAMe9MzDKeBS
SAFeQGcU2DDLVfYcxB69wD2o9a59zf7RN5gqTIsGi/upJEzRwnLG6gqDjeMXqWHI
G9ihFRlWhWJD8hGDIcrCfapftwI32QEtzv7KwwK58sG2lkKL+vKuOs8CczQ3Qmwl
JHkdgwOLaEvv7PoXzfe8QGRfU2VctmQcDLsYjcnw61MOZLigEMwpjdvfP6v7tx+4
xQPCqY1ftxfpQ7n8O4/2ntSd/tFMHZcZUyBlT160F0F1Nffb9JFYLGTJEpt2bjnR
66g8OogcV7kCe87pS2Ajkw+q6TfJo8RExB7XywWAJJsJUXax2iyz/5s1mrtWThpm
9F+LvHeuME1JAwUcETf+Vb+pv57QKuzTeh3Bdxzpt7ech6GoxRu+ORf1CthcqVD0
kSB+XBnaRzsYUSEKmxHCq1rqe/fx8c2Jr6MBQcXL145qDnqhcb1VApgfniw+ht+w
rSl7kzKDJPlDN8QIUUK+fhUkjupWTlFy2StHtnLsFncI7AG+o1jenHXaDqdiTIBB
WmUWWcWVmxjoVdPgZ0Jdulb+V33z782SvZm+PXDOMFGBMquuGc7aA6pY89onNh1I
5DkwpbypCUQkhOIFF1ncG/l/OCN1obpbrc0WMaTW42dPhOQkLigpYrDeCuCDSVxH
NctWjMWhm21+VXrQqkrGdAvJEQoye1VQaLQlOx3iRWZcmh0HtgA1ysWQXkWDsKi0
Oc0SV0+fcpII/Fp+SoxtUPHR3O5NAcSyS6RM4fbJGQKrHgB+EJXNpS/G+8x97rs2
EW+VBzazyKtdeqx4uzEUaoB+Hx3oofzLtO/sDpLxh62wL1TfHTnANHNoFx5KTsE9
zFLIJFrBkrR11nCI/UqR9tphBa5Rd9NAv4fot+EC4VFUtCtgoEgJUwL+z3TyMwtv
sdYmOOAH97e4lzWKqrl0UWJJ8rs0XH/pe1EsPDtJx0qnI8Z10bDrfIiakifPjLUT
KZbSOgPF1iXxfwYLkIYCbGplEHWk4P4W2CO9ykwdyEizwmcSo+Hkaa8tInPow9+/
jnlZMpS0YKPnNWf1bb7otVnNWfr1GnEacVGeLduMaxjR5aMvTc83LL0Sn5Jj1YkN
QxFf3nST4TO0wT4d6RFKwLpxEOMmrpO93gxfvEyPMnWWiePFA+Uj1C2JMVQjbanu
k8iSKwMc9zhDJWzNmEJ9USToH18Hlmw5qmNyS3FY1g2okdNaLDoHTkviec0sauSn
DivDV2Q6I9mY7ZkPofO6uNBMlhPpnEjuBUDzUPDA/bcKp35d8zVLdQT90T9dlku3
MLb3SIrqiwBMSqCLlu6kXN+dJhPF6aA1H/mHs1sjvty+rbzxuLPfbCAhI1KA2ATI
5mtctN7A77doGmmVDYLJS7s6+57JdGn6lX7K9VbIRIWsvcwhiCk47NZylg6qd1mn
qgk/duztcVSSv38DOL9Dnbcryyv3+mGzplTFNyjAIWmLc1mQ3BxJKqHI9+dg/+pa
lWcFHobExodUkWJ/6STspqDuUZS0o/OjYjC2uJHQepencyBSPH9PCA17c5tVGQ0a
VHrvaxWAZO9vpLuqiU6KaqGMs6DbNhcpCP4+iuAlsTOw5l7+dvgE4dU/KpAUS9mk
GHk6WbViZyis/s/FkEKvKkuHvmP/yVNQ0waG1aCc/DC4XAYPYD29xTGDxCZGwIcZ
YXCBYQXeMbbHCe9+kLlhn3vx00y9JuH85EYI8JdsQawH0BjRNLY6PtyUUVRT0/C4
lWse0vCUrPj0ffQxAsabJygMt01dwsPidB5JNmHWWdewBIlDfb9Mbu7uLoaI68oh
YU8TXgrN87teytgWuvyxSZcpmTznjZYC68Zyty1cIDSf54XU6IgRLOSa+Wb4iTsq
OggmfH3ptk+r5C064WZTBxfO3sPrftAjCst1mLdbgrolPS4BCaX9GX6lSuiMVD5b
GFQZq/4noicuponTsCt1ylnc22JiAAMXoeB/GZJt+/dgH9AuGZIeLRgNZL/eIdaW
ssjOrlaFs67NTm2DaY/N+9EfMvLiDi0BioOJ2HHEstVPOWnzP4SY8lurGXDbMXwn
Idv5kIlHS0JzZAJ8Io/pwl9NdY9M+CwWfePrz46RCMMsmuTuSElfc629mo2J15Ht
fOJPEELpjgeyTC6iNJYv9VqLj6kzlc9OLvZSe8NuErYcWpCC/VsfbRe8lo9iMpAL
EOxfXij0suaGxX8MbovujXmZWCX7kmlZkWkK55WFeBfz+oJwDWd0nhM3SxiuCD7P
4llvpIUleUcPyC6J0F8FZkZAHuF+b/8brwIZMy8GKo549IE1BAoO6e3VtcVOQ0gZ
CcvVxHy576kiLWQISvxAkNB3DHVjayLV+KwA1h1mjcXKY1UbrryLLs/v7KXdkzR9
NtMay1eBdvQWZCtoHcRukZI7KSXRjiPX8h1YNr+C6K7Y7pzWpkCLNmjRu+Ct37du
64+3orU6YqTr8H+yTecePEcv+kY1MzzsleBcDD395h9XYjz/v2BYr8+KR7UkfoWn
8BNpO+ClECdPtXTX08ekV25XrRbpgMv3hRB6+zYX7wrSy0rKfcmTBfpSmhuxiI1R
Vonnd9fIN/IsV6RQs8H0mCnSH4R/obU5chzj7CpQHkXmou/CuOIWORtki25sMwZY
6hPvb/Sp9HIh5+L5+E07wa361aaOrfmDUfoDtpL5bGWC6xo6toFVriRQK9/gFZVu
1a36SY9w8aMheiSPTsXdIg/FsTbQTqCaO8dV7nWHIDDnavqTb6sSXbdpVX+V+FTC
t9J0VqIokB92ohk6W3a0HnwuCwiay1n5gjZuZw3rQknBqOZfbiJgkefL38q6zOYv
5ijaW7Ux2ryyv/nxysvn1jiz6TdOu+G0q3Roz9G8Cd7gFiy+CzXMAYulYUWlQOVn
DOSDwu24WYhr03QZJbqctI1KA6cypZ2XGwxNYf54RoUF4AhIf6QEYpxMFOkueM/r
X5L3B71x2xj7DQRDMG6RwskLhf67f+KOt2a/SlpMemsFerqQR3+BSLmVH7wYkrJU
TF3Lvg14VGBDVZtsHSORK5wuB+JmQWbOe+zzM2eGpyySqXIAq3S3wKVS2DN7BHO5
lEDLqPlY7bkHAjrA3+qxQQLYoBO1AumGKWsnFD3hklUU07kerpSqFoa16qM/oN7f
9Jtb0bR7wrNDYvgb77cs8oeau1sCiw9nNlduVqLmTLTG3qh4wEDAfMb18Px8WqCI
YQofd3Km1uzCCFDayLiJSzQm6GTc22/3V/LuDhtPS8z9nyBKRfzgNdqL5x99bHPF
vQL7PI6Q6HBGzL11Oz6ParEe5hxGiLo+1PJB/BXmodPmqp7z5LAiT7idDKN1nNQW
hBpLMh6xGrhuLEDAg64IMJjTNGIChdIMVleJWSiNKajtjabXKsaoVotAUqD9S9Ef
GWqZc5cLLZrMsmQ4U1p8zL+t/OGwD3Hq9aEt/kEcvRArifsYeBhu0mhjeuQsC94J
wCVVl9bve3168WHt1xwSEgKUaht+wS+aBNmatsS9/L7sFBlIAac7lPtBpA4+tHrJ
FEDj4NI1O1vZSFKTNIa+QzhoQeT0j8M8zthm5oC9gLCWp2jl34H1ZHM/kL7G1y8v
TZjHR6VjUKTghT6NQJKpUHoTvrPdloIikPRpA5AXsVJDK9irAWW1EKEMS5nrRxxO
65/vicTG5zU2ZId5wGmxqCsLtU5GjDKvNr4fqyS+ytB3m4tsr690Dw7pzoOgWJPD
YimwqqayJSQfRwYwC04pWm6Gh5rTBYp+9IXI8ZFZPEG3cufoXK+eUzfeEdyeV53+
aIgFH0FSpQqIno2caTBvIzvuY8gPrHD3PcnkO0zrorfmamrX4A36k14daqPWw0Pi
v85w/BLqw8kND9RdKcoYLQc/3xG+fDdaE74pPleObfJy2d7vJztaSMBv1TbUpcK5
wUY4EMvOoGU+JwmlG42zdWIn37/w6UtKuizjsaA8hpLkwNg596aza0PQTTyklaRQ
Mz8id0157rHPl+m5Bd3gJ4YW4AtLbv1+iQm9BeoRc7sh9jGKPFRM0qHr8BI80lwz
F0TYtrlU8kEdEJHkW7BiSB9ditewUBmpvVDEltrr0C7WneaDn455EI3izw1y+rtr
3SBFX+SsvJckany3wmMHYBUkwq4gtcXd8uHas3b+APewytnFWegbBeCOSF+OJ6Ue
h1OfjmGW9XFFdvhW72x46d1EKy2SAnPKCwWmIpxXjGHu5rFBfOqzE/PATfD/fibO
oJ9mFMo+rzHEkLJG05mqLPwWK5XICKbBnr86YRjw+KN6/xzdOE3rDI78Wm4shYgJ
SZxEXl4FLOgjMwBxkGWBobGiReBrqKP/q0K4NE8ajL9AekMcKh3rwktkLu1lSV2q
DipC8Mec/gqvqcPpo3OXrqelPhJMwmIJAgTNPb40mhHK4u4II3tU3k6ExGJx4Y5y
OU7c1NjIFCFLHhbj2hz31MysyIyBiEKxWi2rzZ95uh3leT/a/HqWXMg2Q9M0QL3e
fEH2ki6Bf51YLEMMtYFWRvAmNOgyLJPyG68yTcXiVajJ3d1YWvcwaYKgZ04k4wkm
Ea53mGIVw8bMOoQ3joXyu9CU0bqZHweqfOuz+DxD5W9V2v52W6OTYgkgvOBx+06V
e24rUB5zhUDeKIlhr/X2K/KOo8gNoUA1UXiZxy9tu71iBySG8+69a0GPHS2HZN6s
4KpK64F/5SYOazOotJv25VIxC0ZExo449noVdZ2KJ4w2POfQjrMsGFHXFmoIcBxh
csfW3jD1NWUlITiPi4HiXd5EDP821Fm4WCc25IIGu3yj42YxW7BKAHBH8EF4d90W
gYE5MvkgazS+WsiQhjocsGcaSbDdweM0E/jJjK5R4bn/0f5zumlSqNgE7Ws+gOr9
HmGsoEE5CPhN3NeiRLTiPGPH9t+1Q2ScHONfOpn6CKMJcMPzqCpM3CCahZWxqbIs
7hxkPJDB9yRUxTfRQbyygFKaBzyXdQ7KK2KYTz1IXV84IUZya01aLrI1BMEOppzl
coD8D5LbNAAZrUvDfR5PW0mTC2/fSpeUlkIbiISCBi8w2tfXsLlDOSdDhaAcBGw0
3WBQtWpcyE5cL6QbVxiAIiwPHEXBr04wgkV+XLWb8M1Ln2bQJ1r/3PMhBYlq1UVz
stKJaKDezdToUcDuHL5wDk77nrmxBWRfAcf7ada8eDJrwp4jkXh/JmCXWsSsD4Ob
OQ/CIZFXQNzZykWcVkG/2QPRwmgilGYWVB9VnLiDqPMrjtCnLGZ7WxFKWX1DNmUE
WQRayiH737utwpbyzVzKx2VkGULeS3Z9jzrsoTsT1iLN3HwNmn+mRT+ClZvoqRXK
zKwsv1uVS8zyDTpC6uJ//M/KYLU80AfWWL78VexIL0SlG/jSEizaLfw0/dTL5Htu
BA565ijc3QQB/zgupEaCbmfYYZ0d19kUxqM/Xb+LqK9/MJVLaG/CwN3Qe9RVFCkE
vmnmRv+jJ7Vjxqy3Jrq/xhXIQNoz1xI9daG21zAMCzVinjf9+B6Clort4z/+53T8
k5XE/Tsno3JJYP4vCFMNDOYCTFjxmA/7N70IQiGcwT4TKZdBRk7DCiZJ12OxUF/M
TlqvdxwTZati4hlvbMXktu3O0VPpwUXMfv8b7DFGBtxTwpjF2fO2zDZbIcV8Tcka
MzlXBecIf4SG4x/6mVEiX58aBRRnLfdFfWCrjYxSF+4AGv6nyjAdRyHv01hFbL2k
a3/pZH10wVL5GkCpmzwNd4JdNfw8a3sg59Djj4cLLRjzDsyeWELdnmP3meXQXyM7
jaUFfFpvf0J+86t9Zi+ilp7edqtC/d9trLo5nUEspxgACszWVtzY5JcWPfkbpbgh
gu0hnydYRsyJqe6xEJhuQiww6/ePHKikK14WasOTg/AWbkBp7OhDwGRl8z0jL9MW
rZqLblxtyY46AJvU01M49tFH1ekOy8sHxAOpM27o/Ld/32coDDQP6K2FFL0BJzqc
ZBLr0yFVO/hNIZlzRpZzj9E46BlQvJiufAdyY4VqYRzcr+dzSqcyppev/gm6XTqz
YgMNKFhshlotDVggEEa1M/BmIIUcJhy/C6D/vx/H4a2v3AS7ZSVVtK5Gr2AWaSUP
FfHJWHDu6gEDlrMJEbUrhp7S4WsU0axti0QW/qJWl5pG9w9Kon1tVpbcjH/D2tQu
dVwt9KBTdc+xG5tnla6vSFZ/pHdFdPVArlt7XGXVJCIHlnItxnOnCnnnx9kmpz+p
m0U3dkhxJ4m5pPi0Vwquoe/0ev4xWw8TUeJooYBJn/SRiUecUXc5o+G3UCiwE9gJ
DMz2ZVgNyz89/BKHLP02bMDCODm2l/2MjMiqePU1MtynxxmFjVfl41vTC+xD3Cp1
0icpcNjvhvAxpPY+GCmx3PnRVynhE/iWRXhi3Juhte6KzXHKRPh894zs20qvbobN
W4fMNx/++bewQv6w8d6Inb6KPr+yXZtTEpz+dp9GSHelIp2scLnl5A3YfYsYh7yq
I/djm/QHgSjVq2D3X9/pDPdk7fGGTDu6XYjgztu4LK3LqDS9w4jnwbX+zYrrsU5u
bd5HWYAZL75SWB2hM/vMPxM4lKS6eZlj9Zx0T5XHDozCrwyLlQ2w+RrDpIGx3Tfz
xr3M8KLn1j5r/V/ZWEaDaWpEc/fCWOcvz34fO4qZ2Obdf2csmY/cWWJ6Bp366DDl
DnLA3IZiOtuPee50aSI+emaIb/PK6imMY/YMKc/FdHW/D/t5Cdc0UmBqpBO2zY6I
V/KHtXIv4lTFoXdkSTYPGfVrg+boGfFxVxIxUPmfK9oXmyBbvFWlVtBeVGvgVBjZ
Wi8kNY0hBxswpSB/oAqEdDPSipMePuFOxqAOGbEedlu1K51YLjZ9pbcURC2aAYKh
xVZaaJ03YL3otEuwKR1R9XF9iU9fcPpqU2zAyOi/9egy8M+dZyNTKcYvYSTg94iZ
z58fvA06BqluqipDo3QHhePiVlf6NPLygoI31EoNnlDphjOJRCIhQ5u35VkzLoon
BHwdkj8qnF8JcZZeiQnhkMUH+iY+SlqNxOlZacTzAD31zNCDDmkYNzRbFIqawHSN
QtTr+QkAnbmvw2Bk3/oD42gd8SXMRMHoaVyN+k7GIp8cBNLXZFcrRHW4QuoS9tjA
m4albS3VLGINnMqBVe4D+x1RgCaxI7MXAsn4TUmoBv0K7zBD+wddjcJPkdov50+T
NgRoTLcM4pgRPCsTOxW+hfsTj0jz8kbi6EPD6RUOqYS5N1SYhDR+SABrAPVKGBNv
dLCUkpunzJAsBJvDNJR745RlozsjTrbb7SCS+Gw6K2BbnmKxP499s48PTMwK8pOs
rjE4yOcZB1uyrLEwuaJjrotGSGM3ERWOsHv1oxm3yyrH6Ezy3mbIAGmgqGpaS94n
bD3W3KG6Wo171m/AGeIKrxbLyJuU4QGEKxx9VU2gh154TfLOsNF1AJUuLisjsjZU
+yLrgLO3g3nfc7QE3E2POjRj509CLRIyOiL9bhh8U24NVa1NM1nt/rImbJOMz51z
m88ghu1nJuQuiWQGho29J/LTaiPLT1kIDag5k1ZYSOwvDuRjlZiG3KOHfxKJThWg
zhFbgb7cXoJIdoOrGtnQm4nbBYBB1mvwY9rMXPWCEpQvxNz+WH7YPXX6W/YlwkoD
X8FCen5Kolrm8I9fhZ64aYQEluT8XyVhxeja/S2pyNEqG3GOBk2WftsgFyrfKm7+
iUwT4ELDwO7/GruL0KeTSWhHVlxMmSgzkJiiqONwBMb0ZRxVHm53BrN4gbfGoiem
lUc30SpO0fNDRzlv3AYyrfDUWnRSV4jObxV+h9Ug7QRq0Zttr03duH+jS87p+82S
oHwp/5erbv5cX3jX2c+m+5+1aaJMAaBOEpuFhJOHRP4ZSjhHI3PlVLCMpW2HFgnY
ZX4PRpaAbGX0vH+o6rSM4B1pF+de5dLOAG86H2qncarcCylbYUXwo61NPFPtaQWU
TsdBk+OJ4X7fxieiWHJoIxk5qAB80zcH1AxDq3JA4T73BivPwcH3zBAM5LnPKiqM
4r4eiX4RSeipDz53ED0bRveicBnCIavv8ubHVuqHfC54WlNCZqImyV+7kHudOA+S
uAQBLpj5BKeOlei60nSUApujPvZNUx7Jf1d4I2QAgX9qdgU2H0f4/iAXusZL0lwY
Y8p2OzCUv92J6+l0tH81N9WxH7DofBCAzAfpENO2I10+RmuAuVolp+GrSHoajVD7
C6pMi/eg9GVvmOcQqP5EuE0y/vkmhDyoMEKroTVN3BJdig6dVzbfhMrnA/IGOMif
CMToqLP04G3SlR4Zeptu+whhL5oNa4xWRShIcDvU+y26A6tuQbOzsOJ8VEq4eAYw
CD0Z8c+Wzf45VadDy98eVdNK9wTy4AHqr+RFGccqvwXZ4BVDVQiA2i+ePhBwk6Ea
5pWH7Xd3jpRbKhGDL/2p/NT5tRZYNWNoj2+teM23Z5Z926WKilHQWTOLMVdw7Glc
n3Q6LNhE3DUNlXsjPF+Lipz0TUkSeld6p5vfftx3BfcwDjyfl2Jmi7oyVnZ/3FBh
e6BOfuN2LaeiAaEvDorBCoBCgkLgaRmpPwyFnYl6BtYMsaiLR6z15XXBSgN4M3cO
OmALQhcUq1oXk1xZOgec6HlRRXelz4sJPinHeXy89Stm4l2Z5IzOtEiMORhfiI9w
in8eYR+jdVlqwHy9K/0TEZIPVoR1nWkFCI05PdRj9DaW8J9u5XAmiLfQnHtTOdnU
pausExLJTJlXbVrwmyQHKnAu1462AYrwfx09GpHjKYhNLtVkdlerZV7it8pM07V7
EjAirJD7PMWK25VgBzp7qd4Qvd3+M69tQWIuL8iobbOIwdF5YQFNvo2+flITZZJN
XSk68BF1shy5UWf0tTS70KJuDe+dl3RogSogKaaLN1BdP5wt1uxkXh8l3eHGK6hO
UG7+oe4aq9cT8yIpK8f1PoT2RcNXZd91eTdiMmdvWd2HYyToWhFi5T1bLxjSOraQ
iH51ajyC+Vci9MskhJ6pWNxe+exPXsIuM2/f21KNou1I/Xjw0rsuGYiKFBNqMMjx
DSKpHGD2y+Jk71FtOkIe9GQxP8t4BBqHVC7GG1S47MmmTB2Y1VQii8tMx3lmewWw
kAK41AajJ1v02hq30fzxEpXJjlGDzamhI44mn+l3R0RO2EBQ82UpYqDk2U8xCtrD
7B4f9+0hxwnIC0NKPuuBymldVgmeFTZwDHa7+PnXiHfVTxkdWz6/0s9D3+NigCpY
9OxON4pUqeRrRw/JaWn4saDw2ARPtRTssNYr/JEyPkVk/fkasMsCXW+bM9pXH+CS
Ann4DQCTEN4Mb9i19SQZxEHdfvdjU5QcjdF4CQ+JVWColKU6TtK6ejMAds0Lcm6V
fcwl0IudltOoX1AVcDM8R2GrvZitmOOYQZq+0hx6hRu4vkC+sd8qP5xGYBhB1cQJ
y5RJPGRWLEq25FusdxrtNKNnR8a+l0TuQ2feYRJkQ3OEUetOs0z7x1qJqkQE1KuT
rqbYDpch6kmw/UigOCpI7EYRrEoCk8UbIMYDaFEJOxYV77egupaKEvRVb51gQUTq
tyME1ypyPFcx2gyQGd0oeaFLtgTxcbZEZk5mSsa8Jto8DZTBHzPrCfu7/WIhQWMI
80C87HSOeuk9PoUJlGJhA/gl/VX5nEB/bpYWT861qUERNwQ1BQPT+zie9E+6ARmB
l/TW9NaYuy5gX4W9rtQoes6AEG8bsOvNtfR+4B/6MkYtRvSOKeqbXAMTMBfMSqW2
4QsFA2Z9wn6r0Fzhxl0WmuTYdpuXWf5GVmtlZpjiOOD0e1zOnRJyJthGgIIdinSE
UB2GAvFLTQ5u3FVfIs+ZLyinPnoYBfOyMcQRxA/tVurRQJ1BxFGuiFju3tqZw14g
vceY4ujMXi0QRif+1asaQ1Qh4Y48mBrd/t/9PZs0KGsgw8ke2hx/ZqUiGSpPbJn0
lzla8fjVL5is7p7z2crEIUoX1evP1v+eJ9wi5oRJWRvtW291hgISQ3wFoKcOfSNZ
lohKOTAQ8qQQ9MEGU6kqoWOB1lr4hcG/M8NVx+MMCOuFEqyCimPtGKWhqNR+3gUS
YJS5ca2MQAJJv0oT8Ja48ZCTMNVGdf5NsIdGjTsGti0cLmX93xScMC1CYFM2oW40
3jOuxRzGh9d0D7jC4jDW9zp3HJBGnrrxcMEsdTRF1BPkdZtqAPUaGW/dX6qTUBXc
GTWIadw0LO12bBepuqYWUOXrB8HSPM/vVw667v3PdWya6/JBJO8q4uG17m9hnJsI
/ge+hE2m+Z0CWpASbEhe0Y/3XzvAUaLis57uoC1w78fOssIUmBzwdpSM2unJZXPf
xHrTzdR/D7Jdh/G1ZufM42I/xgUuwu5S4Yk9m5T0FpVmb/5cq8+KLRqzJ3OuLHEf
535z7ll3KK5yVRHyT6fdGj5J6pR1VdFzJJmTk17bu96rpMEyDHklxd4oVncRz39p
slrs3RqOdxI18rTrcEfiR8VD6PFNVqTMncJdHdEpgUOGXwCwLrANAeel2dzGghN/
ExFyDTIvr+9MHB9a3Vf9F8rAC+sjmxSYz0z6/JtngA5u/A9gu3EyHZcV6A+UI/x7
zWE1Z68RVPtcJTEQfh9i7eVCOGO/AcEZAaQuI3AkapanB1XtVOH9Q0iRdotldmz5
Z2edwkxxfOOa/BP5BK4tpbmHgrpdHtbQKr9Mdkq65YpGoIH3yoZwIL+Uunmv54Zd
UtMXAvc1AdfSsK7+boYn4vdBRaqkrFEXHCd23PZTdxRLIbqfhUZ4jE+57Q9LhBCV
bOxIbtC7me3vc6KTKuqOxrjbDpHEp9F/0NO0UfGYGR57IvbfuL1cmjjjb76yY7aR
yAIXU6XRErUlOB/rR4B+exvYdKKbVCzs0MjLXwREhNYMsyJbwr+70af5fjQX1rbu
ILhOVyW0pkLQgd2G+K/9xPcQSQn0JuyL0Q6gUUVuxhGRNJIYrZDtVU7e5Qx0nIQi
oz99di1yh/lh09U8XJUlSlm9HbDcdUpCzSXJrvGXggKrr2AZnNxqCxoKFrMBfZa2
zF5ybyWNdWji8OPrJ5ZSWBOvqd2G33FL5AGBLyiixRppz4UUwoKKqzjfvyhZMDqF
3nd/b+iAj5Apaa06ZdlhQvVGMb1/kedOBLi/vmSCLVBw9ICwJ95hqrDLf10PaqaL
V4cUHcI79/OYuoga8f/02ZGaVp+YXjZH6BfDeI3QuL3mS+qaYRz3rXOh5tFHsgix
Hbo9p8pvZ4RYUnuf14WUWyuV7VIeL4awPguhRVGBt1K7H5i2e7/jJC6w3EUGtplP
Q1akNDj2AdTr3Aydo0VXb3OiM/2yvsXhzwGZO3vjhf+fHsJOCWCO4s810wtYA3Eb
WVcxLY5khn2lwyK8XmJ7+2qEI/SCVJraSwdWCVsdvwlPenHLBYbHTN9sZQjzH+9D
dNhnzvpHjIITIin8ph21JipeUBWa97wLyqpCkMwDEswFoTt3xfNcyAYFPPmz4DPT
MZyvoJqiPtJMzX76Byi0Pg4ZO+fbd5cGCgeHvri6/eqbP1Zuwmfd3VQtbcCpkSqk
j8PhWa3IZtz+gPJLN6gc0fZPnt3IGZKgpt9hT9DGZpNfQPOsAp1BQpDfmdKQDrmr
rMHoUlA2zroZj5EyfTs+85TgkkaIZalSz9AmqJmQDdsViDuIst2PGrMnPfLBe4Z2
6llU9EX8r8QO/lQhluVT5S4f+jD4VaacGbWyy1a1oaD7+ovOrqScUlP4zvNVxb93
P6EQ5xURLgB7KiMjiG0b6xYvQOxjtE7jweC1iPelMBfWnmhg6TNdQXlspOrgpB92
+Lpc0d5xV/inL3NT7FazuOoNXOJEvU2zyznlUhPNT3wT7Zu3Q9e8TaVPqQhWpsMQ
A4Xa7OIbk6iOfwTPMtnv3SXKjXU67sO9zUQt6MabaQvugIZ05iiNLbvv5wilL4nA
ZGz5kVJs9YNgkXwQL11ESh3GHnlFbgpMKw00nSqjK0DqLs6N4kWuzIfC9d3DbElo
yzqSh9ABrUcgFivOv6dzAAxmXVTInXKEZV27dID8YUJHpCET9xdNGyKpB0S9qYHP
8TfJLpmi/4VkD5/pThowk9BAJzX4PezUYq8mYAQX5tgllYBqQyBYjtYPLUN5bUpa
/fao3gJSNQmnbW1p9g/zIj2OCD6xOoLSyRPmA+lwCO8Xqn2Sn7J2wkhRv9884fVn
uyhd7BpnALFIYa4VI/LITvl2ozVMs1qvzkSPkJOA1BGvwPDky+iHiJKq8hb/8rg6
g4KTAv60keb++Yf5BwLiDohUtRUvFh4lmBMKeB/ZxY2EQENLRfgJQq5MJtpka+j6
7kNRFFuNTWWa9sbP80FtL7pFRq/h3ZJENlEJFXlEDSmB2joiZsCRZgWjffjzkpaC
pIAvnpJK07/kWJ+bpwWepnJXit59FtxyXJhaJmgDKldcjUVGkIaEv4g5Z7VdundH
5dB8QQjJrilRG/isv5YMIIC+s9UvKv3tqqUG7L+uUq6oA5v2Pqq3N3BgBgHr3r/R
F2oPRhRDdPcqqCpHKyq3Xa2y2zrxJV9l55LTp9qle8/35d4uuB5QB+qbNXzTSMbI
ccktZ+tiNQB5qctux7jXrIeKIuZ0I/NwKEbbpXwIaRp9VQFAGEHyXIwV+doqYCN/
DMMkzrgEMMj2yYEnDTNp4d+zOPmKoCSX0Dh4NJXw51wLRDWXbERGxQPaY0tvHuwr
CjdFfJjitLLcauncfACugciULfhNJK55HndivmAhwszHbfIbRmGQb5ReRHxRI1zI
xcGRyHMt0Y0nwOfdoVnho1cGU6YESjv5DeeT6OJI/+ajy80+dVSGLpQnAqbLHJcZ
mNHS4DmRuw3HylEANfr9et5jumAJesgJ0Z7Rf7UU0OjbcVKM50osusqX5zdhqwWJ
2lsjAAZXu99G9sv6COzHiYHk7T0hp0LRbmqWt7ht0XgmCorZmye4dL02ovlLbep2
GY3GhqzqIhda3HEiDIWcBE0QBTOsVHNZvUOo5W9rF69snBdrPqShoR2tjaNN1bDy
Lj4L6QMJBMx8MfNkn6aq05eWxcEdmafu1uDigqDgLtj2QfHA7nyKMNiJCRFaCLVP
Sn5VxCZFmEUlPl46OfX1mSZlqh7MX66UkzOLqkZbzOi7jQGjsDjy7INksaUhDIMe
JGNpdm7vxmt5GJMbn2yDXNdTaAcOAg8GmKG/d0cYdXg3QlCSEG2weuHi4XlzwCTc
bmn3qHs1ruLWAU+BKrKvnhxv5774jsj21NGZr5mWdC4QkFdHig0D2xnQ6kXIVkxv
+Vom2FcBOH1Io8t2n3UNokr4n8WAa2dqIN2f0yNn/miOrn8gGB5QYg+q3QyVQJ+S
ebj0gLqtqnweEqCpvKFCVOIouP2VSHAvvqyBV/+DcLPShGiYz7MR5YcEhvSaCG/y
V8Q4Q6oYhuZs12UvHkCGdjqS1sqURINxagLCFR54zDpnjQHxNeKCSRcDCLcRVxIt
XnRxoPiSFD1OjZg6LN0iE9AhyCmb1zh2+xv5JSupfmN4ktzYEpZ0039Ryk1jPk1a
5kDRuGEW4TdWIwib0qYCWXoe44A9cpScX8IqN7u4pAKd2CrXOjedpzwgPDMkLT8e
GpJQK5BwreYc4nD/bZqFLtqSCuF5+Q7kAbiNpHd4gYI2tlFo2v93QNOHyGIUKuPP
xgc/IYD5GuNi00EcodAFLKAxmEOIEhy/dzybTZ/7VCDmntRq6h4QxsDmAJ+FHCnf
HUJxtU8lqbFh/A8UwB0VFwYda5oB8oE4ujzX79CXcVhNAkrzycf+v1Q78ywranNf
wRM22cSvH2M+6Lh3IGgdVSclp0XfbhyBS2G5Mmf3SlTEQHJ4lr2kCCOZ0m8cMO9c
I4WscTSsjic8LQSPX4F4wqg4297Ac1n0gAxt0UKgOaLNLu2gK/NKh+L6pXK8OOpx
0miRK13MlkYDPrFuFT+HfmuF0GGI1NVAQD5GcuFa3zJ5UhEb81CL0B0EOaxaIarP
isIYX7nOcDlKt5+7VYeocCaKFQ+EVT7gOBfzm9lmRmz5Tx5ngQ5KjQa+RPtwFTk/
MwRxWAUE06/MHGsx1/bL9XOil60UTteAXx04czUp1xFf8crpGdgYHiBl5yL341HN
xU8rgJa/D0MOZuRMX3PLTeL9fRuGPKnsBVxgx1Oz4i3vmUx53xUUrjscPCJA9wub
Wu5EO8TJKmZF9GQ/OGDsvhzRpZreRQjXeW8R84U5c+UQ0zmT65Sbc+II66rQCmlH
W3yF9WEZX10mXMMC/UhkrzXviBC9BVUHTl/w6/Rrsf26R0T5fc0Sqz/dNBpzQdoa
VrCTIP0vMgf/hGrwB5WxMFP8R0yLIBk+/qvUx4NTpTeQaP288/Dbk8vt+bdM4J3f
H5avdIKkN1AwJ+rFJ3l1QQa+ROF4nKzteu8p2orjJSAYm+Vfe7kXxWK+NrCXDzl8
2mztp1xNw38mDVAZOZz0rlS/4/LrIyJ24e3JGVEfZT4sTotaY55cOV0XyLeJG5Vg
C/5SiUn9Y+ZAgsdHEiSWnTiZUCmvIARQBDyYMU0U+LqDYOLrHFmScPOjC0W/Ff7x
Bhw5QP8LB0XVvG81z2v3BSnoeOP4X+TzUSd6uklscYr55tr2MN5bxiOXivsSwxA9
Ho6e4JvspUAJ7bEDvAdPaiNluEJCFqtDTI0qwwZcM+OPfu0fjy7Geg7IAwtC5TK8
XSpM8BzxzUxl7HLvfvrtN+Ls0uf9GFCRnFFypdmGbp8jqJKEKPThUJJQbcx1YYxq
F3tTT+lM4+MAMXUfIWI/uA3+0pUQfVYIaFBL6gpxIcb2guk73V/5nYujsRhYtc65
n+3haVxVJgsBHGLaOkc8PlPVE5vlUbCLxtAnZBEakT099/y/8WFuHi4LKydTr/KI
6VhoehoAnvoiIiDpttAeD1lV+xdfOGMBc75UCQrsAzbw0RQMczDdnz7N/2XHWMOW
spnAaakM1rhiJ5TfDcVAJ2TfM+O5eiQEQmnsKy1Xygrc+meN7KsFHO6Dmx349HgL
pisF2CLZmyn5y3azJNpBviGyn3fmN3SUFgsqhkh49Nhmwo/GVBzN8enzamO3q+g1
Tc2F7jUAJgc+P0VtyUG5fq2FjlfxcGp93FscYgvzLhkHBVhLUGa5MGEcMTVN4bzQ
sb9mYsiTuviDHPY2aliUd3e2iU5HtKOdO1JZHKWQY3ShyYwd7QTWhhxtDkqOJR6q
9B6r4/KqODLLJkZbQ3sgwCfgLfNDCs9lwmE/gbhfP6S9qKBfrhJXOOd/k4XwEfHR
me14rGxrRCjCKNiB2dS7RbOl+UCMYJ+eRVRBwa9EFQwyB/z0hoJcMwLIP/DUoLEk
U/p+ANwnd54asUbMCZLf37reG9j9ybbi0LvJPj4/+3ZarxtZ2tfHkYrX2grV62Rx
+QMjZ+HYmxrlA17ftNC1PoCRPfjwIjJWHuhLiZkum21EEoE/1R0O1yR/HoJYI3N0
9IqXkj6eX/6nBpM0xfCtDN+GAYNHcwbAsEGu7FU6LyVZpR0T8zY5iFmSsG7krxMz
0ty5wF8+KK1u8UXva6XdQ/k1hhOPoQjmHt2uauvthy3sTbroN2JeA7UdC/iyTNmM
gczKscbE26ti5Tx1rQkKUaU2GT5doSJEHlu8rz8XM6hUScdKZcqsmKBteXC+8Y4T
1Zh/kjbkrp6RA1+1QnSa3aEcYdryv6w04shC0ugGWspLK2wJN/VAwGBfHTkjdg7B
/anw3sAct7oWAJ9GsuU2doJQPQcYOihN8PHFl9Z/ESELNhJK8LyMliNwhBuMoHKf
VFpmB3GCP/n2Xpp1RR0shfDw9gNgWQYLl77i98OBMlMiNweAtQ9zIjxLv7LCgUc+
TTNG3MCC1xzhQ/ztNkf1ro//RhKxy7Uc1K8JMTlj+RPJJDBoqTmpC4uUlU9hClr0
zwYkQJur9gLR8PZuV9lfdodhrFrDoefyQtnhU+xM+AzwJB/U0QT05tlBe53UV+GX
79AVWTNh5SeMoYBU6B0qn05tTwso04wpOHX/wJbOZZn6VMxsTvC5g6pi7cl/0x0o
Ks0UOvPjqxxImIHwpNRB9PuSoGG8S6qun5Fddbd4fZpbCbnM5ZHifwR8CfkAEgxF
EFoxlX05w/JcKAnVo6m+3TV6g/ftd6L+IyCRTF56oKRl6i4q42ZlFRlmgi0HWJJ4
gqSgvsrBrAMnOozPffW6g/C9P2jkG+93agrDr1DyZZmlmp5JBRf0hRFfd4m/+Q0R
Ww5FIWgT4dzVC0MXOkcnilHcN0k7VmRE1aKjwBde3c8w8O0GiGgY5pDmuWXJjIqU
t3rsvlvtBwpVuXEUV+2hKj6j74jYJInUQfUaoSqpx44Kpz4qkZHB1cc8A7lkgTjd
eXMz48FtQ76vJ9CZXAIFuhb4ujVZKNblT+NoM4roAayhRU42yWbu6WL5CejOO6+3
ByOyYSuxs2zje9jQ0eZLV8pzQPSamBGm9GTU3TowJuOU52OxfGyi+Zd2B3ZlUWVi
7h10ZVAp6/3r6jKfzQydwtV/dzpJafeHEwLQvuaD3VuoSXCTv4TwEloqHJXpHSBm
cW9qQn24lEN5PVK8Ms1O6JWiiGNOcotdvtCTMF28BDPXImPDjL+O+pa61BybQpsI
gk49ewGF2s3Yruvk25h4MF9GOki/abpfqfJhCHYHeyqSZlPkjXjRWfQNn8lSKo2I
7U5QrjgEz9gz96EPlvxZh6PV7Owm573mceANSzpgT9AweX0iCXoizkRk/57mrJAg
29YIW9ZD4xKsRjqH/DKEr/4eLlpsiSug7rakM416599LpkcrHQx/vMt9Joj0ZMgS
KjmGr+uid++7LJBK6V6CDVs1jeNHnuWeD8w2aBbw+J04rxQF4fMl9kLvBHbtytgM
Z8XfubNkClDiyEpoHRrLVc2V2+yFmQG92BnmzoowBylrbXbJiy1c0V4AadL6i1jK
uHe2lslfSbvcAZdLC0HOF7UFEa4AKvEpOjHjkGJqXLPynNtjpEKMHWfm6skZIrpK
fn4tC2XTfwdStuuEpDD00LwkCzD98fN3M+HUiWPE/Kt6GDQUMXHkhtYzyGRFGI8o
578+4T9NlBvOVMZyedbEC3aoU6eN4LvRHVmr4My9iOaOEyGH4/+na4xFxs+mTDeC
ypu4PdYmTxoowtY/jY5l9uLrODQVbwqkAE9Xs0UkP0loom9WB4mpMIGNdKyfZ6kD
p8ivu+xj3FbP7BzQeStbgQTtaYMTlmaBy2qFNbBSj4ZRxioiELRWyUmxdzsWy3gb
668AGhGEryTZiOpcCJ9ISnsCz5FBQ+I8YUdxzWYCvLXC79JRrgSU0uDBgCnJkf+i
6Qz9OpBG86l+zNsMklvb4CFcgEkZgjr600sRyKwlhxyIrekti33L3IK0nNXRWxFh
Aa5QjmEvpYXP1pF7rqPB21XNRonkGcy4aBzSkSGAJ6qAOzBmsvVDFzSj7IP8/e5x
xXbt6qZZheM/ZAIhNk1GX1tobjbDczSRgXzExspTxWI1xHi3TNy/OTXsL9wvwFMK
XZ2TCbq7j6Uvmj+d1+PRQ/I14QrJJYQPDk92v3z3V1+L1/FZ47bAsQ2LyNa7E91e
fJJA/l/qZK0wMVs9sYGAaSSy9kdzVZOURg0OGdvAsp8TqBH4zCSEZQ0EddetSj18
M7Ud+SHnWU3e4ptA6Sqgrc2lm6k0geFWOxhYiZ8s1qSKF5Ngx9A5s0q3j/DpX/zU
gdpc/voj27QdeGrp/AOXKamC647JJ/QeZyMT5Q/QhbBurfDfQLiPPoIGI3D/qRt/
O/czbexnc+ZRtvvqYyazAOW1rZIqwNQJpnJqReBMz+OQt8yIABch9u97TDlAv/RS
/fkwy0z0OwfiegcY2BU73jJZ80s3IQvxoEAqWrN70IgESNjn5zWg72u09JdK0zfb
wyvGa37GZ9hvuL1YdNA8I9we0MIg7Gxmuwrx3reIpnRESFytTJjlQw4JyARL6HPU
OactH9VY7cKdPdvJXboxxB14LHkZr9zYddy5MQDr1bst8EyrIXV0hDv0mVQXOaC/
iTM6epqwWMwpyijCvhYx2O8mIhrBRgt5hMTbYlyhuGonpMeyur3Zm2qF/Tcm+bzW
hFQjVzGThdnRUrOu6lqy5lckIRbNE8Pd7eaz5Px3G7xvU78ceHaP8YFesi9C5oHK
wpdpAJpCGFbVpP9krZxzRHLfT/AvBjWPdz+cF5c+HJpYjyqBEz+RTT/st6TU4hFL
iMbqYlvKX7ljIkE7X1u2I2k/GayeSsUY1gRVv2jVrouqKSbtffcEU3tVk1OSJDbp
kmY9B28mM6vYPl17DnVnftlFpKCFeMHzQXRylhYGxvqAASfe7Jnz6YNYw8k8YJbD
JlxjXjltv2vYoMNeYsqwU67IEGKaVNCczd2/sAkbUn/ClGKpDHzWFpICFuGRzGU6
6DruIBZtENwW2RxiC4l2H3lLH6niFifX6BeUkO1ABVZD0TKbGIfxYfphmGpjayDW
FQcJQEHxr+S1bgrTqBnQ3kBMdtMX7kazGb65a1071wu+musPDL/ygcre2fsETa7O
/5K2kITN/yVrxx2QpcDc8oT2I4LK5g0G4gq9/bmgX1j6sLzMoYYO3za9W4x1gfsa
XyAl2SxwymO4mZqHX0x78bSEKiZzqpBTHcek8ZQoCoi4l/zatkccLsVUlALcuQjB
BG6Yiq2wkx0sGpkbQBUcfSTlOhvYIT7M5cSvhjljotjdJBKeZWjRvU+eTpr7tCWT
vh/R6A8Ty5EI8ttNo6a7ancmhwxl2IZYeNCO5qFQKbxwkTJjLBf2XhQ8UxmBMa5n
xEbfVqQOspQ9CRnEfXN3iC+ZLqj8lAFmt6LkZCg7vqjULRT9Bh4LobPE6gEmln6k
/zVPJnN+9XkFSEOGFn2zwdRruHX0VCxgkscy5V+CY02lCC5QqHn2fiSnlbJVXiLJ
3w4BWuMASaxlDmZGAZxHDTAQDTGw5QYglF5XjMUaAB2t0xDKznMFX8QCg4zON+XE
t/hWYmV4/WDGOjaFDcXoQcAT7gf56PhlNUcQK7TJL0HaDDQ0WFzWejb1j4d7vTVk
rhsBJbJJw3gUWkpzEkvM4YCADI9PRBAL3JeU/vNet3bWJO1K1FbmZSBD4j4uBSul
OHPrFqbMdNnKxOvWIT/2oUOWwn9K47dPFTQuG9WAmu/iJnpKLZ/9qZp+oXou9HO+
UjzNE4BLFGEhl8s38J+LJkVhI3Eawqc83q3vC15odI1wzLXbZg9upCmRv5NQ460n
xWaZKnl40m4HoPEzfCRVMWrVaDdVXBt8s3iMvtu0rNWL6c6rAQJdShgXiw4QMTUL
gBH3St0MQPlvQARDVNNCFSlz2Paxv0hkPsMDbsXBtLnGBLgVn5NmeBNaPHPChOSO
yaaSAgS8BoMi/wsDpiXr+Tjd7xusIcVInPfhCu1RkEQ5hx9M7c6vqL+dxqOiqTNY
ZX8CacewzABhkr4faXdu8xQpBNcUFyAEgHP42P2lOp7PgB6e63fWFScttploK44u
czBFMMXbvJZ15CtMJqjZpol+4sJjMM6O+SgvBGzUQqLt8lizxLVq/IArjUFCIYIa
IanX9RLO3DWgXWQwfKxMIakAOiSFNnGbW3deT+knYyv/00Rmwi06kuwPm/FRJXqF
6s/mEjbxlhIZ6vq0kzUIYQugrYPSOEeIH9x6SkY5QxecKdw3NQwahY8kJ3B/sie5
/pg3XvhGL7P6auSgizbLfiwoYBiTUpYKZnV9QnklGp+sd3813QEJpOzDarn+P51C
ePdcAbk0KLpEG8Z0t6E8/ClyowulaYgu9xJ5fwjJi7x27rxzgEfs/ABcjnIqI8ti
UwDDpe1YocS3eKRLThw6HaqORIST5fC2/85n2EMTPTFeBcJkcd5v6V2nnSkyAyKQ
uXG5GTy7/c5V2RGWJU1C3x+BfsdE8y7zqggRzimSOOUUsJ+YaD2OLit0wp7vCqr7
dnV1TG9EX1lEzNm2F0x0KxD5zUFyYWWLu7OaWRAV5FlKlxo74cTOU0Ps2bSU9mIS
9NUAO1Y3xWfYI3OW6JgIZ9+yaz4X4Lynogz91RvpJsTDmtz00IUg3rlP80PvKspi
7AgqLOLHafTKv6jt9QUH7VTk5AR6hubaVddNEw/y/gtdpOFd2pK9u1iV25Nrcs9d
v7+qKFEg4bfKDkftDjODSHRuZjSFARw8iUHaEvY98kCa/ASnsKEvF5gjziGGrPjH
Zbs7RfHNQSuRnCcl1BHJsEu7LGbfwGWGXxQXIztKan+Z/XCbxt1b79oF4LAOrDuy
QoDSIl7Vzw7wDnXnThiT8K1VAvJXuezAQnnPcsYRYvJeST2jiaxp8S6c3ewxnbT8
X8aTgIQa7NvDglwqcEup/RjeVRjfPgHVUxuwaL6VsF9TcFFHDzxoeU5ytOCGupkE
X/0j9XhbtvJOXzHBPU+y6xOeswXf/lsklSlPabVErMBx5GnCK5Bioh/yOmLHxVkX
uTplqWBoXsRPZJtXp5GdMIurDj9xRPhDDxxxvL4o5f2EA4CTYRpnd0sYul9xolzC
H8zOBkJ0vEQ42svBXCH4bQZ/osrSkrjM8ebLQYN+ZscOsXZOEkfUvWlI4bHi4KJL
4bneMeXnEUKJLrW1IVdQDnqzFNkTyk/NouRdI49UgCig53dA3llOs2CJ+4Mn5hDI
rJzvFh2DzITf44PzphIDEb29sCdHfNl5W7Hi+HPopZm0eobBTx9PaYfJYH9Lz7y/
9QfV3oE3TTfQJX0iDgHK/aZVJXkrlYcHsqaAAxl+P1VLUaT+I1wyJbylDPInJnCI
UOuOgMDO8jvWd9ujQc8C59qHfB8CiuyAqbHSzASQnmV/7URZj4uuCDZNHMK7XAjc
vNGlyoINqnD8aMZ+eMs7uldFvxnh1uyohv2n3ftZBKvDXaTKaFLYzuKFNTJ9CoLV
sYnQo6IhZtvtM2+lh23jzyKCxJy11EAjPUHx3/g69I7hZiR5crlCkkxXnehxi8cd
n6EW6ql2F5HT6/oNbY3104D9BnCGmruNWS3Lh18tq44kUBi014+lSRBas6fu4GyA
IkkYUEWzRkhYWCS6dQ3QVBsUB/NRiv7RqzVxnqc+ca26KdCUXmdHqmiPgJ5Ib8oX
01fmu1fKSBkogX/725zX8+QFCGrw9LCKxHV9X/K3p28ttmc3CA3zAaZ6lCw0XtmQ
nFjq+wHwtlvnz3CV8dENTqNSWIRwUyIoaCjNrM44fq9WOgDHOCBUhGUoTSGSGOdm
Tf3yBRB6YjpV50F5wVnLr6SNJOwS+VvNeJnmTGnIKgl/r5nciMZVdWejn2/SVRJV
FXB8D8XfvSuYev0P3uh0XQwfgcvzT0TRIj6oBWLx78k6pwsbE3IcbzIttVHt4OO1
8vIfbXtDrGbKnjuaGRQkVEDnqtWlvS4LZyS3LAdt4Ym7wnuDhhuSZuVH4qLAmUPU
CsPSNYn+OM1eorwGRI+8LLP5y2St5hRGmh7lwi0mjpxiQTFsGEHdMqA3AdTDQLai
BWKbm9Yt8cREFWX0Emqt7DKCAFh8mC5R4adMxCA7cga4+HSjVigZ55ksFhf6T4nT
HOMcnJJGcZJ4rMzQ9dJ4v9RcaBoWdJWlAoR+N27QvDzqYKJxv5QX3cOdGfXt9S/M
omHutf8aE+M2iduiMlK6LtXa1qKm/oyYwgNrTqfOiiMhwFOR56QpUmomo/I8FMOa
eQcjBg4REGG/pKQXxfAClKayIKLkmsjpoD0IrRhHFFi7lh+T2s12rWIrtXfyEQ6k
cAO1ao+oEe5VVmYozn3xZr7I9bPDlyhbjUkLHGqQ4W/xpYS1/XOwEFDWUAk4F83w
J03fadn6VUJokcU2uasG+YBwMAXJzsn3j+mu1jhaQ6Kad5Qu22NM4nmuti2KLNsY
iduKMtVF7T6IsJ4hYov3235/wKRV2Q9vxpDs/f9+ce6ejD5Gw0+RSExsIXogzs50
pvR0PywQsM1jtnwsPgEi2D9+EWZxfhx2aXU7+JrZawc4jOOYWcq/fw4zQoiOBWs3
lHmwip0/tLV/oyPOvqaj02y2o1uHzgLrlH6ffRsVchRGhAdfViIkRpSg61BYzB/t
IPCiWEmQprYc/FLMllWg9SyxL2CNRYAColNLXZr0wrPGR74BoXg/O9ctDhlX/wlV
TZzH6rbKJOOfNSaD1ntvvJqUD2tRLJVkLVWdrciTYCztlUdGpLEcfz47Zjy+0bWE
gs7tgw3l8nFV679qVLwNVb1GHDwK/0Z0qh3RJzOYAHLTLeEiaPqXkJrX93O2HdkV
BApEbgUUJ0EpFMluKb0HLsd1zOQGnKEfu+JemjA4muYg+C6h+7U/dZFjwEEfSRp/
AspgXxUkyiqZ7zYvlytZRO6h/4w6YSTphbQgmNDE3m5orzXA1R2ikJ2Lkjyn5iFx
HsZKWGQRP/eZgAKjcbud+UXxXSxaT/JK/0OxhjSNI1kEi2AUwFztuocc+RC1H7mR
SQPskaRgwCLOOFxUVbKWB9v4ovc5HTA/KQdHcjjwdBIbGOqfk2CeWAtEyDd5fbmB
BnhuKud1odRKX0aSTRiYoVVlFn+wyRPwpvTCL6mkFf9nXR2B5gu7WFd3yg78IThD
bzuDV//s+OuL743kELP0WAMh3bXRzUU4wl90jGf02d6I/4aEiCBRFfZEjhdfzqg6
LBpKhpjJHjajw/CnqHIHHJDVvYdZoaNDE1q/7iMH3Tik/IWmc7RoDwn0kFSl9vTE
QJOuKvFBIriUyn+fktvcuL6Br8XKjMhUmNk1FQ8CO9HoMW0XFr+tBES8PrUjEebd
uIF5M9Fsncak8zkatGeftnYoXl8dIyAljFs2f8sSKv5WqDA6QAz/k1hML2ObmXtt
LeIbzp1iX3/tqf39tJSoraaMINAhIP+lA4o2FtKZhbAM1ifPuw5ZCRyAQQ5Uxq3t
PoYvMSoYXBn4NIA5Ir5S8KPBPRDyJiCCwYeYgLGV4RBEUq3xETtAjYzIjrMrXcXU
1mkBNtWaO299CYVF5TKt3hLEAyBaIynbcTICskB3sbIj3t6+cQD+RwxFrTZnyWnx
MIUtO2/alPAqMQenpBZLq6Njqrlr4PMSWMmbBeAteHTg4npm2wccSUsMPSdO571+
my3h+JxVnkCU5WAj1tDfB1d7UVhdTOavUaLafZyG33z1DQquy/o2dKgTM+K70aQs
sSLP3Sl1itsW7MtnfmO1fiE/2RTYZJae/p8mM8J+aHDL2lXIdyFvsSIRw7AtPsrK
7OfmKVEyxKo34x3sUbSpebFdTDqcbSvgvGiuISkFvxNlMiBzeWwmAzTWosaqU5mE
20MvRFhKZsBljQorA3M6VzwVVYklTPWJVjJFX8bG5JHAvxb3nCiPizRl9nLxn8Cv
LvrjBVpo+17y3UGNIgD3DuGzQJdOvk/n5/bkwOT4Wkc11J83Xo3IypOuKDupWuwm
DdeljFlp3DTcIjrc5EF+amjt7m5RofZKNZ3AMPA0T+g9cVLJxXPONpf4aPsWbNz8
aXOsuc1co0rTcqOljRfuMFTwkKnTBFMzp+PuIGnLT5JpyZgnT82Vqu4Iz2sU1i2u
F7vaatvVwnPREE0u4vFT0sMoapOY3RKJQh6ZvB8ey6GdXKiQxbfbmpTBl3qVFPi1
o9vZ2K66Bokz9NgIuOu4VdvyBxIclzuDmF1JnAL2F0AujUCJc5S6RHBwgEQBtXrI
nBvv+lNOIrWTuze2Mt2JUsYTNPTs2aurGTY/bPlocD62e21FD2Q2zM+Aei5Gobvk
5g7ApunipWwrYHBZUpji2sLvEy7Vz2PtXsLmDsXIaq1lexJVh9CKcNYud1ptEZk7
NhfNL3DpYHyiKAfAnJlQE06iPA4Y0iXwAUJL869gCw9EfvBcKLyvxkvR3eZ9f1ch
UkW2eFR2EuEQWEmkypNWcTF0cHKkCBGEfjaEnfxfF3wN61l/ZJ3L9kVRne5v10Jv
HHOZNdcKFAvB/0HY0yvLFCZhcc2nY7VySOTaCdgOnekmLoGYPzsR+XpOSHIoIROF
iXnFStoa3b2EoAamdXCGqPMpnk2jYg0Nps8rNZUyoDkfAGau0ifzm0AY+4UoJyAq
Y6UBGGcRwgaB/YwpTAttfv1apMxrBj926qYYFPN12aJeZ5Q4lVD68GBcfsl6Lqom
p7qxJdDwD9HobQP3iSdjqj2E7elKeq1mOjTRsrYkzggHK6s+UlT3aZ6e9HZuNSCP
hYUUJxSvTRw8RMgdXVdD1GR8n97RIQC3d7b8A59aSd5pEubJOT31sch6Z/iEsfnt
Kg8iK22ttlmd2L0mfENrOotbPm29n3gIG87PMH5XcwRGdQiZsETinSL3PiYdHgbD
RhD5wlfrKjf9ea0KIAHRtuDJIn+6rjkNrjQNdG5kalspJmyI/1hzzwJeX7LzGoNM
VbFzAuTsJVYYZUPfrCm+LHSv1QeakkKLl9AbtUCEezb4EEZN1J4bfCnL3lSia+dL
IWgmOfc5vv7q0+nTv9lpndSkjz6+KckGtYkqrxBaxo3O+/j+lSr+/5tWvi0YDsR/
F52vByRPz+llnaEzthA5oihTnxBffkIYu5pzLtu1izbb3Yu51rzEA0B0Iix5+P0w
RwBYE+U91cK9eRFXst8bzv1cizA4SaxgyPZqjPgsnVs0biemEvYxbRO3oVae/aNF
NPixPgbVl8P341giU7OTVAsYMuzaqipIR9MPoRd7t49Vgwok69r3BG48yIjSVf/z
aD9lgWUuIB3fYfh3EMhaO6jkUgkG423r4iNDmYrBj4dD8i6U8Ki4qv8TX/zZ2lx8
Qo+zudts31/DhE85If5oH220J/gg3MFUcKJW+Z4mQDb6kAu4j+qg0UphMnoyJ2hc
shfkcVeqAE11Hyh3hzewM9jdQXKG+xPYQLSVECu81gGGW8yp5WldKCkHHVfyQ/MN
bVZXCFOBNyIy572QmKN8yrJXMVKXxjauHwQKazZ0B6xsq41atdNIV//K6UYz1HXr
BZHsfdjcF8ifpWru1M45tdBceEHQWHiKXLbDrFpcmI6GPJ10IdHPhlodJ8hvXF2r
ITJ0niEgxiyyHoBRa3vDv0KWWhpplsV15nP3++w/Huvfz8sGg+xjdjOc2U0shsaQ
7PcCAb1ltRJTIrLKQy7/hyNmsP+Girft5WNwkquaXbTo3Wl8jxs9CLoEB973qUOi
lYCNQ89QA23rGzIPDosUhnC05YgcnY89I2boYcQr8RnAo/m760G1iyY3WlZKhES3
iAWaVyC8k2ELSB58dUDeomtV774kog8FbuGIAFLy1Dn/W9dyacQ2KlNhEYKdspCk
X+jHFe9H6MHnXKbBAFWBsej1vxMRbuo24NltGPamROv83LF0/MrW+8i5m+pMmPPK
wlREvUadgtzUkzHX/0xe54kI38H0/34mN3vTx5HuQsBv6rRobBXhURvXPCsvaT1a
fJ6vIy/q2JSwQlwP5vMZo4wBD464dEyJ8BmYvh5nVc4VGSkMvk8m5rpQKunkoGoM
S+SrEfIsEf97+prCIVo3Pn36r86JpmNsCltvQs953fwiz/5HWMYZs4wtneWJkMSa
JtAxyX+8640Pk1xpelwGHixiupRZfObxqv00+g4JBxvMxgolm+Jp3k4m6WHrNEXt
+6lOLNzH+HJLfGqPM8/CxLNfTZr8MKSeOgoZSwKv7SToXFvvZ/Fh3d90cOYrnUwS
S3i/YLPHHNPrf3myW8ZFCHhIpoZhH2hQC8mzBtTUjoSdS5EcaHXJLkhBKKGHlJn1
2+F2uBAytSmUOdbgxhDPJ3tegcWSTTHGV+RHAz1eRpN+VNRtxhSF9SgLfZPosa9m
T1QSpebZaLElZx4XWTdcOWUBloGzHet4jYOlYuth65vq/vGxS2fWQCmJWhvWwmVs
yuTOyGdAOn1mYVJoLOLgsXttqh6N2fgtKezQ88tS0zUfeb0l2T1dBLdlntdIRvx6
tbgaVdLf+c7ZBvoG0bN4pzcmsn+1VMD+gb6/om0lnFVbwYgZwvao5gpDJdFoms/3
eKcduykLyE3jCrnBFHR7bK1y4lho26nl6VDYIYVuXC/5+J1RZOtjHAv6SAE/zX4K
hZZh7fg+EBwhkhN26QHlacOw+k0qJV+s4LbYMvgaT6iUGbCDLO/eD+ifAW6Vof07
B5PtZ7398O+aCnFt4kMJZxQcK4truKNOquHrWSUj0VHzTZhZV44KRuZyNjTtY+eN
evne2k0iW4iv15mtaTI0mgYJqZvoPe8k68wn7RWHxFPj5YpUim+vMCV5udT19d3J
OmCH8T4n1gjaoOx5jYQWuGk3a8GXn4R4uN1TRauw+QJS6ONVNN+9Q2ALyCg8nrb0
96iBzEt2Oyn5SwPmp4xCoWNj6dDEea9pX7NX1kOW1EL+ShcXrWeTjGjtrhkxcB7E
1UmWvFsKAxgz1Y2sYi4v2G2AzmMkYyl6ictAQJF8wPV96BhfmGd6RtbVJskbAZOb
IdjCEn1pOwvJhaQ8zLCtdTA5h8blHyRxbFuBpHq2CNbc3EAhWeWI6KDUBxXvUUcX
og1DESvrjrpN7OTTeMJOArAU6GC3TJWxuoYM8xv2AH/ndul0yNYzdYDdWihiUPu2
LCErakhZsmUfhi/WQjNb2oFuKc+L8kjAFM78wqmBawS5VT/8fX3dO3G/VzS+zXEc
5bqgFmW2kO4H8u2b132pd7f037CSGvVieSsXp/5jy+xWNy8l+SKnq6WKQCfIUwuV
lTaAebUxqKIPtLUmhQheRtnfjibN+Ok62bBX0x8W0hjTPrrRoVowrQmCQuBcMRPE
nhHsP23oyYG1PTEgu1ngZ3/FI/GCCgDNDyrS50P4oPCPO6jmyq4ol6MBRMRkndGb
B3tODbvTYt6kqwhxB+Q7DdyaRPIKhb0hxAd46HiBkboxH1fhBRufUsrMzZniqroF
dv24RdLLOxD6Y80JcjAEY2ZkQwopEfUULFLtpQN5uUTK3uxiO5g6Q/ZDbOaT6U2X
UM+upEGb66tC4PTr8zT6VyTMsuFj9ak/Tz7eCnDiOCVDjY5scuB9R+00x0iT9JEi
bHA71RKhdnekh5rDhD95IKLJyDpmZWCtDFSpy7XxttLa9LorCHNymg6hkh0VbbsF
Lfx7x1mBorV4y8K+5vSDB1VQYXg7dSn19QTWpHIfJPPZTxHkGdeBUHfQOFpFUXwZ
Yo7qvvKC1fF3/zukRu4u0U0RJ6szGzF736s7jM5aIpgGtY5HgqLY7N16xg+C70vn
LWqdSNAqugZfSp8QM7zIXSN4v/otSKDQaMTRos1WoXC+CT1hCuXT3kEBlTAX2rrt
s2jNxPIBr56aSRkvrXp/pr4kcDEOMvh3Y86FHpDtpcqtpO/2ih4d0KTx2dkel+Ig
fEOwgMhBK3AH+mjQdYWKChcXoebRbdrChulJ7JTVIZhwCIF+sCMYqvt0bV4ZqC27
yTmDDo0TzW24wknOrS0u3ZLSIXbXW/XSeKd7hj2NulocbBRrIXM2Q/3Fnw4VKPZE
k/L8+yrkOxg6WnEk6xbhk7UdbQ9QRHV6hfEcv7pB//h8IFFgZyRwO1PqN3OvtE5X
PT8YYhaRItEcZME5WkEFbaS2kzHQr26HS86nx3sRsURNHVzw6QNIE9HAXeeUyypF
1ZMtaSnH5LDdagICbK8pRnwBQaflW1QyDgvxkRDv5FuOWrSRySwh7DMzSwUkZ0zz
zdlpEcv7JlFuOETYWOwu5YW0DeNnBmTgjLKrNdW48POCnGLCK/VsowkFs9OtLGqi
I0muy3kv8QhMzi92z1St7Aijpcdw9ui319cQehvrQGbzxnLPqqqxtQjhfZ9IyRAT
226H9r/bUK/CvdB+w9AVk2C7GFBEO2LWy1enzdy37PxbLZ4Wc1+dqIWkpi10FnH6
ZMxwKYasywcj2qr9dIWgu3HAcvqRTqpbuU2wfse45fxOQtXNXScTV6W6mnAlWZS6
Jk2TgjlIz6vz00QuiQsYs3QzWHBcGMzYS8O7yhDGBRdKkFFTn0yIsst7fq3o3ufO
r6+vrrDCcZDumB1FIlap0RLw13l2IWYwmUbF5uL9H7wVfKTrJAakZxBudoNmGMCe
KUHSGb88+Zxvqxfo+scC1EFtpiRr9cB++Rm1fuTzELagxngTdK72fkLRD5ccnJya
L7Qjk7vJDyz1/FK2zKXSdJP7R390GIy7sNPBXvrU2jXyPJAIPKdo5nNSVhaOatVV
ZM/jhhnFByf0TPciIYTMQlFuD0pEfFtZlWQlnkfjjp6AUHS58Bg2I9oqp0BjjMGK
/q6Wwr1AK0THWkulh4KqIMnTGmlbVGbcpFS2lRTyrToEKIOVhii5FQv8KwJ9AwC4
gPG26inxAD013CIQdZSD/K0tVYyeZD0W/2IvjAqhpykVpyJdNrVpnJdfi/6UzM3V
LgEmDJoi18nrxWkAG77mF1GueZTj8+WwIEw7gy+GkNfcHFVrr2WKZayQ1EEgYjz5
e6unvhJ+sXPysGfPcnj0jVhdtQBvJKjPckCBw4tpVp7+z5F4qBOOkw4nC0fHEzlh
zaRM6CS/rqfx1fC9QIoZQeFNpV+SZZhBKI68Z+5cYHl/CLSc/ZBNp+bb5OWxzX8v
rsliNhJ1Kqt57E0TbU7xLNpxb5gFaAoInauaa/EARzbUZtM0MBtZDfrCLkWpH4Cj
h8cptTOYawOzVK5Gncq2SbCUw4GRtDTbLw7J07DThsUJJpaDqJ8iXlyu/k4ghgUz
KCetrdCJSlKsVAl3JnaddkKmmVsJieGIWbIjnKrWG7DlTsCxkPL+W5Gqb2X5wsZy
q1bpxbiqhyq7yJnrlDn4N7fLh7dm430naNq2PjKqxsjXinNYUQg179nrSOmUYSgB
wn7EQ9y+ianHkyX2zGc+WpQo6wAbMdXp8BAkwtenwRhP7XES/mUmPjBU2K2D7EOM
DSVmTi3ci6H/SBhunCBcHEnSqWyZEEWoZTGQnkf3X2L8FuAyPpEMWJHQ/BIG1Cz0
yD4cAKm115mUMQb3DaiOSK2U5z28ncdz6ZqL4yQiI+HgILIWVZjuZ8PYiTaOS43k
PuY6Cgl2uyYvv1akIUSUpTJ2dkksSk5ws8hfyXsDNWZNZd13JlH+4qvrA6RXohxp
7DUABwUeB/xDliT75oRMlZwfCNHXGWDSWJGZSnu03usvsMHoL0e64b/A9biYIcWU
fgS2DOBZPHbUyIOLTVkMW62RM8wh57EkNLFABNJDOIMdMef6fCXjNUr0laucWBl1
AxbwM1I1M39LetDpXxiXm+3aVuh7YgYW2NN6fV0jC2Cdg7iGBPnlopvmsLKnriZv
jIMl+vUpTSOtCc33FO8qNnk5YJFwH7QTaIQvr1w3IQxT3oE3MCVLXkvTJUTfIYkj
MGQ1r++PaRpKqOydsoUd9KKx38qaRwRn7ok152WVIq/uLJvCYXBJFp43ErP0nxzi
CDvSDjSdSiko60KlOA3aLnJp2iErdH9lrVXlG4hTjb16Yf32oXPgVrwpGQwS2mjT
dhMcxjMa5n9RPVsb3RTHvfUYV9LlTClHntP9pqVNLm8rKCmdPC/5iK+uA2B2+0ON
dRaZ4RrRza8R7oHmUPMPJ58HfAYjTth3ZgApD8AoPct0ak5PN7pX7MFTTeIYucNw
7v4v7e4PZSNLGS7Bx4ua/XcgWsMseMjuqyD/lxpN07m9uZyONmN/RvOMe6+DazKd
Pwdv6lsnZO5cYxmRYdcZTmOyHdx28j2U/N3YEiZlFNjHNPnIzlo+j2ms6ExDn8Ah
uaG38U0G6zsGUQNiuEBGU7b0PHU4rpvSRJgLWeJ9Ir3Bo8STs731F9DWqbTj3INW
mvOIlVJOwoNCQbYkHwT/dlcDpMJ17KxTMXR1zNTgweEdH0pFgGyLKY34oPvD5io7
WyDfXWwCdfwPMxDwi4pB7RE2eT7MXzl7FjK/x+vCUUj3/z6Y+wPZRHrCgsPhuAor
XDNwVW4AeI9I31yr/3Z5I1X6J43+DRrprSaidpWZNcptJCtI26uMhpXpsDhxjXsE
EAWdHTCjEWD1/5HMFlDhofMvKHBzAAs8r1AANbbSwvyb8vQyfrRXNXnn3FQx+EcC
tPrWnrbAizFHiuKTaA9tCOkBFD/pE8OAS4ZIYTjrSIgWKXqCbOaXgZ8sZijMw3a9
9lXm9gIw1e30Mas8fBz6vG9XSJ70rpQc9fmGN9IUFGIdgbj7hwxampKjOYxQ8XjY
wwwLzHJTjel4PXXy5+e5UeQhpb6w5uBbUpGboa+nVB5BRJfm/dt5HjIlRj5uKd1u
f+5cFjlpL1bgNzJ9mHcHwEUutUn1nO5IoMyx8jsw+Obu58lvwsBc6nyKKNQiM4BJ
Gv9MB81DdNTzOOotkjFHkiQVEVphfu6+512KSeZ7/80zhx1TAf6mUkew7wmXcLV8
Y/e1LWs/4zngV8q8koUv4qEXl5LbS33vrmKE1KMAOqNiVF93mJqQQxqvc6PuDftK
p7rTmWDcOUlYcDOWHzP758kU6chjisgj9qOrZfnYqNHDS7/YzbZ8rnumien9KNv9
itdj8e6VD4oVhmQuuRtR4rWltIPiXi1zMftIux58+01i8kWy5XDAZzXQj5DrphEr
1KoT8Lvq8To5Njnzya+Yhig+dN9VomATpGeIu1G7liC/0HxX410jj5fODZCglXON
w13L4k60yDlq70k06y/F3qjv2S3g7MFAe2VUUVS9LMaEZ54GYbSnzPsCEeGOo+iD
1sI91T4RY1NurUwrRt4gx/DxjKrSVfm+Lvy+NPR0rZD5zUvkw7xmetyV5EpEAtSn
krZWll3squ4lbZ+vYRgZBGmrWEWgGaqy8R/0+NlJe/R5Y5BcvZgzorOmyoW660h9
KlR9rVNUjElDIT5daZnjPTtWl36YPPg6zAfh8gxZ7WLuYzG1DFmo0sJrjrn7xcr6
KD6w51aMyZ0S0oa8lchTjzeEG05H8QoMzFnbXA7qSNUEkERyDAI8VgPBnzBqIEB0
/0NYw7f6FXYGQA9p8dSuU5BjTFfVJyo01QB+gsANEuZiHGAJpjAx8Tp6Mf1mvWVk
Cd6a3Byfl+IY+ybePT5CSGAS6IFeP5ciD2Nm+XIbTucb6crBIG365vmZ8jDlhQWg
FH7nQa2pUNhBKz02ygQwcUsRnOWvmXxRh/puD+enRJRnmxLh5mYG4d1xYp41+BKO
VQDhgpJI3QKsB/YTJczJBegP+lcm1KfnNLnudSZHazdJPzKS1ssCD5lOn0FJpKro
6Jm7EGGYmomHjPOiJySWbw8u2KmTEjEeTklzd36RfvjZZMiGhOQfOVUeKKkZzt7A
Staet7ZIonSR4Qkb9xqq8ej3b8diA4V/MxiX3MTg2qk63XfATiFt2HOS9ig0qkKz
I+eH7iKSzpvpPYBoRrTwXViJgIBpF3Tvwh6KgxcisEBFgrYqfNRVHRDa0Q4kwQiB
GbPfCMihLlDrGULJkRKaDga9tSeCEve4dYp52u76IBZe7wjjMG+WIGjpYD7UWxms
RKUI2AneBlfJa+1Mhn3EzdutxD+QzqT34kXF8XSl5qeV5OiiFrkzVC34eFq4yM7T
lkmOZja6mz+Jw7Hfd2u6+Ejv1Dc8z6T5mV0ori0LYq1h8OouPX23L1FiK0ZSLP6O
DuEQnsGENrJMfhWBu9f/rVrTwBMoQ2utIOnXanLW2pnhLGp4QhAAarcInnKpDb8Z
rArFUOHvvj6a3QyNjlIie9nANPzUUoTFxEH1mYMbLePcuzxColnIXiNr7o5cksq0
TJ2Ae4iVrH7AnEQAf2q4KFD4134Z3OgHNY+58NGg6djf5pZvkPmtlBVTzwQvDqOw
lLAaON8kPSNsq9d5YAFz+OP4XWgSaP39fCFa9TMeV8g6HkgU8JfL6nekJ4ugG+//
l4vAzeoRqE3IJg1oKLp5SqWsbf0sg6BKBnRfKWAfoJo+hbTagJWA5l9rZoC91NR5
Bi0WCGIuXuOYPx94tyj8zd7zheWC3gwMWma83GTG0Q5aojNgvJioV1LQdg58A5Af
ozZgJ1NZDkiSF69oRW5L903XqI1aaunR89BhKf14Z1Ux3cuHDEkkr07Z/Q5kuaVh
i6JUbcDm5Wx2dbRnFTQY0gYZPuWrrCp5pz2QsVLi0IijNRPNOwV+hDb1i9ibhDEu
Y24Xsc1YmymNZexWBboKdXE7u1e2GRPm1rRCtgidjAxvdU9bv2Y5ymdIf8edZ1nl
UB5JtSiBTppc1ftvBWmQK+H35k2q9Qi1hTM44feV6se1R1zqHrEgnPIVsWw+0L/+
KZqzKYQyqhmUEa3aUh732oU1zqmjPZoZf2J/A4p9RsYTDZpzO2emcPdaak0C5+Ry
+hBxT6be+U3meRdE5tfQRlkywsKP3p7XCZupb6ifCrA7KKV3HtbkZKLk5PveSXLH
DG1fePa8gLftlXGjcn9gghZ+Q2MzLQN3nA6i7uTj0y0UO0axqH1RdeeyUEhe5zr2
Sf+9TW0t5Thyw7sbkbs8cQWOknrp4D18PN2Iemmd4bhmKPPPzUJE79CAdoWDjEE5
/YOdZp72DZsJ48RecHuiMiVBRs7/GfGSPN6//HjBDAfBMzX1iOVFLhmvZgQNKo/E
ELmY1S/aZnxyrshtTjh6cZxmLmjsWDOpcnpFpLvvfYMnrgpomnSFzTYmK7eATWNe
I0pSxaJobxDfbJeMikVVCAXiKlprfXgR2feSRwRwmwErrVy6L+LlZi8InxeMZ0rI
sqkU/cP26DwqLr8vj3TyYJFI2uM498ie/W7TuVRvRMXa+NFx6eA1XQ0N7o2S6Gkp
IQaOHtE8B4aluKfWilorSIMz2SVgEvjTaSdWnajcqOKbNB7J3jY5Nztxfh9Kq8P+
TBmRiuUHLqDMXnhyIqcL/v6xX1J2BnClo82T5+k1uiv20Nv3J0NRd7jTsu7HKuk5
dwOWdH+dKU2C/SozaSoVTm4wgBaJda3/qoO4y3m/3xthDYk0qKddZNoG1KLLOuF6
+deE3GRH+uJlh0wbRPgZq9sZku8MMpiZQIT9PpwuunfMmifbCheyy+/1RWiNW3eN
UQ+NdJvAHR3CkD/sqhlnSisfK5kWcCvjFwM1v0kz+7q9jHKz6CD9cUcY3oxDUkRZ
Q5JO+aR50JIvp3/8XXqMq7b+U2lVpnh5xGhC+Lo+xCJypASj3QuFbshlyD1HIKoj
hPRDE65aFDuMeykWxw/zTM3vTjCX6uQKLBektu9896ZMZkIF3Vr4ypazDwOy3BA7
Zp/HZ2Yltbj0+xY3/mU9NtSuyEgP3JzXoMX6LltehzuEB1cTYSrvMTKXFTNNoLoF
29VkjFol8ct4Z2OfzQTrhZ9T/IJVinC8LFerkuSaQA2iBv/GNMMuM8jAIMimVplm
YeFXSV5pH1GmAvkATB+JRVQ1Qspfxs54kT0VewB+eTQEeENyAWbGusstzx884vax
IPynX6Vnk29bQ9dVMASqF5UYxZlXcOqduGnT2s/BUGfuYysjfy6PixzHnxMDCgaE
05alhfcqJh3YLz+jZd+aZYRxYt0Cb30R7Sw0vcYotfmyrhmqK8HDh+TF13UdmxU8
UmTzle/XoPVa2qTm4amXd0j2RZv/iltvW8nNt+W3HFxzVouPkIRKAgUcZOkAX8dU
+jwyUfa3XUYZzplANEe2rsr6Qu9Rtbg6q0kd3gxnYFNL10a+KbGsrrGGHwFxmvge
RovglUUqHnMD1qyHZ01BCWUcYbMDg/aFExekMJ+e6/yMl8moU8lQUl3MzwoCRThz
P6qc0/dpS+4HHD9WSsWp6u+wIOVexYaJMJDqSPkTo/dbiWhTH1eukTM0i0ANjPHx
Nl11h4dvKerqNvqMmI2FoAOlJyx6vYHfRhiNo/4sxKC3UtYvUwC+3SgkhHJ5fxLI
PK60qNcydLtyzawjKim9NKVsKJpr4jBPxZ01uBMvcDTeTAPyVsrCGoMKH+ocyurL
Suk4imF7Z1EDTs4WqPZOFoBnDltGZAdjW21YZiB7j3PQpDmgaL7L7Ar6J3QWvCJT
EO8+vDwMpCXq5jjdmEqHncq3zneU/98zf+7aZP70sk+q1osleLJebHgNXR2oiz8Z
MgZINJFuq/kDqF+e5inlixD9Y1GISIGwx7Rtm5tqkwxLtXV3EUh+Zaab3lTWiSNq
cawgCSpM0BtpEEnWF12Go7DLWlyriVVmfjvDVwH726I6lrDlMKneFr4HIU6DUc6c
UF5RzPcXH747+Pk/PHEQJEf1m5SW9uulM5y8u7F0cJeBCngKdZsCRZVSHq7/fSHw
3wFXkG7aNVHBto2/aABBUFYwRVHK2eEmglL91K8v+51MLj//HNxF5HcIQncHtZje
6LgJoxZuLO2rs7d4wY+l8IPk/1bBbqkwSyfDuHaCNAEMHBUiHxHWNyjZhdKPLvNA
s+wO1cGPbgjPmzWgC1fbUnkqChfyIElP+H/5YtcLoM0Wq2pzguXnXOPe+P1U8fXk
LBw85suM///+npG2bJkjR46YYqZ3XC700sJ2Qo+4kOyjcgwaooB7xL4NWECYXboQ
yFrZEU30/tElnadsxR2nTXi0UhTKc8m9bxOS7ygEVduYEDLX2qmJZTeE/X4R35Gr
lxaAC6Lo99L6h1TzQaviQV5XgL/e1j/npY+Gx5nUItdSBc/UNyZm4PTJp5eDSHB3
DcDMRAUGUpOToKcJa137/RzVK5vgo+v3CFK6npwbtfPFhUe6jzThvFaryPq/ysx/
XtFypAjeFxS+SCcHXQi/281H/ndHWwVJbRTIgV9jpA7At+MTsRhvQPAK71XBnDQZ
I7Mt6qzM8IwGuSNSii17vN7vhqKMsmPBMGukCtAJl+ZiA7aUsTsu1gugJRmJrM0L
xT+BVuIgDez9CMH3L9/Wm8DubLfWv9/toQ/GRZS3YBbZFiSbjxGNRzmZxtyZaIdk
rsRRC3hB7O8LhLPxhoWLSthEszmNBweMt0iARDJbzFPA5/GrXh89mSWmPSdH+17+
BNdhLIRRH5uupuW+5r4SY/dMPgFxaA8CfcLcn4WOkOuTY5nHQquD9b3Wzw/50dPv
pjPCN1C3KTpa9PgrILGiqUuyoSOob9PRP4u2rvkwJFeMKmbaJJuu/kIo7g060G7w
6B8rIgelRq/nzZwwQ/g+qz2C3oOD3pnxcmYRabdNI4J3jReYRKahpEkPvyOIdYqK
t5Z4WM0ZxQ3Cb9jjZ34eJhubJIzLYMs7m0sp6LNHMg2MIWvPk1BlRafRbv5iayRR
IfFZ7tsSDcY/trbnPHG+ju2HE5RVB/lAZcyZnDdYyiFC8exvkBGTYGlE6qJuHbGZ
zm+LPba6bjfDGlQqoh3IPyw6VgZuiT0GHIhRB3ZZH06mHq3Qd0eMcGvmiCi7TmWq
KesckNfOGgOFWral3Q9wMUhQ1AYe3KyewxvOlroAiIbj5u0J7sB0X3tTxncQiFN+
gS1LioRjIvJfFi+ZUKUSAySgXckBl73FDC5Cxnlu67dq5xF1D5efub5EiZaJ61wE
gv5FjSrrQYu8ch41h2rUzehmCgdijk8qrtiOD0a+wuFuz2qcc35Fcj2WjopqsIPO
LCyjQQUWtn+0pSxgfOgGOzKCKUEMsETTbtK1mXDQs6CoCAKTt+lZ8UCvjaCncOXk
B8cUH7XcVWJ0tHhbOMRq0GqXD7C7Cs+9H4Htr3KoY2/HvBwFVQkry52ncmh0jxFk
Br7Ddu3qs/LkILhc/cEjgVY7+SRzu6jBUvSTX6P4I60YOZJjmA1hse+cwekaMTUV
Z6DnOH1AilwA+3SCB/0HdlYgUIP3eUMZAAlbZpjwlD/ab+pqN1fzndJ0l+aHD2bE
rZpe31+HB0IoBWuyjnN15nM21J8e4+4zWTAjFJtC2Yt1/FXFQnCIlSyxW9tkW4az
sMLgk6XF1iT6UY1krN4uRCA0XAUmiSHrzUMh/+r7zCMHeeLFdbRAQUWwTtYne0Jj
NeJwGQOBDpbK9C3cAhLiY/Qj81D3Fbc4w8XgTvyTbrSZyF0zZ1I1drNob2rPlBH2
xFpchlAkXtuE/nAuuHnH5SdPA4Hkfcbd2z8gFK8uFhnJij+YBdLKTCo/p7QOZlB3
g//MCfLEMQdHNmPj9pwu362OkCyRwseO4LSIi1mysAK5rr2yvC2JiIW6j7Gh+3oP
Vca1pASGS9sM/BqHkZUyxbl0Tk/aebjG49NssE5sStY3i3WhaUtwxpV9dhg5husA
EbeWZEZw5hBwfkH4NWO4YtqRz7J8clrSiPtbo+0G3O79H05lH0AajZlLo88r92Za
sTTYttwZydOLCl8ESjh+ln9OGc874xYCuWTHhx9B5Y7efB3C8JQu2qMucXg6W0Jf
iUumsFfXAI1lOs7nABpkBxovjhAN/SPKQu3ff6uOD9qx420bcWje0boL9yfGyliC
054FsyDyo+fCl2f5Nu/JGqtk6q40QIxpnVKm3oLr2/Lw+IREajMMs4cg9QJlvkd9
9rugjQBdMjl5lL74AFapyZNhcc/qvI5nxRVpOchuTJNA0n59tvG8YIeDnr+rbg/Y
XEotqM8RvJ/R/e4Cql8XkHlifZ0vnmXoy+j7On0O2IXHnNkGQsv9rb9DWkXsLTvv
fc3O7qlo2UUgzhocZDZiVAEcj9CpmL4aER4t3nQyT488tkD5pwS5hH+dfWZqAbCV
GMrokV6q5iSTTblY4nBID5FwXBvYhvBRHeZ8C0jTSGx96roK2COWohuuv1PhZn8Q
nrG0Bu/Mxh/4UAK8xl0dVuXf67pjvz+LhCsooLBlaCKqk3tdP/XjirOtJcDrO6WK
FH86TJwzKQAbdMd6llhUakqiry+bsslQYLIzPpyzyrohwWCMIBlxS7Z3gxMVAawA
6LFb1f5EryVOZOH4DYrG6Ug/XBL4pAnB062xlJVeuzmhYJyc3jv5RTWAxGQFSvvY
r7pFgVC9NFW/WrHRy6vd5uMlgEQovSQBfpYBnNcqPazgU673Mu/EmK6wPPjJwJ8Z
qiwj8HYsEYmPH35zOAsbe9sNeJBM2g5AZxSvpgBGteZ/sQNgPclXtVCQCIYjPium
0dBD/Xb9b55hKk7kRMF1dNpxvvwo2M+LRBIvS44SJzYytikTa5EHtefX0q8+Vkiq
Sp/DWe5ySCjL75QTeb7Bu1pBnmAc29SO7uSMzicq3nvDjtQxEw0XJrSwDH5pglMv
IwtU1JK+Gxt+FrGgNY+kgHBXKg4mwTtRcJk9f7rl1FGYViR13LsU7/Lo6bm+zVMq
65AY9Lwp5Wx1ntvFkSysepDsoXPsfkHMwTpSVyNLRU5YPnd70LaMwILTmAexywPr
9gKJoDLAhDZayOZc419ExkSi1sj3UNwOrav2wBIvBqQ7vY5zQ9GkfMOiD53O4WEp
JBer6NiMm/7J4H100WPj3bl7Y5P6Jv3s2DELLi4ar5Q0/SlVWWPhHcWTj29H1yDD
Zr4GEh0xdZT/3I9EmZZtCl2VsnBgEiPKY13XrHD01AzPMLCWXVRqycndWVsso9Ny
HNdiTgoX8jqEnTuc3QfTw3AO+P/yi8HZ48nIotU/TII8UKTDu+PGT8b3EKN6ER0B
WGiPqTbv+BHXh451xbzH0zPQmzCTqfUS3Eudkg/r533ZluKE+NnW2vAk1jgmHiTk
viSq7b8w8vppuI55NoAuOb/2fvw0e7Ix29OZJWVXeQ1OmjyVNmMXGYL+Jz57TvNk
7byNObVN01pIgkOO0qbOVOI8sm4mAPHvLS8QWmk3RUBP++ZVrDGcfm38lZdvXTYq
mSCeRvPgw6asMmwITQ/E2WKGQLjgzSJgy9RjcnFEsir1cM21lVLuoJn0BncARV8O
S+JesBZWVIFd/9PY7CwsmUkgRSMGNdZigUEQuj1ihnDMY4zhZmLLIQVzi4FvY415
+icOjCbjsM9fVobiOz4MoDvvH0R6rlt+6Q853ZUEpemjOWhpb/pP1gu53N7TM8Db
yZEMVg+kK2XKzDs0bk69Byn7KUr5Cm15wKVDqM49hMF6Trp1ApvpvDisqa5HqA57
eQxdDI7TJW5LMCjtN5qDO2B/SPdnJTjTriRxwJMWgoKfAWbm5U4zXjIz5quebztc
8AqMwkHl5UXzKK2bj6Eytg5mSmOK8eMlEepE9uGM86o22KC0itYRTDPX5oP91PHZ
sIIVrqboFSJ2VZjeJYjN8XTy9rrlPeIOHUhRblnHVBUpzJwQdk0youie8ekh/ooE
N/vCMNraMLk3KhwMGrPv/sjd6Z3SySO1jAhYdZhjdWgLkbYzeIh1uDQgvvJd72yz
R1b1U2IG9zSLoPzTShmkfv7BYKsthHjDcQiCtmxIZKna66dqkd056D2AcyTVSFma
aAP+jt50W2hx1oIGugYnDMR9lC4WwTWX1mGakJ3LdeBwy5LYedHpCZfs+V66gIrk
KmLS1Z7q9cz0LiO1Ff0UiAkAR/yuNti5fQncPJG2aUCCXMwcs/xtZ4rJ3z2auAgM
tWUk8lUeEqITBCZtaSMI/DDq6VQhYXPFGbFw0q6MFPHx3gnbx7CsOl8TnshVA8Lu
ZELQZHGnB7PYsJNBDl/smlMB1xZyNZ6lEDELECtgHjiYdpsWMDkz0Wj8wio87+ty
0udibp1/43sT3asOF5PgXq2bav6Mb6/tJenbuUYUge1InxwAuCEdNHeg5hZJd8K9
EOUBrjlZxxGjJCgyBsZO9f4fsA9rK5AqjXHEAF/cxh/k2SZTSd45tOeN7XvJkQj4
HQWV3NGeIPZsIpB1gJ3Yf23Xyh6Wh203GUOmtq2kwhO2jQLK+4FqvPnuocT0rK17
oS99cDs8Z6JbXGnjSveEMdRKxfUHhZaUKvQicXL72UB7EYo8ZyseQ/agDncvxDcI
6PYsTUs1TjLV0U8nbqE8F/UQvtxP2kwpvALhxfW2Ppxw+pxS3k6c+t6OjS47gh/0
ZEwTEZc6oSToXWLXpM+aCzeXkP3rgZZMIbUlvJsBmPKudoUMswBIHSI86AadCi+0
yvpXi/lCSIADairilJAoff+hutpG0RhLZC+KlfwYLnkGelm06FHfdBg2JqAFCDMc
CrmBsLxDw79uusICVmXxIVnF/LDy8C0lpNgUDGl5AN+aeiOjKHU4H4vTBrnJU8iU
PbRswza+YDg58TEbe/XI6rtA1z3QY2lI+QVNyYHhEsahlOcfydFuRamtQvS15mxX
yaEUKegsdQxpvifkYMmMvwgO46q1jeiYLqiPuowJqt/D02XviTc/xUbNeiosmyCH
NOwIj5fnq6xmvnuTdbyLd4X0Ygc1lw/dWOTRo7jaIjzM7zeMs5evm1dXxumdsvbu
nCm8XiId6LAlZ+6P8f6Z6Vw59JpNkimVH5mheLumUZuy7r3YJPamjUN2nxwPks5q
LzgEHXh8nphW1dKwsEDO1Wfh8zPKp9NkjBI/NmXSnQWuVZjKnbz2105fj5cLc0xP
1MtVeBMLW9Ib5fSDetWS6H/nfuNAVBnWUSNBMWD1uSl1Ol4XMN6HrEXQ2C6kzrWf
HuG7IPtFW5KUF29TO0bOSySwP83yz4TKDgDJ8JJfxSub0b55ykVL8uGyeI5osxeh
lJygCq+vjTY7nd45wnRXh3b9uWKf/PypTsgla+yrh94fbcAYLdVhBmQEPPzei2Nd
ABDb8ZYjUQ3raMnlHQgLRz5oZJEVyU39mrBbnZcy3xBRTeh+hsYb0K0xZi0nY6+C
QmQQRFhGZTbYRpJFC2Mtwj33FEiCRwt5pTPnmQFXg7XQvH4OFmHCUl599ZLCvrbK
yDnz93NDfaBetIJBEh37PM6b69lAWll2KojlY3TwH716YkqpP46OjHjEgEUKS379
lK1Kjv+u/1qy6J31i3VxzenZql+J8EpcNMrRxWoDBlgwrjDkp+HmvgrnJbPUE1rz
KsSO+r0H/pRIszobSfkkhDLATaYe5Ps/Hc4Am0OrtffysHDy5nGayhun5CNa0ZDz
2GoR4WgGgnrEuh2BEcYw5r+cUElX4x90ebx6okBX8XCuK6JO+/1LNzMKOWg+T4yN
C1bV2wZVjijGSTA1iNOp3T/IGmMPT6zn7AE7mdgwSE1Sgsjgj9tvLBoXsxt44Edz
NsFhwvzTtNP9UTR76Y6ICSMomzMe0niKiTvxJQ/sGvV6rNsqNR1RbdO7sVQ8C263
eT7WC3+CAONp5bmB7INjKrGno8kc0A/7Z/5VRKWD0BvW0zNh+nKfdOW7V9MaVCgY
DxHeNuWQngbaeHsUrB3H+oSB4d2Fzy+YsSp/EDC8DtsEiipPxI0FrBoVmSsNMZu5
BHEHAaGBC2KJP570Pg3AIlmsSaIU3QPjXDZL5aKLmurgFbetKHiSnReXiuAWoe2j
Zlnh4yAvjZhlyhxc7tgbVmYTrsoZSeX0CgcEkkjKpwgeMPEFcYdGPTLxDU13d8VZ
R6IzZWZhxLLVdYoHFIawlZMNwh2p1Gqu6+tHN2t/PVrh21Fj9a7SwFDZJ3ev3Ljz
UtVr1skJ/ZAtACbtstxD9rFZP7SGb2D8G4qjD1NQNOATrIHNPe3G/Ru1nZ45lYJt
n784ztmlWlG/6vL164zftvnSzQgV+d92USklMV8MaHxTsoySe1o+GAsIZUneL0A/
LcNLsMsNV+v4R1WvaAS2aF5IkjiZGsAv1BlMo17R+WO3dEDULcpRaHEeTCYZcaSq
SRxGaKxKPUJA5ZtpmYi9cZIzhAIiZRmP1BnlQbbMQaSq267b7RMW9R+z4PDUnz0+
XLnYJF0N2ZL5Hw8MERLrXsxPfbNXctj+XONRGmkQCO/AAHWuJe51JuYASMJopZHX
U76re74iRltoz49l2R99cP0iIIL63mg/BWTy2umxGUGXokPG/bjDhzpwLsSfoCMl
4SZiyd+9Y7Tal1NFfma7Jekun7X26GwFJlAELTrmY8lx52/S9QjJXvelJiSzSXYA
VdaJUlsstGC7n14F3hOfz7UWO7f/iDS3Yg9B2EFJDRT4MCMaG+2LS2YDmYXd4MvW
TcL3+zE1xug+ZqaMwDqgChIu1iokVwhXLEFPzC7ujlWzGI4QnQF2gbphAEwOCuNx
Wj17zLe2flx7Lib/K5VNb4ipcHUnUDBKVhuOxjiHyoffAybAedMcMIZlvrm8Rpgw
/yzN5HxyMyJL+OhYADYnrlwItx7hAL65i2Xb9EUg6OL3qFX/2d2vndT2RNwYgM+o
C3rOJusv0rNXfNzLNpLFmGIWMtfJfbPmwVQe2QAzYEWeT4Do8Mhylk4Z49JtzW8c
s708KxBEP2nl92cTBMRMiUGfwdLzNLMA7viT7uBum9/HKK/dhhTcU546yrHLcwxX
8MU5Ds6zvCrqjVYLCd1M5PZL7Rwy2PEp5tmz5UvqcCliQdFXhII7Ew+rYPw5AUgv
nbJnfFd4ZxsV0lbrWWbmoOsG0VXPq4mGrd4IhROsOfztpPBF6M3YoxQa1gQoGBad
URaPFgG0RA2fPwE2D3bHWCL9fcxgj4vpTZdOe2pWVM72QhALGVNRk0C6uYdYWgdP
Hoa3UPThaxyjCI7VFTFY1lnsb/Zo1AL3JoIQtxgaUxzsJTDRpE1Z7rDsRSwHdbfw
6THxaIE5xLrnxXFONHGSQh4aMez7Wc5dmZ7yV2wuv+D8RgZL1znmEE2Zg3yQJRAg
P6Jt16g4+Z43PgyPjfLBsl9MiJoUK+Pk8cY6GpF2L0HQqO7fJWDo+EgMBwyz5g+6
FOHcqLYipCqmkmRXC0JqgTWdCfkAdRZ5iC3KeXhq6WC4c+gLbcseBl4ymHfWJj6W
D0GXSxn5NTMGmaDyIwh0gMV6+mlXrx8dssEogr+kVoDHy3rFZsbUMb8wi1/bc/pJ
B/611inQqPDdoqy0Ibu8UvsH0guc0tWUY46AGO0s8N72Xelzd71+yUqAeu7yLIo/
/NPNrBeE3TbKLaUluV4rHgZe0pz6NjGiAh8/SceEFdc9MfUgEHnQuiIzK3kChCXL
iuGDsVOADA0Er7BTsrzHhS5NiHwn+iGv5EtmfLqrZOfuw//HXQhaSCFVXrMH5pIb
qG7RQwmUWTer1rNInsSkD8N/IoqcaELmCYyuYWWavOOJ8J7cmWyPAA835oRKubdp
4EFvBLUC8He0IP7pyR9QAMzJnCA1EV+q+t/kaWU4GicqtuSIZCfI/fRCTl7Xq/+q
IJ6ygnK8EEo1Xo0jToZAnL8gkAbU6J7PstFjWZaXerx0NT/D6FoyhnBGTuUEKc3B
Yn9/9en4JMjPPfJV046dt3WD7IXCQssjNC+bgAcKOd2X8zKknHDHgkfUgJbghI0u
XgjtwarzlW/YwrJToZgVL7ZsoNLkG7XLV0+i+wZbcVxUkCg86qjlESKk6VCTyJXh
+L0ULngy+74ghlTx0ucM3yXIyOPpbXOkSfWG3F5vSGFq9oqWsnHYpNjx2zpX3niK
cCaA6f6+XTTY5MfmvxEtGJ0UWWY7maaJbPekWhv2iN7kPpbXOMGd7GX26YwNtHXe
tQDpGnbmOu9IqMWgBeFTMpjOrq2SrVubSww5xo0S9+iDiJgXo0/VHMdiXvxl3Ffp
M0/DoVNkflkBWw1ZTgPzYO/vkPW1fk0HNNHiJOAnRT+cD6J975hPvUDZzGQyamTP
Sv8MJmvaBvJ8sEv8FhuNdbVuC6JMpJx8sdl3PJ1897W9SAdkC/1RrR7TeXKBiFEx
TRkoVaCvww3Qjpc4lFl+e7QoP7uLxiYTbcqOgeuDZOqsAV4VGkXDfzkq8zCRz/x7
lVq4Kb6OXgyRvNT6HBChKhSb0cFxnYf8tCUDaPF0EDYFradcMHTIlvQf86rePX4A
MFBuLk8dkdm3HMYSvaLKCz2kFQBPZnHWzEDeDhjGjELjXooZiManBhzs4POEL7g3
RwC2xnCwsxT4J85cZ7pDzLYkoFx+vhcxB3vD+FEF3QzeHk+K8oO1+HZPcCSykT3R
npb1pF0ajob0aMGLw52iVBjkWRaU3IJ5Q5p68sA3e4tiH3n815WL4NBe+Eza34PD
Y4lj7grakpalat/XJ1EH6kC4mnH23P8R3tBQkMB1z2l0BBAEhF0boP0EDuU8h6QG
wWWgBJ79Z/0SjtCFsOcgsft++yRf/Sn41vtAdXGSG4+JbuViqvGpKKwgAF9YQ2jz
EF95J6Hd5J+f84yz7yVozx6uPX0ohw+6SlPOGQIPZIFtqfNHRvMlqVIwMXf307Si
bnYKpv1Hw3OoZO9aWikKMknB5qHTulwqAh/dZxTxg0v+6gRZ9jGpaNBMbfPdCik2
TgHwaZLP8nZQJMbge5apZ1t84tP8OKHGKpys6BqhH+JJ2itfA6D0Y+WNY/eZoNhW
Xh24xJebufBawrBggqSqowQ3V7oQ/OVvAOlGsSk5uLddG9wjXaV0rRyEjr0exwwt
TQvRjtpqjgA51hCHs91DiLn0yDRGVjrS3OV5DpK4ImmJzvk412UXzfB4IQCHs5Rd
DCmXCQJE9OayETRuWvNzrO3wko3FCbcKLpZ8uZZOVuQACR/uTQdobcfXhXcr26ru
UmLV7GIUCWFh4+RW//mxgu9RXYyI2yfEKz11DiGiZcPs3c6/xuvMjkJGhaf+31oZ
xSXQF+PBfN3+liYHXj5pq45Pu+sKRaSbg4uh+rEkEYeWQrt5XWyyK9ja4VP5qB43
l7ZzsCQNrqHE/3VS3/9F90iegDBXysgLQAhhLhB9GfXy5Sk4IrOyICyzBUytJdWT
aMC9X2NCj0njM94t5tuxODuJ/2YFgGYzTkR+x8ACD25fV3USWj5/R7iNP2OtyKwp
Bc1ct7xBAij74GZBBz79+AlDMoC0cDKTbKVcTOCsIgt7pCe6yBIdxp6RIEfYE273
iZ6y+eiGuurNEqkoI8/kKjgD7EEGpoJ3vRpPYPiAaugMGQi7Y1AklweYHNuFK9Av
nLdgBkdK3jj4FBMsf8b6ZaF1BsCUAPSHWRsI2iPKtUNu2YPllyoATZR7H505vO9P
/YE1Aub+Fx9PnfGclAXbRBdI3+HwQDDYAWeLvG8/Gjxptbj/1jBWMub4LpGSb+Lp
5sIRRyJ/lXSvxDozebuOMmz26QPlN2nM31g25qelBKhXsgn0IbDdlfN7mbt7HKgF
pn2B9POhbJFFheQtgsSY7R+yxbYM0p/5yyzmBPrIFlHA33jqkkWlLAK3BJPcU+yU
01t0De2DEwUYckiq55o6pC0OK3ZHEPk513TruF9EDEvEyFinO66txxl0nlX0p56D
L5nVLGmpR5BKnUNpYGWq8Ejz8hKlF1VElOn9NZ4a1+lVY9oql50UD2R73hFuCtgB
K+r6e+zYkokxuwHZwsD/MuqgJH9UOPp+k6vqnxLQP/ghtRwAjb6+XIGrmpebxnEz
oPo2gIv2ztuF5WKQwiPrYLPrmmhNLmdsQaKBxw/gJqlHJvxEJrsG4AhQy61TCShU
aUjy83/szRGOs30iShhibiElvUlZZ+/sl3WXyH66p3WUqtjujOPulsldpq4GgEKX
DKlTxd/rMTrObXJwktBBIiUJLBdMez3FuTM6mwig0V/dsvQKJ3DFkSxmQw+nAF6B
EWIALUdV/+A7eJMMO9HkqnyUjw6XyZl1oyHymXYVT4FuGKI8X9c9gHPwXPKW8Z8L
M5ATdzhzdao1r3TEZzzqhkVwUh/60oADjSW+a+zrw2hqnua6vG3D5I422xWq3adG
NwVvOOoqgmwLQqI0+ow6+u5/CpeN6raVePpwNRLCO+uk8DkVpB4w0M1pjM1FpVii
m+B2Ype5IaI2Dn0EMDHv1eikA2gE1EabomibUXliuKYB3f0Vwar7gXewjyhBa+9h
makhmsICKuM2E+OPNJgHNArqFEDxTEHbwU9uXbBa/qRVUa/xFNslawTf25HMXKo+
RbpeKBxa216y44bTrspZ1u2olfiEFq7zdgUL+PogF+9EgFZJp5iRgv7oje1D4oSQ
TD5d85YhhB59XPFwZ1llW81ZATWRdp1k0pzZy7gOZc2SnKzgWlSWLB2qZtanUjpo
WUXuStyIlIXllo0o/GM08K/v4mD3HZYt9zbdnb7aJgGOjeqT37E2jv4BY1cOPMdX
Y8I7kyhF00hLZ2QQJ3OYCz3OODqShdBR1dm9PccoYRo/guobspqvMOVlh8ljw+5R
BCpkagqvBye15EftItIB6CnqD1vFB/l5++20N1lMXldrI7+/+wBMR/4/wjg/mT7h
PMjPP9v7OKHm0+zgDTCRWCWdJOZX45z0bOE9uPk0cktEdz8FuV5Raubr/S4Znpmh
X6aRHZXwXOR1v1h19RF9dMqelWOy/mPBZ8B4Y7iM45E4/u2px1+XfGBte7T6JUUP
XwbLyglfPOx/d4DBvWzRzCSWbmWCU4/RSottNUyp5HOFPPO/8vaXrJkGBiFG2usW
vDcKdNpbcR64j9PTQeqsDrPk2asXS+SEWtuHxbclg92z9qJ1Ft2Fp+SRZrskwZB8
vQfQtRip0q5yLgCrQnUHiVMA+zzi0G8RB/TXRaSH5EXQRF4l2kEB/oR47fL8ZwU0
fhdTN6gNajFPFAZL/CoKwKzN13OdLTqPnQ6JkL4ajgRBsO0Y35kbsPnFt4l/3KL6
goz9Vgc6TqxsAbCNpHF0BqoPshE9GacFuidWVUhGqxPUeHxLXKPZWs6r8lckclEn
ipPWLEVvUeVsjxhSPnJIW9Y94c8eM/IYrMdDBOFhj5tPOtrRNiCn9j6tokk8Qwt8
1MEDj5wawjQQj8+6g5YO1vOR3TOSoZ2QHjOJnMt5K5kVie61ZFgcUMsgZCxF0P/S
jahCXS6aSsMwR12vcfpQ1YcsUmHRx3lOme2xR9EtqY9DpubXM0uCfXt42eRqVPX2
N47hoTMNB9v+5PIO68k0SVLqzZZejREJsi4be7+QPmM5gl1BkW0lDSQHXhTJTTPs
2IuqphWRYn5fJmPU8C6BiahOKhUCeLj1Isehky6H7O+SajlDVF0Wsx4qsrHO/EBr
/ErOpU6QE3X5bKQmh1RBLOvrOKL2uopAu/ita4V08KsBOBzZlqtST5t2fpTJQVPy
cQzEs7vK7GsCQrmetF4QElCuUQn7N1uFllqBEcFqGXKECHkkEp1Py9hFBlvbfRFk
6mbMgQh1yQxwKCEYwepeZoKy33qRfFx4Lg64OcZ3xTv6GfOnfLjARSoJpQZCenye
0wsdwm8ARONCpyohiMYw6TT3r7/8C8Sp2qwGj3KvI9KDKZB3I6Pofn+FKkSiv0f8
dx1J22VAlkF7TjaQF3l4WgMiSJgN6tzRjQDl7Kw3lUvFyaw51JuP2fsakGTUcoKh
TRLfidi/OwBQJ5rRTkkN4WyP19tX7Ui+A7nct3wTkfYlz1JQmzY6ZQfLxNkPp+C0
EDRQUwmaoR+/bV8aR2UXRazmic88SLhR/5lsTRomUX6XpywfIy2WoT2/kqDMQI0v
gGTMshF2uV80wX1rnz4feFwm45xWmaljIuW5T/fIoDUFVJqIspAaeKqOC0QgDNyc
BXFaufqLR6pHzSA6jZ7v4rOvdKsLp70Ep8vJDI/j7Yx1MJcdgLOsEmbTg6MUJtYx
gT9JA6NMgK2FLi1yj5b8LGNdts6K/36lN5XMuoBBjGU03JxTa2FNch8VmSpY4/Ju
F5vGGeM8l7DwctdIHllEDVSkeVP39tHU7jxF+u0xN7c/GL5kzFObWq/Jt2q3hfno
y7HNHteVV5BUVy5t/yrR2lKgRs+1eBk+ZQKOG4nb6wT7oOKOY87vqnv7y1J6m4fG
RJWFRzVGbr+irP/M+Zcsuohh93pui35vC6OrEnzB0OyK/jQ9HPSDs3um45ZeqtJo
jvScMZ6Ylk2Dszfd4aEDXoGeVDKy8FGsCkyL1Wz0jAniBZVqftMKe5Girz0lvqPt
5Gg09vVf0+f+FuSG1/TbA/tj0S/v/Z3GwaeNH6XR21/twLoTJpZAaBRxbltz7HJh
RFVOWxPWeMAonpchDcxMCghjrAYBxh6DWsuUWPyVz+yFewZdgKeVGHNFitHhUqMD
vwiQgU/XPo9PyVr4JK9+KmKHAhOLQ4RQR5WYFCtWWnY8Gdo2MUIuZk408fR4vkE3
R2/uX9xRcrIJNcRNeFD0w3Vu9neWHfQXz+OplXnR1R/Bdr63mG9EENOo3wYOuNIO
4WO1w3N6TWCIySslToBgNQtS9es3SMxodbYb7kIDxRERkzIQt+N2Cr1VHCrvC4Th
SxxwU+2nBfupgHv/xg6DvktA4bZ7uVi7Nb9MUaT680naM2aGZv0pMCZ9y3137+Gg
B6u5j44Appoyva4azb0Yh8/2pKbJNlE36ha/7hpu27TUuN4QA38giVizXJJ8Mz5i
hdezHFGEsDIIL7os1Yw5AFRLFWIveaijaIhXgC65pjmp2UeUvL7NFya8zWfzg99a
LBxiYe4zYC26h3gH2RYoNaQpOuzPnRoAyoEYanJ3X0YLh+zSXUuaJ4RUxNPfkAsJ
CS/o4qExbh4ztStkYUn4QjzdIOvlFnIuqluCn1L4/7NojFZ37OR1xFUG6uaxQWLY
8ag00PFa7TqGqDVaJ50HRl5YaqC/9u1l7hzjMSbwyED7sSUF3bWdilmZI8ASoRBk
zHyhacE1VyJ4DLzM4pdHeJxWfHIUDeR0DQe+fPF6+RNb4ZOoCp4FJnNXMFYf+NLE
cWcaMA41868cmjoz+LZU3mEnCQ4Nrx58WkOHqMiJREVfVBs001khGb17EI1UsYTG
ER1yOfBpuEmrZv7irkWZCLJVunGkSMPGTco55lAe99pJAFiMqZUqX9EMb8DMCA8S
RTX77vyzRMMOYn581vUmtqfdVOlYgVAu2YlAKrdT4IXCgURhqEJAcoWl8ryu7iIR
Clb9y2yKYgcqmUHED4uKKEU75sXb8iJue5ECbZDp3acGQG5ex857uwtkdMcB5jLD
Njl1fHnEYd/gwhQcCUqv14gla7tmrezv9lUOu9djsmPl/DrHo6WjJn5n+ZjTn6pQ
8jGimyy20CgAVg3bJ2kW7OKMOVu6NDhzgAEa8RSMKQKOwWTh2yjcYS/3edj1abiI
TUto15QFt8N/kFr7CHkAEsUw/riKoQHhVxZcAEMoWfzey8+1f1BtDjVOfJJyjfa6
MpQanKJd70MdD1Lvd1I2RZ2cRMbc/tpdepRAxc4Onx5lufAhnHI0/jPGJ4BlBuej
EvdFB5ILxOo7+yLy8IBJfqmD0zw+G+qj3yj6Kl8gnG9oXZTB0jGnlHT+4+jZsgv6
io5qXcSOq/nrGbyKTfkT3DuxpuGt3GPYbBjANhAdyx8fpKO3KSX8EKlyhYbaZ9Z7
ifFlCDYtMTPHNuacuGHkhuDJJx19bdDcyNI3jnR3LVTBGSTcDRtzIcuq3FtgDlFk
3cbUUMOazpi2hPcrbybNJObqwIHBe0h0VgByNsGn+L/iJsZqONM7PaOUIsEDvpvW
BjWTYqzh+elB540eRHMC6J7on/ynHmFz/SKNcEdKVbsFsFPE29TFaFeEGBOmLAB0
YetYMUsw+U4aeXKq930n3o+/WTJPZ66245g5seOqUjjBeAuJSmawXC0ygn+u1QOT
AlG+eWVJDquvY7BVtZWLE1bMz3ULnJZqM3faGWvRqUSDnr09/3L/3dxcYpqMjwqk
7egJqszzBNpH/uoCwjw/+YwNl267gd5epLfEso87EtXUAyMVcgd1tlPnho9XJpWZ
JVXvbkQnozF4h9gDL8yH6hvi2ijvIVjCVQIOIG3KpZDlDaasH7qFfOEEpzY6Zeq+
OZuLpKXy187r+nR0qFo8doRztV9uW8DItRn/q0mEWoJVnNj/uKouESY5+zAPFIbd
rXzEm+diKqMLuJzgS/tUO2RBibSLmpVwmXSHnxJQeaL3xZvaOy55GoU9xHl1hzcL
NI7FyksHsbYbx/WPLSgqbuKl65GGrZb/0e/mFU43vRJ+1kcjQcVSrzs9xmUkoq5N
fMuGqa/qJY+WPUvoOaXEZrvmnT9Vjsk3xJoC0YtqJswUdEa42XgCas6q2THbPP5U
XkkgETLN48FJPqNEusmZxhVjrindMmt1RwVn0nIspBeW1EKzMaOB31OlEZEp5ab9
gwgpiAhj+JBCkE4z1KwtpPGFq/EuIPeJfbKLvQ5aQov7u1Fp2Sxq/4Dl13y4hKwc
7bbNUykfyOWELS7nFDMrukYC0gkU3w6FT8yCwnb89AclntahkghrvdP6eP11GtUk
09SD0m224/m4D9t4zu7f0e4RxayKl3snnC95h58ZvO2tITWROyKaPgw/3at/ujnn
QcLjyAYKTYPjl3x+1sNaaJaHNM+PmG9pAskygd/KVw0b49NiAmilenz1T3dHQuLw
pgLWJgGSGyXo/i/uQCMR5FpJeguCBw5O9wprEDi83notV5KjUnwHuWrLbn5zrHG0
TZBpW3OhVXcb3+6vG48ND8UdYRBmgoZaZQenb4oY6zyI4Q8OqdIYIrPthYpaiTab
DKsH15unhpJdgi+uIMEz07R1L3LkzhKUlNbM7ruJbzX4CFKad8kC6IqFA2vweMAM
C+nl1Ob+bcgwyxJXYMXcw1TzhsrpOb4OnqX3nwykLeo+ZsO5I9gFfHfwvwOR7GT7
tlhi9WoMpTecM1ktrfRxB2g6BBMFS3ggaC7bEPiAl667/bqZphRyGuo/4lbu2CLP
oYE0LUIq2iU4mr/cGOEuQUYrGnSha8AyOOs0zbmQ97e6n+SvEOpkJtmbJ/DpV4z5
lRmUuLWSf+BFSkDugbiLJiKN8lxobYBeEMDRwehL+aFclFhGA4xREvgrh05U3uW7
rWuknMrJIBcVOQhAmg+WPnbRhoasV9jVkbTOLnNb8flaS9VptH6n+V1rUSjfQsQl
Xk6r+iU+f8kXkuXcthRTaX/Hw/bsSKJE+EHBnTZLuE3e1uYrtiOir3fM03Bm3pti
7NIksMj1gQqn9O8XKfGNPPnkJx/WhfxXdEeSE16MdNZS9fkkSdoqKq59bvFaAeOm
DcIjfvPn9zPUa0yAsbj0RyIzhz84m5ZkGh459q8iNI5MUQ/pA4rN1giSfEN118S0
8+vRmrOk+NT7NsoZEukGSIXXBKtuMVEKRlI0vmRhjR4X3eoTSk2qpBKB3FGBhiSR
pwJ0lbDkzI26tzBVfYgNj5CHxYnJXN7vZy8xBI8NP4zwWht2E01+sYjYGiJkzUk3
fGlq7m2hHptJBk7SZk+mDM9/F13zECevqhfop6/UzfFLjIuF3wuvYH+rNNYfgG+R
r7P5O8534YWV+F3Bi3YYDTRyT4xzgIgFquukm9879EGQeSgIgsEHtX6na857sHGR
09bp6LdY9/j9F45STJf0re/pPHeyr8MShxk8H6Lnglu+ZtfSjFOHsoH2jL9XhqSj
/kw1ylp6FP5YYEnCdVr1QXIIWExhUnkAb423UkAILLMtwV/Ok7MyIRopwPG27rc/
xYLNHM8H1BQabLFGkXpuy/fnTWwpFDJenZyGN7cDz8NV1Yzr6cuxQCYvjzodIWhh
tTMLbqy2FucUcUr6EY1FnhUlna+Xt0wvh74yxnFspIK8C9cEmgMX8Jw5Oq7/CgFC
ddKiKCT+0eGwNQNXWjAsHVqe/5LUWn3Ibp52MsJ4ghZcM1u8b3es+/eVoSTXqw1K
ido0ygkoPPV3VOXmbA1q1Jy4p/2yhqznd3+xZV7uKwBtHhZDxwMzDP2LQ7TrFecV
3WK/D8RveCz5iaBBLsD7tArq5aj5EV3q/yp52z2jBAnmAI7WaZL8xnsB7svkWqfX
w8viHMJcifROGpbv2oDWbH0LnrTePHRCQMylA1TtpYET4EWjTBOw5Gqu+OPxWJty
HnOM1E/RBQtYvfk7Sx0F8aZtasQHtdo7J4/Ua6tiCBBjoJggpBZNPZpbkYR72ENO
uWeimy328pA1npI6DYTksbPzORgrqa+T43H21ud7/zVn+T/HyKhZpfIKS6d27bCt
AMEwmlaja+jJ6jvDA33xb/YIVm9Dtl3lLBb0+w4gOTLh+x4bJQdn4q2PcdAJVo3h
RSGnKenSww+ljUGriDjlCBwZRIMUYMa1MFlThLq9k8IaeL+7Vms2w+TLelHh1Wq7
OsLUxC3mKslFiNCtT7j/VazHCn3qg+zrJsmaOoHosS5AXSwj5ZizDuKQSj1r6cc0
ibLA1D444/ls22F16BRKvt2UQFjXzCEAYKKAtmIwRBstKMkD7fhn1ssV3iZPImaG
yQvWiv7tvQ/jBMg0E7GxL1SBtQsMNDJGyLqoALbKLY8TmHsinZCgtanlGBmZKmVG
0TbvzHi802IsN3BF3IvpYP+iFYDoXP/k9Vl9TaQboT79rQkiqsa7qwr9f7W3+7VL
uK7JXy9IGPmENk3HYXYHjXYs3ejDfRDQV9FClASG9Psx1fLYkfOKNHPwXuwmL9if
yxfh6zaLok8M+TCg4Aop1f4SuqLeDAdsSUZG/7bakgGf9ae1rxJYTU3mUsqfbNFz
5MSDCYFtUUbULp25ZmQHIxtpeCQsI/Mq9kIn6PCMETkn2T5zOg6s1wZeC8V/obRz
ovGljDa3Nl/KL3S7JY5aVNJvYFQlD1H8A2t7Hm0iD+3n+pQhgWvxKdKI1pNezqqM
y2x8BMMznDAOFEDDtN2pzxkJiIRe2GqgGiOty/RR+Xwh9rfTbb+rkbEL0p1MwrRx
S2+zgu9t/kS4s0/xFotT6KOkt0MbEsfrd/TP9ryb6jOGG650cGCa64R5N+DpvhXm
h+CuIEmZiFWmTl874u62o4THfoDzZigMKzzj9EfTUdrDvyebzbA7h4VkaHLn/yKB
KvRJAlhvW6vnzi3fOPTH3SVuJfCrPvZ7s2pIaED2cjSSHeg7HoDiYj6frmA0vU4Y
ZdiTFCFGDImEDQjVZG4u7jQWwYLzH9le3DKkuYGrdubkIrjrE1DgPiU1JdFQT/Rt
1SNrx9s3b/eicWcwkOT7E8xNzm9FlSf/2SQFmlr4y5IvKx63/tRA6CX73n4CJzjC
hViSuCAJckG+36dgA0UgbOfpckV+9u/Z9ezbEWrBbtEcj0Aniz1PFGpSQfuvVBpt
nERWsr55wQjbcERa/B7s+R4/5nyfAsMEQdVedq7hRBYET8qx5JGwSG1Q6b8NI8sq
V3CzvdivcqmFKqabF1P8oPMYbxZYj1HT7eQmK+K2yiy/BEKYjV44V5xIhLoDIBFB
uQd3U4Q0GP5JvzdegCLEcNpIatNbnQDFOi/sR8o0ng4/Q1v1NBw1fNxPwyrWkVUq
pef6QY08kX5OMtXh6c1fTIj5TcK+SVtvUhMCaZ5TyFR+CD8dvlX+hCag6jCdlmOR
v3brAnx3xu1o6Wn8A2KlQ69omSEZ5g5V8TNqO+4IXGghSgd8LkqVSrhcfqM8SsCp
5ze52m0YXfr4V8YVHkK6GPF+IerJiSg4lUpyJUw7SbL++yJQlfSW5hGvYeLXlW2N
YmtTH5WabO/MbOm967RttF77rNa6RXg1opR4U0OQ49rEcY6FpQkDxtjnKD4fYJsd
AOfQ3IqHn9ofJXnlhruk6DwB3T9Ks4H6TSuXMxImZ7VcjEI8IHB7J7/mqtf0h2/f
DTgjybgqswgcMfh3EW57W1HPsKa7tH85rilc40QqyOLV0ofRif6KDcubnt7KJL4h
uZZuKJlG6l+1N6cv1GcfrTP+J5uBIqkruE4tVndQjZ/FppO4RV1a+SsCbvMZdiEv
e0UAA6BdTIQnGAuQCO0v2V376qlFEycJNvPYtJXDCKvv8xX/nugku3+vXv2RPhCv
lE/ktCjEd0EbfZmPA/8v7wxjOx5FvPQs2RnnvRDaxwULqaMxQ8I7mcUe3hI90XRF
QJPP7tTBcA1/1jwT6Ul62pKLQ5mYdWEpSNIC8rGNPlvfLG+zZ1YMLZt+jj+9dLsY
ry6DI4IKpE1etVN2RHD1ShmiB1qKeVtQ3wPys7PvBc2s2VlNm8xK3axng79xuH9Q
us+2jVJ0LBgy/7oSg+qwAl+/s2AvSoXKR3xq9X89KTlADkFJuqwLJddGxloWDidX
ZxYom9D7sYfy7qM3ijt9o5EiiKfmWFCpkOeeN3r88FqF2aRCKLDRFrgRs7tyXeeJ
GsXPdtydnPO8SsahfT5JqNnUvuNDkxq3hCCUmxYgWkxIUGMMm+Niwnylir8mzL4A
VZDp1WPKBF2GooosYTO60AaKGDbOepL9POPa4vRnoZmJG+yoGL9h/WRp9O5epLfs
8vwaQadhIKM+F5LRUOaufJN76fq9IpERPI92CMQoNejMwsXkFpD98/gspfLsWX4H
noCucij886bLTWDJ3CpHmHVhSiPUt91chJJs3SV2fYyrpciIaG8E0tPG+/W+oBjD
vD5/4sULe1OGwqUNWcduGe6XuFrQBunWwV0i13FJR5e2X9LnnoDf7pJK08LC8/VM
DAp673VB4veVJzsLJg6yPSHMaTx6Ap9ZdbJod4fphh5R2TMMYeXBBYKklmIAoUY8
m7vqzp3fYvDX7WX1hyvdjziBBUWJVDvqrQI3xfSLRZ3YpzetgFLd0S5VwxvUkoHi
7yXs0HDwZ/dxAzPb/YSSXEfpKoSc6Z6b+B8MeExgRX75WTz4eN9o/e6JIclrpgEf
98X6FIuH9kEVZu/8LWjDkBAAake9PedkZq0mIznZfKuUK8BvaLFC5nmAYXK87Qkn
nNxgMtjcJCcQMeZpw1GJ0UhcoJGbQZGtzsljRvgNET6fKf2Udan6Jz6FqIha3ghP
oX2GF3wuHAZENQ6RAwgt3kjsjHnbltKXBfvqZ6Or8i9xgU8POQsoKSqarlkqaEUg
IUGEaJU00Z0qdUAlcXGMJ384ojngGxNIxBrNUIQApt5e7qKIWIf0q/N8WRlRvxOB
sgDW6Dv+u8mK2DVqWt3DScnVqOkmSiDTLpcNaebbK0aI1j35rfumRtKDg9U8WCAE
s/EWwIYiSpVts7yIaiGJzd6nu3E1qd3rKHPjeqaKcn+iZynrMKcJ3rC8P9fO52gN
URWuCtwimW6g+b6TkXkzJUJiee2/qiC0An1yyWcMul+XkpfpVynsjYFgv+WbPKRl
6pdjDRwP+sjFXtxCBU4EMZHGMjb8nLyH+GucK+fxzj8D12mw+cKjUPfxUy10TAw7
ZbOQWEfNF3nwumw8YRIC0WIRYu2wNAPjZePY+bL1qu/1ldKWlYZ6sLrU4l1kXNtD
eIKSY6UjNwt+Qml3ElGyoDVl8VOEipX3aOGLYoe+o64wKJZ0hDvnHKNefXMorJS5
6KMQ1WB4W7mgFX0Lito/UMuqeqjwe7w2fJG1X7Sfj5tuCyEBzXLEcP/39aT0OO0Z
nq7mRwNk+2ifjBodrCm+lN2yaFbdd3izyhXcHWhSC9BzoMxe975yyMdXa2AvSuOM
IbAWmSVcNY7W/ra5Y9UNDmEh8B8G5tj27SuNDqrInhPVcHf0jNuX3V9qqF3xv58i
E6UKFuutpVBL/FUYFv4gHo2rcc4VFEvSnplLwgsDcDZenvWN9AMqWv9NgR+u+ipL
qCAxJ1uvJHQjPBhDk3cmJr23+x5BCeKRS+O7B0bDHBNpgkwurSgQ8AKd/5uHkXKK
vLE4w32mWDHpBjKHWBdPe8Oy8QrDeAAK2wz3ywdVZzstOn31MqiVnOLhWnOxKM2M
sTnaHdVBBkVJm9yMeioLZ5ta3YO27F+0Jrz5INhCdkldKW9wG+C7UhpCmBSGI+t7
sBM2mR7GbNKloHvf/O4RpIZ0iuWS9FhH4amGj1xmQ+te/Zeioyc0EnpJYqNJPXrH
ufv9Jn2xkkKnGqyZXGYqXjJWSvO5zJv7rAgAenZGrWL6QtDqI/tG9HJllK6k730m
3jAi2Z3s8vTToBRnqYvudNhQXgUriW0tTt1pRyZsYh7X2g1RRslVe98MKagQP7+Z
e5AWlvUcPCgwvVy8mTSojdsVCxSXJGUMCdgVYUWXgyvOziaMoCcsz87QSHSXYD85
A5Gizi0zltJVxD21Gdv+etkR8tsPxO0z+nUE/9jKHVN7n0A4LAgjc0+cTLILQqwR
Q+TYSel0uAP98oxrsccZjMfZtkHuhKdYOK7kQx/3HFpRAYdJgNT7nxW2iUmNtWde
nHPGipyDgfQnuYjBqXe+QGxcgXp8glH0TCbh4HEiA2vz79hF048J2oouA8mqeL/W
ktqDHcrr+7YAWVH89xzgsJp9HhjeXqbgql75weCDdcGc/DShpVkVNgMOUApeSLML
y61rNPMOnmoO9IkWmqF553qkaG2rTwugYFcI4qx5SAOeErbtnOIYU+5U5thDJnGC
ZLjmYz4R66zr8UqXX+w2PZ8UVvb8kaqnNed51U78BTOsH+z/RKnGsmvrU1msdWV+
8LUNj57jl9gEZbyruE8rbY7o7TgH37MdaNtrayq742cloSShcemVekSC6v3+c8FT
TeqxVa1BMWX91uMv28ZrVjfPmcn41NdgV0vEHh/eS4IdEM5r8EqSDsTVhS/BRf+1
sDcUIhjrjFY8HgxCF0y4jD6R/IBg2S9zIv6Q//UBbnUwrj81kpdtMBg1fPyINiNd
0ErAGGCT6Y12MQGaPlDM/scAGFqfeH13r6N3lFXIG58KABAuGWaaWilk5hKwVruN
i9H8fxFJ4NDbQDo71mV/iFO0uwKdlbPv/JnU60QdmWVrXfw39hBbqsy3QhyfHHNB
mbAQzDidr80sBnoRnF4EDlHBmMQFB2ExzYjzEVbso7fgPiPlOXahAyh/Ekxkx7oR
bKfsEnx7+KEXyqkuQNQA+AD5vc7Y/ex7AvwyalRVEdYCQ+nShYegMfUcG1iC7/bW
1DdVlCW0sEHlemg3K+wYWcCwtJ8oahAXMyORpScz8cLPEGP46mz8E2/dDiwaRS59
KYFKOUWOVkNxfvJOnVReL9/7RHESC16i7pq+3TmOWV1jvPnf+XrLIZvBt5Hiv/1F
IOhMY84hUV9J2+JuR54neASzbARZIcp2xd9nOULh3B9c6UxgWtnVYQ0ZNyR8H3PI
1Zbca+191pRD1GIY5bwmJ63yAesyHD9nbqtK9LyeH+AYOOtagtAvfXh7Y3L+YACa
GyhjvxbyXV596BRtsJLsPSJp71v9AWEuZ93CI0xV31vsNY0N7gA3M4xGEAy++AJ8
40Nnq/LEeb+aXA2+XZkMxPRSGoAaUfqnsE8sAVAD48hulsiuMo8M6yypjZ18U1et
llub2gjZoAMtrS137+xVC2FnLxND9xHIpMtD6fos8L/Cmi4TSPApIAhKgPRbXEoT
BbF4xU/MWWJzOn2CLRzgZpKM0Spif2V3g7VYh3BdDq19F+n/y5Bvn5KWuM+jSpLn
rkftgLI0Np6P3juDE+/XEuAbtKNMNlnRavOWDnyWVYfLwA5PyNO2/cIUdgVO+kI5
7/qcCF4B4m6T0XG3lH5aoSVwSlmo35vybXrcg1U1iPNYC7FeWWS68LTqUo7J44zc
kMYz1RCGxQq4eF7fUbPE9ZUn6+TZD63uodSViueivWPP8im1awvm32DYIDK8lhVg
OfpQHvb2cG04kwR0gzS9NlvecVzrB5JEEvhCCJHu9EEXqurPMgoXdQLEHvvQznQK
VMhcG/gPcXRGam9bb9yXErTYFDUi9Lby/ehG4oNXRqGewe9g05NWlXg9TYagsGS+
TadJaNVsrmtItnWH1JGsyChoFmz4cvxUpxAi+1c9Y78q2fambD8+0d9g64E7ATwp
4KbpZe3BFYnNs3r661G+ibqkdbdpLC5UixKo3eVNDiK7I99ugyjSHaYJ5u9R6Hps
BI2UjsimUgSqcm14v3o0JBLMMdmnbmsEQMRB68guWjo6Kcwm+W4uCmwk4PB0747v
y8GxUpd36qh3AeGqFquQ6EP8aID+74bAc91u940eV7DZqHfCZEelThnwDb35EdOK
Y3KYfrpVUaNDpzBsfB7gd2cmtVpsScBtSx96T1taoh3MP+mI7g38nj8Sde8k20Bz
hTesUSSMFXA51dsogRSx324tG40uzgUeY/P1gAlbmvkMdoNND76tG9i2vL5Z4W5t
ZTv0h4cg3YX1CQmTKzrkJs+EGUwK1E6puZONV8RnuF+gAsW1JGDup2dE2NH1vEjF
Ixs/fB0asBcud95LOZQHvO6SGkDTF3DkHFsCdF/wWBaay4Z/Nx90qD9vpseXIT6G
Jdma0g/B+G9/9EoSZxv2I0Di2q/i2+eNc/VYSYlV7iEQFrXKdkOxqxM/OFx9lO1v
LEec95qjynl/cZGZ9065Qu278h08JxIH5QpwGWzZTON5YXfrcBCuUx5xuNguIcH6
tOMHSzED8lJpw9xnVUJuaChp4HC0lkrOSVZLI3A/iy3CdHolXVYCgHEG+A4aC3/A
aHCxrUx4SksreS2f8ziOnBdfgFjXywqZ1W3zGe/f8vrpTyPAi3M3NhMw9QzH1pkl
qw4lybt31XiEYnpir0wC9eLERZe7QATTHNAj8lpOM3l+AGa3oHEe4TfkkV3FNm75
2fyBgjQtYnO+kegseMyQ6zCpdEYNpOw+5fpfUpWFIvazUuiKIhz2tYmg6WbSUVtz
gvsmyluUYigACtE4oNLd9bqGVm74RIfoQDDvANKvFwcdmSpvfsS7bSfFEq3uDug9
5TbeBEtnhQ4KwBUmOWKReHnqc3iA0v9pcFiOztSoE4n+kGLWa/GXmY66XzUkyeQZ
3u62te/kFjzhVpN5R2vB6S+mVB4VyWk2TA4ELXRD00WXAAgvaOqiT+7trMon+kbS
Fa911d77a6kGoSsnsBW0R1Ea7+iV4kdaVbVc1ykeDQEMjYQzpofUGErFmH0Pfsgg
ipMOkO/e68PO0slQ2KViQdzZgmzPWbEfKV2KyfBbDqvK9J26GDQu+60Rq82jHEpf
F2eAKx5INVejXGbJaCH4H/GEAw7A6V0ch9J1j1EgnkSITQVl7hb3j9tgUFH5/T96
QOpYG6ZIdYOWamN/I0Sb+81t7eRG5jxABp7ETXvl1yRsOOmXwNF9bEV8fCZR/BwU
4tMKBmCQHLVD473GF4azMpSeulyfmMM7H14kS6L/EC7NNSpIcAo07htg4B1bSNDv
lgunMygY2nGYnS2eaIFPG7iUuaZnBiCMyjCduYdBOovVuFNP24QQk8fAMdj2maaf
Tr4i7wug332ATP2/KDbKVYu+Wy5aMw2tik97Amqi81XSPUBAIW0/BAQP1mJkGCpg
lH84GpXPNaveSnodlebsnEKc4y6uIK6LEVFkeJ0Zg9weq0sIYaS7UDkR3L/wwNxS
hkyzwg02s/aKRKVY/1abaTsHTKNpKdOd7NavqOqjMVeU49NtfT6584lcYfcRsYcq
8v7IZz/KRmYelfbIXibnEOSNeXLtleNLRJhudWyhLP1MOaZathiamsn8qQ9HQqFA
pXK+tcPZxP4SVKNmRsVLzKqtfwWwVpS5WKeLR6K0YunJT2jTExHzewt+QcuB/nNv
2eL2Lgi+TT/n6tSEIIosC8V8+sNkEzC1O5TQahRAx3g2ipkRWkiPg5vyI/MjUHY4
wt0GGBsRPQpAM7KgtdWqIxSF2rIRSOhziNhR03o+xfFI0LEfQOsv+UVItMz2LFtH
pPVKN9RLj6jVNOUhOeVpNHWiHMh91Ri/kwFfRY9offq8EslAeiiiCUmVTRqZwdsJ
kZciEavJrenKm49FfhzFG0+1V6Ka60wc6J2eijOZKLdudiCqpN1EtDDgwpHRhDuy
CdPS4gFeI2viz1mO58/+ZGUfYIxrLuvqm3hdc9fkObtfca8ppN7E4lhrtqdvZI3S
yb2zJfXS31iXfizYjp1Kms5z3iUvZiFZWL8hf+5BRibXeFvDWfiqZv6Rd7gc3SWM
3yfD7FcYE+fyQTh70CVwZk7umu2XvvYT1WRDXTyw7+tsH7u0U9HMFCrOoU/5Payr
2B8bHq1qqGWoNJNoYRV/AZ2nsMBOr9u9qcY2KQFuZmCs8vWG6V14egp8ETJtB6Uf
aEsYjKxUqDQRYc5F3diFx6rbeKVGvvzjPBe66g7m/t4N0Qhb0hmKfyA7PIaEP6Zt
PpmSkrUmL4Im6SEEh7V2poXoioLJaM30ntyJa8wrjwkBiYmREq65B/NfXI82NvgX
6kRzewRVRakXB2cm/Z83pnXZFAkTdrc8eupLl1NGNSu3HH/FdzZlQQb8bkJzFbFp
3lSmN7NDKAp38MHYCUA+y7ykub51riefXNvmuRSvWdhN4ZBkTCVz49PRtwxUKfVJ
ViRkKIhkQRru1vmery/+SOi+KscfJKUCTA2FClZ1K9bUmrKAU+YkwGbtn/QCq0y7
CrEnfduSQ+sPXPJJOZdDohL072ky7N1yveiSqjC1dbCg4v14HdIruuP2dVWKCoeR
26Y7xEhEf/qRW/RDPmE2NmGHkl2QKkQkVu91zP5v5G3VmnNb7SnlXMlew9Q8jf/u
fKcl5LsLGxJqvA4Eo3X1utg87GHwOj2fj93mPu7pmYdK5Hh9UsGE4R3l2fCMAcuk
DNRvMxRwaGRkEXeswbJK8VDu2nE0fuc3o8Wo95jHBeA7+kZHb57vy7jZtwiBxLbd
GeXgvX8tOyZx1csSPS2IAuz/WTALImvjsAwzHXGnU8Nk6ZwNccQ+YkCYNwxX0eOP
e9xY2UmifJMAq7/9j1zigd0sWejo00Iu99oFnyn9RvbZcxBz9ro9lgvavP1ZZuOJ
FV66dNItyjHiUNjff3D1e4E0QElP2Ro4TX7SdWTA0DBrXW2EkvgHzOdjDnav+z97
Q3MSxRcFR4LDYjhCzizEnq0YPxus5c/vn9QQYPs4KZNQMoLBRU/2xmjIOpW/+8BZ
O2jV+LVJPLS4bnIo/2QmEj8ZH+fcyp20lBltux2OuJrwO+bhUOOzRoDnU2mt97Pp
TzvJLlWokt1QfJStv1ldiJHbo8HcIjp9U7P98pcHyHZWJKOr55hCVUhDmDMLUUHb
5630bvBQrEF8laS+F5OP5ZN18hM0dT0e4dh3ktHqlX5lytnwpGc/VW3XTjpzo/AB
jAROndom+WGOX5HHsYAUSM1bSRNDRSHt9r4ghr2nFbItdRZxrpQGt8MGzPJuBdgW
LqshrdE2HZbYKeKwjDtl2b6W308+d6qKarU9plIMO7j1goknb8UL6Gpxkr+Yb9jD
ZD/4sv7AEIg+60P32UdK6myl9tgfRBmSiimZXyxripcKLsGC6ohhHUtGPXj9O4/U
XT9aRGCalnAt5hHNiIWHuAZosLrQrHti1XKB/+Bx86ZRVTmS/mtQP9GaMXrj1X1A
r3VnOgy/Ej/bSWADKM1e1U0Wfq1360eqfzXVDfCQboIqFOzrGq4KYY8VkAs4/sgA
Vo6Ut4qxK1m1FdS4ld5Pb2GgEoFOnOFewDHrAjTJadfKkuDnKxkCqh6d78OIAfOO
MEY6EARNuXVZ7rXoqXMkN6RHKXk6IvRrrWYWm2wMg2083irqzdQZgY2RXKHFYTFy
NxEDb3b22dCPfmAq/V4Z6uVxIhVH16HiukbbLifcLcqwk/HGvYgTE2JBn2dyIFAy
Ui9i06fINmRKa44Tn+liLmPgxpff6YkNZnADt9MIxQrPNgyaXQbj8f9Po83GrNuV
xr4RNNXt5B43amGOaqeBea/LGbVBp0RYlszUJ9WwerINX9o/Kp71B/YZwEXn/mAi
Gj+b2JHQrEtJVs9z54kKEervk4lgCJAe9l4SQQGeVnfyYGXSJ9xoLnw4vPD0WzRs
jhyK0Ka5FGbZOPDUaLlKly4DlnwtrziwZvTuqqwK/gAIENj5qaJOXMFHbcEDKTdn
7c6SJULCrQUkvR71viVLnazrUYZ3GyRj2D/mgyBRqhWyvi66f/2OKjro4OxVlyoN
t9JleBp57xhgn/nsUHXZ2ROg7HpM94C2bSQx0gpJ6VRwcHzXQkIYLX4dgTpAG0oU
qDgo5tqEKYjrxc5NuSRrxhrUwZzBs9VXmfCjTeX5Hsl804F5fAa1DmnGjf1L8Gci
VUlP/3mZa0svbWGDEEH+6/4MuvckMYIV7Y47gkZGn6BJQIAkeixxwsEqjOJFQJbq
YEdgeuKsOXgQYFOcnH4TE2js7/FQe0N6YWvuQ3JFit6yxDefj1JWA/ByHiJztNZI
X0Oc9c2k5jhs0KuBrTAsKiHhUxzqgr4kaSHtsGtXy29j3RDEmTV9O1NNr3fkQhq3
jjPUUFMz8SV8keO03YZliPiqJHroWC3SqwOsGPbl2vcP560z4w25dd4vN0dJlObZ
BT/KWDpPD+Mwh0uWmh2+hh1p30i8A92qds1dxZjiUDjQoyCi8KfXExZixafuPb5c
g9vYXmSng9lUUO9oy1pHtM6YBYmDsC4kFsUZpQqYHADYu/VXJN+EXWJD6z2Hyjlz
/0wvyiQP4vt9mOU3CoJfVu1BYWLJTVbAV1QadNb4V3tVBhemeFOdkpywU7ZgwbvC
w6GTlzNE4goah3TP6cOywMlIGXKazbQuTI9yG+GOO6i64RQZo93BVJMncV3hfN2u
tdj7xkbgy77YV59KCJmJWPWg3rHOdoK6Gii/fnwQ8yLsROLyyZsp7B4kFdGtPlhe
CtgC7LvpKTCuB3bId/23jQzMN7CaZvmkedtJneoyBnK10B+ZwDIZh7qG4OUvKKgX
vKwSTjKtPFQe0qz1svbKAq7YzbbpgJpUHthdkltwSSgdnHa2rlhN1uTuBGnXzJSw
M74JOYTfQSodiKREWM61EZFA0TdIe7ar393iadAvEQhVw2gaJM/goQ7RWe3M8QLt
l4nwuIUMwvcJEn5RBRaKRNLNF5zKvrFNEPpxBiPDdMV7BKCUVXe9iS7ZDmtiq1nX
t7Xi0uflJP/tzTfTM+GkrrSW0tfl0kYihkzoIfFAA10ybQFe4UpHQvTO1SeLDe19
pf9hTwz3/4e6rsH4xT1ySbG+qI6L2ChpnfnqlafMjHTAmhX0y5EdnBTTXllTxL+3
2Ly1g1I+23tn8BuWJdoGsjM4fMKx9hw0NqGAP5O7hSfHntZsmZWtByRxjF9kIufP
84Bg0lXej40D+z8iaJqRHEHxPAzF+GtqnJL9nqc+gyywMpyKZ5OZKNi08IJkQ6iW
dX78YO+8O+BhgsxtpOAqFUDixuxTKLaF2WdLWY3sX67YVB939k3a7mKOMWDqxAHN
KyNsM01pZNABKrNaP9pgui5UR4SOa9ny5n732z1pE+4OUKoLWxGcHiOMedRRRab2
mW23GcIlirJ+Rno9noDjdFsW2DS0GJQ2RUcWe7VnzzPOIPw+kpYEj6fSMVxWwMrQ
CVgnGcPzrvvfrvgOde4pda1I8TTWE/qNXT7WSJ63qnSTxrkFT9XOTbxHKlvbRFDw
53Xkrlp/UV3FPXb15WWaygJe3lbnRulGOyqwLiUWVBok4kW0P/+WbH480cJDkuoQ
L+mS8TTzzjrMc0L/fh2I9K37Rrrfnghl0nKFJLPeag19eLZtnfHyO+nB+b3Gg2Id
DX6v8rp92gWCsZ1kQIl+9trnKzQkaqWZpfL8fU00rAJkgNxPh9fzIV6N1Oii/H5t
iSvvUbvmIlUerJsB3oAXUjPtpcQ6cK7UUiKmlR9XTrPPGWwkDL2quHFwu726EYND
vEwgfyN8iKr+GNrZmSM7yr4alKffMaq9HHidQfZujAzPZfIvYEvk2AFJM5zkid6Y
JOaHLJYCZR9pb+hPiwqhGNWsQXalLkBVJmR8gieV7balGx3+MoDrCna+uATzsIpq
XcxqcGkoHU1sza7w8SOQZ9DBz1vii2p+KixrwNRuYpPamye7kcC6ywYIF5UhnnKn
hGGkHI3Sd4gAzqQfbad+3McRewvK/KJo/unXFH+IRr8oj0r6IeGeRNK6A2oRseD0
ykWDkTXEFv/P22ok+3C01xmi1rwVdOWwyyZHFtG4CP2iWxsHuNUGEn7PM5xfylmY
21fXkPHajdkbxRc796IEtRt52LqkRGrHmBxABpraGL1WL/4xkz4FVPvRLvwCEsbs
ykvEwXfYb+MbEcksMBqxRGyd8qBGrzIldNcVijDya5BapXxEzsIk74stnhQRm/ZE
SWo+LbNVPom0HBb1hVSQ6Dk0trgauahwADajvH46XoQPMDJgjSEpEHbMBeNL2m+1
QC0hBn/XBQMTdupdLhV9gBLF4/6P/SnrFLj4BNnlkDLWJ1tg60+wLSemc5nrRyOH
2NpbvJfHUNhZaEl7hjsZuGAWJJaVj+vtxaTJn8nC5nfyx0I4fkkW8+X8ZmMlJXik
F8ZAHszkaFCkeO7QQqxIqUH1pRB0Vrsx0N1Y8ZkR71BmN6vNH15apreVcv3xWyBy
9BEOm+DXPNaz4z5De0mh09A28UpJveWJBGm4rtiuEJ9nfkE8vW9g+kWzOyu6ed+0
iwdX0j8M/abFzr91yMOAKVfxpXKk7bpJMrndjEfDwL3SCUaSjgRun3Gse1Tt534/
6V6lJjZW8WjAOVTia6qm4nrLuH6g3rVZ2Q0UqBHEPApMkY4qPXXd0nnoqVWGH6Kt
LxGYSURRAqU3oBOO7SOwPvV4w/cblmdRUGzWCbn/pVFom00APdVL2vhcvygDoTe5
IKdKxHQ5JGSJdLszclbbw7nAHYKMk17QqHOwBRRa7WadtwrCeJuiTrrZIC1mEKZK
nYnRqeECBMqJOq//NfV/ifYPjv3MI3xQ5iDwrXvQwVAAqSJSEZZlsQtfvqQzGJyi
GcwTIR+OsPT0uDL7fIOSYtq79sbpLLFSObillvn3GkyUF9vuhvW2d2WMvJ+B/ZX7
CQWz+E0N2IO08DRFcuXGblDWpRh5J41N3GKTueSxGs+RW50AWcHrPxy4v1AJ0vjY
mSNPOp16GkOBC9ywj0w5Lc4k6h+PYWV6eUenCV1vDs6HYxGneZgtKnWrenJu6Pb5
vpATRJaZ0RaUa6m5G54n4eVB1QYXAJ4dVk3ekVvJW7LhYFT6j9YNy7PjTqmqmYe+
gKn9RJOC9MPYwNIavzdZfQkQwzuo4ZEfylMZTCEDSnuJ7OOYBGPY1/E3QQTKHVrj
sJk89Wt+Kn9ItJOOFnkEKogSeNU8OMUyuabx827zNN7QF2OEX92OSM02SiWDh1s0
4H96EbwWUTpDpG+szbB18JPUMaxE8q4p94xuDXrMdyTLN8IJo7CZgefwO5zOGZ9W
ju8+nNm4u1yCFMVHGpljXqrzTyxZO6VLAzxX+EhsecZTo3X1ugu7wKhTtoImrJSh
1rblVysLb/Num1MQpfRXBYzkvhNZzyasHmnMf3YHKYMVHm23hZN4VxiUVt7au7gj
lQQLyjN46kgn5ri11JfpwEwAKxjug8tkQ/XoMTSzwcYVrdY1tmPKXyxC2lp5iFto
sY16fs1ygBsp7uIOnRDm55tFSq4QM9ythNr5rCrPiOr7HWZRn8B2dQ1nNZF7MYBm
g1x+EvV1+dT7JX+ucs10ykUoOKquSdKPxmUcZpesy9Qh31OvuNd/9epq4UTFl3qz
vW8PEACLcLxUvC/AE3k2WflAI8VhJ9Fv+9eRzUd67bsPKbvYYz1Rqk8XB8EJSOQO
S5N9OWTN8o4EliDpDyTT8PBmyyfBoTBDAnNGWNN143cEOUDMCJsiIQTeQIJwOkWQ
vFCbH2Vs6hot8N2FXvZfoWKnmPEK4qB7OxPXh0nhHUI3N5OzmIEuRbtyGl7xOWBv
C00lB2LZxS8AG1XoK5uOOv+zf/RjtNxn2gkBnm56oIu1iceniMZAN8RKodn7KygB
0JvJU27pXt9QZqqXyomY1kNDlP7qDPq1wSZb4dHS98CAPktjfxVR5Whz1KI3v4Sj
h0alEpDVMKb0rey3h6jcEMOcIvzLBbBuwqVgBp8+e3rlyzpWW0i7VRgS3nE+0aqh
GHZoJdkhoi7ecyFzHJ02LoDGN2pUfmMUp5UNbmlmtxKmI8c4zYg+n4FrgrIlUEcP
eWw2Gm7PbdEH+AoQ6CDitBhkF+uu0sg/EP8OysqG2b+ZfbY+FNsja3X7xOohMR8r
YQhMG1ZbdGQODM8nnYmK8Dd7X5xJzGf4D/0MUrv/ghknomxdTmAZwoRKbxKZ2Jca
rxjIF0PkYFuqvbbK0jRb3wmRTxJDzO9zoAfCsowetQAQgSDqRX6q0LftalE3C/EM
BB0Bs5IGB0Jr/u+kjf0pwyqnb9XSAg439yODilxSwyJ7TC610ud0rOhFZv2nzOO/
HBSHxFnlxDh3iZ1Cagjd47OlozANrC3LK0u29vmxj+vfv9juXwywx0WL5UQab7b9
MeN7ui9pCnA4fEGvhDLCggzvl2k1EC/keTv98GK7ycvXntngLPfSmt7/hL9y5d2o
V9+5qyo7A3VbK4CUiHSu/twcSAEsQ6k/RApN+Wa8OflOJrgXwkwB3MFaMwmPOxMV
uXT1P4P9mMKNr2wHGVS9MaKTy0Vj/eTweJ0UIKyWOOBLIENilXvqBd+K/UCVHlED
ES2U7eREtXXROrScbrx8pjyvpI1jaYKoOt1GPUdaPDDp4j3CoiEBMkT3L2Pu5rs/
shagErTS5Z2knBYYmKRpJfAVhh/vu/3dqL87c9vTsl34dpHLQn8u8ttrLbGq4Q0P
dyLhCbhUlb34Q+iLYrBOgFaNlVWNWr1I2vIj1KtZBcTRJm3jSpip4m7xsXotFMzm
xkPsSmuImwl5FTXTt9g//z/q1pRv6N8N6TYvzKepkECAP2uMcLh1+P8pQ8HocFPR
HmPoRGWDbtCPaNWcgBoaC1flLTCxQ8Ms/LNG7l8s3jucVIDDyra6lD8lutGtMqQK
pKP83Z1J4mdLfsz8pKV9tw32e5D/CzgTrfspf4yGN4852xfQVs9MYi/CWhmcKPaP
oys9GTs+Xl0P2eSl8IO4b98y3sBsFwSoYZy/8ET5ENaqZE/vLgLjRLc2uKTTUkKV
8oAXu241yd6GyoorY+B8M2zwqNTgGHzCMEJyKLs2jZt62F7lpqyQibvMptGCxk60
FyhuBUBX7agjoB9y3O/z8qXUDK1mupXeAPdxyAPYINaD7N6lmH7j192WoA9brXz6
lOVePxMpjfUb8VizIYgps83v3v9eaqqyupWe6g5Jez3xDD/VFDZl+se0KhAtMUSU
g99k3LHECJlOF5l4sknKxV+MaJql1wnornkVN586+69i5F9p8h/JWfbkneg5FIWW
Tl3m5X73QCkWB3yKNCXeKRTZ5TiDl2FnHFMO9u1BOJsXi7xpXpKxZ/o0z/b+abA2
3uVq47EY2/J6i/xc+hsjV2TXepkUA4mRA6TEbAAowrrAaTBLFYy4sxpzAoJocBqg
A9EbB8cri/8olmhlU9r6TKTnK+6f5nQNlPVpn2JReQvo0wslrf0oCW834r22hBV2
krMEcL5Jp7LGi3HW7TW+EbOrPpBXwth1r3RC0Z8RAxIbk1ZP18e/hsFkiThAydo8
VmacTVSwf2ufKgmyyUZpLgobXp7LvA37IJ6PnQhFOwKASmE43llhPuScFiWx27eW
/6lyGs9EJE+0wuj72tMyUvcL27DOFTyFgklV4V+sDn9E46bPWOgWwB0uDGF10WZ4
NmbZsxF9JWTJkEevSZ17OUgU4NAsKUDjVImP2rttYW+om4R9/t1HqajwcCU90hbG
pJRxGMsvc+VwCvx6trB6KAs6/gi4NusqhTKOPOrgRcUS9fUb7h5FE9MOVUPVJdAB
ZuWC+kNxqHvUrlPcTdxlNxGLh23OobiW+J/0yWsJbDp2Vh/njloWC6Hb6RtB6A1x
Rin8j58h9kIam1iG503cUkuBVTb6NBFvHrRBI1r7YKp5aYmcTA1sfuS0+RtZd/dr
m5mnjWkfwN/tDyGV2hIKA+qBkuO4ecOkuI67aLWbqvDob2aJrie/0CTBjRJ1ClZa
Tt+EMtV130w5UEBVH59gREB0RZgWG7Y2blXka3HrqM6EogqFPANIlG9MVFmzSZKO
8Th0njrVnswE9B74Igg0zjSq4CWNC2MwWdcDK+PBcPSNn381tFep1m8H9f+5jF42
8qPk9ewd7JC0EMKvvtl5/Z8tPstLk44nHKWNRgqVzgLgYosk7cvK6J3kFVU4e8yx
Sp8lKewJvYZgDe4RNDDU4PBg6/YHKh4TgLnOjSqOflkzWUilaCpEQcYf1bvIS7Ww
JG4kP8TqZAFCrhiPHc+zv0YzrrbzjgrCKklBPDsnQqlOA5hqW87xn14wBmLxtAov
M4bJ//cR/W7KMPEyZtjHuKgHitMab/d31+YrOxCDCfKVQRfd+ylQ8kuxK+oSeUi9
Z55AmxVImLoS7HOpTm3OmLntW8Orq70Qvi9j5UNig9SdzOzQjLwYD3Q+OYhLovM5
VSF8W+0gKSjwe6WYQ0nnq27A3RIzeWt+vVLMZGP2Y/RtxXxrvXif+SeyrmQRD4Dd
ECrIwR4nxrQfyipeFWEMfM/C1qU8VZyTDDi62YRLjkAJXcO59uIfhXF6HaNeaOkJ
dToEtAQz+IMGw+NyBa6l50XTSPSk5yipsTlCkjV8YNI0XfUfrLiqmzGQbF6iD/Bn
EaIEJE86Wu08nBLY7tub1r6iKdniWjglLonIat0E9e+gjDumKRULJFKc/1J5cdN6
AFUJFlU886wK9Rnu147+yhb/mXG7GBasE7J2sUn6nKD/0/bTUMMq0owsNmiqDAqJ
pzpnjDJz7tuB3LTjTxkSgemGU6q47G/la35QL0wEZoL+YE5+cj3jeKNaOiFNTxAQ
9gP3LOt91Sbn8dGJm9gGqJHK+txQNdkSdA92tgTOyH6WLbz7dnS7blsW/rIqZbZk
D9MsqZs56mmTcFYHEqHBjaIXTRCzd1yX/pC9vGUmKNRpWyxM4ZCnlwNaVurGmeUI
y0IFGhuaN1SAEGCAuXdZbieclBbuGgPztDMVi1i7AyOeq6TuLYPVsxGDM/5zkKYK
kuPP5D0GXUerO3nzdnUYlaXhnf3YPsE2MueoMFfqLmkjbx4szPOZ5BY+JKob0rpQ
wTPVdpM9kXebEQpcU9qtMdPxtcRaXIHAzZj8yjn6vgQweCGO9HE3BnYClAuRadg3
ZeqedPEXk/gGDZfPyKgspjj4aLlcYiZtO5exKkzhAKQx84G74jNTS6WpdwFIFvwt
vALXpxp+o71IRgy1GIP9WjS2QU6m0X3C0RoS5uZiDH01eOtXSpo/Dd5ohkmuYtM0
eyv2P8RllDvmj24R7NhdGzc7KI7IlHr/+detGfxJUV+wCQ45aBqtFufyfdNSKoNw
S6KRpP7TtnvfYdnBeTBDff6H+idfQLQ6C/sUdJBlOrjmMW/o6dXjGxU8vGorDTv/
NrQkSZne5w+XjAajue8VLeOOtGxx9fHVkK06BAZ0jnZYO3/shQ0jaIB5Z2voqCeH
xpP9vwIkgMAhufo3VfAbVPLHc90BqZTX4p3ZZ/iypvCN2IWw5Z5N8X9kq/zUO9tt
1U+Csz6PsoFV1pPoxTJ/NnfT8hQ4Nj+wuY7yLsYbp7sNP1DaBWcfszOf0RGByppC
gbejJDGyM09BtJRT3Ph+wyqtrqT7mijEvqKtCBdw6FO5j0btt4m5hTzYgJXY6sEO
ptvf37MGuKF87n8eGfVlFLGHMnqKWkDvi5DyePzUJtyRqBD10+TDyw/LCW/yrcsv
T2V5DO5wWf4MuLy1EUsr7TG5Ln9X/kfRDYKmnMQk3v6yNtpeHVG7ac/N7Qd7Fos+
OveEGKgZwVHBG0VVar/ogOl8A4/JG/ZPeiR5v1uZhXym3GWw7C4Cb/qNdOhegpVA
fPhXmBtgHBb71BAA362kz8bjW1PBPATAv6juQ+wQiwGu/C1k7gdGzHsbRCdExEWO
gzEUrivPNjoZfLERrTtZY3mIiwiwMweSSDMyZPACPdLcXKQDM/baXVDI/+H3Vgfu
DgjI19CcQx4Y+rH9IBipeH2s0t8JieohUpnDC80OCPoonAV37hKA057dlYAjkfQE
XOcXFecmGcLO4OvGf0VyEPoHqjoamOxbiJizamC2KGuBO1wqqDapALi6jDya99Jr
6lOFUQLGvl33qYv3MEi1UOFfKq+aPkEbCqXJmUq3grFd6T8WDdjw3Xtz8SWguBSK
gn3fZSyv4bZMq6y/Hnd6kkLyFUE5FKo/92+9yzazMJ8e2HbiS5sse1FmU4XgTdgH
1t3cbips5V9hUxP566X21z9VnruuFeL9q/9IsUbexvQsUUcZRUwRs74Ia1H3Z+o/
mdsarCTJGeOrCCQl8dGNhm0/YNfpFK2AJOurVTq7wgI+AFACgtgXhk51HjituoL3
Eu2sYtICAxelo+6ewA0XwzZSH7WugrtabmNkLEKffKTTh3N1yqvl4jw+VEO26QWr
vFcA/R7NeeFCH3xn+KNNaBIdpa46r/M7fe02nP886bk4JvueZso4uwkyYZRHko9O
984SFE/W94zj+NNK99mgXzvj8zTOOxVWUfGH6YDP9sUsjmW7Aq0nBEqf16TuAlg0
E/tDTQIb+L9n3NZm7XBXTiRiAbukVHq1ap0Su0SDiVIhXlkDEnbMM3s2c/5oGTJH
B7IVxPSPgRpcCsv75Ro18stIS8SMsFBwKa8/Zor88jL0yyMcBRCn/tHPMN3Q9rGi
8yxsJ2ZVAnYSAj77oNIkhAI9BiBxfodvApWzaspmpi1OCkOOqUh40H4woSGoToTX
l6og9HI9dGyvCaNQOlgDDihMQfofloWz8Sa8izgj1HmGlIT5dFq0HU4MEpT+q/47
ltYM12N1qihPjjz2Aty/OpN6qRDM+ILIlsTekRrSam1TPe3anzEZX/mvSWPcs8uw
NQiN/rZ5K6qaAkTY6X0O3scT/T4OjQV1w5cZGkgLWYXxd3hpYAkSs05cD+Z9c/ia
nbZwcYvKKEe6SsdQNBwBNjVUWqofN0jsz7rLAM0bzBejokMoReQnDmPkL07JVjFr
SSh17Cq+WDzZ61hj0NQ005sNTdcnv0SDqECx8FvV4KzM6p6E6YhZQZwM00twQcfn
kgETfgktM/Z9HVu5tP38A6iAqSz287QhnDhw4qL6mQ2Ycu/k+cZb5xqpy5uBnCWg
Jn0m/RjucElrQSoeRQ3ZFsdUoda6VT5ykvWRwrmmX+NNlOdx5L2NWSRRh2AzJ0LK
h5mc5bH7xOS0y2jidNvW9stkbFcg4K7GC1s2phKLn0HgXRWKJeGeOZSNHqUZLuFJ
OwI2rc3u4Uito8Gd/jwpSmH6epQkOTjEyf/uja+uXtvuglZEJZ6SeqwuA2wp0tRk
RsHRN7w9n9ccg/nM/CjBpfDMZxPi5iM/lij80dwirvJnS9CHRPCpqz0cmQeCMaBZ
3UGq8KVP2LcsEDipzCp+DjMeQ0rreU6hfqZtKnru3n7G4prrSyfVVe7ztytMGGr8
3nwPPu5PISibQq2aR3xRwRWlIvXRPUZQVYnDh0ro1MrxbEX2o2Y0zD1lB+y95/7V
C0pjCW5S1u+iPh49wIqLahg37itoEtQj0LI4geV8yJa83SJQqLbtPu5EQ/fqBEi/
n84p3lh353jn4O479mL7kPuwRw1ZGa7kwrM46AERjoswzaw0Txjs+CFgswfpF38Z
ISZmfHBAoAWd81YlTaupVHE/OXjDZylGqHuwU56LUsKVDA4j1PMDYmFrS2xLNK1U
6CDtbLKT6XQYFS4xkOaLwck9lKjUcVobIELYxVjVpuHHTMi8U7nyjhKeqLhYYXAr
gwFuardEOCk91PmilVXzHJOLkyyokWFrhxZ6KsfFsMNcwzdYhFV6qxk2LdDr6QAh
za3cRqVM+zus/ss4X2lzVFvaQk5k0UeJrkmwW6uZL0e8A8VDjAL9zrJV4jw1CzkA
YO5dKjAALmmUzLB2hygB1FLGD16tkFjZyNA+tbhFYF034C5KtPqwYwMgcEmCEkq9
CDRZTKH/0dnLzcapSa9FkuT1R0joj9HAAQG88gc9EDa8zkpsEg3jvYxzsazvkhWt
34a0RX5pKW6rJEf7vlckY8vUcIalBtfD+mYFQ0IsLLOM/Hla6rgcgBXzouDqbfsm
Y6KqQUW8xPO8slE8eXzcW/ZaUHW1E9GmrkRD1vYJD1lrbDt6k0Fv7cRi9B5eW0FU
ncJk0FD2OGnEiAukKJE+3SJ30+SRBcPY74KEat0cw1ehIl073/WRtLXZQABcRM9L
8FajLna6KXnN3Bm6KGhYwWvTFPix048QpQ4ehGIy8/RzjeqynRXVMOvqNfGYRG/D
KLu9SxjP9RIBwNN3WtmgrBu1X3rayli3HCDJy5VAmw+AP6KUcNoLrjlGqxvHclJW
A/fFsbgGfYdoWBKMdVGgJW2DcHyVflagq7cRL313YXmtmfuw715kKuHmjcSxGdiZ
7T9WVrcRrvpbzrxuh+KkGTiD8wx+DxC7SkxnmJroQVq7kOXWUHoU91hdlp+thoNh
Abq27nkaprVAhVGIIZ7q9dBlba/pasUKNDfkz/jH2FwRFtEDvTXZo9hWVtwVdRoo
Ni/1/q8mqaqZjp7NmHESXwg8l/NSklm3N0M196A4UaN0ukVbgO2WiFQyX1JCzS5f
B2krSG7Ex1MET/Z8D1tm70LUTWiS9+tjHix5bvemZZZHkEx3umagcl1GG+KuuHkL
8IFaExA7iSfWB+kGcE+ROa+rdeykEJvMVWqhMV70El+ku/+jGLzDLR8IYoGVDzqi
FkYx0QlSRgQW0GUF6hZNyuqfLfU4Sr1z5LWY/M4N6xDnTGTrVyXkt5aZH9yin+j6
XVOw6E+KnxbVwoPl1ttbFNF0DU5JPbN1uLAUb6Nxe9KXEIeqN6GX59NEqxqi2mzh
4nzmAtpwuTsw7RBd9hEf6k9odQqPfrjl3Ane6Sq502hE9A418zDJnjSbSEEjsb/u
iOvMfN658g8RF5EZUnmc7gOhFyclsoNqU2HcscYuIhHGg1iJ0lSzIc14+ElqBon3
ytjcavnbsZjfAXyhZvTd0seq9jANECbETtKsmrWcNXo4XLk1W2CBN3lPdtXeJ4fo
bCI+jqnFX5cA5/GmF6s/sfQlqQ63hWlEIYgJvPloWIYY94c4a/FTCRolJZG1k7IJ
LLf0/3DX5rsQyhEt4q+ST6R6xCnb2gIrNHZJm2aAdXgsgZJWfCyE9kRzv9u2J1di
L0CUvJHqCiPsF0BnwJ2HIVLSR53CKhq8a+jW4CMqIFU30Yo0ENKSN032d0UChD2J
71fYrLgz27JfB4WDHDg52jb/7I6bbJbuGg4Lc1pItH3BY1yPP0K/WgFdFNUqghai
Vuk2dHP/yViN57nsSJov6M9sqcinwhg4F44/77dHPQpWGy9SeOfSxqRLABCZqOhU
G5UNA6FrwB6dlY8gylC4p4wazysvcs1e0yqSvdctNAnpS8qmuAalN5g0LE4JmXbu
L21XLG0xFfsMechjyZuemW8fWsJsGI1zGofDbUdH0vvo09yCTRt7v3poRZNoNJYU
IU1dS9l/6mHxT5jcitQETGulpIiHGeHW3szHPo+GPq0Zme4L+7CAj2WPlpCfh9IH
tHRxUp+seDP8CQ7w2dxDADzny0d9xGOfwf84muM2J+WO8ldUQDlmFfTQiNTOWp6H
dZDv/e8nHscWPta+YA0qM1Cex0gX7JRj+dbBw2rQgTdhtUQaVVabN6V761xjTP3o
dcMC4rupxUZWe5s873yvH3Dx2OqK9ImrmMNg886s3JyUuOwWFRLZg9EolLRO+9pc
yi6E0/YdHoiMUdw3WrN9weZxGMBJgWcf204wFKvOahSe0VuaMpl/1rBa00vr7qh3
YJWwsg5I7u/eIdySPIsFJgHfduWsVm0CDAxsfOXIYNkVnajrQO0ji/YsoAl8cd9G
m7tD9RZgVa8aj9JbxwcQkiC1HgVp6pm8PvyXezyyGzvXcsXKQUGsbr9zJcrlpgeK
5kGrLM5keD9S68nUp/S7Q2Kfq1Py8ByT3XVOXu/gvVdhKmzhkox+lxMNrh0NrQSu
01ZSOMRa4dU32eRsbZGTOZ+m2yc3E9zngvH6qbxyu7eTe2cxmqy6LQEljvNT3V04
EEeCX6l4BtrP3dxfxQ+aOqooRGCpiRvr31QshZzxb9NPmZS1El0k4YugyFippIuf
O7yH/peA9AtPVMRSUEeSOJi5X2/4MBEL3pZefH19cKusX4KRrALo/TKqRZ6ulO+B
ieNb0EoX5xZBijNqEWmE03kTOV97sCEZ82OZi796gOciA9NAqYLAG5UgxCt+oHGk
Q1T87AonQMdFj1BfABSawjVgaKBlHL6msRnsN6rhdy1JomA6zH7p31OrTk3EENDt
2wMV+6xGikVBvKr+phMLFENfeRbtOGt5k4fPoyGAlD7AyE+TNJf4arz5gipSBob4
mDEYUfyWP7bFkXMn1Cv2jtnGrL/gWygWlf8LjQMgj3RVBgki0eDSaCj41zIHNbYW
8IsFV6LV0TRV0yDutqg7PtFznied6PvI+foP73jJzJFS3+/pQ2JPKg+IpxefCWPx
MFNtaB1m/U9krF1BQw7LVn+OrRKXRlLxF9C3i7RrX83K5PY9oLK+XspUyKqbZj3b
V2MOTWHksNteEUbp2DMoMqW+SxChFnDlCvdzpgOwyLqVnblfuh1VOzFxkX1mRjOz
GJOut+VZl1d6KrbqFZ+hroF4dhlRohJeeJoTVjPPNYqeKI2QWcYwhjRo+VCZuBbT
IUMrRme1u9cnEGJnF6z6F4eKLvrTlgIXaYcwpkRYgitNT32TaP+l0EOGTqUKmJCt
X8qZDQrTJpks0aHOPneWh0RdvxR+lBVS3LiiiFppO6sZj8glp6vnsr7JLBETM883
AbrNOh9m59YrXeM7s8/yIyAQ0jBuBA24LnyplYTfWaDngYrmoQLpC+71XPrLxK/F
8Yik3Hmdh7F0wSNknaw68L4eE3YuLg2W9mfs08PhFuj4Sd/upElljP+Vu86Kqq7E
wNtl5My9niZ0hukLt9RLUD2mCcTsGDC6o8Dhg+KEd5qhIxsQ79Jdb9m2dQEVvx9m
xLCG5z3SPQDa7av7+0S1hczW83N3JPX7ASt/ygxraHr6taJkbfhihVJQa2y/ZI1y
zvMIZCd2imfKr98ykWwIFuqz9ImRzXLPs0yVDVomW9QTJaL6jB2dWNKhvtL+xA7j
VekqHVSlXA3Qj4vv+YobfjjmIqdlI3fiLjrLBiNVw8MjdZ8Z/53oqgKQSbPoPs5I
dRdyc0z3RVHUUzPBRzh/9gLtT9VKn6vyYLtziHhY1siSwwhgzAzN4F+wevDgygBB
F3vJ6C2CcPsR8KSgjOJiSiF93XT7ny8z+usqXWLmODwo9ktaG9+u4judhmcGeROh
lGsIiHqIW2T1g5D2Gb7BPSH2g5h672xm/0pyXpqlDF2585VNO9+ZDZDhVnONvYUx
JF4Nkv1vVBxnKMTiUobs5Jol1lQTWc6oHno1rJ2xTQ3l4vZbTBO60q+TxxABA5FT
Xs0gUp7h6LRMps69+/9eGTCK71re/yV4esVnptmauPM+QmTwb2Y2se4C+MPw53z7
SwNA1defZ8FfpnLlGj4TAgX32BkG9A1frmzqAxLtjdyDHIaBIA4iuyT6Oya+CYma
ylKIcvODVOpW9MoNdAMF1eC7Y1c9QdsWlbOhfXfPH5aZlh15sR6WVyXjG+8MyKLS
OFJfNFcbtFBgaJdZUI8CGzrosr/FU4XYlaSdA0VMFaudqMAXk6O5cuRWp1On8qFk
VIVlbeXMbiLZFpsSJol5sjWK7W76SZseOlHV8FPln8blvok0ldm5ZyI/hEcqBYnw
V2Zoz+D4mub+35VaF/QpvAEAgEDt5jKwDyLkMw/xxw810nqpWZUGkftpx2IO6gNN
K589p3Gl6X0K1qzaFRoo48JfbouqqpPJcPouJw4KsSmIOoUbP7FU56sBBTifeXju
pN4QGVjFmoqDiuLAfmcilquc1cPYP/aze87k9RHDF1AHK3LRudTDUDrG147qfo1W
h99kof5OfG9z7m5i0EGE+RdHpTr+aNAh2XF/fnCehACKsKmqhHdmEOpRr+Ymv/Iv
lL088QKl1E6oW5zzw+FMomFrcnHsk3rE0ZA4AfPJLNvhvAPqecdTutlKnpiXYe/K
h93lrUR9FcwP22PWLW7vghZDmO0/SeU4AU/iNuWLhI6SYNvy7RIkjG/6bqyswz2o
2xfSqLJayRAjnuVav+50ly1yI4sBYrq68ffP1/+SjpTL5QBe75lVpUwVYSavgVJo
25T9ult+ZqSB25kPPWznoW5Eav5WYhrK+oQbUmX766zdtufUrdtBk3d/V53rVJFm
6V49AoCbRXplHdMkX4CtRSCMTxQHoc+lSz5EAf0qehy1edKZnBzbZeppnkfVAUDW
3MOZwrNjyp0Q9O0Ghw58rm30+7IzCNjcWJEbHa8k2NYTWpYgoivPI2RGLSaBEg7y
nA9KxX9ANDkLulaHOZ3cb6CZbzY4v59vNIzIha6asjmB7KujAvJVNXda8Fi1B1g0
zu2+huVeixiV9cD4FokB6ZwYr+y+RLoTcxERUkM4p4RiZmCf64AU9Y1FHMTbV9o2
g/vSqVu9zJpRyt/gTMNM0KF1p5wvsiyzfByQuxWagUcE6ZsU0pabZxVqur2jZ0jx
2uLh2Emo7bvSS611yj/Vr0t6a3goSxGR2ffQmVj4NppZ7H9/fYbaEPmRQwC8iiiY
1FJ+tT3n3CefL+stme7vX23LcWxOxXV5xthFn1YbER3gdqKithKeLGV/mWN3K+J4
5MopQ/bv7oQT/mDIBo+T4h7j8EceXixvH38fUOv1rQaRqTZabyY2zhOlxocaF2XF
0xiR4Xu2m4JxOa8xqsI2tsYaWOPuGNp9ECo4tZfvARfgwzzk4Lv09/vyhZoXATl8
B7S4GTswjv1/aBCJLgPGzQv2Py+nNP/UPJC441HXKgD65lI6cmA+ObVL0HJzkj0x
zRPE88VDYoLK6iLi6c3yUQUXEy0rCltz5hf3tF4mJxA8qSNxRi4J1p05JRPwlJyy
amEKC5uHat/hVd8PKsYcZhkirWMMYMiRDB76PcS0FKx3ifP7U6CfaQE5ER97raCf
Ti/IHdI64t1T53K927AXI2MJs+/ZKkML15SoNjBwAjH01/1D96tK3RtRRNVoru2l
A78Pm+lBHqfjA27D4UDJfaBuDS4MlOOAzdQZPNnYJrjIMP5WOYztOLgwhWJho2hv
JCaMA12YzRFB5b9Q4hcdhrPy9rX4x/BGVYiEyX3tKpk0NYk4OlG3SfWSMQrUOEBA
CfZPkS6WaDxesNy/q+82+VyWJIdWX+vY/eVFhUGsEEykOT4okCp8W9mrg3xykQEg
QNvRzQUFc1n/RK/Y1KTJPgvwTDMQSGlgc1XrCCqX+b6oAWGiszkln38ZvCg5YBBO
bgwj8Hf3Tq9jA7xy56WaOz2jyun8Ck/OByDaUacK56mOSwLt7GY1LOMHY8OUHTQa
E3+pESaBOvbOm2uXha+53o8jD75AdfXiy0Z2igcAmMeB0JUymVREQOcQ+YINb0VT
AxLvednmh7kmfPckwkw/BxD8UQAM2s1N3el4j6VykxL+lVfONI0i9jbrhmp5jRbS
7Wm6ucCXckgrZ/3f7CfcVi/Wk+lOPfbLlfStnosFRCo+p+LbKKc1tcKiyjpg2ZSE
8eeCLo23dlKBCwqmtnEDMMl8dC6mrVxS5t6dgLjCyiCa3M6p3O9jCqv11HPCrTjy
KNLj0zeInLxf/9rOxu0L35o63kuJgNYK4bQzEFKqeGLDwCAKqzUUwrVjUD0cCiai
X6M3PwUeY694A9+7ZVx8Q+7OjNAqHdivE3JeS8/Atx23zmPFQ+WKDczT/XlVxK8A
O0zjVSBS4GpcQggCiZmUN4PN5mfBF9Y+FSJG+XItFTgzFUlHZIObmjF+IFsYi32d
CLGLXVT1hEN5G4dz3tkJ1K3VDaGJrJRRY8DRH/iJ7pPdoZSeU0ibh0ue2+U5Ymrn
Ta2h6IC4SZfG9JlAoir8FbAN3M1O2R8woxT1/TsCQyycUHF1NOSWXGSyji4upTI3
FFewHd8U2PB5IRg8NHlkM5zRUX7CniUijJ6OGsheoYCuHb2iHgHnw6F9HXiZzTWN
OrjMdVv76Jl0uODvVDC/ZRFTbGIh2MqiN6H/Fg75zCohaui4pNq9DrDdvmkYsATw
D4rAeirkLvYfzcXN2GWwQqNLsR+5mU5m+ov+efMaDzBvg3EoKfOhc92ueWb4emq7
av0upQEDqdhqcFPB+Bth2H+tjM1Wi34ME/lmUEVKHZESpRuXlS57J0KlUTerhSY8
DLVdfTx1lXyQINw7QmpetU2vLn9AOt4GRxpewNXjszIdPQFp8WgRRMCxqJun7kT6
VjoxMbFQBhdjFQOSXnteZ7NozqOHU35e1QhHKA0NXSZ4yxnubix2pQKpDbkRUegz
+0Jg4BpLUyg2vXvOt790IaMYuHfCVq8g/s5hRpQt8WPbGEWiwjuWAS8REZEhfxZf
+yEAkbXeGfPryTx3X2qzh86YcJQ6PeCajs0iOItJ7Bc7hyV4GP6sZaCt4lW8UNkD
bU5PML+JQkQvLK1WN6krXuFf+iSxq2rsW/bPKdtIjo2eW6ZTW/uwxRolYi37c7q9
VK0x1xbMieTLtznpMBIL3EwLYiR1v4Ag6urNbA+T7h87MKVUHm6xZJZtnyf7HJNr
2+OREKDfDWHoxzYaAjfGOD14+1FWG5lsOLuLykG/Th1tNhYwmd/ums4XkVjRhboI
XFpAenQbV6UxtyBgEi3UxqBA+9vN3XtvXomn6uG4AJ5P10xa+j9eFhlLSYFc4XcU
Uh3rTH9AR5I/gZPi81c9jwuE2gzzNbNl+iUMyCqw8Qi8firqzAfdzA9MG/qnAUrV
0hCR6rIcZnlZf7qnS7uJ21PRdjYYbDWetgaYYGy9VNleRbmIzSMAaejDXrceoPpu
nFq9c2QLCZQV9ZkCgcMtejpfcXL2f74w4GW7BXqci0CvorRkU1F6W2wUDk1wxsSM
JSyNgg5C1/R2y6m3mIWyid7hFdDWoFZsADnNaZ0S4iSB6eLa4nglUVEjm2rPTZLe
yZZ4tALdJ6Qw7E/B2h/yCjkvLWPPtncy3rIJgYyT3zGi3LkwqpwIbJFJqeQsDNEq
14ns6eNoIOSIfzN9J4duXtArcyBXwNCM2SiTcjKGOdrslMwztd6fjE66E1puIQCI
RNw6wxdeJN9857IfwMq9Qodx5yE4m7MnJbzxglGeFWwRrhxVcvSL57GhqqaLQDth
wtHm4rc8PVq38MPWAho3+yVwNbUW0AilcJNOxfBJKhcWY9+zSPDxKkLYoYZHdlfx
V4pKbaZ6u28cpdpeNwNOw7599uM/l69BvwWIyqOZyfoa5loa2X6H4gP5ydh4f9gi
6PG/cllMsGFcNLV7RMH2cDzYs0vxJjM8tcvXzhQXF/OcBDk7+7bQ8FaAiQQYcHwx
vP6QG+Qz60jG3FXlCZ5AknS0SgtNsHzTmYvlZbyO3OMjSsNSp/8gqaZpsBC5oMQs
FNF3VwSYtInYEmarcVdILsoKWzI9DRXfQi0G8RuQK22Ar4XKgf9vlzOvlJAYI/nP
9TD0bdmDpatPEGT2PFsxYeL831+SLmkNI+wXDSrKUyT6XGLryc/oFjX0kR7b7/Uk
YRzb6dXD+Q5F3ZMK1wkuQ7IrlMkkTnMAUljF3qh4gsysTiPCkH9i4bQAiJzZJckO
voeaTPEfwHMi4MZj4PVAonpOBaQ06t/27XwA4dBrTEPsZdMz4MFpzOOdQF5+jOv6
7oR564m2r+CXWNrBULd9HACTU6EXz769dJGYhv7pqqU+bHEY66ixm9+TgEPkBAMv
n+E3UJ7jXQYnX2/0ncTMafFswVEFzIkzDFGkN4LCoHUTwk8YX8SP5mV0W/W4oYkx
//3T1to7ICsy9APU8cLcuHGWCzjWCO06+WWV6QOsQWFuNpIryEHBpNR81JDgU3lr
G4NKQ8fcjtxnhBKMVHcVW8xVXvHlgEn22DozBouB1loiXiruBd8TZlKAqkZl6kVb
huxhwOf2S4ulla5pQ283+zUUYJlIMglii3azfEQ2l72QpM/DaslaYO+cO3n3mZDW
I0xS3o4jz2i6bXUAMl6qeeaR8KT7+TuejB8WcR60cVgLqxLiyis+cwn91UDlNts6
kkCS93Ou0lokEzhZV0uQw44IIIvCAvm3lHMgMQWg0NdlM5/m94PYVI5IngdWEs1y
C4KHfmI1eC4xtsjEj/8r6SdSXm0CMegIU+5jUvyc+9aW6utZwdm+M3p31J+SAR+5
v/zhh34XkmgLJoXmUS9s83QViuT5qFvHFMh+xTVlUsgP4CLBFXAo65SrbxW1hK1V
Jl/QrFaXapImI5z6PgYCcSNfCrBvpE1sn+wI0hlED9izAV+Xi8i+BLezEhKLG7dh
/+x0cCqpy1WidZY+xnn2KfE/58VF0cQQomXh3XCPDXxDtXlxt7tW+oDvoUTafzQQ
K/ijl/1P6ms+uBSxXaBqcBsn4l2fyS6Lf9eBFxJQUvgVwedjQU6HyOZh1n6h+sKP
vstv7Muhhq+Kc1Dtyqgxwhv6OpyQBK4+/ASMlS0KXF9czbN0arKT8HhAvmckw58X
6NJ6t31Visgou74rMmePpoHjd6InKLhjjP7qGvCm+VRaWz45f14C2J/3tB1vDD7J
iA/WQSWbSkPg1Yt2s9PYrrrMTTxiHGzzqzaCaWfAhhq+y3hFiTWet6i5L+JNAm+2
0xFwY2/uGzL7xhzmL8SnD+hKadgHs9noCMNhmertl38HWKIKLaD9qa9Ps3nrGU25
OfMZwpLLXrZNlfsnlljWLwet3oGxlMINo5CQ2m3U3ZB3m9TRsAQ+nGwzzGy8H802
BcBmkkyzhdw2XelNGU8KQgFYBmSI+0rVFskFtmq64Y+H4pmAteceMKjY3oa9T+Cr
w499MS9BpZTGclokDVhvafPCHko6vlQKVqguMW71ezIuuVVSHqpzbSV9QYzkyg0v
XVKUKRaUhOF2ewH/ipEfcvcphy+52Efd73ovA6d0vA3h9KQnCtkjJ2p6m8blHBtf
hBDFoeqKqEEjjrkM9r9hOH5ZRq0bpiUqOumHdbaetvcfcJNMywGz+G26T+C+UDop
lAw/v6LsACrZ/leuVp9fE0aIKCeqm5VAJN8UmDpimasajnHh4Tx2sJvn7HjfaN7i
JA2XCzgG7Iq9Nbthz3usCZxS3Klz3KBsClg7Cx7274GlTLO6SJ4SlQ4YxwyS3+u+
HUJ3b7aquR+CLKcURJUu9LlywnxRkYuEhYczllA+FUy6UE7HHAI2ywDAGVBwaPlK
eP8WxM5My074rPceSIMfWF+sXFyo2mxZ9VUitPh+4MvZWR6Jku/zwnxCbR79b7KP
Ol9H3plw1j3Wt8CTwEahdrCKTpxQykr+xU1SomcxNDtrWD4Aem+nbIdvXQ+FwETG
NSOqswycpK6g/OmOi7KGLsx0iYDPPbokyFTpdXx01c7XFE4oZzqD9OfVCDRzgXQb
iYu6fm+oFd8cGwheXQuvgiYsRDqvfHWHUmf/6z87m9NapJvXXXmDhf0IUAdTEmcw
snz9tvlKSoy4XIXeKzn2hnRFbHlKCUjYF7UBiQleChW31fHjTJQE1KHZuIlYAzuU
9oq2KPGF5MdtQR98AyNfRXx7WI/JE4+aMWne871l85qTV+UsZsPUaZDwLX7NK/v5
mhh1/0kv44qOj1pgM6qlAKSZegii9WVi0CtIYqBVq4vEZo/X6igbHvYCLNJVbbil
S43J247UfoN0ocPM95rKeWEz0j3lvILgS5sEuqGM/CBv2176a1EmK2R0ypu+ZCtA
uzbfRGbx+yDkysbumiwVMEJoFJf/FzATTe87ftKYS/aCyu0NBQhhQAp/pXLVUxPT
2EQADN/GDk8gwkrFmxcUYowcYOX8yQpJXWkSWAd3JasaVoa8l5EcZ9ryGOA7/4FJ
nkhv79BnPnjLivz5DQP6RaCLacqQbewEakxhExGiQ9R20tvligj0bquWn7HP4Bok
10wHSSxZ3/eybi1RU9OyGpfPT2CeXx0+ERIFT/fdBurhnwoO1X6gxGKzhIYWpAyS
wcEc4E6AkQndffoWL/C+exEYZn6MyZ6CtdLDbeVk6rvTA95N5QMtTJGN3nQoFCii
uLA0pQaRz9V5RFhYWsl9qrhmf/pS3qnveu34V32h8y9hv/CSX/gtRZmmi7d116tb
Tu5wOW8FGetZtzeLk/E2QhF0OEc21vaBEO2M/5PVU/V4qI84w5uUHuSbzQw5ri+g
lXGpD2yzCCMOql11DgY+K7/ot61OsjP9Ae8FMtUD6olqxVHNlwAWLCqX4uLPyF1G
NuyLB3Mf4IYiSCLJrlM5yV3d0xbKZeYZQA4aeHW/agW35fhuBCBuUQI6vu2NWjcw
ATElRjL8l9Q4xjQIYMO8MTejQbQxNLutONG+cfD1H5O0CnoliRvdWSI4jadkqbdS
LNP7aG3aXIpkqPSYVZFMF/szY5k0q0IcTXSKgNxqo1dsSOTSMgUQ5DTogNFM8OSP
n8JQ7EERbe7g2FYntOucoOh7AZ5WzELvGl2EypTLl/sLs/7Yf1LqO6Q0/8Ronnme
xbVIDPKQQvvCeIKMPgC5UyobNEamcJPJNb1hi04jMtUJwoZP1ZwNjNmfpQ3R10wx
0r4DnPtVTth5LG41x0vCKdtEqjti9WowGVy3yeHkuwcEQE0eZNeNzqsMXSkcqwe0
Dd4zvjrz5DMeaOV0/jfPmTkwr8ftrID9iOkwnn7UAGClA9MZ2ELpDJ8gt8XQKWWN
hTi3Yl10enGf6yF/nHW2De1/AVH+K9cleCwZX6SA9kKzKlViS1JKHCQDpvw0dBeh
bf3h2eNUXAs38PBmMnOBE8WS8itXpk9WK8pNx3/1724LUGdLF4ol2DwFpKA79YU0
fOrql12QGDMqnuR6K7Z9rwTsn7PH5eFdPFK5FcODH4bM+lBmT/fSRXPM+idWm1uh
9HS1kh6KYOS6zxeO3itQdpAPCe50o/H2ao8AaPVjqp2TxjEDFJLxvkKR86oFDDiO
z7vn5x8HIZMidfpQywhVPkIJtbBZ5E19kicsKuQRCB283/o8Hsy7A4sw3Z80li3A
jFH7rbxaLekQ6Nab6nrTNK+ze9Umq1LCSgQ8XOwO56QDoAUQz9fIZsS8SQPFtabR
MY/gtoX+m9Cn8KnTOmjU9bZ1+F8StjGHD9wy0MeiASKAc5hL18/KAx4xw9Uvt1TA
jbK1Yi/U8Pji85/QoFAYZVXFuSyHcbR3qhlJWAXhLSTZftda46ARgnP4YQLrX5lp
TbkY8IxORpLYTkTjEd1qC+RhNfuEq4RNwAU3qVmIN+hi2pqXdH1GvDqv3aLhMplz
+Ac6Rhshw9cSITCxkcaWxKkFm83abJhZrTUcCH4rPMOGLuvz0XK/yL7OVnfLZbX5
yHci3hO90KrdC0OVYV59x5v6DiAJXd5gMQRjqSlqT/dQI57vbwzw8tlJ9oktslgS
EF1ONoxtHotyJfqMNqbyBKhlU3bJ5VnlLHZkdWB+gpIzD/RnIIlhQ5k4HtFhKyqQ
sYgxyztngbhGjsS/tTqvEwlqMg+4LJ4VqjiU//iGm3Un0SVs4AvzPRBkuJJsNgF9
v2DLyZQ4pMY1YXgSPG+EYiXCUmEnI7ZdwspG2VU7BDVwp5ntBFUnCLmlHoClAfZ4
Sm8shbb9GFViB1XdkLYLaGooaPSkJxwSZy5go6u155IVGOi9j9MDGLnA7QUW5RJK
3L65cZDLMqhS0xFHyo3ogdsSYi8wpgsyBMiHPSyD30MvT2wMjc4uzdYfFHSakMin
ftDvcd027vNIAPiJo2eJ6QldTS0o3DychUAJQ+iFeMx1eWltNz0KELFz1pd/iHfq
SrFRDe9p1MujdY+gm3yFNxRY1fYzqT/03gfzsh4Dp+EUthsEUuXMmAqmtd3py9rj
IP1i1P02/r8C8mLiIFvpluJf7vOYGKMVH7F54zU3LjhNz9lItaAxD18bCeR5dIX8
8lkjA5Fo7E6/mUFil+BCTnGsEZx7+es73+wiBSt6rnQsy5zm2ZAd2vARlQZcaSNv
SjdB7mwPnJjBETIT6kys13SZSJbmsdmucrtQDf67jQR0/jSjAeHNYe4Bt++PEZYT
IO8HiyJMGSoodE2kHDuU9VmjekfXcGt/gf43rsMz8KFjJ8YIYTiN9SBn32e89ifs
ceo2mONFCPJBqW90XxSXsDZgQgATVJbp38PmeXmiaUSgGPPtXripiBQeJKyGHLUI
R1oL47UsG3+l7VsaIEOYgn8RO5Tc0NWLeJFv6wWfAhsXIluaMSkHQ9zSbLAMZWXW
JdmyRPyhc92xH64UeXU2aBUojGDvyMIGH0Is4Dt++3ghpfPSdRUH6wOtffvf2FwE
v6zEvo/T+raqqcxIq5ZJvZ5KiK5KDYncTyLiYamqzVmkSbHEqxTD/a9Y1OQjY5vT
TvO964xRW68wMImi3HnpKjpsah4FUIcL7K6bX1/gGypPY8wthOJ8J870lNaL/fQg
9qYXjYDJHNiGAcrGhuXY4qU5w+seWKwCoCiEzAHTl6Xsr4OhoSW05goDZuU5mAyZ
O8M6FQv0wrtV5gNHcOO00Tb7PQ1UVJENhqmC5wldhpQ4j6XizJkX8OWhDIDf/ZAy
9AeAK5BA2S7mb8/tLp6oKNhYTSbCqH+vMSOwGrAGIq44kMOgivE40s/fCjUSw2Kw
1DXMDUkQbqdZfSbpT0vlD6r+2bEfzzN19obLFOZ9Yr2go/eUimSXhEQen74U0ZEj
DTneOOPU9KYmEoosLe13yv2rPzjh3tJuciJcwqdCKZSDJRjm40oJCnu7RhTP/6st
BjhZCCIis475/3BZ9ZhYy6oz8Hm/lZWriX5cYUiLKK/arK5/sSKfOMHchZKURusg
f5Hfh+gAKpBUleizPzMEItgZ6En2M0ZYsdIAklCg5qkFfhbolP/Lk9xP3X/wbUB+
ENew7qXlJoYPnPafbCxRdXVEjx+q1g7CF7pP4T/HeLEgPMKg8CgTVA6LI8rGoeIB
DIXRKg/1TQrS+I5iPosbCGZN1zf5pfDVqOEF/0CQ28SKQlwl9YmDHZtc38Ua6O4d
wTgMTuyH0/JZ9QLc6BLBbpuXDkLfa/rGEEOjOo1SPmc0Xcb0Pq5pubLfrohVemVr
LvlvJ35qaLn2B0kcBLDUgPsthBSU+NvM7esfMnkneAa1CZg7q7qmbvQue5VIqE1X
QRrL0QplhokPiMGSdqArOavOLphzYC6TgW4p0dxoEHhjmLEl5xPsqZzMy7/UjuIV
CLklgD7hMe0xRK3Py7d8r8YbrHPfbdbreGEvyETSR9IS/M1dfNpnUvB2pQFhsYM7
B1uJW7sS6gja86CUsDmgj3es5y3pKMkysJqxhZ+Bz/0arPWxCrW2YmWpzLIorYdi
0X4NAqy38ESQrFhZ+itH6y6KPGVzZA4r/IHcXnOi6A6Hqn8NesP0AHW5X65iYRAv
RQ+xOOxuGwlXH2tH9L0zSkgWKikCjbUMlE50PBx6gGy5SJow0jZZq9+pmQZX6MSd
WOvsF/Wxi09RO950K40136aZNJYATJKVsdktX7ZVi/pMoLhJU9gEg2g981/cmXZ0
kIV7EOtiCWgogRbv9EYJu0Ssna/9OiGGvU3NT6PYBK86m+QykVXtZ3WFmeuQQFd0
TQMEOeKrrqcJANSMusAfhoJx+x5qN7OZQzpgTuFLtebMSHqInV0O5n5N/9lExrgc
lAF9g6YpwBx2o4KJZbBq6kySmRLkJAAw1xoS3/Rem9TiCJcAeQO0shfn6rhpcfWD
Mu+6sb9qfvUOSCqm2pyx8xpmX8eYtpZL5sMttBE4WAY6QkywPKut6TFPmEB0pTaV
6LLmzkqfG+Wd4rjxqZEWGtFmhE+Ci7TPfiISSsy3gdwR1QMMlRldjBzHeEVAumke
iH1QgfuO6TeKXNF3Io8AdqskxXfxKXeznXfHX5uaViuYRdx7XyCYI23WNq6NvPFA
B0eg8khgEkUSFqHXtnkuDwmh6Fo8tp6UEbTp1xMp9NpsxdcOH0V/5Fctgk57jPQf
EjKqxB/wEoTe1DYTrpynaNttpEv3En/VDwt/mgcepzjQ5NJh+z9189XNR8LSWt70
pSB/qpVPGRteQO68tHyn/+6D2LEHSS2Qk+pU4zSRLQOsxRaZXeloSZ5xl8YZy+Jz
XImFZw3xUtf59OYan8/f61s4DRD4W86eD9zqwvUK1lv2lfdXPF3omXq/O9ypAQEr
P9uLqNB6MXAt3vVHnbbdc5rGmPMuo4Sal33z/tPJsdG9hYRcD9vlm/w79DMjFSTg
vMk3asi7aKUkgzxYf7FdWCKjIYC9l2dGCMtUJUtEWITKQmZxSakQzPe0LDE3TG9L
jcoqfOd3yoNgOeytbt/rDBJATocAwwZXb+SFrzIK4frXSSRSP+HcVVDeW0nBx5q6
Gf1vuwwOMeptj0GnbuDa2Cgk/yaR2EpG6yLyVzjBfHdd+EBKWgeBJ3NFcsW5W5vt
h0ni9zTS8uO5hQDQOiqJFYitHPyNuxKQgCquxV4qvcNwQtKKxADpXrI36oOuBAt0
GxxhHKj24FabtD2pfSjGRvY862ppIvsiSO2bKNTXOxUK3/eQnX0xnlS6R5H6NrHF
4f3ppoctbYltUOG0A6zmn3FJqNieb+rEbDg44henVdPi0LRRvm1YeXRFgRM8ENB4
ljTTnpWl04aA6MiOyjVXNeWQDvMvhlCV5N8/A6u18mtK7OlvJUVrzmKmHkaRInmp
oW6HkwLhz8RDvcBXGPidwaSpkoDu/opDGpLN9kBzWrXl9g78EiBEMl3rR2PivMmV
Wzr1kMbjo3KFkdmuXG5XYm+ghCVxzi01ru9o70Z2iKAWiLyg/SaemJSCLfJxcrzL
LL+wPyh8RVSIJicmWnHuIpJiP+9e0bYRkw3/L1njKW3R19FzSqGfHL5U7wdhyy+L
POJkl7+Gpbw/9Y/oOAiINKbauTqj7InCkndNYuHi+tR6osKaviOFyFWPSQYdlPzd
cuviy3vzFf5yuogqEFBh5DMWyRWPkld3kvQn1OQyoWxQP2E3zenZe6wezq+3qrR8
7UZxQPzI7oTaNRRgJwt+ZsJVhyrjtofcEN8ynJhARAaPuaAnTwRHlV+R27dVU26a
9plnmE+ZF9HuBD8MWlUxqVonMoecfDF+ACbSgA8ZYcfWDAVh5xUl+3hoouZZMRG4
om6HQCeLtiIi7xWldz4y4FhRZmykDdAfQhSVPHXht/ULyfZdFG8gv4or63jGCntl
MDLVxFwbLVkmsHSbYVcmneyDOY3I9Sbhrei0BQ6Ve7OgbnHTQt7J6s3RDZ+v7ABn
4Nupn6jddAHovdYn4mtzw3GoPPW7CaWuWMpAs7lMawxdkdRaKpjmvDJ1872Mtuqg
euEkW8bjYNjapQaFn1vRQrIF15o1jGmX8/5gCiDisGQX9L7Su32rXhsaw+aGMwvS
tJluYw/0rpDDuhvaRs+oxlh2c0/RN+SmW+LDrcaDXTUVVmth287tmWW7PwFeTVjO
LjXKtUsbbtpdwOJUNFiPHF0uEewgpUEm2OpojCVBcis3hNpNSE/7t7BrkuFOPb/C
651kuwME/VFggVUdhnu59ei4ArbgSX8a+IOaSjCYkA6EhYKDZX4k8js9qUwqNSUG
sSNzI9+UfznaBtPfKmKxaL3o0ZQm46azNwryxj6CtDMjau6NYySxPdNmgmieak8B
VY7zzWUEW4If/qXxxU0g3bJW8cmVzznRV5ctI+/lLXjhi2dTaHXitgA2RC740Hf2
5brs2boO/ZjAbL7M8BSSQHiMYnRjvEhndLt1NrEMQxs1eWgI4EBd7mIdfGy9tl0q
pOaQwcis7uXzXHC3PHCxar06ltwqkbwJdeNA/HNiT3pjtvz6Q0edTPDh05IQi58H
jrRxQEH2Ds3tNetYhA+fV2xxu7gdMkW04DZ+9tPYNNTubcuB78VrRxrHe6Z2MUpf
aS9snnwo1/JlGKe5tZgJmeyhSJIf5iDdedRzTkbNS2SWgIfIZNUgOsAo3su+GOda
x3Bz4rjLnCQ4ODrwZEw8pqgEuFgCbhqj3ZPqSJS6MkXOc1sVMOIemO53FT6cCsyG
fqXgqcLAuWfY6XwjH2IXo6LWI7h/OCboHil1bYaX1ur35cRGEf9WCQ+W7AhSipp8
9oFJ0+qVjgLaCPSUtAUf5W6jGJS5XuJlQJTv5fo00nnSidN0w4LGsBSX3IiXFPFP
61Wv/zOzeqlJv32NAKO5TJtVYuwQEXRTrvjOFiDk/CB+uilcKb3bml+qR3NvJ943
TG0b2/Yz3SxOur8wqoyPwd8wYSz8IFEDPy1M6tPTaeAUwFgQaLM2aM2kqKGHEMef
5+KQTimLYZKoJK7H2qvarsVwGBY5rrIl+RBOjS5Iv8z6NFmen0SYiI/7OAymDBkQ
JrsUIr/svf01KAfhv8rrrjzj0J6aLNdkrfisYpN0ef1QxCdz+DhrMOC3uH9A7wZV
d0sKzighOU0yp7tYPsSGCaSR27HJo/ZVEWErgn5addfk5I3YAHbl7cWfHHKVyQZu
nCF05JMLn0t+ztHfRWCwVMysHGaYIFSc2aFJwQPC8eN6qwhPyc7SXbk1/JMDnejQ
bU0zbDe+N/FkA15lb5BUfnRuDtcM0RLqZYD7vPNTSuEnTbCENhQ7z+vwX08zxTlk
WV5T0kOzjl4xax4Gt/9vTJ21P2uVdsQEYCcDvug8+Eh9wZcyNXH1ut773Mu6V5u/
3W+noyenhY89SuCSWFVcLskjOPCaesv8DavjgpaLarlg9vg6cqaYE4WkHkqnMPfL
UjYKq7mwzT225OTRjROrPTx1HyimAuajAtzn7mu5l96vlsFNkqok8Bg+aCoKlPvi
EBai9+xdZdtdohchOUVbP4PHgBwQviXmjp5nPm4QQMkEB8CzLaVjdZ+1JC6NzlTI
nQteVOsgweVHuye69RrQz/zi85Mjw36Wt8j0HPcXs073Tv/+Ya+ffJd2/wyx+T+n
Fzzw6db7LivVzxzfmmqEqoAhCQ5jSNXZW3ikBoO0h03fhRIBmpQuSQ74X9xrxMVH
AbE7E7jixpe+l65Jjyv6SIEsjTMZLbto9ItMphsQg46mFaCWDaVmjMFy94kA7On2
Km7fPOCnbGYWoPCnWjqVcVyKNSglRrc6afgq4RmZCf0TPEr+oQe/yDQlRbS6ud04
BnanYKjBW+WzoMmATIB1thpJVyi9P+BMoFBHb6BGOHhsU7CmY3jw+WffykFdO35j
Fjw28yelm7nK9V2qs/UggvaEdpVFQ67SW0fEz78ToZZLOUXhy6CtG+L+wSVkIly1
TO9aVHez/4AZlwxOXmtb9MNGwKWyTs8avUI7YQyMiR6c7mkWS/oiBQycA3mF9GsU
bN8f44PhEIQDzxJYwZzhdIxMc2n7hrcMAG+8BeYi1vqGctbgoDEDwU/CCOIcXiMo
UY2qQ9XC7tQdxknO7VrtvRevpgR8Jfcsb2AAbxpKHKSmkgZi2RwW2Ivsuc2eERLL
yBAsMBP4yuLWT6DiWd4mek6aU4iRcplT3HVNThfh3RrzzhjljaQbSQB2MAUXXXH/
nylrNkuEQBL+27gFXe9yCbOaz7SJELBp6kRMwZgwM/UL+Fhdl+S0DsFBtV2lSx5R
bTygQyxaI65R2uLTvJOK/Uti/kFympPYeHt93NiCbXpkDKZ07zk3sKpDCXSoaKpj
V10AqBvX2QUkQ5D3DheHPp66VahlZ2BqHtra90Ntd3bwsM9JbJFgB7rMjpb8o6Ru
+g9mh0nsdZPJPOXdQowAggqBkL0HDJdDKroKl5tLhFNB87qwzd1OikOaUDMz3oMI
Jult49nIBUzfrxy5f3HBbaB/wA9reiDhZD5BbwqYAZ4fUYUTgDQT/KSf8aVYtbt2
bKpfI/N2UiFT6QkMvt3P/csnGL8NuGI2vcMiacr9/SKGn2naRdCRBmAujL9KX6cu
g3FkeiDjMYFRYl7mh5iA/dmt185U0UiksB9/QlTT7IfMIoEe/WbVk5/ZoazB5OuQ
HXIAopfp0boR5hkGLNpPMZnXzyc2naNJH3m5tUlm5nwR2hjMGX8trsS4oirMuw5a
Y+T3loakIWFnUI4WzcwXnmKZfSuqBZSrq/spx1G3QHUTsGUQWX6ECT+97Ek+wUob
FyLuC+WLw25fRChI5CBbUmRVreYxcN6iLlx6A9J9lk9Ajd6GWkuEor3+Vwroa/Lr
nobp36W8yYzESpvdpUChBuzbLGJeYs1DorbfOHpd9FaquTPptBl4Sy4tSwjzj2tv
QcmeXcbO/XN7WYxwZefoEQrhcP6A55UFAuSukF91iVELfsymqNJ8J5ni+x8zq5uw
UfKpkKtTOev7dqHCvngnVKrAtr88OPmfVTlE4ACyLXgvwNQEyj9kVEHGopjrU/sR
vifXIUtKpbJJAkMEnONTyDvPRCZi+fyj9Agx+OHl6Io/RYHVX+ncxeZoBlTIgl6u
GxobJ2KFIWQq2+HafJjRkXwQAcQtUvYOLFgZxBbFOWqd3qxUSs3yB7ZZKySeYBmx
VZ0ceRxzU4sDXfeSRJVD4Sgk7u1JA15e3cRovfOwiCVuGxUWEM7HFAFmu1t12aXu
QAujLbs23iKJzOhVLkL5OWR2NQkT28Od7Ten5mjqN7G9nlFnrsC46SMavltzlAtk
+Fw70fd0cOuRc4aN81xWFqrCHM+PU6NNe5NNjb/u77GpZGBKCKthtSnqBBTdHfHL
4HGearGkRKpLQHVWNAGxSa9ha49d5PyZRrSLgirWZIR0Y7+2yfCULBp7SxYYsC2g
2ZZrrNzYUedZlgEaUtxucxucJTVeZ7knl7i98TGK83vxCYHKebqMY1aa8c8mW/m2
v7qjPK73JQqRjeWGJBnE6KFNv6LrtIwbZLp355F8Evmutgm6+asKZyImPUBajP6k
vOuOD+B4Ls0dLcL4q8iUGB3NxVOJV6+1D/miwnddPhBLObMRU9TLw/vvkMJA/mIA
r7IrXL0PLxi+sUgpGpctmdJ703DCzwp0ItHRY4/95qud8zvcCZT7J2aY154dkotI
+QjkJDddgRhAUTbmGUWoYA23tbqUfoNqb/sV3iQ73nO6eoqI4J34x/CVFRyX/6B5
dt8NDJULb4wYtZGlrNRuKXZCLvE+dnL5wqgTqZGIZOF4pP1+3xOBezIb1W9wFupM
dT70vtAibMxnfC/oIG0946NeHMFFxFgaCDBk/+Wt2r7zw0z4CheMH5T5FEs3vYd/
cj2/Me9bad9ZIywscFlRnWHhI1B2zeiBS5oPU+0oLjz8Vri90T6KAIieoPgFSDU2
OYRlNz71H7C69TrkXkdlz3h9fa7eSX4W1SI41EkSSfw9TjZtEKXbKRHGW9oyfEO+
o300Go/X+fJBgux8jrLqALSpR1sRJiiWA49tL43fq5QsMVKCq5ZJNcu6Do1VCDlK
e41mL/2Qq+L/7uEIsLh6AKRakMqJtzeDgBTCl7Dy56UwhRIHCBoTlfP/hGahP9F9
IIajRaXCANQXciEHy5hyHKCyNOxMAAjHHGkdPySrdJnjWe6aGZOoTg+5O2VbJ7Zj
BJtbTjYqXjypk1wzj+bsWUFWDjTEGxtqatNBdIRz3eNaJzAW6eNOl8B9uhfSmD0U
uiWpwKy1Xo/cuaK8jCRGzPlMPdqSUBoTUvb9gnRTsYWEa/0+/6FCn5pdCJfY0pgT
KlQ462oJveHo3YHGF/Rglv0A0yE0LX22eBFmKuk/SGfw3yqSq9DodfI/LNbmRRZS
Lgs0TZtrNOarzg1/3ivv8LjTciDZNCqfe++AS2JZgaB89zVN6YNF9LgfaaL84zAp
43Gb4QPdFOiKvV3DwFnuP7Q0cf8zA3dS/EfsOdSI5Z/qeHtjCUEqQvNfMUunW4kV
XDJPUQ1pMCQ8+NUGTj5y8w+ddSve7u5Y3sCoK/9oWbdLy8xD4JUc0ofzX38W80CX
tDrqswgjKRTNNtyMorra6O1IEhvA9GL1Yx62qECFO9VeBLPikn7qVzWEyTBwfKBu
g2dUSObtzY8o2HgWsQE5NC4Ubw43xFwfyn3bjfXfNTTnEYagc7p1SApkQkZIsGNn
rGhMZ6Ha8eqaksbHvNAFMK3zL1dFkBdSQO2CTvf2E+CGEmWh6ZqbcvFrvz4A5PgI
m0UHjKw5/u7ovMoaMEdvO2WsAipomgx/CjSy10J5PXYNn8Y+m3i22bTPVKlW9i6M
QaXVI03qI9u91CJrsarkzQYwpFD9lruWDVep7gfQJkbxcsKTy8MnLRTNgRTq18Wk
C/mLfO1gxaTcP8Ud/cxZP3trfVTNytYfbHrI4KA2eh76YX0iGpTc1o7khODNhoWM
4BUG+JssZAcyGoRPzZqVVV5NapXBb8QVtWCKvrsskfoYZSyb75l0a5RtOSFjU2/P
g2Ji7TuFidRT7qH0dN00YX4qv+VpzAHHXFilY9yq6b6MXSjtc/fSTC9hg3h4zC/P
Y/pUxeSCdmIGb5S+QGT/81HqI2IjBhuL0XNZBsLbpL6joXcwZ0kgviq5jqvgeJcb
O4iu5heEZruHk+CpXu1s7t+fawRcH0cUMnCi8+g2vAljPNLqAsF+HrlFwk+igxaK
/XzPC9SHKHFpYWPe0ZiQRBEQN8lnoqGp5B8k/FNOw03V01GENEkcyay4W76PtWKu
wpKFF2wVQcO6Vez8wAQyXyuITAPYsYdeqc12XAXCfLO+YCL5fDo8Mw3KL0nYW8nJ
pA+xEGza8XegZKEKgOylAl7Pk8lLuWgC9MnDFDt2ZifY+XLqXlmRBpr+QS3z31TC
06Lkzz6nrxZuyPCkO+cCq8wiTeRKCGvaiI0vWJsNEvdir69CdQ2uMuiILYdzBCps
WQ6Fx4xTizfy8PES/WoQ+Bkl59B8IZbBIdeTIV8PJwxSrfmMdyppdO7G2vZQxpbv
CInJ30bdVCMFwMhfXgylRUJHGEhL5dbA2oWzVAHU/FSFkptLL5OTr42b0tvX4PxH
nqzafnIxZG/zYBILzWVAYTKl+swSnozlbe7uzt5/H7JTW+mG8E7vG1yV6fVLG2tE
T4Co1naUxiC9ABALJlWcXKpdiS3uyLWAUJxm+01eiQnBsXCKTOrLrUh5Y0JTEW4g
nxAsv+DuPq1PTVJRgWytTz1bdcqmiNXQO4BKwvb78ujde6vbfCAuF3CON9RJwZlQ
42wxu9/tr7ll3SNS+g6ehBEk/iEwHsncBdJZzXa0fZTr7TjcuBBO+MaKyEh5N/cQ
46dZT9nwywWbDkqv2kWwiJIocVEVY82gZ+JFSzb+OLS8Rjd4198DrPhC8oRlWGZ9
u05c0Yj5jRlfnnzalj+o1rzI6WGzx6J6BQVyqZJvGCOE+cmrGZzkuwA4Qbqk7FCr
w241n3qQ2gm9/CiBBDHULQ3AwJfEwTmMifVsJfL5ZVEzqJ4+rZQkIvM9O+M3LGhD
fwQHM/PB9P+a2KIqMEP3mPkwOVm5CbXJHY4D3hV9G8dEe7VW+Rzbz5NwU6wjONUX
dEM7/WJGpPa/JDSsBB5GsjvcNY5DINZDxnnGHpP9cle1TbUUb6JofeGTBcDbrVhi
RG0+JPog993OlwlAtstTJMRh39sOQtrR8aD9PJBQY1WQSDw3OlZdf7c5zYUFCKC7
L9nawABHaF52bmsI+Vs1sD4NnsIvqzTtG6TPyDipr4QER+FdhhWxiTCl0XBq4rb+
37ZLNkp20kdElxM52wHT3sBqbHEpBooCVa+6IZLlRLjKSvTEIwn4eqNrWHxNot4D
DR84qXfsKWXWWi0KIqHORCPg2hu2D9tBUXo0lYPSEKgNU9odqMP62K6ImoNSS5IE
ZUCkPHSQCutW0IUl9y+cpXfUAKqW0MRTylsA4RsFcQLBlppxujdbPffYdqRzaiFm
WetmPs8H/R8ER/tBzzYuSkumFiiJAxbc54K7GxujCtYl68GEXhZk2zol35Jbotma
xEjHcWr4/W5Ab75KsDXEn7MCdyLpOL5VR60hISbaWIZhZ3b/ojkaf15VHV+QQsHF
TUhWBbK58RmKXbdgLUEwNZl9ECWsXlq799WnWdqHMl0FNKijjbS1Jc1zHZE1nv/d
H1zZizfyWleoy06TZ0ibuJfR0RVXF70d4nLdmoHL+Dg0F+kSocPQmXUi5pge2NBi
yTBVI2j6RpSWmLw5FM1q8PjqOfaHpW0/Q4Q/4488g9HRB7rxqoigiylSaSPxkZq/
rcZmblW4XqL5CJw3dpi2G6Tma4mJSw1+ZofGk3dmaquPRbVSIpwdMvd2i0pCCpH6
7wFPYq3I5jjpwkZ2fEIH5EeFj/1G+1VQZRRvRz7n+FAgZ8T08U9cZg1yNW/rrdGm
XQVO30cmiy6flwEtufZG+b9OWokW5dSsbWWRAsQRD6fSLEC87YMGAnrivZthcnB0
EJLKjamTkSbiAH19nsOU1gwGAbpy0JVhhSl/0yQNla4VJHJ6Mjag/ogHJJBU96hY
CIw4QqejgET+PN79F3P8XO5LJ5FUHh+hG0FPs2RAox30EAfBS0R4HUoEmMv9uOVg
qczx9j6pziW+0R/XNzLLPfSV8xFWBcvlNmI4Fz1SOkkWxov/BsYS3oNPd/BDkniH
pVkoHAqhHwpzeUy57xXIhRXw/A8ouygxXlIJ9rlaTNqbiKD7G/BGm8FT5nbixD8B
rUjmkqn7ze+f8C25xJN8Uaq/A9GOlSuFIOf/1duPBfrJYAmUdLTT9qFBM8ER77WI
OpKumOA624jWqQonAbuBy8PsSU+TBvs1GD/vYNYfHkYR/gGX8+zqCifNQMQeO11r
uBd0xMzHjcaTx2hjxMD+xE+t/2lKv8ZwJZoHj+pe+XwhZ3GvjXjZAaMaV+HCacDV
w4wEQ5ikpMNFeC9TrZnJ6+L4UTEV0bJkJZoK2Aw3vB1oq6X5QHnNeL9HyCJImRJm
hnogHE7DsvYM5NPyrIrXkiPIR/EHpg0hOUyQrGot/TrZwNwbtnc2p4Jk5VTXmTGQ
YKwJVUITJTMvsDbqnUGzmqMBrBrnheCm6DqcS8coJhp+g00rcRtrgCJw4eDRDV7i
0ZDbN2+FUQ8VLkKOadsHXKavQVwHMBa/15L7GI7NWyQPt1mmom99tEXw642hX6JB
za6a3YDQyqtC1nJ7nUYuxgUFSf1Y+Ke34OsWyenWXIMXR08tHtX/ZDFwsCbKvAwG
tB/zivQjudVlcqLunYr7npbIU1evYV0fzgAt615IB4lOKYcVNrDryrWN2x/wc85z
3uh3ImN8iHXZkchBtebDC2SHDXK7EjJLrB36cptiRNXkvOITAsL6IxT2peWe0gGa
D/XqGlaBQoTqYoB3WJoA8DL5Ai8V5PxAA2hYquRo6/yw+kRw2z6XtLMhOzHjXRW/
mtJQetsMF+WQdf8E0Z+0/6V2gNO8ndZBUkk0IPTPym94KoBIMM6YgprK2swVkbso
UHmlfCviCBBUqGFrJc8LC1OheJ/Ui2LClOpY98eRT0rLag923L39Oqp4T39cMrFt
3MRV+CPfAOuSxsgPmxG8p5uVP89rJscNnEq0ofLNYj8Qn61EkmNAAvEwrpHA5gdH
qdj3NfOcpAcur/qHI3pTv5R++42IQKyYWxQdkLpbClEi77PKxjzMukNMuDxh3qO1
973fKN8jgV7qaSabf7pQf1rNjcNf7c91bU1DbMGcBNz57CQ6P09T9uEWBboXdgoN
3kRZ0QKoi7hIbN02J2nlqBwYg6wFKQO4CaiYD8KKbs3AZMoZpQ9Ag11EV2lJ/4Ja
NVyo58Pqllkg+j4SktoreSMdaUOVQ88wbvZWlbCoJQJGLcbjKQjCDu/phZQMUlXb
Zc8EP14zgV5uNnYEqAWaf38M+OW+m/yhIQnaPRM3MAfp6CkvyAOerAoM/At9OiTP
Bm1pIDiEHG5QF3uie5IlhVdV9vE/RpS8eZLExnr5YzoU3p2RikbOlX/7/czBek4v
XvbJNGn1PGF4iBGcKjJ9pjARbVWgJ9WKwSPv6TSn+k3XBTBLo6e7t/qK5/yEIUfH
orO/YX5TfU+1iupn4bDo5Dn5PM698/BKNxE8SDU4959IkHpiDWVeMNDvz9t8Qu0i
bFm7BZYcvizhcN8ojPpADt8Q26Bu3vuhdm4sSaVOv98nt2J2AjO8YEz3u9mGH2oc
2zpS3YPuH5legsreq26rCQJtanG6foGyBIOjvpTTtOShPP8NptPtxlq3hSqci3h6
TFwc3CUIhMmWbmzc8zs2ywhctsl1QNJCB/BWTxHdOmk+0a5cqX1Sas8kPRcV3dph
RwrGg2jNgJgeuKyw9vKOUApA4idjA7hRtw6VDIW/fW5oAMxacjQTUjvXq2TgkP3t
QgKLsxCH2YlB+7mDVqOHGVzFohZT87nJpmVi9S3EeiRMfYD/vKdw/n/ud6Wkinic
mKaxurtNm910BLgh0xjmYYY+TbRNP6lD696S9z3x6WZGrltn9wzQO3QhGdK8UqHF
tyYFDJI8oKK05gDw8pBlJ1eIl0q67SiteyQs+kA43+OAJigDTrwcj9amoP0WsxKI
YSOe15PmGbj9bbd8TuAUENZk3jGWP2Datg2L5IKxyBwBw+v8DZAEC9BjvT0QVljD
ajaY4ZUG3DLZFevxX0KOkkeXfa2Io0EiVCJB7SNHzN603ZoEuINVtY2tXm3EP0c3
T5ZLiasOcyG9qquCDgYxaDEzNpiXLHYA3K1O3qoZ1VOEaLo8idHBoFshoiiozLfD
G41GWANSKk9ACeHbjpKCOSv55eDnb5XFeY7dGCOGThRtyFNrYNxR3kCnLd+IZURz
mjFhbZ3nWFrzPDFh/wpIkgtLbssCfrEKnsiySOK3yUWiWIqoi8hXM7dVQNbrjKx9
xMha9BNKvemYA6au9aEmsOFJhFXWvlHewh99GNjzUysODi+KirqQsiujX9Tv5nSN
xbHKnfWXff1+9Y5xYtCiEsBazCxCun98swSELIJxRpEIIr+Pdn9W/doMiVjj9hLG
cxwi9npu8SiRqECiih6rGHur4ZVEu+s8TEcNoYWp/sigEinPT1mfhCT8VrpbyKaT
xADxnPAhhbJr7YJ9QBz63JvfTEbTVrla2LJEWkaos29ASNKT4k8x1InIsfGI+7H3
Lm5ixSdstpFt15inq4vXAAO0+e1aECQCISJDxZ5pqPC2zxXeW2lwUmJD1obHjZ3Z
wfPaPKj27GAl9EG3ssP0DOMUT56XpHvaG2sstId3+peutGzuZc1GSFr8pQYb4GMO
2gyO24Bgm+7xsXfROLGUpPJ0gxsLqCaaiom8uCTpKQb1PaBTqakh53g1qZe0w5hh
oN9WaXBXm66xLpAVUqx8DjAFKRQgG5+RKSaxWXJKefA/OGJZQjcMO9U9tF99nduf
586Z6I8PEQTBHMgU/kz31PKwR+DJv424p9nE9AWIgmHZmzv+UiDQ9D9trvNrxrjJ
AQpM8UTiWCxWLOuPbRmK6JlFzzgyEEZh8aYyF4AE6jprY5y3zlwYdlQm7C3pXVAB
jsqoP0Cpi3W4SYvLqME3rJRoaEX9eQ1hdEzjYK5gTdP+fwKIJzsuuIBylYqwRGzT
iGYjYKgu+FPcnU56e4F7RkQdjyXvc97A8x7myCPoJK8xdQY11nNl2uaphuSxywB9
GOhAiBHIMCF7RYWWl4GrWcLICH5f/tWFdfNHHoaKRDX7T+BoDeCRjJyM/vyrHpVp
WODp1g0NJZPZe4WmOed1XkAZtEFtqnk+vLXZA/oHVA2Lh7BI8+uSH39nWmgMbsl9
p8R/izfMqsBiIqyb0EnFGZCFAMjGPz8Jz5nxt71wxTPW1OcJ1T2cc2w/8zsyr2Du
GPEfLxydP0dQWZzW5obc5CoTtK7NizFV+XsnoNxJfYLX3FYlyIAbebkbThSiDLC2
Ye2B8H5aBKec5TpzNvMD0vQE8GzlPZoFZXZ1RsB7ZVHrnqRS6Yj/MOHVRArO5rD8
8hluOPIRN/imeEbaUhIfOcx/6XIem0HmwNtwWDKW3hDhcSsa5qIZ5fvR2Gu9LtXQ
FzLYXXyxVpIbAcydHtYQYVd9+jA29yDcbDKP8I2m+gM+vJjvAKfhmRTrCQiGZTSw
2+TIHXw0n6tpZ8CQP2+5tJIutjGTv/D2wvXz6WWiRtPnnssd+qpAH5m7jZVcr1WU
Mq6huaIUS1JA+ylPaNwWgJOab9gFsbCkQle+KBBipny3FK/uM+FLpnryELLaO25b
AREoUdBMILW6aTkkmxWNQvkJRmiX8F7XaLk6EwuiUgtYYymCgRXsxEiL/NZ9QrRo
3v9BrBelp6zPGyqzQUZ5F6gTBOfDgVXQMbztvz5f5Rs3Si+A8c7q5qUe7EN5SMn9
bDA3JPlhmbHIRSwgoiPHAyDaQ0W0kAUjX8B4tEl7bAKVXIsU4LzQ0T3xI+KMO6iu
c5LEv1MNFVM3RX0tGzkkOm2PHnDc+vuOGIGkfPqNX8JeWceqdCO0+cx9c0gELSF5
3OpQ7t4cXtaW4VG0o0Boa37YOku2I9nHRcO/tRBMJqwsBbOHZ2LaVRExKmu+wtQn
jjgISND0PpaffpetYrbOkj7lZEweEDnfAG3bjd3F1ULF5IgMR8eN+yhWxKXNUeaN
sxpVOyBr7AN26ImBTLULVJotHxCOSfHSzEzli3DkQmi3gb8vfK0MWEHQQAAz07sD
psjkARHKq8NsHCtgcIxTmzndCeFWsQ/PiY2OzhASRf8wVrcZMOSvN4w2f1SGy9rV
oEXQ11oHv8Ji6o+gfa9yz3qLf+jtDB1sVdlWjBAgQjd6RuydaqvpWuLkXepojiPQ
7wP7V7uSZLYGNEJGJnsR1gA/OhFABm/qQqQUFAq9N0hb+PXepbU6/RuH8lvDvICG
sDiwRXTlaoJWRzII4b2ABt7b6DJ7XKDOWFtSU9TZrW10p0DsFFxQjPmSbEOslrJO
HuKrd7/RgeY32ghTD0HihwgsCmWQUjX013BFz+NTsTTNj2f7SuwvbnkO6ndMJLxT
8Rzd5e8Lrr/+J3IBcIBmZJS2/ZxBO4KjQozrJqykzUyehQouWrgpmoEWgLZK2050
lK5Ha8dhn4kaqjCvWFPcfxaMprCzRFVyWBSsC5vo5bg8zm7PD7SI4qbJGwZxKQ8G
oGkz0fvxvt5C5o8oJt1KDuSQ1dkqzzOxF5FElnj4darGlboaXyY2r5uZtEaXbNb9
kJ9C68GRe4bAykNY+vzabPjMsLEgMjJA2krA+2s2RR4YAz/r9SaLb52GJs9JyhYg
mxdqfYXleGb5gcDlEkOgN2w5phJ31kRSWlkG51ShzmhdO9rOC0gjqgC6SRgXVo3Y
F7wFZcxmvzE0H8QI5Jn+xmNSBgHmdCTptPIyYb+FsNiJ2D4U1xSTvJEhka/VOIP3
PF2LLm4aEmveujgymd4ExcYnpbbbPVNRd+Qkf8bRpdm3RSEyLyK2YleEoLdSMuKi
4afK+NN20kiIvwqJ+62IUCIq42ocBc8GD4AXgoWzXOP37Wu1NdQiLxc2Gy7oCFk4
F8+kPAbs1AW8ECmyHf5LTZQhd2cGM8Ht8PXDOtgpNEj8Qxghhu2GXYvUGuFnGdVO
G/Gc6XnyyfI5277gqZTcKmHAr6/sF9ueYKJUak0u/60oaxDt5+gT6IsJ8MTffgv9
VONi9HRg4wnR+7EzjghV2n7/4uWJ8HTCMYDfGij9WlYJ6GVjIw7N/IWL+p60+24L
Q+aV9HS1PiMoU//RzPFXE27hkGSK0ZYnTOAvHDYQlteW628OyJpmSblPkw9WZvXa
rB7H+PFpigAIv1mg4S0e0Dd5DitCZSCFP3cWEcFuzldNN15Le9+rmreYKDc5vHYP
3gkoMXd5BrSN6FYBazg8/tMmdFjt8yWeFLJxb55m9/VI7AsnLr+QcYC5P+ph6OEl
KCCZI943M6oyMzcfsNUzzfNfmSPwwLHwQEpPHvKOTYpNDpUUhVI23K4AFKBMHbQN
zfYz3Hy3h3cIyEjHxwste1J4tv72cpWRoag0F4DGtlYSCo8B1s3JwRHgehmfyYKF
td3oHe/s23+EJQnRnfIvuZlTEG/6dasCpD4tB1UUqEye1Ny8prG0RXK76TMw4Wby
QtbXsMLrA7wWaB1/2huJguRJ8W0/1ye8sfAQmwpxylvUN0WZGzzX1lzOnRj4iLK6
tBem7tPggPxQcJyZALwoTec5tcHY542lUgRkR6Qb/SIR8lwQBCnK6lCXYbPaKA33
Nx+Y9mSupcD8QvqTlc1u/op6Utl7TysX6M71v0BnUWsA5jQ0PrBx6lAKYh8dMMT5
geOlWHk8l9SToc/ZwO8JhEzTXU36RI1TFLY/r9qm/wW7YiYEcG2zn3w4KlbIjqOn
I1+KfZ04tp+yFn8EK3+dIqs0yyMtaNINn9StjulfwaGoYshqVoCmiqe6A43O3Bxd
seLNYwna0XRefQTZAWt48nnvw7y/m2O4jKpEzhhnGkrt6XIKzGNGA2xigmjpTbuQ
CxX5fPm00GoXQ7CgHcSa3hYDmJYUOfKFrTScK4Iz7hoOgVjHVmjnytiWrhM42GYo
deSknX5Ku2qa64dL+QexLKi2yAR/HBu1ujA4I9c9inj8fFf/Duk8Bts8IERs947b
xNc1ws+W8luoOsOtGONXeXUEjZ5/3RtrfWfCIdMtZMPTi5LlDLn0MehNOYYhBfhG
DYixdEnbcuXeK3AVwU1tYPD5domLmXtuBflS+lr7uuF9AVE8M0mC7aJlBihqLnxO
0xMAuymSmr8NJkkM6/fnPdgEUIKawef7pgCb4ZQSqCnnh4NSHKyxuh0kB0EZ7GDo
i1PUETnJsutS0vGwTul6O88d5Q+HO7tA91VaBMlByUDapPSu0MVQyjmI/PYoU6np
NXqpeeqEqI1spIpOGcnrNZzX7Qt29QSTc/0E3cdqRzxicd0JMGZIQxt/v7P9QGDE
PKwhWRRMu4x1wzGLWvCEVFIKXZKl/miekZEknd7XS89eQNs26Llm+2AQNS9Stk/i
Y0bKDHZ3+9p8R/vq7ow/KmZpIfGJ4O2y14+Ea+qY/xpJgYYGirJiluWAhnbWmOJY
+WHZMwkHhoBwZWGy2QhjM/puUNKPImGJnh8ZjFRic28x3wFrpFtcwA3xw+xy5q0P
3rS4NG5xcG3PacnYiD9P/S25GXVXp/NbhRqpUigvzuD4ZecXwBoDXye7Xb48PgOC
+uDs/1E9sILX1lP4ZxYdxrZW3HeT9IOaIEBQI0MJSRXaZfzB51/Kq8iyKtXeigT7
hc82iVsFa7uXYZtpViuDwXaHM/wMiuzM1hLNTq++VJBVvVkJ2jY7pbw8OYFybW4p
sFijapjrTjVFJn/SuzJ1p8E5ZIY0IfnG+hr/kNry+IDVGo9Q31FUD9OE61/PXIEa
t9JrkbQpluUtH8YBbNB5REo0NZ4l8jgievJZIU8ATCeb9XajZduKMnjFPQJTG3fo
PG7ijrFQbphz5/ddkXZyPMJot0e0aCBo8jEUUiFCiuBkyNZjFfzBtC8oIlKarKfw
gjDxu+/RnRDn6lwH9HS0sIikD8rBYoRsk6gZOFS7Z5vd1ejhWxQztig2Y5Vp//Uv
WKbEH+upmVU5NH8xAW7wnLLBFFouGirhu7bKV1BMtwonrQ3Q+66AKdH9vwfo9faX
o4f6EbJKEsIIXs4kYxiY6nW3baZMmu+3kq72StkQ9WX2N4XFRHt8K2p00CBjggMZ
7X3v9HrcoCBGOODDFq3SOZ4HkC2E0hZlmb4QBEAGPitGWBt+u5YWcAfBwX2/px7m
nPt15QFA6IEdnaXGAba1eFI/B6ePTHHduL+N63am5JOZJHnwBMAL2vvD1a6kSrJ4
71AiCp1obO7GGhbvi+WRQEC5K9oP9IYQkb62DCmmBu09ywU/s7OhRFggvj0MlIj6
w/k2wiXXdgIQlu8GMiXfCLJB/6KnppuYof0wnxcMB3KbVGu46toBscj+z39+Sk+o
H0wi88G9sI2n7oBmVM96L1OHddVl8/AyytHBpFWgqpPjJCDXzZbpqWmzxTdUsjEF
FAu2iMNp9RL3FX/H/Z3LcHjP2GmZIzhqgtBLu4aUmIt5Sk9VfbCIRF3w9SItJCbh
JKy/0x6NsQ8PyEIllRT+sDom9YnHaYJXSXtlT2UfECoZVDjcbwEsAW42wEuBMs0F
T7IMRfWv59f49OMc17///5IIgR9fF8eml4f/0FfP7MCFoXHMSJqo42oChEcCN4lp
TnGS3kbNqTpKW6XPDW/djgnX5D/DepwM8k0v81QL5dZ0xR/AuJs/5sa1bktBHK/p
4UB/bWlqFzRG5RIMsQkVWNixfQe173ASqaf5IhKBjsGHwhuWzIUAsbhE+jqSdESJ
qNFIzIatXzshERf+l+Eb85cHyuFbc++GbmUMYFFNE5qSyUMy8+9dPh/c4eleZ3bl
2lWxnjqU3CRew/k8xmqcpkB2UW2f1wBQDlNHWempNkeia3STocLESZAwMEZ96W3P
zlzIrCIJf3JapPRLbWTmBCNAL2mXaULbjIu8UdEbTtzC6PKylQGSy6dkvruf/Szy
fUhP7hd02NhnNZ/VLzsur6DQKl4IFOGZhTMb66A2OciZA9fKJPJpaCOl5M0x2TXG
VJAYJiuRfTD3x0HlQOLwjNbtzdmMuqlWkOqlTOZH3+AeHuhoP6GwTd1LwKlvpYIG
J0Ua+sF7QdR1oMtT25b9d2AvwT/6jJBj+XO/fqW7qJWIG0wbYw4TkWasjqV3+v1V
n8mf5E7OxQdeTTkW6qjkipWQLTNw0r/SnThRl82d//a4haJR7vfs+ZeYDl4nu+SR
WelqIyaXgraChDVVaEZ6jjJuMbta+2ALmcylANvEmgomyNtQRiNqhVjFeHFMIAto
8b30jdq/oIMFZ4fM7W/85138uqbis1QlNIevt8heq6E5jW/a7VZExNRSwXVkNF93
x9e8RprTMH+oNOp+lFXZObanprB3pg33KZA3sL2f+QCnzcdJTOrERwQmC6ZbEx+0
+WrmqAOxUl3+uZ4FZYW5x9WdFNuxwfX22IDwHXpT8MlQScEl2IDMVbS02tby+mjc
qBx43wfyIbkQPxiFIwjwxHl5RT6q98SADWp/NdomDxP7LkCAyzQSjaA7rWpU7Oj0
saNE8YoQSWq6LyoLErl9r3yrHf/BwlzsHUC1IjNfJXKK59peDOUKW22WndSNetw6
DQiCBoV3E6nzz/9Dakt8+v7hcoxWd4vNld1t7qbqvUTr9AyJZ/RCCY2v/uUvW1S8
MhXDrUfvAytOa25iZay8ar1aYx4BFKZwBOKnJO0u3T5BR2rIFlTcLbZGvVG2u19a
LG9G7vKRxEVSLAv6X50wDy8+9UrL6SJM1V6FN8ti9aFX5E+K0qqkg7/Q34fOnv/i
CKu7WuXjLgFtkumgYR+OOCN26B7Lg6FTE5kbkTSWoTuXgDX7jhfbVDbxKKxg5+ND
An92z1SIn/The6xaH3pit7JudXuaM4jTCEhROtnOfwK1eVye7ya4VG/hkwK0b5+L
5WnmZIrNfUp5Cb44smIkv3/pO36ncRHWhL7ujxUWBAASKkBcx4siK30HH4hgudGI
WQ4QwDh9KidjuqbXN60Hs+wowWSTiwFmmMbC5LyTjYkeFVM5H1Ej4Z1iixKAWpD2
cQp/V3OJDkobF/+vO3s+2tGiE3R4huUjudCrKf0tOzg9kG1JLBQOuG6D5DaFYIQ1
kpmQLTPP+X90sAKnHPx5Frcf40xiOJ8Ggswpkaw7WCEOm3Q7Lwtf9D0UEtaYZGCm
fErn6oLZpkGFbfTN0mlAs9alfTyzJdSeEFwtJhI/UJa9kgmoHEf7MLx0o6+AUMbf
xrN6PmACLfE7YRLeLJD4HEYH8+ooGGQ70In/SFGromPsT18TVpD4XBQgN6iyDs5G
6Q5394i1CxYadvQAaz+2ZPusbaRVzf4gQEk5fbfRz6qTCqP3QgvAoQ6M0fWJz7OQ
kLrYTkmYhtUPukzrQes7hJhYvNmzdNxOgeAFbUQueztHBkOQN6stWAv2TvYhLOnX
L71qY+q+xsV2qWYavfU3F4hPsVN+M/1CXNCKwMc8biyiz/5HLxWYgriCZ6HBztpV
lplyOoZshuWyrXildel7oVfOUYXgERNCm46aAV14Q8gNNX2Qk4f4HXtJA68GYt0w
AgnzGR/IC2OovaD7tMCirbZZjtLB6yXpuHSEFGifM0PIJ6JgV4541/hPDVQFFkEO
B8x83Fuz0D3wBxfXSjG5jKoKxPCZEvZQn5JsTpuekM6V5ACqZvUsrNydnW1tBmL9
i09u1nbhiTlvm49T7OwQ9251KQD9quAqPrToSGRIehW7D5cUmmLNq9INAsQs+aqY
xKMAK5V5apNjJzRItb97pn7Y15RXb8MXXdw7TonvEgvtNPFctil88FcJCiNkds6K
Admq2WK2pm+TjqA0fKgLHi2R/O7+Ys/oZrhsE/sRVniyKAgtgkxIvb/6ZbUy5eG+
u4M3VofJtHKHcBKi1GSxD/30e4MSr/WSo/Y9rAjbxKy4Qs0oMpFv4yTveRMapdy5
kfq9OInGiyzRPNQEsinZ+DGUnAnZTcA7MVxfZBtFaRBTAkz4GQ9agA/e6kk1PNyU
8+/BAaXJGqknNvqb/QtCXeBHwC0MaK9Id3W0Ap+qejD609gZc/9AMLGcp4bYJ9z+
WCf255efvSzkqyvL0lDY7Hc43uih1WjjPwwv6EDL4S28ymUzD2gBEzkhDQ/3Xw77
ZlvJ89aJu8/QvfwpwQNYdNWRrZAwFRM/Bwfx0w1kZp7tqmgznpqINve3jHYhC93t
xaCAwUdTSgU8oEbG+QB/gamhiDQnnl0HWjN1VxJU0VCU9Qf2Q0gdXHBH946zpvgd
rAsrRnBoEI3yzWm6XhZYsyt/VN5mscKqHGxIs1yr2/atRsG/sRAmuxRoqJszNaXC
F2uP6FGYHHrzY/vj5TJmKTzq0aoRDx/4b+BoBUV3BaERiFv0IqH1T5PV423ezRME
I8k/2m5zbKxmTkLP8oIQlwhNItwI1Iznjb9jft7AGR8uvIlDiHg6jBPI0UIMRVfM
E9BBmq3Jt5+smXKcHOtPvAQAja1z85mIz7LQpRznG+wh7nX8DgtcawiSdbvR1UAf
1nDRnS0PRtiKlhL6cg1DwI0x77GJ5YF+DiRuJOfGZ+JvOlIrjIm8Fam3UA81WLbf
EMBzL82iz4i3jbCcH8ZDA2C9GWWheGeZrvgrMKlBU2v5+onP/QsRhf53qyog1Zom
anXJVyTS8mR+vEIiagmx+4yjdJLNNxrc3UJ4x9NYfr3ZdqwdsCuqM2R7sRP1mIKd
Fb3BCqUUL7MI8h6YxTTiq5262ynvl+SAaRedIhA00OTjUEAyZ0vqFKl7twrxDrJp
hpmY5KPtDPI54a1AxvzNcVuAHgn6IiRXVuFReVzChXgFhrIDxqcacd3P2SPirK4t
IOyiCrAxfeEhMN8wfH8HBX1W2/so7xY5ToTA/jv+IPtqGMBWFhrwlsRTSOMF4jhf
mXmQHmrje/dalGJHyQ+WBiedSd3gq5akgn+ZyGhmObfqjCzm89CpLZP3Vv67KqeP
Nu0YnhdQ5eUwR5S6DR6T/VAnXfdL5CJqjRGXlBQavcFCsWrUpMn7K/iRt6Uy777T
sLNtcm+DC8R382wNT3kNAfIMMLt0L+jw61dzcB3GilqMy+b7rhB0KiH7PRnRWIKK
fd78xWwuEjvtKIXE3uql/ECr02AiEWXXOD9pDyXi3hsy1ED2uSiJdedj2z5FM6Iw
xw7Ih9LlIgxdlRL7oJRAM5S9bymVMCCti2q1qo8u7p7XuGZWoR3kDPzrojcQkC+Y
5RU297Jgw3bheLWaP+rCR0Z8dDd/ZGzpjKHg5lzwbZEqzQU19n2D0wbce4xcX0FW
j1NTMUVyyDHPZqf2R9YIJEKcUkqmZI61+CsZEKlCeDPPi8Ai9UQkkls5VBBbmtCL
Vw+qaNWGF6A4QiPrO5I8L+Eh7QmECNiVhxHWj8JAGGHEqnPrkzTIHzJ6VYf1HRC6
13jMa0v3jNc5z1bh4VKUtlp7xcldnha5X9u1FLapSxNiwmgj7l+BJRgDxTTQecCT
ED7e5c6mHKoRuchFh5IOIdRehNseZSBRjLFeqcn8fcCe32/8UmbF+naavKQy2yR2
qNIpTrARzaU5VDmHge/FO7TuOmGBaQV6woY8/uZlRQPLATKvALwoKzGt6hfAVwXz
EkHBshhP4dRuYHqEDR3w3WfQ/ipxoGpFg4HtY8KpKa4V3h/6FBo11rPd8P6ZRQEf
0IHuGBBIP/qQe+SwKdz65RxSayFniefbfPmnK+IvghDFGILMtjddvcPvPLaiR9yh
B4nuulBvOXGpuTJ8+0V+NWpqIW+H2OlKbUGgu4wRCGjQniJki1HT6u1pTc/8KCAd
kvGzvfD6GsJKVf0IZWH79qdYHEPoLU+ATU3/kmtVtwo2JIkvKZA8+Kut0eIMnsEa
lX3rJf5loYzd23rDWVeghZm9J5N6yNIMKuAjZxouB14ZxoPcMmVSZqjsYFr+Oh/O
quAUaO6ous5GQ0ZU+PF2LYMKnSARol6qMFNcEGniAO3lmK6t2Maf6RLYB14j70hm
llK6bOnczGCRRiO9BxhdlvuNG6DRR3evZLMJsFyz7PcKkQY7AMC98u3EnekLykJe
zNIWlTjBvxCiO2c+7bviJP59c6SxmjEWp1Jl+k+uvwfAqhFuYg4gzV5NYdbeXqSn
nvFPcxfxSuoJRJ8pstQaeaE7ipFU2fVGvVGMct2LKl4KXiOxHA0XKi8vrTf6quyL
J1Sb57oxff3SDAKmEH8c33cYSRVF0YFN53H0VwQDyXtA6NatOnpHhNvA0EkzpWZo
aeOoqgx5cUWMQ9LVHViuK3IrKwXjPw3g8FvNqBlXoBxwKqDbNTffBLP/I3EJlKrC
ZW+P7x1jaZXTgwpUewLALGXLKDMqXvz3w8uXy+8JOXdGwBLgR/TchHYM1cCzJ7HD
hRPYlMBt2lzvzeH5lM5tyyZDNO879QQ8DrtEcYSKwieo6FQqJNRTp0W/ZZdCMdWh
2Rt4kVsTbFdGsgOPP7zyuJGcDfGKKJ8ldphVTvCgNAbym4Ak0upgUJTEUt3gt6fM
mL/qsMIKu7Z3vEbByLHtC5FXCCk+BPAFNlF+DJ8UConWlkCUoF31dCrFTJiKQkw2
O3VrgSMWQeTynaXyc4/K3V79+c9sC/Tv9hfgMjg5N3WsH3VHcQjC6akEuVjdVAGY
9Y9s1P9Mco93DUMZrWiDmrFrhN5IsMgMVntVDnJ+UMh8wA6DPVH0yz5pihavHoxP
5p/JwF0qXHrrsDhsZCCs+oQPOVxzia3O4pzWnQnwKFBdoMoWGJYf34S7wjwQLmKD
+DKCef3T9C8WaoyV34u8zGg1p+7TNHvs7eV6N7sFZpD/pK4AaHmI4LlDmw4sKDOi
wm3MyQMkqrUg2XGbkIf2EKAuwZoRwbtBJfGt2wlySgJPYF+rR+Rb82ow44rwTMl/
VX8VxAZWL/C+QEveCCWT/mceUjrHi72GzIAnBhhxJk0KhSDcn4tEwYc4vMccYkoJ
1STIOQ5badSKgMIzHWQR7d2HEGteE/78Dzq6Jf9HVt67q/33k1D657JZj+naJeyF
Rbf4PwkLB7ot+GHFemoS1PH6F3OS88OPg0XMttY7HR9MRg/GxcFtlEtModQlJ/DX
1niHN13XWc/qSbCVg65p8A+1ExwLy2mAJY0Gos5dtFW6HW6DUAqqbB5ehrgUtauD
SbTw7pUcM3Cdl20nl/VScKSKTSVLncKYSv7McAON2GNCKQBd2vqmqW8OhXaPMBC9
PZ6XDDl/Xg3jNRJT3qk7Mqy58ovX4V0SRpb1fnGY9FQbQZOx1ozyQ5yesy50REtB
N5f48RkcGccxIxxOY87RoWBFtSolwnGhd8CvQZHIDrf4xSAhfAlweTdtRi1wyqPI
/pe/Jp4V9wB67qJzsOorwWuSLjJwUvm8/lPsvcNvetYkk5xqZK1TpU+h31t/OVYH
klsFKKLksXJ5ssRU/srVSKUVBJTG2errc8SVznChQR9HfwEzxOsPs/i+eg8iX4Aw
LH0c4e4Yvf2Ynk2dnBpR5ic3NTmSEOkr3IfOLB70stTLK5RVkI1WS+CKQXzGVj7a
DKAzNg+RJsa6z2izJwAEM5KeT8NEIfyZDohXCoIuJl5kKO1IaHbw+FRiHUb65GFy
rOnZZBI+a/XKsKxsCNBIIKGLlpMOWd4AZT81NZxqkg4ZE7/zBsP8t0JEhRgwOavo
6haTgMVxvnb52zswsOK/05Lin4Cu5wmeKVtvHACHsVT1IS9VoQV8CUipHTYpFrEM
dp0fK4X36rpcr/8exluo8XV8UhMLCxSnq6tFgdW3rNB6VkB+nwO/wG8+/OMZLwTo
/RjX373RfYlonMx9N/VYOiHpmmOn2//dIBhfesL5dE0+P9xoVK0EV4ZPtKgI0rDE
BFBCCt7P49i86XM5oNXF5K9lHc6iFHMo4KHjS+YhoCcWfmuMA5KvZ81+hu+wORpO
RDvB1G9SVZLMTskb1rvYYf8r0Bbd6+wfxKCMsZKpg7+TlVkw8EpeIY/Gzhy7YgvV
UF/H8otI2rb6boacDLZHmUMSDfeYsxniU3WRyD+DafLf/pvzyki9I7YdPNdqb4/E
TCyLI24HzqiYraoRcabJr0LheZjdrmhDa0JC9JakEnlTn/+RlyopMkCq5RQMqkwo
UdgBCCxxsvBth2pTVaLf/Mb1fOz98mKhX5la/s2+6HbEfbDT3sh/G7h4HtYuH/Ey
ycBVkk5B1fzUO7L4SMC7nblhDy+GcA2H0DuchJQDZ5zKelO2XXv3nSaQXEVWpfV0
GvFVAXxLY6P1mAY1NZSR16IsSw3xKFqadajR4matqr0kW1Vke8F4zYqyTtrCUYC5
gBFIgFhVTcHPEBV/GJ9pss2X9k3qQV/lxExmzXHgZOJYhAVWnYM7+PPW24S09qXj
m8Ynl4iCAyvRUCeKJWuO+Fdf7pW9U83ENHMeqCivz770ls1tDMs2Lrok0Btf4ryn
UTBeN002D7Df2OpQ8kA0n3uaK9Ue7egvQGjc8cKRHSOF7DRNiKMRSGgnydBF2q/6
piZ4NNrMqky9SKeNUXnsmUm9D20BW3NClEuALvM/JMBVp7RTFrBoj/U7NJYH/upz
DqiwKNjKtWEmmL+3mG1w1dR+j2Z5dOhBLFK/SjrmMyEg0V4RPp7dVJKRd0Y2iHKO
9iciqhrfLVwyfTLcVkMHquCmijxfik0We5p/pTdvZgjPiTOZuenpq4yi+egBLWNK
JGhmLwOo+ulieW6Zc22HLyv08MLafzJ6nnDJKvP8TqS1LCGZUxMb8MXnIOwtnmfP
934i1UddtT5sSGKcV0XyMHUJUdf+M9i8JhOzS1iPeNvhiuWUb1F0FFZUiPYJ2LuW
immFJTjXtgX+pJfoG8/a7KD2NWspgS1rHfMu+sfuJ+C89JntLCc7NOzU/8v7CSfj
T6Fg/nRQ6a9z0USoGgyVSbn0X780K43e5CxR2gkHlZUGfAyWbV4t8a46XiKXvIPd
PPkIFSZClBPUUV2n+LyJHk76P6nrKEIOEV5o9D5wM4MwImvfQYNiUWEDeGuE4xkE
bWbvI0Bgm3Erj3eOD3llgZRbL2tuB95Y0bj87yDV3y87XrqA8Pb2G8lKku6EDDa5
Amche/vnQvkSPS3iF5fg83JgpAJCDNkuaEh91gzX1pqguwOgYke1mlapAECX8lgY
BcM3w1BCxU7AeSoYvdXVCxO99PmV5lJdhgdDZlJC/4PIiVJNn6ZVHg4o14eLXtTj
Y/8C4q+T3haK346p/Op6k98pdsz6Nj/oupdt1VlZHpJ+MDo9Qr/JvLCc90sulTPt
k3GLugwannk8iVCwoP1TzgU3uWVA+Z0O9ALMHv2wrn8Q9wnsy2wzb0W3C3FZRxlA
26Z1s6ktbwxeVru87E69uJPGUymfuU1mteYjVJSUa/4NYN+APjsX6FLgNtA5FKu3
ZNbobhWOV4vOsVfWEK2ymokrwtwdUBGcuhVcXkhV9Zupq4mjO4mlCcUTuTwavpzq
uUPtzYtxJwOSLmDHb+RtQd2G3TW9OJl7Gpnk7wyEnUnGcCOFAyWg1SEdTmFYnxjq
QVfScZxP2vgxhHZBrueCHU36HM1MaDlqsXaz54DkSXyn8CVglirYHxOkuHy1H/OX
WCDcuNHpLwm7ZU5F9T6Tuo25iJ5mrLjiBRyHwYCRBj0QPKdB1Y/XV80TtKK2Hzm6
NR5bz2f7siqeFebhyuxe9Js3RR/iHcNq7hRbo3RYBq/nRWeCwEtp1bQ+S6deQsfj
W1RFaIva8gA5I8hycnz9akxHIHx5egLOEwR8c2uywLMbXkzFlMu/a7Ue7MPAHoBG
/g92h0I77dnV8CkvysfciCUJUcb7yQQiYH/wT+IvQPr2nz2sQ+2Z1LEE6DXuE8p+
bars0+jkZZoL+peuA9wAjpf53HyZRbqISMEBpkMya5kHx9R7s+X3z4dQABud3wpw
bWdHxSbrd6em6+bKFIO/zZYSAA1FVfSh0JZKTitKDmG5nvVp3gVXrGbTV18X+W9x
CmzoN1axWTt8l6Q0EGyCExgrXZ1nS200UkUVfzJYNF5jasaEq320ggUpQHTrAfJ5
XfPmVw0P/g1I3UQMFrARXDMSRhhCaoqErC+nlUg7OBmLkBqf4SZdQ6VwttKK7wi4
mt8K9WpuLKF7EH4GRM1cM/rX3XtrXy8cHhEVh/IC1UH5/veV/ab8oMUXYSSjUIop
i65eJ5klwtqPxkiGgux/PLa3S7SZ2zYgrUHVBnFkUAykyA04igwTiq1sRWORVr1D
1f8t+ckVqHXhPBf2iJXYs2Y1aju5ntGiBm8FBs+4tkBi84BzS0XoTW7bXwHJg9vv
RDTPiHppl+fwTiaBLMz4bfnGh9d6NEvsYEjTdIpxz+pgdQ4/XPWAtTt4/Mx78/WY
DsaqXVxdJkJ0yYv3LW74HMudARzoiloeM8hPEv2kbiwxmucXBdrw2LCAWBqx2yzN
YF3gn7gFf8B1hYKWqG9S9FPIDp9Xg1IZCrblSJ5qI6Oq15HevYCR7Qcp5JvZdNmH
tebor3xkuW9wjLQ2ldkdWksbWXqMT/RUTvrAS9WwBg+wJ7+f9dof37IDFncEfeAL
bDM6u4S0kM5S8oEWzmdn8kyiarJrxVqnwOa5uWsQeHD4jJoIPjQBYlzvE9EQV/7E
Embs11uPPhoLZo+7hmi6inRM3U/ci1RIxrxJMly8JORzvpTGDA/kLxkTAZBjlRKx
YXihN/G0YAFn2DIrIZjNYy2ZFuOqW3bX1XLTYtVxg8WIzh7cen5avg5mRfLMyVgO
R3JZ+PWQvz7rAJS0k5RXYvkw1KZx8an0/Ns9dzjGzCtBiO/QLwKxnANU+/FbvpKh
XEYl+5FU76twqaTkZGdIPGVbtmxVgxWbJXYmYDFqydVvs1GaDvnfjFdMzSQ1xtP3
rGuyYc2ck49jLo7aAkXPd89zNjjI8uZW3hhWi6rJvPgKEwhha8/VQqeTS4ZgtSL4
p5mAQB7YY7iiA3I5VtRseoDZPWrOqNVtlphySJ9EahN7S7TjjRBRZQM0yuiclQ9K
h3NW3LiSQvjPOKxo7vA/okmML7D6yxsDVqc7TkcJSwpf13ohUu0pDnUCUkaWg70E
5L0uXB3AY57SMzWGTo3mdV/tYcTmwXSIEYRsB+jh+sF87HJlqSCzOXr3kGV27UuP
FMt+FSzFIfoT/vLe+lT55azxVqZP1PKOcqZUocR7IXKIZJ7hD52NASOiSnnIR4lE
kcZ1SG1wSfYIjyMAddGMaI46g8rOuD/qI099iZ4FIFb8WEGrAtNnzhUlSpx50YSl
F6+y19vMe+EANmn+SDe07uLJp/60r9gjQdJNYqCkgJDrc148Kv/nzXxcJp0rF5En
V50czfV7KUmPXWGDs3nhnTPo+whQ6Ftz4NzISZxxAZOQE8Tgvl+o8eD4ccqMBtkI
DD/Lz8/Ywl3CHhB9HtW+CehBM5/XQRaktEfgBPAWr2NTSMEIgdo/2s0/uRFZw0A3
9Fgeif9O/RrVmnascirc9mYvSNj76y4obCl/Vd0AcXhHt+4W59t9nTUQwrbV8+Cj
vjzeDHx0ZywSBb/Grcad6+PQo/5Kr2efEdgWieRiK6O4/DiKP1/zwKScfkY6j9HG
nKh9lvyfFcigioXtJIKNLmB3XWx8sfIguxq/CVY5mSaDqp6AL/QFPuqOuNcTHiEi
GrZCPheU3ADsSaWYO3jDApGcUJ+7c+Jv343b62lWy8fByDxGKqSmsG8vSG4a6+ZP
FCy+4DFLYPEFF7B/VkRWOhQGJBQBM1d6SAwjryY/VfDb+UpF/Jpbgu8fotX9U+MJ
Y6vzRXuhsEx/EcRPASxprHb1VZAtE64U6wxp2uhSirmXw5G+Fte73UsMoib8BovC
tGbYjrxOv2OrqLhOlDqKXYgpzBNLfFOYwQRm3n8iTOLzI2WPxN7nPabwJ5L2FGeT
nTMKFt4SibPWsV9bMgBjYrwK+7DBAtrmqCvVzXCBD3DzS1KvTs/o+ijtDA0wGNGW
5kS8IEbNI8d324xdcZn+VA7Ek6FoL7Ly6QDjmb7X6xiQJ7le0CLTG5I6vRWKJPZo
IpUFvONC7Y6gfnMJDzcKZtCZprR5mDCGYGQI16TioKVEDszn7h4tYOB9I/Tma7pS
BzSBXMyZSDeCuRHZ9G8MxroAKNzC4as5SrDKXESzkIrYr2xNNRYzM9wIzX0TCmKX
yXrzoJPo8hqFbmZdGY0FJT2YkNBbup8wFJC+n7Eb5R9H0Tx1NwZgKJ1WFKMKUlr+
5d39GBNdLSMQhPdoe/nFF0Pb3tBIjXbG+Yyg2lXp67YIQAXIyc43F0VG5tGFcn8w
YS7jpxjjDdjRbWxDkmSbPKFgiGV7/MmTgdT+v6dx8q/MMh3HLSS93LFKn3PSOrh9
Sdl4n6kVzEztfG9OAxejC0e7qYPpsmrEXU1WOVDn/qwpQ2uvBYcrPvOGI6f0aP4U
whMW8NYjX2YQ9hQ/yIFd43kl3t6YlJV9Qxp8uxP2HZtp/mEL4IhK/G6LfCTkLZEZ
41B4XKffox0gk85y6iRKP/nVaOw3CnC4UZwrqyzrgTzr8thJUHiuE8r7gSOC3aRK
is61ZcR17FzdPMhuTy5PjC0VqgmEGJL3GrqKZTZCiNUpHII2T0KIp82KqYuH6V17
4mtpzesxylQ1KBp1inhkvd82MM+XgrruhX/P04Np3zqlP3abuObUi85dZNPpmQ0e
+9zFnWXGgZKUNIhabrQ/RjzL9sEXD6DveZ3ffc8x0t7KrTD3EXeC2W9ejbi/tCIa
aNQwXOZK/5lUh6ekQQc7muNmUmAz8rIjiyeFOr927R9fjFAxyazr2IH896BRjK8N
pUAurRNKddSOTs2+gK00VAFFv44Phx+idU/k54psIPcmQwPiDt23+etp1qmWjoKu
0WaeU0W4VXYIdiSXKAlikv9shehiwPFdi8pn+Ky1J4Dm7mf2+eLG0RQHBiN6ZF1H
G3eD7jpCqG8oWul+pi2LQq6oxFWRQIa2fbiBwUPJ3Mkw2D9xuQfK5PmwOIGEeoS+
/+sSzDs5HyQ3/sfxjwJZyOUNHFbir8OQNIzBg/U8mfuDog8UWQ5XYmB9R4RDvAVb
v6UajFcz4Fa77JNf4RGLyDdVOGgunT2jQrzIiky6nCeh7lujQM8rFe+YbEk/r/u/
KG94D0ZPmkXROw250X9mgYgrQFypIi+9aYWKjAR/sQWpRiHjVsObUJtb0AGvCFYW
ski7478IG8E4eeezh0OWcRd0zn6PcHvfnWLqw9jCXSk9jjwOQnh6H4HXb1L3uKmy
VuwfKDh/KY82tP7N1RPBfVn0STGhqIVA9B/b+82dZV40JMQ8RvzsDC/X8mBN9588
uWCnuZSAUlFd3zAVdh7eFkQRS4VntTr5OB6PK4kN5wVYIut01jDFzUKj6EY6nzOy
WSWHynZasIaRHniUFBwhfxhCxL+Ijugoo4tkXr/KxkieWGpk9SaEK3pkVD8HeefS
Kn1F2N3gX1xzMbQ5efnbY7hL01BH07OhuGd3fP9f8vr0l3k80sBZqjnG6RvKMX5F
/uJPNadFA7GAWaaU7aHZU2v0QPhZOZ/t0m4naZWBD/u9e1Yw2uUl9OKopg8LeSqF
gZ3Q68WDQY6sERYXPr16Y3Q7EdKtfDIMJ6fCDe/s6Yn4SsszoIwkhQN8lKH43ECl
d0KWkidEXevIqI1ZuDFX7280tc/hTYboUTLLqJ4Vg14K0P/qVSvOgPjjH1hWVLJd
samm3zXa9+2j2uhVMoarYtYHCDhGjE492ph8nCZ3e4YwHIrjAjvr1/KqS0S36Gjm
aFDiExzBdZ2FlJL8Hd5lYx7HbgbnezUBbyy8xvMBwcj75b6x2Sx/Lkhrj1Z6/AxJ
JPf7oj++mTjv12KvTKauXuIi7QeUxWCz5910GilbqYpyBhGiB0Wbuh8klBPyrKU+
CpgBETzy6sypoN+vkSdJw18FjYuPf8nfnFAXc2Wswf16oWmH8U5KS8ZvFQ0e/Sid
ahT2gO/4qpQwbi1TqujRlIOJJal6Hcj+aeWMrz0IuDTy5L9TsXidF5sU9tELl8T9
+8GX4FLou5T9aOoTf/TOPSdCSkryWcI3NtUJYEJuhgXibGyj8sCfrW9L41k5vh7c
rMbX8ngK49EGo8EAIO/0x9OpGskE/LMEF6wMmOLNMQa/PANgv/1G1hg9SnoHGMK+
EeL8Q6tLC2wSYvpcLHcma9RD+kN7PgrijvE1u1cKM0rLSXwya2+j+saU+N9aP5/A
8G/hRktjJkoQxkScdJ8xB+n9LXCjGh+WVNgu3BQ5tcy3KeA44xQdY+eKXtlJDBoX
8xMRDDaV4uVXhdemBGEOqKXLd0ObScAIR6frvJsrsNrDbAzb2CzBy0mMgvsL3cZf
dOVqa/L66h0JkGeboHxfRri8T60XdroMLzTv8xLmCc4kNzSbijtnHiq2GuUvLS1M
qL63Xbo7EVBuf5JJnP3wsUvpyXybW07UoKTtO0FxKMTyATzqx1NjmOS1CvKbwJGt
Y84muP9k5c7iqG9DhNztbydQ83xSk+3F1094G1pGpdGPabqMkyTqUC/hXut4WUhv
42v5tVUJym7reGgaNJ7IOIDFEXvjJYZBivSvMJiglqsjA2cwc2jq0qHOBu/Z3ewx
qKO/5uvovb4NAm3Xs2h7TwCpVdcYRSwTCJAGEtJ298WU+d8oHGcvAEQXV89ztXiG
/nB0UKNZXc4r7L+Gz+27/SAOEhT7jzVkk6QD2mOyguHoPnZ47kzS9UgWqqHKsq+b
U2H2I8E0RYvLNQOCDj671qq3NDNa4WB12d5NKZpatXmZaADWBxz+PUK4z2lI7fOf
D3REZe0WLAyJha238ZiH3b5NwQv6Hc8v6kAV3MGGOoJNu9bBmEC9BfDrhrzX7XCZ
EWPr7VUWz5aBh+Y0eE9n1WQhBcYlFcr3g4WEO7KZey9BG6vyxe9jJ9gN8fJJ/5px
Bb8bIy/Ye4br+FxGy5KKqkTHZn4vR39CthwmYo+EvVv3ZnRNQrpoLS040VHlsSr6
yLbmo54HkgjzSzx2LPWiI+YRlEMIo0y7bT6iAl1yd2J9Us0RY9nc01W3v5J3xM01
R6+HEgvMhIxARgdbBKLexpAOIAj5Bqm8RuGN5nskBSknKjk2l/GdHsiN9uoWibk9
9e/vK/CTEEf1t2xawRpsi4CHq6RHxWum28aqBwUeRCqtJFvmVwtrglDAwUxdAwWv
slrzMfqucqHvyAS0gGscQTt9SIFufUzFBWQXL8IGSjEjEOSffTjScEHJ3cDdl6XJ
123dEtZSFJG8UCHoE/9Y8ahVCDMq2eQdM43UvyepOh6vTjtWW9EphT3D4oqohKlK
348V4hNWGD1Q7bUXOZqMrdbdqNirVsDpOd1uzOLPvnfwgxidcf9yKhTu3fRjiPyo
HBZUrgRE+cqAvwlHbzBCAc7nIYuSLqnRMF9jS92fsfciVLLch8CxWzdGfQez+fzd
D6JLNJAureIY7/fX4K1BqjSvVJjVeEuKW8ZtFbPOdY+p9Ms80k2MGzrU/zz909IP
9hqAWWPzxdQyn/ltEWthrv5vH17lAnkqSfrMYySAuwbmuNrPAhFV2hV2v7CgPozR
UJ4kAk4nk2gOftwE1Jo0gRkXfKrMWlyqsRkJFCF2D67XyzYBtVcnNC+XftqwhKB6
WDp+Ae0gpVVmj2g3TZj2thQilLkblVo55RBoApTyFzlko8xWa63HTAhMZ734CAvs
tZSv/9LoqoVNO+WzdOou5qvsfgsU3Jh807cWEknjGHC4L/0j7C+bJlkbC7wkcbcM
ZCteh7WBcY4dR+sEGguYYbLwFR/wd4scjcqs226PYVLajOUie+fcZwHSR3pJovwm
4RcHLpSW+Hqtspkn0EPfotje9n0ZC6qG/L5HbZh6CD6a0ty/ONJkyya9lJ3jCUNW
zJr9VVY9xKtalyu2uZRV7F2FwPH39cBBxgh+0ITguLuQyhEjAQEQZ4+CNLCu6I2o
FX6PnkboJYsqR5f99L+wJJCma80QegwY0aTpIhU7r1NhQV3ZdRpRR6icnwJoJ8p3
IXrOHOPl8qk31F2c3ZL8hMcMtBPfbpz+8v00creDKS8lXZXCFBYcZ2xzeBpFfoD6
gInpujiVvhwxmqyU38mHwhSvTdWgW91zztJW/ZeEkRZkmW1hhpO+fpE6xZw1HLgx
kYn16OgpjZg9FQp/WA5xgoangtPYpehFfqntLmB7dWBSkMaMUsIdD22qF+hLzyQf
Hm5A4z9zgb+XwbuTRgNYX/7t4poEYBt4+bLQ8m4NLy/JKGni1emdk4wljD44f3N4
Xz54/0/Dl61V6OfFeV6OO5RLtpQrK5NOfUX8cjIKcrguPzrs32SOqapzgh0crOM7
Ygnr6yw+oi+e/ucSFEuA0+CqGn4cwwxHVa1ADEB2xFJrOHzKSmKyKlWDoNMS0M1q
LOLF6PlsDVNvuPq57aqh8sdj44ut047QfsH9WxCAh2Gj4wlDzcvkaHLA7XF3gyeU
hPkDIi9grDJr/9Da2uBoU420EGB0tAs+JXbfSntOIPqZHOXU75ab9n+GDJI8jNGn
Qc5a3kkSNLOJzFn6hcq6ghrt84j62R9a9j4FkWucOXnPERKnyZo4TyPEHJH5wxRf
G2lWJtuE/xdsCWFXpvFJKkC5VXq/WI4JlwohUG39okLxXuI/LhWNoE4p78gElgfz
8cFSboOqZx3E9SncxsP54SXQpsiPoSXFHv0T5gDQD1+im+HMP6cpkp6mzqv4tTsy
bxbyrpbyLsTMlIiUkeHGX8i8O0mUrAJHyzfDbDqJVoEKJ0hwtP7os8FL5KYSMI7u
374rXvbWAmXUNjMzBcWkRS7bw7hu4Ua+IOZH7OxvfWCW9K9udfPZpxpoBHKvTSTe
A6sSooL/vi4QKG00Y0EBeutXOhPPAVBeTj7SZHjmlBMHm73NXZ6uhBnRfltn6KlF
h+x0eC9YnqadpeNhCvonRfUdpUjbWXJcI/8pFoT97eNXsjohx7s0lgag/8hVus2f
6BaVi0Z3i3EVmFG1aFPeQ9xRi2JtyMVSWKzRA3RpJ3kDfXK/U8e3KTmMh8SA+xT7
NXUmS+af50gjG/VX7VblbRz+AqPF/vdPnZy2nBMJuq6+wg8to9CtswcMvN4Q7SIz
Aab8VPg37zC+7y43TaZ4Sfz1HwckLQOB/wT298gb/ekKq1JD6nhoEgoZ3wb/SaDy
ticE3MF0WGwoyyPsp6SaHbnErQyNScfQTf6XiZvMhZj9UCxz8rXSBZKSnjwGw4ez
AcLfcyB0LMGQUux6s1pbLQncsDP8fbU1OiyX6eEddPMn2eZ02YZRtzpAyCqil3kI
xYl52oimBN/zzjfh2RQRhutlktUpAs8lXkSxEXrTQxWeo0DdK6843qgfQ3k9n1ME
1goWb8LGXAkvxePJDAYk+1ygWarqUZxBvnKIL6RLUEnF1sRS7+uNV2wRm0aUw57u
KhoF5aZDVZiN4WV10PNxseqf/iB9IUhm3J9uQ6CNt6msrQ2sjOhHBknIWExRw4T9
GnRXAq4fdanRxqMePQ5Ea4lxZ2ADqxWt+88w46UqTVCBJe1QX0lUYpbNPoxaeuMs
MSXac/NtcGHhlox5NAAi6lGSktYCU9Bhv2Wa1iyFBPF81lFnQLIBkJI5qduTLvR5
rc/JKi4GpQUwDOXU1qkhpoBzG0fvMd8f4Cxth9zJuSoqn7evmtLGYX58B4fX8ybG
8Es8ZG/mALwJdxqmOepiPJqoIxjOpearXp/O/MIuNBKEv505AtvcO1BaHn3TIthv
jbAS+wRei1xqp8OJ0OApy2Qdykr73ZsF/m1M3sQpjghf+UDJh1clVp6qc6Jm+AWv
FsW3tR0jVZUkG4xxnfMSQCAvhxjh9ZOmJRoSFeFYIeooHmf0MVMd9D7A7dZs78pR
DIELvH3HOt8aktv17T0h8TbqE1YVeGJDemPKm+w8plEc52IbG9ym8EZ8dc1Jc8ac
Th7LsWbzX75NW3c5Rynk0HHF2ZHpnQ0vb7a/LEmMjhLjeP4V2H/ZZZKP7cTk5BB/
H79H/tB3BsTPSc18OlSb4nrKrbSOydQLUybWIBfUZ+Kkb8zpFFWWAElN7S+Vk0C3
dOfomPkrkpqvPymRTc4Eb4FbfbR7xzOaj/1Zbvb+QP4guTHojFw+Nu5URurVPvbT
5kpLErfCIEZh3Lq3mQDZpfaDV6F22CDYoNgcZAfh/LxnmXS2xHLSeTWXDHnJKGVU
LFIsQ0KQNnumTMmf5j1hOXLZOtmBI8RR5Iwu1Xo15ThvXMGLnD4faTf+l7NzdAVS
D2F7mA2jjuCELXiz/Kpaa9htxz+hrMRjQNDJGu3+AjQ5/S9rnNhvWiPRd90GxIPq
nvonLriQBnFSHDHjmslQ9WKHK526EHB58hsA7pkIG/XaUeX/Ss6KbnjxKOyunySP
C/EZmKy1TahfGjmzh7BDy9ZrDT0jX8d7ivs2i7dcMXDum0bzKErWYO1dvNvrz786
uu8/TCJU/BABph7t+2u3yv0FlBmpBk+TCj+O4KsBB3t4hhSzlITSKgY+98r2SkF/
JlU82ZrlrCDHXRFPLzO8e9IqjbOl06fk5UXJNtfdqb8OfecDRhEH5F0WNnWlNx9o
TgtDQGhLAXR6j615p6YhYGGNdyT7UmO680k547A1X3cbzE+n7o3QTczRW2tkq10X
XLcqakaaj3eg1oDoJbIU2eOT3KUIXbfOgKVtrpOtF92++KhvMOirI2BgZ2VHn/hF
appDWVG1xKJZJlrrRNorNRPaAYv1nSkKS06zNt2auyvA47DWp2Zr7W6H9Xs/84QC
VvhNg7ZNsCmzI3YWclZtBsvMuf2HuLde8UDlDUyLpy96j+fzteqEAWYKHTu+97mU
Y6n3/OteLYBskTR2BFp3vMoM6FSQW7zmiYWFhXOaz2jOB1fjJvZ1Egcezzw3KrzO
V6iHsHY3nlRIBfAKo8KSANX7ve6mdiMyJVE2qRXXj8ehMzJ6yheTVXNwaw8WoXX9
Po+6lh71YBI9eJafyf7OWmiJT7H/vRsA/s/ToJX3roUyWA6c9jnLiehNPJSPOGon
hTX5TglFK3rkW0ttC/SvivT2G2KBrEVJo/MRHX7uJqJmAJqQRoj7DHPMjSkLonFC
pF76gmagvhk9rkKeFf5yrb9vJiXX8jKzl6wAoGszMnayWvTZus0FQuwLsoj3xPSB
I2ZRY4Ok9xGmbN6YTgPKVEPEmcV5ZDVPrL85WymvoDK0A9V3eGSj3y/Plf2uW6IJ
T0GWj/gr9Rx8Vewj5x5O5ZWrF7sYh+IRVVMr+GLR2oMjp9YqLpYqEqGStqpA2bq5
UabpPkOIoWyZEqnYPKvx9BRALBQ60ODMZOjnnuLCMtfXEO/MDm9qH73JeHcYTPb/
2lNAUyfodXGytjcaH8fRb1m/Xr1wE8SOPRoce8Cf0AS0ZyulNtOq/grY5PnyVtDM
hAM54libLe2zYiixRTCITuXODCpv6+iHRZnvhYlifMan+jZ0YQSPJtb8RCqzsZze
NGIObyNaojR5xYDMPgtgBbERQu+jNDXzxdeI5ExVZelvrfDpIZV3cIcB6bzYPPlJ
1BQEcbD6dV5bJUw3wprfb74pRDEj/XplqpKkoezXOg8VlaVixGQ4UWzvkiFumSkp
kN3eC29Rd7o5UQhPBkBMxeCBwHYaA6Zae/oU5kKV4PVo7471m95D0tnrCe1hxICq
+9AFxrmR/shcBSt/iA+SWN9XSIAd3W0+9M1OSpanJT6NUcPWk90OlArOJEXdhDFF
5Fen2mK4eFft9zMtSKIgBnrFywF6XsEfxVrSiYZQMSreX+T3is8ralGcE4A1xDmd
ua2ihuHMJGaBNAt0CN901NKR5CTA8h3KJ0LQhajjnDK9Tf/1El/cZQX0X/iqf9m8
XhQSB4vh+g8KJP+PaPGDCZixjuGXYMRwHalTmVBw2TNDk8UKilvGNQmwO6Y3OSrn
O9WBgLYEhJ0oqTomV8dyOL+dHl2iBTzX2ytoH/bODAco/YPupNFTfXA/kcS6viYz
5IEJtcn+R75os6oAAmwhpafa5dIpKNSBUPbHMtSPBW//5v4jVis8CRPtL/qKiAdN
rFdAcFVIrZDRJfCjciUVZifsD+R7QqCH05RCmIDhnW42w8ueIhywRHWC95Xw9RFn
YzdsJMEtOCecuN9uQf1/CVAzmu2fiDempYl4fhbw5BEFrP5M6iAiv6VtcoY8GLEn
+l94vBKG8OoYuBbC8X9DjzFLeIWvk5dFtn2AIGMFD1u74WeeSgWNTfLKujDmz+MU
s19tvPkTRmQBAt+TtJkDUOSR59lCdsvqia3lgT/O8362QNneipxB6BscUIs5FLi+
ZUbLwqsi43VIu6/rzDBq+qTQMxXcCMqyJYb7uU0dlSq1xneXdd5n1mk3ccwwuM1B
5Ls9UTjMuuSBb7wv9+6qNBdsf5zkwyDoy2OjfeWrUQPsccnzWTnKj67m1tz8iySA
zxbplANC9+47ZFvizzN4lcKcvbegH3kOJb0kpBzplmhjhfDl2u/cBL1sHmeYmrag
3DzM8rC7ZZ3vQMlt7682OD84TBNkKhvpkYSAyie42pcv6f6Fa32mcU9N1GeCRTEx
jJ6QeYJjII0H83zPCAn/WtnFmgn93rO7tTj6bybB0YRf33pQ7AF1uQ6H2EEdnBbX
ZPDr6GG3II89WTPf3LObOoee0alWw7BKVInnzBjhPY2GE7lV5/WW4PpzS1j3gJHP
KuUfYPTH5B3FkT8wAZAtD7Rx1AA5DSi0/oypNG+hknxfRoynKQHXD9G4O8H+E4qA
M/GbMMI3EZXCTLcRtgMlrbfAyFOj/JziBU+gWi2pTI7uM+qEiHqjMxufMmXvMl22
v4MomVNk6eG732p3OaN0qlDPAPYqVBokHa+CZd0bz0yTF30cPD2uBAhLEnW6UHG2
OMETVn67Aq8XUK5OtCj313QUJV8OIeiNngRDRijIDPG3WgDaszM+pzM7wHiXrZu7
n+7SwWu+T6ixtc3Pu04jl/4szgoCzlHAZnZX6EKfKsqAzz2lBVvZuPEIKdr4h9Ov
JVYOW+9jS/e8GizzuUPg39C5GwzuuljO0QXyBeTPlessMtoWVJzze31Dyh2sEbXH
9Q5dAfLDXINK7362+aI4AdCsQnk62kcgQoTEpbfXJFhvAyKZjCOZO4+/LZVH7uQy
K/BH2FUUoyni0xtk1HejXVAA2l/mkTdaQqy4MM2tSymh3qg7zv9beiyNaDDnNb5S
cZ0mD25OzmaaiON2bgINlqSxwfBatsrL7wEkzkep0wU/ZmuekxVviIPysrGdTmZv
7QXrwl+NEKqoNzVol+y9NOl/qFLN2pSKmTyh3fgDgM9cARjyXYJwwESl2NsaU6Fc
InTh1Gc6eFgzFQjEPwSmHGyiNM/y7F3akGE447lDQirMi0pnAqXFa53/+G1NKYl1
NRbuQdh4Wam20uQxuNoXggSq5oOgfD+VROdq5mfZqrHRICU2mpo78rJ88UPLPPrp
xwld8z9r9Kv1s9a9QyaXs08iGSvYBr8IG8c7Tv6W53xBgyXUeIjxPkLy3OFjFimV
lD+kgt59DBhajC+AxmUmq7MF7QVqRqjefxWrEvV166aXMLxTtyDTafYdFqNRBhUT
PByPNsNBZOYKqe3U2qom/fR2MdERjbVqzoSbw7u7SaxNa1TPJWH8OdIQbN2S3wz0
nfSBY+DYYMb8zlzBNAgaAG3AVF+d3cFA2iJjcxAFeblgR8SqEUetx6Hgx+Gxbwu3
k0M+M71MuZ2vmeift6h7Q5XTdFIwE20tlBdFTVFdWhezCkoajSnb0uwHNyDekwNN
fpMjRoktNcyzgUP6qY5tWvldq/gIAoRXRETv91QqXZDo9jlGdJ60aobJtvoXl576
XS2Znr4bcg9ydnV20XvjLd0Y0BpNW0zE8lQlett2F7Co2Rjt7kJoNleMbHoQatro
mjdeX/Nn+OxYAYg0rTNFfDrN20m+ogDdRUFvE4xzcBUDQYO0kaf+frUQjMO43tbb
0y6pBxMbCFI6T9OyHE5FMORfOPzvBDa1dtq4lquS9P4gOvIkYAyDjH+J+NjMDIjS
w8cQr7eCo9T9Eel5RXqQ+Bqz90+lbknYSb3p6mjvMXqv2J1viSATRHEM+kmtN7hH
Ksfofh9RKQrHSlBlVN3wVorn5HJcLMUDyVH6/x78YdJYmMYOMtlu1HbtKyhMwVIn
kQCFFhLqxFnSU5sWegs9TjXDOmO2fj5uBlHGYF4VnMQe0MPDKqYOzSshTFaBrJ6w
VtRRZ4wwxyb+068Zl8nst3xCr4KFrGraW3pVyvQL61GmHXvgn7Oa2y5evk5+qrBs
1t3SWquty4e3sf9NjDVmltVThBbYVyVUNMxmdhyhExFgB6rVF6vSwJ1xAyLOk2e7
xixxE46Zzo1G349wpwgBJTWoT4/KTpZ7iYs2ehNPFKLp9vIxxlRjiu+r7jQW4la8
yA2hWV/SCFXN409l12hjco3er+G5MyXIjVVSv6Cg8osvKVFYpyDX66Db+0xjJzwX
iwLdWq4bYYWkJv5PwOkSyG6H291YH66cW48LSto0L8GnRnX2y28JiUwIlYnfryEm
EQFdnOl0UTp3Qp/e1yhfJqzV3xi58OSsG0HRVv/HADOSzg6ncotfLHi7RaISDH0P
4ewX0QAOl9F+jqLr54/94vaBVC+xKDKqoKw5m1EAz4Cfu17KVkRtTCPEiFD/Mijs
nxmiv08rNUThG3JmTy6Dha4xLVMP0MWEP/lrbUdjrsvifoMZeHJXnyWlWAh9qqen
xJ9ixjxVn7X2ySxQh98UadUPAmdB9t7ZB9KayK4veJ6AxihbLkGCIc51EQv2PNcU
jCPVobgC8Uh+/OuJTYhXem5Q7TfuewXkxem88e9m9/zOzQaI4WcGZ03JFnFW/Dxy
CihJqveCcI8YidK3JpZGAyB+/7Gv74yodVwuLtW3ha0DesJ5O1GQlbmeTREs5Hxj
/v5xPAIU/4VDmML6sYdlJLyfaU3zwdD6N4Den3l1kVKFqV3697ksd0RnlGTFgB1Y
WbFf8dfVzSTqKx5uoofVEXB51yKILEnVmICc3MKIYoiL+ttl9AlcByJ2zpNM3+u3
FzvbJ7/UHe5CzjAT6JbwvaQC4ZrPdUFYhoUVMQANaEDPR9nTNVR9/FTsz/HZTtKZ
Fc5iUVYHPiAglQu3Z3OZeTaV57prVa58q1KupSTg8cnPnhcNFNBhdjErogXw97y/
6/lz1v50W6lyUscqlQVfHFVaHG4h8vXJIkGoFVvQXf75SO0I5DhMNy5sSjfmAsCy
bONpbJuGL7HFuIyrpDYc/BXCpB+bhnsnoNr3BtnwWDFjZ4TSCypsAVOZDS08hpga
YXTBtIByH1no3GiJNvpDlaAdrTuBzndmLbSLukAp0PKGb7QUzegl4e9fRO13+jS1
7wSI2OviH2lBFNhHkQekU+yt1FVEcLx6SQd+QiSOiDeZmaCoaSyXLInbNJRRkj//
4t4K9Rlyei+zP8o0SdLiks9+LFixXAePhe3eDsd1TImjZnxkG7yGiQv145Fl0DII
EsSzcJUHzBnKbFnusUDx0Z/+vBmXxKQuluxYkZ+kPl0IBh9EFIpDVbRGtJWhrQli
9aNV+PXTvUvfvKfD7iJ5o1BqEcZeO+8dz7MCXQYBiSg3wiYDGMtnVIwzkwWDOkFM
A5vHC2I4SYwblE1KFiqIvKzPRoFLCRPn06RgAPSvTR0z7mdEjbRrMua3WFahm5Ot
RPmaYDSY5xra9/J0azJzChOYoauGUlV1CAqLO/9KX/9c2Oy4b0STb2ZEvBV6E7Mo
thN5Gqs0q/CVIxY7N+m/stILegl65nHkW+eyj+gUy/dbhA74gVxz/w2YBy989gTq
Y6JyMKApFQzxP47ckBaZEePoobNhX7tR6CN0andTHYtAK6FKBIUpmfjEFibCSU1U
vu+lLiFknj7Lx4BHvPodqcOogSNae4aTL4VcQ4SNctTKAYoPXF1AL6EBfybBjG8+
HT7dCREj3frfzKJsPLZnNZgkCLafuo9OCmssof+bEvxMkNMWo2M/Ny9+ytaJ8cPZ
ayGAgMp4PhGBV98In6kSE4rUqT649oSTq3P3MvaO4Tl/w85otyf450a964OkpBqI
itnqCD2Z5L96wP4LIg+SJ83GVijE0lkLTOjMJmInhqSbR7fSze0YLa8d+gRxyoTi
yBlRG08ftv4YlHnDP1E4WpX5rL20mc/sbTQC6hSbdysd+RiyDoeWHUJKhad1vOa2
gake3HzWJeKBV1NQCUN+7iVEv9ftD/nohACDEweB7yfIFt88YnoGFL1G+rds9cF8
l1uSizIIl1ES9AX9SAi5OsQYgmrVCGRweeIs4BkQ+R2pWpufkzhU5zY0yTpXkLBw
a0TKIYTxPHq6Rgb4G/JVdS9aNmWS0extdtkkYa3VUyS9gxSlwaUxlWAzfjkmBl0+
q2asdIhdXkepUkNDnU0Qp62pAdFHV3e7SAeBdkG73Rc31nlG0YoY/8Ie4yaUCsHS
8oiNgn+BmhbGCq4qe0EMpYu9GDj75vN0yRttQ4KdGgTruP0Sy7Y9BHVlu4teFNyM
gxCa9Qn6MfpE85XAawJS8KIyLi7QE/eeZBuABwhp2onUm4OUovJNwcI3OfSQPfoF
QjpiHwrZmBD2eJFLVyjOyQ5MP/2e9rxOZpGnNk48nNxnSSKFSaBiOF5uAA8QhZEZ
lLTuQjwsHn9jC/P3VqzmsdC2ngdOZ68vgeCOSsGiPewmqvc6jtN6e/YoaT7FSEBg
5i0DqrZbYedCgHfavFVjqU9/3TXfuOf5Zvk4p00AkG/TpZn3EU2j5SKU7zuAbVea
/vsAH3M3cM222TL6G3ChcRHLgkP+MiNJH0VofvUgFuFNpsvwx7b5sP2dKC2v986c
jC6RQhZ1TzZFmqHQ8hqF0twhviw/53Gr8/5nLfvYsnI7LHdVynTip76sNzOuKaG1
nEs5QGQ+X9TsRdcbdGRrVRJG3dGAYY/gYyfacEqgHPlYTnbzcZpv+3daNYy3Kbjv
/aiUid4LVekbqh3NO+Ydb8f3u1sxN81TPCmOEYg2jza7A3F9kZbjlEE5hDqYTbos
Q0mMrDPE24l6GYMDGgSjpqmpWdwvifBoQqpTdrvPNOrzxcFmtMxo4MRag6znh1yS
6SHu8mbBh6mLTysPEMvmwMl6/Hbn0xVROmEIdjR7y0y9/530217fmVqnyV2gsB+b
ef4Tv51VV6Rk+trSPC6a5XW4ZhOnrn/aUxxbR2hIgbhFvm0KSuiLMizfbkgIB7zz
VIG1kfHzVWItztVOWuYmqqyQMTv3IhaxTyEy7CLfotby9GO17172FatdYbwIghXG
OQWv9+NBEyBE0SmF+FkYwwkxjIdiqyxzT/ciLzB59F+45HOmKZWvYPELNe3IBqlw
h7mqelbYplhCTsgGSpRLcwhW0stmWBnAYhS07oV6QqSqlRKpfVY807rFNX1XSjMy
vlAfN57+5UW2CYL8FyG+lxb1ajO6+MZFYbRnalBwafJ06CnRyauOL7+wJcUAKfwZ
KxLhZGxC5zH6SDgDxECUL/QjR3PDQ+j+1X5cwyAw3i+ZHJGeEUltywjLjnLOJgox
Cvo9oUsG8X7Hf8srpdcz8KM4UCrPHtKXgfAFZJKeoiKYSYEvK8+iLrksYaDv1uo9
Talpa2lqpn9Nqu8WqOXDL1TPaTJWFGnfSsMUwqptd+OXZ2IYUgt5SmPOBuXa4UXN
Srpjad6fpZet0mwGN8Tza91O9/Pkr4+AvxR0LxqwEx+ewME6ufKeN1eueHHNl0Cp
fNi8BSvL1MPsf8ifFdoVkwWCet//x47CkOgNmFCOddDZ/Jf9inQh8No0lKlKnusN
n21JxYY1aJIBNtroWLQcj1SCnkhQx8Zjzo/gsk6vZYupBsJq3xbuQQTbpTdP1m1o
8JPtITcC+ej6yUxItIJZbCwMz+/yoZ6k7O07I+2wpU5FFUKHLTUiKAlZiKMtxsWE
qlAuFr8bZZeD04sQuXivzDaCqjSpP22VG0UzvHDLn+Zz+zmhXDnRjCNAnKL79b/N
R7M5/acVQme4ZnsdR6dqo3ckRyO+0TxlG02nm1Z0NaHgQV9Q5c8Qtpvtn4P2DeA+
F14EnE6KiK8IPVdZjFSb6fRzAAXcpYUM+f2PYSKqSDXG+z0niUBLeg154mccyt1R
/v6hoj3jWAp8JoA0lFwXNhlxRDDnkpvyNUcz4kFhQ1HQYODrNQkLIoGDnxgrdQrG
Uxs0mmSzze3+m+wogGLPONvmp7O67ugwB7jX+M8WbplyRE1aIgXhBqTPzYjJpmhM
z+8di7zSJUhtzBcZ9jqG1NLVd+HneFzKZ9YIiPmQW5JRJztIYr31PGB4XvhCBr8S
ApyYl/ZH9iEv3bEq3Ohp0BqgB4u5GlXWDCES8UBBp1eaeAS5/jhWW3XClvesdHV8
6Jl5V9hifeZrpGSOe+F3kTaTPqGl4ws1TLsigExLBhL/t48sjolmKLvQUqBwNCF3
IM2GxKKvrPLYOOPOU3LygL0pQK3Irm/RPQadtm3nskFAqa2eJKWWW+ViVK/eqKmL
Tg5tXcv+QM/h2m56MHSWWUXMErPQsKCS9hCpw9umQnslkrUHKqmojalhlflNxMSx
VsH0UyMfwwESVYlEO/YQY3yXLaM6gMup/ClSNwdeZP+3ts/CcN/KBClIyB+l4PoT
zH/7ozLr8h8co17DK82sCve+bRurkFh0mqnPKYtWVKnZSCRpLp4eVFCNrltnytWA
T89LULyzF1rQl3tHtgfJhCcQFWkhb6UyEh4eU9Kofdjq0RKa48iPu/PIFzXCXBOz
S9o6DtyFnMQMTeYG/eRdV62KeLvOGhMLM3dLODDS9XCsm3ZQv+7Ol1HRbc7XIuUx
A7aDd1PHJ+9pwiiM72AXwf2NN0DR7pMnDeybwgl7MSBfGsz0eACTRkRPZjZ0pRdC
FvphHwSrqX9FjR+/5R2h+ryFs0dXPIMqzUgIHTi7Vnoj0t5DEVRffv2IdHjk4lyz
QurOj4fCpV43f7SNbl2vAR1+Ek1quQr9AJ/z8v/Oter6uBBa/rammilaPgasnr2P
u45DQTVstDACAZzo63YP+hCbl8FeTQAMZ0b1VG0CI1Jo48Rc+MFBNC5xk+jbrsT6
GHnbJJHGRjDMfHEH7if+GdCXGSzAeW/IT1eGjlNkz0DGOFAqnFLa/z5PzJ8erTOW
0eBVIWatmJCJK2k2Smo/banz35+/Jx2Bt5tAAs8Fb5bwvtXuQT23LSTIpqSrG/bD
LeN9yutRroqbmLrHIEMB8UIRZtGatFyxdMdgwd8yLUyZSM3Da5zyFMtI/q31+BdK
9tRJUEWiL2OolDmFyXgplReYzx39ovk06MkTbhM8QarqJPbDgO37/CSNMvtpwT1s
D+dUtG/aaqMk3RAJgwAE1Z6XSMfk/QzpF8tuL7Rp60Cq0P4zo/d0v2gKBrL4hEkS
oi0os5WXq2JwZtrPoajDo6hWiFXSMNi1G9allytSpjl3S59jH1qPpXNzZHVItza8
8mpzsoJSYetTKnoduoaa8VEN2XbMGdQmyJ+VAT7dwhtM2pzgzDuRg/dGtUsRXNSI
omcIyW9MvYW9Dd4qTP8n3vsa29Ry/5RixrucQkGaR4Ut+dtQlqBYUJDQ3RUHRv0k
6bk1Rj7NHdNckSnsi1HGTf+5AvH/ZedFOe/LavgBmbNKZWJHzFc7QBv0SQKhh2Wp
tL3rht8rlQbq9GtIkka32fGQz2MTUvHUjrB+HJywFssfw+Py1R34u80xq607KzLM
7alMQ7AXt2IxkxYyevonUK/1QlW5y3hVm866NswvZ8e7ZfSc1JccnglvudDgA4Ya
H/JRVos8OM5mLhQfL54rTFUVNx6v8iABeLjiL+IgrzKWnFPOkgQWSOsH/NpSKv0b
XRBAHbIvthyescVAx9hVdecN2av60lMym4lvfFOQhfiPmC01EiSxhjJsCkHY6GDb
BKcBNjpg3NmRPDKZdk1c3jDz4k7sutGpQbNT18gxwPTT9uqfH5SNdxsuOEdk+4+f
gnfl24sweyWBYG09Ymm6Y6j7+YOa0xdlmkFyodTBK1IimBje2EkFknjL7+GOM5Ky
ZoNfoTtVUgMGJkItl6NXbzP8kWnE4XZVFNkgLEuXFKvdAqOUrr22+FrkR8S/en0j
hg1yWG90p/cH3souHD6g4SnkbvM/ywHICPv8zC2nvnNIfpf36g+TeJY6QSq2k9uF
Qq6+rPbPN2alwyRRXeuymdwdJKa5Ge5QdRZdo0MaWnueFDxXihEsDZQXoSU90gNO
N//wNCfkZVHrvlBDwSwFQZDjhvvE+1Ve6wHmcSAu/x8z6afeUAqUe8/7KH9bx3UY
NVjtNv18a1S5MG4KOZWXPyrF7gF6vI3U5EkV7b17N/LnGdMcyERzUhGip7mP8rne
tn/iWMlcR94Z87X57ME61NojU+tfjngD7vgI3UWvJNBvuzSpMqwe4lL1oTuNIm/D
ob1u3X068416BGFrqNeTh1s2wAkuATEIabnFGy0k3jG5eh+f5L1Vb5+669QzGqu6
9e62OUSOb4O4drzMUc+1WxKiOAI2Z4CwPoVzl26ZlUZbHYNYipaT8HdG0Ti0hk1Y
pEXIJ/1NZgQ8iXWUq3f1ooXLJRijCSJC8Br96tBOrJvI5KapFoyydTBxKshSnQZ1
UtWmpL+KTZp2aWhv6EB/4nulG+AsqriAnY0INxPA+Vrx2woaz1+Y+zCFz3pnD2gz
qr5EQVEuQQr20D4Iilg4UcAYg+7YHsui3VK8Dhw59VkFYAgeAwmMgZdIbIJqp47+
PpXqkn813VORzugHda1+6tBklH/fcDKHyHSmtCGdHayendIn/DHyfXSyUc2ukHfP
qz4rVckPQMgs/Vm0Fwa6w6kPQeX22zvSHc2zfzi9PGE5RPNK3Dyz8Z26t1xjW8cY
mKaOeWX28rLmLO1hLQ3b/Nr8ZIhDz/aLZPNnxKhGFXMZ6T3TwCHtRoD2yxH/m8u+
G0G4pQqdV5XYN2LQvuERXwL33nA3KcrLzLAZEfS1sG21zuw+5pgntXxTxgf4hUIB
qjtXbjTD8W93X97BCvskkzddXgRZwmPSq/+gWP8gbYpVp0uo75az2/Wnt7gmXUDN
CcMP+056owrUJ/nvwb5RsLp6GdeY6Jw8ojYB99xhkGMimMFatSpYKmynLJz+OQjQ
+JFwsR/0CU7AkfXLSyTti1pV4/CVo40x+s0lL7qFucKBLQF9q7+oVnmXkxpry7r4
Wo2MmjmXrbTSkVo+e1V/5GrgvV6EQJYBv44m3STK2Qbml5nXcq1E+dqsF4R6OJgY
AbgAvB8K4k7CMeTxiwYh+WkBA7yRHajo/4WUQeBmsB118ulHcp/lQI4VeUbcMS5M
P1XT9dRByeofrBgfB6h9ft+/gKTqFn7tZc5pAlnbj4Xt9s8ARA+Ulgf7ADZ7/6g1
ufNN9UYMk5uLVN6nafaFD7nj1aqfmkEZGS3hShTNKooOKeRu7OxTbFImbBxlhoGh
QKVNF1itH3q7K5lV7Wpn9He4xwpRnz2qzRiYGkVw8z85Lmwjzxui4YI8ZrM2cbcq
9bDFSU2ZOZjhPuUd//KHarJjwe4e9aK35dIDF5vKNW01irTIz3owTtFYjK64Hrv5
MhrHhgWtffVnaCypDtNfcdkK5rZz3ee4t9vR7TkMTtsoycNoJhUDab8furxUJujs
3LwkC317LvyBFZcyuq9EFCFQpfcYLBHVxOqidoPBSC5eaKUR8YSQ6eyf++Sq58Qz
ZJb5tu8zese2BdH3DRYTocQrUe/S0Kk/SBQWOLIzVxrl0/kPccPLqtGGrhUJEsiG
lBjl0OWcUtL0jpsYsUGQwvF0fY3EsjYf9kEh5DKpAvFDHHkt4EMOZm1KPVFlPke+
kMJ2viE7mepzAxclHLOP1ZeGsisroCV417w78YSh11GWB2YPPTNuhlzZA9UIQMKg
2SOTcFx/pm2KSPaoPyEIu+l3EkJplegD9l9BLya+0OeufWeINd6SkzSM7u6wwXtC
gwnrNj6yRzrvfDcSkP0YIRZff8p+DU8Ir0fPLvmCLzdZXwC+zA6Lk7sHNiLMKic2
FdY+lpXo3xisSQZWgr+0515NKkm3NZLxoFLr1x5dxeAgDRd5uHhJAK8z/9Mw6qAs
pV13X8d2lwGKvMrljzFXdRRoL6So0Pyk/T6R/PGXwjiuXjUGPv/sNWd4gdHeULK0
yi8mc3URdjxgUjak4Dfy4tkUkpeoLxzHSXGA222ZuqftqIZPNOYFhfTQtK4JdMhK
Yfsm6llkh1zYDmLFq0beKMJoSqEFOJdoLBjt1KAcDeBrHtv+TcEU/Ue0gVt3Pk1p
WeJE/zaO+WYrF5sqhGNmpaZ+K3/FpRfog+FjvVdcTKmU4Ek941+H/UXXJUjaq1D0
JptnfHbRmhdblcbHmUtWaPPWEdfNtcUJHxYxK0vszScf3bI7DjxjCPKwk1CVHkqS
J2pZhh+bGgomLzMa+1jCWPO4//iD/sko/RPmZ0lF03lLAFC7msda0wR4PLFAntZn
AbRA+r7jeE998C0ujG7QpHp+E47N9p8o44muJollMnTD0M49ji5E7RjuMng6QrKB
O3UD8X0hzgCvwth3eFYcUBhkA929ZhxomwHbt5OAK92wCZNfpEY2JJxcyM8E8CSW
1c7ydaadaLm2o51xv5mKKB3tnR26maxnD7pNBaRpN+2ZDcGaGvIhSejFLUUHcC4H
yZc1StM1WHipnhTw/8RzHMbHsFTTEK9SNSrqLpqeRjcVwV/ySC7X+sBwxNL+/hL0
rEGBuiiQjGH3Kdg9/RHm+S82GHejFa1x7A32KQ4G3X5IAbrnfB3NOq3NgmqfPmub
xwuYQOT2uYSYz32Wl9BM3cbZa4AwqddHeEyh+olPbcImZQ54PiVcQA2tMrH26oWl
2+cPXnd+OXmO4JCHC24Nz7/2WBGh4+hnasj6Y/mvEFh8UeaTL5vYjgIA8A8o1vrG
9rcvX8xTXZr9tgPfIt4mVJnPCZjxGTQ6jfKGjgZeMK8FzhULFlpiuckLA3RFqIAp
+i3a+c9GNWdtZtBcg+Ce3a6DNU70FoQsQulTTVD5Ph6Jy/sOWWBOjHV3fvvWhBWN
/LE3fmklwfvZ/p0kwuxwTTUy3OHUrPyTg6hYfXqilp6OVBmhpgndC780g3wANzV0
lGD/zd3iVLdkkkGxH46EXO3Q7keuH4RGa8mZffeLpxUNUTPxtNTIGBYSOcsLVJ0J
SrV8D0HaPVqJb1VA5O1hp6TWGQQC+0uYe8B+hBnSfK9nOWWdLJw5knPeX6o+uiSB
Twd+AUncG0AqjU3i0paJgWZtEFSqUotK7FPg3+tnv19Y4I4U+CYTD1YjxyofV9hG
5njAn3j+IBDCpRHbhjw3I2HGrFDaZBxYV3RlU/8WOzznO7e9iKpBKGO/FMmJgTaz
ZymkNx95QLZ5Cl1ViIw3ZURD4kI3BWSylxvGFKhNiquwjPCK+hK3JYd1Y85dj195
ibg3ZhmYsdcoEVSIlx+GLWPjZHqmVfFQz0mNul7OYaTwrvRtTbzAGuK9v6ixKs2N
VIXdhzOvTN3xA8T2+TIWCNRAZrgeXsc26r+GvI9vfvtRpi3RaBOxkuSajmWlCiXp
kKMnZU/yuAvd3szKZ8FIW6jQKPY8wb/lxnXg0aZqFDo4fwLCtnK758apqtY39cp4
nKxzrAaxltTnoLIKrlLpw1B4F4qo9L6nqetnOdm8nVNSsJJT/+0FMtDRFSplfxHD
yYiv36f9+px6eufCDtaZ3m5uHbPJX+kbH56Pbv4VVWBGWm3kcsIiZuiwlksvFLgL
cMfmJXDOQdXvEQIX9OxvOckiYH6Hqy8ImyY5ONaiuMLKRI/WYCcIIwYGwJDZaWK0
YXsNKoHQShw/RBVxhmS+BBJoxI/3VachETIQ5K4bZGE4geN5JqGFmUL/SuTReghs
HhRpNFTGFInoa5DS9KGqi6DSH6x6/gvHIxNiWB6I8zkelc72KbztsCUKWJNxY3Wf
om8kcatLc6uF4LTk/+GLPIVoXlcl3ZioeCasRIOkY/YYhrFcjFlLUM7UnAPHlXZT
bUuGJ6S7PmS/YZrT7TwjgWdVqNNy6PV9izxFeIEL5LYF88d2pLs8gG+s6l1CQ6iw
x39UWfomgCOfrxqYkACSfjheiNjZuXkrA3P2R5eUl7Cs8yKqPu1o+asb9lJq1Uv3
2d6vkP9DbJBLUPiM023H1VtXE4oDiaOBg5hTzow9b9O9pG2i4l9uD2sNxk5NTGX8
nBXqgqnnGfxoHMAujgqripe6hQcfKiAjvV1vXwvBR2R9bFeNewTNCbMc+s3GaVE8
NPcR7O1hQK/c30dzwz9YrySHrcKVh1595effL2JLn9VmAcTnR5xzI+VYTLu4ccox
jdEC+2VFrLbFLR39vrBTQ8zid/teGdD0XZaRGM2mrV93OMhRpP1JtxWhSdV8xrBe
h3c1qQ4z82leA9BR6bjLsHpGfNUpUWDXr6SsOp7zOhKMu/mi3nSUXmDUMsW08TEq
YJWV3pvFrQTxLoVRPqxSlZL2IcJiARTqoUdKScHfxiJ926fUU6HUl8zTzgVzfZBA
2ZjmcLZnHKGGlN/BrhKCQlQaFaeNmR5M3qNkZaIck+LYi+qWc89lhLpbn4i4gDTx
+m0cTSxzOOMhIZDMD8+6qco52MjKPQwRsEVJn9gHNQQkBNRvhcMlYGgUwf8QD3R7
4tST0+hLbhTAwr2mRi5m9VMyLijIcDrq3Td4RrRwgKEmQLBWE7MwpvgpXRBjU2jt
51NAYprPQewYASMMGEmwvAJZ0uKMVXhC+l7g6CZcaQ8WvVnYs73j81RWzjyA6lej
3JnXuXJWtHlu+rccYxRe/cPXiz+0amcYbgWtnZAWybzhTdikdM8B/Apsdr3JlhSu
+XM10EXkya2knDXKbcKWj5S/bBFQZ3bu1Bw2e5HEO1g6cz+e2OmxqrQu1u9d2bsh
pjzsjt3LD3/9L2posVpubpckKOViCabnzRX/5hUP0FbvW/by95hwNtnDQWaeWCeg
26wjgr7bhpaWGGji060qlAct1L5EUSSFkT/U+MtNt5XB+c7PM7Gy2WGRzg64aHCS
+jFhFlQopi8voEfqIDWZ5m/rpu/oYBh/ExjOptQtDsDXR9eZgkflwZZvizqXX9zH
5txzv3OWZBM2l+H61Rhu90PMhjlX4Dc3nUgRcMsoZllA8nnsB3v0dvJQlZoSEfno
+Iab5b8v45fDScME/Pqw3G9HGB2irTA1fsZaffcU4Osxn5Uut4Rl3ydUdvZQvdUp
q5hg7eNo9UxbI4cbjM84WBEXJ/uoJNmJMFkHnNofEmLvCqPOqvClV2luz725zojH
lqLo/2ua0t1WlidC1EJPXuGjQelj5oR15UO0Ke90EKFCOWqdbR38RYTPjLS0SYnx
bQwta/DZ0D3kMlmxkeY5VEmBKuJ9yILOlQiCpX4dj5Bp5UIBWIBoA1qakOGHjxY3
2dXZ4o5DzFHCD307uTxti77NmyW4k1maMYEESTz+pkxjwRG5AooO9dG2RBMyPe31
2TEI/6vWxKcKtoFriTqNrz6veBgFICu3x8WKiYS5Dsv8kzxGLbJX5sd8QZnlttpl
YrXMitZcsLrf7Qq/IRfsb30KJfITUus6o30GJ8UD/sxPMiWaIHzT/g0M9PyNFKBR
JUNDovntMepTuKpoZ2QVDgudIFlpxWM+SqbCLjFilDDdV5r84P53OVhqlqnqVzr7
yeLCsbrJJKULxojJe/kzqyk54lvlmeYHQzDaX0tmVFFdIVnJ5QZhPIiQllzMqkTl
oNrUb3QaXHUmgbc0katMtp0u54XcQJAz7T4WyD+3FW7JQoM6wE9+9E9GKw0/rqNz
bJT9eq+LpJtGIZyynFfNogitb+9GW2RPRbPtDTaY7jdyELtAasJxvDIFpaZ30c2h
0Ii8rMvXZgzUWz+Babw96eaP1dxV+8gVR6gQ3mhu1F4muuYUcANGczjWKtEcHO0y
Nc5FUEvbAAi2wQPxFR2QHDXHJiqlPZ/QQIbAe+mhD0viOe8DyhxmRxeLxGw20SZZ
km/aXsF9aH/1LWz1sWdI9YJzFt+gd80ZEKqaHE7pIMHvQ/5JXkdFAyGZeMahKvEd
P4D0TmLJemgHG2hVIFfhJpKEEeD4LSF2kyYlPbNDBruAldji/x3wpghjbrqTGzUu
4/jJUPJNyN88Xm6gToHNq3uf75gp4v+kmN7begMHGrp5kcobk29I7oIOK1ir4vGk
drAuaqjLNdCg0ii0GQ4mhkWF1fIwrDUjJFlijk6Ed/vDYueNtaxaIF0b95VyJgtq
1/kBWBwheMKd07IZVqIE018WdCdISEYanW51pTzgBRb6N7ywJ3SUjta6LULKDXBb
TSUimVzW9+zNAnb5WJjAhpuqxiUgDeOl5CAuC3Vjl4L7sgdnrBd2wCSAMQ8ohn1n
KTadrSPR0F+6vab8CfE65BYECPmOxjcaVix9SHfrd5xQp/6fyGNtY6RTZG9+59jc
tkj3Cwc9ANK/x4ua+eJ/oYbzPKFEJAqhEsioGjoOVxuNi4udefhq3oMPZhGK350r
t2m7qBJ+rf6TysDbamj9WMCDRU4P9xvQsdofyo+GBGZAIPthSnBroMDP2ROFZjvC
Iy5t5mrqCHs5J8RDbpCsWv2MW5Bq7JINtAp43HUKjfDtTqxU4hKQzxIOJUPT86Wm
+3LdyIN3butz+HEykDeALdVNe7NLsMsZRQp1NrNhEvBkIW4DrftL357KCUJhhMu2
ysoLEnjximvX9UViXZ6SEfqL8VHytnNEWiRRaUXt2ZQHQWhJ2gDXszMbzAUZ9Sw+
KaDlOi/gB4w4I77Ulqv1SH9boFdDzywNaVd0CDCetMcBwPP+/p/Y1JMjvOHduQS1
IysSTmNZ49ii3Vre7boqGO9lHsQOIk8+p4Brsfnw9ajx8IAa7zGNvugXKlaNf1Pk
Ue5qHKBzWJWgv/wZPnbFBmkffp2jJcI3uTxzDTf6676lIt3USd5dFHEfgUwlBG6r
vGcfbK0a/oxJeDT1YKpRN4C6hf0Oz/N42PnK/+qJfULSX6oEnfBCs4d79/Fw0qJU
cICeGfvmtAdFkrmZRylzXv2vKfFl4FF4iyOAsszosVUc59Xcck4g0i2UzeYt2IR0
1b8DjecHc+eQ2uxCjF0vqSjyqQaa3d6BppFuMd0b6S25QAoUN9TS9dBIbS/JE6rC
JwYFPJEwxfJMxuLybmAZfXlsG9gEpWif5c18mEF8LjxXZhkSttzZEe5/GsbftQ5A
WdJrg7Pe8Mbc8Cg1OiNYkeidLSSStqXbg8NYq9yLMOcBP13twPKPR6kiuAmkI/3Q
iMhGSGyuxdECKTwfyrkZL4ss5V0tQWwjJZ5OQbJGrkbj1Lcok00tLj4zEEjwJo1T
RopJh02sahh7kMBQ+eqfHanADFO+VpMEfgC74bwqF5xCUHzaHKat01UTt8Xoviem
Ol40Y+jqL35ix2gnF/q1NwW7TGSf9EtZJCcqRvnSxcoA/7MRAsmu2EFNOG9h6yJf
TOmRScGRtKKkamVPrA9AcRoOLcNHTPHhvoHQBetxit+9m4FD+xT2lOJGxUQBd2rq
nZNaAQR4406BjNYOrXwYnt7oeknBjPLr+8bTz+6t60D8A3bVQ5uxc6h0ZdmB2by6
HxTI+KXwkWMdQDgEfnVh+i+FCJjdtQbKS0D89gYdisuOuoqbBWDbuejBi1OClm7p
VPStY8XRuVK5syZAKOvwTiMgUJ41OlILUScfA87SaDvXrz+esMfa4i5ewh8mAJ8l
ibIZ8w5bQT1mgxKgAwPBSqPVhI05me9o9tSukq6uE33L0wcBX9/sd25cGCIzB0M/
s0N1drJlFN5RLgcnyw4npOHEReWFHfSXNvX8l997y1APVQDBF6vLMaVMCHTzoOAI
TWBwUWuhVW4EGDj00Zvn63pd//tYV64e12MXMpHbn5W9pbUT8spVnXrjU+zuKjfU
rCbRyJ0iMHEvMR8Aq/TYN/zi47EzQDv+7q0SFZZyUpveqRziSjttGhjYp/Mkyp72
he3kQHnmJfWCKx4mutEniaKzC4QBUP8H3Iw92XoF2HckPrTNs3pZH64z9/iJXj8W
bBADQQbOpxSHMiR1+5FCsA5ZksKwiViVy8qHNkJiBGiyoyUvxxQc54sLdRFnNtEy
WmwyO5O8Crc3Q7XA9Rw9rWh/cMNM0ldGbPq2VpRkDOaRIjL6a0YfyGiiy/t4UoX5
s7lkq7YKBXFuVtesqy7fybgzRYKUzGOpo5jk7s479NI/UH6DuMS31PRK1/okWSKZ
jrIsdyefOvXdelVEUy+UTFH0oygA3lYvxfjNwpMpoix8hTQ0IyDIvItZbSgEV/TH
mEmso66exh3HYuHQ75LybZV57DSH5PLvEWHsf6+YfKukxbMPDWRWIO34hRXA1j7b
keldMJWdE2oNdUjhG0C55OiBeFcx1MfREQWnpZM7TpnO/dbWFH/dXluhMkkWkhlv
6uPT7sbGiaJQrWT1bbp25lw5UIXNv/F2oBcI9fRrrXSsBiokiCfbiYJx3GqMKwq6
OjIyzizJT/eIAlDffZL8lqk05dsLzrQBmxrT/88rgM3ismb91pZGohwOhUr6mrCD
0BHO3zdVPvVPZ4e9CKAx25EcoXOISX0WJ/Ug/y6iFFH7YjEWhoQsRhzcB+wi3Xdk
SKWbiLlx72YMf2BLbrKjCyAMO5zeEw6o6u1MgE06pHTisug0dWwnGhCZ2KDuUJnj
PwK1DbAP3wLYxJpT/cqFJ9W/IOMFBPq6l3k3t0aB+anBHNFQcO90ZMOBBl6Tu9w6
Z2WOI9hIFMoqFqNujCWf7lYZENoDYMJkELYe/1vpCq7FRJpDkbGdk20nXjdYlgj5
TJnt6H9JbGz77qIqs7BCf8p2cxxHZPmLAek8LUAWqzmtZDxZ0I+E4+DgPRFYGYz/
/nnQuTPdAh6QBVbipeqH1zZTb+sFHshsd+TRxsSCRtqdsadIo+9dIzqcVHn3k1wv
7EN/pFq7E+sv5GCE8Yu9mWa1abd9hy4vSAf9o/M2yVbFYK8Y4gvbZGTQAvBCaTVv
w7vUNfIzLVgFUiEQK69cT09aPfVudvCL8jco1ft8yuykhCOcnspBxIkQBJL/Pgwh
KhVTzgrABUM00v/OfAVrKwMWcP2F9bu2UmD6Z3o0cRN5wcqIfqxgr3/TD2g4KO75
OdpOnyOyi2bzNWlJtjh3uxf9pRa06zMY1fXQhaxZdoAlxyf+phyOHi/p+zMj3LLC
ckUm7YM52RzxrJQA1lzKweZWhaOAvJwOarllpmr4T9q1SFGODu5zI02rd8QW8mU1
McjzJ9221I7vsbt/OmgnsII1py3kVaxD0q6n19hmqzpJvoHvhC3jEmsU/OxXnNqt
pQ4MFZr32lmUh7dpspuQIh7cbX5QlcdGQ8jJ9098SpogQO0jRxsTHjsh0Ou5EH7u
N49HTg5D9ykTaOzlMyup7MABK7Ip0UDE6j2ITFykMPw2bSpAoLwc6PxAInLqwHJS
7yd7ctT6Kd4wg62BNSkspJi5MHwtoBZRjECW67btQakSa56+TC1UCB5BOXevrLj9
U86afe2bgpwy3+QMjgYZ0Geio26hc9P8ZmYarFKaod3cfrTERcp7OLzdz5w06kKo
ZiMIdJNwtQbrDq1+CGXEJCeQ1b8grJyAA7ffy0/iMF6JZOiV3wiOlNM3hzONyuH4
Qu6m1DA7/UQY/KkM9pwLrrTiTM/B5q2rjdbkKg+7iX7Bzfj/OoYrGvAnTgKyOxcs
0lU3dxuREEa3fNu7x+u1zps8Q1jfYc5uN9Dun5FQ0RNBwJB7GseiR+JTcrl7it1X
odHSdMpmyWU/truBXZYIiHtr1RYrJAGIO9rR13C2appw63yfWSq+Cm1Ukmp5gppE
9EiAldN9aKeMIFlPy0NJ+fx1ZBAyWn2WJrHI172pzNgLc+c5lljuKT8lXBjA5R5R
r6P1KDrLxMHHkO/Fc+2s1G0V8LV+uvjkjiFP0G/lC3/SvQ/nReVuy3DHw2HoI58u
n1zA80z/Yu+phpdd0GhgVmZZHnph3C1haDp+9VHCWXq8W0GBbPUXShKJiNUkDcS3
/pFIBX0uEQJXoU/a2z7j+8HRgEcmxM3s1MAY/59Bov8L5reQ2nR8dHAeMY95lMnX
p8vsLKLJ0S9hI9cfmK+gnhBHKc0S42pjpshrwgohiXIvZaXhnTvZWozdCx0HbaGe
faG4Oqt8aQkOgGYb4IZ1z+9Xugcic6D1zb79rGVL9i+60hU1NUF1QpWTHr/z4hUL
5Uk3FueN51/12QT5bDVYzohX4ZqQ0TYRPGuTdqMCP6SlRblPdZFCbyfiImwk2Z7+
jX31xaqG3hejmi9x1Y53SDKKvzdzJ7zPOOE8IPPX4qbMjCa5n1LCUuPookceASer
q4DkvHckMdmYg0cnRcYGzt/MP4hJxkFJr+Hrt9qUQut2rB9LyKfLsy4f53JCyKr9
/Ucn2RX+SW5SvI3VcMjJWWau03m/tiBjegccfznQKWURm4mwdczb2Cp8MqoBabrV
55yrTR4C0BJA4Tdm3Ysf8f1LPcZOitGnh9sAWu5gdmMqNJ/PI214iMFaQwlPvV9a
LroraEmdWZlMxyPcN3evNimROBhiw0MtUj0LF2QOI19OfJ/WjbZOBcARJ4GeH7Zr
2iMOx+vozDf8ck2WNWOaivQlYmXTuD3txhKa9exd9ZSHCqrUn9P5nyheRYU/dJ2A
iy7KLhZI8PGoFTmIwkXa/nAxdHKGtIbPzrWiRPkcqAN1x6UR7nvH9Vr5BDpZBmtd
47I9BpT1NqEFSDfVZZqQiqblcm4HBCRK8+RZkshI8ewwZSKsFfxsnP6CdzItSgYR
cl14smXi18EorESDGxHMoRAPD2Omtd29dNEvhjgq8Al3luU804F5YVMWO6NJMxIC
i4maS3lo+Ehrl9souREgbtVQlbhsKTsDDMHWx0gum0VkC/oIfYHGCiVNiwdp2ZpK
2d9E1XKxJJx+P1WY7vgvItcIBDYQdFf/ts6GQ9tFtpK1/iVpDqQWRuQYb8JDEyNE
fRMRa9OXo+aaYMWkXVWvnQOK6wRUFznDCY7A1RI6boGVX8l/9JH/SBKyhSOt/m6v
kYj5jJKa9wHWONIaQdEcPwDNZB1DWjrrtrSV5nwfD07uFybbok4HQ6r4HDCmZiFz
3v65iASjSK7WElvHShgtKAvIV9Tg47M0UK0Qh+IgsLycdSlWowm8xkQ1XZvotq42
gg8BREm7FTKlwIqXNHIr95y1HaeQGbg6NzcKCzqSi/SaJHld1MNQIdkCb/RBeyfD
vHt4FF2l5jCaAjrvlrAEYPGMv/s00RdnHw3Dq0oiX/zLIUx6iWb5ffcNw7NOcIlG
41NZmnnA55fjbLg3ga9+goRGkT2ndIsbDrTjyjckmHNdsANPhkZlvXbYfO4vJkmS
QdpSkylA3w3VWoAY9T42JFVbSdBVVccBem0X1DOf0Ax5OWHLMVxcn6yabxw/i3Yl
6x2vZKwkUQElT1A96DfFxVtiihMKAs2TBLI2knnPwdlxdWTU9sRYZGe6GXk2P8j8
MgJHyaSX6XVsKZ6Ud7aLhfB0EfV+wcMv9OFdyiN6d7ord5nIfbECE1U84WMtBzWb
NvLvldtGWyaHS+Aq6iyc4UqB9FtJR49ThyWrW9rcDwDbt8MZ/2HIxLfwOwI1mMKD
LZ8dW2zK/Axo5bNU/X883D5mMFcpB5aFkJB+QVQy165fgHBUy37n8u9DPzTVimMN
Zh/3SG7Znfj+Zc7RRpUbUYhzuTrBwKKkIHUotdTVO3AqnxZrKwAWVrz/dcLlB+Lt
7E097paJOvKGQocpQXs4UIcD1hMz5srKoULIfzSYHwwDo9I7FTq9ZFQWrj+ZZdFk
bUj9uQn6uWhMwxtT8Xqq454nt1jupf8twYUkzHrKVLpFmIITwWuFXKz614XsoM0Q
BTAdA7zXe877j+wHzQ0mBg4T3QwQr9i8jfWiZ3siRbxc2Lsn//bqAmM6v4oFUFIB
PIgeC4YCOA21Aqn5KIZnkwJgEOYCxWL4wITvZgnOLy4+mk6nl+qtsFF1atAxxbX1
GlQCodVwME6ipJ0k9jUrO26hQS/i/GH2XYB7T0Di59a5CbzLDUC0UAZC+Hv+hqQE
b54LA3iopJYMo0NoLhwfywzwsTwG4I2FEVQYLXMKz0iCwMYIekL5uNRVdZY1do0G
3RlD2rMArRaNhNX/BibOalgszzqMfsT7zsomfGBC9xzQgqM0DKgsuPVchTJgIZRT
S7GgpuCzPpfOleahfNMVhoGuEFCh/557X6hkiPyYbyLR2NySSJ0mLkrU8kXSrx1v
MzBDjnROxFjYK2wPnhhMmaA0GGW7QoL65LwP05kRclflDXzBt5EKG0nAbgF8yuce
KJE5rU7vjfxyMWSKfIUaDXKd7nm2PtnIlt2tqOom6KFcUJZQjfOQ4MBVWj49hj7B
kDuZlM3MMIOZ0c+1yqX87AOPlM6no3eJpdd9ij1P7l/KO9rUUHutIwJLOz8T6h7d
WSCF7f3qOu34z8WDohFX447xSy8lrFYS7oF3duvJA4+rbGx2bSruL4wWrN+ge3qJ
y6Cus/cZhZc0ziORvhfVi2e1/gxeZ1YcgdGaMNlbWwlIeUevpK7vCqI7Ry4vTP+J
+AnHSmxjH4CkqUY9d5JKjw1wz6/qEGoqgGnCodT9N4Bd8WFyGav00K2lp74bVhdC
eR4103GJ91MnDquMvUwdmGHV8q+wHslyg15GN9zIymkwlo21PQVv414A07P0z8HQ
COAdGShtJQHbksrrJpm70EVgDUXQRzJsTZC0yFn4jF4L+lHa++WMy7EoTm0VERR8
BfwUb87iP5JGfOG8/e+zmY8o/jYGtIsCCoSzc5E2jteMXkPFZUIf4no/84qbSmEh
tYcL1Kja6SbNeClpbpiJtnA7MqYSPyUygOHmWzA8FQ9EOubEWopBL8CIpm9dFLBU
fPX3HHxKjTPEblLGiQHhbXzQhtSod+F7qgON6QrLkPiYcMp2FmCgG03bUHHrXOTx
0z0mJAJPkV5Lb9m0tliw2B7cIX6oj1FsAKE7fR3thE/zgQopmTKf6j8SgsQjFAs5
sW1B7hfwfnvekD4cBCv6TkRMaLE0okp2PBo2qAYiireUgOzivQFb0XfpSCOAvJSf
jVVcmd56twMkYA4Bq9xT+NPHu4Y+Ldrru8rMIOF4oqWLUiemXl+1P4wod0v35Y23
A9h8lvFqkO+MG3e94nQtty8/2w86Y5ofb7EBKCs9DXwXOR/gMcZMa95KLZIHtmVl
bSJmIogqjEXc7dxAUXPz3JjDXe36+3ZaWr34ByyTspRAU4Uvx+Byyk82wa+8k4JU
IpJJNAoYyRIUeNW2RkPzzCS6+PXP3m+J13lbPZ0jrzK06TKAuS5os0dXpCwZ7pL7
Oobtf+tejxZHocmKrZ0OrkMeyiv7rb2JpcyG7U7ZvyzB+JxK5Vi3ktiPX7gnyu/W
JgTlv6HQHgTILd5VJbhG8DMU+v4vOIVxf/T5SdWk0N53Vs9tXYetyqAkAyNNdBiD
pckCyWvlKMr+OFqoDBABV1qOvWn98+WnbQMeGvgP2QeefUjcD2Eltm07wMylIhSI
1CbdxcoyLmrLqLbnfKDt0DnuDQZu+QnzMTkD9FyCtlBIxdMT8mcQ2Y/M2wod6JCv
NdpRo4ibVy3pSpgo97gNr1kQcIc5i5LXnPH61y7FIo1uwCtSjBYl6cRfs6pHoupe
sN/LU6am2QX2L8lMreodWOtv3eeFMbDkDqmYAJeB2I70ifTKDJNquMvyBnZ9lD0X
UwxhNwe5rfHcWvmmLzGgYQh5/odCtMCnjFzZF/r3DfdpkmVzx51V9mU1JY4ZtpdS
wFDFQe425+7VC8fF1EbO62wjjlwDKfIaPrLuXfJLuW5DOIfTWTd3G0Z7cXGmff3W
8xul5cdxFGTkvrlly4gYIIhHJMSFx1XOh3/VXxpncR5j3LpA7bimiNsOOiCIKN7Y
U+QGSoR2VRuXIwNLONmEDyqlizS0dbgbaxRsOWaci3d41he7ON3ksoUwjTovDwqB
ls9VpSEcJV/0nstw5++EaXxNsR6JVjsn3DiMH8yRocLDr5JmgHvj1sELoQef6wy3
BBzltBO4ykzlL8+qRni/3q3dLm/x3WFTMKhda/IkamrCOl1f5DbzFQzRAcyv9fo6
6lXFTwJnFD/Lac/7ip6XzAqD/qxzhGZwlktdmAfdMlSqjz8Hd4QK619bUOmDVcUc
JAml5TT6vWVqe+sJLFdSL79YJ+WINchbKHNK2y47prA0Iys1Y09Qx4e/WJpKpa5p
VQNnFquBMXko5mlhuKT6l7YYR6FDPqUJKB9MfFi9c97lin1ak7e60znuOCemN/Wc
u0CCQAYWGt0ME5RgweNQIlubDk/R2Bfms5K9beqjxf534glLdgQKuKjlszfZjySe
wNJYQak/ivwS6mIKipJrZrl0O68QBkiggh93QFJJxG7QCGJdfTrkyWOZil7qyhk9
kOB9r1HXi5kVWHDXAewx5Ic+5WEOOyPx8hAzl7tGcKv1Hg17DkQyfMBeqUVI4R86
aPC14GeLnFhmM/da7W7uhnddGdHziyzEfCW56MaZQULXZ+Wbi4V955d9k0XdKMgo
wGdsZwp1eP07nDgPtPnCxDfqokPQbox/nRVmWwkVuIEACBOtzg6EQI/MJFDhbInh
dh3Bj/jHB8XmEQDh30ARBm3sCMq8Kh4lKjqmsbQg4dRjUoJaPvRCvwGgwezEVg3E
G2xBD1/uBBPoujmhy6PkScgOQvx8dee4lZQLz0wa/84mCgY8zwqiO8fgnL5QKFRn
YNitvi56DyCoBd7XNKH/TDF+iIUdxV6fUHhhfO3wM13w5cC5Q/tjey9dSFIGvnGv
0EQwQ1k4uonGFQycNcHc8Gp7i1OLoDJcwhCS7xfxVPH7NOnVwEHJjjc7wUgxuVfr
P0+yOPFVMOtR8FA53Pfeg0pN82rsmV5tC2yFlaZiBsbC+8uaAbHJ0fyiMy0OZNyd
SfAhnttfuosfXiUnKeNpqiYD+zDv2cOp2VlueOVxluhQuSpQ1SKCyQV5C1y/Z5FZ
q+G3i0FIwkaGsXn0J6DA1sNE/mtf2ITVNjwgpoNLRa/gZnZm8FWOe9uN/RL5oC5l
9a7qua86y3hPXnSwNtYGt62RmLrVgzGBcsbYiopSUq7nznZ7lshGEPuVRT/jEHPS
5haEp72hndV7RTy3h7+TiL/qiMAUNRP6WF9Oys53IhHdm2l6doCzUR5ODRcx2fXV
AmPLvUZD6NoauKYkrh3GnjRpNxBYG/7uXw4/hjC2tYnl0adN//Tfiqm1J72C5k0H
zAvDo12PyPFU5px81bq5Xb1EEFoQHqo+RRs/Il/koQUy9QYNBsi9/afpRpfoMBTe
c7gjH37yBGCy3hN9g2iubOH6dWmeIS8ZdblW6A/9i3ff/+kryCsEItmsCjGjqW7/
TEwhyF9hjKzSbwph3pWvyWnG/J/CSx0LYSor8nPanUUgQpkR1c/r9ZofOoNE4a/K
ckUjPXx/KPknSEIEPHiuolV2ow40L3wgImaW/ABs+/1JHI8f17AJ2aOuFa0MdWsg
CUCUSWWHTTwPm4htMxo/z2DsDib1NNVPJG8oBSJgN1GMwDteRGOxGtl8wQP22oWB
SiBQ3C1ItnVyg5kdwfyUKoPEaFPc6b8YJVqx+/PiXQdB8cDyYGEPQtDtRom4tCCd
3mrIAcV3RitleDmpQ1bvpRqgQpjaNR5PkMma+QGyyUXAJYPFqYR8nCWZ/vhM5Er5
SuIK2kVaOF15LD6jgjVGbK18MIhvv/ebwODpeGQQwp7L1E+0l9xARBASZnn0X6VJ
A/mDPWlBdTxSVf1CqP4qintq/OAvjsg79P+EdMdr1f8FoxL3dn7EjfJyJav4aa81
7+ialOdK5bxDPjYv92tlkMJp1Ssm2DtMI3L31zuf32KubgiEdWM/kd7CuCjWguk0
L+XSiKgTA6iYt6vjTBhMAT6oAQBEXbgGpGRpH4Ye+z6vGG7hmHVzAEbnqYiwLwyT
iUZ+DQGyaxSn5fYrgX++gaVkTVD82rU1t8x1TEZNyh6x8yAVNwBJ5Yw7lCRVYXWs
2mqMNnew/3cxa2i3xpcMA/YDinBHYgUBXyGta/+cED2CLOwkf86lo7DQncZiWa2h
c9bhgwGkeuwoJJtKfrLYehH5WPF69KkSfByp1K2T99/QqLvl8AYriiqQV/4fHg8/
DGiX0XunbwJ08ilwbCp5PtZNyglVakotGToab3WlvzmiGNofzdC4jG9HvZ9wPzHi
j3hjDupgwevkvwlwr5y8n2yjSi6p0LpPRHvku1HJZ18cDy/rE56VNQYlAlQP6jwK
xSfvZwhnWA/r0pJ6zqSVxzGg4OqzScYIMef0XjRsVMMe+PQJ4fOZkLyRpZJq4p+H
6DXO7lpirtJmi1vUWVAWyndZXCbIxz+2b/Mv9Dk3hUcQzm3UZEzqtNFJXehihdW6
R7fzMTmCI19NvwsG22F+Kf4EXqW+fuy7VGpUNToRPCSli2opKMCHnlf/RTgYsQT3
YinijMnNoO1163iBIlA81VNrgATQTJIdaw7t+wR/wAHsgmrJDT1o0ximXDBU+Gv/
JOx6w7RCEHNQ80ezvR6POtkYKCNIhP8HFkZQV+tKIp3TW4e+/DYuhh3nhgDBxr7L
C099YwzdqpMo4ZiI2L5NIFADIDcnapC+3xLdNrbUmd+HVDy1zOYO7eWQOoySGIlb
RiEzf+YLZYqY4woheRmNQ7+OiLa/Fx4o4jwt1FWf8E/uT+bvzW8MjjelNaPIeCLh
Sge2L71bemEYUMCIvROQXS6fiR3tbHRnzh5QwpFuhARSEKO5xdy82TjLVAhRa5uH
VwgE7BU5Nxn6LKRYHoSr2NDKWgtFT/AFRs5Ch5QBAE6pY5xrUQ07+NpQeFaTrUfR
I0tuVsMm+ZmOTwIvx0B46xWkAvIu1/DM9VfAmDrhQLrhBCltB4GzJUdDE2fFbPGh
G5vuZlhFEl9QDW06I7sPExEw8gervkWI3KYg4P/ZZyNqV0KUx+yjPfOJC1E6XubF
2PKBpte2Kwwv5KZ0DPvGChLiFiWpkSSSRekI/TzDdeN0Ydg30rEsflErrVXcpOme
8mqFY+svx57jl28Kv+7RycALA0KXPNyFmFf+wN2iWofnyr+xnBnJksDla5iu/7Y3
i4fNYvXZwrrx9tHlODrcM8AAMfmy6+vimCZJLwo98R/ZfXObCA1NN+7Mr8lJoilX
ZV6HwTpDE35FQPxXj7hOBbIoSkw+mwkptziU3UOw+8BNQZZJjuQ9SmQqoqaZ9kRv
YjYqJrTBv7aolGaF+onVFthnz6xD1VA9RGqCvf3jkp+nHrYTzsB713i6//dIDMnX
5J+1lAsR87+/V5F46+Vq1zqjfBSFErNevy+dnTeHpC86XyK6qUzKuhwX8gwwCEzn
ZituFC/wBQTed+EM0CEdAQn3xrFKOedInq7kTFipXTVA7v1cfS0Mi0xcbPjL+r1X
XuDOIIaEh1tKe+brT+meYgmXRtMe2CFOV9pzNxkPgBp7nyt5UQ1UEvXDQvmEoM+0
0tqqZ3wUNM58mp9QY+Gs5dMaPzHCUUonDPV95HAVZCUNrB6zAZbTsjrntF3tqsNL
cqnuDvGnH45olKLLu+yBq1zCjXzUomJWhX/cwG3xyz8BMqdotWpz+Ep84dNwGYPP
oSfspW/IrFFMJOFlRV8m3UQ9CaHa/WipNKDpI7bfRT5DbpSY1F2fG1HxfKCTCJ/O
gHKPF5zvLnedoZXkkp31ZUvq7Dx77JS+ZpmDbTEzDrS2kJw0rvhJ09p37gAUGz5/
br9wD8GKZhsitA/ZORbFeG/Ufnu2QZ4kuPSZcyQEx1yq11sGcG/lnowYs9ggGPe3
CD0AqiXnaZG19Lf3Ze38IUl+TLXuDAWbE2LCtkciiaVm+4hfrFKVPZ66T4bEsCXH
7cp4TKhJkTv28uemdSqvYHy09Ff/aDL67nNi75s5tbmN6ZJHbrSHVRMoZzZH0dmB
ebX2vJ7qRTVyqxpljGOH9o8CXz+zgOICUF+hZs+wPMhACB4PHQ5FK13yNp2vTXWb
baM9prxEe+7XbaNSPDRaQSV23U/HpsIjH7KLbHtmnB6Bz24tXWPD/155QweaYXbP
X8srKKYOjnQA7XQ0d8bl6nUvDtrgDapAwJ0igbklxqFDMwf1OBfHrIgAWOHWH7g1
0OmT1Q+K3TwA62Ui8yTdcExcpop1AoChtHgxolZzosHQUi5K/SCYDe/pIxCdBe6A
NvmpkN13UO8LCriXyDrPP+L9RQbFVH93VsfiZRBI6L/E7B/W1Tqi9xwenjMrtnD8
THfLBXKy7cmzZY5rA1NW19IuEtVTKa36ulma/Yl8zgTEeVM6Bg+ctmMVlZ2u1p6J
AQ/Vo8APbow9Vp8XvUwCUk/NgKrc2DRpOa2O0OoV1zDK6yIMkoOOLICTdIc0dlMr
iH11g6+HH73DYN3Y853Fh83yQnFATtk9zYfG+vfFruW70KzyeS6QU2QkM47JwkCB
m9IHsUC5o2OskZ8yFEcWZEk+E1RS3mcVh8nl3urAZj/APgHrKDIpAGQdhEqRLngF
lKUqQlvVJ2nOY/STXvN+pwOnYVPsBIQeiS3Dp/OxTUfVD80fYbjsCUmh99qReXpO
xTEUdJ2z2K3tSDV3bi1UbNr5c2xXFlyflax9QGLMKnb/Qp+KA6StzYipX981Ta4/
/M+kNwgbD0BK19HHJsAyV/aU5duLKLVdd4yi4Zz2FCOlT+5yKiA5G1Vc2iMGx/5f
nKt/esB8XkUh3nOMiyZQX0OuVgqq0KRAxSftk39C1PzYruAjsX+VZwAQ+tnzuyeo
VBQbb5L7jQil/awaWiRCNb3+v8L1XnOw/acDwxFIaqfmxXgKfDqu4B7cmkuytcT/
W6yqVTiu3XuhjKDE/dxejiIdfsHCiOPUwhEEXlqEWD3+RL3kdp+bDUeQN9jr80zK
DA9EMtlowwhWOOUWr5YevqFtUtSpsENKlS62w9YHK5mo8eaRFthC6IuD27tW65hS
9ShLXsn9nerIgbaOpmj8k5nFKwUKYGP69yHjOrqIAXVflCsGy2zQKmEuGlLBS1tI
IC5Pckk2i2u/IZUFKWmddMC1c9Re79oEvomaryMuwagSxv2QZ5ZN3bgaPYxzt4yM
hWojfJrJ7B13Qw4KW7ILtQM5NX9azzAUc+RMlAXWrbgifc3zPetehrjR3kRdcNV+
5HpST917fFwbRbyHTs47VVju2MhMb3FicSQOrOcIp8bCKQeEHJzNa8E9wE7sDXlR
ELFWjYWkKmWrfd76lLrb0UbUv9xywh9Gyr/ujxm/UBLXJcQjbVgdUaSFW9EzPepH
jbBACKD47SDBVdzPWIdzbIX+A77F8JXQstRVqRDWnwa3oMkm8oIAOOS1rZVdSKQT
SC12q3GYumklQKDYaD0Juu0+Xi9KTXOPGoEkZLyvNsEKO+ZlLlNty9BgYMAkM6bP
+AfnF52RyxubktKa6j7L25UGN2cVMC1jp/K6L0HnMG8m2IY3kH1kykUSroiB0D3u
NsaB2SWQvHSRIutOqQ6p8lTZ5jrSjS3oj5G+pFKBRMERD/nFB7T1PSZi+3BySrfR
egLKc3q/gTGkYWFURiZZMf+qT+NzZxDC29ZtSMdn1CFXY0Goz6kb3JNqCQ8yJaSu
I8FrjGKmkz5iUBiK72BE67fAKcw6Z9ddZ/HXsvgNfFhKgEedyWaQksNW+ZfAq2YR
KPgKx+pHZ/O7wPi2PCPujTqZU09x1Hw0Eo9dUj0HOU3tKsAiKA0wtzgYAMQq1NXv
vJwfGRJUS2wbMnTpa6IMin7Vl3tP5RDqts6S0bAya++yrCBXC0Z7xFvMcmNc+ZxU
HWkW+xIYnKH67noIdhsDNxn5vfIO3OEwzJUGvot7xxOWPXuUuJdHKZe+ygu5wE8U
2gMHIX+6ZNDlWmh43jtmbeGoP+v5Xb1FyNLgOXlTdIKSWcDL1tgOg0774FN44Us1
ryITxspTXcQcifuTEwwoIZnHWs24mb+wQzJVPh26nkg3Gs5aexBnuLEJs/GUCB/B
z7YmBFJH9kwihyGxabIQ1KpshIaib0ktCuHdcPscffNZMAbWvpFG1oYQZLI+ka9I
nG3Eg9eWaLmYVe1AIAUyclWiyx5fKEJQfw7Vc7z73uLg2VE6VRjoebebacWrJU5A
AVudpBqd3+0BZOXvQy41dolC3dGJufUFHxvi1Kv+wB0POUnhViZdYnXTbc0m0Csf
OMg4wNcTbCwtkUagioF0qw8HuUslQ+3E1C6yvZr0HHy5EZ+2VWpXSLomdFOptvvQ
HBbXUca34SrLaXVOqTJByaQNraiOwIFmdXIp/Ip7DliFqHdotMjYf85eWCfXMSW5
Z06wM3R6Oo2keUFKLFr8c8lFOLLvpkEZqvDNPEVyXhTAk6RHMbgrvY4SkBdQGMaH
FetfHYzCLKV0cd7HsVW1dnd8c3TU/vGe0qK5D85dg3zqfygjlDqXgcQPhENIQNlG
Lg3yGBnQm+yW59ZGWioZefwbqRYrDmq0Fb7dj9pdM6wo5STmI9rYaMn1RJPDB6ix
8llTyutcTnWxxLEkUaVQItBdTOnZgU0cbl5ck3w4Rx860W3zbfAAseAp6Esg4aim
MaPCoQ6KaUAkbnu+6vIFu8RB3sCCBHy6ttuiLKyxZe5rEDbPZ7mv9dlfzJG+22X8
RyRq+8Eimx+AYJrmFqHd+DojC8c739yos0VpMybKXrEk15sjLx/12PJPTN7BGAsu
bvL8sPz0rm1kKOsS4Tth6TPJPSu0P0UlLBMMDl9zEBoFnKOKQeBXpKhmIbOk7J3a
jCpwrh/VafYa/FpfmXYIEIt6TGFHWOtMGxJGJw0fIAHrUi0+3o4TqxAh3+J5wlTJ
17tMEZ36HBYlfKPQ+EheEmVk5f/rSheN+Z455XjEmD6/Z/PuPSAVekhpHkx31x6W
3V78Mhp31/QdtwMungjHwuoCS1sZ5W5LLkQEZzMIFE9sb2a86wME/NT2Vc9kBq39
Oif+6tXgkwI74Hn68QUidY9S0y56Sv0cmzJgVFj/pLOzzfZJowFJGmSE/dpUMP5e
GddCK/C1+jU5gxLz0d9xuSd017xyUGu4JI130HIozghXdMyBgQPfwUGBs8PSo4zR
u1m0B5k6NhN55uk3hwErJ4BdEswMziS5TbcBW/xLSWgI0ZQdRySBZyA9IdCwObj3
+88ZzzRcjqFplVNss3p7KVS4JPzCT0b4SyNg/FAiazd1jkvkNWu4yo9YFwbze1of
X3OSOrAbUZ39AICDOD6j23Xpih2U42PnrwSe4nWRzF4eRKKL5hg9A9wv7HtNsT82
kdwERUalw4axyJmDL2R8crp/86NYxsQWtuFQokKS2dE4RS0QoMmWLejxX0qS1z6I
E2SEjaP18pX8PWrwBUPlDhzwjVsA5DZbiqGrY3bk6MWnqK0YiAxVP88xa/cQ1aaB
3jossuNMQ1syrw3MkpGw1FLKtGEAb52dM4CoksdJhP6QS4NbJz+Bkx+6H8yILjGP
RjZMhhPLB8U/Q3jvogBkpHcdyiUGoITxi7dBm6IT3v+YvRhe6cbRw4/xX8yp0J1T
5FbDMxJWcn8okm7gePwG9Nu/Tgmmhi9FN3keUYJGPqVIZ7WtX086FgEx3dVaBs1q
BxK9EIPfhGbFWBH2/yu0Euunku94BAldwCRfYTiD//4LYQdODmuCxTEFvCWJdu+7
orwR2p24O8/rUxkbmBKcRpb4x38l2AcFhuSuoxBb7E2H8mkeQ9kx2u3aem8gnW1W
XYkzOIBJMmsP6FkJ1MGscf++Pkwkf9DNiS2LqTvkxDvDpQNsYIJ0dCy2eRxINnzC
Lo/oi+/V63DQlZnFwOGk7uUZ5O9sLL71GArWsxmbBWVqlvTmD6jTyU4HloKiQixA
5IdiX2dcg6ldpC/KMo3FDfkvOsA196/0lMd2RuaGBfuklNdXYC/tYZDGQhH5yIlM
xH22qF+pN+tYLlIXFnPuWQeKVFfbIoAkOz/KgenzIkigfQBkBKPkr41Qph2AEY/T
UnvdGY3DB4pkfe04+YBewZSdRtqkmskrjxaPoeDb+egYCprqZAiRO8K9HpM4uDH0
l5B5yJeHg34GUOBe+CYBfzUBJIrdywfr1nYMUcyK7IugATzJocxjvLclAKn0Vzfd
96EtO5Vd55D0hqPkEvRCruXMSLiL3KhHhc24L6g8N9rAWJV3+ZFqK7XXBu5XV78K
/INV9NrDjggWmI9/RusdaCsPO24om2e81bczDAg5XTZYWKbE41iW+3q7NhTLElHG
3yzDuCobTRfk9RT9hRKaFmjV36buUE6OPf3kXIIxVHkhkZ+Z3JF1e39HEw7KRKKA
WpMtJOx744KVuuUyoa1zMGIXPnL2Sw9L9md7xfIJbJ8sWF6VlG4C/fQKh2IzsW3Y
3IDGluARny0kJMPXpEjjIKyV1h884+UQGf2dtDDnnw7Qmc/yh0frfz8JBHYH+vBE
KKCcsjAxO0sDyWlIwPlLxrh36RkgniLDopP9d9xh+cykokoPmENrBd+deOcr8SlM
3OZ7F18l2xzr58tVxttQsX/CDCHi1FGe6Tgtbg7Sa3nN1MujGLASjQvVFdjRmiv5
7DmmtIfarNjBvTU9ECyoWT46n0BnfpklcV5Nuf9NyKXwKj0wcfik2jbAVAntAK21
kEp4eTZjzK8Df9mMECuvpal6aMEkA3eRp4/eWh/Qd+Wu0J+O8hE99p/FgCgHPAHe
jaDGbgBav4RanDUCNg2yRH0VnEVdRM2VVKK76gP5GhFuagx2WxYhIpyOf6GDsvlb
JAc6gHGCXUEi+QMyPgUOP8ZBk1F4pz8M/aaesF1RiRT4/anNlKvSP0aceUaI1DvU
d+x+HmxCtebt/7owau4QfJ/5j5I0p+Lu2WVoY7Lqd/MEnS+K/PlRznrGOp734gOs
eDMzZzz1LyldkiWJc5seAyyegqVj+8Cs3RDZhk+v1IFK6O7H5JFyh+3aofy+dEfw
pSLiJ7UeS+HyD9lS4wi/0nVWhbpaWsrV6w8na16rD6ceAGjVVol2b4QI8tvJzf5w
bQtc9x7ZD4QjftOYJT/3jvS0emaCZhkFfqADKedlvtry9JEb5mSnQTZnsZRNtZqU
ZTyhcrWv1uYwB5Krkf1Qb3kbqokUS1Gn1mIjQojNaf9LyN5ixISgxBo0RsxCX4YE
TsLj7MgoTxAIIwlBoaQAyxpujpPuDn825UcirOFsrHj+kAEvvHe51H6Y/h5PAfUC
+nc1lWMNdVZdZoJtQnKgAmNstDAI7zIhGdvC2qNZbZR4s0zwSDA37sIqpsnJQWhM
USVi05e+sUoT9XOu2cApwVrWL4S6qCDN9nO3lhcpw9bTzj09Xj54Vw3OUpwczSI3
mTiBvY5SCBla4/EEfBh3M/L77R1apE9c952aCyhljYvN2zGypeUEkQUXha6wLnjv
RAJe6+61Hapfmh2WR8SS1ffB41JD72uAfJRbnfbph6yK01+KF6+VhGwEss8VUDbC
OfQlqnWqxc4mTzTmOwwwwsnYYkKb9zQG0a5ga08JtWQoQXyy42GbJFTgdoWB1XvR
xEHRzGk7xHdbccJcIQcYlNIKuwL9ADpGHa6CpH/kpcDY+jmOefI0jJO7UhYertPV
ik9qKvtXSqgFr/QYF3Z6dWMB7S641y6G4Qoz3u6PJ6SYNIap3jRV9A9LS2ufG3jS
xnju4ZvlHyikpYnB1GzKlvJ5aJWIRqeu0bScetkVu4GrVjr6drt0rlV0ds5A/lxw
sLH02NNNWse8i9f2qtO+uNWgZJBowB3Zsbwh1ZOXgAR4LAad/R5VxtbsipIIZ1Om
c5QQ01xzBLIc/N66g7n1fIcPPGhbUvk95dkIzIbd2hxPrOrrUfBbO1SFrgiqz+/V
BzySK57oEWQhfOrSdtdWxkucS4OGe4NPqJYnuOpDSUT+homca7n7m0uGsChgaUlX
Ix8WIPeAg9ff304zapKqV2eZeTizEGOB+dZizuikZy8fMXVLyoHJzNL9SfficpEj
YCxUV5Xcc2iO3DpAhEJFrvzWuB8wJWTqaah/EVGGYEUd85SoJShUWoEJCnY8PpHl
9ezga71ISSSHC7JoczVMSJ00J8LlgTHyDRuDjOeDhWLgyj9cCPU3XPM90K3L8q3t
BHrem/O08ps50LmtRSkVKcQrwizqh4S6kDCqRFn0zGteHsnSUYqUSxaQR4rNIUEg
PsZ/D5PqjNKM8bkGIlss7nEAD96hIsnnelxz7qb641k8X8RvyAWYPpV/B6+pBDLM
ylCt3/r7ru/JndIwrBKumiF9CCxMgWgBHf2BGTt2jqdUDEpa0SLcAdvbVKzxgJOU
D7MUbLX+AJXxgU42X+Ro9fXJL6JnFZ6VItg+EUqmQtYV8nc3YsfNMuO7S//LXl6P
E7hNczHoBennF78Lgt+DKz1HXNWBNMYfwyJQEUnvEau+fn1a/tJ3Exc8vqBwWU5j
TCbsI5d7KchTbWvUgtRgnX2WKUraflPd6QvTbOW6MvnBJfFR12cs67Y/1VL06R1t
P7RrGjnWAK4eKghyWzjMlSO3aOj9dGSQT1WMRt5JrzS5+hkEm62ANkl9vciZ7H9Q
NJUd27LekniuvYVRXIToLRBV30N+VdP2oolGhj/kwRo6KKYp2rGLu/9K0nBN9ifN
jiP/XaKSM8UryrMWprzrBqpf7FHe38Sj983ML2aFGw/jQRWzvogQMicWTiUTXFZy
HKDFGbxXs+nqNa0tuysjuAD7bpdihe9/Xbl+heeDQGkDDMX/vqXy0hNMlcJ2jSum
25a7JMqq9FdIdJmqx3fKIwTlXha782HYLfWshP0JLu5UH5B7X75Hm3768X9Nmx3F
U3eFPZZKdpBVLVRqV53aHIXeAqFuj1MyzY2C1mnf8p8TKFC2Juq5mtW1P+jBumhR
RYJJcIrJP4GZfP5fIeG1EhOcLeP2ATIVqdQn1Bl4S+uUF87kPNJszk4GjJzsIV3H
5huDGVCtdEXZJgJDLPInJySX83IduW/L/LjK09UbZqgF7wVOYwxKYf6x6FNOJC7t
cA01eP2DIBTEjX24s3X0IIn924HpTfxy/90wKk7nETS3h8ZB967wOz8c9fegANp2
NTF8D9wd8J9ZgsotrdZepD4+CAayYW+hpydY+0e3hJ7OYkwP9Ogj/V2MRPfziSyM
H07larqXC762GFO3hns0hQfvf5C3Iog5M1EbNH5dEdwrCzOUi6cmyIfwRVfUQiFt
5Cm42I1nzJpEd+qzK/DaMIvkJ5Vs1Dfx+EsFhQUT8Rcj3RUGj54u58cUjzoPvrUr
BqrRwcucDqsRT9+vo3FjYEUPty6MD3ssFzR+spA84boJcFuBOAY6LoC7k0janDPQ
5uXs/66kQ1Oi5otVvqJgrXFQbswwBExbVnYzZr1Fg3DLHPrjQjDz8A48W88ZwVRv
sWPu62R4PAqdmwVtw1q0IpMM8+XQZ9XhJqoi1iT+889+MM2c3gbsThTYDQ/iVpbR
BsKP14+9f2rmnDo3IK6xYQx9uP/wo492mHvsSNYQKPANtTqk5xjRh3euB8HX5l8U
OxCWTKeHym0Vb+Se4uEe5RqvAjWgYa5ZjHnHLvRmt4pH7ynfHHXHip7Pat9fAtz+
Pu8BmcjFQ71IW3NoFmFhN+N1dolAqpf4Pgdtsbrc21ud71yktAV/2sl2OhV8yoe7
eBmlPO6e0ZOLM9QIJkpyo8Fpg0qiORZ6DCvLjOglP5TqyYYR3NqZlTYIKhNn3BKZ
x8wOZyrGZZ57Hbzq97heF3DIvo1vaX/ZwYhJei0FHmB4yY5sB9M4ON4tTnqaUopi
XbW1Jdsdt+Nd0JogK/iZEp6z0MzrPGRdWh8MqZKT4ZhnomRqqI0KCFLLWZqrh/VO
6FrOfFLvyw5kCEHMjQGZTJll9PkfKhVvd+301zCEwUAl71OK2x1rWugw80fVNd5d
LGbYxLq+AauwfwkOPtSJ97OGp+Ef05GvM9locQuhm21IY7KbLrbqWmYjQ2ThwQ6/
5vckNwq7TqvGLCSg/T7v0lzG+T5RN37FeOxuWf0hz1hbk4fAgnoW/ITLWkLuDxXD
UNIQhe/kwYl7MiyotYTcS7BOAA/l2VMb/558HD0OQinoVqfzRZwOecDzO7CxMq0x
/vORHOKkIuGQyiV0B5yKjigDxN7w8G6DERjXEb56tMKIsuB5T5fHf/lLEJlNIYAW
rUSlrzer6w1EVTeKB6+LGIR2INr+9RASJtjB1loLgdLb91f/IpZUwAW4WXjfITe9
mEGDl+NXA0XV5Pp2lueQPM+ZigGdHjCEN6ISBNWnYPNECMcTUZuLPojKQJ2Njtqt
vuLoWUx3N13xAyaXfmcC5+MjC3oCnFh6PvG9YAYUjRbJh6g63md6G/obtFrkaXeO
gOmzakJrRRv7FDWqkZ3liaJ4OXChWjUrQBCjBjKGR8SzJd7dDHzm9rUuPjMkSGUe
6HvJRiTAZoC05i3UHlZ+DlMknSk7fyl7Rb3a5UjwLRTvLsPemFVdI49P4ROJpGAm
m1Au9507SzeKt1Fx2EMGEwG9nnV5QWGJCGLT6kPLRWzqRA6lAaNMxrouj0Z2+8PC
yFbxEa6jI1k/1p0aRxXQYIg/oZWk4aUny9YluR5nlrpvML1vVjJoYygMYhXwCED9
FAALXXFBYY2zVBSQ7S3/t/QxUnkMwwFFf0mty0h7Toa6fWPYPp9bVMQfAZEps8co
uPe3mIVZNywMoOSY+EdGZDIAUhicQjeJSGZvdHtPreTfQ9aXHMDxgtbx43wmXeFY
Sjv5FM9gndtPZmKQqFEUh/pdQXsmNE2Mg6sqzNwZ64HSsFdyDUK1VbT1D8D16ADg
C9Jfs5ykMAqrCCIDK1IEcA9eGvEDucFA3x+sHfkmBPC2r6Xvh9/qhKZCDdVJiVwj
+C7+EDpQvmZD06gJSPvepIa3EfyJBQTp9z3ORlNRLzmOjiDHy+VrQ2ASi2L0f+S5
kkWbef8bU+CPCoRG1m2El4n8Hg02CHVyO5ZbZ1zmAX19etisXsLMCn2PZR5iMo1X
MdKozNX2ditrhSVKFj/RJeYpCDkkXU331iGkvNHjdMSxaGYggJ3wRhq4Nczr+h9C
F/SsZVUKMavv9UEX0if4kmbOgDgchMafGN4wxnVE9YYKiVgU0WSxITQV9rc4keZC
nIrYrSViTEb8LgHlX4HsLthN96sqtgqCA6a8fHhQ0/dXjsVmlT22rtO8mhea35y2
p2G6pr46BgklmaoVecSR8j9Qjeg5OsgQIAv7VctKB7tDuEZ2drUVxsOeWjxSLzeJ
W/fFENzNDU/9bKdGSb0OQWbVdL8Lp5UyOoGWc9Zuy8lBFn0DnVag6NUJudpYzJeG
sDe/6PtKXz8TjnxRmm871sw43f/k2AhLMWMmWSMKcyD4LK6voHqMcORNInQxCo0E
pRtJWicSMuGS0MD934hN85MRbaHUrOKMtAnX8NO0uU597YszfssdXq+WpXMCX3Xx
7MvgR0/7U/r1eU6LWMdeRX0NGeJhmQ8iMEtGVcJvDti4hMqSeKILi7k3poV27JGG
X6KK/4q9dFBOGRQkSmpfBmmoHWmHju5NeVPFO6jnWQ3okj2Ut+OdMmG6dPdquPEk
8ia3x5CqPAzpO7tVQxTUMKPxD46/uv2JEyz9rFz9BUDQdSL8WRz2MpWeU3nfk8+N
JgNbP0eEGEbUM2/gTVbatdHpZJ640uzj93oYygM72n6liNysShRzZeiYANjEdsol
refTZEVeWGpNetIRZFjePqRgJzX+2iskTZkK16vFL9tpABE5Cyz+vtghK/Wyoa2h
aQW+x+Y4jqSplhRLRQrbwd4OCvosjFvSPWEaiEVaJEkoyKfuh5S85zmWdv/qVVbJ
eFLDoeqya3sLHU+p+d8zD+9HHiG0H4lnzZ+2URwjvdV9MsPA5TN8DTPhwzU6Lqar
14c6hb2W74Wzw77G8haq1f3y7UStNsH23F1EppR/sC2jl0k27+sataCfTvAxMp0Q
keiL59mXNfu2B+GWN3w18z0KkOc/CXRcQaOdAKkP3FTpxCieHLQPq2nrueilsHvj
lbf/bNBpBvzsPTCZc6JppidVW/uJ9r7DLRaGn1aDUGWxmRdwhSbkinqJ4ogSWCRb
CSLkiD1TnE9l9/r8Lh2owN6dSyIGcMhqfSdH5PAAbmOWR6H53i5bUQ8rVPlw3wI2
HgpAs4mYwQ7KhnBk/2RQ6RouhVGN7M7z0G3m9ax8gOxKPC2jJ8h9/QJH2u5sqE91
tQfyRyO1o11JfAfndLhJ1YTJBJxVFnP/9ZekjKqdhG8zD/GVID/dODRV2p4L7dgZ
znyyLPm68oCNeaXDPc/Vr3FuoG4glKufM65Qbbu4z8ESJhFfg8vuAC41ULoMi7kD
PkdWKgtK/njcaj3b7OJYij/6qjugwywWlYcgymGeF/l2vN913dkqWO61mjHGpd5T
WHuQg+e/vjrDfqGTXIZJEYp7j86QXwuxmsSny9JUarCQ5rjqZFqJKYPnH4yYm1u8
RhHHfavNk4MZv0tx4vFTMbc77RxADaA0vcXAgzjdFK7DiyqoCLXdA5zyZLVJoHxE
s0gvIN+9UPdKQSmDA3F+YjdBWUr9vuLXAucc2hlEhEbmC1voHLGQzcMwZ9k9mZni
B05jHTGru/59GIxIKiydELlNCISgwjZUFWBTHqP99eoFT0+0Jf4MAacaIJxuMeBD
45XjFY56tC5N9kl8TYZXo6Q+oLQHeq7v8x73w384u9C7k4uIfU64A+JfOJfgZUj6
0RdyAGjZtv2lvLzOCpYOboT5v4/ROy9HRS/xcFONFrOoNfY8MC5JgQM3dIjnumOp
YcoVXft0bAze3i+QbAJ5XElrLk9EAVgpV1KMznQQjzQOGq0Eqrv+CYuuAQ7tdPsk
DjQO8IkqbjRnRTZv1CKHxy/gqhj6uZtvWsO8DNqGpaUBOIiwvKdXCDjrEMCYuxwj
den4DQw0tHZOK/ub9AooGqrVM7bESQzMV7RieqY6FU4abJNQ8Z8+bs3JUthN92v1
EaHjzjK4vMGEIyJn0DDQcPGXEcPxql8vHwDkkAulVFEuD4Tc3beK73Seb+d5ys6T
JdMof9TKnMpUrOgS1lJ/+g1w1ZI8USn8C95Obd45oCSRJ9grtYv8moM5Zd+ZuHrJ
MlzwZAe7PVR/f+YL8QkUkiUTfIFUo8m9k/bB5+omTE8qe3V/vFPyJLHLjGgQFTxz
Y+datxPpoq4ueDnaf68y+lXwoz+kkhP3IAl7RpuiaVIgFb8BzaI7tJCMHtXjcxMq
ijQyCqcKbcWQNkTyL3UhqAl6CiRBXcNfSflSom+qrNX9x0jixhMxRm/TnQR2uBL6
x6drWXz8YctzsVMugei8KkatJJtDjw7L4vqv608M7ddSncKUj3cyzGoi6q8156q8
F+T0qSxR/u3+3o3rYwY4p/PpSzsHtDFKZ6RzjfyIom3I/8n3qUc5xtxqjuldZ74o
D1Xb94k9NINAuSqN6Y4RX0Wi641iyTsbK2Ne9r7QrWs/wiWdLdLHmhTqkHn/7qo2
J4l1noQXTfJVAH/dmg9TiSVvHb1USGyNJfSIgHLwBTorucOn7NaqM3aANNvAGbRj
PxkMraYrE9fTD4s/xNB75LFqHfI6iD8SvU6JSsGzB88sudO2LgBdsuE4+DA6diHn
sAUVZgRAt4NvAQy1NcsQxULbaJDZgGx+axYhEVIqZUQ8aoEHpi9bcvlqLXAVKWqc
YmuE/dV7wvca3xCkXPCjl91GOqzE8k1UzPaBIot288rAVMAHejY6bVBl0XUpzZK2
3kA0hS0ePVkRYGNd/sXdnX69gsthYA9P6nPnwvwmVtE3QxrnrU8bzEU0KId+itj5
ojZsaS1zvfMfM7fvAkgijecju3kHjUuYVV5hActOTFpwKENAROCucThF4iTt59W2
/KqtggaQZ90hXXhj9lUUK52oUoTXTNldyNuD1kfFDLakrKc3gzyv2YoZGyafGApF
YgU08+BTIxY+9w3lGPEjjAStgXqg2WC1wcWSC4Ph4uL7hXlgYyqZAF8jVUanlUTP
wzvR0ccMfl1L7bneTXjESpFV+fBqvQrTLSbNGE2i3Eaa5ReLvbeo/TBHQnkM3CbB
pDsuSsrQA+ymqji2JjNtwvfXRRNeZq0zGJVucplPfSLXS2zJrkbPT1nq2H2yzpp9
ZqNc6gaf0FBJm19ftim3xOG8vjsaDYL2AlCneULz3nuJoo4lkq8b09U9/34kyEFv
vHVbOadSwpDw7VqjEa7BZg11LVkCPA1RZJxj/azESgUfo9jkhkqJXkSN2zevYOEz
N7O6ePwRtBi7ddSBHsu0rPhrw438fe409/VMCrZu9e+MF9njJgPsKm/Q6XBtAz+W
l9hdGkYmD9MleUpR0h7Eo7/zn5soIMiw7oC2HPEuIIi7FzdkM+YEAJvIGZU7RTJ7
PE4jmIBdYYBljALSzZoeufCDDr8Ux7p4QzeB49zg6KW0aUK3Bqr84xYuqa6La6/K
RElPTXAH5/UjK7L8SVp8OJff8YX+jqLZD9Y0m70JxqQEJd4j392vPUH+mYYot+IJ
aHd5L2UjLbdyq/WFWp9IDJAucJdORtbjsgIE1dovAtZsMKYx36uJUFWHXHn3PN5k
z/AzH32mQSj3E9ubhIWmlnp5tGFCvFgNsv8dc34P5EfpN4nUBdYFAhopI0Bwlnf4
CarEqRCRj6jX62l9za6Uok7/87jSWE7iruMI3hjpZYtHGziRsOb8M+1nuxicPjbX
leRoxQQ1trPMA0tuf4blrGxQQMpyQzA9piRq9VkhidyChmTr8DMZEkomOV71O2Pg
151j+OnpQ6DHI6CdHpzn6/eEtty66MG0J2hZMAalc8rFzctss3NYc+giM+KsAlQz
JDlahvBT6cs3onNGLvvwvA1wXqdxSDeYN+qzclpmDp1/gC5tu+bNbpr6yIT0eeZb
TpFXbfYKaojzd/x07LhUKT1bfFn4nJDRkIfgyGX40nKuvMeUhvwsAA+puAuvquBT
y8iMW2ZPbwDl+6mD+V8XOMkF267aYqqyKlYjPU3i4H9XhpoDpzoUKnX5p2dPL9ua
4ECXkL4MA0B5rt2vN6D+3sUtr4TPapDJiwmQtONslm4Ah06PQenmrHEjVp5IW9G7
uvE+jfzgfZZE+9qS/qJFEXPXSLZLMAr8F9rkuiAIDSwtkBU9/8pKbzFHr5GTDR41
jtAhpIDKVkx040tNgRJzFr43t4zOJzPlLCbjA1Pn4RL8c8g+2HjDJT9qVIzytwGt
N0iiUmEM8D6J7Fi9qSEfHFsZrNqr+r5/i7SvpJCPv8CxWGBP/prgsAqpbYK+eRE2
nejX2PKRWHxTPp0wtiTC8FcJ1Y9jDQigIsGseYltHXmJxEjhRJvVRzMh9KDZZow2
DR0vUBxqF0vI9uIy6ErWqVJ6RT8nJ1f4TpT1DLF/Mgm6M3xm/RuwJscJPNgua087
CkvZnikEd/JR58fkMxYuTYShcj7OsGzj/08Gq2TKTFPLjJJOUglDrC6LgTolthO+
ExR93Jgp5so6z65nz1ZXmNW6+i4q1K1Dsvsn4S1P42j4n6IyL4mbRwBXi+BqFQ8F
ZRRQysfj5qlOrhACXOlA/ZbCY/v0DnfAL7WgA798Bf8odwjNR6WCxaV6pm73c6Vd
uHXa9QeVkRgPmccJLKs/45alw0IH5L6PQqYEIiL5okj9G/CfnJ9UoObVT9ztdaIU
i63W6cMslj+aj8pdRYZlL4tj9Z6jUkn5Wqgj5Juy/vcOdlnSc/KL05+3/l7J5g89
VY7zFg24LKfggUM2VY6wzhgwZrYu/X+P9hA852CngzO3ZhABkp1tK1AQOb4MB+Tk
IQjgXQXLq21y6sENH7df73gHm4yke17mtHarSmArQr6uIn9tjCyoxH8N4zU+9FDd
tveeUNGBmDYGMW1k9VQtsh4K/fbdiJHdyvpNbDp67iTwSIMpRpnqw5xFLUi8hgqx
ZftR/ZzRtb44vqKDXcdFUewuY+zLMlm3Ja5arKWuyqsj2e+UhMhy4zUEL2mJ8kZ6
xWfaF/Ip3NjbGqBtLBkGYLVZXpciE0y12Xt9Wa4jw8sd/GsFxlDL+6Tc8rN7rl0X
nq/nHK3RIUEZhRAk+H020Fa8WmBImViJt/TfOF/k4/hzI3TXNgWFeoSjeBcY9LRR
T2SYs62x1gQfaEY9kIgKbjqfSWdgNA37EwhVRqJHxkL3K1IjFvX2EWf2/Uq5ZJms
S39v2/MuyPC3HQaetJoyuKnNEOQSpg2jT9lM5uKyYvROCVWJZdUFudpuM9xYssj1
PXzeVfONoaTt1iruxQ3eVaNXB7+Ba5NSy5AyeqqP615nk9GSRs5wVHEt9Oz2nyUR
vLqjuMjjfq0pM83lLGBrJ6+di1P/wDmYKGrTpdvasdgztNoUHnjcYMs2opKStP3L
LXTjlE9L+BEc41UG2geWI5yu/tyP0sddFqnZk/1EiqzHcFzIQmj7oiLQJShMEMdY
ECsmLrVPxk5IOlV24E2qUDe4Uou8GQpDK1qPL0jCnPR1LjNZBDVODL8Rcq9P2X94
4KYqpGr6/i+pMGBwJxUh8P+nDuAPLlsDsDQsx662kvES9QuTAlh3NmCu9nqdAPu4
FrqFWQaXmvHR3Hr/R6Ej6fXCe5a16s5uo54V1ZasaW3Xmyap+aKuZ8w8rWqI1+R9
U+qXY52H3RgyE6jmCcwJzEQXg+f7advIYGAE+kXlHBGCt2kF3ahj1yZykyJc7AOW
NetiQ4TKHqqepy7SVa3M4J56PiRZuyArApqQhORWHSpgXaKpqg64JYiRn9Tt/QZ7
WPP4LVqFOjNYbN61cRfjb0Z38DwJTctqTo5c/5POIEIUuKac7XBwMgwJA727a6Qf
2mBdKFkAuYmPWZA66XK2gmP650qqTWsnq8DmWEHy4R5BYelp64bJ4Rhq0RRrg7Nd
pxKhGKbpIundgQVsBvMacME9tYZdGTsqAToteMpg2FsXeh13Y5qetJcxjC4qA37q
k6idJetn4nxgbHIPv+C5C0ZVvELHw9EXHu0mawJMuI/65elufIN5yH71HA9s8S35
bNWr/iIHphgnE2VwDu0aJ1nBjdaBQpVRHw0X8oTPEuA3dGaBJDR0jkkDh+ImGc4r
gN02O8VTefLOhGXQSRSQzNvsD+4XOXjPXYv9PYG5HAa2yE4rBgWZn/WfdRTStRKt
zXXsbNxiRnxF23wRcJ4copjnXEZrJJQcKjxtvDgdj60RrZPZ541gvT1CygzUD/XF
Vv1YnZTphUN4n+aHdX15t9eX54B8aI1/N+uYxn7UXYS0hfIsiyaJ6ST5ZmxRBbuM
e+ENIPExfpwg3sj44xKfhg90C3pdcgAyAyDPJ6PUPhHun833jwIdQg+7rH/sd7rJ
7sQxUuNVfjJzpJ+2YzX2oNhdLy5/HElAYzBYUcNNBy6mPsX1zHM7s9mxX1+jzgyV
fM51OyUGERkwkXZQ/asKOJP4jacwGXynUx8nXdiZr84ocXxu9VBsScbt5dpsPjhw
um8stVg9zB2W1kGeGwTd/fpRvnb2SU/04QcsKC2vZlkX7UaUvxkFELwXzhtpdoh0
7TUtH+Oi46YBnZAP8Sdnv8Pr/Uztb8qW6+RGbdqQfad/7CZzlIo9twx5nS4h79iK
Cw+vOIDcQ7pU8pDlSvwYU38Hx0RLFkvlEM1zxU1ORoc/kKde3brkEhBlH+sbBU7w
NgSX4sopb/scSIK4+uugDBIResM3cex30/tSECbqpsPSTUuh48ZquZvYzGzBwCwr
TlRaPDgNVtkRsHVME3cHpS2+Mwjy3MUh5qpVBG8wmBwgkTadgEFH32zrbz1QjIy0
ajmGl9lvTaMAoZTjT+EHP7cdK1+GsVkmCpCF20hCZH9salbzzvs7JdsvtdsOO6vw
RgSWcUYWFIsruYIv/70e44H8KZENL3LkEjEAyDhrhSgpQH4qXMzxRTU2OE/XYhAi
GcQtCrRr0e2YyQUS83Xh0olSF5sJ2FdXtU0XQAo3udb0uTD7Q3A+zB56PzQomwEH
2fgMMj0jbeC6vthxKaOvFXlxOilI3aLI877eBoCIbBUF8neJKpV0wOV8trkyHgpy
HMlcJcCXBBiJ2j4XspwUAi2ZBU/VPE0xCyA0R0GFysTApfYI7Pvr2dj7Bi7FZ4Hg
BVihxBATKIlQDfNasiycJD+skrXdS1nLKWKS5zZa7DJJ9fkVzGS9xuZxvdpfkcjG
O1w4jy3Mv8NOJJqOt4RLhYhJxXvkP3276kyzrb7tHC2skOtYbD55Ykt5ONXEm1Fd
jxb9w2xvCaXbOePvzvqzcC1sEdcGMax8WzpT7ZCHHr963ZTk+fPxRItc83Xixkz9
SH4xwNwuduYoI4fM3Tu5KvOAlJZxArIzMHjghsQGLxGKhfPbn8j6KhiUus8Rk413
Q/Lj9eFEf7Y+8hzBFxXsiRaVYJjnS4S5UWanoVtnVh+7UglkKT5IWD+jIu2X0nDD
1+D66qxWzo//DMrK5pRjRdO2bDVcF/kVf8bSe0F1yf/oKicgtxKm0F75/n0LGgY3
3/qwGiZbBPhQJWhw+58kiJCTN+gc7nj/YfkhRB7oC2q4yUC04WyVA7DpLgtnWwkw
zFsR95mLiBalmQiapzpL/J3mWUNIpP63FklIeH2030KOXYpwGUw9romn5C5Bc1Me
THfOOUFXJvyhgIqiuZHrlyosBm1TewNesowXHVTkmsNfajttVNdN3C1STcybuheT
v7V4kkUJ+6Zw/tFDNb4lxdXCL92djiWR47gKOKwPCorXdhzAF4UiOXGJoHSbIGQw
p+EUojWbKb8J+WEDDyIZPBAR3i5nXzy9vEyStZIJN6n2bEnZlvy1plgZeb4hLle9
0Tej1ffZ+fnm/4QrHv1hHY2x1i/RAO+oGNewIIr189KauzgW8bI88UMYZzdo0o4f
6oDO+n0I9qzwP2Y9G0MOsgWorw/dJCsaZG0FVnZl6tObkcBtRcabIjEo86O2jASU
sMDAag4awMdh5Rne/syejsPLidACHUsi6k5OJlY15mU5wFI1sNN48Y1syn/aYVey
90/9O/DKoXMguZv6CBwbZOA3DyJyzoy1WekQzTR0HLDv4pd4XuqC5VI99HWEKEF+
/yArVDDqyIzURzZhN5++/+t41w6RrPn+nei0btlj3dvzksOx697ImfOc80iH9q77
bDxkzy7zc5a5aLECtGdfoj79RkP3hRchslV9DbBviz6etFJPW//RvnYsv0U/vubX
IENgG5trVB6KiSn/uAGUDPg+r6pwJHMAquhLmNEcDXkXS0bXBNE23chOFq7AG38d
byYCvY1TnnzFbNJDSi2q1QVu5iZeMy5wSnIyofdhavWChlvgsVTxRuHYjGzGptqS
SoskHA4vnFLcUls1nv2gqFZ/vBSR9C6rxeOz1TRvjY+SVvMMYLTMimxohJQ7ieSe
7NAO7YwIoy9R+YpypYQUGCmZRL9sYSSZ2QNdAd913HeAFx1vy+6ldAhWkPRzTR2J
/WW7z41wcvWK6hlR54tdZpDMj8yaxTp5+v0IXPkbXGQ/yxv7zguAjiUm1Vr8YpVR
5yOC9M6FKBQQEMAiFMD6lf1BwzKa6BvoEUETNDm0Bo6nECCoLv0m36UpQga9XogN
o3Dfq2zaJjk44DpL9nvTstwcj1dqhOA5dSspEjlzBO1yHOylYLnfDEOVdkcautV2
N+XWXr132pbKNwKSneV4fbnmMp3QIQmOasxlQaoQCntsF805xTUDPssNd97LGG/X
0pmtcCy62ASPCitup356XaLIfW7gGyeksymEUxHN8ef1OcSWD1lHVY8Kr/2h+sUc
jvpqbGHZ8L94is1rVyKlgmdyGM27fr8vGQRM9STmdYw5cV3LrYm/Qni1lAmniRSV
SdPAyvwX27yIFPle4TJEQHQ5PyH+jxGqSHnqMvuT6TXBZDD6q9Pf4wMHu4Cd8b4J
dOMGoebiIru5PC/7iLDfSbhwa5eW2kuRVkBICHgotaJx2dA46PDtHNkVt3k0H7OY
K4B9W9iNUu7Zus4n7yPmp4A3ROBqmXMCq2u04cdOamKLFNv8Ie9MknIYb3JcvUAA
X19FGvGLDcM2ZGdRfuQJH1fSbwBELK/p5ML7wmTK3orAmA0UoddFDB7kBstJYMPG
FU3luSdJn/DnfMnZ1gysFKtIDjdsN/y2xfcb2kAoSx3ioQjRx1q+UfMWR8xrr1Kx
wvsaL7TDtD1vpes6TqnduNE86vCLr4bxbPGhUCJ2O26rnGfxapOn8N6jtFd3T34c
q6b9AtCWiOLsztQSsEW5LaxU1o4UDDi0d96VsFVh6oC1+gpHMpC0eso482PNicc4
ljchmXs7yduynjKlSis0oVdQItPi2TM3CXo8FIGVRDkAHOip7o5RA/kyD9dkJRzC
x3Dh44bc1ljnTAFNZx1q+BQI1nnGWXZGkFIVa6k0NvVc/QA1qvurDr5onIL1ZWxD
QEQvj5ht1NBYKIFq1GVfPCacthua4dicAHLVoeFHK4hQ7+f+gON3+xFARXSeNqeM
SOBweufxXYzXBRQSkZ2Rouhr2dwNhq5V//mZk7mHFnf3blUF9l2J0dMIWI26t74m
VpAtmirN8Ix9QqnxYCHj8ZxPUDta8Kpb+fFiJnEqfWXvuSj50Xt/zIkHbFZSMj3F
EFj26+2hZ47RwmmdicRZ94rgUKKzJrTXpOyLkuyvwmxrKLmfCpyqf04/5ZtPxwQG
lJnn8gM6oFi4SqPfb2ljkVzr8O9qLy9PsfV4L33QCtx7Il//jWoKfoAbRP0UViuC
SYYnkTwD5/gStO1uRIh4P3tRUJtI+St5j9olqZRatp/jbgaPiCvEQJbw7k4uJ8IF
IACXZrADuMRP2t0F4p8NMyb6m1Cy5n9lSkNkiCZuEbsLl4KJcCSfP+WndLQpdEXp
BV4xrFdz2i5m9GO26SLH5hWBCvGeDYR8Jb90R4e3tDt7Z/nQdWDPHaDaQltGdwDN
qJ1c1qJoLfjdvp8A8QOnM35yXWJCk2GiROkKrFg30M6wUALu+bGHvfNzNO9FbTEq
k2MDJMfnUg60kAr91fEEabw0QICKz264jejmunC90oN9K+Tcz3Ir4jrV0+pfiPOF
JaDWT8BtTKtXpVOODx8lWeMifDMvhcJLpw/PESU3jMwT+dFO/ilY5c3AyBHkby46
72c/EWrR6Y+Brld6yMrvfo5B3Av6hG2YfWNKNd+bkoU6+P3HjX1ke8GKnLKbmrGi
oqRnbhFlEXNxlRg2uZnkqByibacNoK0CqelM+AvjzPC1AmckAbxkmfyOihbCWjQU
sf0gPMSN32KsGSFa7OOyQx0IooBz66QBJhyRdxiEkmoyz56LbGrvC1ZjvmE7fcLj
5qXEHAqcXub95ni5nOv0upu9I13z65sGfQg20xPlZO9zsJaFYCnll6xv1w9cP4Uz
PNXjr6RtH8wqILqF3XjJ/4ikuM0jvUx68Ufv3loUXrl5iN+EuUWeQK5t2ZQBubDf
eTkOVfzg9v283AC1jmYPVEGJy18j6Tt8Z/xOf25VjzRojtJKZw27WIdP4dck1UAe
9d7+s1BRrSRttemSPdogE3q3WLr65cDYe90/c1z7+NVQF6mvX8SNQJkHlEoO0+cP
5Q3K8ELmqtTs/sQTBVYm3XRjAB4dZ5MhtAXR3sZfsCgKUSxkI/oXZGUS/xDqYeXA
oxsC/8oAU6ZSiWF1az8o3CbMM28A4D0EJlCzwSoAf/i+Bdoyuh75XQSo9AlvKQeX
v/ggt4H0bRVZJadqEtJbaYOOfnUWUNckRCV/ZrIkTWr/zLMV5GSX3Y00MDU3TDGP
ZLr+1aKSNOc5G8z7+vS7LYutl/r10zvhu78Gvz7Ac8neix+kBovh0p/XefRktQHW
NcCh8ZJjK5m2ckr2+vZgwGKFvX6lL2JGFJj/0MfmcMhxTEYUW06jtR9B843id6n1
YRKRnlAiu1NmeRE5pZzuZh+F+Yzyt9pKwcc1YtJtG4oD3671PUFmz7nTaJeqCEiG
G1juTaR09rtw5LglNO8qu+wNKH5iD+JhWSKAGEQHI6wts5OmQEMbg6he315nTGr+
/B7bKrIFUqnkd+NZ86kZLFCbL7MHD66mGl5fBGKOwkWQw6yokhq2WVRM9oiJpVkB
9eK6EjAYsBB+i10x4E4YYxQIVy4I7sI5YvuODrP8IJR13FtJfc3X4YPXU6HMiIiw
HMabATSir460nq2nb8nXPLhmswA06uriydaFVYI0Atkmcid57VmRlYWEnf4weWPg
k9WZeVQLSRNLpVnmgfOu/6433l0eP1ILiCEL7S6QQf9DIZLhv6nG/7D8unZb3PVG
ATy8xqa66+mGkl/8Bd8IL7nLoyXTElNp1qximLtbW/Ucsm+19PJh+IF7w6AWH4Oc
ruhOFoKgTBboNo9EIqX9ef6qdaMGOHR1kGgGdC6HPYuFy7Wes8yNVmOdFpVZ7kkU
8f56sZ/CQl2rUbr0DjNauoMJdTN9vtcRxVyRnOlSMOjOUlL/bk15kw/iyDRG74wL
TT/CAqnb34F9ZoiX9CwIT0xOyid2goZvjPqMuY7ZOQyluZ7Y6HBPhjynk9TwlBv2
5VGApve4CICpZ957lVA7LBpHDc/Jw6tpXd5AOFrT1hgdsa93OikXSVAaIrgUydO2
CEzbGWjXBz6mWpRvvEibpYyz+MJq/M/BECNrjjoVhLt5oL9qS2ik7T1UcDgSLgtU
Vb/28GA/Mw41PJYT2aMHyIqQ5DbQst9qObOQBfpR9kGSCF8tagoZjmZWiEJJ/I9H
awI9c2N8hPHP66pcFgwlryeL1lITY2WqqzcmPoGlyALYr7/+XvtRgs3KfRHN2HYM
ftR8XWhs4BZ/rJf9s/uqObeOsCr1AzFUgA8o9hCI4v9qJo2rWwKPJhZ1nNtr3Ald
F89wB2YROcLBwAmC4gobKkyOcg5C2jJ69jregfD7vXEN9a+srXs9S6WyyCjghcnN
KaF934Nn1nX0eoRFjHJ7E48ZMESm2qI0IkqDw2m2pD3jPOUyXnJDPlvtXAZPCJXj
V2cEltO0a6I6fIB4nnU5PA3D81IWRCxGzQXcupHYFIDEUluOq6ROfdVe/ODoq86P
32chEDVV9PqQMHxIodAiTV/JPaES7uTYP+abYwxxH50Qrg3OttXLTrMJohgHBrj0
VjHEnP4vOZsdMMs4hvTJclTRtk6mpahiP+i5d9L+wC0UPGMMBr5MFBl2WPfqhbum
+4X8gdKw0bR5ftLfHPa0/Rsa859GmlN/QkI4qoFLHwD+l/QmP8ipMIU14BXrwN84
tYyNdvEd0xU/t1me8NiWfhuMUS2/lkqgyWSA8UWy40EdWY/Y0OU7AeFsQRtUzVra
8mVjSOywCcVZfN3ZpyaElKuf7XZcqwLVTUDgjj02bCfZ0CRvS+clHobrwHa8bt4m
RzlMScc+znJTlJuCiG2vsZu6EqttJYX/TuQ/3zupZe00wAQkQ1IbYgttbbQ64Rej
a1zaJqACB6R2frYHYn+GvKw18OE1DlDBBla5EZzb+IQspOgG1nwwrhMHATeOSVYn
zyb17njce2BEpTS9MXFQDMA4gYCzJqFVvOVfTV65B9lCUinY1ZsftqSvpgZg+e+7
jVp8TVY/M8J1xAt4f+PI9+EOMG5NSChYoAu+ERDj6g+Dcdagozzsb2Z/HJGUvGG4
ompenspVrbAkZ82lAuxlUpRVicf1+novGOtVhhA5Ao573cLdXnBOU+nGNpyuNMZE
5Ah9F6Ps7P6vzg4PD67c603m2uQ811dZoWfSurbAGfzxOOt1TnkVVwLbmt9MxAEQ
fuUV7HeIcFVxXuruL4xNsqx46QzD8REDU3mG9E3AfGJTYrlwpvoQZWAmgb8jqniy
zvlXCQEzQZpdV5/MiFRfGjKDUmIW2OSrYPcZKrSDQuozJh8SPTnTu6GfIZQZ4awy
gYgixtkFEk5Kty2iARYLR01V0+1cTJephMrajl0W+Ga3rdXHtnAueW7z+EDrO8oS
yfU6W9FnNfgo+uzGz/CUmSoNRTjlI0AL0YShgYOQSj4uFfXbkuPsNyUJmfFaQ6WK
o5SdtpxEKChRlb7eaE16WiXac1igUn/lumz6J5Hzlf39zpKHk98FmoCqquYEkByY
lQ7v7TqUDW7bv6Q15w9UuDoubLKB/4Gvsnd6CFZJIXnhu2V8pn0b6vSmXEydQg/b
L4rxuu0jh2MJzLZqF/75vVnJ5ok5XaTxC+CA4zUifVq01cnNgvS0Wn43G5+jtalG
q8g2ABmqAaCjcavK6mTohA3X/bkOk36LQYwFVY2b2lgBbtZD/AVzjA+W/yYAu8AE
i8IcYuEWitJ9bkasjNtP5Pm/vVyiW1CQ9CsZgaNChaqf8AElEawu3IDlcAEMEUXw
PhZ+3ElSXUOykGMLlFqWWNkgBfCQA6wt4y/XEkQJ63Hl07Hjl3f1oQVa4GZHwhy1
F4BT1nqxh+G2vpdRLGG35hXC0YwYvWj39pyQlUU+21rZNjUBwDnP2GGxpBAsiXfJ
7WQgVUDYpfmmS38safvkg0F3Kk1J28kmpINM/5pCtplDtq8OeCoqbVChqUWU/IVb
iuorv8R4fnhhn3wl5iL8Z8UuBIAbM84QYLZUkxBl9ffnq0l03vf29XNpmFXdbFbX
7RxN5vpje+5cVzglfGCVAZyG4UQ8QxJehnBNDlI21Y16yA375DTubQLzg3/sBFQj
8bRngAnWsmPHx3JWPbFjl5pvoyn0nz5IVIOHnfBBwZ65sRAbD3tw3csIGGwoK39B
8ppwNXS6p9QbMwvSoMOaV2zUq3En1weLJ430drQd6XwFVFKAcm33lRuCfd0P9Iq2
R2wPKX3Xp3W//0qBgF7BhyBg0ecEJoNmT09qINpZEtpkguN/KHeJwapEmTmareDo
bXXeYp5R1tuxQjdfzkqD1AiSbY9Vkvqji5/KhI5PNsmT5rBiUiQmPFuI4HsGWBBz
2WDSkI0W0SmslwO8MsUaNwlKTN6oVY6misbTUyiepsKScjly0b/xHbkTQo/ocyNf
cOclB2OX3w9G8kL8TYlbCPQusK9LygTek1YxqmwJc45jCL0BM47AtoSkQVPmcP3M
bUbMunlnWFmHACaVRH0XOk0tCTXSPZIi5DYPvjRgENBXZz6rVIsB0MoXBmzakR0Y
YZA+GVWpV8KtXblvY9Z48FTDd9OsFQwcj6MWJG8U0A4ra7uHklAE0vjyQwJ7pgvi
vX8a3vPJO2DoPnc6N/dw/heT3j5ahazm4UxAUxQzdXxAbTb5eDFk2iqUsYtghF76
01wsu3oW13iBezJx3L381fQWFXH0pZ3oF9dLwPgjkLOeSpDrGbRdeRctUkJD0NUt
HaBD2Bg45E3c2ZtyDFkwLuzXs0gmWbHE6C/RLvC7qXBfXIV1QhrAKXhkd5UmlQVD
6Qx+qvBQWQbHg2mfhuNzYUrucJKPsAYOA2TdiVrSJ5Xja8T6AjsYEjvKBLsTsj3t
eGHqm9AsDg0bCUWstRHu64U59x+O7SOk10MRgRCHQlP8P/G4FW7JDrOvzpzbn+wa
uHDIka7uaZun/yB8je1yXJdiM5LOa+RyaY2JpPd44lcdZGdAyoq56ub+n+tBmjAh
BP88xRDazydIYCaxJUbRsiMhzMzGMBpBQ7TkZ2NmJzVPadOYnyFuwlLTwevPL34n
m4bAzwZ1MvCKsJvr6k7mKkg8mm4gcnZgLxHOBFQu/STPlxxxLZ9h6i9myJyfE704
hFlxseexcIIp+cD6IGJHCh8JLFbuVeITF97/Ihuwo213jb2ytUDpRPt91fYIVpG9
rrVwlUHAc/HQ3Tvw8NOTOew/sX96/6RXzxVHnsoiH/9WFL3WYbSi8JicAykcZpBT
4dm43cwLtawyes8CJvWwzZMVYdvDBkaYvotkegkwScntlafZ2UCClS/ISZq7I5ON
ZqnSMPDiA/Soqf9wxiBIgCHECqiaEOnRKhcQpCt6F4li+7on68oHWGJnXQKdA9A2
hNuEcvgThnUmq9I4M/QixHi4xPftaOCxGYk+z4kVhEelg1evChB/dCDjB8wfugqt
Nz3uKUoyLXmF07FgdXU263Y/aVGns46jt2v6TQ8zZaLrn/2tPOfaZa6LXTUFAP18
L8a25h2Z+JbOlyNjr4HU60A0Re8guwHTGiEk/usWOSKHQA7jFOdOUljUxVdC5Z55
n9achoK9io/lgs2B7XXl0jpHivkbV1PRT+vbmBObvrMBxZiFRoiKFKoktkvZFHGv
jSaOSK6e2oVn6Wl33TLgvogm2XjYt+ZG4raAwUtcfiCY4Cgo745u3jpfy6oDJEtb
JJEeimx6YVILoi2Krfku2X5bXVCO0u4nVoDhTQbEeoTmEeqj0CcxhJq5yUJqMKlY
P+YzOXcH8lk76ujOtpvsAQrbgQFbTcJM//3ZK7FSCW43XeJfFEzaUf2B33mRWFGD
c+KVaskk0IOtlMWkILv8TUbX/QN/8iyTNdbY0K1yv8ooFjFqxHxnYwsfsxVVExoO
FF13u+Wo5J8N/WvEu3enOzVdNjycwQuaihIz3GccZbcvzNKQBkRUDeJtRsClO+wH
bPH10Yx2KsUfD5xeSjIlm4J4TLP3J/8MpSYe2Igs/GzGHV9hd4T/7oOezKCWf1yg
JQrbQUow3immKvYnhS2Uh/6Oww1UfiAHYKNcM/hSo6kK8QvoZVfBGlGjOfPoFbaI
UPFYDzghFI2Q3vcISTkYFpirkHYDAfxTx6RU+mJT21ticuhMyjYbrYLgXhPZ3c4N
F75V0Si8+QqIjNOPmnqQYgAFVxt55pU3+xSpHT3+T8W4+k2nQA86dxXQIUGER4bY
76dQjO+t6ySwm2yQyz3FJEREpZe8ejN9m2EPSKey/zMh6dsiCCf4N0Pm83rxYsqA
jkn3sVkq/Mpfd8g+I2zvDSs0M6WqxEbFPJ/K8Dt2ocj48zZyFzCs39lOsD7uILcW
aG95Re0IjLplTiNqyKyOTc9YHfozJyj11kL3ONgfRft6Yr2o6kZv13orgup3tVoq
/HbFEFGJm0nM2wbLwzJCJVzVVUFqkePARlv8KXpDNGPquvg2oSKnfZymR+dvFZ/d
WdlrHomgnC6nKVD4u43scmezgDqhhovexTJ0zzBiK4PFXquL/Z14vNK89ad1KBg5
I04FILsXiAhnU8FlQEiDVCxY+arybe/OhiuLQT8aezI5d6B3qyJM5zucx19GM7g4
rZOzwfQTV4k3jvoSPTbC/owEjx8p6c0Y17R6AVpl3AF1/2LaB8bQJEb2av7ZOroa
tM1RiIR49DpOyb4EtKXBxJVn2thOZwxmd2B70qYxNo3m+3qap4YEuSQdg2ln8oQV
lWz41dWL+ca7PGITB+K127W+eaLU36hqe7lMfhPYeee7E59bwhJOg88tKLXlydAo
A5acRkdoHp24NhKKFr0nfGi7irXXtXlXGn6fkf5+Z0HxvOXiOzpUtsGWIQfZ+iYg
0iBCpVlH8yRCKCUa7J+wLtQFCmiV+2u9SEFk48lFD8aibCtTUqFNeQzgGsNKEwr6
ulaBJf1l+tTt9fJobEdvkxBuvAVDLOjpYRr8iwy+5KzPruk8RE/aEbQ83BYEM8yR
SGzflCzIBAMDXu/tK5+Uz4UrwsZEx3r92V1FXEHEkP7vHnQ1UW7M++kkVhdpLqDR
QlioNJJqmuni7uczU1/m/SNh2KD/CWNgeMftYYtGPpLy+YK1krKOzaywnVyS+7Iw
RdQqYAq6DQNgVsffGzSYOi47pn96Ld4J7/7jQobMr70WopyFDPr3o4OlWkIk7eXL
sXllJv5uwhwzkm61+CrjEarA5SOL2xiCUjaTvt7NENBVMxcAIJyqSMCRwjDHTurw
lSgm4DRiSont1yq8lwcuuv07vr7dyxHC+fpiGwEns4VhKqGs2u5nQjWNiyijQWbn
zsID8LV0X0vVSRmWNBXbpMwiHZzLcOqXCFH/Sj0is2MPerwugc3N4WWkCH3rxko1
bXIPPJcWVCMGFg3g1K5g3gtj5nAmA6uUvkZClZ8lWqZOsyCqQHRZc7z/rrTveh0d
RS3a5bPSvFnCVqq/RD1Esvo6w6CTvyVwhHeXAJzAllJyltaNqJMSHdCyQpUWYhfS
FBxkMgM4Q1sCfObaXCj1hgzpXRR6Jyj/BsFKMKommK1kW7a47SvUrxpFSs+XWspC
cg9kspGMKk5qk4ukpXTsx2Gt0TNGaenzk+797NCsOkWSuatWSFN0rgKwa9Djt2zt
cOSheVUra408d7oKgPXStWJTuBWex4hhQjPyThg4Rt+Y8n21nndtFi4pq2lJYwaR
9OFs0sCSXmlqJtluHPLrrfrJ04Y4+rsfjPLXY9MwRFBLilezQb9bmhjraw8jAVGF
WSXqenGY8GleFDceBD5Fij9JORXn25BfyQ30M9hpinyfj7aqlqipN7h2wJPj5HNS
uUTMhceH29qQYwt/1bi4eKnh6jEYhN9pHTxWHzRjaXegx6FlsAkKqzsccHSPlJtN
F6BSzVqgmjmAYQZIj8HUK4obnbhZAvOB8dO9CAYMgrqzetO6SXQ3EiDmVhyK6o8H
L/HYejTVsuJ9Ox/i9Bfs0qim4ohDrmQxWIVDPqXinx+ltueARG4g63ZARlWK97Oc
qhlSn3WJKlWIppGoy1HWTpdgnDB3NTmnY3iZH+T0J4UgBB0zem7yak9Jiuo5Wkso
403Rdoe6Qw1NIbLikzAxB/EcB8fLjZmmagRH4L0ae/LZ9t8MLZoLkl4Z//e8/970
zkEUSWVa5UNNXb8xKheRquGB8ERNjI9ycRR1X7CujHmq/l8ZPTq9vPLeGhDX5mnJ
L/bOk/2kMIOm9Pn7MYTLUI9/vVWqkWNz30db0MzEexO6lUReNdlEiLT7n5YtvNdD
VLnSlGW3o0p/iUcz2mZwSrAqsA5asZynB0yaCBi3xeso0TH97wb4wuLFGWImN5V0
raKxrEInmXNA1J05lGBZCpgusVq1fPau0F1GQgQNvHEpg653u4JAfLhBfw7CPz1S
gOmddv6wgROM20oO2EHdXMvlVPRTeh9JLBdZMV7Ug8NtTZ/+9FLjQ8kH+u//mvDp
P0kA/sNk66pYVk+yrHUhVhq0SPzlLQm9CuVxi+CpR5Pe1wvQR10wmhV+brJabxHY
v9YHFr2kN+vgXkIlcW/xOaQezvzKYjVZ1woCkRm+u9yA3OpcyG9/fuERayrxuM4V
fdKFO4Es+qd37Vh/5W/ib8tpejMytZDmDk2cexcSGC78Nm3Ie2YGwPlFCSga/Xjd
0VLO4iIN1xLtwb395uLAOPgT24b2tY4GFz+hr7pGq2adZUuOujMzafiX/YVszGLC
K3srHph9+QPzh4NTZci6yMwGFrxkO0tQFqjke3YxKnfn13FW59R13eJqGo/2QnDn
Ii2M2TEPwb1UkV0am/eFXPCJSEQUNHO2dSJd51fLOUaL+RGu41kCvtCFyZxJytAk
rmVYOGSfBGVFGX9Sf8qGEiOGbnLQIc1S7HBwH5xnIqNGT1YB3JoXfjZfkbxrpYu4
eSlaLltSdpuggAxsE9ZBkeRLBLKaLc8mTyUyOh107f1LiXQfaDCHNtKYJy5uFpKh
VQZrzrUKBCEUF2o6q0UUhyOQJinLY8lH3UmmZ91opT3eSirXhYQAwsEo/oq0RorS
ijMda6rXoXr9CPmQE9yvCinZ54ysLssvZFOAdhTP7mCy4SsRa0zgudDJla8qRaQW
XIVxGHwkHf98Kxqn6oN+Qw/6nlO105SpIjxodMX9D+qS8f9OJmYOCM33zpYQjR5+
kXKeWfpMhup8ExyFAprEDiX6pCxxJmt5UIUp7TziZ43UfAkoZB3/DIqmnS6tqRwH
r3BAeMyVWk6E9CJYoI+H3zliMIVoJitKb0+68lWsMNejsnwh2UlwD8RxkF2DGlya
BgnCVDnuhFuLXHHq+FA2rXVv+RXNMYIbd50fbTUbTFfhvaAUq8vkLdXfYnXBd4gj
XDVQ+/SE8+WU0+UHrdLhxXacciSSja1X6Z4eg1wYN/FmSa0pMDXkDR7uZfQv0ACN
cvTyGdwIKLozTAXm6AFZCk3P5UYFiept89RpAztiIrcRZIar4ILcFjnbC2d/RkhJ
I2ZHJaovQge/1bXpG7/DzBUm72CEQ+b+j67wQvi32QIKQr7VdZDXGFpOF0X5Myho
pc8vpnfJ3QkS8/WjuDYj3PbDhUyfiBGlHQLNva40+Of6WSOFDsclc0Spc6WhjOvt
mALJwD9WhH0WjFNksd1elJ4qYuIb+BP8/sslWoI042SRa2ROfqSNCNsZw72FZiVS
SYt/qX5iWKLVPbab8l1SMbQzwRPIjJ6jP25qnpHOMeQw5tREB5LgCXsHP2SIGVQt
b7+a5k6tpQ3vTL/U5pGBrQKBJN+hVcGdU50V8kef/4PMKzCYgd0VrN9kpU9S524A
fRnZvOo8UGPByRI8GvrsrQSVXnrKE3k/LGk/b4IrQadK8GSDC5OsBP1ALMY/uLjl
reowbrxJPJogKLFxLiVypbnDizK9EbB0EGHXVaoyhDzdEZqvgd6AgiQviV/my9Vm
YpBjXz/EyC60OyA3FYM3c4WxW+x6e3coai5Oty+4P4czp3nnfEg3fitN+tj7aBHi
NLHrVu9vvzGHBHSgQ/4hExvDtTWrdBFRDpeFx0Fpd2q48BIhK6Jy+Be39ER/uDZb
2vsvVDFOzQVvFUJq1P0dNct6rCngHmCE/gUUs9gov7HNPgGQemsMokahxp89S9Bs
d2NS5aWCf5KTANlYU404Rv0NRKxxjKh2EC1PnUKPE60CYSzb9Ai8jOmEfPiRh0ac
VosKUralaq6bpsdNYrcpk/Hbo+xYpq6uPnMkdiQLBngz+TGzhqj1F9NjEC6okVIJ
rH7ar/VWIKVAKO5E6HPRc6hnl70pvcY1Kqyg3FIzOlm53B5Pcq3B7prC+tPHSYTC
7O5CVCTQuZ+3KkwvC1JAC7B9BrTs0v4Pn4ux/L0yPTuSR3VZtT5ER9bmOFElKkci
Yhp5jUpog8PpmIW9cIr+bavp32miGWSb6dOamI6FD63dp5by4X6FCDaf3/3tXZxE
08AvjyQ4fCrpxxf9/DnrBVM1ZPzANUEAYI4+4CwP0WVgZ9U4bM1S1w4htGi7fI02
yORH6vpR1ZUbAhbu22BPch31V4U48HDXcxJAer5Ty2Rev5iMhy0kk0Lz72L6xTel
PYvCgBLzlhyPvDBhpJFFXtDTK03dEIbF1Q/J2BlsX7F+y7s5eZeFE+IYXKLCF/P4
PnnryQ0RXkwL7uZ3R3iQ5PeDlOOuh1LzpdBQZP0KebGyrk0pTyftijQUKgRbofok
XtRNyUpUM5dn9lG7ozP4BLZWKblEDoxxg7yoionL3WuRcje2ZpDaxjXSiLI/nSvL
vlL2Izu9N+vUm5U+moRaO1BbC+2FJ0suieWQCNTN7MOO2/uORpK1hg6jZdqn/yt5
hu76RKiJx6ozsvdYaqgaAc67CusvED1OKNgg/AzqXKYmA9XKGQNETXnDembSaB4+
cCD7jygsN6b2Iee0qVKtlQFYV70PuoBC9QGZZfGrpes0OUVvyQQ1udu0/Bzzq/eT
dbfuyUBRnPvwNjpn0e+E18M4BeB3tQ63Sn0golQ67skiFJjWOaeNlGwnpa1deaYt
YIxXo41JnVChQeao28hPUV5BeX12IT3SZywSX3dRSMqwVX0lq6YBRZ3nhyKbgj2j
mng1ww9xrqVhzF15JoyemH4LqBzz8CXtU4c22yA1E4+GZVj97W5AYHzoSJeYnwGP
v+8lDElEh4q+DszWI1xJO4LucFrtOVquKJTPKigrzo2NoBpLvnnVk8x0Rm+m/cL9
ubCjMHecxAv2MO9TjwMmQvIwNKsZI6i2fCwvZMw3j6ROelNQlyXzqESBXEUwFGik
zEkdefmYdvvQg6hcyU6HqBqw6UgvV2/2DTylx1aCYvxKf51pxfvKzvwum0fL4lT8
ujykRallEn1JiBymQaIeDCCh0nV1fE/uyzQsM7btnCe3Vfk58x51SAecA6Itv3nm
J9S3gqB99D/JFHr7EwOvCw1lAHCT1WkGhdRBvaAiS+4nVtFejm6DCE6JRV0TJwve
ElgvsO6FiHmvsZmTtatZqBHNhNYpfiiEIOyOOTgFy7faaZBeMNXZteyDFYto31sf
z7kd/bb8KtKWqqP3uI5oRelP+8Gnsrp7CaZVP0kCjMgyYmPI0UVLx9iApVfg1VMq
tHi+B3/py09IUWI3obFtCwGhEnx4PFX5WpJwST3fHUImHlPFbrHjaYAtAzB7R+yP
8qWVtIUZj9letz1eLPEevl+pN8L3QkPHFr8rNnjejS3SrtNnMib9Jta6KdonXqUa
37qEstO+5vyij94epLjTYkixHj8slT656Jxc+iVqm2MUiU2Gth+TUP/U2w6jAlc9
xpsKb+SBlmYpiC6j7emgy/R8oCka/Ii64tqroqPmEnlsUbYAKOhG7D2fvWLECKYg
wdvk8D6p645IIsssrtpAjENe15fCvG910mnuJAThqqqdUVRCY0NLS57zXSAcjE/A
3504d7ObOTCGMD2M6TvI8qh8/EW4WewDEpgHjk8gH9kNpIb3fK4WgpZrxQqTg8MQ
ZweaSG0rTXb/g035NWZcUyrsDS/CaHe57i6EzEUHWUQKYAbQQm6SdndmJ3yEsc5H
o1PYd7flqk65NB1yEwd4GCg8DqL9pQugFoH9IRt31M34vjNe23lie6vHtsZNcrQ4
BHkp5Ko0Xr7pTBEOheX1sdqOi+AWJrctcnaL2HZcehCfFpz81Dcrl54F715HSciP
84TzS1YWG1QNFisxCTQ0+oRJNiHJjQ0u9AVk3hpeuKPK4lT4ggF/vGR8ZLjiucQh
3g0FIOCo6JGftITMT3LJUHIrrb51lZLNC63SNGc4F/Ys7+2lNXRlLAwV5pcrlrB8
oEz35YTWT7AxJaKrjHu3jbx+gI7p8W2iBm3y4ovilu2rT78tDFFlPiUGY1dJXGwE
/QXDPq1HNslfzlAyk5Nz1FDnIrCkn5MXVgAepH8cYqJ/vFV7/mOcUySIo0NPB/WK
C+HvxlMC1zL3TvGvoI6kyGot1lrVgzxNeWhU1eT+bimO65sUgPAi44+FokYfJISQ
BISkmiNLBqDiimMXj96yHtf1zldEAyzIY5Bv8x74wiDTMpOH/tU6J0bIQfd+TvyM
V+ek98F+OVUPdcjgw1hopGn1APqFxi9qdZ0Ru/h1lCqXBjINWWOaDns3g0LpBKbJ
YPU/xzzWhiZRH9aC1Q9aVbaPolqHTGnA3gEJoqZ1dBhwFMo0Q9K/vtEQAf2b4NYc
BblNmSajaypDw64PQbpPyffDJpdtwSbkYBznYrmWjC4fbtM0jiLOD8grDlKeCW/7
pHNZbHWTwXSCst9X6q2QkuqnNAU2dj55ChiTZ3Iagc/Av5xx6HuecdvPpMvGFSYo
3LjiM328bSOcAVmBQ6vrB2UDk+VSKo4CHGWk9g9CijjnM+in9wpKXDxbY83s6AfS
vqQ9zgXkq6qCHQ0Xg6aZ6u9QH3c6Lhpx/Ci4641kHrxvLgtyuWZsSssEj1gVMBoe
pF/UIBS3xz+7FipkGGlsh7mIb1f4eBEvD0arNzZ4OfAji4XIN+sjaWzj89amNHC+
QD2cXBjFB1ShoFFVfYyV0sNWHyYcm3+Pv65W1Trh+Y4LIL/KRAJDtv6HXN/GZ4DZ
g43td2CCFgjH35VI9og7OO6XqHt4yXYh+U4UIQf8ddPtfrwQfxXgr69OO2GgWAg4
zt88bflLHiiGFBi7WXHl0K6pOxoSbF1P4dQYRrO5jnnRYHTK8WFM1SpNVAajdMFS
wTkSgfaIXIF/5pOfgTrV+ptORtdLRIvW4v4jIl5u2p0x3q9d4rlovy9MmTM6g7qX
bMBtrmq+Ta2RfIMl3+sjFMa56VOiT7Y03N2qMO9crrmxBht9wGjtvlhpyT692Ipb
6UDLKPdvAEZWOlxVj76DOEjbjMHWJ6UVkyXn5On5fcQgJpbyjWfXMRIrds6Lq7CN
1hVAIso3vhCoDe3lJNH3gTWr+zYpntHdwuiAp1qldha8dl5iOzgshs1E4N70j12f
9u37WwDMJUsFwFQaMok8e/C4XAEmBG4PwT+UOd2j1wZETi0r3GOPsSki1UVQVWeZ
ktV6ckfYBvLX+FuKEFLUkjIgvbSFFO6mZJoIeJ/bGtzf1btVv1xfzSxTu7vnCUXC
qEY+HfwfHkQudpSNNukuLwRtxV2gvCmY240uo4OR1kSJuR9Lh0nQv926YpJEz1lC
EvYE5wD3JuW3QJlcAmUcSRNmJ6PV4TmO/ba4brdQ9XsAa/dNQfyubNUHob5Nn02i
eifASJQME3426fQSCOD5nvK3QvZ9snqhfR1onmZfzvyMmdCvbDL/fvi7hzZHrL+4
59xgJJJuZh4cAJ/XA0tDRMof9WrCy154oqNdEtwYybfVcJKEnZPA+zM60RkpOQk9
zHNqW2kAT+aKBs/sRr7vHyhf2sFVOTu0tgtwS11z31ljMZ/pUV2rX1J61tNKnt5l
KYkY9ypiV83yxn+XfIZBtcRJbE3H68gEs5Xmzs3rfc0r4zE3M2lmwxOifoVL96yR
OfbM1UXgoIwDvgQD1oKGy1q6ZPwQI047qF62Af8lPcewkWowNRlgSQkR1UDZ26sy
AGWdG3SAQu+fD1g54TSANTzWtQd8vf2A91G0H+11jXY0udAI4Dgbrk6nG/ngQ6bX
8ph5S7PDaP5EFh8gzgQZiRQD5AcNms7J9W9T0OT/JD4hmXX2o5gXM4z8St7NxZwr
U5VrXOOlMhjspM/9Mc6jjgBGuVT1DIO8zVld6NfTaIS9gpOHOSYMcMhKZI8muoBY
QN13a3l122D/Uj5vV6SOAAUpHyF7WOgHNSSTojknSNgNTPUNealblI35ZsL4cj5x
E8Cl1KrJ4w1ASU97/TToVU0MK/n4zYeX7YytowxvVh6OqpOu+pHLdruINzzYegrR
Q+tEwkEfyE4mBZohxUB+HbAlZ+tgcCHe4xagdCIIVlQpdj6Sp2Sg35Ezr3SkP7rv
CxMOfQ38zmbOqXfAvIUogVDjQy0gd76k1sRas+K6wsgtShUlVtoP2xZY6aSJS0cM
uzbXlIaUapvKTwOPVtIESsDOHoAPTwcngU6Y+j11MV/oQ7ezsADXlHTK4kCPBWGD
Ls9+afR9HEQNhcq1hnkiPO1U3TitNw+kB73ZDeVQyqWdkssgaPsKGc746L6RzILq
5d9DPActA19KLEtR2r0qUK2ZJ8ktJo5t1m/l5NRSWatjKHKyJMMoazAGcMfHlifd
oGbogv66/gC/d1g29ykCa+mZ4QndaZtXJXuCo3a0cnqFHz2hl78egpQ4Ao7sgSjE
upLAHlwO38iF+4esMFaXhpHNRp4O460nIU+9B1Hb5kJspoiXOcTY0abX3TknMACk
9DFF3/XaT8nyGhzmOv3uRLksPhDl4jHepmBEtGxte59MEzyhvJFPPIbpf7KV9oEF
MP+gjMOpK+vPwzqDd6NVhJ9v2AsL6Ivh5lMCkfO0gkLltgQWDFSa1q5+Ux24ODCQ
9yNwqoDYGndXPcmxCHh4RLt/g2QAC/wCR2uogbFUk7cGxLr8k6AJekgzvRuba8x5
0K4DD4yaxayzzIvGt4x13FdvLzyKpCya+DQdOBcB5z85DtuhDqbtjJuag2JlNsV/
axN952dK5p5cNmpnZEU3akwTcYA9ihxPChc2JHGZ54YEF1xAHR3iBoB1ZAKGoBxT
3P9T5XZgAxGIL7dicLtgSpkaZ75VNYqpAtVLn0wSRrOAfHxfJqVjnmCXtdjXWeBA
TytqKl37h1RJPWgV0maWEh+lrYwFSkBo89LbGRUv7jw6muEJu++tbbdqDBeB4X9E
9Y+5rTN5vJYIs8lbgsi3df0/oHiIxQVizWvYem8IL05woiYedoXFXamx0bieUaQ0
wPsX5a1efrQTDmAjsnn3bba2bxIBhzlsf5V8WU70DBTnqVfbSPwRYJlFArIpJ0sy
HwL3ot/SGF1vMg+jqRTwLNKgD9J6aQDv2lBA9U3HfqBwmmU6nMbVXSczmuCO07Vm
jROTDsfJPZ/cSsHJS2ZHtpd0VczVZA95NjhHw/hZL3+aBrTQlJhcxDK6A5rREVC4
vDgmG5eU68JJ5Fo0QULCWQqvp0qiOvsFb4YXDpMA9/0ifarlIxn4x9kWvgMLVKAZ
swEx7hNDzdJModYQuY21vnRzcxmDLb8BF7DX3q6qKFTwzKaZJdXh2dtfJ8ovj3am
CBAtG1e9wROAzbrspFtbNDAtWwaTXHnU1gQvbQiC7MuCfcaQFjaPmedXxNSr9BPC
DXEctcL729prNMK6dj2pm87/LbZDSUyKrTQ74QojQVR7z4RHmRacI4HzlT0Nm2NR
HGVq2dPtckdxrZpyhQLCrtHFAdx5+CFn+SVpsOaBVLCNke06us7u73YOL7R5dM8+
q5Hjq8vUqyPvt4mp/55OUthQTnsC/cwz6u3AWvJbcg8c/msfjg3K7whg1uRWehmT
6lk0d21r99cdUYJsWh1Fcvpkd6b2xa6W/twaqma9I5nziKU9CZwl63GgKBsVEzLd
Naq69iKOkfZBg4KArAxndYhFnijo2Hlg8/pcOnlwuqdA6Sv96/zxPhLWOUJQcRvj
blqSWhvlAKEicMqvHB2rFKjLUzwndBsUFVnRmCymAD7ugCVgnc/aCDhWLfca0REj
48RJLifUEePM53K4SzXkBf46Olsymos4n4bEBE3glskMaa61QcW3Hk3/2KY2K5YP
OSbtjmK6U6rr6MaDK3AZNlvmUir4PF4Qq/0vzQ0WhqK+240CQorlq33uw69uzHkT
BWJ9MNk3cwV6L/qge13Hz09yl+R7qRHD4LuepEPfX32Q8TIVjSI5HYdHhXf5PxOC
yT58Bfy/2LU/nT14ltfJ6zRgKtCV+5zNAiJfaBSxOOBe2DQJ8UF7lsXpA5esFbbF
PZbRwIOZRNFjHbjXvTbDae4p8xQE9qu8hd5NHgXOq8w317haX9UWBmRiOee3MYYW
bRpEo9CIxeV+QLHdTpPjWHAGO650Q+8uDeQNtD9KdTnC9VX+VBWtb1cV/K813JfE
HdATEbDNhN3ub9H9aJrGBnhVZi9OrHyVr8uQj8WLAYIRAMGj2nWqEF4COgeMgXop
ubZaXFB4xmHPKdvvmyRbdevjCAH2ZeogmynbzlcQpVF2BNcKt1ymdcw2dSzBbChN
M9Au7RK3ELqCiiIT2/j6TsI+6aCBYLY8dGszEJMTkqML5H3NAG1ENuSeMnbrqMKm
xyCUFN5PzGhcJf+q+x3DdAAfLlbpXAdbsgWryg7XEF7t72DBDElwNSGWeNV/uJMp
YrDq55m/sL2ez0URD/3VpF4qs0/q4AYrq6rTBs3p3wb4XIiLbJyHtOwciTGHaswu
BLDJ6YuJneN2EQ9Kzky+LMT+uh6nMu62xrBB0vjfRKJVuojgO2Q7dfPfkzn+lvi8
3hukaYj7410AJiU0jzsiLjOc3FKXtagm9qmOXU+q852uGcyZYCp20oCxmv7boq9C
+GDORAa6b88Ca2vBWCHMKQ1o56pRN9p+fAYJxsWpod/fhHnKuCnxk8ZiNQNTmilE
Zz/RPcG6zYbU0jivRgwgPi35W0ENfgMfkuGgd+1A6co/PwQsyyYagm/E769Efx7l
j/Y26fmuYoL/qxXwN/mwYcz1+OlNFPMNlKmVLvSsxE+wUm/53x9JZQ/aBzcvSJe1
m+J9ZsmnamvsFpInzH8n9BpfvLOxVI8fk5DC/ZhrDN7PaW3qvk6Y3Q4EVYmkMW1D
fYOhQriPdX8EpP6+OwR6RurZZ+wwsrL2liA9WIVmkYCJhLR3+CS0X/o3EcrnWsTI
RZ4no64YRk8/gnXsMUnDlZ0+opXc08NCWNgdjAvulVSp1vqAWdhpgQ1WiC3s8BEk
WMNhl7KQHI7vRhJa+gyQhBzd569khuk6iA8DHwZQ6OHYEJtYCjYRe7oQjypz1qEN
y4HYDIzTOClcxnES1hcAbxzpQjYJmNL5msQhdIOlYIkGpLRmHhtzNWFn1Cz/+WhN
Zgrbt9m6VXp5ykHQpVA5WkQVg183uvCD0lHzUXoiSmo4NU7fGl0ArqlghAp2dQKh
5ovAFZmbxvNdmVG3aMD1lztaM9BTeifA/De8K3ya8gyiqA1Ax6xFhsT9GccMle1o
McrfUqabMWoN3+xXw4KDSU+ozVeLsnmd7H/jZ/Kzi3epbU56JvYTq6ALQTYdjQIR
c2fOvQMQX0tb/rdLU1zCtj8/9K3Uh07yyiuaxjRAUE0mWlKAHgSV8zM+KOPLLvxl
rfDgH7Thiq4CK+RBfsTfAyyln4EFoDQf92XyeEbI2AXxy0mBpzBFuf2qSak8p8V9
F9Tvapq2tAf/ateI1SPZZhkJk1gpuhYNfo0WsYvyeQLw1EAHnhksCQU0Dfl1WrH1
nQBWY/Lap3wqf3ePrnJwITImVKjN2xpcq33xapO84rauCG5Swg20UwoUhNmU4gsO
JXjx9wGb2Ea+0tUOQDhRllT1jLlEl//nqIEYbxfposCFDkTMVdGtN72ZcsJBs9af
oeDevUTbG6IXc6S8CNaHUbqPTg67d4EmW6rdD88yDLTplwdabMnqYcquGX8zLQXh
YrWDDFfZ6CsZWOcDLWsPLDYjP3Jw5iAtVHTzmwnkD0enSqAfTQMfpZ5g2wVDPhOM
ImYg3BIakCjdRV4gd2nhXOcRJbdEzf798aue/MJmo++us5/ipuJqdVs0f7N/vmuz
f0DMNoGPKfXVWa4VrJp7U5w7yzAvlRW7OHJhUXnHKI3eHRkb914B8S1I3yed0fMj
1ER/mNKLvsU0hIwK01zgRxKkJ2tQPFvLkr/T9q7BUOVIsV4WUrS+CkvZat7k92sD
PtNf2zP50rICBHHTkwMVaHglNUWidvGlmQiL1MreLSkrvvD4j/CP/2xmkrJvsZED
7RT/1lpx0s5+qYp7/j6GG3LxN98geHS2C1Ep3VhfCXjEfwc4Rg7Zt/3poHcMcTZH
sR4PJWEzqXUfh3hnevncDkf+0B/ytoRypfL363flg2iSOt3F8i3koIPiDU1x082X
MqJkIhh9t0K0CS/LqkjiEbVOuMsyf8nHW/rAIIONwvEyE4s8r4ukK+9u9raF5kH3
ctQ8XOMq+wncc7DKWjH6HzCRxFTIN6kz9dqnfOLK6FDmkXjO4Oz8ehpe54zZXtZ5
Ma/8VQF10RUnqGbK3KBF2wIas0WEeU4TqZxlNFO934V4GWErY9YygyKbRctT6FT8
2j3TaIpehnczSFLzuP3r5sVTbyaMwG9w9N/mIbABXQcDFlPk6YVOq916bOMc+cFK
NnnjarFiuk0I9lHGTVP9Xc17pTCuUqldHx2O7c7QwywLlwfj3DMwuo1ZH8j0M9bn
6lJO8e/7SZVcfKbCX944PLrhKIZV4zCIPnr6MhU4AmS+nJfBK8HAG7XxcsqZMeke
1YRVIgGgUW6Xqbdm+xvPRMhWXfbhX1eH225bbHQtQ84Wwqh8TNqWQ7rl81fTAMMb
MzfgFccqYWDw1TApDs9Et9tV2+xkipGx6rbhW9Vr0kPhEVV33CmZZlRaChkAMK9i
GvyVEr8tCcWQoYVgG8ysXtNf24K6a33sIIBf3T9N7Fru9UA0H9JGKsAM/crMxRf2
oIER90sHvfNAvV1yPrzYdHwMjlPX1Q/ppwJdxZHUTaKCOhHa7lYOi3PI8PUxjPKo
AEl2clpc48Ljz/W8pbV6lnlyGG/VXJCv+abqecbXmJ9jCf5uXKmsapg6S9angxIp
tYEfmoUYmdg8nh/zkYQkI3BGlJRazUkJGWRU5gnpd+mVb+tOH+NX4ciIFZbTwLJZ
/Jkqaut7Gmvom6lTRfWC4dJYf8lpLMKRduldS/+vrUDJGSxAwPeLdr4bxFfMrlMs
Gv+hZvWMAAPO73ng9SEpwJVsln7quC3aNm1xUHGA263ZHNVshbQoYxjhm7HHiDOz
50bb69OBOdf/KCQobrxlyzWBUpMA9gGtI9r5JIyrCZtIJ9QC8GQefU8toijoiCpl
UIQb/zr9ZKsm/OUdEVC5N/1mtG3bkrUrXIbRtaf40tfOuXVRtGtf6zHSHeOrKMly
qmjgWFpEbE11lv+eE5NmHq/4+t1lcu69KjfseMgoCJxLO3+jokk/Q8iaP8HE+vJn
4VRcFZk8kt3mEcy87+C6MVbucCjwEW0BlE7sTxvKhxeEfllhQIppIjsqkgMbl/Bv
mc7ANNfzKIpjHHkbY21UfHid42vl/jE0oIVg0W2rKLp+lC8dhx3mP2pPjXO2CUGR
FFjQqxf6ytA5gMSUdth38jf5yh/7xz+70IAmqzQ7SrpFKzbroM31suyxfNcbZ2zR
vVn8tClHmt4bTy6qUeIztRQqURgrBR0F44zj+bRmohMbzxsnnB4qPKa1nuILEkYs
S0Klacof36Z8FfeIHJkCXwqMFy7C/g6wpPMIWM4VEwvOrTI0LLbf5AnHRYgy3Y/d
4MT/kP4sWpXauEbJ9NiNUaFt+pBIGFCovQ0BNS3h6/XdGUScnGhTMQy/PiY+edb9
gXpjSt/qXXOEv+YrmBAHP/ke3cB7GLX8YWh3LXWn7n82/z2LBZqjN/jbQmHlInjj
bKRPjmaDiGIzbpkmb8a/7fLmN/k+NUrAPPzTLySUfk+TCJfoZT/o8fh2B9XjmVGU
fKGuu8EirfmT4ND7FOUla18rwte3gAXQoLWNSV4iOwIK5Bh5GpkpXx4GirVqFUzp
WERY5Ckh8JYJ4NbybppR1x1zGvNCNTc1m5SYY80Uaxr6EVCGc4IEEsuNCaTUvBVm
0FxVmrHe0DJrjlA4h7uMbR2rEpi9bJdf/m/DO9UQg7LWrx76XUHKuyaMvnwvX8zu
dF/Adz+sls+8iLbl7fZuiXXxfCEmGh6zEAaRiExOKwOeQjRL0/QXCpzUzsl2dKUq
gx09eFeFdE2mQORu1ZcOLhkxsS30f/4ipcx+9/VDVuXnGX5tV6g/DyOqIEHFHkad
ezVyXyiNhjs2nrB+Wgm1MZCQrT+IxvWObf0j/XUED5xqhsaUkDHW3e+IMH/qBWcf
8aAP42tbLV2eYLWRDB73ej3/GC6LthnvfX/Ls4ILihhmqHv93vDEGHS8+6l+COsy
uDWV8fnOD0l586Wqkg7maOso76j8Z4jR+95L8cYhnfwZ9UaibwTprElWZy7LdIEO
TNjyj5nYhoutsS4+k2GfDGyurNuXZB+byYXlioXCQj4FPO88DtmQAxvTUA9zBLt6
GI3kbpZcqnWd8rfz9QqfYRoVPSIG4gOqID1FwwGqFqurdEAYCVzCNMhcYzoKO8e+
21Y5jiW2ll+eHD/XwIQk2bFQjdAqDBBc8GpDts0bOfaKWKSM4K/bbgDHPp0N1oz/
PCEtTHz+qX/nyWdAz+canqhMF5L7qAcSfu0NzIIuvh+u9mypmT+18Os8FaOgSVUQ
NF/ZjoZ5imbhb+0FQEUlHIy7XI9biDZgzzVhQSAVXuzT3u5jf1NqC0PAnUOtlgb5
3zwRm/4I6phjlohP7ZurOkLTrqu7nnnPUkWjZhxYzPXLmWNFOLs4feQwGSZbdzL0
RsikrjwkftJfKaUMlc8X7L4taAOlyV7TbWpv/9ynng8ZkWthAf7MHwWLHv4esYJX
IV/C5N0HLjAaNOhKxQ9eG75yytzeM4q2uGawVcM5xKxjyBFY/vpR8a5DgBe77Rzy
sS3fITw6QiAAE09T02DkMFg+KszcVRMgC9mmJQDuUrHkyhtsrhReRjYPJh1/GkHV
xvMyWXIpAow1mKUO879sn8bntGcRrhvjw4KbJy9W3yB98ALCy+QRQSEveFfpe9rC
nlcyICsCSTv3+UZMbLgmwsesJaTn9x1qU3k9yEwWgFM8K3jQx6WTYnnyG5r9P4da
O4FZb5lJA70FfjVJxbY0g1F3/SNuK+Rp7Lq7OmT5IAVS//bmGrdN67zUXl36zKvB
g77eBjvupFSDoxdOOJ8+l5BBHEqpG1/Juwqs0oDhGiREpBmama9q7TozH0twKNDL
3KfdVFfqKaD5rY1utWWk1ZBYw2owOOUo7kO6cpQUe26C5VdzeoGGVvQFBKGikSqK
khSMCISrLD3B6UO5JaL0eaEW3it9uN08IVNS4gG/I8S/ClcJ4rv8Zqc98Sx88XYA
LdPQpJHcFNJ5RXzw5J7uulmgl0dgAcT1Jf2Cm8REnyHatp4UT/bI6klAIhTiJKtQ
KrJ8ml7PEYBkGfDj+TbW7DaILcOPbVwmONXczbDG7YTdHwmyodoc/G8NjfrsX8ga
Z6jxbXplbGjnGpE0FEhIwL4mz6lvomMbKTBSPc7+7viSarRgokngZt1mVhFGkiZk
ILfBN8iMkgiHx/zxXVlha6x4HRuSbkarzHeuckMViEfiTg0s/LcIfj9yuOl1INQJ
b4bi0jW9TlTiTBhXypClGz/irRfTavUApItO+3c2PO4R4W+wQaxy9RiyNp1Q4fkv
YmwkesKZgNahQqSP5Z9VCt1Jxzfqv5tNthNTcztv05bM+HcFvzgUZyjoIO5yIOZ5
M3RTPj5rxHeLw8xMMr2m9wHab11BZ77Pcao2ggWI/dTqQAL7XHOcOMD6hMz8P93b
0B6aarL7QTj9iz1CTciZU1gaD6QrorzyqRo50cs5NzsSYafIvx7eTNja1CSICw0i
J3+GgVkD2rPxKC/zMYu6CCk1owoultUZ5YKaVLWAyY88WnG8WOks15jpXALEglrF
yLu29ZJ84S0Yn/YSn37AmnPZS+XcCGHEPHc6LbP74L6oXP4gHd9788hsKSInXcOB
6jaqRTB6j+K2bgzUE6D7qaUDEGl5O0J62TIGiKRuf3eHB01cpZ1kr5y1hOhJHGeA
lWgA6eQcJ0IcJ03PP5+2ZhkHuixUHFMdGRV6IqUTMdDK3yaDdn35zmJxF9w4sNg8
QHlZDyLgF/1IxfacDFuvxnhBXTHjjxQ+k1Ck+uy5rfJojAxQeu8myzNPwbjvSuky
uQqoTgf92qdfIa0fljLDRsdFnvNYdtXI0j9fzkQA0dMIHThtWb7E/G8y+PYgE3SA
nUkITYt3Z6vwXxrw0932AP02sVjNsXEHkFKvD1VdoLMCMtbLOO/BbxxZ6BhTrDJx
6Nlu3aZyJ8TJYh+T066AHlQhuY1+Rpaz0kLuPLhuKLHv0ZHnT1F/WEYuXnx8tp+l
wP0A3TyYwhuVNyDjcOXPlBoc4O0ONHv6nW9JidZkuvfjeWN1MmLAJ6drrLt1H38F
TVmXs35g1qexKm8gYVcd27q5EvJ8Ns9aODUFsre+x30BtkxwbA1vWFKVX5PURno0
S46ZfdRbzSFxiiHZENwkaOPLt6GL8qxnY5G2Tj2a496xUJqUaBvk4a3etFJigCtA
dPLPc7DHy9fK9YhlmqMlLpZ40n5ZGnw/tJ96Hn0Kqboe5LsXRhjfUuPOuQ24gBQR
rjHc/NCOiAOCT8yActw4PdNI3JJCO0iiHXUqquypwPw9VBAsPF2tLVZ69TLsae0g
/0q6Tx52jc6LzQm46EvFhuZjKActWAPuFXjCAICR4FCnrTP1txwvH/73vgcyaQxW
T9Qp+iScxnga6FufHUrHzLCP/tgtZmW8ZCuwn3eHDKm8/hyEwP35QEah9LS7ADHo
KuL1RreiotaE6jFF5nshEajZBXwZcvESfwM1qh/LPHctAjm/oXneMEZRq/Lz3csp
8t+yA4/h4HaEQ/tEEz/yPFV1vULbEJQfw83K+FaL5QZ9AYH3V5igVhQsXhIFpsXS
DMpbx3L26yBK0eK2iXgNBbm74aqMwntgtrYp+fo0FRAc9ymRs5sBBheR6MIp1Pam
abJaveuICHImUnQy4ALMKCOpNw90embYBjbIf2NgDBBN/G5OzHEhCb3fyVfwFbKI
DCwGjHQLdIUPA+znb+JEAQze1/XcPkKb9pcq66GW0wNN4K99Dj1LKs/dA/noOV9y
Z8NIj0IqxPASoEgqV7kzY39ZxtNY9768vMXnN1/mRd0QtJ8G0oKLxV+D+5afjhD4
UuiLL5v9gqiN61ijgPZxuEanACFoAMHYjHUm3V4Npg15r9wxjNAS7XpODQMFpEwd
kxsgAkIcz4pBOWVFGKJXuPalh2x1i11rqYZ8F+n/puJSTBUF38xmD18qve2I4vza
1WM/YdoXnWlQRacwJ/KIUbI4pQibGAZz4MqwPp+ZZd4JHKYGg3Qpj4LhLAyWvCnV
cTcSrGbY830T9hbwJXiGw7u9Q8LO8w08ha/dveOpel9/cLR8LhOaT3SferTX46QR
jMfGTzm1HFwVL+4mm4wTmT8UM1DNEajpEM+vMoCQ/jXl0ZiMONeKMoaoHss6sZ76
qZjbGke3epWHjIYrL/3kXlTb+rYJYb2PqhGI/DIOxUBjJ3xSiwBnGLXVAYYjvE8u
P94HCaFiymL2O0nQ1VWOeI2hcuxIwM0zFU3pQYzmWKYILeJOMVHaezrN95YXmwzI
BOThmrLhislTtSufGxRlAiCY2By4WESo5edySzvVIv84Mfl0F+DJXYEhjbe9DlVD
MtzRGkWzwSBX0JtuQbNdufjbvo5HrjdDN/3YLcMFntUQ39MvlQ5E9cpLAkuaBtnz
iB/zy2X7vVzcHDba9EGZpR8KnrE8eOr0J1fM44paTHSZdqd+bddOXn/c2WVVg5Ws
/VFqyBvf5MYEOOXMhFlakm5c2ehCrNbM/R+tPycLeKqm4KKrQxPdCCFo1K4OBPJf
vJ7sta+Z6CG9yqm8nw4uCx8lp3Mg0wGxZ2s8xQKmDLbwMk8/axjHFkD40HeSAAPk
aK9g4hIHZW5US6RiMzEpqCDQBHQGkPHhYPNBCji5YXgMn614n3oSTkEYdDq6vK3N
0seuAGCBAfwC0EQaMuEOOWwgVUTpl4tw07bzxnukyxE0i6iA67FxzCweQYWL2CBO
/+Cwomc+zW8Y/YdsCJ4t4xaQZohBt8vQhVZxx+RwzjLO6her3dnf4iBLpUuzlRKo
cmzK8cZ4xUYdZBMgkqcr+doD1Xt1tPDcOfkGcdynD3Y6P90/ICrDypt6xgR2XCvF
8QC2ddO7IB0g/jpy9EOA5rgaD/bmIODfWWiWkjqPfJ5DJ57Fttr8tUaLgPJ/79Tk
IzJJPmaREOhvCCrHIeKdOy040F9tb11Per1aJheae+ebZJCGq4/iZf38Aj4ggO/H
zyidoNJ5ERwq1FbpVOhAONf2/PU9o/C5wT1v+QtI1QnWpXNny6wQ9pQzkI5BTsn0
ls1jmdzIxQHoYdAQGQ+sowhh492eJPKU3CdscuO33R4X2DMN0QkWqJlM0rXQOvvh
8f2pNPbW69sSl6UCraSzPjIjkPSA65FSoR8FsrAYUyj1xprdZiIfjmfO5qaZQw+p
quUGN5osrjS8shexq4hdsr8tiK1taoa54KqhrBov7ztvwb8brk/cCQuZwqkm0z4H
YfPAs3N+4o8DZQTuCu/FPpCAayC793dg36zxAI1J9Wbv7V3kmGl7fK4Va6zWsgRS
m8+5duMbEq1PpX7rNy9XqCNBGcNoo14L2cZRYKDt9yiA87Iw3pxNrGD12G5GrnBY
J5DSOKoTecZZhALzL9bLOJN9M321uAYZM7LycYfMXh/PNOL804y3VuzHdjjP1aBE
NmAZBIrLSu1HITioBoawOvWTKeH6RhXtKaybA+iMsRpptg9z4laaOusyZMnOvlTg
6vJq6rPIV9Laj7lH/7kJ9RwV3tkTWLaErg1Uif3OzpEDk7W540OvlIkH26xYuKAa
Wo6rJv3DEG+9iBFGfNSf97MArmR2KvPenZG5WQjKMibpjSBpCMXgZlubqZpzQnsQ
BXyOwwfRsLxf82MT9MzivKffElsy/DgmRe980dnuj1J8y92NyEVJ1fH5RTc29oAy
EuhlV4RlphS/MdC81JKuku0LAUv2Eok2jHOU1ohOynV3bErboIZOY4oYrM+qjbou
MJWlLVY9//OYtmcg8hp6gWR5b7AkE7kH6TBzhKmej6VHEx//1G24mIYPhOpmboiG
1PGNTYIB43w1jG8o7Xfxi4DktKkGFgNZ5HBGhfx6leLcseGjtCRUZZHvjPiRAG9I
uYVTKAt4zhNGI9vJuDuYNkkcTYt5oXlDtC87lkrNokFb1ApLTyPBb1YySPzcRXK7
JMlA9ktji0/LfYZdXOiZkQmmFvyTUcFxTSNTvbMBlYA+1Zm8SP8oK0yVKht+KOhi
E3tHgjjPoMhR6RwEwjo3/0hVboUK9NNxrIkpGp/JpNFgXKpeLJZMIbB2p75ZkKc4
WIrfcc0kwLGU2NO0Xt7dVOT16aVn31p1csg8gm6Qa5y6kNnajAn2rLJAr3VceCQm
6lZdtjo7KxlG5DEDigOxsUI5NheMPPTefq7DKCGpH6a0TFj/QNt3LOxFbdk2VNuo
MqSu+RFTsHz5rJDYd8dn1ztwmHhbnSNkOrqNbXu3vxQw+zUG9rx9CGNLZvjEbgOA
65k/ta4isHD63fwMlN0nxv5KAcTq9N/O4C/0I9SlwOzoclsIUIPPmZwkH53uKbS3
70mF84KAurlrtEDyJzBBVqxTTAdz/Fb/fK0/O3EjiLkWandicg68Ur91FIyp/QCl
n+HjR7ZVIWiN7bNdjXtYGakzpL1JYxvIJHtE8XNDr1wDNQcSUI0Ig8DTxZ5XaAOk
+j/G6IKCOP2gbO4qCIdBCf1dtZIsslnxj5ECzTu1usymnwJuEiQVW5LkTCLY64Dh
5lSFAR/fnrIyxq+UTCQ+YD/LNhxs5iio71jrMH5zUD9LxCt8sP/MRXFrbfwYZ9/M
CoToN71lhnd+DzJpn0i/kPqBFL57uzaYTEV0ro9mV7nfAG187MoyxGuZurm9eqeH
T3+jt+Ktb7I7U4jtFv2CrTL5TuKzhviw/oAxCYsj3TSDaSTg28nvZg/AdWEDEWFF
oBi1woGTLzW3QvBqJKCl3Vlf5QkkuPMFSpCwFvCtvbLT0acI4n7ZZ5s8AXKXEi6J
CXk0NmTCYcomtUjsKu1ZD3+FgvqUQ22icB4eyH7Lnv6wUvRYDHnd56AMmZuU9d5W
L4X22i0L9pMAd19l/HxOF/wkVn4oUzxD7QGAdNC/x7zvlOcYE2aqyhalUIItiApQ
GfhFBIJPtAZBKNiwc0NYCGmNbNfQVjSe3vdfFDGnF+Rk/IzE8XLHYVFOu4JliEt4
xINY39LsEpA9SGAK50VXPZh8N6yXhgJaWI5gf2NrbM2wFh2NtbFwHEkTRNN95hYh
9bc3DsyZ0GXvfjJ6PP/UwIMzDiy+2TcehQle1dbAhBiv6FzP1sr/KAvwvnzlr+s1
Cxl8rjlMm/8cln8ijSvscKmm7L1mQJi0TJIiUGomHcLIzVF1VdCLYcWJO1W60MsL
hi9LV0aKAiofwOIcG9ScIRjbmu8suroFsRZK8R5f3ffNhQ5fbADCOHzzzQt+Qkl4
FxTyC+PJHIat2tmJ/+deJUSdDHD7NIJEm8xjgIzecwmKqVMX/wMh1/TkGzoyeIpG
Q0PnHf8I8l1Xz6i+aqZe8R5+5nFXaz/J4yLqUf/vNc78Lsq5nOJW7gVRjEcxQK0r
DaNni3xJF7F0HcBWQtkOCj3rT+HNdt1c5RI3gEFmFfva2s9lDY84DKcrVsfq1WRH
94i2rGpOTwuYJ8vifyRR0Sb4yZ62lhpWJrlNKEOwIGmDV2F3YxXR5hjVL/ecBjgL
3W0c2AMa8moie3eQoxpDUpA59ezMzaGJu7dZlXa6+eIB2lljEGWyxNiQQq5yQr6m
RBRx1ezmEgzqyBK5o8jkuPX57OgRLQH8Kbej5Bj1OWvvxH6nyRttQp8XjwtfpcUr
GHLdq3PtShCF6oAvgONvk4i8D22p0/LcGtWkl7EWPbzll1kWH4ZHnJBwoyJELG0D
I/5ZOyg/IbMrZX5jorFWo6Ikx6jS9my5InENVER9gR7rrjpR/bezSIFO5yFeZTHR
XfDS8GviL5FXf/b0I5G07qvvpkU15+DkWtCUDtcbBZj38XEnoMGLBy4eAhTB4dwP
vMJR7k/rvqYV0IA0odFcRc8pfCRfNpp4Qh+VjpGsZRNJIxxjE+G0hspGpuiyTWlT
xyLW7d8NL1mf3ZhvlL/A5+ktKj4Eam2n+/OPfjmsUkpj+DAbvpfGQyk9PmE0IMd4
JMC4ERVm3wfXAXKRV2HynNThY3gvZWCWvEVIIh56mu8J4xJ7OhOAifI5/V7fxDc3
1lQrca76EW2MQ28OiFGWuJ37dFmvjbrYFVNQaV7vbjDBUuxGxm2hhYAx7xBvIaKA
EFNx3t/julMt8rFqVA28WwoAjtgIw9uSyk2lIvdDvkGrdqrvpM1fCs9xTJmFTAP9
yD6U4wpAl8BtmN6XfDqLLd07sFWc4xiiyfbnHkdOUUgyD/im2cSGYJK6Zh7B66u1
Y4dSEQX2saluP2+Ysqm7okb83L15ibBNoZ5Rq4lcpCb9cnyR3wmJAGv8sfTNigYo
eSw0bgeyLR7DMOW84eGSW8h42fknRXPRBOkSWiuAw6KoAld5Fuoamz3A85px99Zg
6jAU/Rz+ccr/G3ilNkBTmjA+u0d6xFMcdtm/8eGIv2MAB6GO5gD/5dFFxCKGaIwP
qyQ0NCDYwBJRNswmLkCAIjW66a+AMc4S1ExQOfesucs2NaUBHwWbEG/yBRNGT4K2
wpJkNETQWx0MRc+H8FypcbmmwisAyMi0BvM3GOCXuzsDFR+BusRpBS+zm7qDARi8
ra40s34jwEdcC73IPvScZpYWp8gmDVubov7vOhSh7OyqRIB4TV9qdPZL16CcTjw2
JjlgvDNirSHgwUBSAXTviaB3s+jLCYkiGef/s7RFKazMLz8plGzCY/tqFI5/Fr6l
ot84pBSvi3ORcsCIob/oiK3WVRxEv1hAkFZQxssl8VifiqiThChBypnQLy8wH0Y5
gLUrXqPSpCQAMLra8HzkBX9OsZbrEfnpsL+CjTyeOYiWd3NB/6j9BlRCHBZK3/Ux
DIQNRH5qBFT/7U8bCWN/UPSmusVexyIpzzn2r9ts9h0W09FrihqG4s+f6PSak/IL
Ve20vxuzMdwdpVqK1m+N2e0N2VSGFQ0HuRl6VAqvPiy96rdOkxZkZOToMr6RMEu2
0ouwZ8r6lIE5oKegf6I3xvlbEqQqp8dqPaVOnL94aLDMxNW42WBiPSzNrM+CjNxO
/95s8n+Hhdmo7PHXOlXIgYeB1h7Ho3YdB9t13bwmHdHC0TzARx4Rc6z3j6My9/Ju
FWIwQHD2GlsDlwr7yqEQYA8ePdAsfQ5R7zU5KUMsrsFkveVgN/Wypi+0fSRlCqud
qFh5GFekIQ/lOlBpI8lhJULHHJrfSLEZo7OzMv9jUP6dMk24cVM9IjKIH91tHLNT
tqjMNsHH3A103EcTqkJjPg59EdDUA8Ge3auAhXcxw+omFdeL8VdgXvmNgAFp6APV
AqeGWXO1mMjyKru4jqOVKJn1nkh8GpzIkVeNf6sirKgSX19Mi0rWoBH88I2WnJAt
8SGUuC9u4ha2sHCfQSpI7H06zVAS6jIIxzLqEvGIiHsLHCbp2u/7HGF3nooveLLT
yF3NHBJPnE7U5vdsx47FVUguNdGQHlAdqPitx8AfGbCQOjpq93ULh1YxTcmdsdA1
kEXf3KAMqtUSp0Vz7NviumUNRgppHkm/Adh1r05/RmhB50zXi5qgj4I9RG26ICKt
GtLwbsUNa1OtuXvLqFHYuo5FJepr/noobJ5AUTby7/9quKMqtyGy7XIXuaYKCQxz
3O9/P/q4/bw87PccHSSQtvoclQ3ZfHIb7Lbc+uW9ofdCQViG+MHs+dhfqzd+Jzjt
RQBCU31n2I0fNE4vAFQKdcA+Wo0jcOdufHtlVkHaZ9s+8+ZBGgHOmk1sYfYSWkPg
LdhzoWYok2zcFirHhmaAoDjvM4ogrxT1TqXXxS8YUnPW4aETyIrQOwX0dpPptNSD
grkUcnpJywjyXWpNdkv8C2d44PL6wUibF3PxjdYZZm5bWHJMr79pzcbhn6xfMylP
OOdC0wCn7mWBNHQXCEDaWdXAeSo268z4LhgBrTIWFYEa4lAsDm6Z6Mm8vN7y4VCY
HVoKl362y32SD2zlmg+YJz6DnxTH3jl8gPU9WRsfH8GEkq6R5q5LCLMrukSJbq86
Lz4ZEJxcFMfsfN0yv1iyHJ8U7axSvxEzQ9rn+iLtJIKt1H+oyieVsFcJ+3loze/z
/NHTQ3ff6xmx1P2edldrKjMZTWVe+tvPDsjBQsNEopYdtI2QZTlZs9MXKltRj8Jm
3QowF+n6kRYyNSLZg9ZJgSkhzVoO9w7+L84/CaH6Lfg738uDHqXXYw7Nf5+4eWTf
REPkBUdYsnKQr2cdL3IKMjIVok0zBJk7cGvfICiQ1ziWaV9mGsD5KkXoaBv5AhRy
msSp/JMg13RlJZWGb1M+rjWPWDDqGgODwTBmczgNjUfFemGWP6NTtKfjz11r0mHU
WXAbyhzUHk+D3FOTckhsXBRkhpRj9XsnUs2DB9SvtbT8MRTLGamT8/DIbjVtumwS
G7mt6sRSQQrsFTKgvkVeNTym6tv7WdVHH1dYLIAkfZNxu9RueI98ZUkqb6adPM5y
aX9uvHuoTKa+I4F9CK8dnWnyQ1uonTCddnprjfed1TCnm92LttY6H0yOqIR0YTaH
SV9fHzAiKv3ZDV2qeFGJmxPsQGPP9qk2fh0rzm0I6pzs2J0jE1iWnOr7VrCFsg6h
5Kl/qGNcMD/kfenMJrQ4zS6hutHP4G2/bM8nI7TRMFmwcC393BZBSsdzakV96alO
0SgKJ7yhwxMrehyjfhB4An4aCx4IOlHkpaeNm/xEdol0GpNSZfhsAgHhUi0cmANq
xkjqnffUcEVlIkmrkRJ2sSOa0BYOdM8IL7ynrjvVugBtRnbWpDMGG8NSjRALxruh
h9W2FE8OAEtjDCj29NB9ZxWzBQSuSL5NVRE5c+hmJyT6aEgKMS0YgDWy8NFzm6af
nfqbF8apkwCisJzFSzxFJjElsHacDCX+qBPT++he5yCFEaE/ms7NY9kXbT6vm4CC
Gm4fe5f7H9a58o+YMfPMVJTIkHmTeaaLjPWHtXGpycZAV8cuTxEcjFa9UfJx+mXB
dFi4/qKQmUzbg4lJEQmj6QGrfVA0w/yqiSfETnuULdgsih8T/VmcrPmQ+40RvH5r
JIAhTS9RhT9SJWIJ9EZW3s0kXMbklVqdkqfrhAL8xoAGV8tqMxz5mLKWt9Lt9syd
u8e+ITlmKFyw8yQ1XBwpoK7SHNU0Xd27PKikI7Xwend9bJNh2hHl0K9uK60pXZa2
zL2uZLKDLJSt3WDkEd49GGjAUdy6lDtVMfZm8xijKb99QaLuvC3b7Wn5quTkqvP1
LHHTjSbadupY+AokkkF2XLXJG3KZk2ge2lQUV4S4DTlvq9Kz8sx8cmr8PCY+2kSc
c/TAacSVJZzw3ZmI9uXh8n3qpXwbTYG+HQFsDWVibBluM+bfB7h5exOL18J4B4/0
gaBqI6+e/6uJx4mP41NQ6cdMuwq0s0Iu1qUww0iR8i/yUMk0P70C/CQz0ZGzZ9Wx
rDSIDV42pvtu9TK0XMqhYp1ssUTEO1acnRkUakwcyFtzkaO2Xauo0h0YBaGpm3uJ
KjcCQiiWIXzoAFtTN7ekbxzzIStUpN7xhA425Lyv5fe77azXUwDu9pRIrnosMBgj
i+oiJtINszET4gTrxWHGIQg2RFBOjv5XqbB18PgFYB9E+DqT5rHsNoGXC+4qFNPS
uUsl7vncutDXu/aeAkyOwmZFd1fgUFfMckP3pr/Z+ffw7JwvWto8WHVlJj1duXHE
ZWP7Zm1rozXRTqoreGzPWNYU/Xpe3vR8RynW1D/6RFPOlllf4C+ZK0spYYY3Vua7
DO6zCfNXmW7Q4aaITDC3ImftNWH0dUzjiM8P/KpZ6BULJ4Cf2D55RCjI0ncTUsY/
Nx2e5QLsAV60WihLihk7OxAylpsSiJ9wZVfe+5QK5ttFY3yeRKKG+/A6ohIkJuk1
Ia4xm8CHrDSImuzj4ogEpecpPdXDl4EI50rHxKKICFB4ggfgw08ijKkwRsD4sUXE
R4JFeGyK5ap6drPlGdWDYutVnBC0ado94lUqkr+qHPFIVRyiy6R0AaSlPuqhguyp
nS5owTomWANu9JuqA2UWLV1Zx7ye3OJRIQkFusvvBkepqgA+nlfvXsLI8phcDVeH
ysCM7hHENRiHBhNWb736nmMYpGAcTNZbuRtvps2l/bkRlJ2kJndlN9Rb9wFlTFUD
k1bgEMpHILoLbU3/R+1FdF/geELXNIFRX+XJpwk/lWJzA+KYaY/vTR6+RTvC0YCE
f1pH2hh2dbk6HH2DXlX9vPnn+PGjeSwEK3W6EI0eYPBsYmYBzObwl305Z19AoVf6
PwhuzSi020kwWfjrzUnhLUgU8Y3KGPRlYA6fQxP0MzGNW/04jozg38xUFOcYMlj7
OHUZ8U0H1TygYONHGpKxj5xkN2pduQa+i5FHfkdzo2h/qDutJ4FYJ58RPW36Nc0f
K49i7R4izowksvDn68U3vuIMkPUm6g2BMAYb5owCuUaWUm1pxN8OTHqXXr87PLPt
KjG48MgZ2QgoGB4RUh5rqRG+n+Ay/PKFSl42U34t1fJG3GW7SRrCH5e4LghZKg0K
hoF/UiNIOL2wlE+E1S/I82uAVBnhoapPen86Tu6S+53kMnhXaezYcXMGs/aGRPhh
17T8EIM+Ntq3fsQ2oKUygRH7mvlLewkUmYVIkuUcdm54uU0qQpCDUrOhuct8Fqh9
/E0qM4CDpNUj4STRZbV8Or9KieluuJ/tSU0VoqMo7U4VaqzSM8sSBsYie8KhbYnR
C0yNB1G+ECg3ao6321s5L24pSfmCa5V5h7q8ZLZzvikAbsiciCRb8r6KGzw3W4rl
eiNzHwKrl04Xpz/zyBHDnFWNdzfRXm7VwB2cOW3RyegFrfXnB67TbQ8veJc1fkl3
2/iJB1Lo64OwfZO4yj7UJXeTpfGIxwZUBWvC3mgpxnnY1/mSmFSIl2j5WDgX/qYJ
dCDr+q0O9KoW5yRIM1Pm95O/BSj6mSs1mBLSQsaWt8gaQjwHMXGUJKgrKWz0uIGj
uXh9EOFAoSrlA5iBmpj9OBF2sgpBEBYbzsYT4+p08b4ribZbeM75Dmspsy174lS1
5LeVGHBG1eHKNaRL938oQrXFtM0s8WGVFT2pzRsMRfcew1bV/v8QC2lUYt9fmxdY
xFuETTIBQ73WqtLZPcnZFo8sVHowhX/sqkpLzTmXk3XK7pg+xBqTwjlDoLXH0d9Q
l4S7FVpCnZBx1Qs3GZYm7h9S+CbtxMzrd9VHTBpJL9iF5yNYqjQUh9+W2gG9XzDQ
+mG98oB/oRYq0GmbM75Xtf7F35zCIIxV8M/CFvqXQUWj1j012n/DGDO1d9HA8aTA
w2tS7ZqtYK995Ckh/nG3or/PEJLnhI69UdYL0nqm5RU3pcpe2BfqQ+MIiil6HR7g
aOQ2UdGF6WGtmPTGQDd1sZkHTay/pk2Glif0eaVedE2jMxghl7tka0PUO86LQzpM
A8A4bOF2+dsmOGLQFQKVnRjcgwDdIDtbE61JAYGwW3DgsisjOX8a2tJU5cpPEP4T
tDSMxOUXIacBI9G6CzZT3P6P6RR/6T7IFCdSeZNcOSljCZ+BZPclaZ82nVnBdD7v
JDkFdyq2vI/dvtazK6AKnACSser+4HHZBN3SbQ/vQ6KXHDsH7uLPbKnBBaspjNlT
HHwCsctHCGfsUiaLmM1rlY9yZDbOm1Ku7os+pb7hvkxMJJVqocKU8b7Vvot/POF7
Yqp0lN2n6aOeqS25Du34vJgUkHkzCB5l6fqzj5fFVtmdONN/2ZmF87WUDPPGlvl2
/fP5pr6Ls9NQec99xcYpaZrf59bYUVqNOWiY5IEVt9NJExq1W3yfuOh3UQedSLHc
jFlld9jLq67Jy5/BpbfibsoLehWacPNFymu5lEPNpoT8PbdBzX4fMFZVmzJ/XSrI
cY7xQAIoGO1aZDtItARCxFl2w1kXlJ7CXE9jbn7qawNL66VBO2UgV9AEDbIr/0pE
GV2OYYgaOtHUL0G2IpZw+ygE/Lqe8YuWEH/C0jpMXpOfq9M9rC9nat/UgcSuEIKq
0iV4KFRALJ6oJSEQW/vow0s5u1vDH4njgqI4GHijMyIa1Qe87sdZ+Y+Y/2TF6ZtL
EZdXS8NOvmmbsz2DQFoiCiPrunCe/atX21vmEnTQDP5Y9LTaF0y+8edbOFDBdRsI
lDSxywGliZ352FnduF3+MX88jK/nTyngJRz7mt/APWq50hY4WLHbl8woYlev26Au
mKJYqPve4+83P8qymAhac8TYdXIjPsJRnA3G1JJ0aAzqutlaoADfkmGCg4t6p3i1
dDzSMXhU+VzBLyOnVzv14zP4k9zvyr82YHUP91ul1J+Zcz6OYoDg5tvOPhTavedM
9ARiTB1W4M9PWoRcgWgCY3a4Mha2LBUWgEUF+4JLqgauORHAPQpCKFg9UEoN5Y2w
2tp9FQaL5YYEV7D8dRQn0eW0qlej1b9RDbG1dLzqq5MXMu0Nq0yXNCaU6ykwAnMH
uTVZ0N7CvygoZHKqd9grDPKxoJ5uxTkzm4Yoa+kXbP2t2APlWOsy4NW9lPOFmgoS
5iLb4M7n9CUNEocQkk/rM9ipffMqksS1+2DD1eD5rsN0W+tF72qn+tCA3kGzrg7d
qb9+teyudgZYc9UpgldAIFH8NG11EGYNcsI3WVcy1eY8MCq66QXu44iOBBYVtbZ/
EteXeRA6JeyxS0V5HWP619MOppCFXKOdq/fUssrLarye8VIUWUOqJd3oY3kjf1A6
jPAJu4CUhgkCFpiLyo1ynBwjsK+BG/EMEQohkymptkSyZaKbr2kXUuHTOnZQliQU
1ef5MoBFSkO/WTatBkHoRV5YJ22xE/G1lLpK+xOy6gmPvzPZPPFkjL8LylvBtRTF
HoGwnXybBnMSuSXDFvzKXn/INFkrDM9ipU/q5jmcdGPFGGru4v1R5zqTa5yaxbi4
mkmqgwYgwwxGuF8YI4y4YJM1666mHd7IfPXd0/Pa8anBfaYfbsmC6xfOABQI5zMW
SGB4wlvjoVaeSQW68R4n8/qNWjjyTJEY3+eFH9LAeo4vhWEMbVFaRUvK7FLaI1R2
ZsgCvxyjkXZrZXQM3aplBvcQsAjHqnBxkotDSTx9M6sNZAdnX8znEd2+NusnFJPE
ZfVHGMPdgCOc9eQDBkmcp2R+oY8OvHhlMfgulunpbbP4v+gMeqzXEqddkg2wd2CS
gRdyEm0CqSYAAR3jfdvSg1V20WuXA+oFDRBUVpU4PtkdZdjvGn7AO8YuBGPOuToX
u9okEbW+PuwXqPAZ8NF31sAw235d6ne7qEWtLxdX4Y1MDMDdghxrDSiMUzPXLgbj
Epxm2LRQPBtE5yn14qCrK6l/p95vPOZTknLStWSdKjfS2p0H4TcX2Is0pb1K3HMQ
J5PJFnETqVV1AP2tv1eWl4Jq+BjFOc7lpFWDYdtfhFutm1Ihf/X67cZdEcrhz4SA
+a6dAaUT+Agv4nmNS+AekTCSoMPfhxCGZ6kEa2/tST6hoWiHhXZkiIa7uotFCRLI
5MCZxYEe31s2pUBUSNC9fcxdSFBxu0pEGO0zbB39Cg3W4stqJbP9b2JPlY1upg68
b2aKxnOIGVBYW+9XUlxoEDIJVN1YAO0wvukZ+3QgjG/2JK3IgQ4XWUZG1aMsLXVC
D7KhwQhv8B3A2hlAC5bxs93l+j4zIEIUB02OpSxc2CvSpU9wyUvA/nvaPv+jWOYY
cEaCumMF7E0hNTjMARaNslAhV/+zxqEClw7Ot964NqUkHz1b1AthYd0Hqzcbb681
cDDV2Pqlgmfv3wfOByuYWG6jK2FHncdbLfVrWfkIA5eBD09jXFEXVKlg9oU4Bj+i
mAhvmHaS9e/PZToeEc5wiO9PZKtBU4C5b6Yx5zYPTggXEtM8bLeub7NkuRUitmzm
9OH9m4+dh0TL9njj1jBDzgN3yNl8tHn0CtRSJSPMvUITPj0iqX9c+paig7LDENOJ
69958eU+ZoZtIUD8pGHDZsLnWnrPi5EV5GbQLHDZtjmg7XnFDkgXjY2PxuoAk8P7
85DY3dXDOshdeqsXWovzsini0iutRD51DbBVYGJwe81OIitee9LtR9GoGLyWgK0F
30l1R7s+lJLKdSoB+dquYhQjStTTAp/vBxMFAchGP0ULxkgITHlQurNh7108etML
2mFKP+nr4rVSIjTUW1rAc0KBDhf4yVDTjddmahgu1+HdWPgCmPYU+cX/x9r1Qd+B
N0zAvOcuGUpmlU8+IO+Qvf3Bw/A8d6Zbd6s9BPfY7zLxXHwQcV4Sdz3UihFu3ofO
/vtQU7OguvnN/EQkwPcexuBHYZVZV0ZK1rXGPeW6a/DH9hzTmdUzq5Ao8r8a29Pr
FQwyMStgFXJtT/pLECHr90NjMukq8FlDcrS+F6/bgCNYD/sw4/AUnTTCs99ZtH4G
E/vNklWnBBwpNVWkaQd7aUY0l5Eawdgz4r7FPtWGVSh9bVGwv50LdWD2YM1NZeNy
GF9G332j0tWH+SvMwLokzI2/BIj4jV3mKxVuWJ5y70akJnCa6tc1WOMGfuh3Qej5
U6I5Iu6fR9zdzZLvNAJ0sIbVJutUp4zc47fEvhqtW7idsYgv++vUq8owVvCnO5vg
xtvfsoUzUfctH7LVJZJHBwQWS9v99EDc9mqLx3UJYYOOea0dMz1rQIBwLohL25u0
ZsMd+nK4zGoFWq+265Tg6kj3HPBDOrFZUZrg8/hCOrORBR694O6BN8dKcHJf0nTI
q/hrJ/RzXSJ8KtMwGHu6zn5tvpit+qwTk1QBBA1RYx15OoZ2syjz45lWABGfmRhw
dOFNl+PEY58Y7lkR3mkZ3M17RhNnn+uvRBVfwWLtVgFccbUB/AyRGOknqSdLlXTj
aWeKh2sSelljbdKXdmi4Mt6EztUyv2vWL4QPkFtyj4zr7hhKtsb0hA1WajkuChL2
KK3ar26/im0bAaMNYEOXk8sLI7kMWD50Q4K9slqBu8ChDIgJ0kHS39zWzPd8oVGP
wEUWK8jo1dbW/WKO4pg6aC1pYAGAqzjgyPZx5dVGcM+sn+TwqH6t3YP2YBf6Z1lO
9oA1/tjtFigLoVuGF99VOfI5leMW+v8DpPIIipg3qE4UsblKxIz9d2Fa6ibsAzzc
K4dVp8hdrYkzLczON9/N6NgHVK5N73EitOZGQ25ZAAii23FCfEPbRCL0z8gQ46Y8
kjQAbo412jh+pRgy84LUQ6MFQVzDijXeT9xIRghFSiVHYicHbJebldfEt9sFmmyk
gDZRMa5R+4/YwoIjkA6pMjuUECoL2v9s5FbsBNSxbi/FzTR4I/ptcRAPNgciWG9A
6Kx1DS0DD1/JsIgkr0QPFMls1WaiqH1AaFyc6ZI3cmAt6NE2XaHzBwGjsQ9SU9sC
HwvseuzJjBtKNwLhFjv2di3pPl6OcLwNX7Pmzr65/3NRMh8vFELDMENzWsb3bH9I
YUO6G4sbiaCTXoWhgoHhDdbhSvcc/R/75H+QISQ4iupASrhoTHgnBUZkIS28mrYY
sLB0jBh3MuguLo69Mtqc3ouIyYJZEhESiCVgYlSocLW7zcoJLP3r19W6wC52mzJJ
OQCWaesATwNQR5ZxW/12sE6VY3hvi+LEb0qvULPpiAPal79UfdwZJqPeypU39pdY
XJQNZY5T6QjsNGwAGgtfbSp23MeAqhozi2rdqjlXYhv8fWQ0WIaPQFvFRP4hkuln
uQQNHuaMDAINW4wJ9BD6OqWNEf4SFW/Is7SpqoSTU5FD0JFOqi3cO6vSksxj1XIN
r34G3h2ZrEkDBGvlvfSxANZF7PneS1DAdz8FPqJ2nR4cITymw4I+wEPpc6tb6ya+
8siTKYN3kI5hCTl76BkFBx9kvOdwojWF0h/x404VG7lXWXRNjLmCQS84Bz2hEZYv
jqTww3b1utNrDpAWlE8k5BhFVZc8Ef+r7ZBwE1ZcPFZHa6Bu2eOmECcjPhBZdhuy
EUvAg1ot5gCyjA+D6ufay2dqdsMgQGBR9Xpa9q3sEdfDWvRNt56UZ257m6sWauTG
tMjm7twv0ogDe2HKsayIac6wu0AlgFcBWN+OVyRIbwjoEVQQbY+FiF4UX/tjBX8W
QpzqSFhh2/6JntSGCME6TkdhvlHikGjuC+BHDwMWvZnL3+QiGUKpLDzNClNajBK7
WFsmzXldYzwCzIVl9qeBhr4qYFN+3eSteoMOkh/KHHXyGnARmI2e94PM6jnzaipS
bkdtyldEfypzmaCg/aOzf54wragXuI4up81X1lfdYWGFKcSqLlFb2vWqPbBZi8v7
3MW2ZE7ATCfqFsTImJBymoA/mciCa9NpuMo4CWi05r7OGIUtBEAnFjihJ9i4UnxX
fFW3N4L/8UccudGVCJHo9uMXJ0SM55dmc/J2Scwsq5hDNMHNHQ9ofg0iFxyg9JUU
FfSzLI6uR25m1QTdmtoQtOBv9SzLikezIurqBiCNBG+3tjMB9XWXZtNLtO/0hkgH
zL+uTMKcH4jE47Be0OTPtVHyCXby3l2onnsh9nYCPvDm2qvP+b8vrZoF8NB2exck
UiaZAkKw58ao9sqtiZ3oF/3C/9Z3EjdYbIV6/jX6vj/tNvZ/nBtJqrcryysdLWTd
tWXmkROzaopD2XBOqakoSAUOOcZuAeN1WK9aspTI4B8Ufc86eP/0M+675NRUkOVX
W9pK6dMgx8VHxVbxc+hSJtrntNrTudO9TnRtrP1TUFM0HP1949AG6kQR5NhmJmUJ
q+GQYS6YEJF9whu06wibYnS3n6mpGeDUMWzilljtce7SkQxzv/uyb6L8aS8TQoXW
ERwHobCC0vKvgMmIRnez/ybjgNDiyZyyXTcxPYBnFcZgzsQtT5q18RENHPOVy4Yp
Y2B/PXsz7Z/QKS88lYq019e1oChgZ0Ojv8DXOmcv/Np1vGMbCBJ0VjHH6/1TkDF8
0cl1aFMFtx+FNGOnGdKxKaYAWaY4ziOTP3nJ1wjuUlmeerQBJ5knAr/nsbGui3LY
4l19nwFBS+hoSsZ0J+I9FIHuZqUeROWRK1dwvPhzPeHbEk6pnOqqyy1MzDJx/DY7
i/u4kp9BtdSQLRbv6yetbKb+OSF1x7XcMndEdO11jMrT+Nqq6Y5MqCyTd9mES8Va
mBNeJP7e3Bgujp5I87lVIh3QEsvKUkBVJhQa17oyCa9hkY8x16X5OTT4QlUXSzKA
awIMQRvHTYxbzrpStw/KjYWJnI8ZQvWSscBTaDQe6a3XKmBP/WEtQ++hMf1yDayq
OPGPS8OXXEISwSQNIfIbhHo0eAOn/CZvMWabLwAiOV7y0brjijvuuIPCrMIlTz9h
WX1mypvrl9qOgYyt0CXrGJNginT2efOjvvfkg/OcKEiRKVYrd2VuWXffEd2dDToR
E8OXdsQaUaIWW1Rma1k5Uu1ehc434ZkWvcLUrFM5XiJ4XG5NV6y1afnMVNMXDJgH
QHmSKd00nKkEH9djyk/71WB7UPK3YlX5lmyHrDKQJ4FLc3F602ZJ9ay8mGEFVBBm
qNTu8XT5gChIyVVBqv6gITyFJzYKWGY3FBiDFHax5xugifqCHPHJDIXoqKLTTuGN
YF+xvmG2NiXH+TMAgTjtjrLIiCXrQxT7Z4RfjPdL3R2es1C5Nsy7QURWrZU/sloB
wfIZZT/TKzYJYXuT3CG9OFRf8l0qnASdQ2MPkh/XkaKBayJXYgaCMIO2zGD30z6b
v8Ep+YlvMH6ZZMeGqBX5UdiZKpqpa564KKPwIwEq837ToSjwddXCHm+yEBZMldou
N1w2+ZwHpOBvhsgYlWH2WQw5tK95ocJhDqQV2+vAtIwSHSgfNulSjOyh8CXDOK5X
qxIXouUVTDu+Lzu6DAiDzdWHHvs/LuqHb82wnZbjl3LkqMZgVjDX7nzX1cZqPT5K
1hoq9OolCgZzAIqxJbO4pqAkwfOjgp4MAkI3w0rU/k7IxB8kax+DyJv9SVrahRUX
I9N89YO/tmHQtTYtPAvLvI4HUGEniS6JCnOwoEjBdSZizAkRJK9Wn00YJYMMbytk
mAAxK4GPFEgHTfPiQgkR2cZfa/JZud6CFVZ7lNbYSILQy1icZstS7RkQfdAVjtp+
XFC0E0CO5LNcYTgyrH/k1mBVifjpoqpo5Cw1MPWIZzf+LidqnYoxmTALIweA6uH+
rtGKNxBIl71kzwn4uuRdiImxnnCl8oMKlqicFJTiepLsoPiCXMo+ASXBZ7vgZa2W
4mwOemZdLUN/jSXaX9dDNqjiBtAl61eqmD7zyyNbo4p+jHDp/AripEwMvcMzEEKR
cJ7hAnbQjnopPEcZkQOjbH2R1/sjPkO3hhkj0nSmnFc87gYZvvhNlXvtn1Q9YylX
Z/4fV1zmo1AZUfggct1okF6s+PYsCInWF+5PUKZpkfm5xYCUoDe//vImZr9HC7y/
A1sM4fQGgMdAkb7H2BCrJD2SJVapE58VFpFdBskGgqPEbmDRR0C0AegRTJX8h4wB
o3ScYb7oaY75XCGhFl2S0MbTNhHj4aWCOeRBj5kwTxDFIWsTulTTWO+ihXPxCDLt
dUZbGHt5gs1nKdF7H7n6bkxSbrtXTSRevEq/oeVDA1HQFJmSQhn4z94pMSFGGGlU
izVt/esC3YQJM2c+vvwa0dxE7wLf8l6Pt0iKmLVBH+bquzQ0W2BHiz/YlpSCioVz
5ZlRTDwW5eIvuTN8mVBi+MQYSBmZsaxB1yhyufaYBii++afDy6hVVWCGjwQR4c73
4rVtQ4cCnUDVt8egSvvWzVrzPLlZulg3kSDsLx16dJ/x8pdwRKRjMckRWxUWV/BK
jBcmcql6xsQV9pHUTmVP3yv+UhAZubDCa3LxsLNUIE1l0GYr9ppe3DBII3NbWwMg
/4OIL5KwwCPTmtl69ihVkNqBr3TmoYMZ996eqdO/Qixg4xuOel0eif+9VeMKUPXB
M75TRCWNJ9kGXIP1B5hCV7wRyALIzyv5fjEfca8lFPI3GLz5tIi5WLp/dM+2iHEO
6kU74jCKgNAsii0vrlwXJ2/PlK3SEPqQGOTUSK68NfCjtP7s+6nXhdDZB7ZLWyQS
51/+wRRe6LBiShQrw0qc+UFUv8MSrchED25YF2QaO9/k/vnjWC+w6Y9isoZ+K7+L
LSC47XK7H+LjeYXdyVQoIGx8n1qwO95WXiNEZtI94rCwYJ+bLTKkQHvSuXNsih9k
53BWabjMAROciUjrTlF8np1uIHYJXTNSrciXyy0TmE8ePLePWFRKgodcw+7xpVz9
N6OePA65U/jUMPaB/yz221qG0HjInWXKsgeEy2VmWkwTb7rV2+6ijO7wDL/QkcT7
IbrmdQrKvRAyZRb8VF25xemN7yP4S/74vCtGfbsmrJUrJrsgWQphxbIJxm7udwug
0n0smR2d31dUvTrI0l2s8miJjP7ZT1SykEBmX4weNnOMKuYrUoUXZ3YKv2Fqp7Xv
UmXyvIA+fCeZMdWAd1X8fsk1Nd9QCtvUg50ROLekLpQMGZapbhmo7o/GajOomwRZ
NgqvE3VS3bR8q9LDR/PVmLu5TWPY1oRY++Uarztw6HTM7LVm1Ovm4MBDo3E95w/P
FgOGrLCst54c11CkJBhZGCd2k8su7FLbAN1GTPK/qHWhDyatbx5W1rEPsY+joJzF
cNkrxeg67jHH9d9eob2ueHHpwu/GAHIxfWNI9TSG/QauY/QU6WpevlBpMTe8an+E
DdM2nxhbRXhlrCAt9swDEZAFqYhD/3QPIlEI13rolBvcV2hJOZ8m/rpPPWZJH5mH
tb73ygGbz5rt5zfri4KUtizBaIPIYY1CR/sGJ/dlUtgQQjTCHXvUtZ92QfyjYRaC
TaqwHNAGSz2b/gA4ke9xNfESuL/6bzyqey0aQ8T8kJ04uWA6XmRHKMTEGSM4nMQL
SIPt1bz5C051tkLn0tFcyygVUyFam0IncYu1IRWGupC4dyo3D+lq4DJJeTbecff9
m5UkuikuDo1bCYMh411qcmZRZNdQVoyUd4wKfGVi7jV6hBfrFTyL9MlAVJzpAH45
RAJ1qHyY7W9MWjNhWhf50wZKVFECcmg3OFn+uHh4RgHCwxwqRVQjEyC2TOZNR8ZF
p5jpIZsdjFddq08bOWU0oWjngQn/hPjC0JeovfY5j9NbTMtvOKijcOi7pwTaaCxV
yfDkgzawNESoY2WzXkjD74sGu1uBoALM/wwRCbu7nIWaH+AtgTiOntkuFCkX6Npx
FSOTMChLnoxuhOSY0MW0jL0fqN4UJXsv/+4N1sIpKSqV5yWl9CCAkXKIrAQxav+X
bp7nwx2VYe5dB2eCjzG+t31ylULncU0zvXNROuXSve9/15JTS7/I/6IsvT9J52oZ
KRV+bazCLJF02/Kml6XOfrrDLGSBtxCFxQk4zMqzdwHYYV/8Y7mjc5H4iiIEEn6U
uBYJkAYz2GAgqghrSyTgf9chAaC45pL63Y8UoP4qF6i20+qEN/BNAD2i+1Ev196o
YQ31PARbI8/thlzainFfsfsjGY3F/0dYwsxTfCsuFn0zE31fOXo5My4a0h2gj6Ag
D7b6CXIo7NP02D7WqmN30n75j1blWRTlxcSuvSC3aOfWm79POYvJiyoYYa5sT+rS
4eNP93E+6Ju4MbO3FzK/sGpHqkPMmqmkZDzbBTFm1RJHMuDyyUfW1a72dbGILotr
FDG5wL0KXnkUIUj9UgM4kjsv7Do7KIhHTvO503zOZae6G28Ujrds/JW6LSgZURoo
q1Xv4JOE/SX5+rAlKsraOR3KMSjewEgFVHncefUpqcv32P9sIQtel2eE2Sa29lLS
C1Zm64lkDNmQTsSKGXB+IqxGCNSH9H2gp/qdUf5N7SMweNYceo0yNynazpa5b98+
bSfc4inPprYq6e/BD4dMAbAO6JHS+YnfufEdtQfmYw+rvYTw4mRNPly2XmzATm2X
Lxh9+YM+afocVhj1LYjEWjT2wLYjBeYeDqA8uAGD99XNdoufJ50YYocWVfc7ULYz
qXFlyT5nm+1pLIvOLpSDkyU6pv2cOZS8GLuP1/yHBsdVoLxvpyOUAX3AmRz26CNl
gZqhcBYp74AjDUrT19CAlBEnEznfgIldq1rRSg0ipKsBFx+QeVjkTZD+f145eepV
n4pA2KiJwdFpUatjaNj2CK4TjV3FIUATsKCqQhmGTZmv2YGAePBDNbWIJZmccNf0
Rhw00lBFOjrIHNJDOqDHrZY2LLXZPUGsJqQapaJ++p6XdBxoUtbrNVCqNEOxyg8K
b81xJR3+in9nYIYTPJEmGDcgpW8UUidc9jfWDHzyro4N9Nax2EkiisQv4PYcW3bb
ATjYAYrCFgJjzZk1Nbvx7S5D9E/Dqls9Z1CpnSYlYWYOiLQPriHv0wfJ8bXaBHdD
A7S3D/JxtE1PqR9t//nwqqRlLWEO8EejZgfMsIEqS9rKA2krQDp0mlNh31EK1g9B
IYAUms9GMvI5XuroxUYhVnAm24X4oijO3YmhyLrjXwmKOKnoarxV0aB0+TQpzy3j
/9SD1r0dctm0VqJ6mA78myCW/UQLsiyrdD6ensEUTwpBBaZH67bpt3E6egSVO5j9
WRVn84f8+aCGKtsmh5DquhhWoEZ8eQKnvdugkMSweTsZOofvCtkeQFyX84Tg97Pp
7DOBqlPBrAejn/3zzNizIYU6dzP8rMctEGecjvpwp8r/mcP/WudeKlugmMLWBLVj
+mINV7l7763VMyfmuINlea4ctd1V4vmbk8InXbW58+UJGiGzCYEfkIt8PTAf33dq
ObgtncDElDblzdpS0/q5YBWpNw1fVpel2cBJKToZINBsSQ3jaYSqjI2DwTUaqKq1
w35HLGPK2YuATpJeC19qLog98p1UvgESxYNn45iSgltm3xHsFXNZO0ANiyVlXWxs
XF2VuSNr7VZKe38l7KTk8gIJBQuFXPHx/HtheLckFIpkP+8k5vCgPPcOTmqEmiEL
6ohz28V6R8XNUfmyNCEn/GVmZ76qrumEjbXVJhHUqK/lrAC342pZ03aa5nODshpK
sb9BHu1487WZUSLmw63aVIA+/wrn83S7AuTnuNPLHv1wBygIeeIlG6nKcsS9EHf6
yIj5m5Rg5Tj1oFPzsi9Tbar6TIbdj1RoRirpumEZYi0eYLUOU4/DG30vHyQYJOVC
5gGsyk1qnNQgtQvvfsd62uRSWMTmAi/iiJzSY5Jdy11aWaF/Gv6YO9Ju0s0EoVZG
xXhvkBOUOMB85BPQnkqpmJP/+QBkwZbqmHkXDCmRjDswBaG7L4W6f6p7ayVPW1Px
uqXFKrNBgCy2lH69V0fCf/WxkF4JBVUrcGKps1YzSTLjr2YBZZJG34KSiwT/LQAj
AbTMJxTdGvnFcIk5rZvSR+5troIvxFEOVx9UISLfac/AvqCgIv5/ve3gTQtYMsSw
HiCg0Gq1fpAGtO7ZgGWL8Z/dxwekGRupJJuQdRqjbVbnHV670y3BoII7WUPmcfHA
8fjd8PilI9imtB4MRK2+j9RkvtfBzM/0QyG/66hd0ScrnYCl6SMHMu4pEY9CyFHd
zUjobVG+E92buI1JLg3tllIN40RiPOEYyPMR84BUyb1xLzHPR1BQD6JZFz1ny97M
quPPoOLcRFTfNPqds7qBF4ty10alB92efBbecoh5w9CTQq/+R64bu5Pp3g29nDlX
bxm7ecnlYikeuHMRW+HNPV4o4jCTzydm2VAXQa0K5mhPnUiJ2QEVgbo3AeaxvZup
zve6ewTwswvC/TCmFekbUT1I5eHZxfhvlmJgtNtHezLFauBok/xzW5ijTj8gmK08
sasqCB+1wVPsQ+6vnHWOlRg30IGtpmNzU3+4flEVyoGLnXjIsvCfZFVZ7heKMNmc
/ifVIF51snZsfQtyBlRzZYsgUeiyQYPyEg5rBY2k4GiloxGq2ntd5578sCDPMCux
cDL3zlKRH1LVZWQ7R3adAkPbLVnWvPwsRaI52VjtizF/YP0/lsOPOZ4SzM6Tr1+b
Ki3y25ACKM3YhJroBGX9ec3PpJ7OZzeTT16LYx35cJKSWSYf6BZibl4UJVp/znQl
OUKaVXhhcwcQIw8VaYrAO5cdBtZxPcrUWnROuVtLCjGK3veT3YsL0dn2yFqXYXir
IkYOZ5Amv8dq4X+WPSlvbnLhGL+hOdILdLPBHdn94NEkMFPjgb8CbKvL9IgcQjeL
wtLjFiODGENPX4jkQOMa6ccJU2wgeJfbeBj4dBi6q3KZNRHVH7TyCDUGiHtzlVZp
VZWdDmCr1HsBQELerzwswqUqny45TZFeqHoSiUGzlCiq2WE0HdtPokl3Oh5yEA3d
WunZM6Ad3QKPw57u8B+gLXnOw/Sir9hrOU+YHIilKjdiwE3FepOliTT4F2IyMKo8
DwrBXn60+2gaNROCRbiuibiPhnCUnvFVndPykHwOgR4V25JeVw9lCUvtjGgHTUkK
ZHI/rWh3lBxn9z63K8jxxnrsdwPKvOSVMyVctnZeERlav0MHk6zWAbI1qMw2GMma
plVnlL4xBObOVrJxN1cm+q6Hwf83KQ6KsQ/KEgR82b8tskp3gjZYedwby0CPNDJr
Os6aY6NfIrGBDQRJ5xoAod60biJJGYr4Wv7uFbvEF1nBxX85huHPqL9Yw132/prr
bdwRowzB8bKJUy94gDiStZKVQKAiUogS+hRtvY8FuuBySAsBTtuqO0/AOKqSoXWu
zgjfvt010ChuYbbtnuZ4bdeKO4eIN1B7qzKtMb2PIs0KZ9TXL3TduzZO5XAqZhSV
WwSGejL1kp6NOAEIFu5uch6x7eGIyJkzj7FR3xFTf06CBmxgcAMJZHtcMrbItlhg
0RDZxseN6MVtukhSj/WOJA7MV9+64wpP4ugoTYgh1HXKl6VxXoa9gmYy3T+f+hiN
rTpm/o7gQIs0vAjGavwqxReYdxPe/FdQQ98C2aqewXFMTy2URSD+EAqU/1kWfNik
vmff64BfZBN76Etq0e1EZIP8JfiGHLccrSgFAeOW/90eGjNoj0zZ1K5Q7t7cqvwu
vU/yMT+8VH+M/FDdmRudz4Dvlu6mIs1q1ozdviMufwhEDzCduv1+zc52+PirSpPO
pobbNzUDC3a5dr5gBWXksxMJi9gVd7FS6RRj7p0tCxfP4vhx6OQvzdkk548PxEAE
O8HNQb6DP3SZwEYWvXckB3AugS+aIkRKn/epkDvkbQGT+DLsnVXz1y74qT/nX60a
Ns7OzX83/tdKAjJcIOcCqH76GDvf8kZ+Yq1QjsFxnAQovU9k+BCmlTpgKzQoLxWf
LCwum8EvESSlNqM0JS4tF0/RUBHGJU+waWhbN1wtkf0RzB0H9KqsiqhCr/fmp19O
X3GZb4QlqjFp5XQ7QxPvFDFHPUXCstCUy3ZYm46SN6IJuhldKRl65UMvvI+VHsgD
IBUAsHQEKBpRYC6d9xKbpVI4l/ybtSONBX+ctwtcOXOvftOYmgLVwKacLWmJzhB9
LfY6mYW0GLw6OwRjvBdHCWfbQUGvQb5p6NqRvv9DpwbttpIWFf0E+0rZg+9GP7q3
iAN250vfZ3TtISVCbvfKS/shhDsfag22XSqBRJvvoEZpBMJFiFOlDkdkbh9hPX3G
VO4pvVmP2gEe260JRKu1KStADxnwBfboiHSiea7VGbWl+GWsr0S5S5iMuJgmOP91
zgIK8uZn7LMTUcbmK7OXnEeacGymI0k7/rzpAjqOnQy5PLnfqdn/H1CqNu2moUY0
5Fb+FbSQ6AhWj2x5hYc8p4u71HepYsitvxKfnF+1owOrnESAW7lWvcpnVNmSs49K
NvPcGZM45UVkE22v5CQwiKOT0SdLwtWj3j7RYdRazOYgmJjAzeMZTBDcsCgUkpUb
XHsjz2kgvoxdH336DJ3fz/3h9QhrbKRPobGRbRMOUfqlh5DS6/u8rObjEZ8D+p3E
IZQ0ajrwi1ROte3UaKS4AVp/TxjyaxjroM5a/cfyeG6RZVbeg6gK0LG6r4146BZs
hYeZEMkNWnf5K2g+2G3fM/De3DtCEmUfKzOFYXKyGIErceo0uz7a/tuFaTjgKFfY
kxgzEj986j0M3unBDuBA3xLiB6G+JCJ7SQ6KqguIub6ZhHVPZOqhPmicSBGEXOMq
61pM9RqPYv/eS9Y5YwzH0wk0VZ6uKnsNwx34H7soavUOb4uPs6vQYxphioxeeGP4
XNkE+mjgHFefCeZ0xLtCMqnudlThvwy0C2HcoDUo3yZTU+H7OF+/A7ioQ643TaSw
VB5WYyHgrHOmoLqK7oosch6hvYb9eVjA4IuEknvEY7ArVy+ZQMgUpTWKUmpz2bpI
dOjPn0cTZ9M7odepn50rF4YlwkdHzvkag0gvAnFvABu5693WVYQdUhFx/1aMI68F
QFOv7pS7mAFa1XA0GJlxTo30CBu4siiyDeAw60qn7ZNp8//xr28AdcWL2tcmGoFt
voWZMRnPOExL93EY7KBaEh5RDRdMcGdZ2jue+zvJwP8JTHl/BvJC/Ew3AA+VLlxs
QSH3UKlYPWVfrRTf29YOZ42yhonLlNIVraO14E3Vq0EmICH9Trlj1RC6HmJRAuUS
zMNMT6VRQyyD9Fk2moeTxLzv1aSVNEkJv2yis6wbTgnQDtA5yBUN/7WIcOceGWNh
BUFgJOCrKb4iIgiLcMShKoatO+23qJKtV2CbQ8kJWmQkhou5ALMeozRZIiqA+g2r
kQyyYlBmPXwGXKF5DwVG9lHGNbW5A3od3s2WlV2+FezRnQM0j2oAhsRLxs4Izwmo
G/Q/wyPztq8/AV8W9i6YzkztqoWzpsf1F8v0AtUh/clIU8JgmGVGDgpeH4vn4iK1
Z+H2aCSKKIrZeXfyHiunQQNLyHzwYomPb6py8cjER7lb3NS0165G4cFVxi77Ljy0
ZaGyA2DJwRE8Iv6k8VtRtlFVQHYVDMnYc7fITG6HU/XFKlHClH5XHuRV4WeUFpow
tTl+iqp+rip5hQiORy+NhovbfEn57UUNvCH3MjeRLq8IsL69vWFYAvSyhdo8NNsU
Af3ML1HgnYxjoCbjL/yBCg3SzA0g9YrGsTbmAHm4BUWbdDi0X3W+xcJS8kFiRIJR
LwuE384UdO0ui2nf5v5TKsuPnM60L9z5fxd2jGX8SlnLHNEgISBbwR1xuMIdfGRw
11DlJiWvcz4T9pTzfisriBrjhBagoT+U9ICBKkhdr2cVEx2CnlVaZL0eaw5j37Sv
t6m6Pagft7oauZqnY232+l531QTW0A+IeMmnrPP/DJu10kKyr2IQrh23NkqtgqPv
1uab6XsAKHlUtMGGvhcKRiEPk5p3bl22p2ln43Tp5o27K4IXc4jF2ZGug5BNBr2U
nPzEcqHBBetIDX7suoZatTZS+21WXKGQPjxyrTBdAm0GHjPjvAi5ulMOEeNQ9Gxs
+E6WuuBWDrVJrJv3b8rx2MMSRGbjgpFl2OFjx+YA8Mo9xsvrL/vVRyALKXgf8csd
7VgM803j1xrksr+c6EMnf7b1Xkt74T4exDAKMhrtnUN9bkw8NFHcJro328cXb0X9
W9eyJue4aSjVitqX8b+iD2rxM2QC5l7MKPYtl8jV5yE9CEGS000eBgMA5x5lAcy0
vux9ET+z6kjEJDm36tb21EPpReDZL6MHOMRTIdbOxIZeL13u/ItHQSLsrRYlJCst
Ti4H18ZxcVPz8sOmSxHDnA+z6fvaigOE6bMKI3kEPOZ5Z86NucQhm6hv/APP4cnE
5NC0gzQbxe4iUjLafNWNWmoUB8VQ2nAI/poLjkDR+5FEoJ75PaURgYY0S8zYES3A
1Q9em0iyWakW2deCkty8wcJ+zl38oR5MEinH+JcZhszfn4aefWFXEyO7d8VcKSg6
6bfmhePm8DMM/737aH8yo6Svwt1rpzBWRCIhVCFGxoNPL2mpKYC/t1or0hfFg4L0
WmE9lt3fMprTOUqvYwfca0o64XfidHuwebxOFgV+mn7M1cseGHktDAEHkFVsTF7Y
MJpwYADp00YvPl17VtPRHwmAIjf+7KRPPdDiBR98HPT1baJviwPNFJfEYDry5OgX
WEoAoFTS4909qWobcNfj3Is9jgSSN5Zw0ILOWgwsrc7m8LrlaaiwgJdndZgdPKE2
7E12U8G+21K3Q544aNAVggK74RbiWV4/w1Umw9gsj48teUoa5hQBKfyVVUliVfBh
sxnq3mmMiuz33Bzimvjxu8SJ1jJNgiq+Vd15TJflrMQfIjY06Rfruyq36scr/qeK
cM+f3aDnzyV+BbJiHKuBymor25tCA9F1JMxS1qq/qOVpuHr0ig+tWM2lsl08nejm
REX5WI4u5/3H31snH3SZYMY66KjEkimAdJObUP34THMaBmRutRp6mlAv2490sKcF
vr+nk1M1hxcokskPx/eaK21dyHtGYYLj5fZgBcup3YSCZ8WRiry5n+zZ3cfH/KQr
2us4BlGy8GubTMLgziaEu8t9aVx3C4ka4smB+S1ZOlorixZrzK1FQLn2sbRTQf0S
aae4xJq6i5J6dQJq4Rtl5+tGjQAs2KOr6rxDqB9hUS4hLdDTcQh3p5msD6Pbbwpw
X7P5xBfz2eDFCJ7MZfSUTQANN5jm1cmgdVo4Md4Lj+lnmG2sF6FDpohozvzpJWdu
X6MlnPCJhZynB/JoJKuOZDbOr/TZMZX0qBkzvjMx2RVHlDToq9GsUZKHDQJJqBtQ
ByNyKZNQpc9qI2PMxYEb+9tk8muBR7pLrrOjgcjfe9+Be2Iy9tURsXiau8AsAbR1
ffXYr0mMuBjsTqSoYsdFr/YJDPtbYyEG2mFFX6P9sfHZmwuMuIQdMJoWe7/rZhYp
88CEEEcy57vx/bu2SQoQ4H34S2msjkMO2L6CtkeWpWhBtmWUUyV9z8es6HOot70D
utgMnnlnE2pSzHGLeVFSi4Vm08DMw9W8PmmIx5RLIHvPn3pqan7yFdp+e4c100Br
nlpMuzQB76zLIHiVl7YmZSJ1ZLsYnxOgA6z0AdF4xoN6efKWzJ0dEZJ0lFWlWSBT
Lnoi57bBHVbLImdicr54QzJe2aMb3uomjQPTyhzPyy34/34y8tdhn+OD1lsDcK0T
6ysZD++lAWHV5YEOrnQmtJ7Z4w5U7aXN2zGc9thaXNDDGA5/hmHVRy8iNweN55tZ
JRvM+3rqhwQxZhL1HsKx7+JpurwmApaR2bg4Fjd9PRRFwEQmm3xsjv17lLKinE43
DMu5WIJkHHS+iObQfOnaU5cxVPiRFJt9pYsUMo5bXaQNKeopOyR+VEW8r+P7b7h/
Wp7YGkz94yo1GcGtmRZ5ZJcyzcRHBmiCVriZQycDZC7ml1wIavptSu81R6iUAvsQ
w53eP4IN5hK4kpryIc4E2Y1pbQDs5Ia+ar0Jjg4ZKwRyTS8M2vxFTjBSN0bEBccx
25umoYeDpZm2mn4cDKc18h2rmyRJ3KCk2W+jB9e3HbqD4BMHrx1OUs8JlpaKu8/A
RMGV6N0Mzfnn6lf0YQTho4VFVDxebgXspEK+RaGmi+YaCTmET/To0ueQ8g4EP8Dl
d6HeQXIhVq/DRBfWLJDliw/qN3gMSgTwyGwFtv8D67dIS4ReoQQ9rihCe3DwP3Ke
nJP2hhCJAtM1q7sJOwbgvsRWryI555tgnxR0njJBsgrKLTkQsXq//suGycrRAxwl
3LIlA7ewpYoe41V/za8jjzBYpx/Whr7eIJBgoH7d/anPURbkexsT69Dmgsyx6xRi
AcYNRII6K153pv0tA1wmEWX1p7qBlgBdBy9f+K1SCSAGUBCX6KrvlcGD1sVxQoC7
R3AImmS6/M/AOdFJJUQGQ9ybQlP6RuNBHuvz9f2qqZVkIdEVP/xWLr5Az9235sUh
Q4Tj1tVHSVxjw810w8N/e427TDgN9hbDn+M+N+DBirOP+hb7WAoDAJEp/hOuUZZq
WR9aef0et+t6OmP9JXFGSJrsa8Pk4fg1TxWPW1sEVtEtErHQTcfD3xfkL9nGLJv2
TFkmWVLr26cXrbGYnJyoHuFBnuUX8KMJTHXswx8cqFkTNWg2XsIOEX/D9T45EVNR
8S3okNWKvXnRJpZ1lS3sQnCd8LsMyPZOG2+m3a9dN6jvmCM2Z2SLtj1592HC7Znq
1EHpCZorwlumiqTqbR50U9NGPQSAIzE+dG38hdXnVZO2GvuXMVslF4563cVqUiy0
Fz8waexepqCZlnG012+CGazrJF6d2Z/0Ov0bJ3tHyCu2QUpZTrxd87oC2QtdpsW6
vPYPpx+zFS/8/NvCoE03GDPhics1c9IqNFAskNVww8sWqnfmeNjGJimaFdr5Y5MJ
NPBTQFDe6BnjuVDKGzruYr5Io0NFzuOTh//mPw+bfTktv25urdK44wGBrTIFrkYl
57fHWzuyJm86BWFGDri9gVwiKFZAozKhwMMUX6WxAVL6BuGTCuc0Zzf6YypB4A9R
L4XuqXIfRuz3gj63qoCf310ZIkMRP7ii1NcLZrcGdmYyR+mFalYG1XlZ63jTgTb8
WCpOpd+us+xkhBN7JBZueroqFNu/Pnb4nDEr43IkYqXnXZIg83aCOmZqqjNXEKna
DZPc2+YRL7LO2DWa3uiRrIXhKcNrmEQUskv9IdThbhvgi7Ke3GoHu48uBm3KWCKN
cToNDoSROj230FlV727mo/QhRxjg+P5+6SbMODXu1CdaQktyaOy2x5Rte/OlmETE
CvqNeTNSyPi6f7JTig/JRblERVDtotWReJIDLt1ZoHm6jzDi2vRdNiLvYDeh5piz
FMEky905dWUCToHTslmLmEe280lQJV0no+C0asQybDMf3TkI/kDkmzC3/5oYpiA7
yQrMKJHI0jQQqelm9+oWqdH/rxJxQDOdA12OXGoeNsyVvos0gVAtRzICw2iaJfZE
z4A35MdgbxkH/NZpJzMF1o4Ct7uXeJ2AXshglscjayjul/1K7gFaC/mKRnfqpc/c
0xVrEjpomhA86uV5AUP/3DWCP9sapRbwAeqi9vvtJmbosTxSOGpeh1EduE4jMtMk
powddcJElW1JsXEveglf3HZxYNyo3hql8Aru7e6xUFohnXXakRrUbJLqfcI1JCbF
Wu1Z/gYYYW7JWIg/3tO7+XtIu7RPrO3rLQS90loliXI4nbU8+dolu887spIdl+fe
FAqXqlZ5LEJINb+iYd2ZJOOG4v64tp2Wd+9PR1a80IpT+mpEshoI7lfwmPDo+rte
g2F0FvM3fo7Hq+BByTlJUiJ18h/UyL/s8am79rx0HnItvnmwq17bxhyNMdi4qY9f
wupuaaD19wwJcidrKeTMc4mYoh2ff2/bAcOooIIJvGO3mBZXnVt+ACw9A3tV3nmc
eXAdrXLd4e+73o1ilnrfz/YF8AYbjn0ZqEoX0/ZaNUjKP8AHRLb3PzXdb/ca17pD
XYdCtutit+JlUiZVgkdlWFE/fPXGnBgwuNKhs5uGOhQximMI1pplpmZCa9+l6wgz
70Him7JdIS4YfgZQgvSSNjrbvhrMkDJ2LKy4k0VHUvgyalhBZtm3SVPDzD3bv2si
0+HZ0jzFplBztVn3w5CUtdIGlAfV3ZE7ciHqeYHxHbNG1HCtF8oqODvJG/3dSpLR
juG6B/y21f/9rDxkJDY53qWQC8GBahQ5KhO/6DduC2/VcOFMxtiovWdY9skrjMKf
Z2KikrhOoiEk0Xh7VYcWkmzj9DlZD7iQABH0+iIbYGcFcVTxZ2k2m40jN26NwEtd
jHTArIZ8OHPFsZrV8YfIta4UNaXRdFhI2rlOPCEdZKqYYHy++81+tty4DHQtdtcD
wGE/cQF3mG7j6D25e+hr2H9WLJ0ic9yfQ3Cv0R87yDWIUKKbDi+VW5ccMPYZ233z
MuW5SCJ7vRts0rAPbZbU+OysOQ/l++FEY6DE7PYJ/0fgKwR3Munr0TC4D242iABR
aiPgmBsYKxBaFKgTI1uxpifeIqOHOFOcI1REt5Jw1tf9M1vhmYTVTrA5kHR6aKKL
/5kDroOEc2hFhJuGHbgOyd/octvPmLu0yp8JfuT0KuYPnYT/P8wo8/5DRuqaQShM
qy1xukxk9pbzt8jIUs6MUbOGHQ9AAsfwkXAxsZa/rySx+CN6W8FuxGdTbmzSZutM
i4iRDDn6uzqzhJMNrCmtRcCU2IdIwpVwag7yDRWz86rzIRWny8dba/zGyO65gRB+
XCjUPeNrItByfOFAKVTTfEmjlV2HP1QzEJISUyAhnDuLDTEh8ibCmR/Ci5JzKF4j
O6NXS4/bTv6Me7jyccbBSDWQCAUtrQjnjbxAuh1eYOA/aU63JSw39M2p/wziuEAa
bFPhBH7ZSaj17ifM4legYETX/SjOraY8lRmdqtmQmDZdDms+eBzSVJr3OITQVNt9
qe8WmtQFVAkI1uDo9D14eXPqy/p+ocnv8bQ6eSY/ZgGC1BoHcZlg9SllOUTiPaTT
FRvmb3jB/Gk0eQCstxjFMDbNnwiWhkm09LTutIieulT8xsLTZj02W+zMeKtZGVFe
4JWASzwGMxUpNtoBfqJO38D2OzetkWZjSG/pj4pF5DzY2CAhvM7W2P38Gms2WvlA
6lpT8OR6B47fyhd7aN3ReT2/kownhhZPlhAyzzQetaB0cRs3D2k/2SIcvsN2KB6D
Gasali9do8crE/6qO7xeFDBDVKXyhHsY1tzM6YmX9xD51lYpOHLluPJtf/cnILPs
VSNf7nyK1aCM6KCWu/FZ8SFLSTeKREOs8uxEo62osutmK4meP3dRZkgwCUJSDnZ5
H8pWHZAIMhoPYf7iYGilzEx6hb/JUwnXAu7ijV7hubuc2dW7diWs7VMIr82Mg+LA
AaBnS/MiwkeUpQQs93+FDBFSgR7fo2mXQl+1bQFJQ8lGBVddX4IZEINMG8rFtica
xYWcxfoyrlZJZSCWgfjiLJXKaB3vUW5JnBQcJoq0iBtokjngnlcHWx3Y+Gofq6rr
IhkYINDpObGazpcmJmj5XNmkCQXvFA9oDsdNtTtQyrdj9RE1H84STp1uODqzeMie
JCt0uprhBdPrtlI5jFB3oesxEpfn0lA0amve+IWnYiOInDsKc5k1rAfjdkHt8ogE
KXt1bA8bithx5Fp01wp8MBiDA6b09pXwPWGjNQHpkUT9Z3/tRwRpgEZAqJ5wKPb2
16XA16pIHE/3rpRDRgY3daAfyR8npL4wzk6LrPOHJae0Kmpcs02kXI/wtcZ8MZAi
SKdT5xRA3u/YxRWntxNJP4NIYaR/LZ1tJLlobm78DBrmP1lXflID6YIRSbGS1u1F
X4lQdhgh4/N7aJ0OKnywpdv3WzOtMm7y0oyUK6KqY7pwWX7plSMrgrr2y1EB+6sw
nazofeg+TV7QYBllz7ewzbLJNfZ33mfGYC2ZQ8kBJwtrOMk9ClKhoLI57WZdzmT/
taWmmdkgBvxRxNrwPk0lnth3nrhReXHdT1yKR3JTR6cgngqaM6YJ6kIC6DTi2Ure
lJvXh4M00tHHfnBXt3eckwq7Y3hA2F7bWSqyRm5oS110J+lOAPum1guo5kj5icAa
DI3lbEs3cLE0Zhe4RYjjFdhSPzV1tDcUpbq5pZouRe0ciAuf3nTF3ROYK3fhbf1W
BMqUtX5NDh2e2LZOBOh1Vh2VnwwBgqXBke4OgOFkahh21UOO4EqRU+2qALhH9UWw
dx62+VKAI25kfTPmAjIEA4nlLnPsRt8fTyDd3fNeD2w37n7T05P7SYt5BQ79buNC
Uvz3yXku9/bAg3sICzz8g8L9FgdQP2lEgowGnCWDbgvb2lcVFAETAqyOe/yijFR1
ixi+rEvnLpYwwKao2E1wyw6uZiTrwnpL6gRlhdm0o6zdgQkd3gwB6a6EGcYvqOCB
PCKXCx5cK89/w/4xSZ93QSNYwHfJ3qsLCVm4Gj+TiqVtDlrDXVzEPdF4iHFuzXns
yIzhg0S5sbPrSC1X0dfsUAAu0hcBt8MD6C12h7F9VyB3I+X3Hq51WbTvPverfW2m
REnDRczA8MFIRzNuKJMocGzfiddCRug1EoyWf3obcWsJrWM7qQHcGp5pWoBDIovv
F1atWor9deO8X34s4rEDz5W/YARwBBG6b6RrgssRuqmvViRyzO/kjMDagxqN8kNf
cv0yRCSjjCdJp5NxSieiL4EOQGdIf5sysxJDnXE91Z1UGBivmoQyoqDikMqdc+vG
V+cPUr+u7UvFJjRVffTgApAgo0ZF2RMzoB1tDmvulFMteZk8DWRRjs/feyjITRbZ
mgJuUiwqVoIETjJ1oM77dX4wCzW67cZea3SzGlmcU5CK0twfzkvsV5bEhrTdZxyS
/CG22hdRFMHT888NRJwM9tbc9zuepVmmjKyyEX4NBFEiiWXHNUbpY9E7J11tRjxv
abzBIN2zEZMGpD9f9g9iqzq1zYxp8qZzEOWaFKvi9c6vQk6xu6K9NETa1tcX5Pw/
AoXrA33e5HHkKY9PC2rc8ugvNERqdWbGQLdfhUnWLzk/V9hG+v2JFoEmKoXb74ln
CfX1CFsb3ZYM9kN/HjRkn9bXcsydXoqOssMr9i8f2OhCqyAMAv0Ro1FAaxvy395S
Xy43+Jteurqu+toBNWCVk8TTh3C7ERBsQb5pE63drPowF68AIA3lwiGA9v/WKqOl
l0zbIN6c8LOvCi0Yr9veb6iKKm8LbRrrjw5cvXWPS1oErSfcZqRZCBL3ZZBL43Ei
1HG6oo2I5Q4/g66Mb/Ik97ukBNT3jvmv31Hu94Kl1XIbFMDJFpELz55fBKmyZ1V9
pI6GurmwGtcwa4B3yk1n0ldHa9666cqS4sklk/EzSGRU4dvPMjHHZbPTGVsm1c/p
T8gg/HdUeBLwvCToZfDifypHA6CzgVnjTgNaS748/GX9NoCWio0m74JnpNGicS+y
56TDf+scdJ6APZn2tw6ERqFZo02krWUCmtX663mglTP8DvyiPYUitZyVoeGkNice
EUBo2uJK6u5EXAHvDNmMyJ8mijAERB8SsREEuMcVL1IETqX3Rly0558diFLFgYay
a/mIIZz06jlsOheT3fmARhxVqDdLlBsk8xOUPoYCzmZBFSxNy1gApceEHnlswjiW
Rbxg6mSw+c4JyChd/lQwaqZQpnDRWfVK295RLcdHXYCr+cxjYAt+D5wRwaCiuWiG
lG80Ibgp44L5b33cIhMg7//2zbbkHP7rPCi6Hnu7kplcQIhvA/BKCxsHYyrig1HK
jLuz/WAA3k3pUw0i/ot9yDF6SaJans4Bru2oBPWnU++9c4aXXxmwIwLdmPLNE9g4
MsqvNaJGB73Dl+zH9e9dt8KY56yAMcjdro+hV5CW1HmCKiByudazSl2IRc5CEDZ/
QG9CAWcf8ieLeQpEkNpO720xSA4h5ost4SmIZ4k9eSQsp7eyadPy291o4NxeAZ8G
YAZ5hhj2jm9f+06nqpzNnYbvppX+dK4K2FTfx6II1MpKDd5JzkDEcJQhSOKWtRWv
kKJrKKF6PFWLFOZQFoNR7CiH0xDmZZgGLMvq6hzM2agPGuqPbEQHKv2rci0aMGcm
l1/J6P6drac960thj01h36sQ+/9UO09BHER/2Py43mNT5RYRGNoKzVEKrrHXfKi8
YkoXZ8sl0q5HXcbx2d8SkZx/mcYuafVPW/UnlsiAdwZAMgUv3/MnJU2fAb5Hf0J/
aFnWvvSMu0kxVAHHINCME3/zplgMgT31Ut+6qIQHcSYLYl+GnI5jLEIlTz0TVsQv
POSKl+oqjj7U/lavfGOZOnjAJ1l6vCCUQNERBPuXeKJC14xFX1FkVr/ffpaAT6wr
UJHAYwTatGzHaI91VFsgJxqiMyybMjhkBjBlbtSlbNBlfhXcIKnyT6TIjSR3CmTE
qrQLqLy165MMjX7I3sFBxhHYpW0pQ7fFax20IoqWcbEz8+ZdDZQTJGHcOgZS1bLw
xL8y8hdfdZ33qKUa6cxSfJg61PBa5auNn/bAFHVxja2YnBgiEbvD97a4sid1wkVv
aDS8by6cJyhDRZ7ZK8WKTxrZW8fSpyvG7ZAwoJEnPZLQLmVUPC07RCK/6aOSbYD1
15e4ulC6T2O+1VEY+A0AMb/E7D74FVC992PphB5w5r1vrfgbyUkNMeNeOmuqznfy
Usq8PutTaKWEhfoq2s+feRkFU7KyPNGeWCBLTuzJjYFVRT1VDSLaLhljUvDsUSD+
PmaxiMCDB/9TdDf75AhV6zyDj8i5h+G6F9HBS90GMXBwV8egLMGUhmPY/9b70R/Q
osLAErbTrONgoFIXTxaPN4tMP8zrKrp7IfPjJnRF3DWaHbYwTQSNT4dt1VcSML1I
N8BKIV7bZhVGEl/oWKrYfmYoNxThlUNDc1cGF5QgMD/LaZCGJdRfmABnZpPz+z1K
3Nai0wWWB+Homy9R+ZdZ4TFzScI9z3Q6nTpXbvxhD1ft7peSVYt9Nzf5SkXsh9H1
DCCsvY9wc1lV0Fh94JtsY7MaiIgyVARra1NOa6fscKZSDREBFksdnKXO6ECZERe2
cB4DiQDakvjkk4K6Xk0R3go7ScLcyFrxSCUU7yvcSSEnfPfozLPETnuhzK2j32NP
dsyRVyZIIaJQ0kx7ZxsWe6K2Stl6XQt2oUFY89+++Vqe3Re0OGjT1QMYZctmPHXN
N5Kdk2EcakmLyGobGts0FgB5fWI9/ZWvWp9uNM0nWzRbrHi/EuHu0vVM+hqKcaf3
8cahWs7N972jP2Fx3JgcWxIKsMJ9gy8NZ5OySfRpmDQqhCRaXfcDmt004OlK9Q5E
JC85oy2a1Hpuwog32QVr75BSEDoSuWd64WB8OtFDdXrBw4tS8Cr0mznXrq2smuBG
ti9gKgzvKLRQLzTAeab2QPzswkemgJOVhg3ChnmFLgaHbQPCZI3EVQS0gB4CWA37
K12lFTCj0uWdUbASV12Wxfni4u2kRrV4Abaat6m9XCbxzmMG3cl4l/ZRnnBtEczI
7z5yiP16utn8IwMy77BMwEGaUf/dwa+bomne2QcoUbxLxa+1Q9WSR3sQuAJLevYY
IYybCxAiEJ1HuDL/ULEwrcP7ZXjrQjdM8uRo7j/PHTpBFecsnQdsfNwLEn+ldxMR
2ezM9rwJ/amYIwKQVis52++KXHvhARoJevjDVhp442ZNnMAIL5fPDxqAEH2jJ4Xg
ar9CjfvfBFMcHay5QQh6ItOsIVWoCni+sFH5spIBFLiE4dTirXR7WndWBbe9PF+J
QmGsh4nBSW+GUauhOu9ADjC24D3mX8HnQVikhEj6taGTOJIv26GLn+dYfgWufnud
wn5OpWcJVWPDjTn2LI5Vn+XgRRbxHaFiC8GwPi0saxexX9QdawohQy2IZK+apUT6
4OvqZlABPi7qxVBSE3OH8eCipJGroZUonwhtw5gLZWtUuWX5DohlkKpIJLR6o2cL
dCfjb1Ce6Q0kp40uMm3ueZL3H7jcpTwyoySsoNmb638CBsQY3CtI6f/sHmUtghw/
w0U1bDmvLqRj6XFQAEeLpCOIznvFr1pWokY0727SNGh1uSqjVqh29zHNhloSldcP
T6k88CMJxVPLAaaN7zWL63GgY9UeBDhlZyatRMGC4uxn/uqTnJV5SQSu4iYdmudh
n03yDH51t/IAYvVgOE7dc198cRNiClyHRLq72Tca+fKz9xQRbuVugeTJJtukjUX5
xAu7mD+Ai6JJKECLocJlLM80CjBFcBiLbefTA1Kdp8F7gWsbrf55mQXZMhevt/u3
jP403Q1p/mGgONQU5sAbBbU6MQ/vQitWFJXAoaToJS8/gIwq5Ysh2ReR7nXal/yz
9ZlsH5qtUgxmvDfdyMk/+7hDjaAqz/I0aNIW6+4TByehaYCXU/PT+Qry3RnevcnK
cfkOtuuQUHA657wJ+2VUR6PUAyUNlTZk3Q43YlM/nW3rw0xCMGSAFzqzioLPM+xi
7s4CwIzZwBhWmSEZhrbQ8McnbpUwM2aXlgBM0Idog7XCN91qWlas4QTkqSyXs41Q
k7wlI9C5S0YdQZFlOhEMIQPL8nnzXjKV0xhb0oaMpqTYsJIG6BTArmEDQlQ1/gw0
t65lT6y8bll+PulY/yEufxL7fUHs7X9bLwZpMwUw8s/xFxBjws1K17m56NCXKbgX
qiQsBRqFpBOHSOrXSMvE3a5AhAsWtBp+eCXSAxWsD4E9ObnViahkCvegS06WMQg9
XVTmbkCKfl4pNLOxhvmfjqfE7TnEfuq07i2xq7qEK9Izxs26Zi6vyPeg4MzAXXt6
V8w+e1op/JZTaLySuC2TfqlLcpMzQ8R38XoTyL4kMh7UXGpH2BXdj/AhaGupaLFt
a9nfY71IwF3FMFK4j7+wYDuc7yeIHA0jG4EyK63sEUwiZAE2GVlBQYCgLj3N9RqE
UcFVleazmnUhT+hlWwh5nzvX+1EJ1Oog5TlARgM4eXwNQXCi/qO5G/fVzRjoMBXI
6wGU+0zRklJFrtjlC8aQ9ZGqdp0FMRTbunOG79GDxs5L6b6PPPM+mmFNUcx1ioS5
V0+fudEMZDSSG3pn2u3Pdzo0yxSkF0WObwSSENnwc5mc6SXd4027zj6WHVHXvUdx
AIh+V+lubOcw+dibtbsMHEWoDXs3sJ8pVKM6sjar6BqBBwapigAH7oEmxmpm+C/F
mWaiaD4+yb/BghBJeggr+unzdvKDCzKoY8HJg3spmcsZn4uj68D9MjmaRSTlz6iR
R0QUho8HsrE9mqIm1rBsSOpoma3K4g3fB1belhOibP5jFy1WmcJlrX1vObB+aFk9
gpurOBBho79XrNZqu0JrrJVOl7nzP3D5N+HJ0kdoi1B1GsUAi10u7jf4GwfP8PxS
1YVJRtfCm2jkPs0WWfKmsyZxhGc31nvJKMUJFgZuh4PK7Yh4Z12Ob3oxlWddwISq
pmR6Tk8CNCD4QayoA6O2fKObUZC4rmpXN7BbPZ30rqNBSPAGVZUO6c+9dR+TzVis
XVtmOGczHSFyoUyYGvBTtRTEIk/3y0u8zOHLAO43pWv8d6FBd0TO4v6Y5CgnxwQM
YGBY+eu4T2Bmk3zamXgtvZpsiOmcKxLTN5DDtgiAQjCU8SQ1t5Cjv5HBJk1Bs2FE
EQEEJvS+lY11nYwEdVV2IACYnJTNkX2HdvU/eCqYm2RxT1nWhr8quf+fMLw5ZEju
UHG7lSiXP6K/AVYl0kfS3xZXjG0KczVydUhsxvQ2eGApwbO/LfCMRu5A+SYovAhH
hlEjKkYiQVXaxTJwWDOzZXZWCORliDL4zkMLuMyxyD/kqHLG20YVoqQ4Cj6NiMG9
76Ldui0qmRoje/taZ3mK9C4HRJezxic1iyRdHYIznVsi9P0/deXC+SieukGJNzw/
Ec6Wqc30rroxtVHggw+qiSbJ7O5rYKEIBU9Gz+W2Ln8ObaWl2HbTu8wEmrufLoS8
79jwRzmJKChejVoCUDAJvvOdCL3xEk7cVZTJtYucp8Xot9RnI8TaLEUKobkorApk
lYxKkmMA5ySJrbejW67vz5aDW0+EVCiM5QARpb5qZpRIz8HWTNm1+FbjFf7dF5ej
tGu41/1Z4Zwoy1t26Wy1k8c57JhMjqRA4VszDnCw8BYhbAPQdafPk/gpm7NHUDq2
H4szCCRKYoDIwhjORUTav8+uI7ODA82dArb2BO6eUm24m/5sDhE6LRI66S/Aq+z6
+tuM7CA0Y7NhfYXOFZCMREsTOcgUw1lDZSCieR/aDin1BGIlQlScTeu36Yr7F2jU
bzxzu/bo6otZyIv3XSLud39b0FBSOfzWGVjVLvYA7IxXVBjjvBq9cB03baOQ09Fy
H3asZgfBt4922RPFNgec+Ri5SusyUx4SOCJswVceLTBjNO8NTp8MA4Tk/3TR+CZD
YXFbEg3QTKP06hKByV06uSzVjltHB5FE2XOpwgDuIZ+Ze6gXHhldiTphMXKxnkyb
Im2KnQjsUu90IOiV6YqlAc2pobYdtCT5C+F3DYNVsgPxpSpR7XwhzI/5s8IvEY1T
ASstoFo7sBsq11rcwPLv/415c2amlKu6nmFeTLpH466l7Wlkw/jpC84t0VjWIplk
0HBQaWiLiLzK4pI4eGXWCZJOCZpb4V9yi7LzIIQHgO8qZIraLHfi+ZR8binPLTEk
6bZwYZCAx9yKzCjQsPjVmCuBODTZOTae9osdWroMiTCcGC0NEOQoMKfddLRFUCvx
zLRUJVmdwP2DYOfoQoa5sxSJZ03NvbDMR7vpGYeOWdPvY0681+clW9XeqVcV8/1h
50xnivACAESQ48+i52tGF8J586GljqOcM92+LoG8H+esYIGW+bbIc9sAcutxvqib
yFFpfxydtgf+g6gF9H5MUJLYq6U1gRmz0rQ0fuh0dr7ctHZO+yYr0eOooIrONThR
iJV3Eual46U4k0qo4pICFLZ4uocn8OXnscTC/ycxuRrLDmOdkp2p+ZDUNcmwSI3D
xdZlsC4dmS79a122roo23Gob2gaiOb+3VpPVj00aOErw2vbyj5gUeEKeftZYQiQy
OsbAOg/nbBcdFylbDIN67ymZ2MiLFVg/3zufNdq62V99d316R+J8QG2rEekh/0qa
tojP+lQRPJXIckZb6A/xX6vnqLqQ/ebXtB6L5zhYOqduUytCg5ID3MtSymf22cSR
Fgd9suCD4He/yGvPJ1KTaif6+fXssFAWfgXuG2CeTRS3iVD/q5wH8YwNUt+piFWa
jnpVEOEP6HDRjFrV4gSmFPLZtQOSwDX9wgFCguTyjCbAI9Ptbv3+++2ArB2xnn5p
hw3I+SE3BekxhSTI9S6pQkKlwZJ6IOFko72Yy47/ZfQ+tDUlA2A338o1FsNtD8j7
rNc8WP9LvncLapB2MJfo0uAhW1Lalp0LmmMma1NIs/sCpByo2ChvbIb8vBKSgaCs
QRxnL5WRA6BHnsfGGd9hxo1E6c0qw/G53wTFdIkKVh9/OTjWeidojBa2o9ulte3H
85s15vPr4X5BAALps7fAToFMAeiMe1zzLSBuJWrQ/EzbuqDHAj4q5Ou3hhuTH6Ju
uvQ7fo51nqZuRlP/h9wkSWTj4Cen6eKZMVN0KCgBwD2WlbXjn7ec8uQTap/QoDAW
gjkjIkANlqPT67XGagb0mdZpFAd4YiBp0v8pYgBFW9ebBKG+hDAI9DYV7Gh9kc/D
AB8Mz+iXfJcVqWHxmbmQHvQIgJMpEtS2iaCt1pVUAzoZMXHS5di4NqVcIbSYx3RK
oeRM0LXm5gCfeK90N+iY0psuUJ9p3acqvnZW+Zzg/9Iub4RXCkOcfdodAIGxQ17M
WCqKH8Jyhd/blTsEHbWP+20WWeGZBtItc9bmfcvKjGiM0piLm2qTBicXh172+vte
lmf49p+ocUfWrjjJGLUvMym24FbbuiBhJuXCHBDHrElL0oKQ8Oqi5OPK5RxNTe++
nG3h1u3V96GSkziImfBQ+Wd+6s0qkR406XFG8J3IxtpeSzBKZFgl8nxGkU+aRoV1
S6immfgnvSZzIVo5UcNlStrdI1jNlomcGEnLy+kMzChVn0JqUj8UByMc1fpdeU7F
Nue8x1xzg4m782eWIQFeBoPfcjCNo55dMxX0bimwfoNt0yfQqCh+UASGQUiGkTVv
LjqLt/Ul5qoQr021ZYsTxLy1lKxQZnbDcSUABX7pdJIqRSw3LjSIU0wRhUEiRl0Z
J4tTCWH5FWchBxkW26z9PIOjjK/pEhk1XTSjdOdQLfclqdP5l+CtOTthq5WRh/K8
cKrfWaGKpg9E4u8L1xOLDUbsXlMvckkZrSatUOPPQ9L63E5u89Kb/kYatuJxNuY8
6veyGEOmY3wRBEHUzFhuoDGfs9RfyCmRTqxYophCW6PEdfYr0JzpzWuvsCnT48pz
SYzj8pd8Qk8bt4cLlzpbsGIo9846Bj1B1DaUsnTC9fpW5HCbkaDqLKK96wiObdSg
F1WityeXglKBCKzzoZ7mjCr9sR4Xs1HQgWQLkLRmxnfWBA4K2vwjTSezJxIZ8pHU
yLjuOf8gePUVUdRU7ADo+yNoI2Rtg66VFeCNhSzxurCIGorLJMo4pG7ap1h/Ysri
kIlN/C1gIsvePcvKj1L4NxuHfX9ulMMVZAyp+EbqJzipZDAGy6SltNgSDVEuGuVk
DQhI6h1tXD7w3KSkCHigw+NneXFsUA1KmlVWwbyQ/W67RFUDGJb7uKCEgjtqqCed
sPAZhVPpQ5O9teMdQ9D1sQeJJBywSJj2y6E+eMddAAJW9eCaw2ZZPxSgFAj4ob6p
rcubE3N8/d5rBSuZZwgvkr/AIrcACQZqMzYaTyHHKPG9OMpZ7uerarIDXD3TAydz
0qHvhdBx2f97+y8voAPWnQ0h/ppco8ykWAwsCblzfkj7HqewT9EDl+bJOiEip18l
22yVrGPOFq/HML9H2Cnygbv+aMiJW6Slqn1vPRBOrQ03fvKwxgLfZC4aoMeo8By7
0lrb29UlqaDdio/WVgblH4XlWN1zFhlPcP9n7hy4W+7sRrt+bDJcF1ArXne8Kc9U
RxOjFPw2iCx2dW/LUiDJo2BpDFj+h73KlCCOpaO7Y/sOs4EnwZehYSwqyAwBOGpy
iwYt0xnX9GV5bB/KDrToHUDuViiCzPW4EtgdiuC+dPQ9tgj5gfWXDzSa+MhlYdpz
3aEEhxvAXgrCtRvAtsl689v8l57sqeh6j06GZoQ/I0py3mP4esqzI/1YMy0tn5Pk
5U7QoqTguCXMCpoWrqnr++IbAayCASenVQ54ZtSCkwSneuze+VwVOtI9u//Pg5LW
ly4zHmeo4Qu3J8xkPwku7A5bP/lspUlNXHoDiSIu1B5+bcBJF0kBbERVlpXkMgyL
g2ZnIz2fECbtUxq4kuSnPfQJo6U8y7tqL7yH0tYdl0CgAlPfRdxKOdMxQie1L7kl
eQxEZWFsRx4DAHUInZPwvqMebHwC3/pKxaLbhth99L+z0spuKbRNWZ7CP0xdAA5j
z6xXnsVeEuE0L/1bBQnxRPDJP0Jr7KCYenqHvOb6JbUEQUWk5ivc+A7XDOoaU5+R
5CP8KAg4S561DTgdG0C+hcoAEEJJ6M+zD3SYLQIGyU9M45EbnhYGOqr8RMGv2063
MBFS5IqiNQfSnmgH/j8hGcOID9ybRlx4TTB6YaDKLXMaVBCM4vfljkAFH7q9Y2dn
AiQAHE/d+BRYqCt9Tlz681+Hf8jgXn/58LRWkDeBON0SEcAtESHRPGOvyZNXJ1W7
JI/rWHWqxic93Hrm2exx95Ofwo69OXlRKfv+3IWWOG/kmTbzIYtLf+8Y4F9gC7Yq
xM2JikgvCswzCN4EXb01ajGpOtjEc3wa8fF9UmHwwA+8/Z4TLMO8fErMKaKMFtua
m754mU5N22UJpNEn+mPfVuV7LcxmxWunFE9d89wdots9JoGIsBjVq0LtQEdQ/RgU
WuEQnX3oJJqsnLjTNdoUOHZvWy4zZkOsk7sbFuSR+96b4vx4tSoR0Rh4ZWIfkY6H
pL58SUU3I+1ViubSrXmKGGFZchmi0RoGfgJWpRddGJA8Dl96l5lKmBqn1iKzA0v5
Nk5oDWw46g1tTQ/0KrLrLSw0lKQkswldnP3bRFYnUrpTq4oIpRDYe+hl4jo9BD9/
g8hiyQ4sD6fcCsYLE+sMf9V2vKRbYWVnlvLXWQpsVpgoawv+59Z8e9IRvtIZF0gz
UNZACrIG6+hzMDh/VXaHkgm52nmnm92PMjKVbyGUfuY0+3rqP8VoHvFhnBod+yLp
ETBt7Kc7TaCPl9mhgNkJSb7JeSE2PiqPROH/jpD0xHQy3FdLTFdojh+fOb7LrJoH
pRdWkOax7SnL+hMKGlpZOi2X0INF9oIQQAYB3zRT8IxPPJyiPEOVIhJZHO5cuPJT
fykcyYPWulqEV5jawa0DjUs64VH/O66oRbSYbvyFEnWYIPz5GaRKUz0Zk9/VPWWk
w+A/T+2CmpTj7t6Q9BKciScGWS8/ie11//9D2BglrUATMMex0eIDiVXtwLwyKYrW
7FI9hQcRMQbYtqMo6STpHvIh8A6UZvD2TdEwjXD6aoLwMFprf28LxIVTddUDlGqy
zloroGw3wDGzxWIzohciKwsyJmOSv3iwlQo/uiagPZ1yQKCQkYwgc9GtlmFmNZk6
FlkpICfDJsferoGlpxPnb42dOg+WsgxSYoYjE7CRuyY/roUS0TCqju/mtswJJjT8
HoFziKETO3X7MQsjW46tlk/LzC6oIilheelfH1+YwpwiC7EJalxxgai6bh75fvjZ
rx+2UFSEeQBjhAgMbtGl9KEG3hWOtXJw3pHdCzThN6NKm0HQ8BYjRoGv51c3h/ab
3hQYW+YpHGGxRG2dsG76jJb3N2DfqxVclbS9ZrFsL1hBiFEZPGFXU6HW4C2WFnXu
YEtcFWKsTJjm6LTnNTA2xGz/+jh6Iy8ZPBIWng+TcP6j1U6ibJ01CvokAzX3Av6j
lBinE9yDW4Uj2dAO7G+P8c0Qg8aimBfjdxovWaljhbgi6AUu1EXJSoTD2IZF5BZd
rPNtAPE9O/5vlNAOlOO1Wxt6UgrkThohuwppHNSFVSuhXhJqgYAixqmPkxegrYgQ
Xl1b8DYVpLHJbha4ROLXonp3RFEaF1lWq9dYeT3sBjDp+3hJWGWb7+Txg9BEbJeU
xHmZ+XIQTXu8XEbNxzz7KQ8pwJvtPAmnaD8qaVV1m16KjLElmUdobrhAt1sP1mX8
sf7czFlaL/8LDvuqQ8hPDKtHlRW99d8ll6nA/wTdNalDsINwnBBmPqky1Y8IfgZ8
orb6z71T5UoHAhkEQmBJ9D1ciiiVF/ux8mFIGayUf4IO8EdpSvCg2dyzPTU1/sfW
ZzwONZgcL8y2UfCzmt0rXNYp0LsVvp2EvAd2jMdrqKkoIpkVUVgmfsTlOVks5kD7
xC5amcHfggTVii1azWlabvRv69MyRYJVtwph57Ylf2uwIygVYki6UUDJVHDI1ZUm
FTguxE9mXOPdH21bINkuOdqAvbc0CWHIty7HyiQRD7ytkNDfehH+PLcZv68Dkkji
CqpZiddvMo2HkD5yeVOGqrjY6feEaCVRsqbUcGsfcVWSJBZOP1VObDHXVWv45PlU
6O5tvtDhhwwT/Haqqbaecu3dyn5HWhWiBwPzTRGb5+c+nVZQF04WiPm0t4yvGj3k
PZKOPYdI2daMcRx3jpPx44+eQkCGYZuVsOIPm9zHWr0/U8Y6tese8ARgw0lRSVpw
Lex3AOB1+0m/4p7Behw5k3lurBORRXNtrV6/GarYTcBuEInauPpo0W0JERLsIZZ3
Xb8HJ230Yeq7DVIkxPOqd+8RkWjRxjyeO9JbOcUBrExbUFA9sVg820XxWWxBaESK
IDuArs6wRaRXJigBSoVYIJ7NXWpM2+O84ecUfhEmCWY4sV0jI2BK/gK9d4ttFmb/
WfCkc0m2ranMfPO+FnOFX3vNIAWUA5Kuxor0NTZJdATnXoAIwljrZ3ZYQha1IWoy
iejXeNdUVe0a8cm6pZpZfZqptGaFKWgRl1B8CHhFz8JDYxKMiSOXiAn7ckg2x6zG
LZSkEy8QvdSX3PGZtQWDRalhKQRCCRGGu2PxGolA2CaXYDhhwpefP5rdozrHVQzp
4/kHx6r4ojo5cxNUF9DfspauPPAJXMLiqfFQSR7YI6u/kOowmsNwbIdGFXG3J/vg
bLpdd1VWcmXEkvbUiFXdSxZR1NLVytp9tBWoq89zx29PXn/FHScqr5yiel5tiaSG
wuncswvBb+TE3A7ID2ykIUlOlc78kuCOfm/KR5La9QhC12SlL2cNBVvQXd9soR5R
WTPRMEDN//QactyqAE/02rRvmlfNTophuihfgTW4M4QXH/4tf72d+ZfGoHhGlHzc
IxvYxRxPtTsJ59Vxi8TK5Flt7r2O1erjWThdS4H3IaLl+CEzS/QjpnzCCipdfG45
WJKBi75m6o2GMPNXfn6K3kdCgyo1ViwFoojZKaQJmAsLiYs8XjD92gD5hAi2acRd
jGrRx4A2eMdmGMZpLC4bpXAjWsWYGJparBEyiDIUyk8HMhq78qPc9RC84fyTENcQ
X9wmVe7MCWRcwrT9glGYBCYuFNz4AG3hK7hodQdDLl8xr0baZjUkCzKwZemfq48L
thjgVzhJYfN8WHS21TywxyxnHNmFFIuRPZ3DRm82vcah646jlwrV0VjkCJHLSUSH
IYjmwJ7v5jfu99Cm2T2kHz28Es9Ipxvvfc5lotxYcY6eGtOnCBPv7y2QIV8ISB5k
0zOw3dvCeHzS0ECd0IAJLoiEom45exOaxZBCwpW298EnuRJaNvb7yGFPlMYY6CuM
+dDPo10xma91njqNB1ij1Np5p+FXOEyT9qDSrM67HBKDCZ9TIyYUNUCW57E5RjXp
Ssti7MBMzYJH53k3oTbNLviDOAAR/VDuEBorKSlg4Xs0675Zo/C8Kjfy5V1LTjmm
LzUqcn3Vy85g9DMRoHcPRPq5AUBsZrl553YRzBpB7pIeo/zJuC1zwkYGfzG1Wvk0
gLPsHJLKMKt7j1/RUODXuRR0Kyx389O21T1lbsPYcQf2lPgBETj0zMk1b2xIXJX5
kwGl6VYwyRzpqB6RvmLrubnaXvoNm3EBG5fGI6GsCqY5yRm/VMk8vxNeHM8g9JLB
2xEePQz/CvalKoiWF2M1qmeKEB+wNcUirfYJtTwUCbubSPDpHE5DcyPUyqFaMOzJ
3XU2QYpqkLVMM7tfFdE/ka84m2fJ08eaAgOGvqYfKooA7UdEj0Y6oPvzLTg4XgLs
9BZuSTEoObW9MWFQ51SpYm/k56IERJLMRNiZ0JYEMqf+1KppMMyReXrBkWdz4vyR
9EHRzHNG/5mHbzuoA+b7ydlV2D5lQGl7C1Pr3POWdqNF4XB4XnStvyuaZEvV0WKS
AK1bc7FjPM46xD9ITdEy1V+BovUqhTE/n0lLGnqLqAY/LRcUbWiUqjQIwU+/0HLH
NrZb4s3aWjqwJ1drZGude5ldtFcpvvibI/c2zQPaOoNjoiBp8eHdv7gcW7ztIzzU
XQCEZQ4MtFZh6yRq/0zRbZ+GPQ0jr8qop1wQGSRTdAFCpARzGMlzdrGI2Ce7Uz7X
f4wkzmZcA2qG2OSXWMNR++JQjxbVTuA1YcBsn5yHRBMZnAbmx6BkhoDSGOwoZK1A
cmPNHM//Dv3TtFCd/01jKeIuIC6dn6FOqB5ZHToW7wGBG10Ya4/dxY2UXN2jdNap
GP62OewXBZkkslpi3tb7zDSCf6botjRCWkwSNnomFZJJLWnvKcI/urjLMNBQr3b1
eBrsLaGQJ6phpygHiJfc9Ia5BE4sqbiApkQYgh8MiWmaVaG3YXK786mVAhw/83q3
FxsAyDDl5+Zg/PP3pW6cqNWgjJidsr13d5vPPmKxq3l6/dFD/P1FQCzPincyVHZ4
edYYV+qIzSpVi5RY/qwP0gF44g+TDsVhD0HRxdNKgaX4i5npDWsfZl8as+ulc/T/
sXJQDGGr1J0oe8AvLzggfAUN0NV2mIq9zw2Sl6j5OR7W4cHVelsYLsdM6qq2VI9H
Uoa8QJd9tktkcCqn0HpLeKSadD5A7tpBwMvRsFSzkdRu0aDzKeMrqQpiMU70AKus
2Stey3pvskxmRYYJgC84N9bGlPtlwiiPEQbkJ8pWqFCjFwVxnwR6WjFkq8iXnWSh
IDz06U9NJTCVEslhYKAblJ6I8+B1udFifEasRl2/gMCy0mtHQZ+yZzfV8M9fFhoW
4bUdnJVDSm+KUPpUMgPpXAhCfnCICfWIHOYXJwMhW1vwdpt3qDyw3NTUNAQI9tsb
iarZzARRJoo5CuYY/3NZ+wG+Ac1aR4e91HbYul+tox+vcFBk3HIJLAVgQT3wXbAE
RYektCJKZwT4mtsHmRkH54HiFMHE+VA54nqyLVxhB0w8PzkWK1NINs1hSBgurwtk
8WrsGTxY8DhEOgifL/OmLyV842n4AUSsCk/2u9b0/qtsZ2qQ3LgMmc7YbHof9zMC
SSlRn8mrZBKkKKIf8g2jNbocK7TpOIgnj+zlfDEvj5c4ChKNL1iiUu6+LeWkJnB5
FNbViPUWh/kyozia7LlyJhZaG/KaXYob+La8/rHGXzVPfob5klJRWc9uAewPblso
7q/csRORzEC/hFWeFkdjhHlv1matz02zyJDNgFc0PpiaORbPtP/2GRdmZAQH3yYv
2zFhg+3TzUibBRep0lP8T44OgzR3vQl1mHFPcBiwD/jXWxzZs4UT6SchCmWifUGp
MNByxHmWHE2muTiFucCsSaMuupozoE4k5w/X3z5UAjxZQlU9/vOsLNGvvF2GMP6+
VtzWClK+87irhMXtAuzpzPrk0gv3NL/jsCfEubZrkbn70Q0kvekFfCp10mb6IoKj
I4gtJCHbkx6N/9efCzCZYD74fqRqAhEhodk7ewZdxltnI/kOBVawzCPr1pFiN0dB
afZV1XoUPFHUog6EbFkxRJxXaJKqbU4XgLrODfHfB4b0UYg7VGiDC7rM62Nr3qqF
tsO05YKEXmahs39ISCTmVEQjhNbpoT4j4w5xerQTV/5Y6eK2NJ9O8hq3UhfkBWJ/
YfTGa0OsKWHa20Q+ac+wDvia+EiDvRj2rYHOzoc3/W14Zjl3CggmnnGVqWOpwL0M
T+/uCd8fxzWiccdJcomXPJwAFozAKz9Ynr29K03dthXUjYsLexaGB3IIWllL09a3
iHSfknQ5eUiSIHrgc1Z98t2y6iSYyhthgnNZ56KDVnFsm82C7X93zM1x7A2CB84j
ecZrf3emDhrWO7zGmc9S1qVhb1RDfkZU9EJMrfVsijNEhTFEh6XZF4oNyYi3Dm/B
JIwvZUjVE1k4U3dtyuBDmDxQhhbE5gQfN7P1pLRrqJHC7q9N0Z95xJohxfhepWo8
eRF9tpvikvdnW2j/wejj5FpbqSfjnWINCcktM1ewr4HP9xFCu1Jfu5pD/5RusyyG
ggtTPZgD5pNhUGnU/LdWTjKWDhPOdjNF2KBE02SST/Gm1EkKoFBNblKH/Trmenv7
mznQkn57GDFswb8qpULzEBefVmGAeeBer+OdPHrD7redpRSGC8Yrt0HocvNPHDiN
KL75SSD6VTcKeYTus63Cto2RoJyBExdrdtIapG7wGAKspEt2TNkyD0srqkGTb50t
qG2nrjL2fWuJrxkGiaDEqK+/pEQ/O4OFPEuuRVqdtWx8u6YZVX63YPIPNEw+aEf3
AtFyjh15/58IWPArEiJbg1STK2YXHSn1oXGgfdvwgiPImaED9mnXsV6wuaq37IYA
QmdLkuCL9ZhQYQduMRkSv7G0m6tK4V5Vv4IcTYXAfwbzH7DA+T2LHt50Dose8hnx
9uHtN66FErUtFYZcjLw5wqAWGN127n915jcyxeJUFagUkO0mox2HlGNH4nKfiRwy
Eiww4Sypb2IAB3o5C8TRJQbU319c/RopsTnkS7Zjb2TJi8aA97CFDgZc4WxvaD7Z
y+PikXp88cIj98pjGJfRfMlYLOOyP/ngx7Z6dvHZ5iKgQU3AIlSWDy4S+AjHsB7G
6UovT4APu3yFTzBy+m/rkiv78FUX/qgFShALg8i5RyFXjHBpgfIipUZhrYA3Ei/U
NhH+cLhaT19zOgamXoJgZmLchiDe7nGLHc8peGb6lerikpAhYavS/fR2QANkoh7S
4WF7ZPyY1xRwIk+YuzSg9yPNdFljpDX/DOvgBEUbuHbhArjLbInQy1q7whY3b9Mp
WfpkCDtBLcNzFmZB4JMKpVdLmjNLVBdCXG4SzG0CdGSFH5rvY9PTBW2Xfi4GPF7c
rtkmTV1Oyn2a9IdNWKYGYuFYLmoW46Pv1DnYmqKDtdKqWhe7Tvh8AQkl8OYttcFX
4A7YZ2SJX9dkmn//opofljke92s8Hn25zrNxO1kW+0A5XL273rYzwnAmKoqgQ86w
wsVrFlDr3O5DmNRc8nY+b3CQugQ1rXJeJvR9E87xHxANDvHoM34ttgNDvkJErElS
u70IEXSSkQYf/yp5SBBF8dmVmCpCRDQq7Eb+43O7Lkni6CWzisEJryP8KWnt/Pi2
F3e5W9vVf1mRBgPT14inOr8UKpddYFqA19gT8BlrzwQVa5uLtzqlAbtSbfpaLdO7
oxpLiFPtoXtzGVRNhxu6qOwiM5wQEkF+9yXxj6YTSMLvH8UM2xw7OMkB1iH+qm6c
6mdwLNd38Z9P6steo/ovz1KKP9zVhTGWEVt95xuUvFaYzD0kqYjGiR35R836wT+Q
Qr4whxRxmL1u9PV30tiCatGDY7TPo0Aiej373yxQXVb7MDRz/TdN81XRpHwg0AiL
z7opM6vQCSmkSezXQKcBwP0zixK322cg81e3acQPga+Jj44PzxPLjbbqw3R5bqAR
snI2BbAC8lUr59ltHtXutuGt4N569vpKMrNroxXhVhB+4d2lkib0urgdj8XPnmYB
LAQ4PyxPaWMQNpaONv7C+UrZWhV6tpQUyFnts6BvP/YSygzcog0oORDClWMxfuut
Ry/vtD8L1PspairWDOYPOdy+bmZe3glkldO7OS7kj6E6NNwN8SoSVxvHbRXArFTJ
KFinUapXtHrglq9Z//tVtoNJgBri9z4kBaHEjHKGanzPQTMD3tVlxIcDCrfLa2kK
toOSAWjFTZSxo+ivhEv2aHZzmj0Au+CvAkXNd0YBmph7U4b7QQxYMbDRgfyoqve3
BQZI5dg9dRYo1bp3/6CaNE0VceHdhYRrqWiAAx/WQKNMeX/Bhn8r6ySqkv4qZruX
mc5R0ZnfGYHfkUbbpvvXWS5FFpgfpocZZ1tH2yKoBCshjldxQ5uxSw7SxV5P/vAY
OhrtcSkbPftK/fGWEV3ZxylFbP+2ewNpeqaLgs7lgfgxJmRnD3oHhuPemhetYUQG
oarIDzTU+13m0n76jlMlP/UWxVWcWR6oJ9N8w5P7TFsm3sR6U6HqMZ/4w31rX/qw
imjZ2RerbLK6c0atvzjBFg2/nSV4aQt4Bu8JmAvqocPNXtPP9taMvQuctY+nsXcd
Wv73sQWb8SyAGXIp4XCnPveNZBPt1IMCZADP9R6qSxr42tKHeCU/5AKnOQsVU5je
1dJmbXk367A1WvR4TaSSdC3ABjG71DlqT4Oagmy1hCCf/DrPwm6PRlOwHW+YEs9m
HOsg+8/PeX+6CDaIJzCw6FBTKWQQxtli7TB7QjAax7mgwc5EbcW/PaBS/5mTWchK
vVgLy95mQvNAYEQ8gbiY6AVoVzVGofLFp3ziUlZ2YfyiJClGh3Iry/Bl353y1gln
NAgIwz58tQoSfqSS50s9ujRcv0YH8WiPc0whO4tL7JRXBtAqbHxLoVo8ZcGYgzAL
s802t36d/N6Gb+TMsyPFfYv4kLXDiHmaxZf1c/1TsCYgPexWruM254pw26Hzygwy
tQ9XvL/QVabzeaibFctNqqCWrKU5tTkCrTPONWIUZNeuTY/9ega24Cb0WIPPzhAC
qrS+k+qgHdhb8Pv1zIWguwghGagQKl82Xy6NCpK1gstXAoB7H4hAJN6JWfo8meaP
XbcAf3KBcUMIC1kF7+chPxFHaNqlIk+poXKwRGUNX+qW5GToH/ksC9ahIAS71TVz
HdSGOcFWTdP8stX1f4Pg84ZeYhBBxFQ40TH3wrpx9LvJmPnB2Opdo22Bqr+nzcbk
a576EGUMRdKq0jzU1ukxnwG0ZBzx7YSQoZKbdSfhZsOIiPOZ8PAbMeKnGAUKZ544
fedTfNLNaO+U3IaHiniprTMqzzzDM8oPw89GhNqW9oq/OBHF4lTW6DEtyixMUfRx
VGXxePmXXUH2n3U0KRw8a706KJKfnFPLgRa5ENoJTAJyQXBixri744ttrER7fbgY
QVRISg6u+eC3BBvDtMmSE2Azy6JcFlym+Nn1O2K7VAazD3iYlqg61iNz9FSlF9iq
EusowS2BgffQDFC2nbMRk2/9hOK0mTDOc5Ra6Fs7jQyr4uE4UGRT6ySFWw6vfhxx
ppDwi1Daz/JWlLo0KPXfHrxSUZ7ynVeaZ4pGettV+35+fkgprZbXxpxOllqUDY6c
L9rGHAb2nmq1v9m10cAt8cqbRWARObxCBR3Kb0Bl/+6A7OCsjr+zcjF0vjMewJZh
R8RTBdw4H4Z/PmI/wml42P//31pshk6iTzErqdRPahQ63lKV2gviE1WpFNb+zVd2
3rscLaFJJ8N/MGL2pCVxA2NXZ9S8v/HTJy0mqnTdAd7rvu/n7PGY/Y3eHPkQh68N
8ZFRmLiNt5zswssfH3qe1a/NG9ZJQxILvirTylQG31CAt4KueMWFQ+cAJIL5EL/8
vF/UYk0SX/xKktj+s30E2xEKa92e/HQyj1rrexTWzkdSfXvfQETp9Z7CPCt0wFsp
3KbgnfkprNGU2QwnaPqtXALZNZOsdxTomkzcqpMbQUch/S53piN9Yd0PVUb1v2Uz
Rb92dwogMm/vnFCv+6z4iLi0ROCe15NEu6C1JmJWEP4BK3KlGPLMN0QtlBZxBp+r
bN1U0VJdUJk5vHX0BAuKMRnpx872HKhd7b0poAnjdkiQEJi3eoPTXcasImRZugc7
kLlUKEar5kWwfhBOmk1kZtEXZgelBQxLZYogYyQMIm7P4QA6XBesZU4W30hmTUWv
xkomDwjLYVNXWIR/F6FVH1DyMUH6OON47/ca8WcXDhm6hZA3d0Y35PQuFVdrnDQ0
pHceoLpn6bt+0bk/3iipLDxWgXZifgiAbcIBlQWKJHP0J7LlJy7HriBUcAFeM+q7
hkMgWyqTZLRcA68J4WgdvYRzETHw5c94MXUM2stnbt1K1KLI8A4oYyuQbrcxuKGr
F4z+/CviwS1MJpVIritpxKLDUzn/5X92Ntk7TsT5F0kcXtAMHsRnT7j6YGr97pgV
ThwaDoWfJTmdQ5VwehZQplS6Z+2g9oVGWclDITvWeuZPhex301scJzuBjKgWo8PE
L1ExVQl7hMH34Wt0I+ZsJFLp/Tm2i3sUHnsYEIqbYL2hDNfgFlA5e7BrS0zJYxuf
J2OkMskrfHM8GhU8TXk5Bm8M2rEy3ZrA59xo1YPLl6TysbRu3+rMrkFBE/mkxwwk
mSDuM9dM0FvSEbYN0aK54O/No1OdHk4tGUaSLu3P/KIBrWpOUwuSOfoBCr5Dg0hy
5FeQW0rriv7y3JNLeyRDd08GaY5DW7fnOZulD9b+PsK9OXymCMEZMB19JAynbaUU
S3I/Z9JNgR0y3ocFV5SSVCV1kugM2zKvE+kqxVcFVgFMA9bVcSc3zzJK0ituVr5/
mam9skcsLZLdvpuHqQsUw+b/1/SxoL3J3C4QAqcxnbZoR8bvNt5DIrGfG9MjbJMa
TocKHYLEZjvUJNtDZEu49hQWluLDgBc72oHWEvuDotlSz8vUreqEUZiCvHwCevj5
ZrHytRWBZbFQ1dDSRtcmEj60FEK869S23/4nbKqhJ8YwjQopxBBNQeGTeXhgY+QE
wTC/ua9SbnJQa99GrrnKFtgqpkCb4RhisA15sbqHqgbJTKEj6pnjVFmYwfze57er
wfNOcXtlhF5YGPQZ+b/HPAktf/eykruEs5cuvjqTai/lOMXtW69nF8012J1FerGL
EGUdGYTIpENNxAc5JG9hJJI7BQksV3D4wqgjTmmD7featbCmswYqLh1/8GkrF7WZ
715oo2c54+lvdm0xT5DoVH1xBufW3IZGAaqSEu4Qg4gHjb62M8KiMiLjSaB8Rx+z
7q+Rm8oSdYytfj/DmRfB63Zrbcz9zvaqo/4DqFyIIabd3TDucDZtQdDlBdLVU1ks
xXoHEEC2gh0wAx5G/XW5Ij6e5wWzK8lyt6FvlDbUI4/8IPqTY5YGHqBluVZxonQA
h9y5kTLL86xIEdPNSBwzTEBjdXQkZMEM+CeOsuSr6YNUT1zXal+vCUjNedZJs1AF
jUAyxQHY4o0AInx9cB81IPTnE7XPypyokcXsAp5AUd/IomZZdDZZoxLfsnv4th0+
h0h7RRZGMvM6UqSaFuduLz2XwTzFtKdsnCg/kJP2UOFRXHRLuu+eMaKZoBmQktL5
Bti00JLoedAaE1xMzNBevXShBBona32wr8mR7Ea/ndoylhwCoL0wkC7gheYf+RTn
WnM+vl0t0oB7pAOzeaf8yb345i5sAljkPNuPFHSWVd3A5RhLfl8vgHvUj84DrGKk
FBKBnVeyRmSKMwvYILeV04T3vTd7uhi7HAbWAVk3Nk26yG/MNxCH9ZratPOeuuG/
FF9gCmyDBEbSB6YAAFPgWTUNAdnizhMXmXzH0sWW3kn+psLWgayslg6OutrDyOXO
qJZ7CzHqxmHUfKXz+ej+XMQfBwUQc5nbFhcxLtpVSugi9F2hXZzbo12DfED+Ah6o
ehgkMjGE9RnvZDcO1VaOWcSAHpiTbRpkNvyCjaAZ5vhHMu47bDXlKvoFLyJ767CC
xNccm+mNbNAg+95jEYd8aj/euS/Gcs5cSuzFifybZCg1HUUS9tV72t+KZcbF0fpt
opYlRxxnrXqLSgpeYPAywGXpv7xl1IKOiq13ki09y783lxugYD7fsbYEChC0nFEv
YZkgfx0J7MXGaqiAeDVlFlpEgTjHdG713YUje00DVlQuC/+tsZsYPXbV/bf7Pk5n
wXvfGSqS8NUX7Ov2BTNhrCcBAIK8hPNeJFm4mXQgX7X4wlH6EvsZD4VBg+Zmgatv
PChTVSEx7IMqBSxHNSzm9I+AgUKGYZj7aIr3fCFz92EBvTskUkMOKkS7KmdQ7Ybb
/HvbSC27aF4bMiN0B/U1T2H1FJ6RAsjt/VUS8LxQzHNyQjOlU4y+5IPHlQaOmFZc
WJgpoLKI74TcPnzKwI3/6QTRj58nARqvat600SG4ol7erXIiGR0rIY2XQ2LGCMY4
HPLb77h6XbrzZyI5l285YsXg3iL03WExd7kPy0pdWGGpDnVfI3JdmANHkZfINg3z
NGsg7/6OFnBd71u6uSdQuoLNs7TgSFSphu1GIrjcLinYmJVb0uIP43hBgFMD/WKw
JbsVRdZ23pgL/GvL1hDu7TklQHhyU/nQAsDZouO75VRPGMG8HQrvDHbtPUvMhAok
3SKKAnLfozb+ABsuMEUpqLVIn7+N50fvgaaEOHZoJ34EQ05FhBwuTMCGtZHhEfMm
lG66xMk/62e2t3cljeFVpydepkX8M3o3yfH7UXS6UNc5risFpafJiMhj0rRMn+9t
+NI83TXVxgxsSN1eoF3zGse0flxggn6QU58R7sIeZvpdjsCVJ0ShVU81jNNg1eaP
IwPZQBEOyB+NHKL9kBIoCrKCkCcdreqlihuVwoliCNiliv4tStFQuZ6k9inxzVXC
0kilt6vaExZoS85HOrGnGHCE/CwuIO5yUI9WMg9jleaMrjKM5l6MzJSGSBw9LJnS
Pkub9sJjgBCgjrKobVqysCu+S1TIdjtSBH6Gn/Wb9EsIieC+mDuWB4JoD8MM5PBY
2GILcaEydvNcLh0aBgWonnlL7pFw/0ZHw0Ss/hHMqh/yTRmfkHHvi/SwfMlgbI1l
OZqWLekv1Tff7QY1oWGeqIC5z7pfif1TuJqGE/cGZ+u04QvxByJF+OXLCWEGacTp
rZL5RbzQxUTEnr33/Hmm96NuxLjCCFx6RTT+TRyfJe2qR/IPrgjAt4WhsFV+AVGf
FyOkKQ28DzpRs8DSDiZJYMMyLta1Nyavbl68tayn0W5mgD/wPLYLaa108OlsACn3
jX/dSuwkA3I3yBmDUTWtGIF/B+QmtfqI8UXpytPhbY59FvPDCGJzzSSzvFO1vBl/
VtwSAWOA7UndIGqEmNkgMq/LjKiCVaUN1UtUMHH7rBDPKLEIOSLous0PSNTlrGH/
zYUzakceG65By4Cd5sUzXrk0J5ajiuzjT1mVabSLlYnRSES0hVaZk7IZNwehj1xP
X2NCS49BoQzz44PiKisfu51ZkJzhkJnub4YW/2qOHj1RANG1ww0x+dvyM50XC6RE
XUbDSA8V4gQu6j0QUhbKJFmSSeLpqVawyKDfP1/iC0Zkw8FOd/C1JMOdeitlqosG
glSn4SqcF6rnI0sBup14Xgc+JHfe4kA63p056NfHQqhbZdq8EGG6cx1PVLPhvR1L
ytF3htud0Y7o4gXTnTOr4BAeN8L30kDqrWFQ6lLOJIANhqDHmPrt1SKxbTrE/Lej
EHeIEKl8Ldsq0oLJazHusLwPi5+a49FVjOZ1cOzqlFhk+atsC/hYKx2Zq95PAWn2
QADNW9hOUn7ixlehO2Hc+q7qk25aSGFeer9bVJ+SCiOKSdA4lLIh7qE0O3vAL7at
yMgImvrWy1uLNdSHlW9foVwjQ7747AIn4YWvruzx7D7V64BQ9Pz1pbiRZEqbMxwc
ZZ+2Dkf8mR4U9j+v6e7TK5B8U+D3O3hFYLFnqJ7nnrEJi1yHacFX7ppQL8VCTelg
eOG0hKDAHurMBOCc7mYowDlpk5tOshzv47NHYF5I7lPG8V/gQeVs/xZNgTsFTZv7
ZzRZgUkgMT/sbJzTD4EAB+2lgLY+m4WqZyPpfw6nriRQy2+xzJNNaSHcnBVkrDiw
nE8R6qAzCLjITLuhygmyxJfxFaGnYos/w7ZDdj7IP1eax3PcsJ6wiLK0ZxR96ay1
4YC19227YV70qgn6FTc8kSCCN4+aS1hmRcUCPVhs7vs9yAiY+qlYPy9Glp5C81OZ
FReGCRCMAsCcu5pN+y9ju4RVbb90fHXfFEW1v0dRGj50B1KVuqqDElWtpVyU1gH9
QmdN9EYBVc4RsFa4mxtLpLS9exUwDatcudOhfgutEMUWcJWsEmZiDoj/o7BEQYGc
rGepJe4EVEXW1THQyUkk/0ASkHqtGkHC9tY5P4g4Xe/Qmm1X6QN+gyCUzHWKp//R
strWo2zM0Oqlh4yYkfgw+h7BnLy0PNVOgx6vadNlrzAId6p+OMmgXqSzY6upqSUn
3tnr8L+mOFo3MxYoaOdwXdZwl7Yp77hpgEzgYFffE2Qq6S8pnKccukxvC/p52loh
4gtQbYWWBUPV/qNf1xbtIo3HYOVj8K2bsbsan3A1cJuu6vSarCQKWxBBbxOaY8/3
TBYoe4j+OaYO03EnUfZkKERO57HX2sujXr1n/PRtodluRH0H0E3WmHeWlDUteP6K
dUllBjpMqinrO83SNReBvFdU9kOApoolvB5FE7hCHC7zlvcl8fvKENzFtOy8Q/LC
f6nYrGOoXJ2ZPaNYS+uPqzpQF0eAVWqFFf0gRFrD3LEAB2bqflcwXj6cYVvF8v5p
lUmmP4LNocczhvZ3X5Rbe2nXC20Xi+ZoM9zw5H60bWFYUQmla1bOnlqe+QoYVylt
QymubBeETcpsP0MgIPzft0FYapHOl17N6am+egb3TSXqep0vJTK3sJtNzcszUjTe
JpiMZ5d/H+FdvnwSXzcyYAw8MnVcvC8qLgxIBBpDkq5/fuTf6KzFWyCOUZlmEOZz
j/VdDGOUcH9leFyi1WAFO6ZNFJgSvU5SHmFfwBDumP94Tu/4PIvZZUFk2Fxb5zUv
DBk1+KZaI+Bxj8iIMbL/ldFTrclpdj4ivFmwosy0gWC/f5039wNC04DURBLoA3HY
8Z1qX2Pdarq2vi93g4W08u03RuUplXwoVLN9Srr9IgRDmIhTm82nUUHcJbIKxziL
QlduP+AwaNPtzQwCK2un3U1E/Aej6gY4Rc+7P+zrQogsg/kOX8bIpyVAQSO9ZfSZ
MQtprwMLbmhAd4a+aI7gXQdi2DJoF6wsz7QfgpRgGoHTw7M/T4hSHEof9aRfKtJR
wpSyMkHMS/yBzWMjAIay/w81jGeF28JPtvfYZ2TDrC+7RbBAfcHh0SJu/aaMvusr
2YM5el3ZsB9QIiX34LbkHy9vm+G5S8QAtPamQ+fXUNZ7RSx2irHJy760V+CvU/t7
SldNxxX1d/ZfcRYdmvGC5QtK7zIn4YElYppdenylaKssPLC3+K/Z0ewZyq9R66cT
Xb1zMGlHUYDPj/AzNRKVa2TZwFTBXtgxYCkOFVWLN3KybTp41YohLrr7dDcZhQaG
RisUUlXwULV0GmNKWeAXW40Q5SaZ2cQ5ZyY4a/aum/Riwc3H/fTkn507B26L/2WZ
Dj7BcNe+lxQl4l9A9WKvHyqC54WpiaX675qRorS46WhVFji8rJIDYPYd08qb6aLx
nE8Xar5tzyBCQIBFHFuqID7H/WVInt4m3mfQu8voIFN78tgN6oeLEqGPKbIgTmW4
Tmli0VcHuR/VNsJVu/d3o4QVP0XHqRP0uWH/qoIfTeHXFkoeJMJIYCxhTkXG2lC6
c0s3HiBCSoonNUweE/ZpEeMMT2MmLuqJiRj4+D7RWeeQ1WPtIF2TKnhIEqZL5zU5
ynl02uDWLWS9hiTMjhOyAycckVUY2eqFc2CDAgEetvhE7yAttN0dRO+mLkhBjRYS
BXWVtPRRPSEc1om6tl8Q3H0yYwntuTuOepiJrcTzXWXNxsA9yzhsOp93F4Lo5e0J
qW/bIRRzWt5vkQiLSApvF1s3ZZ/0y75wP0O17+vHZ/0EueI79W7DbcegLhvVDWr3
XOIiJjMTmvEvdHczyq1hSkZ7abdLY4XfoEPrGH6YZssgO+4mU4n/WRvq8o4Ddpr2
74IwimEvR0C8fD6QAYDk+2gojdj+sPhB9iyXj2yBn5M4puR9WRy1+Ms9q9vksZxS
NeyB3c0ifECvM9zaX+PLVKIuTDBkCl5bU78gjTChfpFUlpcxhLlUopcQPRESg3N+
NYAJJNRQeuy6457J7wk10sHbmPduvOUTOEk2vSN6GXaIZt93G7wUoKtmO1BNGO/7
DSo2n/S9GdzrqJuzKY/oEhzPfnxD1ruuGmTUMEf/lWGiObkB01qPKGdympbd7Tif
UdHTb00lYYKnx0fI5NHfh+mG0avZmWlO8HkL1jP723CmEhM7AuevFgfbqbWChe1T
teyNHhgd/TYTYfyCzl/qFgkIey3ekiq94E4O5MYZocKT//GwjQUlNM93NPZvEdd4
3VJpIOK5rZB6mrkZfMIue/PGZSMd+tTZo6aferWQQ0A+iWVeor+0QtyaIJnBHAho
FHoVfOSH34SO3jTIqLAW0Vbk2SatIdP3QFk3ik2P4ShpUdK+E8q86XU8MpWzjHtc
Uqd75X49xO4qRZeOHVL6NIzLgtHOuIzW5L4VRZ0zF5CtoImbHEaOoRQA435E135m
aVuA4oIMgLFuKyZW1JU3nEdQNNqkgJx5hD9zzC8iCzQP8vaAoorcyMDdrxSR4yBW
5U+bK603DjAlVybHS0gQn4oTPURMWLav9NtOtdMee7jKrzHHnInk8DvT5/CG3/my
UfxJ2HAl+3CWWa/26qPrBM89zfWhzXIhBQJGrhK0pPu+SzC1g1wcd3W1NzhhXUB6
xSu24bbluL01uXZOisHJiBLRjXBUhRTsT8LYjxgcJNu5Pe0wDO618cwYkI8ZGAFC
1fel+MtTDdhZW9jqtd8x6TOaxLdo6NysT+AtVHU9Aa7EZqKodgzqpPDGmiFRMYm8
tjqXXXQ7erng5i/bXmmEgcGI43njgqA/CEwsr1CtooL4F0d0hR7fWHsm82kaNcTP
YxsWHAywbsj9kgdP15ZsJY+cDFVJav9OZvjMkn05+n1BebNM/+5qSMXA/nj3aGzb
VYkqrS2f9xTeXsSbLuwlMGzPE5rn0eXDU31zcE/MytAhH0OAh4h+W0b/JIh/ZXRq
AMgNcMy3raMxjzxDFkjEg92v9oHBcdLustS3m69VjxXcwm8uUK8CLnYGI0y+wfuc
o7hhpSX46M6d5p8Of0vkbtnHgIH5rQ00qMkpXZ7EHnA3IU9qtlPIGkQDpOUO0Mxo
88sTzM1SOs1lwog17v9f/l4ELd/1Zdy6Vitg289VBBUZuv2XQsWGChHCgcsi+dJU
BSIxcxiXefMpkrIzZkwoZdq+BAmIQiDaTTQAmQvMKLZSFtM/kULAR2uRqFPCJ67E
CU7CWqJ4GZISuJ604EfNo/ycyZ95zbfAD7gGGd70QxFcIx72De5+iQOGZnzYrYU1
jbiJmyNhmK9CEJgSV355OjxrYeqOT2eaVUFyDEYHlPxhBSzMe8zkqb8ev+Yigh1Q
tWe7/qza1s7RigVkynM3SbhVuZ3C3EXHhqFmWBjICdUDfFX4yTASmsg0cRqMVZ/I
xQtjDTQlerQdFHh6CjYv9Up4PtqMJUPj0GJtOADJP81JI2CYwNg8A3H+2EG4c+0F
IHxpcQmeGcbHd8LAqhX3FtEJsJEB7pZXkSj7wZWhnKOOq62+CRBqPw3E14yF9Ckb
JVPnE79MUz8CSQr5TrdeX+Wv589ubIc+JI8ZVND2SAmbxCdlPl5ZkFtd4tpKnqzN
6UmmXg4dBllwZeUiVVxy/b27Kg2czJPQXjJYmcw5JUJQA0RuR1BxjKRold+jXunv
BPveb5XAjkQS/WFJoMeLjJ+gOHs29R1Oo2q0hN8J7vbbrgC6nFve8Y+8yqDT5N/s
j4L2M5KUXmP5Js4wnxC1Mfxu6+QttgsH/Qyx4d1Jco1TRvuiuT3hQQGlJw5wUqmr
lPGRUIbLYMnQwS5lrV3j6Q9qPN+WlidepDurlHxKby23RD6YIGAVSoSDIoNmA2SA
Eznqsv5tx1JkcT2yuPu7+2Rg4A2ZOrINJnaGjq02ldsv/r/DZ4dcvFsvq8dZ8aQq
2arCc0y+Q2eVXcYzznG9BH/FjOoxb1HooKnbN/cPjXxtWYTFXbuKQSYdMex2DF7O
qzy75F69ZHFqiaJAOZXsPLTkcZPUZ9GFPJKdmlvN960stpq7llV6wOqV59HxSc3k
Ao9spMSXgegk/8R3hjKiJVmafx1a7RokznwiN3nlE3rA6J0xNg3bhKtOjWS2syTu
LGhWIWD0JhYfBKK6yoVIsa5A2CSY0Kn6ThxaEVfrr+HWUY7UAwfQkKoRgNwqxJ09
KCGz8smFFS4DdIb2776KM2rGqRu3ocQpfyT95xwTor0AQHyM20qAXMxV9APK790c
TLIq7jIAbJ4LfJskBUSrqPA7FIfKvT4hOlJXBBXoVre8LoEZU21AHSslbquYK+hU
IK+x0bT6p3MEbXbJoEVbCVFFdltavvU0qg+iVJREQZr5svp1l70qLFb398t7wBgK
/YlGMFRhTFVWJQdv/hRiX+ce/y5vnmtrgGvcEUgE07qp7w7FK59N0w0FLrQmXIsb
xiUaWEumD0tidecPQ/zDFMILZM4ALfGWqXhblUh2qHeUYlCQB651qBu/cf9y/HiG
yOSkPcAdPhSnzEf0m4raGNuN0tqz0sfsVw9bA3halgKVwZKD3xEkcgbmXWZjTkfB
qAXjm7jcqN0c+7HIS29DDTmdatDb5xVHea5BuQERewneaERIpfjeHmtTkbXdFVx7
MnzRHiQidRkJsBAuCEImObOw1LCz6B4GbD/e6x5yirHIurfUCdhFc71l+AYsXdJ8
BNzAE/Ez9pjledCKRAGN8Sds2ROUoddFS/H0bXbwwo0WBHhWJ1jE411OZkyX7kXu
duXBvXJxHuI7Gi3j/pMgiWRmSy86n/eRw9FB/6+goRUBkObR7Z5O3bf+6aKISpXu
0HpGYbq/ST6VtvhyHCKgwsFUJdzGr8pjrN+UVfKxF9exOhuST/E+RNb6/gRz5YiA
mQRcJcWPy7QVG7r48UVVtCpRbQd5wAWxitVYaYYzU4c0TEESiREba4zZTnnl1bd3
7IXiRFFwDx+2Ycgn8MexFIwnhQorIxZF4FvDLNSSrNFSyUdMuYJHkYDU4FipfplG
+VUMQ6jv+ugGpFdb37Cgd7Hvn5UAG3TUSioXRT25/Ls5egbjsrei1uVMQyLLwL+K
VcbHNq/DqR4RhMZcsIQIdq5tWkIevmICEkgMBe8GRL7TBmqTIn8XY4Tm00nyy8Nt
FeljVtDtCeChC4vEu+mgVkPBJrjYQDfkPAGO7MUzYKb0lgyxPp8/omOOpj14B5ZA
Dvg33rrtRlYTBZI/9iSJ45klVHMO6Xmw4WzqqOcv7mk7VOYNCbbai8KQQx1DUZii
tYV0mHbNtsEVlCJhzNKWitH6qKKm7Thsb2E0zuyeMWmF/Kwqhyqfny2qA6reSAn0
DRNZ8yeNbk0i2qwBVU+QvvK/NOJoK0zhCl5Z/gwF7PuXnTWTNe4iUz4GtZ2X8R9X
cg/xZHSC72QQ0wjhwLydiWLS1l7V4vyUfb8EQUQbn8GnJyN+mkrmJZD55lQBv21B
VbxB5uC1ObS5rwHsMsk/tUhf++RYireQdHPpDQyMtL188YvyTSzyZstk+IJ09ZCF
RKF1BcVLQy/dSWN1RrQyQTcJTkymTYW/YPGFIfsbWseTH8g0mNvK6fiTAfnFomt2
I3wWO6nQKGxxverezpL1g5cWyRK6Rbmt3HJNsy0wtYG5Ge6ivrCze3NjD4RSlI0z
zkdwEbVvzMUCLjwHJmCF29nJYZMZoXjXeD1UI2zYuWAtmoOWXrmvRfuJTSWDsPIp
uswr6dtlA4JIYwlYIPlClAq3UZ+MWrRMyIw703DdPKKjQuQfxr5mRBjCjNoS8tSE
LObWJQjfpyPBfHvaTh6MJKq98mDVKOeZX5qWHTX/Jw7nB0KYwUPREdr2khMG1rhZ
TWViudXePIDLxoiO70TiBKKQKkG8AD9nqCCylsjGbF6rgCHfavtPKqg1ebxGsr4+
Go2KKkbZH7gQmQ4PDoC5XPmWx9IXIo2Mmpg3R06ShpQilMFQprkCC1yB7ioOWFsN
n7GvyClXGI4ilHzkm0uIrCoT45mJ0rrRomueg7YhxnPPS8vDoPzAqVzXmwFkiqMx
AEw9gFz8eFmHK1HnGxLIk1fDD7INS1D8PbzNCoboPyhFRTriBknfCL6JcOEMhWcq
DZXCE7eMS6ZPPebh21rlP23FypVzazbFtTOKAsWpKZXJBRkWTDsC2vjPVKQXtCPn
2zCuhR7LgFShpffbvy+JFt6qzf9Bcq8xcMWDinKz6f61Wichj4EhxXZGOI+FOGfg
2P3nIn/fWNoFOiCIQ9hjpYU5WaFQsGjoXafB2fEAiYTo7PVJJ9bcswHtmoq3JuHD
xygXEQ2gnDhpwSwv94cbcphlpJ41b3xC5qIp/1KP+gqFKh3vFMyWZdyoypDEINFJ
OduZ+BJeMab+JtJ/Tpfnu1/bhwq9wswLpHjfI0SHS84iQaz/DkyhXE9DkI5umhZh
d7ZkkDaPgBnKXyyPyHCja/4LMRivl0Lkidf14QEyHiwrb6/hkyrbLoDQDeaf4eB7
f8S2rfY1A/VGwSwfiByFTDMjoEGMGhNHqIgp9F60WjdhOB0H0BHBva3HiLr+SZRg
BF/VmfBnUrE4hn5Kn2z+v4iIj7nQj7/nZQDmqjzADw4AaxNsEFCBBd3qoJlJvGDP
4QVudYUCYCwUTHLqOX3wOPjcLdWGGJEBtZLqnuT0pa7R4URqXIyoAztBHqR5UhsE
8QWY8GSaxgNyxjk/LlNpIiBqJbJ25xmfq+WD5iYjxIEg4+xF5NTkkBeGXjrdvC5K
SOsG35Dndu1MMImxWHKmmXdPBUJRmjgUi7xGmqO7j2bwuL0e/W0wKSvAZwwr0/mh
vgEbQ6FRf9Cyj13uoyTEL3IK+pmGH1RK19+Ju43GyhOu2sNVBWEq0okaGpTgOuqH
pHfdxp4t+mk4Ad7pY+pxsc3ZFtxREzvmB1Em4b6YxpYGlU7siwblTc3Y5eQRjbLe
HQ8UMgxYAfE/WmUaprPyIeA2INy58Z+p1DvaaIr/IaZzDKzT1GlxuKMbXW05Dhqp
19aT1ml///+G39T1znBPg765vNYmWM5FVpgssqcLFI8y7ov6uhcPpaCeIa/s6Pli
8Oi/NNxR5sQhuH+0Oull6ZsU+j0YBEgBK4oOzJtQuhUzPF0uEJCxMlbAkWbgheDG
40nxPC9ifv72qFGm9Ja8zDSUpX2WndTabuvPlBgAT7EeNYAXOT/k1PANkxY5Ik1s
5m3+L8JNKjwRW1zd6SdMojJPp6aytav85ocazozVLhMod8urprM+Lf/u5ctgtS5F
Wia/XI+bmPdmq5BQ2c5XIiZWQi8brb2RE5RB7Mts753MMjZlp+ZM94nxzr7utO5A
2GyPgtmdh6qHAARdDca1s/W+RqgB3V6KKJAGjl882OBGhYCIFd1+UH0zsbirHEQf
+FxlYNqNa5LjS1oMrW5uUZQsq9kdUzSX6G2VPiUfNLrA2ObaIiUOUOq6/ICMlTV1
4ecD+vCRxc6iS+YE8hXcxZ9Nz+7AmcyxOaMSXKVvWv39nAwZ7m7LHbxnMWqzCowl
azLmNMk34H/z8MbnKc050zFMceHV/FkyfnLH+OvGOFBgB3j1yctGWJTLiM3nyf/X
rZqahbcDtxqXnDmfz9NQ3Tn4HUOGohTknhzaN0b6g52HPHMLWgcGdMqILzymeC6h
wEZakSbIiQLZ6rvgJHnm2QM/dy+Q47hA1W4R/d25TOHH3aeXmflsKouNrWqylsa2
XsBlGf2EobXdDY0L5KLncbtEuRlZ/h/z3YZuBpuOyEazSdXN2GKVD6Vfu01qh4Pb
+/MA9GjzSvLg7sJactG4BFoUp23l4wyqV+rHwIi6k67MSBxwzjZrJLQFF20q26KS
NHpv7uJto08rkm3jIY7qhrBNNSEfQaexT0E9yOy+a8kv5RDFSN/EyOqMGndWwbC8
4MNMB+UlLwRJIQ4U3CXGnSfgzj5+8zPrMzic3siIJY6PHyuVEVXxGNIBid8tyX32
dKqimxzhjpnfrAZq1feP5Rm/HjBz4tNFCWf/KrqD0iCYcTrbeq57f5LpSGEwiHgA
QL8Xa8Ag9wHxMQllVS/PBMtfQaoNFzp9SE78MB62CrmKFSjBDA2yuZKLLAAndntN
3xZ3SELiKCwEcNw1W/m2CYnNtrEVq8FrmDI9jmCsNZiqmxrLd1TR0hv9jgtygfeT
TMv4mGMXOg3kvJodiaWdEchSwJ9Lmla2psPcxSzzx84gcW4Nv5oMC19i612aNm6R
KKatyZtxf+wQmwuiJ5UKA6/ddzd43x1yilewM3z91qC0aWoM6mmUIyACgLnSS6Al
e6ssMh/uSnfXaK6r40uuWmlwU30zxUqSF19MtbaLYv1zjkZWFTrud/8sA6CDgdEt
CS4Sb/gzxnBo201rq5bwFjLC5AN9ZqAS7o9qeMyN9WTiygF797/l26Hqyl5PCmJ6
nSVAjBL2VdLPTOMqDCCEDMK/xmsstlrVeRtUWqjsm4wqD/SjOFSeS97TtmP92aUn
hoCZDDmwwi5s9soGIQCzoYRfbHXxz9jX6ldjvBnqbJesPJAKcQJ61gUaVg/M9W2E
6+q/VwG9mo87K9X7gpSVR0anXty7uvJxUhQ/hFRroZkI4R6zQdDw95tjRvVPaEUK
nzlpVkxtJHF8w8IamILNpsDdLJT+l1CiQv6Cbsb4lTQ/N8s/dSXOPsMv4aoUSkJw
beLQY0pIWSYbqcRJCJ/sUUzg+aRQOgPY23vTmTTLIDAjlsqxtIjstziS2ZunXV+L
Mdx6NoNvvu8YZLGFwRLgCSr7EZJEuvVvUijw8XkS/A4kegGb1GWYRp7KBvTA9p7A
SWg0iG62CpSm9jtXWFUWnS48IO/muV1b476jZEOVPeRxzOKZEuWH5wQfhuC3rUwm
Mfxubu+TTZFcHbEY8XblghJ9hT3UK2aufiRiZlYgNVdGwx1BePIeyMzo7a3yEF3r
uuFNPyTHWiEeMX4Vlm1cqXtdUn8ZZC4+LBlOLkr5Q3Rq0gFXzK9AxXj9mSFdbLki
bnf9Iy3MDqX9I6OFPm0RZonkjapq7W9ICHYXh/YyESj57PXTNx/9Rpd0WvhcNn42
xKQrjV9yI8wvYTxDHcjK9JgVYyXSySZ+Zoo294sm7mXAc3Ol7O7WOKArglm1W64f
t931ca50UyLEqNcbp52yH2HW74cgSxPadzWRVKFhS52utdRFZiNptQzUI+FBrGvX
duzxOYt6o6G+HLZsw74t/VDs4Ijz/qIBVB1+n6bSmZrEsFb+F9mCcoP2I0vt1aae
PZ9tvPfvnVKFN+MjaaCj60kc+WpGwFs/LYZOJU0Ms4B8zD7h0e+tr5MktyG+OSco
TPcTTdTOBKq4pgklrFX5PuT/dtBEICfNo152JViR2/GskOSYxRQUemrhX6eCshQz
JWyzzeI0OparoQb6MvqNteWThSGoLnICpFkyv9rUNaEv3qX4/CnLRs6DAAYpJFWV
xzxT7a9CEZn3m0zdIbA3jwX1iJIp34r++JlLl3F4zA7OI3nFhFu0CL6OEbblwoeW
bjwkbisBOofr6SMmevoeaiDkf8D/qwkW8tPH/ptLHtABMTpkkan3v3PEyRdtOYgx
RiTl3k8z/ONErMJUQQDIoJxELkXmwC4goBpSoRx3pCwBZVSfCgjKdJgVkn08AFT3
FvTtHQX7HG5RKyjUQxnac5x1wp1pM5iWzaS2ymUeBE4WUVTUFbwxzXCXngDfN/qW
JEfF4n7mulMmdtSCOFwrN1IhG6o076r4XIW++ZDUCLHuChsNNriwjP+zvk+pbcoz
NCgdhjAXhkHp6ISpS1ykVvG3KfaIMVMSfveDTYAURHqIXQkTa8YtRLrfzXd0WEbx
YDDxJhIlhnSsyfxHDXH/mAtVc6BvW1VKVp/dPEVGOdkNqE/M3M4gjpkPUmwTMJds
7TYWKoWbZd4aCZQJAuHNqhK1j6lz7iaeN14PAHJEB5IfvsYhuweVLYsEBO2LNJ4F
aTJA1rEkQt91msVYUt1tDf8irhYIpjXd2wuUaWJQnagBA6e5oz0BkgqIcTlEQknH
LmuzCW7Hvu9Srg1eI0x+lf/DreIFXRR0RWc8aIyK63/dZmrCmsLqj8PLvkjQHDeL
wQPBPdIk/hoeHJKyKAKVqknO0Eqz4g79aPkJCv5tfvmYzzYtdB6Ga8a974F0f8hY
5dS9e5+zxBuVJl15Sh3JR7SQwqBqj7QBZLhXrN6JFjCZ1Vt2XeD2iFeFTJ7XLCXS
bzvBOkUEt+9WOPdPABMjkakgecbFxPVmCQTkb++RN06VFvvmq0+uSKHXnO+NTUhc
R+lX15bfqJUvFCALnD7jECzoUm6Ecrp5QbESvyqFhW6KebF6+wlsBedCerdznXzi
3egoxgrURoJZcYV/SOrxp4uR1OOV67JyTawBgmH3Qxci25sCFfaDL1Z19IzVwk8q
AXiXp39u3sczf22mRC8xy6HDtFr/ojzGSTIOxT7OIgbgkTgpNhuxyUObKmHRwuWL
ljnFuh8+ZOtD3oeMM862Gs5FNOIkzDrXop3HkJGuvtXoQL9qRxNmc85aBW2SF/Pr
/LazzTaIoTApBkriFa6F0oHqlZhDTcwIuGiDFMFFBSQxk/rKKC8hcvNVW8957SCo
S2fsjvFGcuxOlZzbC29yKeinLGPHJjQtL2mBH8KxD9HVHFHF9DfEgCTSkyGEZuhn
TGO/B/NicGc4TwsHu3S1R6ZaSuSWABlBr/2uHOsNQtdBToeFUROzKE0wQH5Ypvo1
BZBn6S1OjNIlDYbHdX8+eskaDgcg6+eZBzkw9NgsGbL8Bxtjrn4pLCfdFUs+v/2H
g7ISz0gxpTeNQ2VO/I4za5QTUO7awYaqh9FmAfn5kCRKE2raBjvzaMCeFX9kPWDf
u4iAEUjbxIXliSk18745441FKBOg1xGVC2i+7E7HQr0xxJ1aeBYiJMc0plr7HvW2
DSfbq3kpD+Vwe5TNPKA6y0YRRPLTn2V/mKrqtF5aQcDwasjH68B2BBJ+c0yCc4zc
QVf4uUUY/VAgmd/l5atBTEPvMf5mKFVruO8YAF6jss0deCyG2QvCXX/OJZAtbvSM
pXi2eBbPuqY5c71kxBQaPL2bhTEfO8OiQLt/SJSbJaF8IEuV1ksi2r6zCC36eBz/
l2oO7Qq6j+rRssK2DRJrHbA9uRNEh+VNxb0xPLCAMLek4CuTZHgsuEHsfiMNrLMq
Otof5Xk5dgCmOSszpmOVd2D6qSR+uy4eM7P2cMxpv90lhsynZfXdsXKQxYlFb1nn
cBRS4dwE0cfMnl/nj8lUlcBGY/rzZH9GeM/iaFx3Uk+XekZZDUNsNwK82fJQn6s8
7zXBCTRq9sFoXvsJJ9V10bpoT+deYkoD+1phwf7uWXUjkBuV9PHms+GYPTbZifw0
n2rxNpltsBQM3cw6GA+/70k6lSHIfKq6Z6YYKCIFv0FAH4yMHqBMB3mdwYHSAe3I
fZavnzJF+guDxEBfv9ON41ctB3+uIx4bCBJWNMh49kTQrDarukJJhUrQGRRLHtjZ
lm8I3kMLgPr4AZ8qhn8rECLinbAFZxDw6wGDRBrCS2QWBwM76dkShSzYFX1xUukJ
Xq6byNRdmxi5XWYSofMRWR05G/nvR516PtbktWSL84UGrbPaBDZyFdLVXXpUIhWD
ZO8MTCd9Qfp4TkqShZ7dbA1JqOPOmGZfskBtEPXMOFWIs1tJZw5iMFbaq98xM3hQ
LpBIi61RRCZgFxMwq9Co+3kl58/P2MVLOx/HqVp/Mhl5KMgujPZF65cIn5SmRV/I
4XFMM06gc6/7H72Z8VJ36/kzOk8Mq7ucQ27mVarp1UZ7ScLd8F+il+hN0rqXCFb5
4MWv0HGgx0QpgaPuDZG2Ui3MgjRb4LgwDJdBmEhT8vKSEBmpgJ1iAzFbEcjiW5qH
OnRwBx2mqgAv4wmUMsD5d+A2aEuk+Ihn9S8JUHsZ/YTYu1MfhCrQjivtpxv3UN/f
E2J8atru6hOrGCfgm5pfw05SER1iMRs0hSX10vMnDMRFS/a0hlbFDMuKmsdwZtMC
07taim7OYxjN8Hay7x3EmqullGDDPOmE00sV/EYE2O5rsCQwRs/yTdYHAE3MzD6Z
0b5ubeICm9bYMJAAfsSH4WbUey2h7Rht0xBwMud1HQsbT+HrU11V1DjVxFKAi/Nz
xT0SOiC4kwgszKCyWWX/sDa7gCjeUF+lqU0nMgTNZZSz1V0MlUpyT3z37VIgfA5x
1viInaK27B5GRMffZHewjbUlcb7fmZy7a+De9UYsn03CiLZkJlAoMwZUXW1POPEC
S0jCmRpufsG6LZqNTXH2a0VS5GNQs/KbFu5uI7HhLsAXmZGMJr3WQWZ7LKyXob0l
wsq0g2qadzz2xO9sAb/Fj0ALNjNQ7RH8GofYt7J3bp7BBcPj3k+Pz3JWpvtLQI/l
E+d+Nlop57kzljDNbjBHFfFOXc7W2Q6EGGlcaJ9wGmUk0ca9s9QJrw2J04nbsEDG
8uoIL/Q4CRgEtkY44CFYb6eNSYAJ+7p925jbPQmqq6NeTfvBwhekcpFE18eMG/8u
DHAX3uvc9HhMF9wRadyRJeGYMwQfWpL3cKy9yfFGv6tfDwYZVqAniTuGTyem32DE
ZBdmAkyg/nN1+4JnEo552UCs7q60Sri1QxGDNZUjD9DyS0DODvsRcVMpTbtzIh4c
pP/pj82QwM7zRklJgBBwMILICEK9KZXtUZUzrLv6pZV1uK2cGD9fWF+4tJva8/8e
ty9RtmdbIwHp8EX6b18hCQHH3SKA4fyEI2eh/R915GPLO99OAamhSanoeDVrNpXV
+tXyTP1ukRdMvG2ZbSeHNyPb+114B821Z8NZ0upmuqvCkoglQUJG4aOs428ktl72
tHzTRdKxXr2tJrrIG1SmBw3Na/dTMysMpmeIO1fIHoHzlEQsDSexPJSRM1QpQMiA
+LAFjxcHVKMBY1E7D7feVDfFDu1PLMF6kPDkHgvQScahtBdXQJ0Ou0HtwIG0KMsL
qwt5PA7CQ6ngmKKCCi8YNqR9kmhX9WemQufevHEi6a3SyFKti+a0go8bzpQk8hdN
lepNUbB9fisowmJJMeluk6zOQQLgZZWf2EjoETl2CYvdNQr2SJtp4z9qfo9WgKD8
O4fr+zZtsnzT8apfRbeIh1V+PrcHDn24EHPf+AzYTOAJ0NGK6yXOtqWJUA6y6TkC
qBrvreYFXPJV1HVxNdSJY6ht5NPOwqgl32YyPaFJyElttvO0IW/vYAMnu/5bhCFg
pVk/zr5p5EFLozBgdNc8HQBil0VyAXStAyMQxkLzGy/dmo+/JHftbtuQl07aHlKz
0L7WfaUPUKNedXO9roaHvbbASQjo89CbunzAzTbZQdpbRUymltJH70q6SejKlwwX
GLKHpcBh+742ZF8aOO4vEcE0NsMVN1JL4GJ8Bv31OHjWm+ufMGGnHtQeH1SqaM5R
HzaGgLJk7FQR0gP9NwZN7KsNAfsvsRfrQ/jFrrk+/yk1wR/tvX/4QyC7AOHJSxN1
ETi5r2sM9q5i7d3dMKyfLW0+MP71ZvMDpgXmwZqmReqI9LT73T/VW0exV64hLSMA
iC8ZR4EKL9/guRPjNlYtTwS6V4a76De7oYGJ4DrO9yHteQofTZX4s1b89dERrVTh
EaTCw1NhBiY4JyRHswIMYxA0kxliwptz0wueelZg3DnepKuOEn3h8iSZQHs15oL1
vwRuHgshS/45JpoSJdgW+AuybneJwXz5OvxasPqdB7SZ0Sr4OFYQY6/Jz8hJ55yJ
LKDupycAQ1//yWUcOlH7f2PSsDLbYh//3gJDoXidF2qtQnhr/puBJ1MiHEhWMrxs
lV83CsPgN1bkf3i64HiT6nX/dx/Hmef67SqDoe5Pbw7O+Qfxk+69sJiun4h+e/Zj
oKDg8xwlN5/6Z5yutLPzyKftee5xIIL10n/6BI+Hut1QLISnaEraT5BhyymtMYl9
vJ5C1g8zUS9lia+XUY//x89aJULmBtreFElUtgZWykkkRODzdYtZwCVZqCRtyZSC
ZltcfcMXDqBDBCdseHebVuOrM/KG+pwC5xm3SAQ97ChKLmZHZ+GFC3vgErQFOCa7
b8KVi/RWb172kOJk8T1XeMMJQR0piUjolDJCHZrGLdrBeeFyWeKpnMTqachoHE+w
Nri1ijp+gu5cb0zLWsUxby9YB7kw1ZJnCBXRlBiCmb8joDg7Wf9HXYo99VKXz5GT
bT/DhFjQ4hS9ZtXYlXFfqOj0ijkQQjwXabjDlh9aA9n5KNyxQdrkIWOBg7ikgsZ6
JrsBj4JYQcmhWUDauA2Z6ahurzD+u6tMGi3n1100NV5c8VtZDsQT1vZ09GiOQuTf
t1rPsC5W+Ug5JpYtDUAg3Zf/kxjGEvjx7cmp4ndXh39G8ypWmScwXLjmzdr9e5Y3
73dM2F2W+9INcvvFzEUyrxhwQpL2v91ZrFxVNGhA62fFWzciK3dWxiHR7SYl5C3K
FFTqCDudRjo6qKd4GZ49b/NezfIxk5ApFPx2aWVudsuOOutefaO80DHBsYTqHMVj
pkiMeanP1OeXC/i0XNneWbMRmPQTMCJX/JWf0OaAGJyYp7JNBjM5kTRn936JrXuN
3iV7Ptf6B6v9OUS8Wis5cgb204n9M2jCehR12IlitmnCpuFJqM7o8x6j7ArlCU8t
LG3aqq9xWRq/9CFzcEFkDenc5yTSXLb9fuPoTVzRdTHCc0ESAALbzIg1tcwnCDXw
nWUnWBBKslqb7ucmzdLGNXERQ66CjShNOz5be/FUhUmm8vXJvwQBDtG1Oz1o8TDO
TnsPtP89LAvbZtVzaTE7EN3cdgWjlkFlT5JpuGanAzOlYp1W87N99H2eY91DejjV
XOrzbI7oCIqzKIJq2PXuOwKHrRe8GfdnRMddcOH7dFH1GSrVQLH9hJo+vQpXAMrg
R/K0NNvikP9Apbds+1J7Qgxd+zsDlnEuMZLTDH7cEz7BqK3n6YlzekRK2iuafX24
VzypOfasivKedzjROll76SNBao7v32ZCyxdnpmvoqdONHMTouqVtSDy77zZVExbD
5h+PfWswUQQln0m41/OX2IOBxdgSvEdOQxJj6C7m5c9/MG+lTL69+CwRsoFnfIHr
9qtzKr6nzzQjFMIrEdTMECLSU+dW0RkjX2T+FN+1kwFbUDBB/Y4MP6V5N4uwHcqE
PD7h+Ynwg/14ZZFQIGD1Ab94HIRbzkW3iLdt25e/xfBFJ7BaPNQkCg1nSgeKDQjY
/jft8gsVMHqtfpnoijx6X0+hFGiXPJa7brMfatofS0gBRayjYYzaMpEkCBR3mXDq
43LnjO1jfKyCliUyTPovrV3eV95e1rhX9uofOvOlHyA56hLaeFY8NEpD7Ek61/eO
0DpTgvOpWyUPXCdhN9Y55qrZu0NPe0qJ8hVPvI4Ym1Iw05ns5NJe78EPqAWyzjPa
eZ9PrHC6LEpRr/RqofIvPoD60OWSATjWdA3E5341pBvQK8DlK4+ZdpO7Q+y9xfS2
hdj/G1kqJLS/N0MgW5gQp7LNF0ouYM4Djg+Ls8I7wUBrhcirvNevBXWBjDsOy30e
Kuz4d3AOewPzrv1Dp9JI/l58ot+yaD7Rdv92Hz5Xh3ATz2wRMkWuadLZwen9ZTTi
So/ayexjyyypYGYtCGISgcSnW1mginPeljaUQbp3Xr4PM6g6D1qwZup8pyk66UNK
fnhTdgEiSqYLlYKuM1rwJt70IhtLW6qxe0NjaIwlQP36zL01jd1zDBOz7vzK/UEQ
elSIW9ZRttHNbfkYk+elVlX3CiXjZM1cCf7Q7O34+k1PTzgtjN5KHFbqaXPGOjYh
PkqfFQ83mAN6s5XyxKOhzeOc7t6p8LJh852ETXR9zoVKLhraSEj2qODNN1/oXiMi
HhXAfUrDfsr4FXmaMB6WquQrAHBrImUi/jOh6+EADy+GPqK4/rmsuC3tdzZot4Gd
/0lY1DeTuVWgMHQjN5t3N4zyuIe5g+fHZvCNcQjJLHTHtqsC6Cf62hA8mDL3TEzN
8WqP9TUu49CS+D+g7PEJRucOORAoxGHm71U8dOp/7erNpNeLQbCfuEJRI1bxJ53n
copvY0inkVGHC6vhkUO/Xz+ITSUIQvb7bY34N5fCYZvsAJ/yQ1VUFgLiOHjzR8p4
q5AbOgy9rC5YGHGPMdxmGAs6NLUYg47lTKnHbhZPjImduArrQS4KJgJ2EITm3nkw
Wb5MplZFt+KEIKvuQH7u7fkD8ORpuzD23mURFeTacI/P2ZSZ/Luwd7WrhK800+bW
doeL7ogrSDp98juiyhtPVTFHFXY4Dgfu8g9QRQ+pvofB2pasY5NzOVmq2mm1ByPe
SXBXtoKnGvieNpE2vCbXqzDwFMgwepY0Py5cncH6qVVZZAYmndSH39SL+rYlFc6v
Azz/4hl4wb1LIsj2dC5OWc57SZ0wikBCGXS60/eX496i/EiDjuyept29AgY2yScz
pBuHM/67Mx7DuxBKvfob+1FK1miI18+EGU5WW0q67Ub+tmbzd2TbL24jDGiEN+8k
BTS94D0NnSAbQ0ERkglm7K8iAdvD1BRe2D6bKpdVP7D76n0bJauKm6mYanErYSB5
h2y8LRl8WiDrizjMBc2COb+v1E1DcQVeslUuoZ3PT5oPfGQ744pVeLJUbUmrnHP1
hdHFpqRrJgV9ipoyR1KL7EuWFtRXqKNg7zVQ43a46G4A97bpAzjpglM4XYOMZFLs
H1u0S6rv6d52txdU/KcSdxcLgQzDYKBTuZeABEwWtr1ljH3RJy4RWciKqzC29mhY
lZiKp/AifZXJHvSOBk73LjIAIQdtqCFzCpI8cKOVdDGr4vy0onxK/WB+ivXfrBME
mMTKWmwPXCPaWgyRkbcZuHX7qd3jb0VC1asqm0KVEKVh6Azi5fXt2FBg4hiQsjxO
n6a1cvEqB5PUJKJAV6PgqlRbneONE3JgXZ8vCWtsY07VzUU3jf9RifyGrCbL8Vic
YrFmQsEZllgBxmrYYblhOofeOOPLXOYRNbWTC47FRKiE4jwjKn9EZYrDOj+tsq5o
Z7B/GwolGZPrZFXqbSlcq+gIvUdNSdvmDHUtFHHz5U8Nza4RQ8qOB7ZBPC2ZZMMv
jPPsAXhwJJAFLMexZU6fzTIFcWTndKy4p4dK92gw5q/lvKhG1HLJB1LGqeTV23+4
VOvWm7xfCX1jpTTMIB5rrZSsZMjDqg4OwRJZ6UwcaEVUlYvzdTjIqs5hGXQGuEQs
UutBfNAWSpAOWUJMuUqHjsCUQYbKgFHC+olFf1T4xwuR1fYVHKj28kRRx+ayHQYr
6F34NTZxkOcytK26uKToqDHJhPuEHYEHL9eUaO/e5DdGvypwKqtT1gJxChUYd0u2
8AtERHFHJYfToTavB+hKfUoeAX0zy5ccVfQIWw6/dD7Cl4gz/aYOa1xYpD0qGDv8
6yKoehSK0mZgppUWX76wDEsivlX3EE17BXSKo3zEmU26IMsAVaSJLPlrlDJ8mIaq
Ns9c62pAo2K3TzZi60SHDuDdUFjniT9tjL5RsCLJA6xfp2w5zu6jKw61YzC3phnM
eBaQNON2R9tfQgRVuz6FOnCMOEx6+jwwS22qUDaQUWa00a9B0rWtJmYEEyeYoOYD
FaoQgs+Fkm+IM425YKd7SDmt6cSWaAbVYRxf4dxzi0tvdWQnnry1KUrcVArd5Za0
skbiXSfuEEzqg98Lq7OCATJUS9Wh91QB+bmNiLwSytBsiY5LM+T4DNX/zvhtqErt
h/aQeKBD/HxRTjQVrzLP8d3qyhF0H1PBuCvm7JAK61qg4pHc2EVkuldqp3Ekmurw
z2rbIlHSLNjTY4CfRjvlHPuic9Ytmicpr5mA+stTC/F2yHzz4XPihB1tJZBZFv9B
uHBDhNdgKoKfN2f0OERdUEcCFBmgBS5vd174s3CrSp9TJFV/5/DvctN5Zd3KnumQ
9SaOjh0Aw6Lavg+2p0OUrfWfZlM3FbY04Y7lE7NGBfa8p4B/6OvpKcOKJ0RwtfC6
fsDwO0G2C8JbTKfvgAEOrLuZZ/n7uPl7WUI2cWtNb/FqbmwAX1rxD0C2x0oMsoJz
Ovv2QvZURPZM3YTQLFKUblXNa7+DHkKTfNR7puUGf2yh4XUhbZCn/TGx/uUjq4Nk
VzXiyDiFkrinSEtZO10KsiEIa9ar8a/RF+sE0Q9P34ygQ2efT/ktAXbZHvQ6hw5g
bXc+N17JuuasyiLF5QKVOWszydvU3Ss/q7Wd/IDj6JhxUtbcZx2DY7pskTn6Ofvm
CQ8SuBJwwhRqjZaVJ2DoTFnHfqjt+Kr0Pmug0NYn32nTfUaovz+NVqe1ElBgPDXA
/IvaqkjoYWJsKP0swR9ergZZTMTMr6QdQmXV8joskelNdk7QMGjws/DbdkRRNXtC
WYRpuv1JeihzzBAWcO1J/UQloMytPIVSfBzXTgdNqsoDGfiLP4MEmqg5rVp2jHku
YgcMXi6R2OPmwtfs2aaWERaZiaw90CSxEWxXEnPr3n4MXhLL5/ya1d0CjEQ/KmZ4
c/f0kjIekP8ENZuKQU92IjAXu9uySFF3IUJ7MEkHgRorng+nUPeFMd1s5oEHcnV1
Zo80T69XpNx9lUenpwnY8QRgBVj1D3z0qVvl/Bygo4pjKbFe/KtrPsNZh1coGiD7
dqmLOHncpsVR6/UEYDbCZCLmBR5d/mHgrCcsfxl8tL7aEJ32u7Ff/bLFlT+mOka4
hac36i3m3dMvfgc9bIJFGlTeKZHL0NvWMr0G9zFDlWLN8wJGgJiR20fJ9ivFP9V8
pHPmdb7ZRya70AvciuxPPDdA9R/ScBHFanuU5//TZOV5CTL65AiJSBJXL1+zIIcN
pAD2T5iSFyYFxBQEBvaV6MErf0tGzhX+K8T76tuz6AzNf8XMMd84AF33h7VyztKx
A08QdgmH9iBoqTVqW75lQSMrhUbbDTViwsJyIPUYqFrl6JMLElT+G0G7g+cu4soe
CJOPbhQ3O2aHrYCYIi4nCXzEHhNAGnI/AqOIHwieIbjz8gVVJQFKBbOJ+DMwen7J
D+G+hZqwCmp9oOe2NPBp564rEoC8eAFoXMbY3XcysrhfsA5gMSpxMp3QIjjOQp7c
aKOGco3Ofc2MP5dJKIX4XqyWdWGQV0+CF/RdiK45dTw7vC5RE/X1fU5ALmHzL5B0
wcHLHcQuCo7m42qNpTkkXRXXAUqh+4Q53jp7/jWkT11gGcolT9HUH09iHCTaKHpA
0jxxfSW4Y5vN+cs4fz24FrtaVj3IkaApX7Brw2jhCw8m9/eVfvPrBIE0sOzAZQa2
HV8gZtxb97SN1JjokmjHafTzlj1a2tODE6uiOG1CsK4KZzXy5GNmD9Ay2v8YjyL5
AFVilSzdDr2TZdyW+ews3I1LUHy+tNPL/6huzDmIhsz28pgKGc+B6K4VCOGV60Nl
tlz8H6L6Ixupa7qXiGcquiMGDTx5yB2NS1cYMrQGo4bsSVkBcF2uuBq/j6lpnhoY
TETHLR3qYP4w5c/ZzuqniFyaSYdCVroH5KAgc2kq2m2h8b4AB832nFLbeABApUFb
HMsmOutM7N54FLHu9Wx5cP+h4Nm2z42UMJaQzxE63ay1G9kRYK6Xn5sUiJrxkLOP
uXD8py6I9O04NrLnWsolCtaatVGWhZZLYaq5sjZRfADXtmd8ayuCh5gXlo6S6RgO
QrnO84Tbx9i3cqhKdmwohK8lSgYxZlgkpP8eBFips4Z3zX7Q0EiI20BwWitTZwDP
J9GuNeflSt9oO9WeJEAFIUkXgFWcJQi0x5fFWbvtkF2LlzoErN6GxsJww02f14jy
sMTfMTsTpE0gYk+XzgVJfnJq1L7Kpvq6IhdRqEcDcoLN2vECqPdcvVcclRxk+xdl
y+Ld4iuZUq2SLnGSY+3G+33gbf+yqmYoZRRB9cJ0gVZj2parIf/Z6CHXVjz8tASI
8ZS3VFa32Y5RtqQO2FHsvspc/fA5VkAzlakJ6JCy8M8X8epPJK7ifrnGr8cUR2Ut
dgUla4BmiAuQPjjpV8pOE56ccBKF3+mS/pNDODoSuX3EOKYtnflTVNCdZxlWorOf
FBxvji+vTSSRLzEIB3BCOWj9Z+04Aq2YZNZCJ6eTa9MBIilyPOhqjgfko3tC3wRI
4YdLtLTl4l5JtkHQe9lp9vuPrXxRWQOuh4uIahCnGUXUkhWzevrJH5ZhVntib6Eo
kUf+l/gV7GvXyT7tZiWI6UFbxPZ/IfRzr77Duc9NC4ZaJnt29qd3LZRBot2FJG5z
Kj4Jgp2dD21APi4wrLjJjXViLoyjwg38fmAi3a8y8uZel+nlBWH58gIRs/enTfre
rTrXidhx2VykrH0XifathGIXqfCERfeYsQsu7cwiMNIRvzKt69VWLqYMMLWOlbaP
qhbAwIO+3EQK/Vkl1cDe+EFQWHAB6Umhn6IbGrrTFu2m+ZjXT0yOOMKHrAgwhqSI
Xd+nJhesOCIIMfVAEuKN4fxrv6/kRM/cXb+OKBJCq4qvy4VulsLSRPn1d1eYERYB
6GRNBXMk8oHEXIErUkmXiOPR+a0xdyaCktzGVBiFJHs2WBRNA/Ly7Uzs1abs6ret
/Mxfb/+vNZuKTtaoQWcnPCqzTgwWWjIQlhuYWaiRKzQ6OtWsMTKT22N3/+D7Bbyc
XTeHJbj03BazDPkPGQBwJlXIhxtjKswzwicIUeHIzklBXLhlwGTHu1V3N5UmtelO
vEFAM1Zp/LMNRTnYFPNW/mE9wFeHlMK6dyq9ObT8tIxJlDwU32BxNH67iI/GTbT9
4lpAV2BEQiG9gM9HwnIgVq3VrCahS5fhjLuJ10ikXt6wLRt02Wp3D7+RMSSkXz8J
C23Wdyk5kyk6FFievdN47B9WptTHHPe7rTRmu1DKpKxpNHbsWYS5gEsrvcxdxp49
608QLKzmHrnYzQFrm1e6uz16WqJnrYqcXOmu4njm1CDJApeZgSHOukcRQ5dn9MuJ
gDQJdqvm27lU2mmRIQqkxBZ/N8p78ABxfwqtw48+pH7WeIdRyUTzKFpo25Gcx37b
EnSa/Wh35rxxVJhmShJu6Q1gajapPiZbSVGglvq54KpzXgyfEN2qZ49i2v/wdyE9
44P2OwPlrOuwDj4kQhxdy/AaL9x3gf4eKw3Nv/K1gbJ91rxoqTF/ic/WyitjRxqg
VYsKzDBScYgPt1xyDYqlVF4NwzjEqWOWb7Z1SBRn8lZEjrqvoe3NTzbPDXdXBPCp
LgwjGBMqAFxXH2KGyY2ObDh06rFZE/HiJqjXdC8W+WZ26Sg9ZXz0Ayc4tw2o6amQ
diwiMPmu8vB2MhJTaLyGwiWZ6dohXinz4LCMyQXUxYjcuyQtvvMpFopU4fGJTifX
elqjHW/qSSPWE2mpxdvsgsdz0YrJDDElzgwVAQIa1lOp3u1PHzJXEv5NbonnoBfg
VbnekFqzDsml4xL7TaKpGmvw+j4SM4fNfGKit4NWDiXd6HytoYUGVilfB7GXkyje
aeQEAxJZTORvZlsMz/vcl/m4i8jEQk5QFmpH8Q3CqTj2h3+E+v1dBygWFWiWBZAx
J2yFhoATnbJI07onefPx6rK/N4PaYMzhoTQJcZclMQlUxlbnYFIAGvQgPgb1je3A
R4c+10RSsnWp9qOkeBVgSGcOV7FyuD6CCO/cPjNvwtR1ZkCXz+2o3bpOfBs1rtc4
pR94a8grTzHMduwl3oWFIVmE5F9qUtL5pxzxxaQIJJmd9AQu8jFHrK0c4RncHgBT
JpjWBM5eLJ+6fC4HBJALt2J+uUHXYtfizHZEXPlIL73+Wivx6ftXuReFc1Xsh0Ys
9bUnG2Me9hAENNPBDBInE70OjOujh1CYrb14Kn/EjFjjalymeBEnNFWm+uvtf9qJ
ygtGbUb1q1+brVOpmL6NeZWWFTw09Hn4fjHbLYCme3+PktLaCQROC8dlhJ0Ppko1
o+iIaWokH4qyR+U53eafArW67D5uqByjasXvmE08acoxnXlT0EUAweYKnd1ye7nZ
mfIYrmsHtsAwW5LbNDBlQw6xullRG74HZxxqSM5F3ca4X57410Kt5oM5HUM0Lsbn
tHJLlOhS64WfaWYPq3olCLknxGf5hkD4fjL8W/He5io8Kwe/l3W9hd+M4dgvDfp+
NfP8wYXoIsj9r7nQ7nbuKPZDnenysVCQSKkGgOmCvK7Gqj40fBzbQaS091EL02I7
tXlnasEWrL6cjJ1S3XK/xXo+ThSmEwL/2LE4X2MFAjuDUoxFcrOgFFf9PzjRvU5X
xG0ieVbRFUwWMB/9D5zMRjjBIgusErVvz/Tb/t/GCaa+VA/OWgqBvPTsYQcqzK9s
bU/+U39RH5EQJawEY6a3JDYIpm6HvM+ah91HGwJQSPPjpcGqWtuG1cHDlcjk3A2T
SSxB9u2ShxHfkfcsSgick+N6fjyfBDJPDwrcNSxDG29+vKCY4OqSlPZ//rxVt4aa
XPtliCPCUQW+eRkt5NyOKPj6J1srDIdBK8rDPOHpqZZXNDEGM36BNOIYBjYVcIzb
/RLmpzQs5TYExh+jB7+ck5154KQ5HGLPCrWUDIUbGfLesPK2pUkH9ShjPfNGutmj
uqfLmaDZxlS6fJBF3LYXt3PNUYKEb1BQKB/vX/0KuThWOii8GhaFvRg0dC4GlKaK
HklS9V1pfvIDrGwMNu5ZH46wkL7Sdakc86A2Kvem1DRJCdJNxhBvQ9dFzAbBYcD/
0ub+MrfUW2GdNGDxG/tUIrgsUWPJVtBUFNZDQ7/eWTAcO0QiwZVWoELUs8Vef5FA
OjaVmJ+03Erv5vmNYpPMPtdevY/+XUe/SXnEMm+jNuuVHuFArHvmCAOgTruV5/xd
aaG6Us+Tk/k8Kv0mBWhk7gewGhHaTjn7pCg5urHCBnfeytJKi3c/P79009m+Kn6f
iDuTFHN1tKvEcvT4SqY+v/69XwG5RVJS5v3sPlh0W627A58yRFj8W9eL5e2RESCd
qeM4gDZSxjCmIqgzrUlRvmbF3Xb+jwTiUKPpS6M9plWNRXb+cg2Wp7WP2uVlF55x
+t+hqI6XtyNXlQtrxMxB4P0PsZn7ikFrY6OSklY9aRPrk+mBnBiUTP/mTkD/spmQ
aYjYsvK23wPtYLYSZxM6IoJObfiDCoJ1pVtr5PfPE5zW/hjcEgVHh/1h4nUvov7h
a0RVp3DxigMZLNvbwbWJiEi2o0qjKj2mnZAmBrq+kDIjRIIVpN4EZiibTQLhDSOb
IrKlkCTVOnujWJ2EpFGiyta8Ygw2fnpXff7RCHUuyBbaIoMi8ZCvogMtbcmtjy2I
YSaQ5LEt6d2A5P+H4QIf+nFNRYAoiBEpvzu8Nuul820XPjGaEJexONHqCOVvp8Y9
UG64HpDM0yXXbxgxfvagLcfxNMUYUrdQq0oV874Uj0KLpBlLDKJmYFXflqjKBSSo
cqTpjBFhgAMdFqEK8/N6AR4v/A9amvWxKiUPA+2nENBpTVorCP5NSC3XjPrRq9Mz
+IYQc+1BPMO1/pfmUiq23oflAhPzSC0ftPkcjbfakDfUZrwQlEIyXfDy6WqhMSis
Xa8h8C/1HQYpZMmkSjleBXI+9Ibm+0RAdM5KwvCULE4Xord3vrKKxFyaeY1jNmw6
zODKskbBcQLWGnrNMpSWGVE45h9r3YrfbcKWZor3gwTmk78zn1o5Lpg8gGF2atbZ
0RoyNJbHycXnY+BFh22w/1/3SHPOPn41HLcmJ/vcx4al++n8Ka6y8Ui8IqIVhdcA
3+6QYLi84QCa9FAKpe6rZV11E0v4kT0ObRlJGFqqFifOSSsEVqMNGMCjtzxLikto
oi/J8W+FVWsdBk2zl0TNi/ipyEN+BO7BwfGlSg9iCDCz8BcM88AsjPSh6+6eM/JA
o4i1a9AElgP6mDEsXxGfRlm32XykeTqMD+GNjNlsdlHfmtPrHKIL4/x/GX8wKyjV
Mv8o7vADRV0KjLo+wbvv0EU/4FJxrCbjjINbo+kOIABv4wTf1c0i7Shn0t3a2te/
OX3pxsLv8ECUrh8GI4k5K3uacA3dc0kmRZ7t2P1oUuT8iFkWJxrT+kyumZlbovjw
7CP6wAhNN9A9+zrm8p3RmCMpioHq3LqQUzwrW4b3PEFaqg0tRYcQNNoySmKVdJqG
oYyvBnvftZybvNnQeIGpK4sbGm6DPNfpt8EbTfPSXajfGclT9Z147Ld78D/jZU+O
4UX7b76SNl8uW4gVqyk3U1zQJWfKsKJAsfJzp/KcNpjwrBehZMceIkQGBDVYmOi7
qvRcLmwdzDr1atnrmW0a6YaESjesyEbECZIhjpBUZNnEGFZlZtNIw35FHOGwNXkp
mEeDvTN4WRHovhBboecTUSJa4EUFMCOaH0wJs+FSSNHBTKz6dunzCrnqax40v6Wp
i9EjkyUJUsCqtNFS7EmOZ3L/vMLCmggkAROpQvr5i/f+0gXsTauY/PcMUIWhqKB0
wvVBEs1XPvcZlIvRkcAWaDC1V+TSwMWHBH+rtJJPkLP57s8zGsaZpxTpYFRJXJCg
8LkL9FLb1Pmlkf5SU4OQRpXSi07aKNWpsfHLyw5KnItH/GWhlpkrcbF/dU6a+Q4l
lr8eiX+G6oSajgsc+DS3Dgz5YdYplSV9KAzBgE0v1hCyNyRzm6/aGQVplZ2cdXdp
Rw5Wp/qVMEVQNPLma4+seOwKdryS/txM+U1u88/y95H7I9Kqvc2rusEK49WsISBy
oApaLke+NANZJZ2YZMFKCoc5/L2vySJcjPpg3shpM7i4BmNEgZXEJ4y8aJDjfc9t
Pda4is+8SI2o+cBFeXEXg/PvCWdcI6xlbYyt/YR+FuqTYWtLSmGziE155rlTPFTS
sbYVEu2hapixwHfjHKCw9g/LChzCxuJlsw+7Fw2MoVUnuf0Evn22wdcbo5zjprUi
cDS/d5r/nQAsFfPax0Yv5j7t2JFn+mqD//kzu6ez28C4vCAPTFnCxWUQN/+K1xMC
yFuEG/szLQWsTeWUPVmcCguna7V0a3FLmuM3lOSOofKSUr9gtpwwaLnmZ9AAp5Da
n/qRPRTLcfPafeP8Q98Bvp4L1KpQfb6dhKLP8mqM1Z0faOzmziJVn8lL9W397sI3
QHwaEJ3Fo+CrsDLjtx5L5O2kDeTsspuJLvHJ3R+0CAcGDHFMaBQV7mB9edtij43w
9NAiFM6EpioT4A4G33YLX91Rr4S4QXVERFJbygdSBjpadL/bgyw3Vw+j4h9YXifS
bNw1g/ploufSxMSVCRNJrGy1OL8yi62y/yQ05goiV87EmdHxmDLdOFTSfyyWRCaH
1G9HDMiN/8z0OEDa+LXSSKQuGJcsbPVqy3ExS+V7nOk0nJVYiz/lsJ9pJq06Opgx
eueKX0lUXnTl+1gwPWFQnJ8WoGOp1/EncPj5rT+IiXqXNqwXKAbS1+fzaDhRtPRo
PGjVoqKpfgNVAQlFtrQzKlvBmU53OhLZ8I3OVp5se17UhhKi2mWR7AAx4KcEDs4X
lT3/uqglKNfkggpzSRlUrZKpSIaqy11Vo3X42fd/jOGrncsSqAdpaj7r/2O9Br4T
JOAyWefaB2LLKm2Y1e9HQLBYNX3csEHnVJB2rTgKQtHWQbMpiDqpjZ7m0gLOpa0z
7WpGC6qyB8XiNYP4Ez2LewKsc/qPk4Anx+fb3F21SBPYIwYOfavJT89oJ32X+h27
1uhSUsI4AxMoJaszoLc4QiFjJk4vwzf6dTywGnw3FPsYlb4TmgsITZF9iJrGNLhM
HkaXP7bkUyLKb7RK9iEKAbHxwh30nJ1baLdDnATpjEw7S+un+t8Puyx8Pq7Gnu9B
FJxcPud2ayp5XobDZmo8hUV9KLU6xx0nzMxvnm4WkyIIsiFto5bVKQakrNQDqkIo
9uZKexsYfavVegTRjHWVm092ygx5g4VeKdcgCr5xY1kaRh7IPfeOh7Uebf4VwRX2
77S6HnHuIzQDZ/2dk1Yej/a6S2tN7wPSPz/sRSrFySPO9bDb/FiLhTskmV5J+N9m
XJh6QubzWsP27iZ5DlSjwWWkYlDIJkIKDRHl+ZQP84EYEGZ3ny4qhzOgNElGbvUN
VzKFCMju1LxGXdFZuzka6/OM1EB9tFht4aK8aNzMuIlEfVN96+puXlONfMjQBFvd
zDKp2sXGfikEmMDdJKci6zSb7xrz9b+M3KUDgpItu8dEnShxfoi2aZbLaQWs/R3O
3+xu6bQYftxLzE0SUQpRi0UajYuQx0Ik8MADOcrOQb38ExZW73FUWDWZk86SqchT
mdqE/vuAS2OHUo03JVqpm8bZ09QSNTBdTUeTMF6xCZZak69brbbMrTq8cn8aj3sL
NXJpk1ATBxTgSKOAzpf5IiFnI+pdn1+hnmliTcCXFB7mY75Igbg57ar5pmOT/IEC
sg1qSSRFnq1H/5vpEgKFb1QlwbOR19XQGX2fWUZ9E26qGX48KzmySKpMmtidmc9a
Ta96btDMQaki5wg31aJFMcAK6pKELrQkfKmnBxFysWXPMFk2YAg9jpxf/+2JXijA
7QgXEc8k7CiLK34eveRqtnbp+VcojERfueyFWKczpFKEWIz1pqae6LYMRGUQTg6B
rexxi8V6G4HXYfRPyHdhbfVNZjwhicMXVMlv9fiT6+Ez8CJiyZZoTUWidCYPWnH8
mAYAeUKitLFa2j5nT4IlW9tlSfIdTNyC3P6HU1HNkMNs36FXlTg2kEsJml7alk6R
6UvrC1bS8RGXo5N+n/yf3irjGvlepgNacJyMux+DwIz8QbLeuKdz8bzDYdGOHete
x0lQikCa6dcS/VzMWS/Icq4GqFiR6JwY7pJNxvnvdDqnvSqmZqG3dLIowasSmsK8
gFPGFDQ68wE7QDZdYWJQZtcDAvHjRcLu+tf9L19u3HhGkcoshlNb74vJwXh3kS92
u6SbkcLAtyN9SkoDlr+a+lFeRnL+o8YuQ6nEn8Zr/ARjN4TdMq9J1Ht7clUlTtUx
qtDtj/PY0kznAQDT5oSCmb98X363BxV2dj6S2dNOO3BdyXrlb9bsGRkHSxgHFWti
FQN9xeNGwZk7KtC66JpLTZWP04iSea92Tv+OA3cP7XWNJLs7/GiKIobW/BMXsHFV
wUWDD91YPT/7tXPi7DJetTmGm2q2Ky0lRy5fSfmb63lXQSOkDg5bisWQSc70Y/uL
5k9mlK6IX8puhL7wZr7wEai4lxRQ82OD1NQew4bUMfWykhwCXBpHhyfdO04tFzOt
ZyVAlB5WjqcRaZluPaCjJYB8EhE5qMrc5nXX3/sMzZI31oD8SfsLVTHEZ+U+9aqb
AuE5v4kh+aeFTWgRafcLSJzK8i23DedkjSHhME04Ra7Hm4ybjw8Txhq/nCjuJMIW
EShxFj83oCmTIb0dZybbmkxE2Gl+2yicY4Llsot+fO7ztcXDQYf/A8udlIdOUJyg
9G2jSigWtbknReTlGIeNpHlTnDih3B7T+F2sa/Jh1P9AWUUSewv0K9SBptyiQU+k
EcL+RRXv26V6NAAivi5426oRZlk+EB3Cw6Ix5T+N9x6NKAD46bTyCP55RfJacPf+
ICWb5ZlXdYoXKgcpVI9bzn/Pue++dmnrIJL5xiHZprVA7p/uazeG4zZZuTDzizma
O5Wxmvgbx2ZLVsYZYScHuDmpas81WiRX1q2jY3xoYEnjXLqDXduxAzpiWe6xcl60
ggq0iSWhov+ergRlwbYVxr2fpqETlF9eoYPXrWhLO93ImFDc/NCor/uI8uL6ZzYD
7vmfnb5D5w/sSxe4fac3fgju0j2Jjfd6FKXeEd7dQb1NrBw9qfGaMPtU+w2y4tiN
4m3uYnICQHuS5RTKG1rtfUNtwiB0JWQn2MjqD4Sq+hgMITBwxR5SZJCv4xJLY5/E
fQ89+Ufubm+vrH9l5FTbW6Mk/jaT89JuqjAPE6E1FQWLo783Bj7hA8ySetLfNX3q
WpqHsLongj+0z3f8/dm5FQ8Wq2UdoQg5OtYBz6EB1oR+TP62PXhiJkMjLhi5SOd0
dB+BM7gxcmFlCFAf9VKvWixy+VkEM/DQLdwiOUTKAKj5l5NkOEcKHc5IPLGTQENf
24svdUIRhaXBn6B+l6oEeqaZpO47HRnl25IviBLcinkxbfwfbXycTrOD5Yb0fRnX
zLhIGUfClr0nQzEBRJkX9T54fTF2HF94Ed09IDmbu1SiEQSd+KiHL434HxD/J3pf
nzG5SBi2mSCbub8y6/5Xsz4LYkREeQzaydhgp+XNtvZyzPD4E637rZrxBILicEBJ
pmoiAYUXQGvp66EOZGc4GpqjulIWmE5vI48Jt9n0S4zSFQoE5a9RKyWrgLmQaUu+
2/fkFxEk4NFDYNaJLY7I2H0rXTd+X5cOAn3aKEgzWet/UaSQfylrXYnDu/7Z89Mk
OOz4BBZ3c9VlCGgLXj1XR8PNpLLOdb9MLsWFMnKMwxG7xwYEFE/l5WI1ydlfP9qU
OtIXxsESRQrR9SdlgUntOXSx7pxDd94utgvtLqKFbE3rac2WF1mo9BYVq/zsj3G3
DmYGm4tEUqzf3X+RqH9IfvFrRFGDWeNRx5RqxTbaltX0dAwiKlLfbDbjVR6UOSJ3
BoOmLFgQxHb9nbjMkBepKEZqn/3mKv59NPFLiXMZjAGGR31pde78edink9H80nG3
66fA3AlcwmmAbaIMhHtArnXzTzYOjhZCME/DgmXd8NPU0z+fxpk06EUL0g+TA9hs
vhNijxMqfZ1NT+lVTg5P9bxRiuS4PJXeFfBt40VNITP/MS8mISTZBB/ewtf81Tv0
7d9Zal3CdwqNP9bMhU+2ob7OA5Z9ZNVCMpQ9LV22yoT7o0NlLapvQ7uSzMggwh7o
YJd4Oy+W9qVvqHQb/ExpzqSflWKVhPKtvP5TvdYCtln2jLOauzFD/3RikWfXL1AK
LXhuCUf/MkXshOdcFdkeiKZs+fsoHmNqY+ga/SDQhanB214E7+Xlksr9/iPXCep7
JizIjULEcr+8FG1iW223Qk+lEIdcGhjPRWTJSfu6rJHEsA/2p/FLm/z++2D8Dz8w
t9VONcI+3ZWXV8gRz0GWVcPWkkxl0Fz8VuWaJeqFqTe/or6vE1qlVwLAPoHOQr1o
F9XcpbJWqXBmmZ4odZdS5yHjJppu3I+teiX4K/HTwNG1Rrj3Vr1hjHNbo6lGW1OK
M9KrMGR2TtRLIK1wY4IDPxd6AQP2Icx+Nq2nIHqtShhKWxjl7lEmVSqL/z1BX9MU
ccvvTHFgeT2YdbFXGWqmWxlApNwefLj1MeJKb2eAoR2XW0DppDcjCN1pXiKTS51s
uUc5wtQPRijWNV/y6b863r+j2w4t6E4nRNqWkyUt+lUcFq5uFtuRlguGHvAxBBU+
AEGxBayxshSNl1T6/ilV6THYGe98BvMEPtjXPfFHgl45F1BBQkLueJlTB+f1SUJt
Hm/rNmSRpYWGNgrFOWEmNtFCEjD0wv1eokZkAn+TKJVp+XS6I1v/dXIYoAJKU/nC
zXD1qV8paXAd/wJAEKiK9RHh5TntyHADmcG8LZjWMmG11lvUWfUiwMV4iRPAS5hS
MfbdzQVoznRE0DWZMcmOhcWBtFJJJGjgy2RYwD7bXjwFo0jiTjwpCjbVF5A7t3Gk
zgUJ4pogwNXG8Vvl1kXXygLoSptJLcUCmNOpSTcKezLpdXHBXklIyXqZGXBTTuOk
W6LOi9EKgSP2mC4YxM8/17zShv44XEResNdmFOMXZe5DoEBNpv1TYiH7i4bCi7hF
chiD6Zi/9oATfC9R6lbRUJITWI+DcLebxf40fgiWIrca+vK+ZWRZjl/KONwynyAk
gNWWbyGf36Udy6PBOHNcVG1HPzYoqfmbdAcCICuOMkUJ/jXLMHAb2oboZD+PQyjZ
0buYw8mMKPeeyTcdEhAtv7RJnYzJp4x6N59UEszt14nZGcQQs4zepay/8QFrKyOW
MqV7HWQwIEX6nzehwRRaHUHDq6jPEM0II7pY2NOQkbb4rcbBzi67M9+/mChdZQ3q
D6TUtUWmDd7ZDc9SpzyET6/ZQGsF1obBwIeXADm47Ee0kA+Ct4723mAcfGrFAyjZ
3k2OZjwFiPw6WdKPAJoaBSW/nh0iHpio/NPeWXHCBUiRmk/pvk21rlSJUfqYk95p
opQiOTd+ZDmVGr23yCG/6Uq2MNf44u7NCq3jaqKw3aqTP/GDjE6SLggV/Hz4E2w2
n1TwInDHoWZQrw1BYX5EDIIogT3orLspDcDzwgnTHSu5ssx4vxs3Lt0CYUpamCbW
4DuosdGBbTIZtLnHHr4vXzCZ2TVB+EsmAr4t+1Kyvo2VNXCNCg6SJDQPihpwx34k
aXpU6Y9T8bVGH0pWuAKefLgqxx8QyqRuNAJasLtPNsA9WvXIqlZ3b/m41Vj24L8S
amjtEaU6x2w99XfF94j9NFtwCgs6nkpg8BDeCzez0YAh3XDHm1jBdUgGXxubrW1d
rSv9MtqCfg2aWvUd6ePtm9vIdoMP3+YKxom7Nw+g2H19HN4eUwmAQCYtUG7ie4Yr
Vfwfvlcen5O0e9UZUCDNio6HnhwLH09ZHyQk2JiXWdQPZC0CzDSZtOE7IknZhqYf
FKZhI/lAsl6HVGi0zWsJgTz5HXYihL07YV5wgIXQUVTaxKb+45xTwOSn6G9W9f7l
UfwkG+j9OG6C6f1Z3eGW3HiU8xYiiaUqH7C+nsp7GVJ4T33lu/ntgzZvVhhXqhIV
7KY4hHgljnaQO0a7Au73+zNrRdopQhjnLgowmwoBixSUj8jgmrhd+9PruxacfvGW
w4vR2KHK78hRrWSz6Rw8PBGFuXSRTzLNRMh/myC4+7MmmTmVCEwDigEAKlEaHKlL
7PjX0srpOA1xLtD9+d8tYRGMkFSdCA8rV/FkFydpJQUcUj5aDmu2thYvx5dFuFHF
YnzB1yfqp7tHbhG2l/Q09r0Z3Eoci47OQv+0soXmvefdNIQRd2Yn/Ljvtli3OOJO
KncJTobE/6qJ2d5zO24gB0tyPb3765NqF/4cTpn++6JtVJXVQwp0OnZwvBVS9oku
fsM5etFAI/vhQ9QmVESKXHoItQ+0llTzOd0L2NpoY48HGySnGMvaFZ8OdSENA4+t
/mNBGUam1jMAIyAS771WnCK70oPKuu5lOqSp6Sy4sxyehBxyahcMokkPC+Cv+rpx
gJaotAl8GakERS5VzNxI/6iLGVvq7usIokfWeBb/9mY/+9tEogUWuiXduA/H8rmn
t+SmEPTzsfIGLD6tvVYYMlaCIEY4fSecawZ2XJGD2bM0449/9shaBtlbtPsrVF3T
hTY5MuBBqL+vtKhf5pO0A0VnvcYY+kelQfvGPDRE92zqOcq6jODUZaYzGU6aKER1
/o1/re+t52BVln8ZYqiIIsfSL0Nb2JeadJEyIORrv8cKvjsyBY+2G2BEPBKdwvsF
YB/ZWpQ+x+lGScuvxUgS5+rrz4FPtXR2Qpk+izX88/6+UMWy+41BlG920N4XokL0
2sv/UWD2kkylEack1nx0NxToNmYMA+mI9cNkUm07+Zv8wHuD6zXlxhkKm6g965yj
PtHMxdHh4OsSEjhMFkCpb1bAOyd8tZH/jlwOrn2p0z1X0YXAICXNPCZtZU5AcBdG
gJcG89zgkYDeOLCs5/ZQgHcSb2M6O3IwY0YYfwXXAjlkh2oq23c0frRW6KBzsx4L
SD2dVGi/jyAFkc0MCy5hKIKaGjbBqDU7+x80X+ZjdhMT+V7k+7usyQrP6/NsYgzz
cOfOn1Qo+F2c2Z4roSIhmHlhHyOzAz7MiOUT3UJJgEJCI1YnbtOzsMLueEDpFOC+
ArbnIVrri6KztxAgmJ7dYiDdQTsteA3P9osUHR3yIxrSHbv9+0Mw41/2pkGl72xz
V4kNNA6F8AXYgtgb0B9heHu4t1FbqCq5mH9m0v5E/PVtweakTuAA5X83+cZa3jnQ
4nFUbG+yQSPmx2ptDwVBHbUgJ+l1QUOo0v05UHpwYeIEb2dlyGss493mrv+t1ckF
4aj0jOACQ9sGgijG6kxKo3ixJIIGC34Gy2krBVAjMW2vpCKKfrI6Yfurus3AcUiC
GubRGfBraNEfpfLqNJ9n1JZ/yhRIFYfQSFf3hc2/VarNKfx2mZNGFM7GV3JZe2M6
7phFRUwupBTcUP6/NC+AGPD3uPI1D+gcFMqrmZbG8nTl+4skUol9XClC9ymf7bz8
l7tTWgcLiEvl3mJUjDut6zvR5tq/Lm6uUAJ7n5Jvf5g83zVcTLL+5d1FpbJon0Fs
XNpvRgYPk6Te4nnDe+T3N3Q3fqlVgmUZmS7lNiB5jS7qrsuGdec8iFyvOxZpuuSN
hPY6SOAIfvMyOh5hmZR0hgVxGnVrEToQHC/nH+0ghkeA+yyYz/kNxqYlkMjTF/68
H0Va05lqgim+7rV8DOsTn5atQ6D7AbPuqwH6++gXc563lbIoWep9/T2lfNK5VzZc
D1YiJnNXY/ZFw41el1VRuvYnZXei2rrYiJRUpfNhhtDs6gkubLEOeAEnaYigIcV2
9AWadTn99U4m0IlngDarnTViVZbScmz8xbpaV7lFNInD3URakg6W3vR0TWIdkFeo
JhfggqX58QEwiAL/7Cq+OmH7bmlr/PJ9BL7FbfK1SHLFVCq42cSF6Bnjm/q/yKQZ
iEduwM5nOCm2205E2biXGInck3Vz8Vgx/FEn+YnN9GhZdVBE7NAHHovz+ki7Gz4y
NcUKW83bNHTDQstU9NJdSSzkweJpVxExxkNPy5rYvN0d1QrWs0mlD2zl59ECzycG
nYhNDRvJsKr5TMyClyecKdrPqPw444cndEuL6Jr/9r154/4Qh03tBLqPSIEI+qw7
Unmep34QfMzbhw/YsH+Jf+bIn8N0eSkiaHmUYDX2ro5eesrG80ngHExiarryinyq
a76dbB9UVsEs+v8X0C+5omyCYoMLjC8OmZVnIDoY2mCBtt9YrYyQjXWglzGx/4mW
PM2nH9w3djuVt5WMFvf8WMaXASGgp4zQ5l4sEmT8D5h4BJPUEwiNC26ELPVdSqE6
GeyLwbM9qvtXlDslNPnocdafzIgOQw8i+YW0te0mUJC32aV9vMvb/ijoCC2M60dG
uk2jyLMGG09jS9tyPIf1qI3Mwy8bVZZp6Yb/e7X6Pbc8PJzh4P+FxzfdfNs2xLVa
+8ybgCcZPMPO4rN6sbihGTnxKcFL5W3FxkA8depYoQVuFCkL5hVhJpYSDvdnzcTb
5HGO2+ivVGZMPnL2+INvniIuUZYgEz/oKlSafjs/NK+9JxdDIO3vq8q2iYtVq/XV
8mvVQQeAGlo1xpfyXmkADCbdFVRTaXOWmYpSm7fEyNyX6SqjqdnZtfxhbl2j9zc6
un9qXH0UzHxflIsBhtrlqJSXxvSWgfi6VTRMSZysoX5mDelxtini/b8oxoKPXian
gE2zth2escWi9DdOPYX2QgTwtjBhzPBsrCA/nsrYRYnBoXdXPstGH4Lkk0QHJ+jz
zou09VT+LRIfbgeZTDdfpcC1OJ+UP/sM/u9N1InmZTGp0Xmo39hpwlBm77uTidvo
FttmHPqfX3682ykyCu8wVOnKk4W6BpLADQzmpl7VgKb54l36VFU4P4oA58fo9xhD
lTgt3XRNAte7qXVspUlAoxa/wlH5uk9RR75r3TaO8MMDQiqUnw1CGB+8PbUXlWoy
A3sEuPTV3qW1ZJT7Pj3kbNUuLYIB/P1ZEsME16gDyVxTA2jEH4gclW8/IX9c2mXJ
bN5Ec2Ab+emAnAvtjIUNRTefoIwN5u44a6JDGuhxXeZBPBiiPNHN8MTiK1vN1Y3E
qLreIFDCwLuIzS8lxTxeAkxAceLlVNN9VBul6tZg6vyTJfeFpbckT2yQF79JFAoI
ddHJfFknI8/oNNzC+XcACwv7jxuMLyceEzhcYf7NlHsJ9nUa+PbznEh1sbm137SL
lIHEAqbAeGD3uqlP4bfd8LASgvgoCGy1vai7wuwmAUhZf3OgK138k0FH9rtLndRe
JLw897L3Mt8vYlyGrMYR4qvaAhufOCINK3T2S0uJg233IF/veO8QvV4BHrhRh7Ec
OyFZq2u4cwOqxokEIHfk3cxDAoOOysSkNdm64KQmC31dEVney0HBJ6t53G+MdHGP
1mikRWP9zAfzRFUqb3aAU7PWQObwUyz8zjfpYbeN2688Ymom1BtYYH6UkvkQfrxs
0d9aXBM+k5YcDsXuy2pbkWS46E+Y1pRW5/J4r7xhcvRkRgf05sLw4/omFiiPk6FS
IDJnvNqOUEJ9ZJDy7IOEznlugbeLO+ovjrSd++Vf9wPp2ZV8HtkZWDnqmmX855EC
iZcbpv6iK0zzWC/YcUE1w7/9t1vpAkkGPSE702sIR1lTPJzww9dRqJ5x79k+w1/I
R1+oJ0MVxBC2WRyuJYefIavDaugxb6geZ3PnNy2FoTVk7MiVtTpZ9evdf4GyfQgV
3X38xrnTBn2vASzU235QjUGx1Ey0ev5Xxr4Q+kqi/rCjLUFl3joI7J+92MGEP/V0
is+F+TuYG6AIT7fKZaEMvmFEwOKt9yJ3sk7ibD0su1qvWDVPDa18QIVHGX4HMobz
osJNpMHCzgQvRv67YD7T2cOXodaUbu/VbFRm0ifyTs1gwqL5AWQwAdnay3LA9VY2
H8H3tV1TIH9YiSyaOiuYd6EIwuhWa4Yo7RpzvwK8fbkvVbk2xQ8X29EqpkM/SXY+
SGbfbiuwFpmuWUF5jo8q3t5oN/38jEmjNaLfAUZ858G6nuSR3IYSYzp1AHwlViN1
nndTEvl3bYCrimN38SVcmTrtE0Wzv1muVFcPS34aA0dtKZTJKvaqpVn5iHzk/R5s
TsHKBkAAAP5R69q21iV5oFNrbTMq2lAfuL1I6j0dnfUrlkcMrinrk0ckRFiCK9cT
R3+SVl9I4AND9OqTtPvy1GFBND1GY6qB4y9r8VFpueYr+xZle/2z19gFfxH+0Ir2
QEu/e/igJfHvI73+RFFpt196QFAJjjivhZtcIJC4AloNWHHN//r0y/dUruQFZuH+
/5zIWV4016+Vp+Yfcae2UVgPvVl32LuTznISBzrVSdN2V9+9viuWj4+oLGgmXFqW
jWPch64/mtCr1XfLAG8n1MHhUQtyrMWal+pjWOuLfkg1j3XS8dchEtTfYBm4jo3h
eFMCXGFdzdFxMl8IRdRm4zHqNUF82EwVgRVdGwODkFASJenxKlPu3TVkIxSLzAwH
l3uW+rTJRmlHShjbsZgkdv0UGk5Ue8g5uRvWvdTSVKMLcu14fTyyepB/4XOTRaOJ
jD81+iU3YR/kOZdQxpNp/FM4EwxulACmZ+haQrIPivPguWEtzzojvdz9257eSbEX
FT5b+e2n80UWdOGV4mZ/lferGdcs7m4AbKCZfXhROujCm0x4pmPytGeBDrczzBKO
w+lq5Xrd2IQg1bo9b7YoS4mYCoCmpom+/z/+/2vdrarL6mgkcvo/JXRlME+/0Mrn
+Rt/KCSUuwKFBlP+WmzYQIsexrJOwOJA/JucQGINL5SCn1EkZkQ4+1emn5EeQ+DO
dsIeQH17QzGz+Ur/4CxS6Xs3//3F+57mIOAJVKqCP3GyNRSMUEDhoT/hXZsCDN1L
12jU/RsvGaj3p2zpV+3pr36XEgZ64MA2Lu81wStZFmeIz2wUH4J6q8mx+twRu2Sc
KNWa/O/CCiMddre+f9Y0Bzt5DNvr0601GCG50AfrxrEBasvhKdSC6CWSOn7UbIS/
9KU7P4DdKTqDibNEHjEfJqMxoTqLZxyroCGoit1XNYjOYu+NNqeXknuz6Ojy59CK
B7/6/TJgxjHbayFTOV4Pq6Hp927uM6q/9IQU/IBLfDv2kIaEeMWaJtSeV/ncaiW1
num2E+I9NCzlzrkWgVAeqJCIByUuLcgYzOTOOpDhFWdhv9j2j/G4yeQHdD8G/WkQ
+A7CaW8NP8TkLLIsNytAsTFJQkDC3svWtd/sxUi6JC2w0qOvwCy0/7N0GbuZ3NvS
bCjdnckq2g/AiFWEe3shbG8wJQ5aLQZVmiwPXtWr481+H0Rqa1zEyJCAnEqNDqvF
0yTuVQJU2ULw8kiN9QweN+a8UMR7In9UEeVYwBPBtGa2Hka30sKDVcrxuAoENvQN
cIUPpw2GJ52RWUVn2XnToOPE4ZOQzrey6CURWPp8my9j0rdwAgjRjP9zqdVSbhaO
SrQ+8PVwUvkr11OgM+zQgW22+BYFkX4neqQ4MTMyZu9NuxIgP8B7XzxKZxpW6sfK
0dPzjYfH7F8FWdMabVSyZNO6DxxA+9Xwd8Mnjyiay1R+Jk14d3PQ2XL9gc6lMqUR
9S9BjyA3JuS6tuJAxe44aGJ23K2kdLOEG3DaRoaA7hL6AAeTPZhEyzzYcJFZYH45
fAeLG3vmCYzbIyPxFcw/dA0DuungNcIvRltn+x4KPXT9Iv6UXuu6GkQxmBU3wpoK
SkUbP7+fUpydUlTfce7FvgzcqWsvHigutBvmJj7viO32IROPDo5h8PTshLp0/8H2
aPs4fNyWUB2l6TdPmvchZ+y3+IxZ642s7n+6qpAbdrRrySK9hKEfh+HOnayHFu6l
GE6yIt7SXtfkQi7wkRVGW8nu8jEK4KrEv+pslfsL4Nkwz9vQwegPHRf79mRI1QPh
8mQmcem1WZ2Q1F+K/1uUXLFNtAF5YOlzPtY6yb1v9SxbdfilS/8tq/rL1RN9lu+8
qxe3YB/JooH4Cb7IaK5NWlQXQA/rF1WcpucD5+pJRBwvbQPpT/PXzisFXV6NZOMu
mbpxpcT2S79SPsXCmWiOAleq+rppljWTayGrllNIVykXlfcDzb8/h9UeI5KgO1lA
/kqah6QWz3Ttc6wDwppYbUB1ZWhifkDcvWDW742qQP2d0S3Rc7W830QlcVP0lN5j
PKiIRCvg5qzYLjurUT/6XDcXTXRig1u6LN/InKtKNFZTgdqiKSQ/2IeWAn8VYe54
pZkicOyP+odA/71AEZJbmlPSrzfUw23TgF3TrtGAnr1i/oDmf7144ZRNcQ3aUuT2
lm887nItXkntw2+8O54NutNvGBchb2ZOZsGCQWLUU1t2q++0++E++r2VQF4etRuP
qy+0dvYWGmA/WWlik524gzC61n88hL6rUAi73jiHBJXaBM/jO6+RpTRhhg3x/fIs
PjqPW07JtTGQav9aTlDVH5nkxnNXTADBo9EiMmjF8yIU7ZTcJJatyaG4tu6ixudd
j1x/kXD6btMCN2vKH0bdyZdzfM8241xqOQ1cE6RvHp2wQkQHYHSNriDFIllG7X1j
9jO2cjrBqDoDD2XqIgjQZYDNGgeuqz2mtAVCf3X7xaSh71ThrWAA4Rb62uqAicQO
krtWDMGGfAF49KhHL9gnRnWx91K/EfDSzXTE30VfrNerFH2jiDkanY6V4EPsz26V
GOKB3NWxUSJcwBtuygZNwoGX7a5G1PvI951e2BonV1xL9sDII6pZTSx8O3i7t01p
J7ZT25c/rKirKOE45hQ2w1omaCKy3M36fpGrrxBy4fNt407cL0izzKoelTb8IkRp
mleQlQp7YguI10vg3Jb4CwCW8uxis9aUJ5WnsPK8GQF2eZRm0/RlBlmAvwu6bIEM
mdZS4sNL4/ITxk8GnLK67Bu18StfrQNmztRft2NmMApRIHf6JqId0xITCvvScwKp
XVhMiXgBTOosvJqrwcx3Xzdk5MXOTtxgSL+c8CX87uMM4D3xZHdXrlRa2RvhuQy1
LZeRlhEc62a+iwHYUCO5KzDYMH+PNuASNXcggBPt5aybaGCBckaxGd03Of8wxKOm
mUkiZZc49KqIj6uz/3b76njYF6oNaIiEGeK7o9SBYeUgH1pIOnItrX1sSqV7SyzS
GMETuY+dZtOefzsNdRBtBOX5GGGhDwwK07+xkBEVtDvEZ0/xUk6iJ7Ly4WgRy0Zj
TitQBoA9s12dvqmFzjUUGXxIK9et9i4GYzUeHAgf0SwOdyaHdQTSkgmeQYzazzpw
/OryXYxuLY/ethqvVA0z+201aLJMG2G3AjkHQ86WrGEw4lNwhkai0FtbyqOrzMp5
AyiBwpgzePXrhWRBHiMIGS5c7050wNU/1VrohGd3MV3peseUFy2OtqmVhiFKIQ+i
QRBsoeWM0GQQ6K13D8TvayMe7oaFUg61qUI1iDJHYa4yLM7mEC68nvT27h+YDHu7
e0CCotnhpOwbfUnvNVZjOD6hugokL7G35fv9unn7n1NLTbLeW28IyayzNHsv80bP
IhfWXNKFTNZ/MVDin4oJSPvit8BBW5BLKWLUQ1Ey4wNGcRwibioR+q8rb/zcDGEd
y0HRyh5LrsQ9GLoB+MbJtrl8ABpzCzsF2Ya/gVdnTu7i5gF6RGRt00HQo+uRJDoX
bObkYq7JuLjo/bwKzsNr/TKYg7JtnnbGdsUErOGlJcd+m7Qjvi6grcChVM5YvK2Y
VljDYivSLP3URBLlS0dLLIhKitNNRnPhTr6vzWMeA2Et/ow5Ort7O9H36Yj0WxuJ
15/PPwVAEdLsURRWw9WvOmSD987LVic01JlEH19qjf5qMWRQT1J6DW/L3tqB7ppK
jGOpyXoWlWXpmLjxqeSj+EFFTmfjkFaXLhYC2drM8HHe8uSeFQlcfuPsm84CT17U
E7rREiU6fM8/oueV8/kG3qdSJSEw13R6ByRKaowkHnWY9YBCzzu4Xbh3SZYPdcV6
iFzd2/sVfBOotB1oMFWrjmabDui1RseS4Sras8ETHfXU0BK4KP03Kh+tnLClKhpS
OKW+x5AIZ4u2xfWlRCbPMxZIR6oPVftoYy1+h+fmtCSAXJLYJnnf8iNwx79XuT/8
FRDOz5oCLTfsAn/Xnllq0v66ar5IfGBhLIdihhpRiWogjGHDw9F9LX4Dq4Ho2Khl
4lywlI20CCwlbvLAz2agUX5CU8s/75MY4n7V4eUsyF5WfBN3ZiZY3x/ijj5gHYSL
eTZ8Hz2hFPjpCBAcwMT+t58EY+7V5mjgzi0VTgqDVPT/EPaCn0wGGvjurWBj14JJ
qJ7wxhwK+DtmM4zkt8Itl2nxOJPVGw0hlseI+2HwrIwpIDmBkvYSvzEX0Dqk1Z5X
ufb45iFXqw9GyVsERD8WQwOvCgMvETDMphLMP4BxkGKeKNIxoU3r3uUDNvavq5J7
z7GesJuPIGoEViNyzjHSriU7OfPBxrAKmEjwtmfImHMv8M1AdgNfLQIcafjL5mVU
yGSplBOH3UdhhjjuCxQwHxdeTMWu3X0bTZOh+wJDHv0ZAysxNwfhKcqaBIs4WhLa
wcHe+NKAo9hZvXDGMMRtpkOtbyVb67/c+5n+Ga2LwiA3+cvblrBRJT4mmCgsCUl8
7Y0aVJiUNWR3scFSaIA4xZ2bbI2vQCm/ptw/l2f3YZr8HM3TaxUEBYwFDcxh3qlD
eGwi3tYQW0A4NtLEon6L/WlRN0JErd3b5PDMKdIOh2Zl2pchX5lt2NBFwlihXUp4
/xojANW3QIbAn5ksC/+PpEJSEOGEGr3dHiLLtoGx1fFfWL1IR0mu2qQN84Au2dN+
It/QRm3pk60w9zsFb9dJA6ALgAvhK1GwoAZZAvXOfXPlNn8UdiciEQbIxnBWqvpc
tjaSiDEohmYVrzwvIZMm+o8G9p1fxSG2Dz8zqirNdgrPEiwguD7egsxzgO0POEVQ
uihyMhZHCXnGBNx9kGw77MYd1kJXWzVQ6ZTy2LgyEE2eVkdjGRlfYe5+0U9+5/1X
s8ShEo6wYpI5UYp+SDyOdG2IE1CJNomGmzyivwklVlPSEupnvEgdfxTMCtS8ly9k
LGua2MQesc8s/IvzSF+I7zrKFZwTEBAlSe7eQZ57xxezbD3TGAeOQSDKLQeLpFUi
Fv7232Ukf2ELJb27rj/W4uZfXpPhY99mX7IcKnTDSuYUt2BHTRvAsneERYlajk9o
ElikdzixO2nhKodmfEQxQahXLvgJ/ppJab+ey+SfxOJFHXXtDUVSQaVIxgKZYrkx
1CZtNym7zWG74gZTBWx+VOqMttTZMgWEebE7Pn8QKzgMOnu7ZzyqJaKe7iIKFXqm
2VlaHyaBpO/AwEYzDarrUNYi1VngAj65tF8TwG1LRzx4ub7ugtZ4WqeQC8Dyb+o6
anjrB61Hpwm64wyUv4Kfa8eg/dNKRh/KsVDbklwoR61mPnxQ4q2gj/7/9HF4eZaL
DEHGDy5e3pcql/h+mAtJCzg4kcASkTCgay+ShJCn0lNgLOTja1+1WD1izMkzVlJN
IV8dUyzWj8cdynfkGBwo3teS/eYsBAIWumYrHROp6L2a7LglC7RJQWOWOToXjo4X
wSxUwr6FTC1a94GzSJa5nlRyUVUg0gVNBEhuSgAFVQaZZV6FBUo3yBjBBrc6DwAO
99ltAX8IXdb2u0kDJjPafKQAMyxjAC3QSydjQxXK90c/MRl1MH2zGU/kKADwepCl
sOFxeFML47yXtxq6+N+QlqKuLAPGGqGzwedUXSP+sRIfZckJkryd2Xokj2Y5lEs7
hvIGOQT6aUBAD34JA+6jacBc0+ynItN1gPzSW8Nv0g8fBtKf/KN+vJ2Uraye935B
riCmx2tOgK62T2aSh6goqCGjzS0e36fNHGfBP5xEF6B+nJUiY4T3o1YDKK5mGSzd
W6ZLHoLrDvMRfZ3QxNZ+ILgTn9n2tOiD+CXVTQRCIoBmAKc6RxC8GphJUcl56N1x
Aj5AubB/3fbpT2qlEMKKzCyR1S/ZaEYafvbNPCt26lPMEcL+52zaM6CqSTFhzESa
22hWq52bGJ14prmbARboF2LK+PFFyMzo6NZdaxsyw7os6g7tCd1v7+or+uIsTJLB
IiHFDK4Kk2afS+YZUSQRHHwcWj5AV9cwLM6OZDhpl8XMgYNHiU1pePIVTtO6T4Fp
87SlRT7Vt61gdiPhqF2pbDsWQ+sgG10s3e7WZCCRU82VdchDmKYn8isRdjdrZbjb
NYMD2G+nVchb6YKpu0AyitWHbs6DnXt/AMTnZX5yTd62mcmv4XPNQoPlyqx/glRF
tvMlwmc3YpYPpjj4Z+xUdXajCnJG/T5S1as7OYzY6uvz8l/+JrMMD71PIjk1Be0u
No1/GHzzuNDrp0LtC2iQMcwQLiJDoitz8sJovoIXnAFHWIEGqKatNrOZT4YGzAoB
B8djQmQiLB56YYPWtQBkEC8ejOSLtaBdLzM4ydMjAE/2xso/PrEdzcnjYpWjWagb
AVcl+g584o5pckOU197wpbE9QltzjGg+vrLEvK/sEMPWhPmQmAeEpxINNUDyyHW2
y/K8367PrTvLbM9VuADSVInDJz2bRhBYiAtVw8A4wF8gPGL+L9+BN4PXKi3g3+ly
C7xePCe8zPsXUbebsq/6hvk+Xapzu7Yscu/Oz6+JgH3dhtqfjzmHPusuUJcEvEPM
rpEjQSVh6V2SwyWvEW1/JuA03wrHraLGGrpDi6dfMSvOunRsUeh968JNJ/KY5To6
cGtQSdhDyMjZJlWh+B5VbwviIHObEACQBFAPcFEUiQy6gqZ7gIzo3M1jSZfHGS0G
od63ulffvbZ2pr/n/o0KQonIITVFtnCqT+DAIFdw5gYjy4keG4hsIKMF4h6sNxVs
se8n7IZdi8yP/BZRKQlarpsyldm5SV7mwFqzHkVx25M/soUVkm59YMsyvQIsul/o
0dxoKAhdPkwqheYTJswMTm7FQUsCRDc9yAH/j24xa1R5zAUI7OgOphrC+R+YTVH2
wvPBf6/7dd2gCR/aHjDLm2xA39NOV8vgYZ2XJh1WmLQWBgJPB6HdlxKrQF1pMtZi
1qQyBEk+/NXl5TaTBayXpF+pHbccWyg2uzjCoN2qE78nbcCRckv4zahIHuEGxOfM
pSNaxxseaWuvlyMhi9Oz3xU10alVQqg3zDfv1CdoglC4Cdiltti27WFMc7ZgrKXh
5wZ+/af0RYjNYIQouuZLiiDC/87DzhL5HD6726NS8XoWiBHMoYDdBVqEqZ+29STc
NiNlxAn1O4l6rDf95CFAj6xdnvt4037+Cglzg2SwlBPmV5sX3JY3uxjXrP2M38yY
rJVGsnsQP/bea37ML/+Rr6EDNtPhg8S0cdDVDhMn9llzZlsrvQjbTxjIpkindvOe
nOSiRGFqzsJRgmxnxozMpgWX0XVWPmmFAE18bQ12/M9PqSFfUFr7yR+I7QjcK4VR
8qAoPWy6Tuh6fT/e4DsUUIR5k5Sb7aUfIqpckJHkPj44IKBh6rtYjCBdNmN6UNhC
mFchKxh777Bz/dxuIO36JFkmCQmQA7X2EFcEjheZKCyoPHGx3kw8IONNGHLccstb
4tlzsIsw4QSMwAJs9FMzKKBFoYn3BrFiJRFCBnsQq8shUsZ79tWN24XdF/F9uQ2E
L14vP/OwOLJzL5q1sMFGSNVRmSDKdUAZIG8UOcxtOgfoepUyL+uRIy3gF6whx5SQ
jhDRNeefecsuw58u/yS8/eqJ9F69DxxQf2rDtQguF7VpI7vCtBuiKeOP8BOKyLLg
RnYkrvcmZkfwhY2ybuf7xR3/UsQ9oKiRC3geMjBpcJszoFEna78iTnu14VURlxLx
AMKWcZKf/ASt9lwA25C4EnoxHsnbLlnk/iAyoL1vO5oxemmR2hHcKZ+hWTLhXkL7
h8goxcUdU7DDKlu+Yn7Er8h4GqpTFWLbhEvzvg0G68MwklxbuxSk2gTE9hnufrM+
WE0K9VekHai81hRzbig4aVKeCtzSUPrVmpsSYh2HS5W9AGieI6nzzlXvoQj16roH
hhzr37wcVdhdQeHk7+K9i3C9iW0YjXZoMw7uUyntQl+vlc/W+5ejqdL/aLepnbDP
S+oSUaGkrZI2drbuJeqTjSBU21cJntLqd2hSTASwq1MS7RRiPtikLxf6EA39oZHW
KTPAPQsBSLc2aRalobCEl9+pKEnbMWSOF4kFmzptamcD4y0/1RmmkRBYBX7kw3j5
ktj6Ru6imVbaHVAawNLuTdB7C+c8OSutBQEShcTJm5p1wX6wAky69JpHxIpaY47B
8Jm0mKd54u9ON9aMiMMepE9uJwh5OyziRa18gkQAAMsCACqrm7C9TuH+xYF3l8qv
fITnq4klaP7YlO2HAeIcDi67Hc7sTUy/1SAC0o+N8qKDlMMv2ppoZVejRTck1WMr
hiSWFa4EaONoFHLrvnOLGUyDnXmI0OEN2CBV+Va9uQWE+E/rDwjQLXEn9ebvBm+e
E0946Rs7Ei7eHljoupOL5MBH0MxZW89bpDEUsLRfkGmQqnmOLKGk5ivbaBcnmH0q
fqFTTdAPuHCYo53c++bpD6Xnl05yo2bRGKCw9h2h5F9c/0th/ND8nSFQPeh065+h
OkLRg+rCDt2pPsUFn9jwy/2xbbqy+QgBtDaIb7oAgqz3A7322KWCc2ySusSytQbX
+VJQcKmKMX946wQwz/t6l3dlnHpI9qDl58Sgz6Ff0D6C5hFGmp1u2Up2EAcWAyOz
SOONRbDzq8c89Cpyd/IX1nv7LAar9iWFtrYYnvrlDRoWl2iJ0rBjeFLnMjY9yyej
G3+FxUdCZWnhCiIYe58MhQQTydoHpfBPg3Lj6ZsuPu0vJH8FLM9rbnt45WIOqzjv
twh1YjUPn7RReRfEnLapLL5gYIVfpFHhMlU8XSOmLduLVWFJX0OR570sJdNO7010
SigvK+Xq0cbd0BZCJWlAW6olW/IJPjtg4ixUx9Z3pd7r/7stanFKEoDv/cNb6xvm
dB6Kxg8g5V4h9Ev+k0EfLJnx3FEb/QEJf+iXemBDivIFwpQO7HOb/EIoD5ZKU13k
9xlhsXxMnIPxKpqmmUPeTjKD2NRyBTvUhIc30+0DT0ECXrLgGPruR2qSCbnud/iZ
YtWRQgc3qHIEB9V5S6oCAAHI687kDoyM5INIhbm4W+Pb5NekGYDXMRWwGyCJ0VpJ
zMRJFUd0HzGdvubXuvZsxx/V93mvMdus07cWhi00w8BdP6kdSzBCHAzsXILnJ6/s
qIO3GyIrcgU6J8ThuQhpi7Bt7ChNFHh554onwXzx1CHr9D/EPheBr8w6JX23qIJU
Fhu2KVck4rV3BbDqt36i2k7CqbRforxPC+jatWOaWzMEqnkX19zAvPeZfceCSQUZ
GjOM+y9B8OiRD81rWTqxSB2PxqR3ulr6/7PEN51vTeCzrV2R+YdhXjuTemEE8vU3
7T1iUxNHZURRMyAVS4akxKxK4fVdVrIaycItnm6dZNqwu8ONMmefl6ESxkek2hS2
9/rvKRyfOKM5ForX27eJZaMWlXjeIVW1O19aspCIHUjYYZvKnVqSdXytfp5CsrYL
Mf3O/e4kPVcgYR5DxunsN6IO2DfqjrQNCZSHECygI5UpjY80meiSSvhNs6hpYH4h
NtzG5stIRAtP3+mb/IfyBDErSBzA/itj2mrzR63CV1iYar9vh5AxfxmNsmQRPDEI
aDlTIlrcKgkw4NdufSn/nvBwpn5mds0U5E4jaY8JCMsecsSG6aKd1XSUKUZSDH62
xLyq8XTgG5Tbftnzx4hhD5Uduimnc2cJm3+HDt1ijh3aXPuiXwCSYa4AmZxQIp/F
Dsw4sElamN18XMIGXM5Y+4vWINz2qCQ1kYbHIhZCZZBJWvnsUa0FcZJuMI6+0SWz
IKfi5smdDpGFkVHn2Wx02uJTJU4r9pfM0Vp9GmPANkuULpJJ0HMW+BHVAkNtFsiZ
XcE+bYIpx1S8MJndZbuiNS19DF8SEaR92P7jf5knLaEwtiiamkbuAR7FD/+WS0+w
RKzbEAk6GXHCVWUY6dkEgx4dbTLj9jzAxhITND6naSnZiW/DZ5uBVdD7ghMpX0aU
FXbpcPvZZ39pg/YyKFliSjRE8qVGW1hymqzxSyx8JwMq3GPu+YLNOwaWvzAkZGqa
N6ChWLECNqqDaGCPAke4E5EURBozOP4pfNZKY5IPk9cpkkU2Mw/3CLT/L7Jp3lra
PzIU1d48m3HqgQ4vpyO4cQmB7FBpHZdgRdqSa9tZnIEpKQ5Hw0t3uJbyCxVxdIxT
2/PH4XmvUI50y6s2ZlYYjoHH885Xt+DCCSBSp7bTGnu4qgjdOXPeUwp/BhWMfmOY
Nb2ZJvd8WXUt3Ehp2NC7DiywYHe/QUOhot/HTBj5crWOg/ot5LtnsqWqcpVhzt+g
UOt10FHQo9k+Dn9UzrHTZBWQGmNcDABPgq6Oy5Xv8WnJ8ARGI79r8M7rBlldDWqF
9POwflhIWQm67snqFuCEsTCJ2yaXf98TozI4IekMqNfA2u4frWknOa4zHEz06xcG
p6BJke4Dtz8g4yuywmhabl9Lu0/eFIXyVisU5J2nymH33LBtp+pH+Mu1mhmhgXX9
5ld7dpVewgG4E5URovD9/AtqEm8+aQYXaKpNmfepNrjZA4wW28qUh4TMe8pPVIPY
UC+LWyLvYPPfylbcZOVM/v45aBLThZ7pAp4sjZv3zz5w0F/UMEKITwAdqnCSL50/
P9i4TJSfnnD/OhVJU6WGMeW+n9/JLrTejcbExJlRQ4WfXfJUmXF7MwWrxXH5mu6a
DUQ5ksXcuStWS9rqvOG0+Rgg3M8e2r8jUw37FTbJS1QXGBuw+ZNxwPJ1OdIXUAgU
gKQeq6bVGj8blS9dEi1zQS+ojJJhTMMr372DluPPosAjZ3LQ2t8cCUQ+0ndSGcFz
e5VgOdr5xTgx+y13QvRCM+Y4DuH02Dyn/KpVtNwf26ur/Jax15Jo6Ur93/AbdwsM
SoY0UWbj5kGijFMrvQX+R/Nq0DeI+LorQYimmYvPFe3HCaO6iBmzIXYckI69wXof
HPJ45f4nTB92HcAnbKvAyyK/mQtYIUv3a6+IvoVfpqyCrbyUf9MpePwlZ08M7Z3S
Q8th2TddfEIAD21dbwRoEtQ9zUcPKppGc2JS+JK1Cgyp9SSKyTaqx+rlabY2uWnM
hrNhn+xAcSZ++DK43dGJwfzvDH9fAstxNuG4RbOxZAf+qK60qdiwuJnZwNzM/lw7
oDcWZyD5FiGd30ga7cyY9qJsVreyTXp/o8I/EqOBKbkVj7MzM+gc7MCD4ro2Mavs
lTz5soyaAMSQ9JJLPWQIZrUP5r5m+6efQt9cuJBe83sJS6DiiqlIycv9fPV/r8Ju
MJ+I1zamCl2jVtsyf8Q9/eNGPRyp+8PhlQwJtPMVOmcwLYi9CEEbS+a498qzZbIV
SItcZedAnW8pLRcd10D81ECLEcXQojTrPhJ9D7EylNLmaBW/sOWcUA3CG7uwfHXZ
sDsi42fpX67uKjx60446PrBuFO/8OHjOGqIwupGGQhTmCR6l4K7PF3GrtSh1dGM/
qlTpd+Tb4kxU52CBQ2fWr5e3Oz2sGk6pD801oyV9WA4t1dfmwhIENWqOZlTstw3D
B+/nc3IqkSkEGu19bMimRkhpiIkA2TmaFrWfQGAZkX3FjmRRm84LFCBhCAGPdW5k
TGJyOtWHGEmnTbHj0I6amAyhU+x8zipVEhDojxi2r9quTjfUyF6ZDvXHaDM0pja4
J+2+3L6dmFwE3BprL2ArVlXPmAJMtnxaMHbeNuE2pDokcjEj4JpPsHVIYghO4ZzN
HoLNfDr2KOdDZXhBxstpG5ufox2lpE44hmS0F4qR+WfLxacixfT9NUhB3YUcfswW
XxmUyq7Ysl66btgmWlPcrsBtpnCnbp112WQRngQKw0twT9hfQnjvzmOhCAIFL0ra
bxJYAaXNSL19GzoCBuEq+o25aaiuDYPzSoyey/s1mnZCoJB8btFlbFsy2QTMPH68
zdXqlV2cy58z7rP40NUDlQynaldP5hkIG8lBGdaUpbr0+vmPoJUBNUoVUR6RLpSS
lV0XgR/Hr2g64LNbbU3l0HTZRd234xd57Q9DTRnaVIuutqinm4Y/IT+kG8dp5bVs
y6roH5ZR9F2yLkRZXjjE8F48QQJIDJgG1nz0QBSp5sxyZfa9gvx6dbkNbwh20TaF
Z9CDMfIQbQEk6qU6/vxFq9YLxVmJbUn8wmK+IszHeQpPRk5OAYAeLYSkWXQLXkqm
Ge2H1ldatmwdpI/sx28SqQNaTJAS574GXibqh5Z88/TCMq+5fGbuFd/ciHpACMtx
x30WtkmEJqOg57meWzVAwyxvcJ9TMOd+73Urfk6z16KYcBcSo2PVpkrAkf094aDK
MwM73rRCbNHOX6LF/zAVa/nlSkJhcTwA81cV5UK0UP/8nnwI820mZwfDpCKceRTn
s2NoCNFuNycN29CYtim0i/lVXQ0k/q2oYn3dLsfUMFGPdh7MSGe/Ic3W1oZAO2ED
WpH5fSQYzgbyGv81L/heL15kPs7dlnFuBwSU/9mRhRqkVT5B6Ythrq4Q9Vckebz6
mf4JueJeKyuEyuXqe4JBbXP6Ys/KlZEk/940k4eCYjX0r3N5pcHOcifUKn9Mpf6v
ejbbAD2KfJYRB+MGQA2s0o1ZUbjL1eOJnIXdW13wRaOgfPbE23deSA9lJxkTvfpa
iRZ48WIthV4T5MmSRtpWIsoPksudwYBWfJdzIyjodIxVYeicm4KwvcjOWkst9ujw
COA5s2GQF0+DpE2yQRk21npB99t/cdpIW9SJoOg/4EdZ8CtJ5iyEoCy8ePc3ZJoR
dig4zgBpk2UUiPTy2Ft8jbBttia915/kF8VAbuwUmZZU4h+fAaRCn8bnIbCjJ0+J
sIOv0r+bds2ZfbWpUkSJapS7sp0tE5Rkmm+62rXKI0wBlPAkeaXZecqNeYzklFWQ
P0yHYNrY8NrQLaWRXMIbkCS7pu8yhoty5XFdZEXm04rIWrGbJyQABaQU9/Retbn1
M6doVRygALS0CFZgZH3ZNW8gGvVjCbs7Hh5vr8woGn7ABuXFtmF6gAjuh04v+hox
mfHrlgsNJPvU9LU324ag4voZhmgxmBbpspbVzXw4n7Paf38eVAk8p5trFQ326dsz
bB0tmKjd5t6wdXjVqbbAJDp6QAYrfjrHh+Jg9jWH5B1OhGEQZwbuOYq92ve/fils
VJistBcPer/sfouh78gyl4UJ9TjMPRU6SX/Achw23dxkd3bGWOaS5EBZB4XVvW/F
bwgsy/BK3IrKAL29ienWHVPQHOp9VJP2+9Nci0Pa4aO0JpAFoGHY55ZveiyBoAKN
XxfS/2V4yYmAAs5AJqaHSeTuIYOijate5hFwasRcSw4UxZYy74nXmrd6PplIT8V/
37lM4DtZqpmTgSjVX8odTb7xsMsVUEuW8291o3mQilWjbGmThPaKjVBWelm+70GO
iAnVPodFFOZohQTt/Zlp4ldxz/nthvrTsbRFY2JaJ7dd6VhNx3JcPH0zWAUpUWmz
iSIMca/V8D5cjJJTgTZsd7U5xR0Bqv7OPu+boGIF8m6c+pRIfAF6eJ7BxJOXbsXg
aYpuMe8MlPxFa3Uryk3rzx+ACX/S1DSaEiiN0PKhDyoCnzqsjWHhC2BLFTIIXgtw
M/M4wstoxORq4M+onX7wWKnLdlhH3+xV5eN3YXRmp55G0YGxWhWmMhPpn9zVHaTu
KzmwtdbkqgON4ClIke9WECT2gmlux9UcQugVVs0FvNI8mQJa6J+jy/eX1ZP3E6yd
39sVhC6NEjoIKUzcP7KEtUM4yOAMIPIz60sWVZrwdPLbtXe2SXMWl8sav2dZ+7UJ
PKMNhoNcZLPo7idKJDL86TiB4gRJ3YKlSkvmGl0EdKFEIrhZiQcZeHhieQoujm04
RjDoVyRCvYfi7XKQV5a9jeKw0Mje9w9+EBr2+Rbgx7+4mLmkJ+73yQK9gkAkjbqY
1iWyHno7cOaATu1OCDg5GkyznX9QtI2FR2hd5Kzcn+dCLfL3swPeIt1ZIRi8gYEp
cM+3mObHgja65nsvtl2dytUFYwTDdiBb10wj3WxMdK8Hvc+0LBfZMeq6syIRUtDN
Sv0QqV6hCdl0qfb4LF3GfaN55Y59gkx3kbQAMr9b70KBn9O/+hE8iFJoS2XIv6ZZ
Mb1dOyeMGzqdoejbi+OIspJE4Ds1U8pnPrxqhKqYW/yaOEvxMDPjsU4XoRrmGD9g
q2C64VRCsdngWZui2WQuOx0+rPyIaAwqt29gb6PhVPDdr69XPxy5pD5nb2tikY+F
aUn32u+7IhnbY8UDvw5lz+AMXt3RM3tlC6qAEQ55pItvgEFybsiKElyb3bqRCCCY
ysokBH9sdE4mwfyGCfMkyTJ6XtHnNtvEwLzj4Ne0QImtbWzo+PChC/bp9xi01U9h
s06qj+Q+2z1vryyadIg9mQU3i2hAvVx9IwVyeGFLFJspITrvHVcU4IdVJpWFFOW0
oZtnc2K0A6q5mw+6heWmU32rV8wzLWyJ6UAOVLnJWvOoF9WtJSibvQsJ2/GPUDpG
z8NWch6XtotGggeNRyj7wDp1PU6PxCbtDDigjjuf3coX2dwRskyWNbIgIKN0s8Op
5dhl3t2IUYAAS8HCYzIEADKRSoxKsWZcJAlvGvArzW20wRH2dsHU5w4nHTrNe9Qs
NgSxFaTrayEWjLDkjuUK11uF35Hgi7zhdmnpesf4xGkOK/7ifPBoZ/CklraBa1Ab
3X8pZBJ6JdoCORlqjE2waEbIHVcO98zo6NM5RALmAnlJir7N8JKVqOaO2KDPFTDW
xOCa2WIvYuduMsSjaSSoYQebgM5Rh3mDsuhXWyCPb6NLM8TCCHgHC96wQixRx493
0sOsUZGcNJ6xAm39uuKAh/GWiQJeEtIuU545E1RkK7SXa56ndchLqem/tpcoxYFf
DAJ6pYF5Wrf96BF3PzYq9dc8UCdgndfiqH4FzUoMKwMZMEOjo/0Cs+SbFkpng7H0
jipI7gusPgIZcWIxYfIXwU3HVfVVysO22zGNKaCQZvJAzJ8QQpiiciJhUpwKbrOR
vWkmJ4prMCQ+JBcqKSq9mIcjA5sGI7poQIc1ZLB2VEInFh4lZEP9TZtmt5+Dfy27
1ScBYcJLC2uMTsNWiL0tDg7b+V3KWoYNyIGnt4RIZxJ9RhGyiIiEkui1KQ0eFmt8
PSQHD4rDD+nmyMLjSyueOVJqgayj26D8BhxiDsIxJQLtqGCG5BAgU3CcDY77V2AX
ltglmHafu+6pQc6ilUwqeSwk+Nksd3neho+dp8eI0FspeNAkGvPjpjiDibJaR2nw
ArxN1pw2sGmOz++SkUSODatelH64LHk0UsR2CS0ZA0WNWG27Rk1qHRRqv0VQOvpU
vFx/uIA0i1ceg5r6BHXB27BC63/luZWlsOUaTHibWk31NN7up/dpEA6bq2dOZq7x
ikIHmGliru/UPmURs6LrhGb/a9061L7IKzOoLpXoSNxIbqjkm140SBOZk8tnfICe
VozPvk8xtt177nWJrFHeDSWh9BBO9WzmHBJ9dTVTVxcFPu0RO0b4WhtWNFoLTHcM
FUoeOoq9DKYGYFZAOD8EoNMeZ4vUpSAabKy+/PDhCB2z8Hd+A5nGppbha+P7wbAz
NCB0/dEzdw+axZ0ZaNQ/eH/XimVxeNV+Ueiy8fXRxiPiakyrm9msZc7ciWs82r9P
0Fcq/z78H4rmqLoLNeKd6KEMo0lJcTa6MNgyuq/XyqSmr2Vt/dWoalbeD2jTwNnH
R88Yb9t706G+DmN2lUB8/dV+wuEN0G075GRTTKRT5Mj1t5ZYX7fqtZoTF/Yl3V7n
5cUKrwtsenJ/BaseGDeANHL07QBB52FZ8ELFByRa7RfmHW0v/jkh3VxSUOdCtXWP
SgBUeK0rCaUptJ+VmSyffHjNTFDNGGPx0fy0IuLV802q7Xzsu997/8IZTOM2ZibN
SdgiLpoKWgROIcFN3UnZvunK6ZYNthj3oX4HFsX+3S3EK4O3puaH/ZLAdhkVNgpD
PG+MDd7tjL2DDzhNx7PWfCXwt3HjPtO4HUowp9/kPIhLtlPG3J73CFPySj7gXqsT
1IeIZWBmnFSBXs11tY9meqSddEYO2I2ztBt2LQP2YDa/tF6cnuc8ECRT1rylkb/0
GaG1hPF75CNfrjOm5SsUtJxjZ4HlkW3lb0RtuhhjOtdLNa+dVRuYlEI/1zi8h5pD
AlWmGS9jOQmDSoAUSyWsXVxMP4pLvSCkrWPyXhN7uvPXwVm27tDx5TAw8iU10qFR
nDT+1+U0pUTNhY4fr4AeDcKlYkfCrkX+q+uSErpCAJ8XqKq2qsDQ4lyxL8UqGOmT
/Q583ndnsncmy3E5ePVZLSFFdWCMXK+XWJ2UgXhG0uUEVyc37IZdd3F2bFnsfdy6
DcHewKo0sCvUjMeXV0TmOgCFpLcGKv51foNYw382MzRLRVLjEAKAqxZtsgHHO05C
cfOjs/l+vHRIzLBLX7rxwJiRn/To6iigeRwBaXGWpey2TPyTdLkGnhqly/ZulSCk
a5HXtFq76OGzwO5qs4w0/GITcy6bxJF2dlGxGj7iC2CTGU8UEtjh6E8ZopleLZR/
eHiw0dugpzQoxh/hd4gO4wi4fsng6dqG9IGxY+BHVX6cYIPv4QkHqw9z3uipavZP
g10NDxlJFjlzizjUWVUgdbpapSswlixzbAzsCMc+L6rN/yPZ93ULb50Dtq2m5VEZ
BsZAv4cuC1F/XL7mps/rb4cqP9q3VDr26tJYxxPCa6ehelMvQAmo5VC9tiCibPxv
ID+XKOvi+ECIkiJ0wmHlylTVst6XAiFPmJVDfQ8bDxwnRIJ0IU33yLdkC5HVYvgI
SOt+5DiPYyFAQVLhzbiT8j+tSfNU2Eri+u9mJxXd6L7wAXymp+avHE2FDxAazdD3
mWCiHtlcJfuDraDomMmANsJEif1BhxxCXb86a0NwDh6uiRnQ4y8K3jtpxJNUxt/L
+ehezpkRwG1H/3mjZML2WA128UpMY45UUyvjK2LOkhQYkB5FSxmk7DXjpufWzJJ5
bPOgxOtieQ5eyCzVJ1NnCIYbxDggaBzJpvNvmcKiCBIfGxtFMQkbIve7v4UgPROl
ZT6l8r1uPsvqJZH0vHvut/Uw3cLVmqFdC8yFjcy2FJP0tFHs+up7ea/uOAUcasrg
D3t/f4hk4jvJ91R2f7ZBuV+VrF6woGZdWu+t95BmkSSnZfUHY1hvZbOz1AyglReK
ukOCSyKG4kOe7IF8I766QccompAxwGj/3LVTBl6syN2Q68LJQC0c3wXbrJk8C24Y
VrR8GhSTdJIc2SuopBP3xzmMRNXqLtAqzI8ZSWQtqVpX0EoES2QGkP9KyhF87rgs
nZy4eXKvWq/HDI12ceSt1JuHoP/nXCy3dvPBM6axne86CzavYWqJfo9X8KqpyUKW
rRoZXT5TCwrm6xUmw/Btt8wMJHI9qMobrFF0eOgj6zv6sBRp5vuVOZAA+weNC+ng
UsmuuSzQmRpqp2A7Sg3ZviBlYSChW8KIGVjw2Yx9MY3S1eueRXh0FkYO41A4Bdwl
eYB0Wx2shTJ1dg21MvEkjIPsyVjg0q+EICCVyi0CEkxGYwqvr0ei95i8dm0DiI5U
dyH/t52eR1wHRYSQ1srarnLdPkpua2t5D4MgzcEJpP0nsoZQBJnq5dDG98e0Qq5D
vSZQnvCbLzl+enfBDuUANhhZZZ1/awk47UH8yFLq6OcScf6EhcLBVBXMGq79ppHi
iZGDDgv4QBGabt1Y3GtZSkft/oJx4Tdtc0EGM5rqfncKJj7pHYr7hTAkzNFwDkkp
XmCiL0oQIf7eX27bxfukIptXn7wrRkKFPVIJXAxPc3ib3nujSfimGqF9Gv0fbXj6
J4VB5hWflJrem85pCJLT+dks2Y8EAuKwApPUJDm4aydI24qXkySq4zKM2V+Rde0K
iKyMMgnblbNwUYVnSqoHCpc6FFRwgJz9m1ZA1cypQHG85dd92BxSzmGi3J06iBLs
0GXyfPKMsZSrGFxXnldxJANc/GbtaRXPJqOq/v3BFr/H2EKJZNzIfS3wCgbqScXs
eXWf4Io/5nbgxoO2XFxCvlso0gJhg1UG/H0VobTlsAXORAyeb2x3MhhSpljcCk5U
jXiQczHn3AIee/rkh2vjUvqD3Cs4Vd2br5dTJmaN6JGGO5LR4WxCc1y52Nkszo4B
OK3ASuL7TbkCbs2uX+eQy2NXQdPBllAUOLanfrA9r/Ryw8WLT0rjX90+KGjyDmkR
i95/S3yXGl3nh2M/1RigmAgt5NqVXshuNkdXsMJy5/pU+Tapo2fLDSoMm01DKNgY
6VH9Zj0+W0xrFo7VWEdomjRwxsYC5FUfk2LvPjPegNhWN+o51Xcl1+QkrHUIoJ6l
S06K/j5h+OnApP0B7P2qbQA5bvjvqivz0SdGyl1xSh2thwe3yxKAZNWpi7Snx0Ww
7ZQC1BFqa2Ru2CPZpkSv8bnlq9QtOVqjsZjQ7r9iTo9J3uK2cgwwbQkhTootliz3
OkdLyfE2bcsoB2KRitv5wOcprJQMVfmeCTPf+uT19tzJ5b1+K8/v4BTIBvqjm+fH
mI2hk9gbAfM9U6zPZxoXR+BwngV0AE/uWfz4tNuHRpAehjiRIxp0iu7XvD5bUZU7
QvFd4ypZxdi6h1yUbts8mnuM8ZBVAlmQf/G/NVQQol79ozEQewBOw5SGQ6hWvxIc
qEEzSz0w6x/2toUOxhZCWC8eDeayE/xcC4PM584ZHvFeWLwiC3rD+RamTCmMhquM
uDsp5a3HLJnlE1gtCkjUG279JlNRL3+36ej1+Lf8Gm+3dN8VZDr+xRXKe3RtKroj
eyQxHVYU7ZJ3Z8EXDQVSajktlrH9W/RLJmuOf9P8v2fFI6ovqHnyxr0CKUF3ifFm
fPk2avP5b9TAVdYpi37qbtS7aiNlJNrWXqFSdw9yZX3ph0MDlWdJEtfZxD1dVxej
+qm3Qbol7PkrCaJoJ4nM6o8/AD7zP0Pu3oWjz67CV0E9Ybty0iXYuC59A3OjCL1w
du/RZdI29JlDGh3kgcDTLfRCcotCvuZKBDaXeBFUVcx8YTfoUoskVxmQ3w/yNB9j
GUA6TAQG3PonlMDsz1mQpVZKoz7zRQ4m3Px5GT3Jsdp/v+QFuq336Jyb8lU9OOMb
juYVGG+IMl3ykLnFhZdGXfSRedVLcafILEV2qvKgJqn/DGENsl2rKiwjeUcQo6uf
dRlXM+rYny7P7dMRLp80A3wovzhgqrBtycEmnipVo8xvzcFOZTqZvAUFK/DJ9LE1
KRVntn944/lymtC11lyj1xqDU/8/9s6Pa2sU6mtSROp/jB5LeaZKO51PN5edDKeV
b2ZJ23nT4KPQGLbJxTjtZMEtaePzbe9P4olfJ/kj3sScJ0M40XbrOvAYF7+TMkrl
L3G8O2XJUXSrMzdqZyHFJRU8D9HmNeXgEQhGplHWKItKAjYoeRJjpiSGsRc6tvv8
7/xCfGa5fshfRfxp+ZqQhE0nYI3yWk4SklS9eEQY6/Q8NImmWgokXHAuV7oZKwbk
/iXwjZob4IifSUKxHaq64DgvKIeswe9nXfcGuAdQpKGiirxWCgg7sR6fhqTYenNS
bZ6wyHx+0kwKrdpUn95zuWa/33UvRV83FgyBX6M1xPrl0xjQC3VRRyY/v3m9Nwru
/iRHS8ls7vOhhCdwmu4uxcuPfm7rGbCXTu98AvjWGJsD8neR2dual9GCh4F4K7eJ
PSLNxxaKGZcT8GiptixdgGXV2V9iCJf/ZeJACeHPfWr0vEURTfULAqflqw9S1pWN
4jjlZiMcvnMAeM+wu0+CwmyBAOl/zQGVcPPS8M/Lk6u1LWOHMedNDZaSrhrTtJJW
tY7alt2x8CUZIZxGhNSbaLAl9OdEE95XEmq423UBsqx9wK97gjI75b1qzwhdUvIg
pFs+VjFreNvaP7y4/29mJVXw4oSh0lstH6NEfEpkCwxFZYFf8v7S+Ta6fYS+4lVi
qmOQC9Q8FJpNMvHGih/ZgxUxDPDiYCRttxOX0I+0X4oy4QFxh3HUtwX5jy9Azv7P
pQV4/G02wGziiDAl0vDaWYaBZJvsVcjNaJL+8uqYxvXNZrWjPv+Ler+/0F3M2gZC
QoyXx2dmKunqDP4HdaJIg1shXxJvcYXjVicqtU/LzU40UGMSEHo+lP6U8OsR9S+E
Ps7d1yEOWEKWqiXRvtBAm7GHvGpKFMKChr0Vcd2GvxsmoHd4n4I4DPEIP+UgDGNN
h+j87vHAp/Uo15vD8GT2GFDhLY65yfFyPwps2tO4ADEDVdWC3X4JThful/YALtIB
5MF2MoItAlKl9QYRrqialCvDRX9eehTi+UMkNpvD3DJHm08xsV41hqZOR+0ry8uJ
gVAqRTHjB1P8qMXzI8ttFDzQJAl0ff6AzMgKw1zRPeqnrFjtFq6a95bUkNMsh7iE
RKDIFroK13Xr7WcTM0HhtBvy5vasN0fx+pP1VJayJR5U8NtiTyAVHCPPx0q35+GR
HfWf1iwnnT1a+BHz+S+0aoMZJK75Os9+JSpy2E+sKAmE4N6JGRjr9U772h5tggls
9Eks/wgtvUN0OYNt+1fzW51pEy/hACnE8DFS9FMQiiXDkwJXFE7z/5+N6aVg8Ry4
bNUgjQz/SQJaFenVX62g6uXzKXT8swzv2QE1xPbRrY/JwPhxtWdyJErYLQ4qBgKq
AF+4ZTTHqThw/ojYgk94PO04mOH3c5x4ubzU+DnBZxXmHvBZDGIy8+GEYo1v1PA8
WaQkxH2AUFkMp3crNfuAMXaaAV3VYL4sAyI5yZXr63blidQKr6uK8H+bnDkckfml
FETxnHpniMGHsypHLlESjR7vlWd6wouQmZg6n7HR1COqq+R/J1yY7vtEsZuAuQVI
Y6Y/ooQPtojSCXpI7fl5n9BfB+D1ClZbtxEUIoYgIy2m7zYjfMfwfPN+fG3twV0g
W2wexSJM02mcHrXazdE4cFl55R8AoxiCKk8jsUTkoLEnws3GQjj7xjWIJFseP3gm
D9BBL//JBajJhx3ICHzmA7L2b1wipy0GhSoN0mndyjGaR6bWz6Ig2x+pSHnRug4N
dTbVpKTZWx4hdrvh22vhCC1ZCPDw7ByVIWIeLpKIPAVWEBUMolBAOQGFtIjlO4Gd
CUtMEO9b4KZkISx/WqB8XsSVsCB9eBgxfB5My8j287l6L15KvJgEtEVcyXoQJZv4
ssY6mxA894puhcCBto6T5Ht/jLVSYYdJZ3bmT0HVv56+Eg3o2lco+mxB3JlrJ1hw
l0FORpRmVzV/noIhgM4QgiLxrUUtvXB9k/yacJggA++Up0ffSjRlA1JQ8FvBeotb
88m4T08FImdmvtPJRCR2fTDP/6SxqCZceVYkJVhMGlSR96Weu+U+nVvkpLiCSYMQ
zFsWP36XqY4vEofqDbhXaxGxNmG7ypVHbciD5hy3aWCBsthnbSAOtnJLyq9cy7x4
ncfyB9f+MtwwEwITZjsBqrrOndRNVgx9rvo0h9sNPPKo+eSfa0PYIRf01VjTnYJX
qKmLeBarkV7qfUJRaVkvcI7uwfd2955jfZeZPOBqo2njqt/J+NV/oxdF79cb2GNS
qClV6dPRS6Xk3QJ7usyvcM+xJEA6WOvSuWgcX9qY7dJPn+c+FS76GcQz7QPrHY3v
s1nyP+tdkAJuFqN+ru7/2kg0J9m+oH7ybUxTT78Whn9dkmGd7alPpAmj0DLJ8VOS
Hyj5umJAV7ix6DOi5VETLGXJa4wsSE7TjQtP592tRcGgcjw7xyChGWK7cQhO5fCT
f1Sdb5GmbePg7osXAq7pxSXXeC1VkEz/nJkWzGp+FhrkAApCdpYDWMc9lY8zDq3Z
bFVZQj/ciW17Ws4U/z7ivvYkvE288zAww+L2RE/eZPwRhmGQfp9NM0nKQLMAx8aO
/HHbplPCqJ8+SlQhoZObQyi4Ywz/rpmbc+ZiSLnhLYtulF8OvqKnBHMNRTGuYCww
qnoQO8HLmBh9CYXoHli9UbFO0x3XA5UMbeSTO6dNWxScsFU53WWX/+35CRX+OXjJ
939H/PlstP6B2ZH2NIQpeIxI0iR8WyXIMwdkDC0KxetPuGQ+NyNnAaWtu7zlF4zb
x+7fyMiumXo2DhL84jCdrE9ZvZEgVgaWNIUdhHIhbd2NsBSaM/SjAvapR5bpvNfm
4V2BgKhJDqjAdsDYtaYgIgGsfB3a2x7m1VX50TNYg0HOORR4hUAYyS6u8TOejRRB
T5Jbx/cAN2g6UmYNdgm/jTMsd3ot+kPEoFbq8j3q0QZj6D9wbo6Z2OaGTjcQLUnL
2zBs/PCnb5cmEz7fEaYHBhgE3mIlXwLyalVSYm/KC9TPg25VkUbzdzrDdKgUTwB1
bDFI4r7ys0tK8r9kuxtIC22OUt5QRo+U5wEVWQ7AKqTpDEnQcEFRYydWSOzSodf5
0kvIfV+Mi+i5//u2JXdqmS0EzF6eQCUhX6AQVI0b63VPNsrsYJ6oNGlE1yQNS+iv
tBm1vIIaLJFy8qeNlLjcuNU8y+k1Gc0ZSL4RJMbqyY97wNrFXyRs2oWYTQEmSC5I
tzrw9L5hXAkDLRtrQHPIbwcW06UwvcMiApv4NHu/ecEcPOPZtPZ4185im+RN0fgU
i1zgUgqLp3E8uHzHt/1JVqYr7HN9cliMiKY9OiNEsPw3nAUVsYEoIpOF4J2ghkQn
OwoSMVdKch3QDOvIgQxBfOjYsF+n0wp9EyvRlwFtLMvrB6DaUgbpFcBBGa/gk4oj
K7MbkpePylGcBhCMQdEGc/AmIiG4CTB8Dxe9SVJPS67Ndv6nMY+RpAL14NaA0TJE
DVNVeAyvr+aofXPFJjHldPDrHqyJgGEwXTTDEzn0P1iOzGIianqcgB9oKjdjj3aw
7tNMM8V9zmiUdI2XOcs08RElCGtZJ+QGyNE27UMAdS5Erde0CxnZbaOGUxzQMoY8
AwhsTK7+yl/tTIPjNdO2x0KnMJb7ap9f9oLKclTyOyHZ77WUxQamcXjsl8+NBS2D
3IBP/6xaqI9vifqIPbbw1tYgxrianwaNuYjylZ+IpDpli+2k5XypaiHZcmlU5ZSq
8cK8rNCzrdQwisgmSLp32dK9DH+OUF3P+vcc9554pQ+03vKEbykdR5wS0CP13YDx
k2BopQhJE6amgR1TmWTLUlc8dkHUmCZDd4FJyCXKPEjOum1yxLksk8E4H3JLy5uT
jLylfqsPR5wEXly/ro7gJyY2ApLulkWQ+klEVx47Od3MSdlG0yM8IKotm5TwCREN
xY1B8yA9N1886uBL5pklzEqXPQLAjcG4EZfq766aPTaWH02vga2yok1hDxRqJUj+
ij++4oR7ylYBGbfezqZVX35h0TFR14wXD6afWZrzEDAs0x7LB+ZLuzN4Q66PgjF2
PenOzvd01HBRlCZ28ZJidqKQ3/l+pyNPogABlA+/ryAChmdNRASFbl+ad5n8g0c+
4Rh5Hm/kq+X4dWZt2WS1RAeT3xxbKcYQUkZq1XzjW9wLqOv13ZoUuyLISC7Q/rEu
3vBzO8w/j5sDksYgGNhv/XLYpIa4+Rs5q7aaWMwXzJuErBXjgS5IqeDyNO2K4hJa
vjXgx0IAny7wiI8DL39uzmAnVFbiq+b+qQcMXEbHys/fBuFDi/8plq+5fUOXqnqZ
oKnKRmsQVuF7LDPEQ1KWdclhbUdNMU+aQzDiQJ4E7clMAHreezQHU27pRsI5kFK3
9REBed2goTUblJW1pukeUeLtK4Sqsm3GY1OyUT+dOYt/uJYpZ8BbvVLBt3enGb6m
5FwW37GaTK/SHR0ftlaQyfSA5Zth8sFAENaSHcREFanitkqF7/iDdXl2azqYD1kX
sC7KkmWpecFR2qj3ugpAKuWmarS9JN/t48ODddveNrppfj6DhxS6LP4S5zJUjkvs
0Ul+wOCy2XnqN744mnrJ1qiwtfVGkrPL/n23jqBP2CKUyoxKxYam9Xcj74h+KMjT
XkcAce3ObdRnptjcDPAm4YOa0YXZXHHYOjMwqOGrNZ9/iEFWxr2mReQ/evvITZfL
wmH+MWZ75GgP0cZEcIXW6eVHStnDBlapriAzhWSiP5ftuGTo1TPosatxVeLWh1UP
2LClbxDKyWSC7sIU21Fhb1F5Opf4vz1ba+njLhVqDU8REkEtLzKK2AE3It1dtFAz
CgghtQ9VrQVLEqvaOrhp61uo8OnYrPtkqydB6ghFTTXR5Nz5el1VHlPkXbpRMAyd
HWdTHsuG7vEbmKO335jWZCUo/YaoVoeSK78O2Vn3gK0iMltuh0aXlSvsEnDGXQnE
kbK52Llw52pN1qzmzk0roNPtoDRsRzohbLMtIXCax2pRwgMGpzhkFgN4MOkO1hKk
QZHgqH/G08I4hnq24/GyWeEFjP52pFTLvonpm/F51Cy+ONc0DhMDHCO3RyrlmI0l
j35jo7tvIDsgmLGNO5EOe4m6r8CK7m1TfOMwHa0ed8EchmtdmommGPmqrvhG+u7n
K3Tsa8LH1tSBduZX8n1+oW3MFtcqhTnkUEchcRWzWmtbayds0plH3+QiZ23KyOEZ
RbRkfMf7aueLkGUpDqmUX2kCIaDJqdZ9INvYEWwLCCggxzBpNU8AY+j8cCrNBVq8
67GuBg4jhETq/6vq20FmmqRw93XCEbB/p86NCNO3KKxNDtvu1PlEN/V7FvxO9/1V
1EVbdOAqKtrjaHGf/YgkGi2RF4vH3GCkzgvQfuQ0XT24Yug3AfsYvBT6ZT+nbixr
k+xPWyrtKtxq0g4JvFbuQWzwXcOqi+Q1VuCkUcMrKHKsk4E37LfJx1Prv3gBpKGS
oJHgX5M2ihzg7vrGw2AevGucgab9XZqBueV5tDw8wts75e/hpB06qLLqAOS5+Ui+
ofGfAKYP95Hcb4Zq3dfsH+naPeelX1PMxeSMrXdDCDRH/1tIFBdf1vZupPpfoEda
vQ9R8f7buSCELlNbcDfQLDSc4870Qzs6SV/6PV2ZLM7xTVuVS0+OQPJPGpchg+jk
ppo7v6tQGQHzj86XigNJXM6cQnjoX6ILnXJIflIY5TPrDGN6uZRRlpq+F6tqdwCm
1niFW9z/QRdvnYDLq2fuq+FzQ6tdbiv/1kDnp6TO5zLdVuMQVzq7e75025/KSPSC
y3vgCK4sLLWmnN6GTEjDbfph5XzSriestPz7QFA6sU6KpwZaF1lTSPJYcIMRNQGh
YuWz1OV81clgRYSMf4UDnofUI0NbhWkWGc/fue2OmObaAsoDVld+75ga1f1fsZ7M
IkJ66Dq61J08oHmlohuCzStZPEQ9+injX0XaUvnzVBkP38scu60b7tg73GT2hO8h
1q+oJxFTjB3xBxW6pN106kHg+tdlWzU8cmLcPc+WapTa78uR+R56pBecF4oxbet1
gyzmbj3mk492UvC2g8g9vQuncTf84gmop/bedcactljUGcMdWIh/ka+5cjC+2p8P
MzuQPmiejxEiezVcglnfx/BatyGKPkBxEKrpywKbB7bV+yd/x58LOgjM238AMdo0
9CMvBSAgyfu67ZTSxcMtxTYsTroq/e5t6Azoo1+uSsUhiH0MvF6AQ/G6B9q0EfD/
LK5kgBR/eyOiilGNuz8aLmysKtoDhzgOYsVaO8njlRrrkr0zCk/98UolwLbF1RrE
C8SYhVPyJ4gWPfiz9VXp10lLgp4sQgOCFaeIkBeOk1ADAT4xXA/6mMBWaEcGc+Le
CYiaTcNlKXfwRdpVhxw/msrYRVyS+iL91/qHObLAOPqSPgWs9BIqIUokG/Uio/XQ
o0mpDAL52WfxLFy9jFaxu/HWy6gUfrvLUeQK/3Jo1HWzxPap33dzla61jwA2FDVT
L4BIdihPwDM35nGVd5if0TZw9THIvIErrIRZp9pWJbx/kZDnO9F2vwdWF6ZUIwWL
9tS0Wf+fyJ7jvopNeq+8iwyGJuXzRB+t5gTNn6N53BPkbesqxAVbbAfZdt5JpNKp
MQcUy65ug7AnH5g8D3mFyHk3MKPSw+eyjkkrjkzdT9r/49Eiex6pgyq3dXuNuSte
LGsvqwiK/2Sjns1VyEvBTWQcW1d/jHWBx7hzPfHA6krIBw5NwGHWMREJmCa6TbC4
YwZH/YI6jxSRRa/CTKXH7mI3ZRn2VlHzoDdEwTC20rs7l6zmpGJZKJWdbsv+rJDz
K8UNfJRtGtZe/dCZIZiulZBRY6k/tvtgi+tTcXF11DUW+XgiltrxenVGY+1UvJI1
IaFo7d/5mmp4OhVdGTUwG+yINqmXg7tfkFjygdwq04AZ38okoyzdaYnS58SH0vhB
1jLzrX/jq715C4uHy5uJpZinVECI5peCE7k0weM6h6Tcb25brL3bLKy30+8eW2RQ
9d5tiRBggIQgh1oChVKqcQbxB1xo+fX7uhPcxYtBrs382AXnCOBb0r7OG3fYlECF
mY+6gdOijA5z7RORzzaRMcIL+gmpaPHJt4l7/p7oI8Y8fcjMdXPuD7rpD064vc8Q
iV4gHiplRfB9Q2qDl/xSmLQMa3uMjEaF4I5bV55LFyhcf+0mFNEt1d3k6m1Qz3CN
KBNT8Pa7/eqLaUW9yfRvPiadOZPMIOLBbHryCGf7O5OC2QLaoFkGeMWEC6tMGkOT
SmOLIeDEUy7hpMzYOlGtInc3KnXZMSF1SJObrTkPOekmMstpZzJ4OCtkOvTT7wwm
V2vr5IzD66i2oshjPtP3Hl5h6CQbuvt1Z5GDbaJiJiXrBn8Kl/da+6AV9NWcPEma
QyH2h0IJwrIYlF8FqW+50YlcsnJQotpQ9Ha8O8yrP9RTA8GOVw2GpHqJzxUUsHZ7
wuzjkspXECs1rjxdgQ6Yf3hHd6yb2QRL/F02JrALo72d7hHiKmudXRIaUip1yhmC
QZuNLywZFZ1GoG3m3qXp7eDJJkqzyc78YyuZwJaPpNkH4/hIVWp2E538xCbiYD4R
qLNT2ATo5nPC4yiRMYXZqVteD1qYoVUK+PqbV13Pci5iZhMdSL2ktOnPPk+M2oxT
g27fSLWYK9o/UwCxQABl1vk42mEOZl9nChFnVeptXi/bKLWeu/tqGlLGZZCdBn5x
+GqLT/KuhBpdZPCjtfn5+mBnI46hB12UP0iAtqcCIqrRxabv4tOGi6Wmx5xtBhUv
hDa31+PO946Dw3aKJXmh5Mm7PCFsEtcoua+iL/xf+iKRP6T+Wfbd3WVT8YD8ub0C
i+t0iqBg+NBCIe6KlcyfDbe12/yiE6aQQsXD4vgE5sk9qUGJ0ckVPJpX0eSx+AaP
Ww8IB3+IqwDmWenUbF0T4WSfAgc7vKmnwvtIdUEQvpdKhJ+FEIHaUpEEO3EwX7in
mcRg7+WWOfaLfbp94Ew0VazJ+KLfruLBTAC8QWjMRiOAY+9COiYCskss+N8vr6x5
kTtNivDQXM96KJhGKrzHXcGL5h1MhcfmLgkxCG0QY19VIy1ru49jjqhh2xJ8mYQh
0bcSwNE5S+2RS+odZRZRLgvBRzQ7Ev6kYYFvY0bzst8j/F2+d183JVVsvL6x45BB
C/jMRzL886qy9vDPmnkSOlmp7R8U/APYGUOBTEEqXZ6r2ccu6XXB4gvGUHpRWL3x
8QJp4tQvtTu0uYpriBO46LH5mdV/WjUXwBAx7xaHDxtbdsT/6Xh3sjJyg9r3Zys2
pEyd1Jf5b/RZIejvWtlMoNXOIvd4S2xaaYJYXNfPGPNZnSi6pJ10nQ4URHUcV3RL
+Rp1OE8ri7LjapAYhWOR3J41jpT2Q9xxDoJE5ysCcUfWR+GUpdDFBa0wa2TuRQFA
ekkpFM4iDtL0FJfY0yggpC3jtwgHsKip7MhsSYlcDAMIl+93pdh8PmnVlj1Zbid7
BCoRlSkOm/7ryj4JKX749y74pC6La4chP54XPHkx16cPwxEbyY/ohmFvzNKXyKAt
/96WhOeQe6cVN6EMHKHb6Db4rA/eLuQ2Ew1bTP0mowSzbO/mZiS6L8nxzMidhp0z
O3kYGQ4GHXPCDz0+lMXXxpVsEe38mUedVfvgnFIz89glCVyrqRtbaKJT1IbOzuZ6
v1EcoDEofETHVrj8OsQOPoaYOUodYBoXQ77+i7CLV/GglwrF9Z+Kr9B9bpITDaVj
6hkJiyV1T89Y/W3srW9FuCbcHER98pWF3u0eSaIEzYhh47qIk0n+7wMhxeLnAgpr
USqRhIzlSMdnhvsge3BN8auMwfTrJFg5kWeUSoplljM9YMNfic4+njHt+vu/JHah
lU+sBHZp5pwmAkBXZ/cRn08gIijib4fPSPmsfcYCqr5jvTnFTWybwZn0KHIsg9NE
GVYl4We8CCGtGD6T1IHza1AYuBSLmHjuNPmO7LwwJY3YI3LIF0TCkS8jGN64jQ/T
uR/Hlmp9zlPo2SV2CmCwyYZa1Pwn0nLFPw+alUx4BBQ2kxfBKn7JyFdraFnfzja5
YFX+RjBmMPMACvnymej01R5E5lfSFE8UzoAcN5zh4zMHsS85EsORo8OeloES3/FT
QAllPM3l5Lg1rAOoOUKmtvid/6aRExJrAgeBoImN4iFDCLkL45ph0M37ayVot8vH
+/E2skGmfFXBMHSWUoydlqheBMXs2piNmBrISLt0AXJdrp9V9/V3COrvJTw+uWF9
2J6QGcGLI7ICg21KRC0W6nkkcw+oxtetiAEYzM5O3D3HCKPSarg/8uBc5FX+vZm0
Anr98D+G6BDZ2hx0Z2G4ZNUii/uSnOswC3rNOtcYjzQaXJCTGMX7PsGqCmIacFhE
K1cJTq7bG+lAWdH2NWVVuG4iAnLHqQMweqgCR+DJHj0NKNe2kaEnjSGgOo+vEZZT
qviqNu8OqwoseLvIfKikX1eLz9v2lvNIQtJDnuy/WT7M8vS6aTYNoeCitxY1SQim
D3mNSbnDZTme/A3rAbMj4XJPVSHFAmeFFmPWjSkemAst59B3bCR8hMKuVlAiJwBR
Y/jwTUUVC6aEfpBZaY4/LHfAZgN6+pPkTv+ByMDt5DOMPi7ZthzTenuRoKrXPhIP
/9bv1mubGxB6VU4oOwE3hY1gAMjytV/U+MmCOwUbVfjUdbWTz8lMJKrjqkzJwt2Q
qjhkb3JJfBVTMuqFd9unPsRYdJVq3Gq0R8Hh3u51CPJOlIY/lzLFkeBdFDxx3g2W
mXpU+c2vxTw2Zu4K2zCK1O9KMIkK2mvCPCXDpUEvcOp+Bi8M44cRn2gNnS0yu8NY
mjPGuWUjW47ukXanWp3DPWp+xvqi5472ccNsYaN3VdTT8yqdRA2dgg7f8L+cxAfV
l2AvPFO6HmKzRdikogtBweUDF4yTuR5LDkLNZuOKBYhfshB+hFwTlJ4PF5afy6R8
M8aCmP/+Dc2DednGvzLcZvHta1rV4UlGiYT205Z8+M6lrm5XIz5Um0skVI27zBBR
KOGk1KvS0dHamCpcWnjeEcSyxZa41oGZKxfhlFap/IA9ABd9YqEH9jIBVorTjjr3
V+COs6XwJH/rBn9s9cUKm4iYJ/YAxYwWvBNvapd8qlGSsY6G2xC8F2MYpq9zUHMr
yQLeNUFo9ahBx1NGdvCtet2xq3jfGADBMLHYWeC0iMMLqO5B25WJihgkQyK0CLvK
h4kg5SAhIzi4aT5yciU7ZQafGpBztCLy+DwAP4KC/y+BY2xsSnYQT4clhsXzCaA0
6yM7WGT7FAgWHVgnmCeMetd7hs8w/Gr/Ysx6xsmRO7bsZYzoq7Beh3qnMTqrp78P
6Xulj24ySB4Msft5EJL0Bg1fG+7g9U/Sc6mTWLu34VUUJjsjYiiIevgiucCgZUjO
uyE2ry3/+LvS/U/eCaaZaW1p7K/FzGgE454ur7GQ7SuXYKq4++rV7xWAWFKMABnp
bsGYmER6q0raLgHMSDPHykfjlkdT//hI3hh/4jUQgw+NZkzefvU3gO5DSWZheW5H
ovzJPMeRg5ahrSTPcGIA28Eb2WcDfnHFAZc+/03wzec1NEuMLqjxX/naD9h8gv+C
LpmnUSDIiBxTXGNUj9lgJ8WZGEmNB97jQ2R6R189ppWd5KXiZSrF+b3WPSo0CdAm
pfM0qdnu6es2SIXopKtz7WbmiY1KDp2jONg9r3qFQ/PyzXBWQ06F2KUKVhElUEir
O01g+AT04E5E1VJsr8hWtR3ujDVHvbtagDlvIKL/YZOoYcJGmtnxdOhPoZh3eNy9
hkg0qxQKDVOANVPQutugIYTBH426q6SLMIhY/wP8wFBmQyEeAIT7jP72s55quKzq
Jhmexdz/CBJt4Hf4sTesFyn3mCJVV4GPXyAi3wYp7zVQdFHzygElr6xIbG06s5Cx
NVHH1AbQ79js4A+2a3DD5baRMS5wOOyTBsJKBV0S5tqZ/7A4AueYl2LbruuUpyHL
C9M9HsuSDhhfA6tC5NYolbKS/U2SxrVF/M+1ZxCsqh7OpzhiJBuJfUr9rpYAanm5
Gm+k73dWImckLaKuc5phnMMKMFGU/gGByWDs9toA8XvNa8oYplDCbiSif5L1k0sf
oKA/3S1Kd+K8JN1ut8RIO9Lzzl65uoRkNCqMjAEefLpZB7OR6nAzIo67+RIK/3Tq
ecewv5OaWXLAFEiBkFwWDnompd6SSSIaLUv61S7iy0DASw3770x6A9WrN0p9DmfC
H/GjnpPPFTCazODsAExM2P4rEohI4QErPUB2kamp+J0qM2p4ALUXNcMLUEsYrP4Y
4CgE/fjPNxA5PGUrIogcBf/6OunQ3zp+12Py33bruAgDkWQQXsEIm+NdnZ3nChKy
PuzSjE55z526tS6Kq6OVu1OnqzNnBOR0/NMfftIPG0WNpJ/7sz+geWuM+n2Ii+rQ
9r4lfb0DFZ96H1RV4vUpuvHugjMw6MSi6eIdKh1Rjp1fpRxOJsia1c6deGMnpEJ4
U869n3L20YMuJd2nkxY8JaLPuo8RnQY1voRai5BgNwmoycO5Gx75ckzH8Tse/giz
MeBae2WCzrNVl+DVfkhps4tacaQlIfkRbHERrNpO1sjWyEPRJl587xUWo7mzFGCr
X5qrFY2ETuZ79cR5reVozqQFRk/gQgSxK9NNPaR7fp4HMN0oyj2k4JOEg09hqizw
oar7JOq5uRQDbgejVOOG4ExjNjWKP6d6p6zTjvFmP745l9gTlj4vCmVNuxx7HKot
TKtASvvld3jMKr3ptpfpVs7XbVbBI1JrIZ73K7BkAfzeRhxOKa1QdFGqxcE0a8Go
bPvm0QNWvSrTHAuDzwvmKoLNLWqd+dNmxKuPtJ+KyH6vgy46uJydh7x0TNoPSkgT
1SmqcYmmh3RGOqpBKMkq8r2K+px62T1QSSldVfjtsQXrA1H+SM0aruYo8XlBGhZu
dGyboKosv938JbZ9an7KLMKqYIImgFQPYEKgEnRF8nK6tzLNbh8eqvL0boFCcpxb
SIz34jlJ9KylYXUDvbSkNJBY0BV/Xxv/epe58RZErGLzt/hojaO3pw3gu3rTzYvu
SOZTcHOQlkMiujDffs/eMqwKNYeMj6vDQiGJRwAiS8KaV0AbE2SK43htOCbQItgx
M4QXlOp6w9qaYuaNcomwll8j8QXmRE663qr1SA84a5xcKUB+R/XbP+aeh8dYLNC5
vzXnnCiT9LaGjdcB+TWHsJ9ovS5IflMkdwkLSD/RuLVIG1yayrWBKFoppVE6lnqL
D3QBMVFDmsErJlUEJNZkNX+RrndeOnpeSV+7kY0Uf67JLU7QUbhcmXu7YnGSSyl0
1BLq4R2MmmD0IQRYob570WE+kARFYz9fgN74/sOoGWbtfg3wxHqO/4omrS4jJb4L
dzZ6IkunNy7E7f/OvsxjrJS3ICLDjZmGp0MbpklSiwXOnaBgXcDE3Yc4YU4cpDer
p0LXhpfoLsbbeuFqwFhnbdZQtjU8ssUSFTpV0wFHr141TiMNX8FoSwg+PZEkvYi8
HM3Hb4E5iFdRGkSaKtq88Aflt+eZ5M6zX2JRUc5qIlAw4QwpsZ0us2ypheGQOYWp
fkl5YttTU8rmjFF2memowpXDm7r4gurJmjQ5i8ijxhLSxZL3gB6+fMFjkSTzGRly
aIQSXSxnCPljqO6UwI5NxOafQo4yBEWwo/vcszlg4nDgXxsMCB+khN5zzTaBE5Z5
1FmG8gOww8CjaEe65/JntkFghoB4MyskuJyby6SOEfDranMzD6RZJmmQwZziS0ZT
3slobXu+mK7eIXjV/plrlXKUBy7DU1UosLM5atGuvGAIvk7qFFctAflSy/an7CcI
BJtzQk/8XUnGTp+2eAbA4x0bhzvet+DJH6ug7q7XttenZqALVDeX6V28DqWvfRVh
wYDU5YKEWhk8Wg8iXrzRlpKHIjkpeeMgjldzyfpSt7xIx9gq0C10CTX3xFkRzWDI
QKGG7p2ssFRZWJTZX9rVQT9/cVpjz/irWyeUk1sL9LT3X0T9mwydt3ptarbyyrkS
pSARxHlga1tYt1qUP1Hp37xmGGUnMcG50zm1/z6G+13PDbC7Jp7humWJptYgCXJt
Q7txb0Vjm3FGegmgjD5J+jPcnsSJ+Z7hjfynE97o/BMeqf32b3piCT1AqM7LZU5a
OyH8kEyk6RlXQL7XDAG2qWXxSmdQdo7JyjgajV1uUp5LJ/3Un3zb3zDu+HARe9JF
CKEQDBZxxAmVTaO8WYTMjezJtPR3Ou03LSc5bUOEDp3h5coDxShB7ds4YDZH9GrB
8u3oISL1ZGuFqqbR4lLDjlxSo/RmLWT5dGPtz01swCGEKZve48DL+en7gSGwmPV4
0m7lzOyPQVuz9fn+qoH2BtuqzKkssst8I8Xwib/PSnOK3mnY36KGa78htNWIT5Et
5TPYuhsBeCeIcHP8NGjRRkoNpRqXrgRTO0uUU0CIvjIe5I6Hrw3Cc8Gxhpz6umUy
NNRDk1dPT/34f7tbXqTM1JPBohcJ3MNX9bbmIknPPMqgodjn5kJnNFz3mWvLtADc
9JhEML7fEpyCp8qjgze6GbmCEXnWA65eWCC17a0T5B0b8/eaHNp0/Xa30J84zs9d
Jizay1u6RBDWqmXH2nAM808nUtofQl3U/hdLetGEVSKv6Z4nhy/ZafusDn2wiI95
D3zUzgc8RxY2BMLsLJbGnjilTTt1V5aoqWNXIRQfvzVOH2kxqrlPliOKsP2acFuE
g5FtTV1/kJzSOcKcFxOEx4xdDTR5xrcAJbM2Ye2zXMUrVKLSeCPOvnA+F1kdRYiG
PDbVfjCBJ8dazptEd0MzhjqNK3qRkpmlh4WgY3gpBEDBl9c+2CSlpBdHfCxSZHRC
Ae684E2+c2WhSk0JmtXP8IWS1Pq6oXZbfL7sYVZuBVAwIVcEI8IGauyB6+iXIglY
3dVjOsrQtqcpJPK4CjRmg3U6pdXPUObnaRU3fLOhfv16AmIAg4hO3MezYOqE2xLu
KFsR+mq6PYWeYIlmVvsu5+Xm+Tj6K69kcMsVQoKQGZVmQ+EzUxoN0lV24nJwluVg
G92Ulc7qonSVMsSE9NX88jXQxVwl3lrttUSaLiwA48fVp1Ou4hEdhC5rEcZuDKYN
DQmPWik6dCA2q/fOhQYZQzLsViE/MWfWLkLBZhuOG+sYV7V+SQTCx6F5NebhfEVO
rj7j91Zvxj0BTjW7OOu8RmTNsCYSBD+oWdOOBaCQA0OjblpBqwMhm+aKrIBTl9Fe
WpU34f0zbV9PawqqkHBOOefmuqxFk26hHmbyq11zpmr7rzz2LtxxjnFuzI8cjJP8
NQaoIASIf4spU2AT0zZbJu/hpnnpSth6zHwV0ybH/TVLxewOtNfJjEDHpvE8MwV+
Nf2v3ZusVTbFR/ZkNbA2wkhaEERcAMmwcDVQJ7mnS5s2MWEznk/2pPgrP7hxbl9x
YRZkTze0J8ejgpfhFKEfnCtxtjnatrvfQKvCaBThzQFTAO73gbF1XBOPRkGzkBeP
zsTFgV68M5+oHEphaKnkLDMiZna6kxwHkZrktN5uYuaHWW/xo5ILEFr5pzBnWIav
YBTZdYAumniz9KzhEnUpLvqvxYCbvAT2CxsWsIA0lBTbNakLiXgJRmBXDlJ4kO0b
4va/YrPOw0hxxs3e9SpuGZwmfnsQkIcv1HUU9Q5fTNL2TmWqubEw7AAtyPZ7RMuS
PFsqQ7SgiVWwQVG7ZZo2iuqVR3TIBlOBaviiTX+W40FoKlEmmuIkuapmDP2QQhBB
tXo5GWBMaZiT/lfiv0YHCEWnPwElXPQ2c9U1kSK7RCBuHmZ1pFVvhAURspTNJ52B
hZCwzhdz+yS/Yi2rrPVlwpt6quQQU9dSDSlNXU5CTfUm6McCTnlmqlwLxwxHAR1f
6xL9QncTbzhFNfdlv5ubWvSIaswqC29FS2bNqrKR2Ok406KbT/EmzeP4lcUc7/mB
oOCqmUKC+FEmfcNNpccwhkX5XzGsmWVQgY4QUZr3FQ3FYPAVDPGyEI5ApJM+b8qK
YBwVwrud8/nnzlZd6+pgNSAfEvHe9Z2kcMC+0iysDM8JCllvjriZeMUQvtVNcYLx
0j3Yx1H+u3N3R3VkVCX9y/iHCGPY27zTp4nrrylagVpQ7N24nxkuhUPsL5rc8vOT
fr1PEWPo2rbkkkmgwe6OZnIHPAao6SnZ1u+Mxp7rjwlIpLt4zFUxTkQFYquGZQ9G
6HjQKTIi3NNKF6hKxJdF7wqGVR3Ui5ZbPjkplUN6bID2Yo1xXBUY9jKLEgn58hO6
K0LYbjFTNPxKjfDvTd6zfJeN80GB0vzLePgyGTnjJJDDDCBM0Eo6A5IoTbOdZtBA
XeoSwUuxW3fNTh0ZARsHmfbwPueoIY2EDuan+TPaP/kDi63V336XHDPbJo7plnMg
FxvvvbVnurRtkIgfRkXCIJFskGGjCqiNaoH9FOGcHo/WoXXg2kbYT4qXakFlu7Io
NjVT2aMQILH6x1rl3381yeBwKCy2Rp7R5KX0EHF003hXHGHawfl9lngVZO46lrKW
VACSqymETD4Bv0B3Et+hfvtJ5IrR5bjCy3+PL5pR1/FylMzwq85+XSbuqBRuNlBo
+gyPFDbao4W2KG4YbHCRItwZa/bxkrJum2Sc9mmUzqHnJIZgh2l46Mxr0U1iQMPT
M2Us+Tot/d+nTe3jGEtoxMcb9qA4YVwN/h/vo+a0eTsL3jDABGIfususpm1X4Z7f
dqi0sSRfxUuZQlz3vNDL+W5MIlqb0w8+MUBiHVdyV/L0/WKauW6PFi7vB7cHFfkA
/U6t8i8g0kti1VwJmeVbgRVGE6Dd1cAUFqNYVg/tgqNsmvyM91Z+JGunyFkKH2Jl
FzYLTwN1THIZijZ1lYy4LbegHG9qb6930V1vlLVQeae/VR6KPepRAtMYM7QTVVES
J/i2aoH1qFSx+PrKoGM+HYTDYWw4iI0GyORpqIGkJ5l4CLfihfb3MSITiHRgykl7
trKmKuuvn6Uu8aTC9FwP7KiaIAvRqe8jgw1K5hViKMtZaEJ9r2vwZejcSR4tXawd
KkG1nTdl0ydRgp8sUXPoASjEQ67tGYa61xTUHVly/+hIcIML+alq2P6JqNf+Zzke
OmWkEGwgKqrOGVHrYUj2K92AL0+62WsfJ1x6vz3iQogyaXR37tALm+FNMJYHu1pG
y19slGZC1CkSgoJ7t9jRhkLMEbhV/9MjVe1Kuk+uonkPDF5MEnUSFx+6tihJwbh3
dv3hCCEBr0Ug2iLBgYD90fwm5gKNuhtE7Dt7KQP6hJwc7B8RwMjl/anpIjF9zJPh
kpwPXpIyN4suYd876oLUBw3MCg9TIvvBFvhYBTXR1rM3WJriuUm1z2HdA5A/VM54
i0OfnGQgNg22ZImemaAOW3VLobtTFlpa48JzW8cOZkQ8USJhkpvZeey+VGLjCeqy
LcN0IRPL/UitXBKYJhglyMhYRd5N3bjHeQQLq1DsJW5sfK+NPLZ4j7xpijhUba+I
LJJjtAMWcmvIHP713USwt+6xsgEC3coGX2o0hV4ZOrZaJmW3Lux+GyNZKaZIlWLt
owWQ+QbvjEQtmiizK6ww0GV1IcCTdkQuCycstIbLAKzfNfbYsM04UVzjJDCrKNu7
mKY2EVZeOSEiqCjQUZF9ZA3sJwwcG3z83QC04zIePSHvDzm1peDmC6cEhnW216fn
HDAX3cwGeqBJsWAaBQfJdDtHyWbWtGYUh9RbkhF0FvpK0ToBLx3Dh7I6fhmi6qnh
WKmMF/nydU2yQ6C0mkTBv4glue0B4m3ita8W3t28xRDGh6yBbvw41jtlsM5tM/44
YHQ1sGin/IPixkA2E9Rw0NCWbrQ1fZ+gcEn3ORSb6zHyLgmO45xgeFrhl6dbae/e
ypGwc4wlZj7Zf2/8KnR90QgZ7srbxRDiY4mnU+YhVJVEqWrFd5ViC7xBRvw3LhFl
SU3QNteOeuBCZFCji155nubhHR+otC0JzM1GsbE+YPdMAT7oWk9xAMftyhGRsmIS
RIX/O4701clUP9iOkv1cW89jlVCuBaceWOZRxH3WrV+8X7oPz9Cg5aqq555O4Fx7
3XiUT2jiXetxcO6Kg21W5toNGFa9QptmBHiglKTTUNByqnZDmXum+uVzkSJ0wzs9
7kJGZbwDDJcM9baUavpMstI5n9u4e1fVrlie5z8tXoGuH+ZilaZx9gSSpT3UOLVM
V1IzANL9643SXYl9VGzsO4Jtec86gx7kyVHoLoH15OWXBj5EU2Ee7k/nl/sC7BPy
eV37lL2ZFjb5vwA/QbrlgWlZZuARgY2xEPpQuCHjLwzRrwPUQeoKSFU00krdp+CT
tK+sHvSpuk8q9cTXyauPfJGygUlt6S/YZ0O1zGrifNdAgSmuJqThTr/5+EvY9gcj
cgtcv6ftH9BVg6AAjGWPHtSGqT1/pjARxDjpiwWKokZj/fvZR5wOT1um5JUaj6yc
fe9SQVuquztRMZSI55S7rrMwTNd4xTqCtURkrhgg9YpaUJbgd7gjKiuDEmpcN1oE
BrFXU/SYGZwSAXoIdH9fp5Nes/HJhP6G2u92XWUGZhlNcJGj1DKDR4CrrboVBAmp
8nh46wiEWDlafwDzanof+ldprg9tHw17acfYmY7d7s2gwfeDt6xvK/WATofKgAAg
S0NmJ5N32X+mbw9p3hYIO+L9QSKV9UfqSnMbpyDb+5JMw7N33excVpP04+3z1FsM
ntj78prdkPK7otCLC11g/jztiQcJuzxWRmtmS5ptxX3SLBWDC6gqhilKzn0sbAor
qI/8+Rj8UUsrJ4M2AYq+W3Z9jwWMiATHJu6WOBuXgPD172T/klj098rtDDaOWKQ5
TWOYmGS0Yyjsm59kiPb6Td7qmxuZ9sB82nz9CxXWLjYE27/YI6kJHnZy+jKyXq6s
IS1R8LLfgadCk5lelNuezF+2UdtJO2rRRovwd+5qCXWSEufXS3eHDic1fYKdFsTm
1Hfck2c/z0wwKAJQf0fMxi6vc8AyovTDtroPc/RYZy5mKhdfciOsHMvkdvB2hdkb
M7de5u7aoJ8YPy5HSgjUxhRN+srgYfj5AZPYrdlK74Ssr0Wdgz41tyyKiWD/18Te
n9o5ZvCm+49qlQMq1dljoFhBWh4VwEzkafZ8UeD9BYyGVfFwQtAERMYAuFeWqz31
Yb/RUowMEg/Y/sDN9n3VV+Gb6NicOWQWAOH+bWa1x8TpVOysvssnVn58jofcEkrU
PGUiG9gT9CIYcrYur8iP9iy4NFKofILrFtwjeRT4/Ot3feun9+U9JJ0tbuChPd5u
NnjFIz8UEDFcBWeR0sDHQM+7r63Wb9EHOW+CEkHDyTZBNcnubsOw+z0pJTEAEznZ
hIseJoXZMLAedjekPgVKCpaktEqgsindAAZfQMInt9auGOWuzMk3yAsXOo3ZAKJT
7nWqk2NeL+z35pB2u9mOUl01qsm26RIPjpOuJPwJYVX2rug7i1C0E6jeC74N1gZz
x9d8lYpKuhQqGG+aF1Hym2xUJYE5fWAYBvZPNtuWN+Bnjz8X7x56lQiYBXeyJm8W
9TBi8/40fnCUodCruh9T3UMzrHk04luAP1DkUeAy5Yyog4mbUOGeZ3EvsJGauEgD
92fP+z5pbGbJ1BEwOWlSpmbPTvWHRqfgtLmemyEWMhQbugQ8LJ7ZksOrD+JicbMz
Rl1AFu/4uI0qGBWIQSF2vg25X6c6aclXrD6O9s9XjyLgTWn4ZH/FlX92I46yH20U
3P6OTCm+430M/KOxeyapMETtJpa72t9NOEUQerJosaAs425ivtmlSltniOyo/23F
PZTijQYi8SW+9VadA7NZg/cfm4997qElKxHw4lf/aFsg921ivVRhtCqYUL6Js3UU
Km4GdKrkbJihkBjNWLt17aUqIIU/RtTDS5+Y7NV3QNLcZdR/qvQpecMBI16yMN/I
QqySGL0k/h6n+OynitTlOjysCvCUlmbSWRAeCA6cPCgxK4HJs/jnl2ZP7g7c11Nl
Me5P00lV8VJ/MYhNbaIqTgVBwrl92fbx2B6CzjoObnByt8zblXO+96DKU58eOERo
l4lTvXbngmNXNisNmYvNrlNHiDqrZV96/n662XsJsGpOGGAwhP6zUi0DcYKZXMXh
UOflt86zvXJ/gKj7e26h/Ad1ydCi/t/FWVOv7yi4rqDutJc128f33ZGlcxrmuiCt
kGM+3PvFsfw3t0dgE1DBzu17gKdjPDaXyzHLyTTCCW++blgotdMYpvvIABqN9BG1
qfUJSJnj8WdStmEZ1ZM3SnkNdqcyKTu4fmviYSuy52Hh4bwPG5xqP1qk8TBbxS3g
/vVXwyeAQ4uuNGV9tu+z/N9for0ng0zAwckYIJO02ifT7T5U9ahcfkaG4nFHIupc
oG40UrtR+n8FMgocPDLEI1QWxqOa1fJb1qpPK07H+GtAgEfwif+MFJXpGaIfotGA
3EpkIpIBY2f7IQzYqOPrfrkpZjasWMMp80SF1t8bqObLKOrjcRGGXexD6qHxdUL7
eEq285paGCz/VYx3k3XjXyDp9VNvDCBXR/9pltQaejOXtVN5GgESnu/chGarI5J4
b5AK7/Amq5kcU3u2p6ZAnCkdRaPmi9UBZ+rkYZpXKMTu/nDgXfPALAwdKEeiLR7y
kiZzFt+Gs4chYICa2Y/QX/V9Ey8gMdTdoZ+pxjcos/3zupHYWjcTEhUf/v4g7Dg7
DQEk30ZONBf6+i3MnclC9Q0cpxVgZn9JQ85p4IN+Tm6GPiw+4/9syDIl09rXyCzG
vH0BjMftiGydEgw/eIYuFNlWx+Da8sn6xvOBDfNJMB5jM7ye9lib881avIdvl17o
GjGrR/w7ol9Flvq0SQSUINNvTx6KabCZNwNhsVaLpyHGTY5msL3RqdcaldGPEj3G
nnp5Cm3O5BxjhvvagrOWApjRMDylY9JPtd+TXT8pshXA6oHCuCGciZols7vnBMDm
AjqD/xH5zwOqKvwR9q9Av0aiirz0sVfwTNFR3TfiynM08XYtmTtpRBMX2osD6Z8c
ho9wMak5Gpm92+Tu4EI+sLGehR6OcPkmQyo2p8qrPuJ9aibP3CL7N0e+USGJNvmu
1hOZUy4ZD74soiHm0T44dNRvWbvmY/i5oIo1M1goQa/InRCcvSQBygq7E9dDawIb
DksLCARmOV3ff0ntQNtOm+gy/X0cSnZ99nQatA4aSwkCM7FptkuoT55XrWekGlrG
QXDKN8ZLosZ9/rvfV5Dnn04Cbn6iLtjVa57sTZqVyPw+OSjA1KH/C1n7eCsdB8aB
bPVihIt0UJeuSfCsF15n0tvoEifIFQqgwphIDez4yKpHDazKivIO9OwGh/RgmE4T
e1Vwebkm6bMO+nGuCW8JpjIzE1NnvP9SoTKOa5VX60LbvmD9NWxT5By6jot/aEHY
j35u6qIkaeApE8+8tN7teE3mUqfPNYhs2x2A/WshlQDx4i9qZ7PbMT9MLbcY2wQ8
bZ6U83C89Jy/hOU6py4FXLvd446154FCAQUJSS1BFNEwJhQVnnxVhqQ7i5Da31k3
eVth+D6jw+/1mliqiMuU1oGTd6gs6Y9prbn3jNostNCodkZFAAc1Ci/7qyWGy+3+
N6IXUXQuoAkFbnrLdlwDizrdRcMNHnDq/E+JhVVHO2h16LDmT1Lbqrvzoym0A0D1
fO+Wa7Gc4m4FEDOz61NWdCn9Whid1hsQ2Ab6kVGBD813Jhgm8ur0Ejtfp9amKEch
bk9pnUZ7Lj4pBpTY99/7mV5SDQuOuyya/V9Fpc690hCNbDv7SmtWKXvt5zw+UwwF
kNywTygqP2uMLUpLphl/c96FZvnSP5S7UcJLeiZjAtzCcq248Iwo7Lge0pTeT+QH
8+eeCkZxylDZ3skUmm5VIKcVtTW2Ek/GS1+07YBtJJaPLYrvZ03jtoL+vMEajSuC
v2I7ld76SANqUpxPNQKr11+yD+yyU7ieJlz4SExhMzYbldLGO54ojJ5srde6kEox
SapZ1zcvMM2VNB4O1KQxJitHS2uJ4Di7JU+TYV+TB4pxr59fsWb6GVl6uUeK49eA
4p3qjQgMEBUMmMw6rwwjsX9ZtWctEV0xdk1RQxNEjX1XxB1/V8SAz+/RWoY5tfKg
qtixoNjTj3fwuyJWu9XpyriZXiEB5rdSJJHHfnDT0XZPGLCs+x93daM5N9dNuucj
659U5BDTmvvvZnO4NQhLgpja8RUlx4itzPID7v93MW8r1DrSAEHfPnr2M2KSMSX0
TlW8KV02qDnPYkZCo5kYE7NkmTFTgC3qM8N7bnjKL+LvSwSmEngsRpwbjcRNZ/oa
Nl+KGMztRkF4n0/60wotY9lYFzXg3RoOZRxjZp3KLGFioo9X2HVaXedpT6GQC4hO
8gXKQn9WksamRP6226u1PZPhEsF/0QLLmZSmG5dGRccDILt+GJnj5gA8/nVpMH+l
XU4iize+rMXp4D/FI6UN1J1LqSsLrnh85XMBcwwMvD9a+PgbBdUEXdGzmhiNjJ6l
tnQHreiHj9I+eCTScmTfOxRE/mdf2ztcgU+j0Uk4CSvOHp+VpFO4nTPqddcUg4Nx
FmCxHpf79a3V0to4L3Itq1E0uZHfjAcZefkGk65GxvgcMTO0xNIWP80hca1N42iV
ROr6lU0YEBk2Na+iLv00ldEtxzBZukX8SvcZQjjoeLivvnAAt0oLaQFnxKnx4OBI
XfbrF6k1hMM0Aw0vAsbnQq2XLUPGvWTG62pBoKG0lFKZx43Hb8jrb3xJkvFKUYV2
FhKCKYTC0+R+9ydGFXy8TNMc4mvdN18Mg8pcUdXtd1yJNNjswS2c7VgqaYJVeAYZ
9oBGOySRMtavm03/E0EmMyETmkffyyWjkAl/ix2gjFrv9NtDOFRfZRcTkCaIyx3Z
gC5t5sHNfoemh0CIfuxIY+quw9HPTXeZprKGQfMbYt3fBv8AqbPvI3DdbRSr9yDq
nN1mQ/Ze3oY/ekQJwQTF4wlrbcuVWmzbwKyLOvIJ8kHXl6+Hkzpj1ZSE5jYA6rqx
bKnxXPF6U3ZIktm22CTtj0FEPh3SKBZHSD9uJvaD7EzbuE2C4ZlglX7nH1ItWxuY
h1GCt2ryCqo/KCJxD472+AP+Ngg34J3VF0fD4tMp3NsmO/nFGLF59+GKazFqb+xV
BLxfkFKhLHVQkTrKuQjzXi3C7Nw5yVgVnezGvDh7p5+bq41KppD5bmFWSUPk7CuT
ojWwKTDeRgB/1zpH1Dd3mXi+MqzCvsi14emQqfip1J6CtKSWVsvaTBPduqKWikNG
DWZO9m3Z7S8VIBJun6jOYHa2eqSbYT/UvzAzqi48Mslb53OaqC4QYfkBZq9018Tc
Kr6DjEQdKU47PFqEqMdPElPlA2SXRGLBcfmtcfQW+csleou8nCGx7dVXscyeOE3m
oHkpHKfQAfXwhRMyZ+ekUH1Uf88YPHQeCLcvA+L3VfTbGwd79uaslbboOS9KjS2K
JMXxMzvlPvWIq/yjP7hiQU47NO+0jV7ylmfwDQha4AZ8pwScvERTunsUEqHlW6Yt
RtjgQaBFBxLi5KnSLkK73IKsfF73vDGsMnF89g3zDb1ERX/R7HDXRkKuBIQezQeU
owacp9K4RfG8lT6UMZ7Rlr3ik80URaLR4rjUqWfxU5XypAAimE+ZaZZ36U2vqz+q
FyTs6/p9I61xI8WjnvRscyeHfMMLOM0RBBkufu5y2zEeYbf5kc/OG0K/XVpLTole
6qmcEOJ+tB3qIlSXevPaxuDB/eigp/vMEKj1sAGLVWrXIQIHGNMC+ZOSU7ZnN5PN
uOS8OheQrwH0bWjVEDjAwSqQLO1NpB7+lj1H+HPrVlXX1PMIvBxF93JLzA+5iZhC
k4qY+vIBHcHZTCATGINeT/csuaH11SzxZV+vnlCPMyfYfYo53GAPxNT4xJZjE5do
tBomSjoYE4tcz0hiSVQ51U7aWEFfyRV9S6n5C/zNmUGa9anJ2TOSjOmERYwOVn66
aBbaKIXwZtBkNM4Q+iK4kUJojCZXIRepgwlpswcxwwjUAnwKrbMkJ7TKJQCb85oF
HHnE4oX+bGR4hmRrnXIQVoJ0C6bU0F3u1frpKTa831a1idjfNn0Xp7jk8VJK4V8C
CYt2efQUfa2lJsJqxTfVfr7at4quEATd2hX7HvZF1dAJpdCtBKzfGoBxzHo6O2er
L+JL4wyuwH463ZuHsXUOLIuTBJc2mgB841o3VlPt0KhmVLh2p4mrPJ9Fn4Kvnfpi
9fzt8HI8ra98l3Oio1/BwCaAysmrvqH9sm9n7aan+9QI5kbF7lgsnQ5M2I24gw9F
uNS8SiSwavprQnGwtTofKweSlAn2fkaEimtCOzp9+cyXTht07qqkC2LTPW6LKlPg
o/c6RRBEKDOrh/1Dslz/5GZmz0agHGaKWkJ+QQWB1rZhzZk+/bkihZ1J3WZJf03r
lHPv5PRmax9uJ4lPWYul2ln17y+q9t0FqLsDOTN2VwlITugzeA/xty4BucXRaaml
QEGVmpPCbI8eTaq8wJxQkCqiewgp5jRdlLpKhoh9/7YkF6EtZx3sTofJu+szLp8C
ZWxlg0LRn8XmtdpoMTQ0fh6PgYEulToEzMzf+1aT/MZ7t3RMQOo4jDqkzePkzgNb
BuLZbKzaeeSdMibYVV7MbtEXgy5Eomfryyjh6/+HSYHJ3O3XxwxgUoq8lPFollNZ
Ez6OEI5rl/q1pYd2uoDyomfbEqVDTI/38kMm0oluMY0eAsKLZQqHf21blUo9EN2N
WgalqSmxczGCvExN9UAYhkLDRB9OSPLEBXYUSL1SzFr54DZT7LHMevPmoMqrDGBY
7MLbZQDmc9DiycQRWzRBfzuiMS4Fe5trzqC2DkwRt0XRmPuwE0bz27RCaRT3JBHM
P0m9ys3Z1+PStjCA5pWZITtsGTycBjF+WU3EUh4FZ2TwnY6ftb83NNWVTs1QWVFP
KkIh46P2F2AkZLEDjrDNEXn9uKBNqQbflOWYqM3wJu7VMof30qdmXNCroP7SU2GL
8KuspULLWL94rve3PC6Zm3yHrO1AZ28AX23UV961OnTLXkbZGmJmxpKWiBYHsbLP
kixVLNnkHfPplvt0Qbkf/0WXOO+7AzTDv8Ia6QnzQ8wZXNGQOpNLC3zhOCzl0vt8
yZCzHvUAh64XQrD+G/tEJ0EJE+uG7xqS7H310TO/hMto2VcoQ6XBgPu1ZHD4cmMR
QCMWVAl2FYFS8yP+pCVcS1ZbeaXm9lV6b3yudnK66dvmX3Qf4xkgpSi4g3kxXwoK
6KZ3FzvlGp2XM8Apme/3yurYY0b8xWq7FOHuVJZYX1oErra3AMbmETCVZAUl8jfB
rtWMsitMYrbmXdg8BY7RCYgGWMtg/JO4+FIZ2yLqsIMFIZOAbumxYKfUnVSaRYre
sVhk57q7td+TU8hm/MPOcTyZi5c1hhwCKKQnvGSWRozD7ySRfkGrFzlCyBTQIYWd
uR3mSEuOhPp9pp7otQZPPRIVW21YUrL+19a4beIYpLOI5JsC38ZUsbpHNOC4Xw4Y
ZUabJW2+jmt6r8XSMIes2HnDeACczGalNIWm4q0bCOhoWMh1aiqkqEsYnhRft5wu
WLFvY2GDUmFyd8GzzgTUWv3k4UzwzspFEy96xLNN2Nup+l+yGFq0/FwotlgvZnSj
J5snYMOpOanSkBSOA7/6fk6pRHWKYCz3alSJwdupae5j2Su9xOMxJfhOsSoG04I6
8jrvir/Y8BRXrMAh1A8nGggxv4mQLYbDxvmUcMZOppV9GuUPWkEOkyMWoD8Ig12Z
a5sy6eruAB+WFc5Kkg6x0ZqcEDKzLoVXX60W6XdCzvX7zSHMD8jihN3p1/T6L6Ka
L+oxxA0OQjspTtKNnwfBf58qNA8wTGkg3oPPvwlGW/D9kFnb4eSMMM4MYCxD9fu+
dzlj+m7wnpSbEeTZBHnYumWkx42APCPsPIlp7YO6xq0RIHxi8iYlzaejQbQe9tHn
AYGLkFnT6PPVluGYTMrl5rNELr6Vw0+NawtEOTghxJAz/m/3UQy0j1ZvJ7xaZhzG
dliO+1VKjEn3gVnYZv3tuI4dCcqnfy9pQDg2T+K4Tmqo2hQU15D2ZIoiJiqaSmpu
JL/ZT78IOCTZ8/+T/HIiwjNzHOUwN3Bx7VgqPcFs8CM9MeK4D1Y4WJC0D1gU90XO
+P/eG1afr5Aet2my9nuwG2EwMNa44KKQT8vRuPfEmIsTpYPUHDrVXOa3p6tqqeOx
0OttgyIBCQE2WIQ0zT5RCW6e3CZWKEQdlkd70XlBRjdID6zgaAqvAS5liEZaNALR
yfCUumQAcTfEcntKXwLRfKiCiZ69H+PYubyAYfmVJnQHZ2e3MMrKLyR2yMxgn+iH
c78Kga9MKsK1U3JGPKMPRUqEQYJCGlPy5KGnLkymEnliIJm1oIQ4sZtBIrVMk6t8
wApz+BR71bQxnH5TjrEwrW+rthk8QRoz3Pvr88hr67Ops+ebTzDvLpQ6L+z0LUKZ
jJIcS0GXLXKkvw46257oVY4RcwdUBB2PUjHgP9w/qMS2s/59TEnNArEHnSClG050
JE3VHE05AioqNAPe+oUxoES8alDhcoJLgjDPOrRw97sBv7Ag4Fl954qlrG8DCQLX
mJrKOvRjMhZ/McoktVRSby7otQthObUAU/3hR3yeSluebsin+mQb2OXfkPl+HJpa
v7v4QwowwIVeABhnW+v6D9+vxgx9ndFkXoA0lTNB2JawaS7L6jPOZ9HYrcbFZlH4
8Gez6jBlHnHauGxXz1IvdFIreAy7q68PeLHLExzVbDWTFTxhox4+zag0hLDb0F3L
VfE/bWatx/Vq5W2Wic7mfHm0npgP9dspzTFflY8Db/imvHtgBRvF2961Pm+M0fkq
cLQMDKfyEsjn5AmGTGZOiIJrKA/6lTEti2H3/Afgu/83JKlF0+yC54F2X3/rPRPx
lrtjJJMPfavx9DZgCNt0ndkUUrhfO+oZNhc+fTK1fDeGS2gZMJAtX/51SyjcsU5F
/2fSqopYk/+taxspPjpQg8Xwk7OIyS/ZnBexQx+pqUVufxvICJXFd1Ra6QKMPvw0
6rKuar8J12i07ZhYgvE/etxZplnov/G5hENcWVhoiMTDKTYBTaOBP+t1bPh/Vw9C
2bpH8OSMYjccm7ffy1wwsTmjBlYNHVaTW+ldo88vLa2BCpy4KPstrXesiYGFXKvd
jwxYTkYXZSoel6tfYcd6PyiR2ihOlKgIReNSwq4Qm7jiI5aj3c/SUke6geOFDvlt
5s+M40cXJXEV761OMJfw0+MoJo3ino0JWaHEk9StRm4XAsg4JWH9xu4oM5Zqdrar
zlLvaw+VIO+ob517uD5UX5jzweV+hIrIRNuzOjo4t3YcAdkUmlzKJnQ8RzzLkeBC
Fhe/18AWDFBHDsMGQ8OgkrsiebOyHmp4OxRraOQYrBV4oiAB7XMehmATCTGv7HcI
loDOlaPZ/bsqv8/sHb2aOJy26zBeDneS1gC06j9iOEgKNhS43qH3uVCui9YQeTPh
LoLWXv5QmERhCXHa1RXWEbcitUBUXisd5LfEYBHSfzDZnKAgniQiRtSj5gQ5XVrz
UgxyalCMfEfQHRLfTI2VCtMUe20QJeNAeqIdQBoZTk8lOdeCZ1t/haYoBfUJ+m/d
2nD/aMvQAsV12RndNaskm0gQZv/OEMCTAq86fz5LzlHrPZeTAZ1RcUv6UfmThhnE
A/yXcHZ3bvVWJdh0AEdOa9sy9k7ES8fF2lBvacf/GbPhtGIK8PJA32XaQh0nnybq
0Xu6gPomez2tWG0D30B1kpDcnZsYxU36m/4dwMgqYUcU0NcoYCCQeu4ZppPHTzQy
bWsHdrBgBXoFh7n+oJDb427E4dzFxjTDufPYfGUIn4zccj2AEEUn1UgMeh4TsL8d
nuCC9mOEZqFNSrOwdLbF30TImU5d/D6nGcdm3pnf0UK5uycBPJUr6iulp9dOQchu
bBSD5Uiv4zuQxG5ud6BoPHQA62yrAUj9DuPzQypg98ms+xpXtsQ3aGaY10dG8KLk
xsHkNHmpoMNESZZWqTzFnvu+3hiWv7J1u/RL64K51nPVRp7p0Jhm00yNwJZDc6/G
SGuZdPWadzrNP7GEyTYFx50Ld/bThsu6WpuwsyUj842cgSsnpFEMear46bvqwu6I
K+VqRmDV3mMFJ1YwVRBZFfCaOArCYH2xCCnOZodnA8AIk1Q6ZEWWQV4eGWeZc5IP
bniSHUFhpmNROhZyM/ZybaQsKiRPkVN/gvcOwgBabUx50maP3tnhVr0r6z/OC2TV
EHdlGkiEJXziMnXPDKMrErbpGWyLZ9aFew+zq+kqUR56td5/Ai2Eq/I6WnnOdBPk
jMLUfOW16nQmty8k5ufAtIa6DOlGja9X7qFw351dyrTdKHzW4KgTcTnRCSq01hnU
kTO+OJH+gXPJrDPrWTjVQiU48OXV52FmXNNypKwTKYBi7LhQL3ZaLteBvTn8abzT
FyhoVCcZt1oG/w4GWI9QifeeSN7rqXt1GMqGJhhac0ocb3mrN+vhs/L7xOE6VFVA
6VrOmyqkKd+tNm6K+PwbRFkzW7cGMbL8KStZiwVfsa2HKBp8CBgr2AefJEVj7b+/
gJsJymAW3Z8aaWDrkLOKFPOrRTZInCnsjXZ6RgDcgQzkm3yg9wIbXXWNj1ymnTDg
J0Ga39nx5WZuIYd8IqsLjyI1AI8lo0Vz4v0PiUKrEHOvoMrwfcCipFSEoVa4Ugrd
W4sp/EmwZkSYmlq1w2Tg9zPt7UhFKkknRBSHML2ws8aBRXrdeWNRsFzmsYti/UEs
ylYl+za8wLAEvv1w3hdchAmCSP1KZpk+SE17B1M8fHcuoStHSV7AMYLpIVnzxf1G
Ny+dpCN8z8Vpc8r6C/m9158QDLN+IjbGPEbjbbuDD6XLK1HeXoNyaAENG2XbFne7
WlPcI5SQeW+ZX3fcLHmfuy8BFV/jJGvV2fNSLg+MHMcM7Tv+GX+sRxwLHYvBEST+
10hFzbB3Vc/ogYYV3yvUgDtDuGiJL64YQ9ShLjW1+oTy+kb9S9oEV48DIcqqgttj
Ni5hGUEV1/ve4IpLThAisQF9HGFarWJtPHRk5TCypaNF//CSBoFh58uqyTnEzJxZ
i9e43VdxDbt1Diocnd0QEoFTy4Hg1EKyaizb8cN5j3ihlqMkrZcAf1I/0XUWPxbP
73rOw6B5CgazPOE3RgpN5rUZdJI5npRZVRiTGrhVTscIgvGlDWl8ChdTks3VnA3W
P9l1Y3DG/aGuv5PD5mHBEYeC6AAQDU7/KzM3+wzR6LPDPvmOiL8Lk+2+Scikwrxo
dhEkFj5ppeFWRRr+dcJkd67ILkjpzL7Yfbh2LIzIYRYUUj3IeAGndct/fmMPLya7
66YaNI4W42LYm2CurClBV7r8zTwV9MarbF6NYBQS9xNJE7rtyTUC4pnWYedXUQAo
ehCi6ibamX5Cv7UxglfFfHG0pm2RyLQrwUvRk1cnF8EnMV3DL5h92v38U1mrPKXU
9qV4KcLFSlxYHYWBj5fmLZmDG1O9P5I8zeByiXMaOe7IY6o30omYKY19F8Qa/tmZ
fV31SctN/UW6JGuu6lzgil1d08NE48kdbN97wm9jgg1MAt01mBtvRTRlmr+ktlYt
qf2bHJfvSmR4y1SzAULrvLeQKh2n/uLXg4q+REge/2hV9/brgRtio62HeJSzsz3/
I1xvToZEUw+ANSxNjnkAOnjKC1tcFx7Vgb6UnfxAsvGEddBfyarF/UIX3cQj6I9R
1QRezuscg3vJ9Dism9AOvINVtEr5vrMnmYhslV4P3BSmb+KTsljKh6i2Wy9En+Aq
6QWg7wM48X3wXmXTxSNd/Vvue7Z63yLlffpCVodgQD5LXdS3nE0Fu2BI5cKX9kHb
9yJKEX5wgAU3eV00vIM88r7qjeVaKv8bvEi4oxJD73iGF25/kMJ8h9Mf0ascrCHi
3CzFNRlMkmGSOsslpS1u+uBs4ILzbHc4lzKSZJXBVok0CZO4EJj2S9uxWy04rmxg
Y802I8lV2zS6Rqx8oOZQ7I57hf14IlfCIjs8JfVpX+5BaDslEILgS5D0hCFd3GIX
NKFE4LLZV0ysJYvVpow/Est5sszTNhFM8WUXpdJS28BSiJ1z9odvtUsR3ThZK674
pobRuTpu3omZoTMQVDNSL+v0g4E7x52FOH0NMcn++654gIRXmtcuO0/0c/X7aj3z
v9EFgtBzktpJXbNYxZxfCtjOqgEXlcqEKHRjCFSAcAKXlZlo6+4o9HFHHFewSlY3
FqwpRtdecEeoH5CZQ6e6K3OVQyWv6lXJwNGIgT/9Fi6gZ/4t6TOi9I35WVGV1vSw
u5j2m2/PVTVyTtCZHdjRmh8IkcIwj1Hp8fBIf9yXhedDmB+mjdL5EOEz8LaIA6a2
1VRVNrwB47mQEmeRhh7mFW8rAls6aocdURqZFglgV7ypxiwzlM4Hbn/8jMQzJtFQ
g0BbNB0RPtmwUJFBjJs4+gf/kA+WOAWmMXOUOrsDa+5BUBCev/PwddjqGw5EmnYC
Y8S6O5y/fgebvC1uVidE2DoNCA+hiyW0tns3zqr9XuiFzZsCRkYqgoDaBQkRrR/8
9GFqZzNZBL9JNqWQaTrMQ5CiThMDKnHKOjlKUqSgbsQBqe0RPF6nQCK2TyN63SBa
IHAGrT4Fz/NOjyX02JivulbFp3cc5IHslp4joW8yQ3BmK7s9qqV1Tjhy2YsXPDmD
HjcMAAufGc0Q4/SkDrqfz5Qhq1V3K8kO+lgtrL4PtQ1VmcOB6SA4t9gUR/XUMC7l
ksTKsCfKpMvdLyMX6NOYFl+hAh+mmqcEYSnPwcnXpeoMvzDc8BEe1zQ9sHdwoy9G
bQ0zwioS32e3LJnvCUHyumWgVlM4yYQj2sJb+sYgJKc4tmhpqMB5wSzF30WgP5ug
f2AmZNI/q/634YU8Af+87EHDjPi7PcZNsx4cmwcdLlML7uQNdOl1NFNC3xuwD/km
NERm+Q/ft3dGQl4dhQa1XYCnvEkMlTpJKUg+E+OTt6lawuR1u+yY8Fgo55tYOBa+
RfoFG3TQ4e7Gnf/6eWCkMjgCW7GjcImD+rFcg6ogmM8Wy7AlDta5G3woT3tUS+L5
AvtgNGwk2AjXoGTddUZtoCCwgdXf7KSvPLz0tVNE281PzZWfkYX7nXbhtVBurqIb
d2ytHlTeyQRUXkrC/F5nEmrHKAER4brmIr866MA8Z8Px6WREPTxWQWAr9Ng8n687
VEGZu15dbnSoFniesbkZOpnJgxR1rz0OpSXiq3Noh4EoAjiHMae9ttdWJQmmOWXN
gsSG4IsZQHTo8hkFHjvt6le+vr8JMwyKR42PXP24RK+nQ6xdyOrSnZrkx7nmZSiO
QkuZ4x/PhyZMeSRRAJHbxysvQzl6AZX81Wjgx+02bO9Xr9aqs6h3uzjL37jIf9VX
wB55KXbYQvdqlxp1vMbEI5pVFnrPOLW9rCSCMiSXByTJ3Q0phOBCA0ca4lly4qlQ
hcktia4UUymbziq4GJsbCx4Vwzd/idddTjbSL+dr+BOdoTSdzYmE+JlOmMTtMV7m
UfgjWRT5UFfTKWyl/+lDNcXa+fnD4iso5yy5VyYCyWq8XrJpZimGUlD/q1OW59vy
ieEBLVQ/ngJLRsuygutGSCRrgAx9o/Ebvxn9zS01g3ukz/EH/c0fuWs9aaZtSMNS
E1siBVNzF5QXhqNFvT5MY2s4Uoja+5IwhWCG0RSlm2HV+giGgubLYKRF6iZVoHVo
ubzKGpLqyHxW7X9kmbXXWtuNG9BrbAB+oX6eigCFlHRVW9fb7KGFE77q1YVBruyT
0luxklIq8PMB4h2gR9IrqWmygFb3m7xp7wx8Plr9VpS4/gnt7HxzuS7RMbVozi58
fZENIlPwwMayg+6IU7qA6fE/reDIqsLApkONqhvuc4Zhlmw7+ygBLT9GmQCFVJiP
9I+16MlYuHAKlVaO65Ch5uiuC9pGhOvwlXpGXbet2+/Y4JjVtptqrEbCMN+7phjo
nSWLb763EYkM4FJOYZ/MkhXfg2YpP4x6yqMYLdzFiV72br6ldDLfrNEqrwWTT613
iLU5gVFYVdJv+iOJKdEdUjb5xBHhkqmxc5Xh7yQrCDIRwHmpeJNElEWMuqSxsS75
65vzG8VgEmOK5q2/k7gLxR+VVNWPM7hz65uCebKgDaOTihDCWnIJlc7dgG/c29bZ
5a66ISjyvdsi4ikrBy8Z5sPDiwDkv/aeWvKZWx30rHkpLD1q2zCjFDaP5q4c8L+f
5grBaqqV7Yq5vuB9bnXtsqcRsDJUVAPA9MfrHR0L1loJrPwPZjXFB35MpGvg3avp
6m/VhLm95qwLHtEH0PGz1K9bhHczoR2X7rloZtcTBlTb3tSObPxkbdDdQAO1xtAC
fCucfC50SJlyULkGR0DzmgwDY+OUd5fyvVSKvT6W5ORvCf2B/vlINIBH21MfQHId
bXB/nPG+q+sU64m2AfZTAp4S5CPiXGkQMGo9VKaY5y2sn81SyMTHSO4z5XSwDUz1
l5rjMU/UzlA7g25FZZ8DejWKwLNTQQm50HKJyY0BJol1ydq+XID8cNaAFBUWIs/O
rx6E1XzKDcaQctBzqo0PbXXSl/njgoqiCWd/N74NgQKzZmOpldWZDoM57Kp9ZnKY
E3KRHlg+i0wyi00QmUCoF+8pMSlrhk8f8JRMAFCZtNj4+k/8pkbyF55xJ4Q5/2aO
Ml+PS7y1hdIC6flS0LA8ewjfJTyjVvEGKK8q5Kc4WVe1VLnsNtzmLcoD2NbYIOep
Eswven7I+5SP7PfeQ6XGSKZYCNJQ54rRwDOOY7BKc4hbejlLgiKVQNAxNPFnzcHt
1lBnDgPpL0dqFRXiXCjmfPlhSB0VjSYjAq1I+vdCRwFyVeGVNV3ofxFo1HoJnGEr
/lVJ9+ahgzVYLDXOrq23Ti9p/3hdSGpCcIWkqFUPljpmiYKTfnK3i9DUFrgCY2jO
Kd4FRzzMCYtfm0/n2zHFCg2aB62+VItbXbvYDnz4LRseBpx/LAqhI370tVhuPZkZ
9Eg9Q9XhhTG59Zw6W8rkhK9a16RWbt9emhHt50kGgsVpJGH64yGIC+/BAjY7a8Zw
FP5wnubuY08iRMk9q1VO3KvnCS6q9V89j8Fk+wIKSPNOr4orZrwYlH6otD4qlV7n
N8zdGC9zVc0tJzDN9PpIVkD8aqeW/nVFYNvPUYRPBevm+PjBtgJY3wP6Ol4Jkg7r
vaLDES7SgR2jSFazT+yWfAgJKb/2caGYDponN135v8E7JWr1v8UADOMFDhUj0Q1u
mQXzwhl3a4U0OfAWLIkVkjnOmU8DrChiuAPgBusbpyvYqQmh7ikOcTiRoMTnOBaJ
bJfGE308jP/M989Z2k7rPx5jMuJbgOXvrzt5AZUOUsJodIiqPKqBLMhKva7hrzGg
WtCsyygDZXZOTRIncGddGe9Fo+UJUP6DL2we8JLVpsle46N708wTaeXscFbruKt0
gr5+qDr5nsNAUtVV0Xvx9Or3gpb/HTsHReYdcg/NsmF47gbUMNM9/tw2PFGRDzSU
N4eVHyPq7c6ddwlsGWBxijm3vQh7mLDxfUD8A/n8EpqcZGfbhMrkjjbHYGE5lKxq
y2q7Vhj8l8Qu78eWiYDzzVsmeQ4KMKew8KrdNeh236AKAdCoJTS8UO7dwB2L8k+D
1ooXrh1VbgYEszrhC756fJLhJWHcKEgL9E0RQBw0IEGETM7ohyfCMyR/zod3toFv
GXwvzPDf4IlOvKi71rh2PNvBM7ud9cGL4OO7sNFsWH/YxaYZx4ru+d1+r5YUXTg2
V0oqq7l8Z7+isIuIv5+B0Lk3UTHvwl4ByhVcWfFrjrDY/XQkG3Wq8RYfzFDILDjI
yL1EuxL1h3mk9nQxcHx8fho3R1UzsFRoTJwKg7MCv3CQZZvHZcGQp0btICnPH1XL
8G7LHw5grukvpgYuClgmLjMzd5VSgbTp8UMWfrRH6IizZfzRefaGcpnP2tf8PNKz
bKkTwzr9xweZ9pkkmV12kJ9gUpXMRI/9qNEOJAcvw1KVLfREXTrdIk7llL1Mw3z3
BSpwDTyxf0XJQ5mASszpGuTK6FjhzsuLx7zuqBBn8DBFDdvogkkk60BBRacAkVxx
0KNfVqbg0047i9u0/znGeMdV+QpDmxteKAqfn1NOx0Azg7+byrfVjKhvvMorWQ7k
1upqkTeVwt296dREc4Zh+yrCXP7twknN1PiFjRTG5KeBWxxonkSzyeJpRW9J4ToE
miTzvQCrU9nCDoIQ3s949c+oh53egP4PpIjzonrH+cDmNwrqRJfo5EBqTWtswyo+
qKRUgc11+MqPBMRP/u8dZDFwpVir/3lO5umMuBXRK4AWn2/1G+R0bKuq4WmXIoem
NeVBB/gvoShSa1TQ2tedYCQiCHXPwuhVhLEAVK8dqPC4oXtegiNp0JnDhwpwFJ1/
R+absiymhhyJASVhVX487n7YY1osYQ7HtkCqmYzkZXkIZKKsAN+bLBqllPLN5+Ro
crUsSdEmDRJzE+UIJAVN98e1lX7rk03GwCJ0u6qqeNVJeD2eiKc9JW7+xnrmCnSN
sSMX1ATJ/VA35r8GWWQYUoee2SUUBQvqUyRjT2UP3smDSpF8VYuMEDnCH2iz42H8
04QyDSyuahmrDXJmgTX5VQMgNx3gEqqPFMwHmlZ1M7MG7ltMvvgeLbyq1TRk2Bft
LFEJHN1oPC/fCC0ZwzCNVoDIA3B4OCfpPe52AS5uWpPB6jqcYuqKxnAdbbIRkr1/
rPVB8EMOoiFIfMTCfO+Aww42z+2BVanYrxVqm20EfVIX5mkMtcUOphdo/JqdJWjl
Wclh8hG9wl0b3FOtNhaLbO7y+o9aCRVcCCyM+74XPii4fWfNv1o7bkj4KHJrgry4
T5x+e3njXxeJ/NQCsw58YGtuc5TgppHHx7NxcVY8IYNTxku7nUAOX1NdRsH9HGoy
WGh9Izr5qlvZ/iPwR8YgzGLXbGmpznWRWZRyp7HaJZXCAHEYcQsR/azu3VTb6no2
+BxrXFoiyBkEoxwik7EP+OwcycSaYJk2DiyNv4ch8v42JvQqmMRkWC0yARYarsMn
tMEtEqB9r/3QtrOi0tTKuKbFTD6sfeDzE1+GQ0LyZwG2OxH56/KvpNZjY8vj8YCp
pl8jycMBMYgmJeoewdXn/rKi07GSSaBI+KMPTh9yjg7ZMi0FpSktMYJp7BLUiK6d
XEIOSjEqgxI8bh0BEJuaZNGX7uMVpAZ7MULbYqdojGTvpV83oQXpLTAlwZJBfvc1
gOhOGoZM/4nwWA1alV+hMBYm6mzDSs5ISWNKjK709ZCXxPvfTS3Po1eRiYzOBXT9
v8QsSgQqnzq03xmM2MCYB1bqsq7P6+lAHxmCc+Xblqvpc2MQmrd4flURxTqO83fk
fZcOFD1BdUbkQ3u3vMlrvTzXvyHefPFpU3gDU76w/giicWXEB7GvXkK5crcOlMnN
UVb/6zVqMteH535h3OAaWPursUHi4RXmo/awmOsJOuuTjm/jX/9+Ri14JO6SgAIr
gFbXpAZzHu+1h0YH+oa1oGGadLNQJBNKQZwlsu/1+/LKpWpiwtcKFSzP+i+dWIAP
2uz9Uk7kfhbEH/K7ThFG1GrGXOsBzPT4+lC8sP5PrK2rGQCwtAtvlVO8meNJGE6j
SG+6XgQPLZh4k2ZWyME7c6cocVZTEpEiYeBBtvQLVs1mX3gF83rINwsEr9Yu4eYb
FAFgkTRPIe/zVHwNWKGmnzVBvP08qbNVQBsfS2x9jBJPqylPWHkF5La4dxU/0Bvk
oBMi0T8+qQnLVUejuIRHKxdYSCs8Cj9DursfzBpw7FOfFPHBYDHrSCwWQT+ro3y3
GiKuZYz8kVoZTFYkYWAA0gHS8FbbyIaXsQfFXToeWFYpiE5+sqt/JsAxp1SpHmq3
nWpHP85FfK4c7HuAUq9Y6BqLHRBozN25ZSi7GEZ1KJR9BJsOdvSMRa3I/tLG+NAz
k8O/i5YKWJuE3dRYQfQEmS3CM1qEqWxAscLLlkL2Iv7l+UEiaUxMbFLyGWGszQOz
QsaZTeZ63QTPGPApAe408Ujbn9dAHbWRmFGm2XKvKU2wQUFUvPn2VxwhlBm3SQXC
Bmr7iymb0T8cv8GAskp9ZuMMo1ZyrbDN/+Ex5XaDE3JGhlzm0lWwKRlSLTWo/S3R
vmACYQlc6XeijQ9yjIbNb/RI/729mEC2WD2BV75YwjPl0+58iwHd2eqdVYPDQuBW
Fziri0poCkkvInoj1LaudrjBWkETBoRa/QY9LO7XWOuiU8e1ftreZIYsnHnd3K5E
GMzwi4mxBxSR1TLWSo1dWywlf+xSexOSzJ0K/cAwJq2kJjReq2SkAV8kBadfQUf6
aO2qUc5nVFh7NIyNHBec3HvFvxUdYf/KxFPU1XYEpjTIg/5De+bVbBX8JamlmWNL
OTbvPRi34OwxWCTuUI5xHrhedd6XOdZhIKdOhBJTlj1GQLAm4tuVT95B8azb1VFO
TRXVfHJEstnz/+pmrETBFJVsZpGllecYXYjOVuq5nYriGAdESicJJhnZYo5dsgdY
BQyup2hXsjPsQch7GftwowR//DWhbiKMoX3TVNwkwUCT2bBKQs2oeceG7yDCXhHD
L04BogDAwkeXqOBLH8awVJ5kfHCn9O9jz+TAtoEvg1lu+l0CavlahQEeYihdjHnj
BgFP8Iexziah0IJSQlt3jbQSgYUiRL1OVpxfPWhhy1K3mIKyi1a3MDBpWkeLFs7H
Hn2hT7muM52kFHMIMh6q7qSgCJaorkBACaYr0mJitHxjwj+mduGYhWDJa/0b2wgK
VdDXqsdqCJuKW/1LS5N9UqZtXyO8ZdcovhHMe9q2dnht41ELuBAjHUG6utyXVzO3
u391YIcKCbmSBXDcjxtT91hhqq9qJCrTdArKN40w+ik8hkH215CoDU4wPWGBteVZ
TKSvB2oNAceIjDlYJfep8ICTdyDEBpJeI7G2Ft00AsQob2bzRtdmySLexZCDWgXK
MCo+H+AYRSHBor7i4B9BooJAuBllqAW8nTBSOeSyPJm4yvZdmxTIluYU0zoJqkMz
mwPI5YjXGaom75ph6wqv8v/ui/UQuMZwCD3/aW+8Bzn4o4t8mAVQbN5rFzQu5l/Z
6Sy+QwcjVP/C0+vutAjBGf+hvHU+MDkM32Hk2sgN13yx57ts3vtq4A+8qluNC7BH
IeTxgV7msD5XlD4enmlnIyd0LWzjBca9wtJbtjkgpwKcshWkHPuVzbOk2sT+Q9BY
Y+rYGeB2sMMlGiTE4VAhtPQsl4igWWKP2AyUm0eluU8XjE/z5/tG45lZK8vPKRSA
mO8Ze025nqRmrU414oCiroktI7ynLjfWI7ycOhHXW1WAgOE4rtPQpknHpXBZLWVG
cKateP45JzkS2PFUDMBZEexSt6o1PDEccJxp/uyFKCsU44HInYoKOuigK1wxckqp
vfFbKiVFuX+3TcXbBW9Zh8G8zDQZPdzVL2LNPgUr3CoQz+fbF5mAMT/HEjqQ1JED
UfjspNW7npo63As1K2z69NpzItNb43NSRJGSzTL1XVjCjKJE2JHjxRGBcD1NNolE
RCDoDFCrXHaZ7UZ9MqDeut7qdYA149jDQU1m/avO40ebdOzzwWRF3WEoxQKBAO2G
heeDdTF02+RC9o4RNzy6iRK4LVIGZVPoA6ZmGsdpVRlfQfZxHyaylSoEwqC9sYcO
QRCu7vajdnGZb7Iqm9bLLmw2kXVTv4l/DtOaT/rl7jcRmzoQh9kJ3zyx/rNpHvLc
W9ZQoHKL0n2eYvCknTovrsjZwCjO6UTeiOhzIQoHPfNFHy7thCtbf2bVhRGsjI1m
OfFQAvWEoOf96spbP22/ulNiN8xXWb4zqLbeqpKVKuPLsNOSbLhHQ6k6K+J1JluM
uh80Op1uwQUYt0taO+eDZfVojj/TYSFlyJlSq1nGCIGfvUdn86e2iOHBCGXjuuf/
Cq6hLARdQWewO761G3rtsuAvLqTIouE7od/N6sFPc2k41jbCgkkQCDyUy+Xd+O21
oMpCT3y3xn2y/Tn40SO8mMkhtbCPaLxwD2RDuvyUQt/rf/mN2aSoqj4KtNPDfWwS
FEUuGqxQhw0qd4nB6JIGaCRNK7UTX/du0JyF3lirwLW539EF62G1nA62GcdSbVWi
fkw1eQP16MfBue0Za72h6Ic7r1vx39Ld2ImAtDnQ/WHvvWBXCQUgdgLoGrb8tSA1
KUQarL3WK/wKfQaUwSJaBLA1aDKSGeDEWgAH2rfx6pg0ELxYjHuK5XrMmhw7kQ65
mvEW7jLqcLEN4Y+v+1Wvukh2AmJQRiE7SFyBCsIjGhJICzwhUTnM4RaKVxsQ3pox
QTkVD+DmWE/IhxhRM6sOcfX95RRrWc1dhTWICn5oafG2d10MiJRzA97oKwtPzxOt
XnEfAIta/ge44BXr6MZpawrlR1g6WpT8IRIzeOWVaIVWzcYn3tSHXIbbU+HXlFka
c8Zm2BG9NTBpmz7CgKeO7/3vv9+LzZ+t5G4f/zAmO8RJH4AEujWjrLaH76U+1Or7
GBzslsD0jhsupSCbFKT7KvobLZW1I6go1mYjBQ/W0tejO1wbkNTFlS8LGYIJ68KV
DmU3/1tldBc6TqqFV3U3lpQNoSRlhTc/2JnvIXOPr4R9woVXtraL95TX/y4EbWyb
hlmfyF2LgyJTfAP8llm5r3QIFkglLF5XtbcNwAS68tMvRTICVIZSUvAjo7w/NMA7
WkXeDyRu4tAk4KK/PLtwYzyZ87b1axnunuACj/klO3ygF4Mr8x2djlQbKd3B86OT
L3cn9xlluHgErUfXbZ9N4FdcB0dlE5RIPIAXyxjops95sQzN3ZTig+vb3R8HNntE
UeEo7+hVtS1jA3Qd/qpA90F8m3e2ImbmPCQU+7wLkxJNSd6LwpNcgsfmRwEYQgyc
DKdmRT/Z2jKWberm2mYkcrorK8JZDs9QRvJfshWA+toXujPi6ggigkREl5BIUZpq
pNoV0nKsecKceitm8kCKYMM3GErVd6iTgCKc0dmNwMkDz5bSMHYe1mM8g/x++Q5/
yS6sgEZrHL+IH3q/euM3YImJu16+LpJXHyqTZWL0fqw5mjWuGJSrTcZu8NRlE/WH
Be8w4OCHstnQE5j9TQvOllVk6LrhCq2ag+gFugOsYFwueD5nvcMCdAls5nTCEig4
pBveSJ9yugoddRvt5devtswJgGpWI2rjC4FWCcjSJd6VQ5N7YT5U6/STr35FWAcW
La5oL/uD+bwVNPEqKl4UsPYgisXtNg5YKKp93F2+JbQzfwrk0+PPlcq8NP8FimnR
xWEYjerYFpiZMCjyM6JwlhCaVpXmX7Xl5os/mwHfUDQNKYUnSHVfGM9geAVkVjaP
0Oz67YucQ8heH8sW/LvqvgnMN6zrB4d2NXeDjpd9H2WW9Wq7MaDh07yNQc8xW+z6
aIBrXeahPEIU7OgnYbDhKrmhmLgkEYnj5mj439/s4WWR1Yo3jC2+ugjJdgRDPSYb
H2D4tWc44ygsC5dwH6gR1qDj3Jcf99r0HPZ67HBN2oETKDUsRfxmUZyR3aUiegP5
afpaAsVAROEH9ikK+gruMqf6w9KcCzElSgvzb9SkMxV5CGQf+hJvHK4WFJ4cPd16
m5nr2yvynbA23OtNRTib6octD0gqD9Wy94hHVFrODrwpuqhSnGRcgU1MqwpsO6jz
k1yzCIURnOAkKOccjSpcLcR0KW84kc8dm2DcUpw0B0twoHwMbwtK9FUxyXDaFA/e
HKeVbfIs4MjyGp2B7Dkbh9dm2zR7oAPe3dO7J5xZgT81LExNhEiGOvnVR99ctO07
Q/qhSUtZmtNlVuoA6At7h/eOvEVNoT4OxQk6aZaODyJVC6Zb9ZwL7AxHYvxpHB+j
5nDDT2rN+aKYWdc3lr4mIX5ZdFxGVBjssrRsn3NXdg2ybHWvxyUyUdRl5W1rjCaa
pYDIdzuGLtSGYLRWbAl6setlch3txteLyxk+pwoRaxVxPv/IFNdVd8zqkYtio9Y/
Zdt6LmCyWLsXNxqm9ytcEsw2WONrGvt8vI29/s4ilq8hewWGK3usyutF7mEx8+z3
opaO+urJ4kEgOrpzwn0pCxuXmMod1c2rh5NoGwoF2tH6y+z8kTDO3tyoeaKa6eXD
vfF6CYkrUEf3cb8pEecDcYsX70bAHiVgljXA5NAm6nQEnTm5ipcp70PePmnlWB1C
ONd8WqHmUsuhBWXZoSsa6kp4aKmbiBlQBArOGkAyo+Xu8gMjn5F6eCe9LDqDBHRF
xZCzLBMuPNP5VnBpx7XU3j2spAH0UdeiL6Nennshhpe+BY1foyJZ+UgJRvuFIo62
9fBr1nUT4wVCkQJlbJCZnAu+I6ununIw/hzhJSSXkQL3Zeu0/MwI2XlEwWESeVd5
6DoAOQrgm6DAS95Xm6DlzCpSgb3HsGCW+Uf/KtVnc4H+M0bEU/b2JJNlXPPuhKvx
BV4Rrl9voy9F8moM1kMLaiR5vr6yWqyCYQyzm9D13YjG+v773r7vTXDVFfEXVztZ
a5E+3KGWPXTc++u6hftUjPnTojECaIA9+B023UIXXyFTlqMMLgR1Tnhdot8By7H9
G9WEHQ05nDsdcGfJzc0AQ2Qw7yDfq3qHjyM1UCqaSQnah5pMefDEg7PWPMnfNyGb
F4cYkBFuKzi3kmJlUnPNqvR75KQ+zbv/EhqbHwEoTl4uXKm5mrGbV1HLLQzqgZPm
PX/r+OGfqiHt/bi7bUaPWQO/r9R6wmd6SUUYjC/KET0FEW+QNs//n3LPjsf/8/Wz
jw86pUqm0snoLCj1uXZexDLex1MTX3PK6WkvQGlvtQZMBtRHZTTTIydYMK3PRfi5
KfBk4jjprUQo3onvVGZqjxWm/V6h4DLouM5RGQmCZlpMFsprJqgJbol+r8jYjxoB
U34TsX55jqc90gEI2/uT807Pn5vurPwLDK99a9xTJa2j7O+vXGNIpNUSuZv+qE8l
XItZdxGJmQjsBSqKMc27JhDErYpwQsY4kWvlJluk9DUQLjMtcDZAFy9L/6FBdS1A
y+p4ib83sf3MKqwRsnoCDFbzlSDkkEKvCa3TI7TtSd1Ic6BbsFSMOtKBB9ARVf4t
kEnEJEgcZeXlL0GAPMbw2KlPwj14vtolbGh71ckd/YuCs6qs5tI6v7L0zeKNe71n
HumGHqi4jVbJPIzmsY6Z3cbP27i+eDYZkiZflMRu9FvQ4xrVOB/9v3Tf9YVjhFNd
MUmk5wI5GQ9OMMQYyWC+L6cEeLUiPTIFr19t0sDxR4H97A8GQWGx4tYjluGLzKF1
xR5Ssn65Yr4rkJnDi5bIHR7lhZuGZmzaZGsYVPtV+HsuhlYsVMEozzFUf4MI69nU
Ny1VmB8O0UMqMrLfj6sYSxUTuDFA+YrfWUWRRn9sNxD0Ggpc5n7dYfTY223+txDW
s1Kcf0Pt1RjuY4I2aTWwcVIc4wog5GrJzJM2fUt1an0dkygjEpWbBD+3obBrv4lW
Bants/WbAUwv5e0Rx/qe9sTLN6xmKcAle0sW0hQh7e36lTBQ8eG/t+862JjxBGpn
GVR6p3N8z9XjdW2/3j8C1QUwpB2iHgyM2Aio1ralVHBTCdTB7v1+trRpWJlusdw6
L3OQmyhmg/oors8Y26RWbNRhAZEfeCtWuh+W5JMnSEzWamefIejvrOykQwKeNDlF
psSxAQvTyJLh6LclfUayg8UKL/0JMqsOkJ5xDr6h9hma+vW/vBRXYGdpHkIwjt56
3snhLw4xRrzGi6XfWSu4/5r5HOF2A+r9wc3nSTkWquI/epiK5TTkhX7UYbiMX520
maw5SJa77Dw5Gsn+eZ+1FxqXCMD2MNuBJoA40VxW+L36Efu/EevfMX6BytM7oj9R
KEBnhda5I8PzKC6hEYGUKMZ0MDvhVbzfQTnK2SDi3fM4Y3n5BsFo0ejMyp2Nroer
vUuisnkBu0GL9cMd6GQrF4nxr/diMqyUfWqwy/b4zGmgKAtqau4+jBTca4wDsl5m
76IoJeLnqjdPcjEb/kddpII6uLGyqq2a+jvIGZFeWtNwUARKa1pPXyQ5kEFfvP/p
UOj5xTF5LdgpJy9k+9ubNIZT17WyahWq4MiKpu732Y+oSrhIDHoeyaN+jajAwkcX
8VfIEXvwjU191QlIV+roF9by+JzlW0K2YCdxFY28QXFH0k2wwUuWry2CPcB1nbh4
BEjSjQBm7Zwpqx6zWKlxPOyXDgArnSZqx1sqN7JCGK8SOTgzzOrTlcpD4yyvBoKb
LD3EHm0MnFaE+C1CHwCquA/IUJZ1Nbq3pW8hKZ52p3F1yh6Q25E71JpqnYAw3ekU
hXSOb89qDtR8atMlZyjguZahNpWyeUWwYAVzfTVCAdCuFcBMs9lQlKV1sXjqrLN8
TU4JYMSBKMcXZ/N7M8kI5l6Cv1kQyKTbYvFeqfXTo4SxKSJuIGForhRzL2kW06Pf
OyFIL8fp+skr4HrtZqkiLiRhAitvTlJi5wg26WUUXst6jiOTmakFrkxzGP0EZDkh
8Dk3cU8JbUKpZq1ah1SM7MTd0kx2DrJ8zOaauN+J1GlzsiVqKKvRC3MIYolrMqup
iYm4mduu6jcvAJClr1YZETUE2XVikcZpYGj4azlN/vKk2NRlYT+H4QBIt6SlarF7
h+HOxFjiCf1g1zorJCnOcg6KR2i/cE+QH1YG+qLiHVuqu2SRwj3vI4PFPUcBpDsl
r8U5Y1DOeR7d86o6n5npH0ewNsxkX17AOrtgsCjpFLxaIFDfIG5uKw+RqmrVySoU
ihWNbf61xPvEPKicFiGU5pJojQX44/zkPkmmnmrO9YxV7M4OXqF8d7WStNSQ7wnS
xSNyTC+NqIRo/CPiVuD71USXZXK+c/lwL9xs21f9WjHrZ0zizKfGa70JwX4bwpI6
3z+GIdoabRmcv6cv4i65oawqopEfqZfAAvYTmWs+wWP5DBmlhbpspaUVdI8H4mR+
0eGSkbl8YBY00GFAeOVW+cy885SqYKClv+EnV3hQyvgDDHWgTG53Jd5RA0ZcToYk
je2XzXXBo/CTg+rP6Mwh2Nmt0OoMYgFkYF3GyQx/8j1KPAf/nJY2knkWFLLhKaUz
6G+V57yCfcL0dPJ/gEgfQXBsA2goJTy6SaYLfUIk0UhHKd3q2ILVn4OhsBqcRyse
zFdG1XQKplysAHu+iha2cRp/PFoXtSIbeD+PuuB+EvjeBLhk0OcNrttisAEBMr//
+5POUlnbiJ81WU3tLVV4U16SV1edQ+Fc6SGTeWqHAw2IfFT8LWmjYpHF/JVv1WR9
3ixHmFLflXxsSp42ItKMxguX9jJzf2rejfCfELOF147CYdRp2mylUcRzRETLynHz
kbMjrWxxlrbmE9htOLw6m57iM3BbTXQRfzil04bY5Y9fUTNK/Ts0haGnbrzyJjXY
WuoxXHsllr+cUinJD8w6bPAUnsKgMgfFxOmgM2IIubWYOTo5TyLCMflmE+A6I89N
FfewBNTQwmZnOawYHNzU1ihVYiDWT8L32H2YJ9+gcAsAfJhRpYo5kgzRm0gkC5m2
/BNoci0KlglDOWXHZdgxVQP3qO2Aw5MPsBrDXaAmdn8SI8FGxAflpH2qpTtfnhmN
B0CvVdW3Hm0g/vg1D8Lu+jmBOh5JQchCr2HROvUuSS3i4RLckuqIGLnpAShnhcWS
Udv+2fkxEdo4THlS8YxTFV0ChidxLRi6txQIW/4tLGY3/EsCVMIBui7NK8Mj75zt
paDpc/6SCqrB+t5bQ4gY2ZasPrwKzpKTuPVLaYQp6+uzXueyGwumo5kEHeKi9b5z
dxdGxE4MKeFQOXlmAelPsFn0928ykCFkRzG2btDQVikZA9ECbSjRDnxNDPVD9rRS
C63pd+vkAKbQAV4FX0Kl1elRmuJwv+76MJBCOCpj/1d6/fY/OokIq4cPcEy8qqAM
bSgLCRhOKHy043jkUfapU3BFcHloHh1oW7nzuvUpCyHa+BO1tzoH6HHHTNhWzaI3
e0G5DmHg/QKeWBBE67thSgLX93S9+HqWu+/wkUxz3/FnbZjfs0YFk4GZW2P6ZK2B
mscm83M5t4tabNkAURcI6OmRWh+9gmq5JQhMNRiQwJUm+uNXMDcV1R1t6l1Pn71w
83fmygkrR7+wYu6WWI87BysWH530kcvfS77JRJIfkP3FpQwKps+E++y+iSJfrt5e
qVF7O7RBgsZNlHNyNCIMP4HPMiI6nZv+te/tsm4yDU0ze3KE3eNW2h3mvPRTLBi5
WV1kjEALcm7FiehnA+HViuW+qfWwFQHOLexuiZgq1wO+lQBRZ7Ur80vbBmdIGyAX
vx9SwXy3zPoy6sUmHSZp9Oqboc5d+V0A3CPFc8fD0UPMD4old5DsDN/ZxTQVh44/
3cMqXdTKCzKFwk6ebT7GpAROEFNp0VSkdeKFrz7WIJMAI5TiusNERUrexriiFcf/
b5B42eTJEjJ6kk9uxCJAF3c0YZmEpfixA/7kuZSEd9Ezjqfv4FMrO2D4LzU+evn2
TzehiLzt6U25sWfR9jUS8Bo/4MpmxlIkAoIzqCUgj3SbUG3KiHu2MWSq2r+TiGcQ
nlz6gybMD/Qw+5yC6xiR/siKT3Jv0+vNQw2++I+3/5Kby8Py4d5fazQgwMxhJeSs
Z7Xvo1DfYqSnjWVa6y+FgBXMu6UbWaeVqLrxT2dUnhFf17Y/wc7xpNKzyjm/D/yy
XgRaZf+FlFMDJIrPVR2tOpANlOI2cfazN4TwUbOERa+z33bzVNQ07JbHy2TyFgZi
7uTU30e9DF8UwJBZR3l165DKcvwBl++ejt4FF+HbCH0OuhLOjiGZfLCWIMeD+5vR
BAXmp85qtbeDV3XfEvm8KfYgLv6QaMb0F/YR8hsY7BpxmPMzHZjYPsuwWDXgJtBj
l8r4/pqDFhcJ13nITC42MjE4t8RWIPc6MVV+nvXk086uS7fKXBHIGproIwCynxr2
ebUNnRKNW/suAQ96knG3VIbamMQCgbcZaYHXXcxMolZb1achP3j6V9viMF2z/QeC
Gf6DwB/7J4MRyt8xJ3ZTVNWzrMPry94nZQ06BzLiSUCntgwgZj71alsZvPWWpTgg
mpA/SBY06kEC4A8x8+U9Rz82/8/5iejGd/Wu6wUpf4jVpf6vNNv4FqE/Oe5BaXzM
R81zzKs51XSwUOwRyaSSRboqT62mXb/D5Mh413FaFcIQL/MDjp0avP3rFORWr0Zp
KEefym7YQHOTAqm4erORnoMvEUxu3t5KfxAwc1KqOYMcSrnCHLHdeFyWjnvkbhPV
Gdzb+C9fZPcsZ69s0BifPH5rIV6fvYmAtF+DUbkEJNdmU2Q4p4yjLvql/THqAmmx
dcml8d8oJIKUh/v31/eFyREqWQTHgO/2a2jDiw+ad+3itfhNWeq4usf7NDE4eoax
+j+Eos8RLuxubmJ6hCigRKsvJwOJnROA3zw5XTOcXTLaDKEb21PwAjXL7ypciMI0
kzp73O4GRmykC9vYE2CqhjtbStf1C5ZHw0KGXYfgJ9GB4XCKlzmfg6YkXgwE3ZHC
KdTiUdwDRS35y/3wCOflHq5riexdKiE/OHcl+QHVAk+9nZTyyK8rFdcjSxkVs9N5
ahqf9xddYf9Xec1lvqDxqVTqHGy+7kQSo72Omjc7WhDHH4XqIatHV+Gon4UxLC0D
vUlDJI8q/7Ohgw3OoNhLtOjrJO4uP7LD6FzERnbX3i4AlB6ByDctnhUonmhi70iy
DNjm9yS02Rv+hfUlif47DmrlELH7j7OeIQWBvj4a7msLXfqF4LriU+ETJrh/9+O/
VgHRQMb/FBDQYqL4xbtufH6EPBqEDNbTWNp+4e8F8nIrkyHrq7ugVENK3dIyi03M
E1lPZ8tyLvax/kNCMz7YsqOGJhWkMzWnv1TdGGzLAe5ADnCrJtyQtNmVuhY2cn8L
poriXXWwM6Ugf6YKTb32PF91zx9PqWekzGZ1U2w6lrNSdUrjJ3zJDNLoN/8XGhus
HZxd1bEWeBSWDzXewy+IZXUStFITmZlP3Yni7CJ2UU8+vzMxKGxzeOMIv3owTCah
F+ugSoBzldsy0VRQvpsiKWIwLs+zRj+DJAYP0nGgS0Cteecsa95HCBQsQpNIHyjy
snZp1Vmbw+oHJ+WM8L1x65nBTZZVuFUMYogpelgiYgqF7ZD59kP7zowA9T864d4F
ZRplAttbYVVxX71U0gAOew+5Ku2JNnfX+86YlvJZsoUbV35N2+RUe3TX26wIVZVL
06uNOEscdSW8s/vpJu7/yDTDi2+CqK8bNNwYgXg4V1m/CEGgui7uaRLF6zFfTdpB
bj2eY9v5dyJD0yzrsaU9mXbIAeBCE0wIMxBdXTbgv8Aqojrld4BRVhXP5o6+O/pv
Uu6lQW/Q7WGdNjrbP2urgR14WEcUcYMA5jmr1LIJw4WfR496r7RoChSYBJWe01NS
uysl7LXVgShLbcWIN0PyB1nTHKJMAZL0WFLT9VbKF5gqAZXMNzbx1PAS4Bayc3b+
zGn3FgzlSV+lLLKgAOsU3be/slRb370570An29O8kDjV2MQiXh8HdwiqDbXK/Oi0
STr8WJCLLHIKv0XmXJEe6c2PAp4QtOyI12z9QBnmGkeni4EGQtMBFG1sFbNhQOiN
hX5HkOFdu2X8o/nJO/fG922A4y/hvYOkezVFu1+wvQharapLj7Jv1GkKyw87BMwE
RR2r5kcGn9cpro23dGXHqX8j5+PW7XIt71eIsb93aINpC9YDjkY+wfYNAsoaGbKD
e2Z62iPIJBvS1B6HY1kI4A3ENcBSStjkwtCPxg++EgcgvYNPlkN6IVqCb5tdYdzH
0xknZedDevpMKwNaBgd/bCVk6oNddSy1HATJgYco8b2L6ZFB9uj27GH0V+RCq+uO
1SKXIyq+lXpSfKQxZ2vSqA383fLVDzhFDyqh8vG/1Wmpl5HpusG59C3jhe7SB2V8
uyWThpJ65de9OE2qJq9BztBoodD76qlNUyKjhqVzx5U8S9EVIpz1yUM1SVo+E01w
JFVH1z6yKAGZ23R86dteUtmrGA9C34OB6cW0or16m7ELbKrCn0AH+SKdqDbbTajE
Naty4E9ew7YEHeOUQO9g+L6GqaVWGFZE/Bu0WMEKTBhJuSS93WBm5XBqX8hGoiLP
P6UfDPSSQYO+MBFtyk2RSqyBoNi1C/AdWEfq0s1wu2quhFZMusJAGEcMU0HOyu5O
et8n/L3DyZdnwrndI/niZiNrZq2SpgXJPaUo3ZE71K9KjWTS7tPGQwWT6svyarUl
Qa/QV1ZcabtP3LTWSkmFUEJYn3koDWiRxd4DUlEGEXr2+IUMtrcbrqd3bFrE6hjQ
2Ta8QvyzhmdK/9qxpXxxEalS5dOuo9841zRANwncHuk95ozwPaSdbvPZZZ6Z0nOY
WeUsnzJbvJAhnmgCtvg8MetHd4Qwq55Gvni12fWFKd2FTzDTgFUPJJACavfVRBjx
WJbW9WpCDB2XvW6UJQoZM4UQSWQQ6oCF2zZNkOsv5o50xEFjQpME4R8AGuU6RCus
1Hv3laEk7VaMqfcbouPBVuLrwOcCk/yBSl9ooMApyMiU5IOyvkmIUvd+ijDlUuLQ
vw+r/tLC+AHgRSot3ds6zW6OALZJtO+dg0Y9aG3uCx/6aNfnp2f2b1u4yEntOxoX
9HGJNMCg86evEjKCoS2JyS639c1FkK8CjO2EBFnHyo9Zp4/GYpdm49e6lYBf5p8b
fQos2jyUZBXmcqtpKwP01E2QEv7uKHN7FfV8XijFw4NSIukh0763s23nbh6v01If
pryrsjk5iRVHl+CTfT1fZcjTi32JVv4iVyO2uqA4HZp/LltVeKAQkxT0LERYm0cB
SchWMrLuTLRSw4LmjZENbTuUYlFLbaEXQvcHdA9NRdmtnHMa+ZASK1Xet0HNlf5E
D2jmHNadth0I5yy9QkblWNmJJ6Aw0M4ckDJH1edJw8ULoAqHQfkbYad7DQRFLkfD
xcKPcopKj5dYYX+TOIHlx2mwXPgOXVzb0zk3TNr3DHevSnUfn1rZX538mlig4dv4
yMSI4PDPBs0lk1mLbwlBlGdUKJgpJ8SKEDumjQth8vT4Wekn2bgiZHQCfuq57698
H0FeTfwS4qdFfiB6xSViNy+Zu5HIA64yztoAS+Q7U7yqOhuReb3lwJlkx8S0npyI
cVYQvpp0vBHxtqZzj/alHWgwVEXsCvUTXTbsW9FT8iZxjyi5unV/w92AABDHd7hL
C2+FUaYsBxURzKqc/dMEu4C9CwLuve2tV2ChruRH/LIwpRBz0PaLINe3RjK98bKk
5RL+s4Ufp2kxj+VsiIh5Sa8XpNoCl6Fn2ehYk/MABE7L5S5DSVzirE1lybR4R9bb
HNgBTbQP7MHbqEDeTcyYziSYCcMNa3G1Dy1QJIxTqktz342aJlt63qeWbawzc1Lz
EMulPDmtc6mWOILfDQmifmhBWMzTbxQpUYnwdng3Z5Xokv+AP0y6REVU2TRv1pOn
uxJgVqSf7KAUxEEM1JJ2c3aqum3m9qcIiZJ31uPhZUAI2b04ZwkTroXLqFuW2Tm3
O3fxpOboqGrr+uGEHeLFjd68cU6x+MXX8V9PZdOKYXs/pYme/Uyn5EM55o7G543x
BKPT9YxMQ5bSDQZfD3/LIQTZfzDSXeRGgDpNAmXRbrD778/7/maHuGEx48ZHrZyy
uDkOPP5wO4wJD5oHpoOLN8G5r8QniErrGtiRTqOBRqSkFcqAL8kUqSto6a8gM2RC
YFc7T7fI32tGIKpu5fGC5I90N7xgOquNdLHEC+f26QGUm1GEWnbBaTDPoBJS2My0
+kUCa/DXIlGcRn9eR6nQRld4zli2WfE+9VowZUdQ+O1a0KfPpvsIOP27JjAuA57L
LtaOYv3NGvZyyJwX2/kHbzD7sVDTqOCP2b8lCL4cVnm4MaMXwHq4EhTu/DT0og/L
JqNdvk3koNdUn9QclROSgNC+fr4m3F6Ho8UbIMrswsz9PIrcYcOQU3GzCqSa+L1l
iToYb91J2F9UUCzfnUidht/zOdyqpbxia8zKdqKaSBFiclEIzfWsUdVv9Zu5syPR
VvA0dbXn3KUhx+IgiZOwX0hjHB4L2L7n/d5b7xS8tGNBENH2s3ZRh3pZHk617P1C
SKB0IUWEIrvBc1YNX5EDx+J5Lh9UvrjMjd0RHCTYqMuRXlowrOvqIT9Tuhy3ECzQ
JzENhbtUBybSxNkfWZpKvpym5JEPmq0dpoYcSyvLELIXWXBpH2tMBPZ4HnSpJxed
XNbO9E4Xiloc3HNgPdJFfvJkBE+UBb1vQrzQ3LBmvDyEawgs+mpNPjnTLYprA8+S
OPRyA3yJNys9S7+3J7J0DYdMq1UbGCnciW+UfEoyE0FjeOuJj6xH+oY8z1Q7418M
sYu5X2oxFzjEc+3UgnlDcHmgU8ZRTKay1Z0Fk/FTJbsUvga8uJ0jqDrP+5oaFsNj
7Nu5smZyDoBm5CD2ZVL7KTkfEeESdLyPJiOGJ6qzKpEG4WXyGQg5/xmuY1VVDPTN
i5YdYdnXfwAFTEEFj5obHu/WHhtgqtJ/gYwtYbVDzFnlrvYOZrDT2xL9MO6+NfK7
L4V7H8DdgyCCur6Inw95PKJIEHa0HEjSYa7YcHAiHCdE16Hdb3yWUvUAEAv9M6KK
sTz7p0VqGt9xbynCxP5UmegDchDaODYYKOuUakbxNUMYzCXg6XAyyxsToX+ZsC7F
XVhYHXFvtlS0y7oaU5Yoad94T/l78tMaLOVrpjUkz43au7q8JTzjP1FUBy7rvaRX
jNf7OThQf0OEBVzm8zhErGBSxPR8+kGVhDhNIGDXqQVgMWLhpSXznDjfPId/wank
Sddi9H9P76ZZtTGRxSlhIMrUMYhGaQgfW/Pd3gJktq/5uHKlyOwa1UYzlfsVOgb+
fZm6uL+FI29v3YwgQQ3z6dCu/nVE4u+jNt9ZVx2jKgN9wDUxYurDCdZQaz1rAhbl
0Av0pexFscM+CLTk5l1Le6qliGJV2BP5NqmDYk0W4/kE7u8HArW/9QlusiCgFHX9
y1Yo5vlXYL7kgFsc5cUGbeV2gDyzC3U93PK9IEFHx9Vk3ag5NvFB3deaBADL7T68
vP5Jj06fC+nfB9l2sSekbUPA6jCZU7PBtt46tE9vLgyseb6uD1PoPdXBqogAnV/M
loIs/9CMF9gW7WL2pF3Wc1FjFrf0/mm8rE2Dqo1B43u0SEqZDPYosdRdkUI/jrp+
JVJ+KQ8+Wle5RqnTyAN65ygAeSEE28PZHi48Rxf2OUDkd3ux4HHl3NSAW2qyBwjY
74769hbb63nO1AmOtB0auK0WOWzld1/K8eiH/+lniINVzcP57USak1c7+YuxnrAg
fBhpGsVCxowAhe0vvNkL14XSo7z7t02vxI6G9Dolkt0nCyhfpRxTFhES9JIvzh9F
kJWZRsN7yYgWf6eSYaqGLEfs7dTcNX8tMu4jzCcbqwpUgJXenvwI4OkG1LrBCuU6
EPwoEFBbfTZcI/z2wDJWOoe0i20Z85SmdC/CxmDNu/YvHGmoK21U4C/JIYRE2LYG
gwaENOGfXMTQ569LqF4VRr13qONKvIr+I+oqqeFzj72TiQbGf8UIaaHz9o/cRCrq
/z36eXTFLNZdU2nFjrTZwL3vxSkycXTPJGLWdzg59luMvREN/FkoBmDiNfCXNZOx
mvVaBC1xtN3upSQRvgGV8WIKxP3a67HzBA36HO5/hXo+TYl/yDWQeIOnq6Q8Hz0w
eh/l1mFebBfKZVWSQBfjvWBtkkg7Bu8upn1lLvtssvHgaNXHfxZH2DOvvX7OuejF
SxjpU9oMIZpD4YsMxC0B7p0ka/LJocRVehMllW9ZE9jOvxhooesmnLvFoQM7FoUy
PD/cVEaHOD4UEbTd8X02vV5CBmy5t58kgUAq/k79KVjNbWxFLBKsfYMwl1gICPGr
3pFdXekSyKQ4HNVlmqv5Pm8TP65KYBIRfiKBGW3wvwMS+HDrjY2y7nDMk1k65RiD
lpDKUzBqtY6wU3x9QLt1ClWKnxrFUNCRtBqvszlsCGkbYT+VunvO9LOn0VWrKymV
qroLyU1jM2WflfZPoSdr5zXAIHENuhtnqYJ5ewTcHkTD+x3TKQhGfs9FQbKnQFDA
ybwozWszCSIv0f7/pSw+Qaqnhf0Qbdy2o3DYAkYT5oXKAAVfnxjDZT+usoU4V2Js
liX19RoGAHeLGO6qF/a6e4Hj66DzuHmVBTMMhO1IjKqOmRUtEfy+6HoB8RvTgXyu
HapCyyUNqgf3BwqRah2r7Z5VN6Hrv4t6bB8pkBiKyRhyJKgalVGGhgi0C+1IdmRB
YY/MVsVpacFPKrT7ny/yLXhnl2vmje9VNYBSWXMnEdmC0P+LIZxPSFyt9+HDDJ/w
LYmkXWDpOr72+bWyvkqP0+vLpa5fDqPcOzQe9lncIvQoeeExKyrHnUfFrO2gW/IF
B1V88WvizKJey+DCPQwv7POF/vjD9qbQ62diK6gpX0qEFF9DtQ4zosZE4wAKWTLY
9f1/Nf5SjsX4DhJ0vYPvTlVyOPFvFdax5sydW8Fgi3VYPRjy34+KVCFfFkHbukJj
TWMRbLqJ/xw9Q3f0vl4qYf0b6bM5jqhbySlt8EPaT/L2D9BlP25qPIhe0KIrrTaw
UyScFHNUsbqky6DZZXvw1WFz/jtlYPLVJDCP63mfhOUASUdfCCWUhE+N7I9sgY5U
okqa9pHQXFIe22ap0qdbxXnt0S9mRQSUUiMqdSLFM900dnwK0ogSVeIcmEMIeQpW
CiplwEGAbP4Sbc/g+p0d4AtAhsKOPP3bEuwoJ+tjOPwxQavmLPggrG+0+y04+oy0
MIsae2ix0aW9W1J2kl7VudgffRf4268s8stv8erVkKbZhbis9Yh0gzlxzvdQ4uye
lg6uar9cIENH8vYt9UZtXt2DmoSea+6PQX43QpGQF43k2eEkvQ2eiswoccp6lX6m
j71TEukzlFsYcjZDrQidoD2ef218C2Lj1sRC0VW6y4jY5kxbsl+2Y1WgBlymH3Hn
4bmpp8PkXq4RvCOS3KzHDPchM1q12d5SLfAGGUhnG50WJPay+v4GjldDjY7EUTnM
lqViMrTstETv7EWqSlVnDlZEMrtwQHhdB16LDoKqFn1iuMeNVVHZPC+2jfkNx5W9
rHHuPhe/6BM4hN8pDAQ8UOmp3NTx83y2SDqEuac0FKMCQgjjkUkdJbnYHhLHstGb
ONEIC/vMNyj+ymglNEFLHQwCtQYo4sxdRnujUh1KeIMsc3KelRWBDPz/5wt50TDc
7EyVeILe0WIxNUgb2718e9yFou+cBGL+IZUZMzRhAgGT+M5ahFEdyFkrDvOsuRWc
KM5Lbi+ZBA/j4kpyQQo8ImGdFCsdc3QdyGm3pY4MWyMnJ/ROYT0jvHdA38GD11xg
ltiyVCR3oh7cVUG3MGrjVxnd+DnUbVACa1Qw79JvpDSl2nRudldOb7rAvc5P0pRL
3ukW8M/yAnpt6lOm9oxHWF/rjlTATbdwrLrsj3FcQ/wmcg9iRXNQHgv15WeOYoop
9fsG94PkHf5pcq/cT7vVv418mFRgK/eQKsdB8MYRA+oq99R31SUiOivB8yhFRQSj
mAM6KeRYadVkZwMTLii7JwORxVrwB5yYOTSYqupr1AxCBgZNKx8N3NJp6Ei8ZPQz
wQfiJfMjo05bFOwGPWAf3yhxoY8x9+nvjyjw3PJ21S5Ctsg5IVA5rl+cR4NXEkc9
NCMDzK3QYk01fvvS0GxyUSStoq3H4vXBpzcEGdAJFG5cTWpSG31JUEebjvBbKg0J
QJ257HykM3kxpDe9CTdCVF58id42eQI0REOkeGyFp1MUbGvvQXy5VNL19NlSBxKZ
SLIIz1gFj9xb0JS3+IyQUgtEBju0HEh2NhnoOlFuBxZkwK2u4V3PNxPPaLWt6F6S
zqP8KbxmPmRGDr/b6llvuARyfdw0VOO6iyNNuzTZP5DrL8VOHXFyk9bmehTQW5tl
RVnrJn8bBcOW0TEm1bjq75qmgGzFw+atMF+ErtiXbOEMOeUWeNgasjXDjSpoBeAa
4fnPAGPBeS/0vg0HoiP8T2JT9ZuhQyxnlAJ8yHm8ejEOp9O8wehTWsd5fviwQxaz
PhpJN7WksZmS2mafB5qNcb2JDGcaprG1C3DDC+r8D6qrcAcuRenR6gT8T/mKTs1L
CN/6zdOqc/YuyjUTLlhGpn+OglvWp0vWiSi0gcgiUMju4CTQUygLrj52rqP88vfA
tn+U4bgo7kSmekYIaLwjG1Tkd/3QaZr0FUaUi1lAcbBLuK3+F3dGTrzjQHDoSGGc
cxAmXiq1g3Y3ILI+8ZXz86Tfr8Er8ST/d+ID3deXz23zq2M9jBPV7vE1VR84jH4A
PSd+RS3kaZ/ytMo95tt1krxz1K2BbHE4YCVI/P8O4l6xaw/pfKBbdNovSV0STjh5
gBchrQ/B5apbVE7C60obIL/Pts8JZtksyeVkOGSlLTmNVddAiIup5uG4ZGxGIzcV
F2G3O+Zee+TpgMQVQafht/x3sTfXiALe517fX5tCO35LCugICNW0ej75iJ04FS0p
ph/bmBOHWlgZMQdZHMFVKO0XMFSYiM5l18W/dV1XEoOXBD1WPRs/tdWkzbaOhur8
jwzsoxmGdYKf7BG+Glf8hjOpfMW35yarFd1piCrmaC2HmCZQFmlbtbH9IlS/4viU
nJ1Ar2JxdKh4yYoNjc/s5mIf/NvMW+TXpWO/nKfzdCmrdzBtNjkGn1XUINW4If4+
+1V6iCOWF7dYleIm4LFY2eDnd4g9qSr6zBMDFhp/pESNEhAXNsbtBz2TcoHb8iKn
fpErTSpDU82jELmHhbmyHa4wh9feRcj96bXxJk2wXILCcFV8OIXn7NZsYfybSPdV
382yDb90sadbJCeQKs2BODjB6Bo8CVoTytiNhi/clIXixAYZ+8//cPbPnl6tBpaf
POpJU6pzq9z3HoNmfOQ5FzPxqwZLr66Ni1iD35KZN1BfdnsnMDhc61bxwQJhC7DO
76/yCf9x2QE2YJFpzy1Xe5/5fTydtRix1F+khYMetNTl4E+0U9AA+1x+PiK28NFA
qIejR9IyWRcr6wjp6To2TjMMDAlg3SvTivDFj2gKiRugdNes4H9bRIbQKKiLYdTO
ygpgqMVdaxuUkHtotDrMqtHyFc0dadTP/BEXIaAAoYUbzE5X4fCTfI4YGkpJJdGz
PqXgtyhdUr5+XPFi3s/3/VFuHtShj3iu96dgXl3rQlOZktCU8ZhGwYv1/GoS+rMw
Oaw+AGWr85KFOXds72CV+vvMnHYghDjDmUJSohdDggZFrLfkeqYvkSeV0YrxFCle
WG0W4r8RW8Xn2WQW1iTj6sLUQVoRLG/OVzWj7VBh14OP3rQeysoSEOAnk3M48Z4I
06H7+vnR/dDkBtsoxaDkY0xxEvhcBQtbdaqZDRDtIC5AkBoFyAe5st7aHIdSl2aJ
P4uZf3tZpt3aT6ZNZ22vbN/weqvAhQlx/WNJbOd/su+AhGJD158EAf0q2c0m99wg
3d5tL0H+CVBHWiDd8F8q61l93luBT7ZQzDarUj9xBl6cyRPEzNEYXQEsv87B7JI8
KNwbWL5grdN+IwBtSPC9LabXPZGOEKH6Q4sdUnxL/HnYtY8Hd0Q5E8CT/LPE6BuJ
VIHdi5m9isI9l9n8pwUG8exzYXVDPjnwqIsdD8sL3RvVspHpPSB8XKPPYmYIFcqf
DEABEIj72RQ6hBBogtS6bq85QQUuWE6d9dTlFSFGJruSxOjA3xMeJa1sidCnofkr
Djsk+9K8hj8MNuNcmBGL5tZwrXf3/NfQtlSuUSifUY2zEnxVn3dwgZRI8FGGzIHW
h/Wxvur0UkrZki4eBaLWTgtZy0Kdv5tQ95vcX2hZ2ahYP/VbHRvUJDJL9wGJmJis
+eBx1xM713BQ4x4h/3BFi/pPgWkzdN7q9MdOokKhQ+60OjZ8swzTFaR6uc+rBYhp
o+VwaVOCBtMJ3va3C5d5Lsn8BfJVx4cZyqBrHKXLPlT0eoBrlxHCZnBxWz44z0ey
NSoqXupcocuURO1KB7VFsXQotSguQSlCK8iodkEKTc21JiM+2taVNM3XAJ3oEAKQ
tMkpyO1gHNoBRZDyHIeezz3KxcE1LTVLGvzeMT4GTMs2Hau/vn1aRKEfbB5E/TCk
31HM9IikAeEyNIzxzZOjnHPc0IepFWd2IrYGrmtHRWoL8dhvoxqy+zXc3pafhfz2
gIhXA5lxtgRuhKVRWfyUwsKHbfKhwoX4xC7KmFeqcnDlsg7AEWTfB3VNDpYw8p5Z
mCZYypCGmvjdUaIDyIYuRKNeat7Z1fY2N5C58Hqu9KxWlN8TD+3l+ZVYEb2/hYyz
pEaikxT0ftPFji13WTvCK8SSao9PdWBogNCniKalH2vXLb6gSqTnZtQ476exfPCF
sn7/To9MjbKlUAVgdfJz1INmZBcjL7jLTCft38O3XUU8Gls2sUHEVWzWx6LB3zVk
Koho+JWE45ASp4tEkwVUVCTX1lsS+qF37wZSzoWNJ9jbUVK0QzWEU0kLqVAzrYcI
9fVCSl5IAFMI9reP3tBuy6ymafitUAoUzpapHu0drH8gNYm9HNnDuXLUgzNTN68n
MYf7yCEIjO1ABBJ4yZXJu1+rRn3EOSvOaj6TM54fgDY45tMVrTrS6kk+ilGRKNkF
6At6n2JfAJHnB2JHr8nAUnP8QtuCiZImyAM0wetR+D6LEPJUCAvi/ABiCYFZ75lH
ghw2UVjjz+rgTAqLL3jaHzEzScLz/EGRvEKjN4iwiDaWbScUzUCJAfZTGu1q6kYb
Ai4xLp6ZNKUT8gRvcvyQp9XOU5NAwoHMahOYbRVfSb+tYPoiWYIGb4Z58KiP7kXx
h9FfU7P76fU1WxQqjdWA4QR8AaJ/xvhFpF5FSIw001QU+y5Snh0J+56bcmfXxE7J
3DPb4JziBMOvqh2j/LjifriFuXtXk4ZjzO67dx9FW6cLtBMUGpRe+1/KgcyaodV6
wIl6PFRlTYp6dxAsOxjMp9HDuZyC0HN8vbj7WNGzbIYJ0MfB2Zle8pjbbnhWSUXr
2iT+z2yBpeE26ZdSfsSN/jOC4/RkhpauIUGkU9K9XDNeKmVZCTIQWulfnyav0Igd
qiV4mStjnHKNofQdXdlY7PEEoC2tdVw3OBI6lZ9q3RXI+WTmiWAm3+82V8C7jA8K
TMb3v5IoKHTjst+GnTvfUVPs9iZJffcIC8tNm2fBUX5FaT+OJgzRrJBew08r6PcF
kmqzCNCNNDrjmGi7fdcEXWDrsFOup6r1lWvw1bPjL1FqWT/oFebLSfvfKvLFMoI4
BYWFXDgjoqmmn5MWj5nMNFsRjDlK3AetSh3CqiVha+32q+kocyJsm8zeEq+KlYi7
2xMGVK1/EdPGyDUhtkO4OjWp5mCENR0zLCvLyt39u+4BAgXTWVlVR2fz5rM2IyE3
XBu3i3ZwsRE8Td8cBP2BBv2gbOzs/7QyX1rrBBMESMpCpGvpYrhhDixfR94LMcZL
WJWFfMxEqlDRph6geJ3Aac8SkadaeAxYuJdfA6mfkY5e5stecoU9i6nnklJXAckV
WmcPNC/Y9ZO+QXiJyj2jhAERpzv4f5DNZ2R9qwinsF3XpQotc/hWwzrC7bPLPkWv
z0LN1ZvAMlbG7prQGO92chUFGDRJhWfO38/M4pEOi84rCaU6UFqslEz7GewKu3uC
JwWid+vpqAZYs9kz5cjXV1nm2J9JeMY6SJrpk/T0GTrk5KykTNd1fzz2lxS/9CmC
64JaLf+OH8+r59jS50EGRl5g551ntqZy7wPBtxTofttBHeahotOapvZ29bbNAHH9
wwbETLTHpdbvTMc9M38OGL5G4Wya9wUSdgakzi1qIBQVJCst1lo79XzT+jDPv2bJ
vpEIVzWtr+OGUzpHnSuH8REHvDDiAmZy8Q9FOBy8JTp/SQG18slqm1O0fci38SOO
b/fplbkyqcbfb5RqVwIqRQ/Hmr5Nmqtss1zII3Be0ykpouCx9cbpOjCuKpjCHwpr
oztA+Wh9v5eUqP85TpxbvTaGPJgAh/Q5U4RQ9o8J9d+snO7aAIKKfhovj3g7csZO
e5DhN6o4l28eapa7XO+Nepos8OUMTXo2GgBbqVtDqpo7rgyPyGfo6LvKmgM3tUkS
nkuRusrZFE7L7cXnKtnCuA8LyODKfOrthTJd0wfs4ayaprO5fDB+p6AYndmJiac6
AIbwNiBZjIMTi+ohvxjqk2sMi70cy02Be+Xrmuor72oqiXUBLnhXM9imZPkyZbjX
4+CKjtYgojOySBFZXkv7I9Ro9s9dwDBxQk6DF3lJgJ00cOsqHmAFDMjfk9p6ZL0D
EYuf76DG6Eo3XZGlO3fwyqw5TlS3nzYEnTRsfk7rMLSw18GtDzRQGUKmuwGXuFXQ
OkwxPlz9FbfCAB3chHswV8/BSNHG1TtQffurpb1o1HEA1JSwmSPsnBZifO9sQbrD
IcJXw6mim1xIfOFskz5lM+O3tR5KXjPlvC/G4Eg2oZUB1bY25Mhj5CaaTsu5Oaub
xe1V/wVT3vjYV94Jgf0Mfvo+YsyY5SE2ZaPVHonCFYPhenCwQW3Zu1xBRvC5c1o5
Qr9hdugrI77OP1w6APVeftDgL6Vo/lXPlAYbGhQ8Krp6iKm+7F4ZoJ+sMkHVSK3H
B1mmy/q2EKSVY3MLNMox8Skh8iwt3EdukimyPwkudEWFOleLp+vST05gGzUk0BF+
YkspUiMISrNOVJxRz5z8wSpWH1R1hjf8tdOab1xlw7vCGlRViM5rZid1xA/ZHL5U
sNZ0CGEdSkFKywAjIG4lSUxj0rk+gQtaVXLctqtb9paPjnKg7ReGfMSV/RYWNnbz
PP1I/oQYwSwLZPF5vIMWwKvsW6n8egiEqIgxiVNV3sbWzxC3cmn9UzzCUiRJfCa0
IO1nwNyQ7TiLvcM+JwJP9w7CLSWFD7r9QZSMxvkLfftzPmev3O68j8FV59L13i8r
M3riwYlPZduG/R8jhvTdQUFfb5qJG6l5CczSEqEXj1pnEUAkDkqCuvycZU7eIi0B
tbQMK6CMgZXoUgoU6DNqd1OOEKFLG2rqtX0cuAxL+hPL3e4nG0FYC5MWWLO6o2px
HmUQFcchhn1BY9gtXBRGc7Po6RZhChxEiNHU78APW4VBT4FVztiQGiYNvpOKIUht
qHAixUXl6+TBLqen5PhVDB9By90Spmuet1Mjz4HSPqnTY/duTJG9cXBx+qJK1Dvc
SiZbq7WGf5eXAxoJjDZ3mb9JUjQjtqLJNb5pqOfdJFDK4zJ0TNt+llU+2qtzzW0x
jSqGOVQHcSi4bB2SjOjE9dgrc5nUHSVykSoNgRo6u3INu09Z5veoXH8P9lfXoWum
4s82CbzTHpxNaPCh1HBaJTeF/jTdZSU+5wLZ4FpU0OQY1DpuJsG4WxrQgabtwnKa
7/yRIf/Wj0KOdM13ps01R1vmHp0s0iUBYxHSYxCxlNkoUzXCJVXTE+d5uH/vnglK
Ra1VJSPxNIWjpiNQQRLSbExeuBydqaTchTfkqGxk4DrP8Ggj2ymfqNT3X7Sg+8+f
lLp5NNm+WNQ9cZFTEGXwNOIgJUAk5CCX9cb5TnXM6CNGqkFZN8leZOx/aEo42i9S
wCAjdhEaX3s82fylr/62YO2vg8Sq+P5tGNcjr2gvC+4ddjJypI17sLWggFCqYb2I
wpJ63ZOh22L5IKepKbeSgaZ+rDJNqxt/Vn8ohcauzo01MYbdKsvXaSWje9aZeur4
irHoRuV+/2HqCTksc00b/EtPKBAdAm/JoSbEvCexXSMs0oKbhBM5djbUSmsHo/ra
pAGnOQqxQ6iIA9dn9bg5KtMs5IO7D6MPGENWIkSE8zEdZhH0T8VL8NMAZ2uxobIv
8n07IqcUBc0+uzfYnH24D++ic7pOyEp+N0NVchxwRxG08CFVLG1bp2/GhlezchN0
cLRnEmmvvh1SFwik73hhQJegzzxj65K7IrfqkqdFAaQwU3lsqqLbbqItUW9qLMP7
FDY19f4gMW/w8WUcJdnPq5mHwqngWTWFDykaIUeBAA64AryI/2NvHDRC6xMMwc4o
Q4RSEObYyA8KMO4T8yNySKzm3q/aq3k6hPaKNFsD2duqiFrsIapK7lV77tgyOzNP
H3JD4quITQf6j9sDs2towiXJ0RSggqD/JSjLACf1p6nk3vH1PwdmN8/rutvo6WJX
TWf/DYkMUMnDS7tLRCgIqcjAf6hxzogsm943Hj1Yw0KyrfPl07cSB0SWqV7L6LYw
AofFxpgTg3iCi/V/dv1XNSgeqjspEb3sC1IKTK7KvHi/bdo52c2nAzR0A41sWuyn
bE+yRzk47ipaPbb4f/ScQtWyAxwMj4oBC9oRFEzXvdgE9B4y9c3o7WR46K33SFt/
+6PcXEqHn0KdCYzQ/EvC+ngTZeydBgnzTPSttQ4+Bz/hZ4S8WlAvFNnAVwLDfpOE
bCyV2OD2ad/YzlGuUHtTU/50WfiGvml4X4J53ZWF6NK3W/q+WA2jVj6uhsxTg1O9
KHgQq1X8pDRsvbnBHJ1ORG2+xHSVe3pfs5XzXTe6m6x+b4qi7BRtEXZTYXQUGbrw
VSuiNZczIT/eJMVGf4cgp54hQ2uVcYbodRSpyumD7hXS5RciDaZY9lrd4PtGmxvR
pxk4lxBpzelYp43FwzfKJ72d1b49DPlGm0UPyd5w/YAmSDpFYKuC4vhmip/TP5Zq
auEW8UoEuPoL4VTY1L7nzf2ASG3PtRSNFeSSzIWfZV3VBG3Svabd+NmVPY6OzC9+
DhJgV6bdUj78YHW4JDlxDGIRpPnOUPSto/e1FUN5HQmsq1FwgS2ak+enMs7ab8y1
V26xIwQzAN6uC4v9iJkNXsY+m0ruHql+dgvx2eWxaXtGQoVoA9LUa5cYE+7PPvC+
MzCaHHyqe6RaMjbaO4IZYmDx90GLa60d+cndFwrk8negr7YQ8riDYv1etRB/f4lK
zp+Mrf8+tNKmmUs20NW2d2lmribQrU04yuADtFs9jDhnazAZtbAl9+aXX2LQ0TTq
sPzsLquE4PskvP2qYHmX6WYkI9c/+NvlmO0Vu2vyA3tfD5EqqY4KHxdUeEn5k7Kz
w4hUDNe2hxqGCVij9LzK9A4QhIkOLokqu7bMl484MvVOoyeukjaZ2N1bouJyV+VY
tTv3VSO4ru1HcR2jupJtO72v0sAFZw5Moh7vOf1f4XnIcM2R0WPnulku2SL6ctp/
qNRd5KYJN2G2I4F8h/uhOoL3IVxDQ6S1c3QGJIu83ZSA667SMrUJcsRZqecq1RVo
lLRSPlNS3I4ZExxw8TswEyVpyHRdbdWdpYVP8ykBadvB80hNon8TViq7FYjLsKtR
MCliz+dU01uBkMECaqGBHLboT2fJYNxgGmIufpliYNDZrUnlmrjAQIeszoF6AFvu
R7qnYVO8LVp+bLBPYSYu20l0Mk2+G2BvchtPrcRx53LKvAvz6LPRPfE3BCYrbdjp
Q+p/Fimp74f2WNbMJwMB/z8PMteSGRebjEcQkRL5JX8HG/WN2Mkv5ePFii9+VRL6
JXlbYbZND4cEUvqOSTi3PhGYJIWY1PkVygQBbVZXSU5pSIKkMcTMsLxGY/H4Kvv4
nVRFsYoG9AmTFKFc1UW46HM1EhVZz+6+L1irb1QK7iWONYotyfBzXFDxjHdIc+Lw
oB95bjKWTtpGvk15K/tFL+rDjd42OY2HAU/n0HCceedgWeEsrkdAS9ho71t/B8IH
fq+/n0ANOsYHb3uEX9Nmb5tX0SGuX8vzqx/8QNZOgNglzE/1r/Fth4iVvyYPmas0
KPUrcxsy8POtPCVeFaCsbJk6qryYJpbPKaoLqYLiRK0pexOKAP8q826krrTSJfjx
LaZolb/xEbR/lntp5ntFI+L8SFjkloIvpyliSU6sI1ywxq9kGMJryN3JsKU09lQw
pOhSLYhk1Ovk0rEKBVtnmAYY0h7yt+ZHuy1hHE7HgYCL92G1X/sdkNqjE3dWNvu1
mUXa77t3fOr/xkyPub6ghybJVGtl8mSlc1GpZJzTaw2H3J1G3R9kPFElWL+PnOOJ
GVhnJ55zKjfunjDN3TK6UjFLaSZ91Jw2mMmwZVyMHc1564TAOCodNEl+Tq9bdTvI
LhgGyvezANvnnZ4pRBCY5l2Pb/nkp0cCofbao7ugLs1164aeB+UEbdYnTMKKULqB
0jCP3KgMDjmoHWiU1tHMhG1NOEK3RjnojIUMV+1KYE+cUlNh3xQXP5x5ZGvS3u1R
y43jl0r5ezuxXL9i4bcoInmdIT5GNgIAMCszKl+yXDvqVMilav4BA/0Dc9S3K0gN
3PNXWDdXm1jGGLe6iXAuvDybHaXDceLjp2ZPqgwOiaxldAmPUGJ6aDMrgxs8QWKw
Ve8HOTihIHupS2rHFbBYDhtGQ/ufpjj+CI0/mGNOUWSiuiVvF01+qXjNjGLpl6wd
a6FcM6smRVr2Ud7/G/JhrRykxzaUd3Xbfdm053Xq3P4Dgom463cgslYy/R9xeY03
+ec+hJSkWiI75/WNVvxDIrPPah6Kt5Q8LUq4ehseo8MPrWqkAWp/0z3SP1Mb8fZ7
ihLMik5GZUK8gSA3E7mZqMnPrEQbEG2PHOD8Shp1tSRYPAjKU8t59ZFMgLpeGrI9
ULHiZ/ymSrZmZ+jJ37iTZNeAel7Y8C344ofb1/np7YcSBD8KxvxAyEVW21fDv9hY
ipzW0JpYPz6b+b0lDT+DvltFmcCtRb0CrPeDbepj00F4pvifnGeIUDnByRTfkftf
v14x4wQFuMGhBP3LDXuD2b/TBuM3mQicjUPq+hgDV8ng7cai+ZXI8tZdUnDVz72i
IXs/shfhHSzQnDMrVwlHHEK+UZ3r7MqxEfflMsRAh1HEhKX9C9S2GTNJUxbA7050
D1uRlS5lkhGiodGq8Il0CUg+QIuwYEuDdvLxNxwo7cFxMsXQt0qIDKN/R+iQfI7U
GfiiLB1DaSESRyMmdIPtc7fz5dYledOpBOv2uIIgUauKmsPCM/VsR07DQGIR6mmP
0BwaW2bO6XXNFz+7c29ocGcM4Jay546m2E1q9IivqsU1x+uFSQJUGJn64C3D17Zv
SLxDERmNWHykPxVBlybhBuuDpd406463RZfmVGuPkj4wXzJ7Eve5FmiOlklM45/8
mRl1+gOSiwcXXMun6a53LstbyaxQuFo39HScyOb51nmSyif/eHrSmyNzJ3SsJ5AS
YHEB0icE+uaJFTMR1wUsOXXhuKUNZpnuVF+0GP7F6L90G42gxxGx2QWEnRMqrSa7
q2Nl3WyIFNcyCKF7ML6L0i8RwLU69MBbxKEqEDl9efL7/oJhppyPwKF11MU0fJCs
QGR3U5S/+PO2pAaPT5NwmZ7zK3Bq2IbsWll1yvMn9u3WbMNDiXLsqUYLI8uKQpBE
kXJl55COVsmIMZbAK50dd0bh9qZIDvMmeSZISmuB9zawoIJdVNXnuY9JwwIWHpvg
Z4sLXqY6LKCNwk/F31JR4eLnHh6xAJKeTV3afehlYceL5jzGVeBiv1Ipv+qLRvHF
UxiXwW3Edloa/K1Gv8C9ch2eE+Y4G07bIZw6jO9c14R06x6vsZCamHri3RJ8O2Ci
QJFP1ugKwrWWhJ+DMhkrwxwXwkP4iMem4IY3AVziC9tf8ZrG75skd82yWWkuShoL
ktIYmalFLC0spyKJxd+ZGDt4Sfj7tAhWoM28q/dacQhaK5TwtqAKfPp9t0SMjPWX
IholKgfphmXu71pj/AGWqV73fzMFhKo9/RqRyvS+vjwvC1zWH5ExQVYDWYPBHhLS
XBf1/qjycxXTv6L6BUkJHZxuqF8hOSySmpNHUnrDQiQfE/nS0VyAEPNHLIp7fgTh
OMCYMMPTx+YCKAxPeYETTZQAlBS97HQ1s+XY3Rj3r/Q7bRBjSmsU0EQVAepblsr2
6o7OpYa5c+lNJtmo6KmjmTBghIvwUWEIcrjZZhc9MU+Zl1fp6922Yswwpmo+v/2X
o4jRBIk9W9C+SBy5gnZBNmanT5f8BPPMXc+TEJbtY/oFXTOwSxgFYtLattoO9tSu
J0EDyDRjLl4MZYJh4rhPK5+dB1ROj10o3E6YpMbkm1kWHfXNVrKN1gygUOuXSJ80
YmlTnX07w3+JHKNlt97Sl3IS1UwiKX5QHnS4ScrVvRt2eyIy0xSeOXVWkgy/aNoP
4/rDzjZB6syeCItjdXjJhHYK/n+gJieDwWtyImp3bNmy5JB6mzwSc+aLOC8WcysM
gyfnGvc9Izy1MN55YBp/DkwwPAiFicJmUkVYAFbAhPx3uFdTVm82TN1IzvkSMbK0
YP9k4oHpVjAtZV6BphmuNHttW6iaBXYWLGsKXuuJTSMxGmxH/ZGHtbqPVl6hl9Yt
DhwwjTzJXGhDBQ7zlbIj13m9zXR0yC/3Bz04gkz8Wyf9J+dJdV0tok+SSBhhD8x9
aKDAJNHvucG2DbzxPmqt5FxME2NSDku+4dUBRAPZ4mEMA1+dcD5v9YPYCsmak+8s
dEI6iCTzrVJYAnvu3kk0nEMmXi1pNSDq+76v0S8100MbTSJ1zjZG12/hnAFrxBfI
aXuN1hyX1fd5/jnzm3IBnYXfRO4OFvC381NKCWU+3mzjPFwyxpSdTUGuoR1LZSHD
zeZAiVuzYgruNJAyrxyyMwQkLUpYGNTT28K6Eg7hXzX8rg9++j1DqGp22ddGTR1X
0GRvL+p70r8HOzofbpX5Ay27i8Xd0cRghmdYuvq/7XRBBS3R4ApQyJ4pfyC/XX9O
Flync/oqcaAEwJLYLHtiLixMPqWgXgfjMSdJdGbpT9i2uXxN3uWvrXZzQ+i3B1JH
J/lS/cTaNEg61JL+0l20aRIXJjmJIF6nE6xXqTzpZRDXZTV2O9N0Jg5cBwMp0PBU
9enyPIWyYWYsiA68Y3oPJWScnsc2HAFHMnfgfA3TeFGdz0A6m1H2/SZpGTG6u8fi
YlOyv3cqvFL9VQJL3iosb6Vk1J/wcMYqJqxGfc73h8PyAqGVAVo0Y4eEZ675CL9d
kDHm1vXS9WzC1K1z322qNf0LEVddZeFX2yol48E42VIvX0hLAFPx5zkZnWx2Go3G
3pDGFnbTUKyVBKN+FOFWF9a0S/oIxTL1lDQrBe7Bi2w4Q/e7Hrs3/9y8w6gXXYsJ
oa5MO+lpP4en3+SXIx0WZhKfvU6x4Z4aX8utLyY01W84w8VM/EpELEQ/F5Otxpy+
DjpcNdzouGXMXL5GLdzB1ooZnJuDh2LWdYjD6S3Y2qrTIMCvMWaYGRXlj/45erIX
RvlzR2CrDBbXDEeztef6GZaCCEoo8NKqhp6peQlPtMQFsZ6a1dYGKjGPvAxaNxna
SdCY5RnrY9Erh79C9GyZfJ3eDOoMi0V6tv64a3QW9K1EhtJ9lHvBicgUZ8fg+eaH
nBY3RodgTUa2fEVafLORJN77YWi3cHY+W8E6mGoXbkS2kItbJUSe8V5DkebFiPj9
ZrdrSVnHnveS7dcx/ZL9VBfuRPJql7xet/6oWRW6lnEQ+OkfF6QkVZ2WwZLCwEVN
abVBcPpNlctFpexX8p4vzk6vMhQPn4ufbS8LJx0ibZoEgYZzzupdjqWKoxDkrdiq
isbpp+q88gK8C8VNnSjFxYxXxDYowXtc6YQIyH0nnIFNgvgPLJ0Gk4Mh8AOGwcPT
cutZlHGQbqGLJXOtIglNh4yYI/vhb2s3cQ1gyuT0PQZL4boEz3j8c1sJfZfQRxVs
lTLPZoEsfk/ArD3YMFF6XKkutiNjYotkKlLQ6DeIsU4oOYidbFE8/n0h7j+INTED
dOjxy+JLifPyZHqCxwuROCtVNhL6rAlkg2LjKh95OxbDo91RAVxNdF6FJrgOx4iA
ouL8oHQthedSlCynFSBBvQSq/bpJxAOLCyZ+YotG1qbY/++N+ZNSaBp5kW0MkKRU
gKn+wzGcnEdzvQYCis3eNJfBnkHLpRkh7MWpfInN8M1GKyzfqmOP6HtcBR5ddlk4
niK0GNdLVcfFKgczeDGoPm3sIqrZXf7PWtJ3GB2Tm/8KQou7QXiWpGlMwSAMgi2b
zB6dcsDMMQzdM/2YDOJeBe4AhZ4S06e9p3zPY75ft8J7yeDhSAPvoTzc22u8nuOZ
SlH44rNu8Y4o0y988l/gsyD11AIJaIIPRpxQ1n2RmLmbARNmboL7r4Rwx46elgbY
7tqbXmWoSToJ8Oq74GE/qIkGDzMVqANTIKyB+HQ3ZbU3nf9NBPSESDsBi9aIpvK3
rvKaLB/hRcKmmfIMBVEuMBqq2bxoF7w5h2zNpbm+juHZmTCGwxsDcFXk13g4B5v+
R6iqY54LbCZFkpJt7EXNGd5kjqGp/3N/Q4jaurS0Fty9jQJKLDD6wttoJCw4etGx
hUs4f1Dq3Iy6u4WjFpLOvP1NP2RgGve3grNbznb8/TH9R1VuoxHMkp8aZ33phKXp
K1+8mP5m9H95UV/9oVUJM9RB0zVZ8gdfhW2LGbsJf1V5m0JlqjXd9B8VUjAZ0xs8
39CzuZUt55J/2zapWPKH3/4vV7z59jWQyDB+eSQwx07rkev7FN9qAo0hmMsaOqKQ
NtrmkwoSTU5NFxPVPdF/zknMTKzvIK9oCponeRTWb9L8LGqqoHOJD+MqzaZghP/S
ty8TS4yk8kWd2YlwzhiaQFgGoqBoUJZlGI7qwNbtphnV7vgkeRfi/R/BeAapX/SQ
Q28k+u/USlcEk8ajzrsiedBlQff+Sfg5ES4rEPmb8fFla9Qeq1FuXMH6ODPA3mXf
ou4ZfjAS2TCmBg/FDBv2cL6hT8MpkbxyhzUQzRfSlR3xHyQi243CESQoBQx908Nj
vWynV13j2mv9g6fNGZFH75zvN3SU2xvPVnDErmQbcO/BNIVlD509mAmcJ7qY2vBx
SNVMP4f/1laT5PzaNy2DAOoG/7i/m+Ko78N2jQ0gO9V7ViJJiK3C2umlzC4IIeDX
HiiFTMVFOTgWD8sxxczG9O16IEwpDrMMV5jYSAP2DOiUpNFx5IYpPSk0LH2PXCK5
Y1ILa9+Rb30vMjBU+6USt4Wjwg9hgVGLU8ufYrMJzh/7eiT0loNIvOqFQDSwuL6T
5t0x/sA2XBNrA1u0d4ie3jSgfyUy+iu1qEM7iMXaycK2OJlAHC4Q6nA3T3rk+PP8
iqxFe/deNTJc6m53gUsJSlUn6HZ2ITuBd2E9xl7owWjHcj8+tNp14WLf2/XyU3Ij
MmyuIP2Phqj8BpqQE+MyexGMD54Yp9Ezq+itOLwRq5ZB+xfS2Ul9PR4VTP4vb1mg
MLUOP4jNz5n/FSX+RVVj7CWnCga1z1rjvn+o7U4TJEvIhF9Sq1USOZTLcDgskm8u
1nI2L363czs4sKS4MSo1vM/sM1XvhmISkm0QqAhYM3AcxIbuXDfjcv4yefQ3QJns
cHD4hhpxrnscpoayr3jhhVZiWkgtV5hosEgLzM2XAAxn5N9yYtbvlu8VkN5Yf9Jx
hCLyw0JiX4rbcVi7PSVJW3DYS2W9gdtqqMUfwcyP5NF5/n+lwRHrSEV6GPj4Lvf2
nbaNpj08P8+QAMUOzIVoD4fGSZZuoRheHz/fyH7XmUnZjUM//66Pee2d7NhNqH5y
dXXvblVU0B91w13LZT2QB5yXiR0D2JJzFscL+bm4MpfKT3gRlN/sRxdZkH67gfV5
P2U5eL3GMBem5F4RGdx5xXc4Ds24voyNZVc/aWo7oa+XdwxuGQwjw+7KR/SSx3bk
Dt4Q9OX3m4UY/IZKQKKhGLiXn0ptaOFUV0AtButHskeOWQDYLiLT5NAk4ugyEEXq
k9zr+ljDiSoJFAlen7hif56KqADlAUuHHxiTVSVjSk4AhFZ4Isd6eW7CgS7+HqTO
1D6fNKueGoiZB59vpmTF2hPm1uRXeOL/Pzc9nlfgaOP6ASnzO4bIDW2meHYCQHPq
GAn8uxNNm/BlTeg5yXOfHkbag7kced8ME/fEFhBAVwf4Hv+4ixY8DtHZBRv602qL
JEFUDTB+caFRZHczwmJ66xoHGQx+1Q3D8KLUVPXrF5mM/EOceWwphRclk6hiAyi1
LK95mFSEylohdt00Za/PI9SAT7EF+iDWi9QGjc3nM4cHWXP54zW3yHz0pqp5+mOf
GrzwC0E3WBHlG8859wS+dNbJ8DLJshKJiyVMXTQ+JjOX9PLXsykxYoPuXH/n+M4e
dVv3hb077Dvi9nKNJQjLEDFeyOLA6/YinwGHrLpAQ8xVplYypingPxKm9Y8ncJOH
l3rF4ssUh/KSD1C72oucRROu/v9FTHgFepBAXGswoHoYQTlNFZrI5/mwlGtyQpjx
nqoLoNIEv89ufWDLEEe52nFhcHBA3X0VaR1782Ebub112tU6trUKnog233FmySkM
zkHajeUPaJ19WFi2yIdFQU28HFshM1Qvm76jLyzjJeDQeI2SF50rizWUMtBT09Ua
xSqvFzlxN3RNN1NX62hfFHgzaFeIMEC/+9YQFF283M3GUf1yoTRk4OScCjFCtHbV
SZpHRMnPuu/UPUPVWoBdz1l483GTdhbYFNYGUHzosO0EODxHDzRh6agN3wbGjxs8
JTjGOIrnzhqljRPXM5UJNfwMv5dw/84hJLbjecpNjYUYOqX357G94hAr7JaLUjHR
VYagYmAyqc/9ciuocnstmm5fehQao1OXeQxeRuRDadlW2eP4NTe/q/XIp8gtEios
CiahLFWsjgnl0kxrtjSlbzZR5VemFWe3aTAyLAMV5UnUWgSuoFTIaQFEtyMuhbk9
ntIRhap0vqymR68PNu1/SeMxSW350ZHDDiH2muHv4bXjghRLDCaZLJ1nliLjn1mp
7kvatQymuvJ41ttgwWn5CX44IhjXdM6C6pYkyQqGEpGJ014pVyagPNHgm7AzcbWQ
3zjBwsdCK9wEh9HVRSjcr2M38KEFAIjpQ29vTd+7PJ7dw24YN9PDbkb3aoSLkKR3
3gVMIjVJmgc4oDWUjEH0YI1BJjJDU2sWZrCkVkaT0nh10uYnPmLs85MvIkZLZiDz
NDegC7dWJGfQwg9Mhz8T45f9q9GXWqUXMtvY7c6kEVWp/1n1r94C6AVlORS5hr8N
pSN3kj7XMUZZQOGdLOb27YYCzKr37EcAInr5vdWi35NvTx42BSnFafUvX1nZzzLQ
+OI5ijYS+aSsTlVzQkcqeLrsbBhGWNHBZDHNCSt/yYCy3nra7IHbJQg650mSYqyu
D//+btToQ5FXI/5T2gorHkv2INe9+TZjLkbrnoDWHt8odm+8oiu+hM3YXW5IZzRt
ACf3gcE5sehKVOFWsU6Q5IVzPFWe1ajnm/S1BiryahF7Y+fCuKAiA/cj1TPl7GNz
Vhw15rSIEKU5UFm9yLGa1Py/ZdhioF/Gr5M18lCFfFNh0BslecpljpsejdVM/yt1
IIqSXNEd0JKR2tgCqmPpHCt9qDhTavVU34sxH6vXTYHjWHabD/ghZkIQMeTvBP6Q
oE38Ju9PwOBZDwwJcfr5Mawm7EbDy8trLAnxXA+gDbBlWn/45eXmRmKHGRss/0yn
SU+fip+1gTegsaZUHallVZYOHEl5tM+dEbzaCfB6CZfKtyNXYREetP0uBJbyUGGa
xmwydhgwdtFEFj5R8Y8dMVLAtG3pU5jS5ax9nIU4vE8/w/iCXpongWW0w8Aarpn1
iOTq3MAaVD660k2OALWLh0H5txbDQPMJHQD+zShB7ziHO1uT/s1ASSs6N9JWfNpf
IL4mvm7s7AN6JVuerwWNeSeublJeafjYD2tHcKfdmc2DsUgRmylTo49v0UDeAZuP
14yhUX4mKftkNwnHoUFflCb7Sbd3x2Pmcj8m/rbfncQLNk7JQxv8e9H4uOHLTfmH
kqi3/vsQQfBr8oD+YJsirkNyG4q1lIzDhqMxrZrqvAcbOhmrYUL9jNGTvydboDGG
P4G8NoNdloTPjwkk/dyh1j3GdnW7cRue074vTv6dnWrYnnkK2duKSrwEax7InV36
YcRJujtBptnEFgxY3xpGuzZnkf72KcOEAdYUIuZvaxYuHBQn5P7juv9c71Ydc0QS
Pcwla4bVGqFF3rWUUJZ7+pK6X+4RSu2EcaOGt1ENlPuDdQxZCEj+00T7GTxLHm/p
u03TBP8uYv4+ag0P4pSk27Mgvy1tIhNH7O5KOOQAIFxQnsCVcBlcE7rpaIYjizWE
fADDdJUD0P+Q6eKK2/3c3t6RVgn6q3FIIiuj3KGnDm328jQWJuQB4KPEbstPtwLp
HfNbkW4HoFyjrbCf/FIaQHUTibBONlRPEL9ITkTfzggg13KwUr7OP8hMGH6Z3xhK
f6nQ/WqlvsiRHEKOtBh00BxvFwH5AcZ1oZi15ar9sdyxEDEJOYNW7BPhk4lruoU0
CH/2pekBVl3D3IPUK9WrzArCXzsbBySswQLWmRdQ7OL1mVFenKVrIMgjCxpD/M3E
aWYG3CQQwPF5O+TEMvEz1U1pmB5mfQwg80xB60weC9dS0eZalQa+U4kkgDEwo4rh
hOMJ/ZaFObxk+exmlRs2pM+B+DKe7izR16DRRzV+bf8ezZkMZ/zJtLUClv3xqBJ+
H6mE/VY/6lQbVbdFOkzcZ8PTxu0TboSRxO1T6Dcbmb2e3MhAejbrukZsTcXve4KG
25z2x3qO2fK7Yjxjjk+WuLNTCrBaG4K16dTnHeAkiEBPfZRcIQHKBnFDk3YYmNW9
bizi2N3iGYvgR1povPcjrlyjTCDiyg5Lf/ydpgiv6/LFgRSehGwbfxNRh3ZE5eSb
vD904aS3Lrswi3i943xbuVCfT8jqPp1baC5g4RwO5Karz/HPGj4t6iVno8r17y+C
b5BzOXGwMKEQ4jO1bkM0MupIhzOAtJ6flslWzLLQEruUpB9ont9sU33yjy0msPIJ
y0I49Y23JxTvEog7rI5H7X/x4JHQX0HxFbvh51Po8jD2slriNF1q1zv1BOHLispx
cWTrylCW0KbYvnym/gSOGbGBDjw33cK8VwK5kuKWDz6oDKiTT3YA6+77MJ8XsHTl
00JJ3FzIMiMLQl5QK/+w8duGAEiKljQ5suj0iXP+tNq+W4J+Ng63G0oaQaiNZjqf
e/7sAU0cC8dl7ESB71q8u+IB1VUki8WJ1PZ+uN4H1wt99lu1OOSDEnCystVx1cKx
xgNWVJAIcykXO9FRCI0GEIj9pSwlm7E9pDm6gSzg+vQiWDaH/bYX0XkwOKNnN+o+
9lNXsU7stxrB4uAUWyBmre8vaOAWQVNiST5QpBqUmpaeWXodHXL9d6tqjUSbrpA1
yyWLEYiRlkHrdFR24RWFZhTl89kX834LygDfjYlp6CxIXdI5FvK4t8qpHw/mGbRS
gHUUHPEshwBwsCGUCHFRAgoqbZfnA2R8sfLV5t+Ei0T5Cxib8KcivI61jHtXyxSE
bVutP6z6yBuZ8/SX65PixmFyRX7pDBnBRObRsbuQP3C2F9bytEWi5Hs/fkUEslUq
Q/rMUU/z3wKF0Fp3UH0VLvesZnwFousP/DfmjJbDLZGruPioj1aSRp8MQ1+MZ2U+
ovFhn4VRr+I751+AqQzhtg0+gCs+3MIPzHzwiXyE8eLzBAYP4/8eIL5bBO9+/eXQ
mVI4E2IWgLUn15rlU1jfmscMUElM+b8f7rtInmWpoGe58EAidCOAx6vbHd7hmNNu
bwuJlDUls2hOfsidMrolslRaeJQ7FvdAsCDR2Z0qfDYpr3he+KsZs3T/5z1+C1dP
JANJFw6ivg2SKkn7a7Pu324ZfZ19QDub+q/y54z4G4wAfjyRq2UEtn5sPwq7sYqa
H3ZnjhjvbHmL7gc1Yg3RUPMXlDdBRj7n+AiQa49iMtmF63e9liZUxJdeG1dH5Yp3
nMH4++hZ2b8z4bbY7at26dB0IWZ85wcMmtfFycUCcYRJNXGVX3esfA6Vw6Pp+9RA
3+T+5TtxhEQ1TLDdujCdVegCQhLWwl+R68a01ZZVcVZbZWnlRVDwb5GXmjFnRGrN
OwwTd1SjnvAt73EMnzTulywrOt0F1RFipI7373pKV8a9AK71rOIOUgBhX8hXc3Cp
zfpFoKVA/N/nH1Ew3u1r3WQOK9KBYH3rj3XpljZVHyHl5xsbBX3vMg6Hq9K4T8+A
FQd8z8VtiWtrix2qe2VEuMhC5ZVoS0xE0cOada7gImbj0AOQCKcGeb1LLbhqltKT
NfVJIuux1/1oTdrk/tzbRXAgpapz/qqnoS3UfIyb0qPNl/Wnijt/iUF4ijPrH6Wh
WTMoIxgbu0OJ6WhTTaGHtrEhK19FKrJyMqzkKSInu5hBrWndw+K1ZH9acXmAjUtL
d20Iu/bb665pYUOy2fnWLVR9wjVZFBDuWrii6/PwAOisrTDHlTTeMlmwEvf0jmDV
Nspy0NuEdYp0lqdtsOvCIYJ5DAhReeuwB8+0XUsnSBZz7iahcWoIoh2FDAkzPouh
lMnPP4SRqZ3Ue9S2CQL7wUnoH+9POmusWCW7DPtFNUS1DL1VpXXbpH/fk0cwInIY
ypfHlV6hvzl5jyBm5of2AKJ4QyMOhiGrGlcOR9bkjKMTNlVewDY3u23p5mUgbbou
dIIpQjjZJBqE65XXdjJmKz8ccp7Z90eqnE4kn3ZER8nFcJutK5B/qjbdVY25siC/
HLOnZdMh472eO0d1OfZtbtDfoJNF28m3Sgs0hxvbGV+M6kWfZtBwxdB9aNxoefIC
cRfvHdXbASuitqXthOk0U+kk0gzoiWOLdI99BE/pCj1v8SBNqoBfEhJEmBAeq7Kd
bNj2TxYgI1wgBKyFiGOI7dzM+zYvyDi/MlPrGnUZvUqtiN34kUdcA7Avt5PYQ9O1
KFdhc7wuZNFjGlNglKN/GkeYk9LHG9wDbEJc+KlfIxeMAvHZde9HgZ4rUeX/2bUy
v3OcNxuoP/h7M+lM20t27Q6qocY6ME+1cx+COYOGJZVCrPtHK7ZFXjiccrTqiYZk
gZsTcQqBXq9lurx18ND7D2k8dyKJL7PgCJ3hcVEgLxdqRkpUe5ob4/HXr/nAk4s/
+3sp25SrcyYXc8MEk2jJorA3nJoqps3IzfPFJ6dokdYAkR12QIbFkbECjPMbMQPK
Vn2XVaP8BY85BB5l1AciwZNR0OONvDcGbGC2HefF2j0t2pjfnTAW/kEE9qz1O/J0
tXD8KS3gtFY1ygCZ4gPBNd5aPLv9u807bWurtHwSxI8t+mBSHuhUVahttVdf/6eL
XfpoRIfsBtqzLT8rPz5CNlymZ0bZc2giq0DkLm/vxOC8SZ5BCj52R3kR+1HdmUyC
RJTVwvrxbUCC61XqlnKTUF6yUlSfIxk2o1DAtinO63pVYYMHpzIZtLA+uBoWVxVX
DHL3V5DhqAk7ympAShxTowK1gSh4jNeDkcUhtlnZSRR/zEFaiwaUauNOgpU92zZY
wQteSELLfFABFYYBfYI6dTpK+nEIOQ4ap9fB7uE6/lusUheCfo45klizsux+4EeD
VMRL2K4QBBDmgYeVUTbvhFkY2Uo9Vs77DWuDpBS8PnEPDtJeRe+jZG0UIyVhXT1P
ZqIETq5a6dciXKQxLmc5NLY/Qq3GLalBh/aN6BHObvFdiAhS3wJNc7nmNeC2An9u
iISZauX7sBsHKRyZdCMuKS1wG6DyDTMgWKgi7FWzoXDTPPDEuTwvJO1WhFEDMSTz
n4iO3vZPpqSUFPdR2z53rmnUtgc8DIVyihKFNpl0ERr7A0XF05I6am8muNiCnAHR
cQGaK39C7ToT4nehcwvs8kPOdKwLG7PMI2lHK0Uw0I1ZfXFTskoOLkYkGx3E2TaE
OqwyAoDXEGnzFA2VLyeaGgsjAQU7ZDicR71gg40qwUzxw5r9iVZ36F8F+30ubP2N
v4RIQpBOKOx6H3Kyh+tnXPKOIITn71sn7o9a2bWSFpx30psdxTVK87/J+Uu4s2KV
G9ojZu5g0OVM9Yl+CIbocNsQSKzCHXLlrGDfyKbL+ECLfCOoidBHslcYNHGpf1Ey
BAqomuyiPLEMWvkNRQ9gVxROfcvuNtlqSPIZkv8F7LZ5mc9dyJYltq4lGBVTnsAi
um+pPihjEGnfm55wemNMX+ljv1/MvJ4NCmDchPqZaOBQrRMfgaosTqGTQGMtPYVA
B8mKposV7UWlNAtMd/Iqe+1w3vdHYPkdyWqbGYzVSAfwZFYoXCe7UKA+q01R2yWs
uFinx10YV+PZCC4NxtJCjGPFmFV5T+oO9VNIXtyHc7BYBRtd/KF62cMBQP8uzyWd
H6V6WBT7wh0iGtkdmPm7mOA3UPKVs9ubVtA5dSEdmB9I3Z7oFIpaq0lqWZJJc3QB
Rlk/MRQnGn8RnCaOeJq35092HmFiHVOvbFb2TmXkoFZUH4+HvC3a7zGPnJV8KSEq
Yi301epCuOHRqQ6qP5DRmC+tyQcFH1+BqPN67/2XdDg96u5Vf22PZwq8iF6krJNl
W3+vbLXIwDXP4ZrgPvV+NgtcQ12yG5x6HSD1l2UMA8qvzWdBWCBs4TGROy6EeYFH
MINetxxchi4TeRogC7qfhDoGqX0K7PHPOx4DRTgdiez4o8gridMiwvJk1qk+ferJ
VEfYkWKk9v39gtOWN57bpW1S22G1yxBE3xnQO+svR75iKoH+NMoY3HbZYxhxqRgN
0yVYROlUHaqr9qe0UCP+BTBZsKlPdHqSGWM+Z4w7CSSS0Wqfd4uvz6FV1WnB16kv
zoItCw+wQquvTABJCVXk3L6IkkL2CEtZ0UKEHTNuxay+6Qz6lp7lS4pwYxuwFLjo
YKvNQ1ecS5noFXS3MhuYnhGQ3kepIXGM7w9AnJNiuzPmpoHEvYGYj8Ini5NNShRo
rd/WXtUnGIiBKDddMNVuPr2imoKsahUB7YnZ0ZO79FvLV4tsfxX/pRIHEiITloOj
SJ/lhIxDgaOKuqEVRJMXEx8m2b/+UxxPSzbHCZne703i35igfT8LZo8njDOVcget
4V1OjVOLU1fxFQfLH+1y7FU/+E4K/I65D8etmvsGweRSqSMBkp4BgnxcgUG9jdy7
hrrzU7BvF2aBs5N9/UjZLlmExcgVTMqH42VNy7ynIiYfH4NB3GG7d0HquHAzjxfJ
dcWMPVpfTdyO82IECLFgbAQJ4YlueB9YDkk8DCyqM8hDUZh4jMP4eeM+fZuO09Vr
LiU8GJm1+tgZiV+EwXDlfwT4/QXCfwOL3/DOVenxkz+PhYuuOc0T6LdytFpRBqZw
d2s1V2QM0AJiVtOfAaiWicwEoc3Sh1xCRpG2YOnYVWt9tzAHL6En4ZjhWx5gKQVi
g4tx9B/9Wh3fxScJ4qh/M958Fn53lArjyHGjNXOxbnAy3X+KILj7mhSbWoKnL46s
MLf4n2qgL4xw7cSqXQf7tE4D8yxuMIJdbmBFU3MQi0VvHuO8j5zBWgUyh/Mx1ph1
dR8Ra9XeC21Te41Y2NG0Dhc2J4vT6RTziegDXP9D+fwbIlt/zgOZ/GVuhtwcZ9Cb
JDPIVA0kexXcy0VWRgm6tTvUfLeV6ql1c3RmbM1v68ZHzViko44hr1Jndf09JA4b
L0Uy6RCWL9WnXdoIpc3Vg3c3amNcZaw1pIGNaAAHpoxARMwpJsR/Omb8Dn4g4OIG
BeuUJcXHOXUdUyEgUmNtaXpQWK/i3KBkJbqmXwaQFxiLmj0BmVNlLj9PrQvIFJWv
CE8oDqoTQuFjzj8WSF9CyeCrP0JujBU6pPu9xx6HD6NOqsUV7YoxESavBd/7ccxK
/5pqPNuC/duaRmHc9AbYp8fRve8icCFJGnh8OaR8DajJAaJrdRZjEUvvlDZPbGbg
VkJpMFef0LSzSuPu8b28agqYJrIy6wMmBgXtakza10/GD/CDHrR//S5R+v69sdg7
FHvczTsbYOL1slvPuGFxyxcOiszlGJLlS6g/DGJ0E60lSi/x7fP/tzOmtrP45x1W
patnuW0Iph+hj3Mr675TxP78IKY62ELhRrpjAgqxGBsOcrPY59pdlCcHnt7ktT13
H73uRhX2LSGEnmaJpUFzAwdl67RBWPumFXLWYUqLmBQ3tbVU3tu7wWOHS/Zr50Cn
3b7AVL5E4BIL7I52FuWcKCW72m2X8KZhZSmAwWX6Q+esEVeeP+9gsl/huESraPXs
Oh/flUg5Uwx4yJSI+D4Jrp63kt8x0HlMeIRGnth1reE9d+X8M8JWoM80xLMnjES0
d0GRdC6rli/t/EnzSQA5eCowN1fxieg7uC4Cq8cC0gU/QcrELWLxxnlgvqOCpdBO
EaruANnQFK0jz9IlveeAhhAfRMt6/hsfBGU19GWYU8T9BkccU2l8P2PxhQu5g4jG
H+53BwAtGzWJt4gOWwjkhUnWBh+EPRdTxC0K/v5+b0DBV0l31i+z25TrrRihmyhj
g1a6Aver2NmPAaMKEAjm8NdDYXHsv0pvcDu20QwlLiNvCwYosa1EQdekhZZTJ/hE
l+GQENzn8Lsm+pO0Zajo0SrERXTn94EfUJq0+84lLkuCccTGGrdv00DsdZ1Kbs2z
xDe550RowVSNWwIM+vdKni+e3W46TM1RRXFMQlLZfmhirfU8w8251NlRP1McvOrX
vO4yWpayPzXJZplLKAtj6waP9FceSQav3qkLKf0kRi53OCIWMCsjRgAtEFbwda1U
EnpKREYKg5Vf3tUYdG4c+PdUTEPBXjuVqLCmkz5UZSQ5m0XD/GDP27+YTjFe6C3b
WZB1HkA6ZqB/x9RVIKAfP6cC0oZsGGU14GvM/hwgtzZQ5czBgfoMQWE+kVwusF/8
7dK8bBm340Rsxcx/d3x16ImYQGHa6eqGLZXSOaa2pybgu9337NUvTHSKGxW/dyhc
OW6Xymb2E4zxgwIIcBSFGq+RhHk3ANmn4FPjxAr5G+M3Rl8Rwzk94Glb7q2qxYsF
m+1qLMyYx68FlC/Bonl77okRBa+O0rHXr8ecLm5IaMo1q9w36cx8l+xBk5hIcF3D
jasnHTAQ+D4+FGktQ35ablu1C6+F/6BdzLwGHLsSBOhFFHFrXlXUA281k4ZwX9Tr
MMsv9Pf69ZGwEZanLH17C819Wae/2CiFstbv50XqHgnZ7M02v7jz42VHLNJu3VUC
MH4UyJhnh4rZfm8i+0sqLtzi41Astn+BOZIBx9v48eLxusUEh7dw01Oznm8QcSJs
7w1QUJ+eq/8Kmg/KCQYPpFJH8OGaTQ10ZJP4koOdGVI1wtNkRjYmiKjYCopgjDHc
5mMJcOs2qKA1Bc2f0XoQTRENkr6mWQ9BXg+6UVovAt7320njYn6TgRbUKEGU4uOC
br5upRKY0qBVyzR/1E5SWWAU4dqS5101mh/L9ILoaTtQx+ykx8eJ5SC15SSBSp7w
HdC5Zj2NraEfDrl0fc5qu1kPmDa/21v4lN1BnGDL2Cg/5QeFNvMw3Y+RbxANTIts
31kWtODAiwbvxnuHvHEnJdd8a7IIisbwn7YbwBAu7Rk4i/Wr6hnBACh3eYEoCJZO
NHpwHB/Z3OhEuNDffvoZMr37sk3D1JmPPbLxitu9qRCneeJSumdVr3tlf/lH2YvG
d8yJ2o2LudTuh5AQToHgIcN+S12UTU/X+NCuOdwRQldrGek1apmb60A6xJ8ZuplC
ixXVrFnOWI7m6wzYXIJiyz935QB3d1DFKpxrwGMjOmSfgxb9RH+4lzZaN9t3BOqn
IHvkX+cmqksk+keTZJnisOWM0JedbgMZl87WlZOQp4pNMNxNZxRUukj2gMecfPqN
2K0+njly2EqC6NJzotDZRs/5NtOjhN0lwWB29qRtYI+p3OqVmARRtPxXImHrlkkY
WlqnYMwpAIpyirpYv1oJE5vE+ehXFivoRo6dBYkVjWCGdgG+vde8D/yZKCBkjmNF
O8ktipQHsdmgojXOWWRi8e3OoDyDE3BzVsWWb9FhKp44/vYenJ6exeY9WQspWpXo
uKJSJPMFHflxY0gEehN6th4puQCZ62c2njrLs1e8fJbK7LMuwfVCknlmPdTHJ1pZ
VkSweza3N7e6lrmgsi9xIEE3K/QvYtHRd9MODn9NBaMhKVEecwcm+PuXeM7BZS9C
Ipt3pAx929dNVt/47588w01xQ4rHVruGnrQmAKvWoG8Icq5iyqrGnYomlRq5Ck22
OVPxfc6fcD68YxbmIU++38s5J0ET23jiw+xzuxnTYUq5wbBQNUBQp15U8Np+pbMt
nfYEP9AGGchEXIMaMMC2rA1SWNc77MczVwPzQ6O/EfMP6/fer/n1fIvXeuWhHY2l
PTEuwqWaRPxduHGKVfraqxDoiSUdOkitVrk3tL6cz1LJj9skaQ5Iyp0JeWVgovSq
YCJXjs9ntCwX6X+lPNmIDTs7BX0YEzAmoxGttcg6bKdpZJbZGA8vFPvltdfAQ2mN
XeRSDRKasqJ2Iyw9d3kvgIsAGCM51hWJv7EFYuPniDI4moK6YQsfluttUZOrDUk1
bbU1cys8ft/pDdcMQS7dkAFK3DavcY5ucNGSvPMCipmTFoH7jg9rxGTAAfmYje3x
2EAB/rHEKSp/vb3jMDBgUCxlioJhrS9ujQmkZsOmyrqKFZkKSuzJKst8yYznfBVC
sPHUsVJWcJ/NO0odvV4u5+OL3WfVBdmKhxIHooCSEcIWEIMBeYYiwUmR/DopdCWn
gLcT2HizVJDbGiOsfWMIXS7TtgxLlf+AvHPzX0bm2q9Q6F/5C0LSj9/OSyYdgOya
t4ServBg3207Z/rRPtAsLA3n6h2m3Ew6h4MAfJTN5HlYQ+0MfbmsHcKoz1wrTb43
3f46jGLALJBJzEV7HG/jlnOUSNCX/JYKKQIQVAVR/hbL3PAZ5vmTQOtMu27HjKD8
xwDVWQsUNIhZcnjZZrfMEkGacw7adtj3Hw4ZzUqmU5gFitFW7h4AaSxi/O+ckY6Z
SQ+k6TNphfiBrYncyHZ0n/4aEeCGMAmOsVVe0kloMY36/y6QVzkQoOoPa/VOdSqE
SBwj54fGkePVuuRmIwa1EJrcALxxGTopYJRrWXPKcJDfEcZHl8jnoerBQzeI8HgZ
hoU+aRXUseVre84of5j35E2jmEfKW11JUQrgWWAyNy8qfx2Rq4AeqPqr4s7MmT+d
wlrj5xVOg3X4B6xUHr6CFWwFpwwBAad0o5dnbJCFHvvXFOEOsna4uiGhNUYg/LxV
Crtw5HvudbwJfBnlyGRbslUnlJ+ykxgyCRQpq3dKt3ue2NABNzCLBZjK/eicdQQF
haIYi6DhkCqFzuF2lYli76LZd8SYoowUFkFD5dnEcfuuggzPoQfNM42vjEN3tU2U
PpgEhngJALW7bgHPdjf/Zxbi5kpwu7lRXz+bRImH8RmouXRT0YRbm9Y3KtvBjxqW
+zKaxb2H3ACtCJstLrsHwDNlYjMLP/xPyeC86cULKgrSkBAYb8xEjOHGPHs2+N/J
ZYG+knkhZIPVsRGwY73A9InEJk/VardZofJF8sj5QDopCh5XP2YUrLk5MvWtNuPA
hMrnrq9q+Z9dmqHnkCTTrPiiJDHeJi0Acg1AtXoUMUUIoG2eFVTw9beK25CJ+ENy
MJlwMEvPoDTzuGtoNvxqmvbSPmoDPQ6g+gTyDHITgODFVvKSf8H1EN7YX7Mn+UjE
eP5B9DNYbW7EUkBlZSkMXwAbrtvTIF4+Eq0Yu9RezFA+JRbUBcPZpDj8yusxtYXn
sPb0j3SYWaJjX5Y6Lt1Ft3Kkhj6nkpp+cpnawl7DKIlv3BkZlPVYZrbxIonolFz8
v1yK6MiKYiDf5MafPQowPj6Xixyq4AarKq5Vd7fpX+3BGtbvI59K2R1WTicvIt9X
YbPbbOLgToLpTV7tRUWhiVyqNNnED6CA42C/EtBScXYgJr4lTZRxcncuQJ9wC8T1
+u6M520J2I/85NQNj3ScdNuDlU8cAcgOp+oskNAyEO9qpgOBt7NxlZd0fglH2knC
A3cMBdwiXspQNmin2OTpP8uAUelfruk4jfqvYAXW2x0H442U+OjzNOw00aBuKhVz
ApvLPfrMnq9ef7U2uhehMvM/8kbOcNsVwpDT24/SsBCo2FW9Luqo2VqjB9j/cxCm
FwtYL4b9OjngMqmlS8gJoETAU1E23Q3HEhdcA4oJJf/Nwf/EBJwYKHsuzs6zT+Uo
tIzo6SWv9OxQC4GEQBGVBbH4vrzX6krxVpUVQh5iY2t+Pj3uM1M/wwz6mN9L/D0z
IUOLF7hHaurfquViaIj54iAPD99MbhttqCffmHjjuYmT7omtPu7ad56KiP7fEA5m
brGREr1nFWin+qdi1Kz4WI3erOgXRYqa86MRaBUg+9PubEkSA7oJOJT/uc3r4fbZ
gQNTA2rgfXDgAS0Ljr4NadHY4RdUp5M5ML7Ir9SCHvzByPV5iWFHnbsT0fGpTnTN
5WC/KRDQ5e5Z/UxMTrpkWKQoWucV8cCuESx7O63dN65OYbHaL67HwBMILxnLZIiF
pF+tQfU7EN6a7myLLHjqOv55gKnulYWq3PxJXoLLmvPM7859HqvHPymksQAiPtmT
bavAKwekGPNa87/GKPxGfdW9k7l9i/l9DrwRBXTOCxAagWxEKzOENEUoTyrlhxcP
vH0mzet5Alb9I1hCsumQ7eD2i9eLxJsT4P0wYlPwzKZ2OufaNmHaAdxZQOO6T7Xy
EKVGAee70JSMBcSAZFqdC+YYyTJbbVePMhe3ugpU9XfiETg9HNJZ801DNvnjsoxH
r2TPIBgifiUSD9GXMKAJMGvAo0QY6T0Th+xNvQ6W8NofzjTKfI1S4uxX7XBYvGFj
Pl6+EGLCS2QDLdI0Uc5WBG4xI+nVGN3vyYpCC/6olimTxqURb2GVPPIZes8HD1uO
VvFFyHiKBoqh+qOdUrnCq8pKOlwZwKfTS95lWQNT8zDft7F66bVdpEFss9UyVAaO
SZCrOJm+OfH79LPMTuYR/D0diM5SPBcYnPgwsANHoos9m1Susr3v5kuqQy8NmeCB
lHdmOLmf4em8fib1HbKgpE0w6EnnG3DmEiO4DSLNEJAjC1KeiT3VIc2sBItNhYaP
2EucmGipP5NfZflrNOrZVscQekneTel/ZaQalbRmJyrAEQNpUxmxq5PBQKY0DvC9
j8kLGX6Rk3ql4MTEx+OszkTuZbCjSHhejg9CfBFb9/XSt6a/LGB0FeYx3B2A/tIM
8t0Bx3P+QJCSRxkl95cVbk1PM9p3VXe1Ftp7nnP8ny0Va6vxxfBFsJ4AKnQFNkca
R4N4hhufEPdr9gN92CIpDPWrAhlHj7w6Zw9KZ40UPfgCubOy36SoH4Vfy8+iUN2p
ZfoR6xy82HkGTeyVBeO771AIkXGlZryFQOLHSxWmNoXFyV1GTmhB06spaIpSjnKI
9J+hjmRtZaEMKKFpZaqX6NS409Wz3nEcMOrX9UGHbyyY0zdUwT3gO15SbEqFPbta
RASMrPOS+fXtFZYASohIMbp63Z7/yKOTnor5cWTkN/KRiYwBjW9zze7gMoxIR3Vm
Cp51NuMPTIr2VhrNW2/aT/4vpKGA88WiTxe6znzYB7n9YbuhnS1WdiBbbJ4gTFcQ
4RCo3TPttFh9pzsUznn/m9i2aeF/h997VIzQ8JCxCOpU8GSZhQQDs0n92ibHxva7
iH+TXyVxXlYinLBovAExM/obhiS11XP93Ze5+owWmFjpYZIb8/KrG9HvBowE1qp5
8i38VMBCmG7Vi+ssKVwcWHVWDUqixCSGtcurh7AZMXaxXTkLHOSGIme6WryJfKDG
B12in2MBQdpszYC1+IjyaA/2knuBxAzry8KVEENJnoFPWCd92qJUTd2ShnGmzmkw
StXvhWoJqsp+3v7JLF+sBkPkuG49r3H1pARbwK/E90tewsZLdpIISGytp+Ucf1jx
y9Rroz1ekjyZFpY2IglA42j7aPU4jJNrA0nGDwNrsjo2UtThwTCQbFdq3w+uMvxD
jl54uwMiHbp60W5syYKCuKZ4k8uMBCQusEO+KJAeU7KJ4Xf9xUBgVrbMB1NgIinc
CJQDQhj5auQLGug0HDo/2wM4K2VcaXgf+9xgfJ266OlrnqRCt4ofwBmiXvf2GRCk
3RZATguIoTdvuuCM9LPuUAlwoapYBlu3jLbs6IeYpsG1A2pq41uUxK8P9VGW19RO
vU6GuDxKQfDi8Th/f1Ou3ZG+SS4rf5MtDlWS3BFnWdtFSa3ZOf/VHzwLNj7xENgn
wQcWZUbvuM3ahL9VXgGxxQ8NNz70rq1ab1pOhpQ/ZMnS86f9lhgj/qdmD29nUBGP
eYa5bBCsmO4km7Uf/nvFLc3p1sngxC6y4NsC90AhTLuC5oRIHGa3JDQqUlEv27Sa
fXQa+9AdTIPZkkto8B7hA7tlK8qNq1cp9rCi6+6ppBedGoktXiqNK88+fgMxryKc
F/AKfNNtzDD7OyyVTaBeRnta7r0+f1e3HE0wORvGiQx8mGu6avDCUYbomEParuPh
e2YL3YJzkuVGslwzJZhisF3XlcKcW/irPR2ImkUpntOZj1/VFlrGjh6AOOF6HodE
WWDaB4wXRQhf2ZrYdYxI42/S+/bICxPlW2BrenLalC+AX8W20FIBOsm9LEST0yfA
uTShchsgrLohduNRSL6wzIFJ9//IWL9yyJgafXBtj9Y++XJsWZ6FkjdZCa7N6+UX
FCkU263bROSPMsDfwKwIbHEdZUXmXA1S1EOK2QhUrXj+2/bFsXmRO8aRdSRt2TMu
0tMRARQRMLr4KiXlHfqBzfSR0vuarw0zLmD0eIikeyBFcha2IW1gq10J+Krq8Hpk
52a2LPCDY9xdn5Z7qMHSGsaATZk3pDEeVD0j8AP9wY1tgn7drchjc9M8bc3Gyogk
K06fuM9nEmtXCmzMC6GY1ZTvIBU2H4goaVBdx8pFcJ6f747euqLpSKgYhts3Nc65
9O0xRXM031FEFBsjTU8KhPb79ibpA8dP79A2DDrJWaXAC26pF0+gm0a9LMQTYKKH
hQsU4v9/uMwm3XsGFIrv53xGCv9y9Fo1M2jmVALzT61UmyEnQQHBhVICVDYQl+Ql
SzahZr8gIJZxwUFBeGELz3yBLe3wBFbq1JiV1DKOjDtvmbCXTEcVuEVk1S+mFeC3
Lh5XVNfCbfsrKdF44H9Z++nCGh61rrITLmcBxbFSj0hq+868qaLQ7Uw5ddTUN+FS
9Sg/UeSiUGr60z9ECH6iXLBYS1h5+Uxbz2ko1TGHSV9fCDPfhK9CbtCulqCEm0Y/
B8ZM0aVoUHosoojP0NRCTQEuzfhoj2IQEpQDM2yEpBLH0Eya+hVmsqp99FdN+EU8
xOoHzxO6R1HZlJMlR/mwohEJLYeBg7XL3IT1EsB5t3VhSQtUMpGEgx8H8LxAjYGV
EA24aJWFgud7CQNWtxItboAXLiYRHCX0Zn9MJBg+qo4eh/F/JEmziSysrDXoXxsJ
B40Tzm+X6pwuhdw0OAfzoHpjO59Udi2pa/SzY93aHwHWTKvBnQFmV6eG3iJVrh55
+AfhCYb0+8VDVmUv0B6u43r1nBzjrF3rQnMNK2wQpStBWoPFxUpFwQSPYyYuHMkP
A3jp2Ups/PvmoKYkhWGIdwq8Lmh/h9oZ2FqxjXRD+6pMtGO0vPdKgBi23AF+ln4k
OwJFEFJMEDNppSEZUz27WjMLY/02/YC4X7c8TuX8K48/fT01uaC4AUfWDEm9fzzr
dPLsb67aLawbdlxqnaHJirUys2vBskyTPYdbhd9LB5BQuEV53v/2zt4X+Pw1WXyb
Lf7u+fMO/k07PuQFKsCBK4XRvZtw15e3hRFGqQ8O7N4FLy6FPbvX7vJ1bGzCUItN
FwFauzW7QJy0SkQeXraMt/aloSZYyC+WBbidYoZtCU9Y0M3i4ECPBqA+qhx92UGe
hapAsRGDa3zarFkgyxwImpYdw/SVwy+8AO2jJs05gPcqIDjhBbgOEfeX2TDsB95W
cyaodh47VLGVPEYYKkTgDNUYkgShC8/OmGoOw7aXfjyIIepmXaJ4seejmb8S21oJ
zZOntlD0CQUnTfjOIPI8N/IG6wbB8GSIpupI3zcZhuenEfqSXqe/tTxeaicmTnXb
iH/A4mbY524+Oe9ioh3IXe+FFWlxW4hCF/0AlF9gpu/1OwFbJvsTP8ExXFTp7+CG
uCj9aLgCTvswrhT3rfVdgCEBQl5YnhKksiy/MmKCDc7eEVQkhyBnzlur4vBKMdWn
nLlurHUM+3GdgjbuxCbNBzR6TA5Ll1d1S2unT2bMwDrtJXEMxPvAmXS/Ser0u3k9
ek6q87WxZom1wh6+H5lYsQWZZgTubwRd9QRHpQJ/aUEcKrYI94QHxIwKrvE3ZYvI
e/0PzrhM3Waj7wGZTB7NEPZBO6sa4le+phZWdiwVil3WAUf2Eitus6Q4t/tUABqL
q66zAw/YXdUlDrDEvlv0xM2iKjbBzFCYn4Vwg5EXKl0phDJVWFs+BbVSQe3tEUBz
gfLQqrLbae44QjG5l5h9u9fLkweYpjX66ZYpbP9+9CD95Q38HbCtM378+NSrCUR4
p2W/hPEilW4RmCkMk80PbJnIk24Hmq0+fIBzDp9A5p7ODkU2ZaIQLqFxEDd7NYeT
BHSpHfgX/73e+SltP7hTIKiVHNNp3O6I0s8Na4h32iPu4rvxZnW5Z30BPWqYzpEl
y/KBv15lFyWmM0Ejh/J69qYAocKKfa7w9MHjgb2yh4sDxqoUU3DSIkBFWi8+FZeZ
meAo82esjCtwL4ZD3R3d74F7Wb/OOxHgszDQvNONrBJELBT0J6cnEM0mVWKSwjdu
6cYvuXzRG+hg0yE6v59VKR3zwHzpliH8LC8IqKMV+K/mgU9HaCT2uzzp+m095jwy
o9sq/gCwiVogl2u8dEi+aCLlozh3Ctpf7MGW/0euCYGgSJgFFVgp8DV7LDIibxa6
SmkozBR7LJC+WK6gCW/zDElFgNhKTAax46eRanDEpPx/7e8JBoLn85AUfFE807BK
YqSHjuxnZzMA7iZBDwtlAIprNxgmj5Nx8P1MZdOOvJj/DNBqYVJo4Kw2EGGjkFSB
Q8Wyem1EhqpDESTw3PxjWsQ3fKur9QcvCmVHcbVkxfPfFBvNzscV3yQI+CACYHpA
NfxRxb/krj2/dKVCR8o7mGgccvkBEhuQDFfzEE+RT0ATQRQX0ep0q8Ya0XAijhg0
ollHs3gKtRdLOZF/wS6wefzt8JY8A3wJiAwjeSXEOK4CRn2JAbQtAyeQ+ihyikEW
l5ZESrN+iFTyL1eyw4xMD0EtOzEZ/iwxCaqm924bLmOsybDrNTSM2woi2aWaLt/4
ti7elu3TDgWzDyqMK/NgUfbnPW8yyrchCa1OzNhw0Xab7HwK6UI3LflPSObruWkR
h19Ut6OJEQcPo+8jxnshdi+0WJjtEAT09N4dZKYrnlR8eOsW+HLN2si3Le6OshEQ
tHVUzDnXZrrE7hszj+E3zfhkvvDjhqjvEOwejiiLcaB9p4xek6PBHwqzkcJ96oKe
2WEkhSLlt33mjE0xK9qBhuNpqlkYKz+XK4m3cLb/Q15DV5P8Y/tbUcRCiBQUJhgZ
YYv0fH7dB9s0XZUsoTeR97A9FbgHEFRHSmfpqgvjji7buvX0tuneTSkiKaLzf3Qo
ssZGKIfXP9ECT5Adrr+3psm6s4Y0i6q05RFK+hdo8z1uj6LwS5PBAYeSQoqK83+1
D1CzzZt5C90k2qvXtjZyZ4968sXJZEd61ipHO21SVwwf4SEVv4uzQmnyMKV+Hm38
FKrm0hrowAbbFvZ+rll6AXsedhopUNMuvaffpQQ8HQE/EqZSfLcjMMiTw2LJMZ4A
JOVCKMsxIBQRbkp0G0Y6enyu5dHyKKTqpT0CfKx5Ha13zQQOH+kwkets1zoW5rK5
SZaZHsqnJcwsrtBLeGHs0kSS8uTYtt6/p+I7eetQRx+Odg9XaUvJSrZISiPHPu83
BMPpcs6EP/7IDyrYXRlftGhdWahpA/ebp5Pacd69ALny2+obvom/10zALC0zRQch
4cTPsvpTL6lUz9+WGBbXV0YBxlxPAjQ2t3ZdahhA74EYf95VSpPJ5GPi/XVZY+OG
il/crxafvjHfTgIsrUydIVcxQFgWNAMf5KLCnvYSnfnR9sgcRIdZjmjOi+OKTA4a
1oH6zuRUaJpolle+3ZI3qdWbNZxj/MZv7Q0M4gxCljDJGvrXRKl7sK47SYO0w9ub
uFvNOdEAyT1iuongmZos8e74qTT7ZqJ/rcgVgHRBJql6QURbURXU2K2tVLHjfxTK
VPRXxtOKrUN9snQHm+nSFYW5JHvMf54cwwM4pT+0/SReuL5F2UQiiU+l57G5B+E4
TaqqX/uFWurSWx0KcesCMtYjhg9kBbciConDFNOW2HN8IBgb6lfhWuBXrZjhatyb
sMnbOLta7y++MEYrTfGQ0A==
`pragma protect end_protected
