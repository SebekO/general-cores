package wb_fpgen_regs_Consts;
  localparam WB_FPGEN_SIZE = 60;
  localparam WB_FPGEN_MEMMAP_VERSION = 'h1;
  localparam ADDR_WB_FPGEN_CSR = 'h0;
  localparam WB_FPGEN_CSR_TRIG0_OFFSET = 0;
  localparam WB_FPGEN_CSR_TRIG0 = 32'h1;
  localparam WB_FPGEN_CSR_TRIG1_OFFSET = 1;
  localparam WB_FPGEN_CSR_TRIG1 = 32'h2;
  localparam WB_FPGEN_CSR_TRIG2_OFFSET = 2;
  localparam WB_FPGEN_CSR_TRIG2 = 32'h4;
  localparam WB_FPGEN_CSR_TRIG3_OFFSET = 3;
  localparam WB_FPGEN_CSR_TRIG3 = 32'h8;
  localparam WB_FPGEN_CSR_TRIG4_OFFSET = 4;
  localparam WB_FPGEN_CSR_TRIG4 = 32'h10;
  localparam WB_FPGEN_CSR_TRIG5_OFFSET = 5;
  localparam WB_FPGEN_CSR_TRIG5 = 32'h20;
  localparam WB_FPGEN_CSR_TRIG6_OFFSET = 6;
  localparam WB_FPGEN_CSR_TRIG6 = 32'h40;
  localparam WB_FPGEN_CSR_TRIG7_OFFSET = 7;
  localparam WB_FPGEN_CSR_TRIG7 = 32'h80;
  localparam WB_FPGEN_CSR_FORCE0_OFFSET = 8;
  localparam WB_FPGEN_CSR_FORCE0 = 32'h100;
  localparam WB_FPGEN_CSR_FORCE1_OFFSET = 9;
  localparam WB_FPGEN_CSR_FORCE1 = 32'h200;
  localparam WB_FPGEN_CSR_FORCE2_OFFSET = 10;
  localparam WB_FPGEN_CSR_FORCE2 = 32'h400;
  localparam WB_FPGEN_CSR_FORCE3_OFFSET = 11;
  localparam WB_FPGEN_CSR_FORCE3 = 32'h800;
  localparam WB_FPGEN_CSR_FORCE4_OFFSET = 12;
  localparam WB_FPGEN_CSR_FORCE4 = 32'h1000;
  localparam WB_FPGEN_CSR_FORCE5_OFFSET = 13;
  localparam WB_FPGEN_CSR_FORCE5 = 32'h2000;
  localparam WB_FPGEN_CSR_READY_OFFSET = 14;
  localparam WB_FPGEN_CSR_READY = 32'hfc000;
  localparam WB_FPGEN_CSR_PLL_RST_OFFSET = 20;
  localparam WB_FPGEN_CSR_PLL_RST = 32'h100000;
  localparam WB_FPGEN_CSR_SERDES_RST_OFFSET = 21;
  localparam WB_FPGEN_CSR_SERDES_RST = 32'h200000;
  localparam WB_FPGEN_CSR_PLL_LOCKED_OFFSET = 22;
  localparam WB_FPGEN_CSR_PLL_LOCKED = 32'h400000;
  localparam ADDR_WB_FPGEN_OCR0A = 'h4;
  localparam WB_FPGEN_OCR0A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR0A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR0A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR0A_POL = 32'h1000;
  localparam WB_FPGEN_OCR0A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR0A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR0A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR0A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR0A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR0A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR0A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR0A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR0B = 'h8;
  localparam WB_FPGEN_OCR0B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR0B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR0B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR0B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_OCR1A = 'hc;
  localparam WB_FPGEN_OCR1A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR1A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR1A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR1A_POL = 32'h1000;
  localparam WB_FPGEN_OCR1A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR1A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR1A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR1A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR1A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR1A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR1A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR1A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR1B = 'h10;
  localparam WB_FPGEN_OCR1B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR1B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR1B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR1B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_OCR2A = 'h14;
  localparam WB_FPGEN_OCR2A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR2A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR2A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR2A_POL = 32'h1000;
  localparam WB_FPGEN_OCR2A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR2A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR2A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR2A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR2A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR2A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR2A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR2A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR2B = 'h18;
  localparam WB_FPGEN_OCR2B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR2B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR2B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR2B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_OCR3A = 'h1c;
  localparam WB_FPGEN_OCR3A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR3A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR3A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR3A_POL = 32'h1000;
  localparam WB_FPGEN_OCR3A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR3A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR3A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR3A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR3A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR3A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR3A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR3A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR3B = 'h20;
  localparam WB_FPGEN_OCR3B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR3B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR3B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR3B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_OCR4A = 'h24;
  localparam WB_FPGEN_OCR4A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR4A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR4A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR4A_POL = 32'h1000;
  localparam WB_FPGEN_OCR4A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR4A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR4A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR4A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR4A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR4A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR4A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR4A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR4B = 'h28;
  localparam WB_FPGEN_OCR4B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR4B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR4B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR4B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_OCR5A = 'h2c;
  localparam WB_FPGEN_OCR5A_FINE_OFFSET = 0;
  localparam WB_FPGEN_OCR5A_FINE = 32'hfff;
  localparam WB_FPGEN_OCR5A_POL_OFFSET = 12;
  localparam WB_FPGEN_OCR5A_POL = 32'h1000;
  localparam WB_FPGEN_OCR5A_COARSE_OFFSET = 13;
  localparam WB_FPGEN_OCR5A_COARSE = 32'h3e000;
  localparam WB_FPGEN_OCR5A_CONT_OFFSET = 18;
  localparam WB_FPGEN_OCR5A_CONT = 32'h40000;
  localparam WB_FPGEN_OCR5A_TRIG_SEL_OFFSET = 19;
  localparam WB_FPGEN_OCR5A_TRIG_SEL = 32'h80000;
  localparam WB_FPGEN_OCR5A_PAT_EN_OFFSET = 20;
  localparam WB_FPGEN_OCR5A_PAT_EN = 32'h100000;
  localparam ADDR_WB_FPGEN_OCR5B = 'h30;
  localparam WB_FPGEN_OCR5B_PPS_OFFS_OFFSET = 0;
  localparam WB_FPGEN_OCR5B_PPS_OFFS = 32'hffff;
  localparam WB_FPGEN_OCR5B_LENGTH_OFFSET = 16;
  localparam WB_FPGEN_OCR5B_LENGTH = 32'hffff0000;
  localparam ADDR_WB_FPGEN_ODELAY_CALIB = 'h34;
  localparam WB_FPGEN_ODELAY_CALIB_RST_IDELAYCTRL_OFFSET = 0;
  localparam WB_FPGEN_ODELAY_CALIB_RST_IDELAYCTRL = 32'h1;
  localparam WB_FPGEN_ODELAY_CALIB_RST_ODELAY_OFFSET = 1;
  localparam WB_FPGEN_ODELAY_CALIB_RST_ODELAY = 32'h2;
  localparam WB_FPGEN_ODELAY_CALIB_RST_OSERDES_OFFSET = 2;
  localparam WB_FPGEN_ODELAY_CALIB_RST_OSERDES = 32'h4;
  localparam WB_FPGEN_ODELAY_CALIB_RDY_OFFSET = 3;
  localparam WB_FPGEN_ODELAY_CALIB_RDY = 32'h8;
  localparam WB_FPGEN_ODELAY_CALIB_VALUE_OFFSET = 4;
  localparam WB_FPGEN_ODELAY_CALIB_VALUE = 32'h1ff0;
  localparam WB_FPGEN_ODELAY_CALIB_VALUE_UPDATE_OFFSET = 13;
  localparam WB_FPGEN_ODELAY_CALIB_VALUE_UPDATE = 32'h2000;
  localparam WB_FPGEN_ODELAY_CALIB_EN_VTC_OFFSET = 14;
  localparam WB_FPGEN_ODELAY_CALIB_EN_VTC = 32'h4000;
  localparam WB_FPGEN_ODELAY_CALIB_CAL_LATCH_OFFSET = 15;
  localparam WB_FPGEN_ODELAY_CALIB_CAL_LATCH = 32'h8000;
  localparam WB_FPGEN_ODELAY_CALIB_TAPS_OFFSET = 16;
  localparam WB_FPGEN_ODELAY_CALIB_TAPS = 32'h1ff0000;
  localparam ADDR_WB_FPGEN_PGEN_CR = 'h38;
  localparam WB_FPGEN_PGEN_CR_ADDR_OFFSET = 0;
  localparam WB_FPGEN_PGEN_CR_ADDR = 32'h7f;
  localparam WB_FPGEN_PGEN_CR_OUT_SEL_OFFSET = 7;
  localparam WB_FPGEN_PGEN_CR_OUT_SEL = 32'h380;
  localparam WB_FPGEN_PGEN_CR_DATA_OFFSET = 16;
  localparam WB_FPGEN_PGEN_CR_DATA = 32'hffff0000;
endpackage
