// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VxpGSyBfOCo5mUq0tGLSnWPB4Y+0XNwf7Y6K2qWhaXMzLzHgRqLLPp3WXnEyw9zE
ceYfzGSGZ+9g2XwOsvp1F/JVhXCMaCWaj2N9/UXhFfU88Fq/ZMey2lKxyPATN/5+
9ebXEbO+uoJSHkUc4IayiNmEdNHyNl7YjVicoPRQ4l0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31744)
+Gb4gVL4Qzyh8K9GFHQmksRogR9d9+J6gzFRAG9H6AK1+k9fD+RO+xr47PUmgFGJ
skF+I00WGql6M2Rr4uyS/jE9Ex1OUe/Sw71t0Z+pCimA7YSRI6YI2Ymt2aKKBtlf
lIpMEdH6k9+QFrUOCZItv9iscNyEgRc3kZ7gA0VrgVGa7rDP9v9pG7qwMVPoEhj0
J1gKKY8yWCyhYLXwikjZL1AmxNU68CKOYxsrfN54fnvHKL/htHZch5C8MhD+9gi8
PjCS5dBW89Rc4uVzLP/15SOdWb2KQ0aTZAmHhYxgW6DyIutMDSVw1TC55eczL19+
iYv/rrvq1lxCwmT1RwUCNp78i2r8gJvahAhU4H64dkFRUBn4GHGXOII1LIXVM9dD
09jV7xQW4Ek1LXCr8aOf09ICkI6FxCC/WugSec4VVKZ4ucDuYFhx5doQZErh0f6B
4X7cBa5pi0VAYzlZoujglsj4QrkpsnwvZIxJCxGzRU4qzSXhYfSzNf7jwjcYsCJI
dvKWwKPVqXua6kQvCPbI5ZTyuhua2NJ5S6UfogFIs3r4msAaNT65W2b1ybQ8RJ8a
X3SxYj62vAOwNJTcydEPnC8vBDwlXLSXeGKmUNTE92DMl/b21NMY/wtxgtrt6rde
aHzeQ3h7Gt58ZNnLB8D/Gbq4FNWYZevEoyKGfZ7M+2EZQ1h6B3Hdi3efZlVnKmqi
TslfPD3VxSo4lgnZpBxfZbPH7wBFGfqwcU2CLCPShr7jHJz2OC/HQw7emvA3DRE8
eUWzBfNBSKOHDFvBw1tDZWcjU7RX3KyQV7/6bJ2friStFhDzcPqZEctgq4ayNuM7
9ACPo5/678qT7fBv1HZ5T6/liIw2s9VTHEfcKqGROwaqZcuCQndMEp3m0iwvFzDl
r2JFsKIp8tdoPtjS+veObx2mTM3vJZDOR71OcTl9iST8aWLr0a2B47RsGMC6ueie
dXYUvfbGma7wgnS3aW2XG3DDtOLVQGL8AmJ5ZPvewvXbcCUo/3SlQPIthV1sy77L
y40SanzGFDDXoU8AuDZewuqUqHSt6xbqM3JqEVaFoDuNIYTDQBzB0/ZSH7STXjCY
sWLB69GmkqP9rUBD28ok630w4o6s+S3UEMs6ne0vln5yGHRc06Dk6rYkc6V4jmM2
4GW5qxCHBouDP2r+wrU52DDRNU+DZYwF3vF4MVY5Owq1mBI1DkNskvzzUOY0J5t0
Aat59BvNLfXGr0utoIlRAdlhaBJEYEQYNePloZvpyKCpWUE+b9TBOieFqCdAQJnn
cJsTLBHjONSTmq9AfpY9ZD9uDzbRH7jmlZEDZk8/+iS9xE7OEH5Pg0iYmeuxZ0M3
7daADY0MQDfMtTqCpqYVGZBYZ0hl/ogspUWSc09x0vhVIpgwBTasysIyv8EwVt5o
uYkaKxEn+6o4j24e6VhdGcQUEvuLfhPIXFz0gci4Uz1LngZDLk4FB2lCEyfRhMJ8
SdLe691s6EqvopHG4XaU0SGJwsBkvN0U93B5hMHblz83N1gFY4lsyuLgAgU3VBFf
ShBTcb7LCaDP5ObfiOFZeCFomGWjJt36IOV9WG8XYbvc4pFhgezeFnbFvRNPJRnT
pb8DiJ29lr4Sg/MXL1TS8IYRKpc51kt1+jUoOUVc3J4rYE5UdjvuzeTpOurrPSqA
cBvE5rcY6GYL/QzzJZqLQTwoxhHYlq3yyyl9Mvjw2TET/gHT2pmYtzH4kckJXohl
2Icto2CQDtdQK4O8QO5CM9Fo+wUH076j1y59tGryycbEkqOlC46EgAorYDt8sgit
SYoQn4R6xq7NHG62BQSVa/1RkCVkyjvvgwvittsebZ26rrh7I7K7kB2Es41VX9lB
Pr4rkg2g2SfvYHPRhDfV5Q2zG7vwHi4ANqSR89qfLiRcoHG8P5bGzBzHcqgtDAHc
4z5OLlyhSAFnmfQoaAMODFIRSKGarvWHEWEqSpDAYUofgmxsTuvzEYeEPTSlKbuh
ZDRBGSmuR7B1NsXUIX1G88+zgFZ+I0T3SSss28XJO+m5x+lAZsX7a5MuxLsHX0FT
8JVOmjCKtf+B4RU9cSQSgWS8xfYRTkApNrjhfJAG7sRDC81d2jlqxiPPAmm2koPZ
TlEzkA1GTopv3y5oOZWvlGEGqdpfLKE288+3XvMKMfQV48rVky5VZbV2piBJVEFY
PCStFuP2qhr3qi4i+UT+Zk+oSkNIX0Cv9BNGoFKGMVljFYLdKCvctd856wJCgICy
Y6aA9+QXdpZ3pp0Na4wVR5G7CkFg1qM7vnC/uTeikTSmtCotLs8FX4Zuq1DOAp71
lyUACMm2LPDhr+HTTjWcg2yN1En3kSnIr8ox3bbjeyQuBk4HGLRj152sLU5D9aiF
iuZByONlq/wqOyQsndfjFEmPZtrQklrTDtuIrWeL489rrakC2HfMkiafKQDIfMKa
C8nkxTLo/YI7mRq9RkIJN4y13yaO3WOIq26ArTC92XyyFlydUstmmahVK7oqsyoz
F/fO7VGxtE7am6CDbcj91gKz3QnWHQ0lNzWdaoDYSR9FLTAbYSKH/MBCrN3wWhmJ
9CCARWQ+zB3AsL/q76ftJjtsW3Kt1q7d4k7lP2mByQ8NuNpB1v/k7hUlgvc8hARl
OVwaaE2266dfxLmrBLgF9PBS6fWgxK16HnSHQK6RX9dOmOzjtI46oCv/ey4rp+sE
iWBx5a7Pe2BZ5oOpwM02Cdvd1PB3I9nArErKgY3+8vdl2dA1cA69L7+DOCqLKL7A
FDYF9OPHW4NdU0FvEkQ0mZg1GieTnZh+klkiLvGW027s5yfEyd5qgkvnWufGxDcF
taVSz2WCfkoOdnbf7w143wLg5iNLYGLrkmFZHr9BYJz5lmpmM9oO8LSQhQL1xN1L
YyeaF2G3L4eG8eWbkFU3v5bo+Ri+/z8412xIWbFeKT8DpthGcnyCldmlXvSay0qT
kTksYj5AhLTbtD/39A5Cr0xP27xM4MzMxdipHUVGg9hVZz799yLxvpj6YzpDjXHn
+Elu8utntB3pzH0QupayD9xFWVK5zwCnPpynaokjg0PzVopu1j1d4eOXMOggnodf
HjH+N0Bf0M7I34hghuuHg8nQmk4ZZCF96oLUyBbLnY0PyBmYIFfLBWz2PmBEsq6I
t4QhuiGJIGo3PzS1EHvXDpfG6Yo0dTEekeheNl9Y22392EAwN0WI3y/6rrZGJqpj
3ZOWl57xU/LJSNZNWbzrFJeust37cIymWxG4lV3mwVqNJiycEjUX+KBJEhffWJlQ
97kof/uxwJzmzRMXAKZnV9M69E1yKaq9H0lIwFh7d4JOZP2kezfbm3VkcXRXNam3
a/igNFliZ2EloqgPetMfAhJvk8lFhCwDcYeltMj9OnXi+BulFM5Q+sEEENgwliGO
s1ulryN478xN0yv8XFlqPUnzh+lbN8vkVCN/zy3EC2T1ow+irobPnImOP80E+WZT
nB8VY9d0K/BI1fCg1SfNYmBgOuVClmQe7qui8Jp/C6UY5APVzCuk/flLKOdhQbG2
7Q3RoypDLSlV07PlAurhdhRG5ZhQrn1ARFJJctZWUZW78YuVAIqNjn1VYWn+I279
PvAZXnb5dmHA0qtXCeC2vWTGtrPKU1VAv0DrQ6Cnq0KSO2ayvcOmNteNFUAJHj49
8ksfc1eY/0qVH2J+ZUFQcIlAKRHQFjWbpTqlkYHXDUEarGwhRg/hF0ktpBU/pxxq
dsjK4SyY6VlabkgtK0aT/K8OLSYbQQz5fx21B6EU1fUo3DJDXKvumGo6n+Ooask1
+CxZyHfzi5sIXUIdpYUkZq9C1UBKZgMG/rHnNAloXOpm3OO7uOd9MCCzduF0FYCF
k7pvw7iBJTaAd73Xyd2m+cFsHWNQoGtG3Ul48xvraw7zI5lv2HBUgKF/gZdqXizU
cBw/T5XwU7EHpfJ8i8ZcaU871UoLhlBQubg9xGFyk09c0nuZ9ArA5Gpe6fXfY+3r
KWUvdCHoz/lfCJoJNebuxje06PXGxJ1Lkr9brosYW1BhPgaa+zoQ0gC3SIbKQonq
5qAGpvRC5M1BFnJ0H46+UPmFrW7H2jxTaAbd7c3jTgfzCbRpLFzpXC6KfXqBr/s8
7IvYkZqxhVvbJf+YZ7x2IfC1WEXkIAtzANkwoKnlh4GvQioKWRHa55slJes/Hswc
DZ3vnI4SmZXArnwtnMnjSOrXkw/SDRmpAvSLaAp39jj8S+D/vVVUn7uofdTTabB6
CIPO392qrTdKj7NhuqQkaiPIX1ttmkx2LvYZa93CbTGRUO+Hr8ufmFlJzFVKL+ei
6XlX9hfwdi/3XEwirZzKNBmf0T4tSYs07VqtzeOql0gEnSs1a0prJ45XG0h2h9tU
bSogERjgJs8eDKSxsqDbbF1rRu+rq+rtwYuVuAg0gZYj9uW0fo+jCRGEe6y8ju81
enaBlQIKw1AkTt79uIBdTztOVyGvRNnE1zjo52S+cw63QQ+uxKWFdNJEsgQvJZ9X
ItbMKFy8JqDza7BCG38nKm4E5XvOS1/ou6hyqEDvimQuandBFtLFLPBI3fVgNn+i
nL4RmVuJSqTWbCUO4Hf6CGrph6HdfOFndpWaM/WReiiL2VWw2LpAx5khyrkg1wCb
QdROxw3bjYKruFWVw+0ZkRmH6Cd4frS8jAGEREBSWXaFbgZrAX4S8L1J9BKnKx/Y
DQidlPSd7K+jzS8spGgoMUlfMiV5EI311NplE4glK9EVA8X7/v0nzazfor8qUDto
F6HjtoQP+GPvyDTOZsZlzvcxfOvaEf5ELxYlfRsue+/KakvfMygXWWpPvKr6+cRr
itw18f2TujgLx/t5d+G+1+DYqsTJ2XEQQHNbSAiMkpZvA1ACdjGML5tsoyX1LMXQ
/SD11ZG703RVaDraYWt1N/Rug0cmotN4UhxFfiQfrY0PFBygCMhyMt+PszoGMdgB
quZqMjLiEBSwfk9kT7Wc12/hyzaO/+c/cZHHLRTyDUsG8SOWX71IaS7X+RYixqyS
JtdyZO1CeoYrxGgWkfeNPlLOm0UYQokIIQ/HwRm4iqs3NmJgdzFfIFORC0ogjP38
gpI5h5uYjB8S123KHOruMGih6JCJITZW6qScjwGaGSHtySsABgNMJobyL5wXSnq0
jX+dreSpJlDa+8enchbu6AaVWPXM2e+DXtcFOoMGtbQKanR7S5h2sKIsaZlgvlrR
zNulJnpAN72GUqKHSOHg/a6r7wYb2053ctP/T3oe5thf8jXiuML/PglSg9E7/RLu
gKYRkCBOj/uqmO3Jx2WUFGQuBH1iMmQp688TRm5rBLHzipMuqZT2oOZ/3CTUEXWP
0eRIZpgen7tUVSVyud45d7kOBewrm2FLqfLvwax5BH4KiXZ6hq/FUhTOUOZXyNE5
MKE92jrOmXOQAybyYxoaovbiZx8QiXkjb2CVnKFV7BowvjkUgb1ZKk13jpFMmXNL
j0PwSzlAEBgJzDO0gz/a4ZccSMw6jFXoWO+oYATT7eFnAAF9MATgyQzf0tPHwVSD
oHcCUGMvtUlr33jsByvF05NKteJLVGjU0ZCm+zNVw6VDiTjfPIE5fOgw5QapEaQ/
Sxd6jP2605oF1qcVTeLzXisYrAdSf/zQ+vf2AbS2oXd3UKEaJn7w8DZIKnDSarOe
u/EyCgkME0j6g5SZQIuvJDz9HNValirzQeUibIMwS9Tq8thXE8zNpA9EDCyDGjKt
yxfUVNfAn+hQkRISkCUFgbFXbq+9I3C4Z1EjpgQM5EmwwZAXfXl/Y339a7U3X6jN
7COeLlHWSbH0PZGlnUEjay6jqG70ErxHurfoapn7m46yQgMIyuEbqvW8amuqfUdN
GPSrwMRFfzmrfWqhmpjcfIErD3gVX4dgdRYs4hKW8pbGDPpRDPHydtKYZfFxZvOP
dtPpEQMxcsMvS0xlTUR0ZAimlfJ23C5m13BfEmouAxsppDMAAztHYBQBTvD0irLA
tyUrWMh44IEXOjmXRkKur6Z1aNySprOBfStng8BgrO0TS7HNnOj9zt4UzQJhbv6F
tNbxuclQNwESuGoywvfOCunZYRRkULtOuqIEszTgbXH0sUl3e+iyuwosXTJhJSV+
LGi9J0/25wAR3mLRB64zuxZzaUItM6akOJjOjvHqnxe/tBOC5YFWW4CNtgPAY/hU
AbkRcLqXvplAv45GbkvcxfHigbJYK7enJgbuKKDqk1VDOd79PI2GpxRhyBcV3vm7
BVTm6txixWI/BxKywBo0xNfcYY76Ih+RT/nD7dAd00RNy2ro0j2yHfuhQkSFp6mT
gYmRwZ1YFZLvR5Y2NfQOAlJbNQJ4kicdQghOoTJzX3hdv9xWX6MH1vAE/6P3wzOx
hLfp18Zqr1h+309ceZUikIrjnmuUjPWMjrBXldsYbT+gYXbKH9chCHgVNsUbz0dv
976NsokiN6W7Uy6Vx+xhjesg8t3trDmD+wYGCi7kvXXzGnAcX4K0XNCC13uwxMcY
taaDyR4l8Es8ivNF7/pAfwMCna+vp9ubUMMlXcyhq8USzdyumGK8Gb7yXx1AHg3W
KYLToUocfIFzqIBjrbwEb63nrRtrcMZTaiSYxXq6P3w8D58O8OuKA5tbU4tMKvTe
dS4Kiw/P776MtAhwBaTgLx9fpsEWa5KHNe8yXYUbic8cvdh2NHPXscDXQJMrcZxd
eLLiDmtpJDz3GNa8AcU7sh09uoDZqg4eh4sjLB/i6YpUdBLAhn2TC1K6uqeyk+pl
PMxDvq2wZm6lwG0HS7PpKDXBlCzUCzfcA4p1F1Sf+BWRdAzCJB7YQnzk2iMhWk9/
xwYoxqZFC6bNaZTuId3xPs7xL2ZyY5qfayCJkFxpCjHJn7NAy8u2uRU7kA5FQsHw
sNpN7YSOSeNHDKwTCFE9z5DymTg9QNULb9YIwRtAyen3GcVE50/x/7QG1pRgcqcI
16ZGvnowU69uubAqFTrbcdtyEtSrh8mTUwmHrwAN1ivS8Upac0Ui06K4q8xoKuuW
z0WFoH4KmCvy7c8Kih1FTy030yCWfezLohRuhk6mwclErKNN6FXkAwOY5KgcU2op
5LcUqwtSoY1GE/y2aM3VQs7vxqF8i+U4InWcH2W+uKawknnxC+hocOhnDrKG7m0W
zy9CaWKqKL43QzpoMxkC81TnICMsBQ3UZd4RQRBOUX1Bf6wSb/kMPDcWMgUdSb7y
KoRg4mkQDlXKk51FAbUz+fshUTqFkQY5DDMqZdzhEYdTsI1WCsA2tGXOC8aEwLuA
4GY6w7BRnqTih8O8rsUNXpXwAfgR7xiHF69JUz4wO9mImRA/BqLwC/pk5PfYNEBa
7FxGMZvIMdXB72GWnS9WMK2RQVATyVYWFbkMOo3PKCSJi32kzjr5HxIXlqMmTNqR
N/RVzuRaPbykkcq+nMMNwTjuV8JBUO0V0BNEiEyt62S57BZmAV1mzLxXZjwKnDXI
CSAyePDLqlRUR6twfwOZ0xfd6WUcxrod6IP6a+QvRKguXqKZVgrZLTDhxTMWWvju
QWFUBFeN70WUuyJ3RkKkkVb9mSspeKDCBbuvzpkXP7RuHpCljIJxSyurop/EzeAE
qPD1P7BGnVCdgSFcjGGtZTfG7VoQbs9TUEJNui1Dtoc6A9FvKLdRRlO+QhHGDo+8
/71EUUZBGvY16LSbmlIvjCH3DUNFwAJJqmsiboCNjb4RcBpGmtLExKd0mTFzMvxO
mFj3skcsLQk5yrlYJC2mPameKH728alleIEWBWd9GtEYMXHEgNQsXES3nhLmGQuT
knllt3NhD6mUl+g1MpzPRTU9wPYPlSbVFHbzNnS9GVS+XXibPLDNoKjZpPfrii6f
VL1PpW2r7CRz+z0iAkwfcUrt/BB/VNNdCNl16509x92uo83bBzKcE8elPVJzoDKV
iUmnsh4UQ5i9FvgyjphBgYSrWhuJ4BMUrDRzier870/38WrzsewMTQDWRTgnREnU
+deJAaYDVWI2DwW09WKDEwGxjUVqKlXE8rhMxlqWhfqY3io2+jFuV6sxw18LDmjE
9IeCSpnJI4hEVInzKc604uHWxuAE1vaWsgkOO5nUGcP2szBXamcaLLpAF/n9cg+u
xUmc02nX7zVkYBcFA7Uwdd36PchFToxKVXKCJXLt68zYeR7HdVWYVNgZfF4Ot7lK
12hUGjHt7o8pReuXXq2EXvfeqU/nXHS/ONIRTIiVStWEAGWcFA/W019qIoidNSDi
qaCdp59893l85HkK5ZauGu2td/VkTMJBu13wqz/8fcoQAAzOJbDYD/xTTpzxWBBp
VYq/QFMq4J62Uv3W4+7wm8mLN7IfHRQbCqHFpFgR2ersmPqOhhhSqxXsMIkIP8g+
ZHvw2FC5Jnp4f4RcO7OMcxmZlA/wjUl2koAlSte6AJyEzWYmINahw4cl8bm7cyYR
Wnw4PGLexKxDeDnJPqIsWF/jEED2+wetKtMe2UhNWLqj5yNdaowQfXxCbT9+5N/C
Yv5uDmSFqopH5SG/JVPstNwL3mhO5D9FyqQh2ocudjZ+6YdegCCXzU7WksOd8TZJ
HOguI01C4cTTfstYqKcOnFFFIKNXaCKgauZH2Il39MQgZOBG6mbeGF9RDfNwTEGz
MunhbUTXzcp8JBOGzBnr8JEyzhzdMhRRtv2YvqhumgAgd55qaGBzY+Q9qbFzz79Z
Fg+ahZZJ6SXCI2DbOCxLgcVNaFifYtBvsqnNvW9FQkvGN7FK0AFXvLPUrZI0wvIV
nO6HCOkvW+wYKT7NHC3JX1XPVo2w4zhTTwN/EJ4uKd+2aJoM1p79mBqzwHixnvDQ
OnjAd5+qsmJXtHOENfh5+QFiXzQAdTEyXVD5kapiwEtdjY0+2Nu1ptuDL2IaFC7e
z9lelsm9cBXgsRRhy0cBPUYdXQvVm/7NMZzBwPQeIccwd9vwwXwNt3GB21yoCyLn
BwUDHK26G88pkmJpw2VmZdmleYsf6O2QChayaL1WPkzC+d6XlTRLaD/lANDRdNcQ
xhvRc0NyElRJr4CODKmr0/9EHY30gwAMEty/t9K9tbh2Ep+krEkhtW1y6DGrbgGB
q9EhIqe+36AqIsQw+g4zdXlihe8zBE4MxxVfcWi9ddosV2YMCat+NXYwVzuCKcz4
5E0f9OWDekiXr26PAayZskbMuFne6ADn3Hn4+xEuQ25Y3HI8jFIzQ5/1nU92YSgZ
JeCHLonDWA+gPx9bDinAya7eLC/uSvRWOQV38UiaDnxy0LVnpX+2OvydCpdxa5os
rMGtDoShkESe6MSr19OOwbvderaN/6erN8zEH4D7NGnbYRbk4RZAzkSSu2Wdej6n
cECD/gkplUlEtgKbyCyp+Iik3RXd8TBPHRk+cSP5L+JMJgb3eeQObgTtJNnm0X8R
72ItdCMQ28HhBChDVp5UBSKOYObCehcKALFV6RG5SWejnf5IvCCTk+pZgCX4dCUc
/eXFcev19WEnNh91jJRNNAtF5KLCH6OTpO/+cKF313oRVcnGhBgNXYkZcrj1q30G
l7hg7xWU9At7GSLyfp4mDvsgOlY1lwg7oD1baoQvoEJK9Uw4gD0m50icbEm7ZQD2
Yl+UCGwx39Zwr8XcdIErMUc5n1jFlLS2L62wRO6djI4DoA+cjdeq6jXpqLeWARvA
/+/nRNeO99uXL0VdIrab67CMDTBpPxJewd8QQkJw6cQeSMJgSXwfa/85g8h9Ml79
Z7qKEOIENlS+JPglLGAryVSjvKYqkpcvGr0MAQToIGi6yOC5HLLpCfuppDOZODYi
qG6Aonih/zZlLs+wkYl536NitgeMnbeb4e/EqBHoWawtdPNYsvQuwnfwRgVysFdK
N4M6Bnl3PgDMRc1Bdrjy07tIhowxfruSIFOfusOf5CB39UCfjnvfp7gx9Nxuuebz
k1JHjFpKSM6hcrzcOpyfIGz70RnM6wDDaworYu3Eahkg36OtAA6rNMq4zLxy0gzW
YkOvG6LZcD406Aqyk5XhX06sz438zA/FNGlb6pWs9EztBZIpdt+J2lbYW6Vh9qwM
E4ZQuactH27YSsbm0h+Eniq02HlZbyNFMJq3Fm45I42Uab0rD+SxPFw5Fzo0Zf7S
tQTPubxHpqHj2YiRyaNxahFFq4ChjxFITExi8xrFKLGhr1kHKSPIMtHTXaSxDrTz
D8CtAfJrkxMvPe8GVlR27bc0SkvhsLkcQhseuzjzaPprTxck4Xasw5moQ8Ivl8PY
ULRwB1J0lioiB+EhN+YgT2aMw9b/3Zre4XJ7gVoxOtH0gU0YZDcIGfnegt/KG3nM
g87SpeWkSXUVkLDyVaHex5R7E3upDjUK0ebEFqZFpur6TFjQ4xJTrBYLSHskF4U7
DFwBbgtCcOTUkVIVCBvjRYS6dgeXPQM/51166gAPEQyr0YjRmB4pOPOGfx6iabCy
1kQCdnOXDAfNbdb1aOpzCIftfR6R0gozknR7A/on19w1db1SbGripEoT4alAPkWI
Omd0839GxpxZE4zZvvZ9nuqtBHMn6ncBoDOFf9VLm1uCQd06qM/cXytBbp137Pc5
RVw764nWc5zVvx5cQHS+xFKdn+aHj2drqRecsPVZhTPfZg83FQ+Vbesu1Zg4sbyI
lIZ+pAWYCWcZYhqFdCxAm702bEIdpTSecYnL5E7FdLVUNI9WlqpGS0POAZ9m8PgJ
ZE5VGvVEryRCkEVUnhJu6moK1kBO6iRZTAWYcdhKoXc1jrZ0BTa+G8ult0YIklZD
NdQtABmSdKbw0rhpUhuTC45Nlr2oGM09ipHITkn+W2XrOjDBFLXYvXQ3QaTf4BXB
UumnugPCpmu6VccX1y6TaYYQiunPi0VRDXQXOcw12QIumn4Mj8ZzRcE9RBY+X4vQ
BY+sqMH0yGmiRtusIXoCFbZoniU4p1LATFdPYpuYHXriCorQ45xVo/aE7ZOLdSyd
LGuueWdthXXROsrLMv3OHVgojxjUQ9YPyQQ/ToqephMRNWnKx6tdfLscreJ87r8V
nXGg2E6/QYrHwD69loopvjefV0Ji7BbxPMCGyV00NRBwb/EBtk6ACe8+mf2n7ilO
bnZZBIxf+F9tsrLSIcd0JXyK8npDNEI3TX11UfpkyCdXn8odIu5qlB3DHxGNm2Dh
c1ehHffwzekK+FQfDcEDAFYtVydquKbUWT5mIvQJKyrqDXPqqbE+IP5zb8ZXsbyt
moPr01MWdpvhrxcfO6VPwkA9CiteUUEHYcXBfkyJ79ppVr1alT7mWHPoDj5VcgRs
KR9sDmu4SH2rp14H45lbgHSw1UWgb+8hno7o+g5PmqQQhP3BdiB0K8fNn8NseF+E
yemmTtigWG3gNavIQKsOoNkU2G0UVufK5ZrU4F0XQbPzdR2ZA0fcARuDKQRv0bFH
BhKoVmq41hyQFWv/FRKl/bGEJNntSwoP3FrYb79Cxau0cLvyMaZH0wGkklGAHa4N
xKFenKkRerPnepMe5zh4s3kEsmpDaDNTzgS9KipJ6B2auRQZnsVRpo8kpqZHhE4K
3RqLyYtdv6l5lYES74O7Gk60SSR3Hh/A8Oxnx81ui2/jhXF69VQST+2C0zh0VGhj
YopIC8nT3OZrKXJvph63FsJ6uhUSRBl87jNjHNyB1KRtvXxnJtY1SlYY4JApOogQ
mAcA0xKRydal5OEWxpRkxUTXHX8vlyQVW1mohdmVsoibBvNhC22GS1hqUlDCZiqZ
YauoYiFIFq3y1GY91loqqg6mB9bpTDgT1WFd/OMOOkYx+Jr72SNjltJKXmvYOExe
nCMmgRrfI9UgTQTWq/LYtBCArt8jRG1MqSJqVAvNGG/50ZG//ivskUqVyJ2tn486
knCVK96troVuFfPK8uoQncnE0GwuMM19U2W0TdOxTY9zksJHGbyTylro/3M+zn/h
RZ+wPEz4SVeAXWH0N7jaoZ+mzKHVr7TU257ePKur1kd795spMLM1YHfRGCCSlhxh
HZdc8d1ItA7AC04HK8WdUhdXws6QtS6RkSQRGhsPBQPMv2c3a5I0BnDhN8HQ45dB
288qCWavbrB1xdNuxkt2iyxMUjrHen6o7l8mvIFEsPFEs9P1H3p8mpOG8MIEJuOr
hKhVT9/+tJPCKuNeK8GYVEB5VXFPppGWI10eQv35zNxa2KG7oAQUF0Fx1MfLPEja
41CGvdoOTt5L5NBywZSfNmqewuOreK5yfXVEv2zI+/nHaAYSpI+iO2wIVqlhd4QV
gI/xxCnJhmEaeQziE3AHq476mSEeWF1M8K/zjnU0jhKZIw2oIpT8qKtY/UgsvkyD
Atxr9YWL4WYxSOf3u3C3aAry/9Suqpv3hNMASJI6dBe0noMzR9GA6exorDATw7Zo
W8epxSYPF7+1sH8LOW/T6XQwhh8aexh0NlZtzPtSml7Cat2knQdTh4qm4wfXRmBh
XDoSDG3P1ysWdGaIxusvZ1723Pv7znGeWBv0+DSY8pvIIMo//7Y1Zzxt/QtqIQvV
+Biv32pFr8U/Xo57SL8vcqt2Lu4De23E46RkqJiFnefm6pjLgW/EhueKR28PcX6Z
mCcK5ZKKi/aysmnG3Lvq7qiIzQcY5C4ILrlqcAN8NQuF4duENUfSIsOHjRJDxbTh
taKtIkE+4fsFZvMZd7TrJ+eEwiGg3wNROISq5WX/RDQyJOMKADQSlrEobEr6UU+k
n75rS6K5ZascTOcjR7HcvmOZ4/sJiVxBdqWWv+qCb0zfYJHz0bq6JL+dn+CF8c59
Z6Sph7NpZBpV/mi0KqirZ1WMCH4DS+fUPQeazKku0Cbu4yiRpBVGSOvvL5vBulZp
iSXr+Zp5v73iwkf+QzvlTtQlFVZLFUPZO5ZL52gIIBS6ggm/n4LYG175luSXJ0Wp
azU3Ay+1V4j99gN7r4C9QjTTmw1Xpk0mU3q42QBKSFmc2SiC4O4REipxXWmgjS93
v9IvejCUVs27gYT3rnI49AX4WgIOwSgxaVI96mNGqKGj2gwy3iuSa2BlTcQXqcyC
H2XHQKa7Nxuq9hnxuStQCIH2bHHWrnnS5E7ssxTKp4UeUzo7WjdQG8XgL20aztTT
phyO4yBf4ABijooC9LmiANsdtbIBzt5o0WVKIrCGjOmE0txfqf+CVzMb5UO0aprP
KvxWYk2gmuA/ppp1apANyR0Svxo4IsFBd4GpJmLljMQIHResYxLLvoaCF5Zs9Cu/
WtivfVS7k90D/I6RzoXdp3pvsMM74rnhHQIXhww3WEtalXDHLagDz2vJu9JYlnwy
X+pffD7EjbkVMJ03IXzH+LAEz8t5wLrW2/80gFwP6m1AeFiCYeiwj2YEgSimkV7h
UD5FtqTLHEzWxZ9DfE1AdUvyCuJ9BPD1o6pqKgEju43W7tnBtB302G83unrgAYFW
e+IabQf7Jf+jtc3JtYS/goTtyfXS9T2QDR1h9b/xWWmcf/TuDtuOQbJH0sk/HheQ
cmjU3pRbQGa08SNRiljw/OPry9xUS2gCSMAONdue05vKGctFGovHOVF6wluplF/N
pfbMpDb7fvwLQow6yQkEVxcjaJ8TX3aTzzcUGD9X0iMVfprophOb7+A2DzSMWBR3
q3CSdSFZXMYwZ24M2cv68VtB/2xbYoOnwfb5ixCtJ8zDQ2ILJtteJQ1LVkWMnoql
+s9e+VpCIwlNaYIqLVHZ1awA4YDdVAyVBt9AAjB3fpGn6NIAd+8kX0QixVvLmTSc
eZSndZ8JCibRkoxYy9gK54yQdr6TK8GLckMSz2/LFP3GO5jZDr+xyyd2bHwQh/VH
ihO3yOLJxWrJI3GeE4spbruLaFEX+DcB6TBCbID3OeaD06/pjN8QgzI0UFjpsujR
vSEEDrHt9SfAvEXAQ+VIMq8Gxy2IQRUESTD7xb1thZYxMrtsmdiwSfBxlWb/n/tI
StEGg/3HY7xE4VDUPH9mn7U+Ge0NI9tFJjWZWyrVw6r3XEPNuEJus/DOjz+iqQbM
pogHHGqQ7exmrXAqWDS0cGctCnUjv2z8a1qAAHLhzdNqM9cmaohuLiikSY4QD1yE
JQmVsOg2vUD17u3MgeBQZ+w+QdkubM+8S6HxlvKdDaL3BpzjmetoijK4YkUPEInp
FdcTg+cpy0S4sdFi9LsF1fgrSuII0i4Yy3ZK1e/ppwPj98ahTtSoB6zju12w5Jsf
gq3W8YpUPHL5nUGV+9ZEeQvYzXUQhMPHZ66veQELqbTdNvvD5uZLNPmS+SEb9xSj
+piYPTisUgjHT4LFHjzrY3JJ9Uornn1NH59DFqBPtlYVMjlrh8a8IsWiqUdyFfUj
LWehI32OaqOyySVYI1u95COTUmmodF/fl3ODYP0Zf7FnTrTmVnwjCBWslKalLeRn
7/JMKdfmQ3NKaf8Gwg+xeYpv7kg1A1JMzscX8JMW+yIDAbYHW9nTTVTOmGqCvndr
tX3ieP88QtWSOk+DkLle6Yr4Nem7iIWiDhuUxtBYz+4OgfNinXw5cNzlBA0qZg7S
q0HMQlM3GXIs0lLVL6uFLbXr9Jt0jQ76tz1ejeWlhxtmrZampQ4NeKi3/n0IJXQ1
B7hTnqxKhCtqGos3UOzDAkK4RbhQwASyx2+3oHNfXCjc5hG7pp7hIaMRl68l69La
gJYmZ0Lub9HgspPBWZnYp1xRdtMt+wwk7NWIRDt1g/xBF16ZTD64r88Y+VZHjIut
1p5/Aht65Sff0z4vJjkfMIjUhW55ryecJyHW1DsvTXBlhYIYnrVaK/axkHmt/L0f
UboIGTizdeY7OI0BCOtuVBIF8gCjmZDAuobmRMPGvLCEtfQDa0OWYyQ0hmqoFDbD
3N7cesAJIIPJmxQrUUSlgZa4P2/ZMAjpMrqZaPCFTEMlIu38hztCjKT7SfFwpOBf
AJV8tD4DsPd1OMzKQ5B62cXED7rTWTEgv5uDRD8FAO7V9Jv0/oSXdKJcTIjRyJ43
aYUXWMy32myy7qYD5wY3zCaTNLuUHGhR2kFeggPlFSUF+UUrAasqZ9v0SLrBAgm7
AglSw8U5rzT8IKvxCwlWI8JXFr84J5GvzuBzDSssXiOyH9tCKTLquZVECNxDntYN
fuYO0ufpjo60QFjXHcIqUx+TlCQDpEm/Cg7mWvJT/LF1IkzIZESiSbPrZCM2zjzO
7H133Wh+TM589kgekv7A/KbUyVBvjR76KprJRLWQA+KtHwh9xm9kEbYJEwcsivxV
CD1dXZnGu6U0Se7bCRT56ClOG8ZVS+x2FYOXIRjBPgE2XqaFEIVcMTS1+G5OgaKi
JVjJKKzWjelORETsTTKjls91ePHJuUMvqe9+6/J21jb7UxVgXkw61Eyvomp+cG5e
A6rVpoIj8TJx7OogYOQPRt3Po0//KzGXdbVESQfqwQoz7vHfCC6YicyRT/Q6HUdm
JzlPHlvi+MlK+UN9Y8JA70sZCFvx+eyRslQmSnSEGTP2hweN9gp1Qv7XG1trNVb2
3+tgfUbbobrvRGv4DkrDBVtkIkDJ+XhiTgZsClTTqRhcS6zkqy3Abj/pxiSdUKfo
BD1fLfEr3clFcUSv6w3BOyAonJHxIfPaYQ+QWxlEYaPr3acoc9tVN0puEmRQmOS7
XTuw5Pw6sedkFyA0Di48T78nHp666LcEkIXQ/yU1DUv4TdpHTBcToyqae4YdlNr1
Bj2vlhjeucgG94QfGhpB/UxvP/iGTOgoX1LfWbnhQpKnq/RZtZrFJadm2om9xHIC
dmNh7FerPkqGBTzdWpxBebqdTGP9OqjGXqzMtUxlzg7GBmH7eJsTMuRJIxpOZW/0
alLRuljbTl8EMMGI6FL8HOPHLqcv4gQZ+FsCdLAjKjq2KUy6jJfb/JKFFfaQ6D3U
wrqwGL6y5uexZb5tydFWJH1LkJpGVgIxKQ35PmlSBdQ1fUT5/uP5jIB3UrEybZOk
2ruS3V2/NGCTHUEZfv3OMxIyvAk2qrGCeXz57CtakyM+FCiHsCYS/eZk/yfAnBo2
Zn3CbAxrSHQI9cjWh8zLczcBrY0HwLi1+VWnbm+cYBMgnyAZhVwmgLFJ9VWqM439
XTGHm0aQHkLQtuXjLopmfrkl+ypkml4AGvZBxQtpMTTaY0RlNO8Em4EdO83XyrFS
3/3wlCaNWLlFyJANBVGlTqzEcBLHRrVdojfSBn6I0VgXI0pUlfjg4rnTDp1IePlS
LYL6xt7P5UwB7DVtZJkFyfJe0r+IuxNK7LmnXvQa5xXoTH4bdBNvX2RmgbkV1914
8gxEr1OtTVHsiIL21MGRU4LyQlZzNJRPE/qIf5JW3Etc2BOJnhJ2+ebOOYVTT/Xq
65GefcR5diwoet7CqtwYXBYtPSUItznlAWBD0feX5t7D5i3CKr+yRpWu3cd3WPD6
C+VQ4130fB8Nj1MWiXQTDVTUaVZ43KkPpZa/Iya/uf1kaKT9OP+6KiPXaTeDqIbW
jYhRezVm4s8LqJ8nThgV2PI9IolDEoW9pf6xIeGAZk4Mm9zQrgXvbk+gWNDF8G2G
1sIPO4+QNCYwtIBK/OF3ymCDyiepSvCyAHQm5CGYPq/vcHD4CeKCNNe7W6uMnIyu
VYGKBqgYfr3HVm/tiiJpm4qkfOXEC7i4Q3Omz6xSeqs9s49KMBE2rn2f4eWDeOQ4
i/pDV+B7cjS6i4nYkoTZesNrhRRXdZNRyFZUH33KLzwtrFkNL/wGjC4hGcHie7un
XTrH+4zixWnJyggJ7JNtxfrmgMlx3qPTK7/PqpbR6hOXVfQeWVJ6+WVjHagPf6Qk
RGMyC5cjk4LiBgO/5+mh62Ubi8jj2t/+qTwxtzLWnbZDMA8GZPVDPb7z/L4yscHb
UEM90X3IR+h6AmzEzYc4p+QJt6hGMf/XUdaWfpQ+d4U7WDP2w/6yrxODNe9AgB3D
1kGrQer9NzPDI07IfSxy7WOD2oDzxK5SJcwcoYXJ1xr0aD/qIpdSU6wWb4m9GiU4
SMkhzpk/NuKCCueeH4ge2vEDRt0AjLzwhrgQGQ40J+/flSv3ulCGCGz6DbMqUVEl
5aCEKz1TYhep/ni/vJU3EOELslFAByTHUYboHCikFBI19NEzDTxqvM9rVOvBFqPP
9LLl7sMpBYTgWTpXfm9BMMeE2Czqk+TNQtgmO0ZVDRJZ396TVEg56s8Z07R9EVFa
qrGcjO8S3wPsG/BlKOEjcd+dRf4Nv5iGfo8lBbYJQa8KlIfdK71FMCC4AtXfzHb/
s7w5oco6O2WvjGRLPn3BWp5fFNPY8iYviRPc6W80J1+iw4NIQ4HulSSbFRD8o0x7
39K9+y+06p++qgUdk8Q8jRcgx4jDUSAw2Q8CR0nvLUEaytOvRrabJcbos38pWHCE
qZrnjKLViWQNdxTdRKwZAR3GcuqMwbVmHMavFGCTfDkW/9pEgI5zpO5eBZM3cR9K
FstZq7m/vGQcG/SyB/GhOZ+60GganWFDMq/kmXVR857eJ7YYEPLAvwRrwFQd7oSe
h7dIXDEYLtba9sne0/PX1HZ7XrW/TcJrWRav/qnMsC0MwFIZOnq2QBQOiBmXkeRg
lvTyDHG2GQE4luktBBc+YP/l9JJ+0219g8iCbdn0KZTYQ31aLF9r7CQVUB1QM1VK
0iKM35cW9G/oUdXfdHWT+tNUfTXRQfcBVyBhszvy2X6qT9nINyik3i7czT+YHa5Q
pJig66bR1EhAwHzra3z4+cW1D+wX3o7RFVOvV2atA+3VTajuU7LjVbbTgjjdTLiO
NOwSUKi3f503yiXxX+iIhCaeDdrj8Q6VuTPKh8GIhIkcgI98ldqmNSW70/ZY/K+G
987VG7A5UtkhjV97i7hhO8kQmI5dotaRyzoOTbDwZ84BJ35H1RE3LU5nTT+KPak6
W3wmZAzS3pdaLX32inELSe5XmNuL/hdtc+6zGdHt6tT1BE2pMNHYQ78GGZQQeZFF
JH+8tECYLniQfNFtLjYBK7TC5j5uoqHdbuQA1Idamth5qBSjbhrHJlyJt/7htzJv
FiX5TIW5NKHKqnGAM0mA1qMt4moLm2hRtaxcIMeSMqSxbrxR8tKB8qMRNT/DybJr
eVppo2IL2zQWiTP7kihxjZQIFU9o8dUkhmoRZ1x0Hz/ORlxvTm/5o+59j6OnFBaQ
Dg4BwqHO3SsUKG4okbrR7/vTXVC4anPcusrWYoDRNMtbU4zbrJ1XN6g0qJBXJ7+/
M0UO1d5xSdDkKBbU3+xyvYDBsHHkxgcKiRgQeA+Z9PxL/Hm2M3ZjkZK9qhjbN8aM
gXDvgpLmI9PHICo2xyUaYEEk6kTcCQYCNA576rsswhpqQ8hGCp9X23WcnIfNG64g
2gsxacKnbnkW5y6XCrGnx5T2H3mYwLXpczxxwMqOeTdZV7Qo/HtV8dtZeis2ZnIX
VMEh0/h/qf7RNMWonQ0lKogRLgLsW1hAqRlJhnxBN+QOwfizvh60bHuEnnIiQT2/
pGXT8xvdYNe08xs3mVqBsdkRKqilGxceEPPVLr90Q/axF5JU+RLE3g7Igs7yQEdK
5Mx9SWqqWdMdAYBFbfaFVJZ1pTMilMmpqhePVMFUMFblFlVAcPJmgpt/E5eLNfXl
Aliw1ImA38jNq0MCSE43O/cQqGm3rl00fM0Caedcy3ROvqYWKCgy0yY8yIAh/0U8
vDvpQ4s6UB5/f0h+tN+825fQ0hADUQH/3dEiLzkkj8kbu0wthEf44ZbznudQWvHb
OMtblcDXkkY1TYdcuovQJWli8v8OXK7Q7PcYPtmU57Q1LfiZen0x2ySbxUvyZcNH
CaeyeBpu5D25JexIZ3JxRWdMYiNh/djdjdAjw2ZvTTduP7LoFHT+SRgragt1xC0g
YBDrOJFMSmdvQEHZ3QROzFcYIdWOWw+dc/wMj1RAOS8qhmvNbgWA+2KlKYiAgWT0
htLEUAWR+Xr52I/DbdkmaDLdtq5C5BBJI+XJvGDf6PJaAyftEbMJ85hYiPvvVNJv
mb7STMwnBHsEfhCxLK73urrLkK9DDRZM6ejPgXgQmkgGOCXeDO8IzziKZso/ywTd
sbU2cozQvPSw/EDwLkfWj6CdFX/JRQKUHc2ryMBmK2l5DoiqR6hVOkUm++jWgX8X
GFHezoIaLXOaqI7eFc4q9zlg0IECjQkvp5ivsnRWQIoE+XqrfpXHtWG9bseZIMB4
sqeVZceYvk6XdvZcxMD1cOqoOUJzhomlD6WW/r0oHnBr2SQ8p01wDJn/JrtjJJET
H2h+9gkxJWBkP/tQCxzSvJw+Asj92VJxqDrj5DEoiMsj8XL0KPU5csiO6DODJD2d
HlH2gCmTcQAGY47kwCBfIKHePhDj30kCY3T87yyg5zKrrjfJ+LiOmcpHCBcd+LT9
VE7NczeGOVmLAiLE/I/6Yqxfyv00l+06sr3kvg3YLwDU2h2QzHSuQWNQZucgr74C
v8lxzHgbnd+PxBHWA1GrPEDBaTv9j3W0Dg5+kuSyJb3dt3ASMamakZnTCuFyGl8J
wTKbgLNn++wuYd4IiEG9MDcozBrLCC/yDt2a3nRl9edma38b/8SBbHhZsr2eSUb3
QwK8W0uifIe8C4IDyTq2CTal6tMTALcGcrv84tIQNCfaDfsyNotyDpX/dXKkIQbn
6MU0gjso0pHqR1gOYQKLEuSqlAEicZ5qMsxyHBLfxR15PBkCOn0I4UYilbhpwR8i
JI+lGgyRSTJw8LRZ6er+ofdHrTtfKQXfK6ayodHm2PvqJCHfCMRE+HeJZQbcdNhW
uDi2NwFTYQ/7qZlK3r9iEPwn04b5oKyyoqAtlvHn74ki+f7qpdsIP7/bZYaXAFXj
WIjrc3UY9DYS77CKxP+794+/w67PLADDoWhBeu5IXbXdvT40mBdvF75fVrG6Xwhy
gfSeuLKvlk/KZ4yr9w0F5dtVhSHQ8Sv2MsjXRWkB15aMOVdaNlfXwq4AZvunERIB
dZfvMOqjJWjPVy1/96m5Bq43/4MDs2t/BmJU07345m0k9gZ3x5TMHfZOV16EYum9
pg8dFgbCj7ZKhiiBcMS1UGgHZckvuA9UzuzGLBwp7BhmocPBDAE61Hdhku0cOM4t
oVHLuMRNlUoPUtMWzTNwYDOk8g5XddhxQP1JdgNoqvyWqrZ+2mtstyORfnCDc8BH
+lsasLtir/vwVvntHqipIeYscJTl46gJs/ZvST0W0QlA45gx3aBRvFF/Ta0e5+Io
WOOYjwrJ7SmZ7W0uKvB7UFJhkmgZKs1jRkWXdTfpbR7SlujLuNxLt9c12vgk3sSv
A/DJ0+PJWPwdYIav9mCrFULDTbCkRGv5dcUY7Q/m7YeY02vJhR+SFrC7FS8/jGGA
kPh1sCi/yU/iRRHiJmPDclv9wuYDDEE+1kJKtK06WSVWX1Ws9JPGsFsmGGaXGQLI
wZMABnJOVw+Fs/QH43g+0DgS6A24uzEsCc6AkRYQYZhqv/2lZQjhigSdbt1MjrPT
t7YAfhExhtuq6mQDEtGEeNCc+yB4LMJjscQnrYdVQI8TO8rVW+8YO4G9MsFhFoch
5K9BkJbQb++iaKlAr6TjT3h+92pw9Ms1eV1kApmxPBclL0FJFMliSZ5ehzW/6a0r
C0/eDot4oGN7S1s1NOBJbKfOT6f5a2tWXvDNrP68q8euufe1KsulPESaKehL+mYs
QJU2nbfc+9pONL0AwUgu2MsdiMs+DAO5cOJ3o9CHTWixMAfKdHSQnAUtNL7neDWi
AhyrikzlHuhMBeCJWw2f3u+afEqTzuSG8ivVDGWqaKfsO5ToXp3WcTkuFCHA8XkP
Hs4xO4+a9/GrKe/y6u8Y0AwB0y/Aek2rj2ac12cglXaFdtN49XBtD1nVltwE3cL3
zNQn0pPegnO0+4RQYw2d0qpHEbdFIU4I0DNJsLBKIkAgua68TlI58vsIMtPRXl4h
WCK3MgyRn7EHthHRLIn5hXNd8XyKjcAOsLYZP+jQ7FKaAiGuUMI2xXvagvTa3xEY
nHrsj9afqL1b40/N8iId1KQD20pW6JxKXLxofe6XBzirhbq7V6jfk/W0x81eExty
6eWexSzOeQayxdNL0Ixm+i8WI6UmHA8Z4Sx+bk/hzKeUF5uL0CmJZuOviA2eYd+b
y55+/Hgdw3wPEOZVvC8KFI+r2jBurALDwNwES9umxPsB7rqnP7aj67rLViKBkqpi
XPRJq3ruSHPsERouoCZ1anVzocsxo/vWDMVz2gNBKq5vX23cab7TDWCHBjWJ0vg0
T3jDxv9ewDJuP7scVMgRy/6dI3HfSVfRa2yWpgRXGZRygB0DP659190RpBr7BCA5
diSUAUcwibqH3q0YI+MJ1AS/2T1oECxbvmt5K34MsWx5D/pJjR2z5iyhp10adDO6
jqDHDtch49+f0mP2d7v04ziVqT5R36TBuRrQYpc/N3zltLy8KY3Jm5+H2hKSZzOh
Sb892nbc23ug0mMqcSg4goKt6ccYL6gBPXeSw3efmDDHLUJPRXkekz+khAMz4bhH
lq1DcpVbiRMXPnIY1npAPUyyvBCKBMCg6GYfBio9K8Ue5ADcRWo6XJ4ivxerBjIR
yZPU5nSzsVn/sK1LUk4gBaWgVay3L+Uio1PVr0f+QfmZabtLiAfMIaO86mhlxUMz
OkRCTXWeI1bqERaEfqc9P9lov6CMIf7sDny8fdOtz7Jt7xU82m3OslDut8H3vogl
xaNB+cUzVCXPh7bjQ8Am4wci/ZlxqNFyJXi9BcWQNJDOGHPUuMnHC76kc99Xx/B+
zMr8aYjRC9t8re/51hZent5DWAHc9kpw3jdtqVyNL4GK/8ToUV46Bo2bEM6Ub5eN
060Hz9xCP9QR0Iv0QiCkQfCpooXnQ0NXBmhnW5CGcDr/ZxQ7XZROGEbSyt+HyABw
kOndwvpgCgAXDRPY4pLLDlAzAbxu5ruyGvN4ocgRnYn2ft1SAaO84BUtq7wMzNIN
7z0er/bAdjFi+Qc0izjipB5Cq6GnNaE1zXXp6Qza+6hP0P5J2nUstYtY/SQWOc5Q
wmsJ8KMKk9Tw+QdBJDMUhpjVBxO9VJs4IecBYYOj1jU5dJ1opIqoFTwvpfZra5lx
SBJhf+DjmSbfEbuk6KJtL58PpcEz9KgyL9JzpOakqf8dUfZBuTBtWaaaK1JeO/5V
+96gzWjeBpc+8nv2cmfQk1+SJwQIwvZ7jEgX7Ld1UCZAgjhsCkJTvLo6z+qNBwSc
I3qptH6ckXhG6ym83rlmUHXdtyFJyq/eBNddBYUH6oj6fJLE1+L0+3m2PbHy/YrH
HzDbNcqFM4LW0ZK8U16b5YalumRR4h0EcSjDoA1fayUXFO+6rnHMzXW9qajTON6f
Ia3GkXbaUFPdzdhKV4aqSxcxevcvunGd5X/8A+VyRXrkul6nRJ+3fv4shlfTgOY+
K8AvVKGRkwZBb+MWAuvt80tfrR+CtO1OSzZFIIGHOif/FTVwPa8MgDxXBWne7oCJ
6bs2ElYEVYTnG91nF7E6vbSrxGIvh/39GDxHsT5TotCV87dcWKitai2vsmNsGoTr
tXQs0jZ4t0VYbh8GDSlSEAdOjmFWkMKPR5Zc27FWJ8F+zkVbYCE3tDFc0qV9NZ+K
zYnF4PxQyrDqiZpXcDbhzPBhD8TkynijPQfWSZwdHjZ4kXCA6RU/WMYX97D2LKro
Eza3GT7OJ1Afi76enZWQSKBHmnp/musZuGlhwJA/EJ2M53XIYf1MynU+BtVw/J95
KSohAtixQlKGIFuAGUJCTRIzXDEhi2fau8Q9wl2yGscjgfV9OAEgYMr6oaGPRfrI
zPl720JoWgr45MvxOMsGGLxzLIm/woVORdhZNLKQkVvNksrVO7JI0UdD/p5dAs++
J1nkqClwWAvEMLWuComk96xpJDW5CsE3WG5OdZXI5AIZb1VJW/IJxtNxr2TMtqF2
Gh6y49IrO6ivQrwmAixg/KfUZsj1oyKd2ksL6daF9EkeVZspOCwUuqZJRboKx2y+
CsWe3bckmYH4pp+F+cT/Q02ikBg6eLGgea/QhRXzYhVjsJU7HRFmKgFuaowmk7m4
KjRkTHuY1tVM3FoBPNmR5QD4FkLTRX+9yRAcWLmrKtfRnItAw4iP8NsQJkUNHQDi
mfRZARlP+BA2I/SIuffOse/ik2Iq2K+u37fiXqVS2r2QWozeA3naFZe5HXzCVlwm
8wdAGRTkDt658+npR8nQC8SBIvWWd4sMU6nrYosfn6odnb6b/fdIJgoQCBuVFSUC
K8h69qQXO9MitKv/bjOmpD8xuQh1c9ZVOnRCilic8xH9dvsGesSd37ST+ywS2OO5
ouRKEGeZEpAYl2q5h2HO2SOKKPhcvsaC/fRffqEMS4Xypng8on3b48Zb4bAre+OD
loT/EM/sYl4XDFmxXwdsXwWb5cQF6UM04KrrXnXyE69d3k57lJtYwf0ZvwHGRywa
Xx7uUCtWbyynAlGqC78Eq2YD/ATIykQlGQabdKTeKoq0ZkuA6j/nHzogOd4pIYDI
lBRh/7Vxx81SyZ7YxTkzqR5A0sheD4TDx99VtfpFhUD/9SeBkoc8E43KKjWyhaIO
69YT/WfI9dolfKWysTUG+q26va9a+iUxg7K9mAbehFNLjHHKszV6awaqe7KXXVdZ
oHYkoO5I3w1q5HZI7CQ8Ab6381EiC6wWdqyvjURd6ALvMyNcivx5CQgG0M+ZmZKK
J3ROMkpxQKrZU+fhuptDuskJjVf47FvGfsYY32WV8ogFdqWRYkiKcqMAHtwcmcmQ
WZeg3xN8BL1uDMlATT2NoXeeeuMHSEoRqobwaV/W/mEVftY71PLrYiTfhaN8xAt5
QO48kZhasF2HHJfi/xndo55NWF8jyEiIalksO4eGbASvrS/IYBv35oSnxyOEzYhC
asJ6E3f6hujV3U4OLvQUuRM9+M3f+QMsxztsV1OK3+dQ8xxUgX24v8XWzDcT6gww
4WrZML0FugQRLdGuUhN/4lEGza83hLt/vBMup0Ay2V0i6FwpdjXFxUpay1BEE+7z
NpyiCbcmUEnIXPoAyC0zF3lPNoMPamycCGyjW5HyUREfb6mDMOObj6Wc03cp2sGR
XVvXbjsOpcL2gY5UKiK5hVpIKrtM7PtPBNEZdPhy+UrCYs5cZplITKWY+saXN3vj
8MB7eXNNdvb6hau1YFkoOZBRN3mnFZUSs5ciFqQqv1vp+l1a7lXxn0vE25cQBV1X
LpXDuh+v7l+wFP8ovWUvRjvglzcDe2u1aZXl2YjfsGi0cfBnz5C1+Qa2V55N9XQ8
TJHBjkK1CIvnTEOKuvqNETqyw+oJgBOY4EnYEmozSqW4k30onr06ICChrNGwBWi7
fdUDzwXL1DDWwSj3x7jFeyOV2mOvSW04HJZHwfSITTqPtdtJPDUvLsN5MoV/0k9/
8tFBVaxgaqxgW2igh6dExFOH/06QHVOV43vV86SAr3pdYPGf0riwqLx3jqFMiI6D
t82N6aJkpQ2iTZVg962c4aD+i318awpDxvv826aAuLK+yMfQLpzfeL9WDRJBnvST
uX2lWKsaD2ETgSBoxJbNsyrF8Lo2bVes1kfwYphqrfKdX8cjrjLqGuZzhblQBGjG
pu2HijqD4DeEn1/2h56CvOZhKvZyG9xBJZ15jaxdCQfXQze4byEvaeowv7U4K8gl
5B3A3IJBG9gxVpPwOLOvSsOoebkpam0Pc6gqotEeuu02RniSrEmxJ6X0PRzaZxPf
ybmWaISkXtkadse8v2+nvSZXCaaagfkOfP/PeiTIjqUiuGcxCFZrulY1kzt0ihxi
lGiGb9lTKjdY1j9/DVZOhjsVRwnnrJVELdIUBReeotoBCNWTv3aZsXuSfWfEC168
prXdi/oBYb4jOGE8VGjywSmbnhS7zNZLN56dhecPSHYGuwvFtlLByNj3MLUlsZqS
h6Ocz6BGZKtHlfAnB/qNLiDLvLvjMxcFwy37m0hLWmQ02VChAZHxFIa3fzyPPViQ
ElrwutmHESG6qQ4tf+Co6Q1QfncCO0Q4GrcgSynw0RqR8cRiFYNQY8ckTjAnETH8
YhXvGvf6ARVylcfSPTTFT/6c9zxjZk7gQh97jOpcfFb4aR2fiuDlW6m0Dim/EUYj
D8KUEaM7IIFuTcwDy/MrHHTopjuHiAf56V3zPsJn8oSCYefMPk2BfAQKy8GvwCoZ
jjYFrVaupg2nohUqqJaoWDElkElQUeH5lN03qWqCX3JpEhvuXN0rtIHJDmUbW4Yx
6ycU96oXrN0IfiGtjSxm/ibmHZKrQJvisoTCAYWnbsybDdcFcQJ1DeMxgXKbTcPl
HQmd9Opam3pbp5TzcqCpI+jqRk9RNOck9L+sJYWuey+13wBOsIGY4XpWFqcz6g88
uK0EC9P0AycWOlQTsI1qBU/iWaJhzDUHRjGfbxJa/O7sgAXaLxYn72XLOcELrKDv
nErch+NeT05wZ7Ku8RgVunBN7GZCKGA2/mgON/PvCsi2TYWrxbLrGYPcbaEjQIyE
wuIPsDTfjw+NMhTJLzZwPt7GQZ6eYc+B4wBc4dbtmi5sfk/QJCBqSgEaIfrnEJ80
ELMH/ciNFbYa4ClH7ThWzK3/Oo79a9gpHZReZDp3aakp8gd7A3Dc2j5DG8PL+bKV
AqlqRMoobYgNgfPaucyNQpZZ4p/sR9CNceFje3H/+CMMy0AbGBnbVzj7OROUJdI2
SdP8nemzWZHa54UQS6pneW22+dIz0NWpkJLCzZMr2fWtpsFGu2hZTmeloXARCuqy
xFf4IzWaCrGJhUw7Oq5W6cxgKMq3W2hdzrqkr+y6qZMT7if0T/i53cgMLTFWyI4X
2GLxv0DcMIsf032gsOPamjBGKvxtUB7lKRjsK6Ny+fClav4r138voqmRQEYjCzrh
u/RSy5tyUW6ODWbXhM+ObqXe9FRIsrkg6tIQ6yVh09W7MXxuxFCCyt5gE3VmMV4M
nhPXuz+0ALl5cbFLQ236OoOuoYLDykBvJKse8vB1HF4XxtgyT7ShFiafixrrCkq5
iEo7ExcDTFMkzPyFXpT5jaYSJxgOe6bEeUNFUPhAiX9HBwm3QuukKAJY9abcxvaw
eFcBBNIVoPb2CtJOfX4bojc4JS+vfL7UjQ0Rw3L8Rj6GNkUv6QYQFLI/YOcVqTPF
ddIeMsUJYUUpDeG/kK2PnvCW51DdB7/yCyU6J1kVKfHwjEA2py8Xzvnn0HSXTr16
94ujC86RfR0geZsQqIQyBCGMK8Q/mGsyOqkP2Dh3fnm9vqNafHvXx1g0mkC/k/P4
ZLSt9bXpipMAA7eIcZZ/SX+l8m9yvCgMxBuddz7dJduBdTCtOECBWmlOoIGUaEqj
hn91WZVmKi95mUsaHRik05O799U1yQdm5vMoANp2KfisVqlYnaKIti6XDKuPx+1s
qAcSnlCZwIBoJ72JogcaquVBga2o6JJSeIN3+veEYQqDcy59Ytk34AZjUMkwphk5
gjhrYtdXJMfTP0LxIbzD4Ds+U/RpZ5hr+nBxxKA5C5v+YmdkV8cRiUXnhCDhVpat
vUYMdXX3kiYR7VI9C4yOnCoRu0E/bQgL1rPb7PXIkN5uyLQRLovYdB+jESFGBbVv
XvHYfjHQP8KXUY5KVCem7oyS6clnR6lV3uZQ0DHNkdtmpQq2fvx4zU0uPO4tQKsg
3xCu3qPa3xmdQrJwfE5WYjcsKjwwueXdbZpo+b98AEJp+bHag+EB5SxWOY29+Bo8
fsOmaryynFjfVMpzGciS/8ePGHA6k8hNeQgfT3zNzP5X2gfVuanyw+5KC7+/fa15
QiHHP6cUWmbYjsen7U1GFb1FWhnpmIDVz9pGzinUeG+JGHmFRzZV6gXt3SA0ejZs
7hQBSubHKNkq/1w+uD4QegPkimVctEiUct0i/nezrAVXyQ39qups+VjF3ibCYlPO
Flh2Oy5GvWySq/5kkr1WxHKbwzekG4CzkEzZl5bBVQr1oaoPnPuYsHuZLwS5XylQ
4MTYllccD+xVityCVThOm5oNS7zVcTM5sj9oza25GkN1pZL7DR38tKg37wZBaW3s
DDBv1JA63GZJvnYv33TWVl7tvZV2lqE0uvdVCWaw0ELe0cg0RHs4aUzbSEieWREh
GE+V/F41Bi4bTvwfcGw1csfNixf2SYucv/fucX7jI+Wrsqp2ur9p7FNpas2rNADA
oJ1RfH85Ity3bq60jLowXhh7B2awrzEqOnqz1pMIosu4X6ar1TwbSVE7WW/aqWZ3
QtsWZrc8ud+Ka9oKzhwEg8qPmWYr8p3mYMkUHG65tFQIUsQljK2yAmYDscfnbtvC
v2pG56i+yamYgLnAVV89qrl2xkMY5CJx0TE1FS+SGFLGjixGojbNejCOiENvir6C
UjNRtzevFC1PkHOwZqgLgBlJ1wCq3bYhZNkXZHj/H/g7TSgQgk0AUjxTudJuCohd
Eh1TTyjiqviJopWtwzMuJddz1LuFVe0iEVlRDxRfJVbIYXSmnNeaimpw5j5tqb7y
ppKpmoRmekJAIkOwskYPiIT1lL6FF6M17hC94jyOdXF4XyR8GfTRqCEMtQtnx7p0
+VRoPHOYYToqcXU3MhtjlWA07Wgo1IPsZi6I/6NBoYJUVnk5KAiyBVkaWNnXNE5v
0UrMZ7ForVDXepdxA9Y4fnbJcU1psR0oYub6ciEK8wWn1NfXiptvTSJ3CYL8qpLW
qxKMBqjWujzR3yfondV2b6bfJiM9Gngvo9lyHVRSFUZdCQZ6bFDMZWlIlpN0fYuz
orRKrBRll1INRaI0sOLwK9qH0/MnBfzEm5LYBbswYO0G6XRZ20l4JBHE2FuxU73G
/8vmAleZCBMXDpP7/2W8VRpoOcVGpNrGW84lY+pLcsWwn5Ad+ZngKyDqcO1rahuI
lX1H1/l2lJeKAOisLcoGCjlIGX8XWVtg/ziqFMCeQVk/PRWILlUBbTLwEN1Mt8wF
nctFduQV5qC1e7GNrh0s2MncLJxq0CJ7yt4Q4XniiIuL4sl5/tkZtKiGLeUZ0Svy
ZklNXwjaOAEn7rSrjGnVN0CIBUmSdVHIcztGZLa6WnJHxnrdUh+Ad3K+FauywDLn
m4kbFh/9lDO32ZLTIRk+nbIX5haA/gVh39UdAy/JCp+0Dw/b4BQbcB7XFDPNAZfP
G4fNpoCuRNvbEFyz40rAcqoQkxRk64tfGMGbVTHnp69R526BCqyPp4jtrMDxpu8c
vq463sbttS4W8OVmq/cbLQD9PRqU9A3ififUc0xhxbPgh9EgfxqoV/yk5C3fgVhR
8qNAb4xLAug2BBm9DI6xa8gmqOMFCV2nkSztGrcbbV060A97B5P7b0EMwbLkjWOs
Cdt7aHjgSgwuNuzBwjAMQfOQU5iYHxODFrTh+czKdv4Lqj5+oqAIJny6AbUyYG9Z
32eYzLoVrW01hyJHANOq6eW3+PX6zBUbyb7cjpMctWDw+259dtdPUTBVT79xEHeM
juwm+uoWg1E1X2zYX6KioLldYPaFkL5wEFNNnNMZi+esMdd9sYM5wViYl0n7wlcb
hLclrSGFT0esK30uyjqGNSqcQJxJZ81fSBpxHSNafO859Kgn/XX0wg2Lv1m9eLpw
AVMlBgp1v8nIeJDQFPMtxRKcRe8Lnf3uVXd7MWMlSSC/IN3HE76AKLXGKW7b8imb
ju3s8dYmVikSIAAaR27aLP3tkL/yDMBFP1xpxW47NXCajxh0yW9hgjMuGvF1THSZ
3wHrG+SbdgHJQBDrDEQe2bwD9s8qhuC94ER+/PP+AmBC9diDAZKFAZGuGGRVsnsm
XDFcNz0EICwKfwIPyF5iKhBLT6ooBp/XzPrRI9eltLFRkxQpyvektlpfrPBYX0Od
lQeZBawS9+7tomlfXnp3ZvibLGeGm5aCdiYWa4TqdHgXD09zI5YDTtbG5uKT0BJW
L6kJSAxAShZui8RQhri4GjMtH9HefJufzV9ClThdb+hCiM7DXOvjfCn0Bqw4SJBv
mcSU60OgdERGBlP0eaDyPCGt19wPT4BeIDzBC/XUqJ3qwA677yLU73CcOvXj80h2
o4BpGyKTCbPVa//RNMcRd3qC0/SP5spoHFwGLWKLoDdlyMz8Vn7nmJNWLeVsl2N+
tBK55j7w6ZtDHlaFQ95whOV/NkK0cACAJ4LsdhEo5HAqOwpnYHx/lP6WRAAEaniL
a1L/y4HUexIGQCZy/aTDEDaim9iafPWTXiCvQMNwkW5y60djEhfsuarjN0quInix
hzHcOZtGybKVw37sAOFpM+Sn9sqdDF39VeKpMV3xVrRSXeyFo2sOJDXVsWpA5hQI
Yiurre+fhnRAvjTp3JIBAJb300m3VoOnxwS+npi1CbZmfulb2+4XGCUs1mrpi1ZG
gT8U2kMO/ScslaEttsKl+cwqTh5ZSxlydIgHsFgRWt2V6WNb2RQ3TD4xpOhRarnD
f6l2A5bJSJ2B2tQEPDel098ryyEwnkZq4XU9/Hc9lyxrouz6wxzhCl0kGjNF1w35
juofHp0OfDCQTaFNAlRaq+WozQrIA+1fOD2kzZ5QEO5V8/sNprL9VRx/kTAteNhZ
8aEPRyH7CQPKV1e9NLwfluOzMWNifiSWvJJDkaNoitzjbdn1jb3ZN+AgOUcxXp7e
l5EPF2JnzMCAT09Tzorg6/sYITABVJxyd5MDWRL+WcZXDY3RP1unncKnocKcOEqf
oajBeRD8/gmn1nPPBO1dof+7tC3/SF+rnUAtZGZkoBZIXhp6myv/FWYsjmdSdAbS
1+mxvR/I05NWaLNQjMIzr/JGWSU6iVYTOmwdtJoM5XBNmMNg3ZDHNNFvD96kbISg
g6zGd8ZModpCj829LlXUdNF7o/yEbZ78VY4WwNRiN7192M+ROrDz//XD/MF2TR6j
FKSGkn/O6+rBw7kQPpPNJzWjNLX2GwnMZvtukK6dqHoswLm+rOKtS5wk6IYCw9Su
Hhs/ZsbMwNMEjBQ4pM2Nn0qyr4XJHnTtnFLAM/tNby6UdmyGY2D5h60oEBd+dHvD
E6/wRLdBpkyTk0emXBEjXJuRwzUIsSjPRUtKESErsWWIAc0gWxuZARr3hQukul4c
NjvPLH4lX4H6zMy4/XvVT6fmJA4enRFTL7Gg8hwRIblCDnWU0Y85lP/aC31c30Yt
OGbTeKEA+OpUVRF9C0c3bVlWir9ESPWihfXcdBLEVCqUgo+Q9vxNp/pX9A4YPNlu
VJicjV/hNgBZ75HhYNC2ATNbZVIC4m+FvZAUhFpMtSy9qN+jvrViy9VsQFT/mCrx
2vvR4pAy9qaOkg9buT/C53LVZqu/JvFv1blxGyMW+dyYeWlzpUcXJNo5WLfYVEA4
yFr8LuLVJWwyHQw0of+ZpxTJcHP8nPEQFfW/u13FLdoZTbbYNLAz6Ttwy3jvpibT
pOaAEAZclEs9wVJqFI0vJfJLlV5gligW14ceVCv2AMtp8vD+k/+uEHBaOprwa8Xb
9xPU9/Us3V3+isNkc5DuXyE3W6iK9yv4SSVSWaT+i70cxMzbVlpn2wY3UtiOE60D
I5zwgefqPMzRB2lzKdBAnSwArBpVTebg+gUr+Xh+wTVtNWTpZJZ2XDnhH6vNuFTU
Fh2UsY6FT7C3ldwTCYTFsULPwC7iN4BLyPzKdX3YXilsdMRFwVa8ztsg2IW70VUs
BolU8+92YiE4YzTEZrOkdjsaz6z+c9GZzBfW/woelWBg68t4gWxg4ZG82BCbT0fn
rg68YLram4ejVsV/BEMPXDzUyagjtEuItHED6gR8rudhjqWP+b0gKkYcxiNWiqHp
GnXsRyqgk9IZHg42iU/PVwWq+uPYxdjtp60n8zSGSfcnO/OvImC09DTqi9osX4FA
Psh1BOc+kXbk1eGe9liJoF1YK/JWc79MvAnQ2bVJv2XDWUMvDIn8XRi+NOMlu7t4
Vm4dU8xKf7HecS8XZmfeWl/QuT0QksB1Ffw9p5v3vnTpRIk6BGnF3Oxcd7r9TLzU
wGehooJch1xRptM9jLo2Qm5acNUHXoR+JgTnu/Sg1/Duko6iMjAxAyy5+iFbN/CV
EVzwpJRzq99Lfgqll02xSY8rc7+ZmiBf8cMeUk/dsMBs3qqGKbCa5nbAmjVEKucW
O8jM77SgIXFmMtzwgCO5znRPgJctjuIbdlMu9awQg0sYSliLU5OAiNvTCrwLyvIh
98sWcsYmsogp+aVLojmodRpd9l4Z1NVcyGKqZAnalm5vZYk6jD9lfLtvb9y1CAlE
4ZVKQ3qIAUYZRgmEQEWKVTGDa67KnGzwRvgojpK0iDEq+QtE8xRpDwscQLNBlvLN
Bq6fuQo9ju21irDmz6G2zuaQQ0vmJrH21CGztrGCrPvjx+JewgzObA8xeQO89c2w
E2Pq0UrahX04KIapOZy3mpT/m2ykzkEm5kOz6AxE3CI0bAK/TaG9J2daGNx5X8cK
GCICxIC8pMNN01N7lsRb9EHR8Cy+QHgPhJ9t64Zo7Tj69LxvTx0RGxam1LXbHhPj
+e+OsmGFkxqBXX9VGBrM5GJd+CpcTqb1EJJyE4bVRVdUcTy9XhpxzL5Hjz5+fhKJ
rD0gDW+kCtrLfEbg+7Ad29EgKQI8qUzQjyBlZZ7CbH5bebopQ5Up5pFlnhm0IO95
NwY9nkfNwrSpCX/zD3MgCps88xxJqh2omS7C20340d51fooJs2U11Oorl7y/yhCq
HdzGN2XYZpwGgk8ng2tbAT7Y+AXpMCaaC62HjTMgUnT8z46WPgzEYenOl85B6bLN
qnj16c35jW5Yv3FHsQ2HXt7xg51az4Lc7bemKW8toJLb5zcvT6iHXSUdkBf9ippI
xECYvV62DTaRXuNY6Q/M192HHnn4c6JFfuTzWMFkA9PI5mb+3SAui1Gr/PmL0ZPn
3RpLN4xrSBtiYSlP10Meur6+HBY1pOcB99/AGwUxV6gCKQI0luxqH5yKkfUhhBp1
Stbiqp7vODMnj/R+yIdLPDypnFYNDuLwbgr6qaNU1MdcQWiFdQJeJ1PW0zUMt7E1
9/H+qgbS1HCJvlnD3rW27tQt8h51z8PWQL4uyk4Ib5eqqH1sEJrq3h1TGFlJPk47
XGWtAXGxMHU1fHrE81gTmJVomvPcIXDMDRgXvK63sGyXK6UdN3aFJFGZE4aWvU5R
KOB3WbJjRZedUhy9HWyhjGwmNjikohqWNo3VPHN3GySwR6kU8QTgkCm1r8wiUdmJ
+XxbGLKf1PbBA5SyhJjeMDvARYo5cPyMjLuvd83KxnTNI6BZMAsVz8PeGnvZJEW0
PhA6E1OZTwODbIW6kWeF1F/gfMSWcqqTRfoOFPmfi4nEoURRKNpG8hvjzVnptb/T
RA6k7cz40kiaYaDw38Uk1cJOj6ZPE8V//maIok3Zkkd1QtuG6q29bQHU/mdBh96L
4e2Lf+PfkI5wNZleLAANEuQrQndLR5psDFkTblDm3HElEV76vwL4bEYRsVDnX+vJ
GBt6MaJouP4SRRifEKHucntURR9iTrfH/oYmMKZYug12HVkWEhWP0Fy2sTctf3my
Ql5eiSeYGa1M4uE9KnYajh4wjkXgN6CfwfF3mg0EwF+XuEoDm6fxjGTWW+9Ygw3f
sp2tmDFaihXu2Bz+gJUZAa0q9nJKV1LmbOkJTIbi8YlASxA5J8feZ6Wk4qeJhOsT
4VpAUoKFaPmpSkAtp5JFLFzk75SMMF+RHpgJzZw5KY6XLzrY0Wq4P857to1v46Cy
an+pf+nngKty80AZhWJaCT/9CB2EW1gaVV/hz7jxxWgv1uXvgLhF/u47CNRyjPA5
wAA6U+TqAkXdvR1nVk9lx3p/5tTmIGNmp8BIPRPj7/ehQR9FcQWxZkhMRG5l1u9n
H51BWGRFaH55Zm+ZuqWN+uWfOqV4QDQLk84/VPE+xgjXKe477+b9+o4yCH4Almhp
XadsRL6cbJQUpup/9mOtzAgZN365IYSbbLxYVVaYY3VstJnnYbCyXLoH9QqO59pO
bDJOkJ/7jkt7q/WKESmy+xgjwXsGwCrxmdgHxHrY6JJipdXUA3B3U7gr3CacaTJR
S4jTOYU3keMKFwJo1i39L4dQCQ/3YWy0MZJRmBhH6Bc6Fo6fbYlSQjisgy0F4ZPM
IwLB02ECH5G0b9BI6WzXAme3CTiISdodg4KFNbyU5SjJ6wZk8y1/9wiCBXkSdZ71
5b8aKZRaER5Zfm7ZVU730OR+bnlryMSm73jdEi3yXySf0r5C/7v0A+UtM550ZX7d
BSrslz0EJlcv7OVHj45ieg39QNNXKa5jAQbiO9APcUf7khAf7NZQ3gW/FiMJnM+l
yNjC+bR4jSKz3TNg/MXdJNLSFEbKn8xX+2J+LJ+yZfZeAFufSSOtqgbAQUEnjtv3
eOFsuG1T/2FzQ1VAdNBHtkDlp5QPjGHWuN2Oq+93pj3KmnwDu6UvdwrCz0/869jg
w+F03rNaDZ/12uTUiiTmsh/j90XHRvnvr9bHa4mEyOVVGWefIRvmpUR8MLoDR70l
mkyJ90BOGdeq+ojKRMfR4ayA57CYzdLjjDC3RJaq3cq0hod9C8Qwc9faZjyjL22s
LNam659bQophhEMdVWckmz+GBqYGqdddkKF2pV/8DxyrsqpwP4bSjf+u3parFUIh
1RAvdHlpOsEC5fbs+GPbmjbTOF3J5Vyi1Xl95++o5SATz84yMq9dUzhtn3sHFWe7
3arfm8xvafxBu/nxPhAlFxmcIYx4baIgLyFehEj79SYPWx3SLzsISJwjKM0FOxii
RrDkbbSJOD4n2BF9KyzkCZmw8xnirgX3hjG0Js2aBrBtXjaI4z2PWYe8Lv5OVN2O
0nYMpl0J3aaw8bFIzkujZ9cVKuHaFTJWEAL5LnJ05aP719JeYx0lxgxLJluaxOIB
x1uf//4LoRTlJ8WjV+HCUH766p0G+0MFbXWDx/zBN2xuEvaDGL3QcDR3Cg1lD39e
vbqudtv0uv3gxXTKAu17uQPmuCALeVSca5rd818iaCjrCQtDyDbz+nQXFyBj8kbD
9uIK5cQdIHDOio0Zc3t4t9qYFhMj72ykLP4KOInRqqrttKggrpvGtELxdyN4a+Df
V7ZeJChj+OCKKYyPUh/9YM4mOvsoGY53s8B0wfChVDA+8HD3KU13digO2BCTFxd4
eDTW80ASq9RzGe0VUzyDY41gmuSF//IXtP+o5AexENDADg94mRlcmRMs7hkJgYuV
fb5/aHqLzmumESrYppgSKJQtFsHYTDPZoUlVtd4FFlgRyILO3PP/X3D1FTblMKkq
OU1pkCxh5sUmLmEyjLRChcV0O9jw+duOrQuB37Je8NcwqTCle9RzbDFFKArhtS7Z
1NtJ9VpGwMDEfLn2yVKlU5WdyY5cwXDwBLngLdQwFM0jWEO9hLgpjgupxWY9LV3o
/bIfIHII4HytcqbDPCsMTK1Rt8U0XmHrGebp0ohLlhy/N0qWNDYEPAtsYzPqcp2j
qkPGJUSnIoQA1jiDgdALLCTmeyIOQM56iT4g+sYBU6KYob+zDfgzZvZVVsOmfbYL
ZeaGRWDa/d3KfetyTCmo1XOlLxwzrwuv4z/B51uA0TKxeyDafN3rUTxTtm+zqm9N
p77w3EmYafDObpeRasNrSZlMxTNII7/8SQbrZqvvnGVq6SuVLEJ1aq4xUM5iadZy
hhtU2zV9p4Xjm1o3SVIjdVNqth7eHvxZ/cETH5nHsA96WfHWRMPW5LMMzDYmvyU7
y9t8WsdP3A7AkTGkjQ+rQ+y5IFg/TVnruUz6fGBarBHr2rBz3hIIWfga0fV8Cm3Z
VWCR5/as2f9X36xbkSqZMLmANwe7JDHBRC/6IleQsPsns7+M6+PZbncQlHSx7MvX
U3WXS1UkSbIA6vwvuJ7keCEG3ab9PrQZQ8PB9a4prLrncgt9Dl1E+2GzzJw4hYJK
QtKI+GdW9afMPcxPcHJgIkIMl5o0xwVz4VEy2vc0YjXTsfY64vAtTNG31mIWZgwu
i9X7aMi1rRCNOsJSg2uaa/IsS5OnvZeSUgO/FZRIzLvRxQJTFZPnNNgpiUZYd+oH
7clT3/eGZR3yHC97GMuWICBrwHYCpixddowRNk5jAB+lPawijfYw6oodXCZCT3ZP
RENAEw85u6w2h0sBACKZQgntqYV56aLDV9q3ATh4yeDIgq1DqDTRq+/qM6v10z8q
OHG5fYegC+kTh7BFl59nT2sGSJtWwJUq+SRGW91yx6JT2/k2DC6g1ucJTbAJa+iG
9gMOc+yS/P9ST5RM1ZpyipySt6Ne3H+iG8g+0qsQkHpie/iQSsGbV5Xnw/SBEPU/
kcClhtihgGM80m41EOPbX2AF+X2JHw9uboTd//xgtGo/gVhisZuUSnKau4tVYlIJ
eNPXopHFNyDSdjSijceZArV302WLrl0HWoqri1qqLbAYEQgLhVV83xtXxCE/MKzg
GGjppNNPPWp/rsPEW97cCJWCSLiGXWq8AESS3ZKlg0qwvDsEvHRbTEWxym5DlqYS
LsdmZ0ZLnOHjKlPF7/m+coOE0d1zo5SrM4MkGgybSriHxH9JXcjiLEjEp/10R5pN
9hFaYJo654HB2tQjKuAmFStjTzSi/CGk15N/fES9OdFiZKSSfWXvlrUQOZIiccy1
rUXsWnV+I8u9gb4ZedoEs/B5w+n+hQwuOrAe4mkdBFp+adELoXP8xs3CIBueOBCe
SgeRS74x1xmA1ph4CcwxWtZlOEiIbXWPPMhomKSQ5rgb/vTDysSZ01H9GMlosO8N
IL2K4wcIS7hC2UZ9+ZYCfQnXX47sN514712z65AXRNs8ElGh8LO3AFulaVdvDKrB
1AVncHYQbe/7F9DOOQoWc5J3jAIy/keKk1wtCTXJVNsZF86b2YVXnuIMDJQJyOMn
OB52MySvBnFi9Ne/MEzVWRHouXzhH/8eT+HxdDjaLaKPPaHbkBtP/WQ7FpA4aHqg
5InwiAoqjDdvJPsVi3EQzOJIVEQGerX2cIfa5I62XcByGijyovOvSXWgWLEyPyJO
MQ0ifLS3kVj4yZY7XE/HcxfXUK5qtVwm8nGAyQ1kaydjKKvxCPAjOuK5bgAkEdii
0tw+upKTpgghTuJDEI1Dtq16qHxbr5QXMm4gAq9izcdl7vM7Les3ddznUYTm9zgf
mqB70d6VDb1osKKRzON/GuGzCuOAqu66It4HlW/fdA64IIOUHuaso1GLAYu+mesy
DdbpC1PWPLcFzJSiqPKowPqrYHWDUTYlAbY9zopVo29QTpR1wdVIicYY3aHaSZii
0Y872rO9+mpzCF5fbZYf7h0Ry40gb1mby3hB9AZJjZL1PbGjm1Xa96YhWc6kqhJX
QI+Q9is4bgHOFI+89Uk70sLNLNZUp8m3gxXKSXFG74iUTp7U9wi3DiI5W241fKXH
57dN1GaAfkSPr4MW/hTwwcPwIIyGbHC3tQit+hp/EOGFM+5lwlq8wJ6pNCCM8ux4
iJNRBHShyk97x2FDZ6ymYRXqDxx91hHvDSRrFjtMaoEi6osEW2x0Iomrzgy2rZ9u
jJOa76siCYwMTsPQgng6zQVaC/cL10GqTKVDIZ5lG78L6ehOozO+joiTsuNKivmw
qOs8SkYcd38IyKQpUrNqRF4gsyYCHuEeQXahHLUjSrmB4ncjD+KnweZMZpaE1ItG
ofAw7GXi1yQOFIVtJ4cYajYRr04x1pacCj2Pg8qZC3slawUFafaB3FeC5CQJdbjv
qKHRE0wTRnxTL5EvR+6dvpO70+YOE0ojZOgfFCBpPSI8wxfsKVyCI9BgumawPySq
UaSCi7m4IJLHtnc4wfKhUBrVVcqSJ451si5Azkoag/z3dvXc5fON89LCHRNgQe9b
HDn0d8q/a5JUsQnNBsEJLT9BVm9OgD8faOA7oj8CkAQkdVxuOPLjUMEnqe1pkFV3
oe810QTVGg7rT2FuSiPWhO1swEExfyIZ/jqRdNdujED6MAkuAbKGuPjgUi9lxzI7
hSXSQZMJVpbhU/2QEDHfnv7aTFImdTmq8k0SLd349tOaKpPZ7z9ayMho5QIkIo6n
8/YNofHyPGTzwzbDGezvbiVlBFs2lpl5vh5YliY61chsX8F3OCWFxCAG4cgVOWY6
mITByePuVP5DROczDTT7Ya3me9b2QdVkGCG6JD6H+z35RMOZ4o0f2bPz5pYisw8x
CM62gjJHiYuyMxoFNCBvLzLMeMMzKgA6RgMD4YszDwHO5mu1kwXi522CxH2wo9B5
UrNw5U9amB/+OfKWF1Ff+NsHRLJ5EcFreCLCT5k2j7pODWELoNx3ZZv921+s//7u
xAMDbrDZsKQF7XKAUYEwOXe8HvMmjfQ8UjIkinzqig45ZoY94s52tbu3tRbKdPQ8
udqad2cObluwTaXDdZHUc6SrsyP6/Ztr0uDYowHXzC4JS72Mw6+SnDE8WbZ2hA2K
PTGjO2HYOIYCb1RXc9mrcy3wrUhr/g+tqawDH4wdh80MateTWZTXxZFObFvwaFen
B0JCut4NzW9D+1xcBxzlGkVAHkAvTRACxth9nLq4pr4WscS0q0/1AHMtWtM3jMIc
AuMtXCOpVpepf0Y9kpCSpQNDGNl+Pn/XlE7/s2xdmuirrvPwxhMw/284hrLYKkF4
iyp2IRIwPCdd88OpuFLUw+6B66IlyWFt6bUp7pExlpp1/IhkN6lwcODLA44Yoyq1
JqKNX4VrHWUwzGQneWpcXg5IaPp2FKYf5484b6N++2FN8TdXSkQOKF4YWk8jMR5l
Z+pgc54SYHq24iZATDJZF3/2LEdsw9+12HAzH2jlmzLUUkkFiTNReiYWqDsyC2vZ
gng7nJYR1Z+xyNOS7OyI1kZxJiqmDZNXl4MW3v0vSyCx1f904lxkT0GkgO6GNsNp
ACpey6YXgB0xOrQTASjz21STz7vEA+Em8NjbUAuuiQe3w41Rm0+6zj+hTi9qIYyu
s33+NwqArBCK2/apjMMC1BjLmxgn1HYJ5wMIma3issS6uwNcMF007sK8kAQMukvS
4GgeGka7eFBnsDclO4HfY9dl9C4Wi4VgNKzh3OSXZ2/CAPZtJIXcY8oLCTxRtHpm
R6SS9zL0/Q7chX8rq0CxsjJqsVqko64ECxscveIIpW/Z9ifhcneaiYPxSbqRkblu
CT2oVIQCDbGxMXOy4UzSC0Xp3RzIyD5fc7X8dAi+wK+wu/vdcXyVY0XLo6yrPEEF
Owb1xU1np/I6p+ZyIfrC6mtDBxs5iKvNCUCe0o5fQkKcuI+kFoPFN7qnqk6+4M/P
btNc92oX2PI3CjbJhpwrVDU9j+zLhLI8j1XT6WgXnH/AqLJDZRJOT6DF/WRAdEtd
upJIj8+uNQ9VwtvmkCO4+uYBpM1FnAFxYOdymExtfe6JR6qxQ/bVa//vagujWSIS
yEKvYVMxNVjvtJllXf5OpLe2qdOYi2iffE692D9zgIhEv1ADlBj4Jj+8kNKFKphj
NlMV2eaVBttEtSMTdiWYHtmPYUEPsSOtkEyeoa4cMNFbEeOWU0sDz/vXTQNNIfF3
bdr09lScxTIPm8k6FjDsKExwCY3reJP7O2gQdJ8C5SdC03uuW2jQqcBuv7Zm3sfJ
dRvatiDBCAVfQEQB47QcdQSdI0Rnqtqo/5cfcoo/gN8xaTV31YbytYxQMAPNmuFc
Qdgt1uBzSddlxkrRstS+sIoteBSI8LPPjX9KyyMa95zBaMGpdg2QR/MFqM033qIC
yCRkXMbUjFws4ZaUTzE1xJZds11ZMfnzt4P10iW02KDCrYn6oqr+rNQYVCIvN+vI
CPQq7VmHVWpwPJE5llS8cU2QgwQFE7/HdfjfcI2TUq2oWF16BFeIKIKrMrXSfadQ
Fcl//cneUtUO7ZWZdGsKO9NQasQp1WpoteH+sDQYoBs0VMPEOLr/2bPb5qQiAJBI
6G2ZxgkAWSVaQfpYapSIdX1snzp75+IYpDubJDRb49VkXk1ojZVUgucmz+GqozG3
7eZjbSkm3eH/YQ9fqUYCyk2as+Rk4mp8cxPH4pgJF5cAQvELgRB/J4cMdAsVCZZ2
Vb23XCX9wLPjUdeOVHR3LrjCe6KbBme12W/ds+wP1MSaxRTkuUzrAyU1rM2hXy0W
ZoWzwhvrMFL9T0eMz16pCSNxDeLXAN29rqnBF+jatGI8XV6swDH9W3eLhdb9pXYn
YHBBvovatavhZIno5uYy7wZHnd6kRtoFQVHw4yVlwAf2+2gFUEAaUUPMFYYEC/Z6
e70fSeA4PCpgzGT8UvK3TYu44W6g4UaJGBgmCsK29qKHBxq7fjgNYnFGKkFo1mY9
RW+9UdYeJlixGXRHxMyYR4SNADM8+fNKB8Pubi+VuhXjALtGL13DiRlXqo4a3Nao
x/5aAAmmotfN6icy7RrOS7JZ1TaqKJJE703FIhXKRzpY0G2+ji8WAoxE/JR+wuQA
BWoZCVFURvxxGAgDZVbT3c0r4byx06cbK85ytx0BXt/D2LCpQCZcw5rhCb1bWzM1
sUGHh7DmrnAhZe4K+rQoYNrO5kodT673gWwmFyimr5EMKPjyV51IlUitgDIgXF2z
8gHbDiksWemDULvvt/6Z8XcdVQz2c21AA6CJRHP959+xNqZ8b5K74t65Pj1djxkN
0pjw7FV75VgoXLumY0AryAe/Z5IYrpkfGw5hw9jgrkS56lIggII9LugfPzVTUXe1
/x36GnihrdfV6hSH61KILLJe90vioVNUzxe3Z+JhrLfGcQ0pLs/3HymkCPP9+Dd3
y1G14XB1wasPlwMqxGLouns/LB0roAqZ4gBwPX5Skahkgxivcbv0KSge5RAVjzGd
8LxVP16/bHEPEJ3XCLoFqR/o/e5HUdX+7Mo0iFOe71b0n9ZOw/Fe8dAU6bDUKCwB
Ql/tVB+Rr2wR/N188khP3A3Q+tQnxtAYoSWFnQO1t5Nda9FkFqD/8mdNVOQP/iOD
jUdAGw4JGFIcB5JAdb8STOmWcQUbpexInCY7Ahb6B+5vDVEEhooWM0wl1cRbEmU5
ebrrw/XQ+eRnGM8y5rGhVsP0jreeR4+GWcXBEi00hizT70hiQFquCStwKVvKc/oE
BL901kejHMbEmtQUVm6qK1WWXFV18dksMEzM6sqPc01F3tU89RCZCf/I/FcZfOU6
/7VOGiuAiK4rFQPIuScKyToEMyx3l1jUFlfVZPtsT+inYSHcY6xRypORP7B/hOlp
01hDr7+tLwScKbjP2TS81+UQXyt8QSHkyGBcuVvFghqynL3HfO+HGNFbQ28pjHvh
BdIfQ8zYN9nQS0SspBnYjYAUe1IXdwAxHTZb2fhWoLzguzCwi/IJ+SI1lIp0ssNB
tbAE6yQfZVQiZxMGQDV4YUfe9ZZMXJOvPGLek/anI+Yw+dthW41bMJpEHcswVhTK
dkcRuG1E0mibTttDHLNOzxosApsx1CvI98Qnl87HTJLbrjm9yCc9O7Q9Gl/i6OE/
vYQbUboQiU9ab/l9fDFiineCVK7sLB1cwIAEeC4dl+SspQHiCtBR2SJxQHHFWW5F
nlxCwzglKhMdB/PfkD3tE/eEz6yv+SqRx6Et6GnKcKgA4n0ZdPqhfEPafs2pG+3C
kbg/ZCrOi4S4U/Pz9j1VdFTfDSSNbi1lIQgBdW6mlVuPmbK6m4POnToy7eVFdN8c
x6GTD30pyEJxnsgS8w3F6rZYI9G8qKOHRY3U/6yf/gqp5iockXMLsJTJSeEGihBM
p6/VmW3iVm63S8UbjMF5dLj0yf5cne+J917DLANMa6dLMS+t6zhFbdVmC5CC8R+K
jfHyejKFAR287kf5DsgR+t3MB0ZGIBVxkbspMIskQtjt+DInwmtEUvrj00wHoa/o
dudeg6tEnszxMm6MocqCn2WA9eMlEa1m0R3V1wcg97CzQsP+WmsyQcewmm+f1jMD
Z8M0k8nL/VcOO64itq7Ou0Zy8ma10A51Vi+jh/khoLlZ5DviZ5zYDxz66SJyzBXm
k96EC5G/Fp6YYfXN9kno6llI5WT++51mjOw/hgYVw1IKL0oeLXXZ985PUg8EhaaA
I9TrgjlCiDaiLmmQtwwcCtIwJfpKEr8SeAS+Fwv8xizVoxx8BicCLZ6zYfn6CPgN
cboV5Va6G9XDEjA06bpr5EMo6V+fUBtt/rnouiAPf8hCoDxyuMJm0QowAlEBU21v
QixQPP6iiBg+8AHHF0G0dMFEJaOOgJ0Y7Y/KrANyApwL18NlAM0yFXvn/qOxKbM3
jmfMjgJCnESTFc6NzDj7OXB9dZJUEa0kiF9nZXi+REfXM52h90Be7GODGpTAIQBc
VM8HGpF9jehWk6D8aoEZO7wfhzJSPRJguxNZAhrtSnOJzhXQuJXctGZuUNLGobQb
80Psf6UVSwAWi4F0b5gUWxdDlIwRDzaJ29tiSURutUm/A+sYMNJ8z+lCvizx+XD1
UoGlPglWI4WX1U6ZNg+2NVQRpd2hMGPL8HPHFiScepNTM4YjkcfnWeNn0cUQCn1L
iTCbEFP4ve6SCb6W2XbirZwyXkHT0LUBxrRx1WHQhkJYyqlZTQ4SdgX6HsK5tR/K
I9bqaw0Bm2r82Pn2DezjRynXaRhlHv4NGspubs5kq0ZUGcryLabhaVcjexZeJjPa
dotSe9nfaV1UQ4yJ08WUtcWCJSyPam2RouWfApl96yYXNxnP9q8H/6MJU/C9QBRe
449MV5C7WtHdI02dxh+Mo3Dxmngrr19UK+ewGvCHSlu/aabiAvtv6f6hm6VNMnZ/
h9n2bBXw+02EuJZD3bj9wgTzbwc+wQOUqgqREZfj6Tx+cfb1wZJ1Q20+xuRQJ0Ww
aPrcetJahUwyzvSKDgAcqdGJ0VozmHjJwy0vdb5Z0WqjJaNCaylGE+Qi7ik6R7cV
Mth0ObCeSM6Z+3NEjMCFByjhHQ3YiD2ffsmRrxXQ3utXYybirNyGXo5b0SOCvqvw
I6aHVFE6JZ2+BJy2K3vcbYdku1eS/K7WVJaYwHCiD8yG/rDeuQAKeecoxx1pXMv/
TvJv22wLlLYs2I51xP91Rs3AUqWlcUlPIBZaJiItaQWmyjxIoZcJNyw2nGOANlOA
uT6N5M/R+EGHxQ+TOiJWd5w1OzJ5WgVyBQZx2HM+776eKuX0AM5SFB0rC2YkXtdx
TCPa8u0XCw0rDGQHymDuogdf0aUWTYCBWuVwHR9REntJMywBUQ1RddKwqbd99GAX
/mCD+0C68pqL3V3bUSS99aMn1icoPWSZhO5br7c/SngRGmc9dCQfHN0rUls8/cXC
5F+T+hD+rb/e6gGVtPRmEp9f+NA/tN6HUocdDz7Zi2vBkdpN/UMucwwyH5mpB4rV
WIAjGouVBgartcAN2aQTHdhMvxhBzU1bvdWc+CoCIralBWV0u6uu4hXxusc8VeGJ
7RQqLrZ/hn4TlErm1qzgwxawh/YwRyYybZ8f6FMF9e52+Z3yYw6g5WAv8zOcFt5N
ykRSovq2dStTl5oGU90zyAOtIV5iCJvH/Ip342SndgUlrYJ1zz1ZZBghI91nV+Ga
gQUedgAeNM3UtMkxIHRRdzAc4yTz1Wce20hKaWIhgyo3MvI1I4eetIauFLDAea/e
e/TYDJ8P9YJAP8TQd8AW1tqhO7CBV9dYIzHHCxzTSCuM2tp+UnbktsPvngKl6lhm
WXkP7hhtBuVQgHFTqks3xA==
`pragma protect end_protected
