// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:47 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eDxFEBgM3diTIkftm56vGvvF0WmHG6u1SbzSfjkRUvgHIHfm65EYKN3hMRD7mvua
+Ynwk4udu6fwX6p189KjvFuly7SDPqhjvcGIEBxvHG7fx0CmOcuf4qV32W4xWbiQ
+pG5nG8BuHXB/BaO8ToaLrpZ+eGmm7Jjt0FbNItAMgA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4112)
VHqZhM/vxUtMrtNtvNnk8eg9hpcFXylho5qd1HvkGPPDX+4MR0G1I+U8SC+YCnOi
zHeHKf23YOdacUKKTUZO0sKLg5a2zOo82QkhlFmglThl/gN76ptgbKo5N9SLrYy9
PF9dfGjzfUHEhCKUnQ5he9vrN3kvf5B8yey8+XRqPw4sAthJ7Jw4rhd6z/kcvrNp
VPGvcImPwISo4zNyL8u/IbZk5FhkzhBa/QrvEARFm6mAgw9R8oEZ41AzkcKekKwR
4ezgXdFAaOBpujqFo8pmtzKxg54bVCFfWMap8WCA9Rh86C1gcg/JDeZPb0mhSJJN
qFW73AjeKHpj5BoCgtYtxHQ0QFy2HRa4sYLQw/uATDNkIJjM7FK1dSSSSOWS8kdA
n3j6+imxrdTgjOBwZX/nEFiBZ52RbA6uDCzwz1d3SFnZ81Tux9MM3w6P/BPe6UEQ
KJskVC9AKIsqP4RYU5TC3OamXj476wrXdGZSgaQVg6NoDAQuyabcdgSAyHKM5Aze
gTWYepEwOzgY1G+qyOSzrML8nJWik+e7MWuE1TsNp28W4Hyn1EtkZH4JlJdMDyRG
Qb3ah8rWB006dkbffZKS9nht1a3QBK7QTG35yXfK7uARzz0FRuBCWl7np8LJLXRk
w6sU+jKvus5XnV5qnXH/zhuJil8+zsy21vJn0VcgedAk9nsUg3JECRWWGGl3YdSC
MmNLO1/uSz28TH0uVupIY7O2TFc6HdfnwdIV6kpbi0OM9xIDHzznlKIve43abpT5
8lBLCuufu+33uHt4zMxEfQG9xjIOvG8RsK0vLvtIRBE1huTLwdLx3CRAtxAARx9q
yDcVmOX/+V8Jubyqp/zvP9HWyL7gt9Utwb5/KWWxdXHbDq4ytnS9hS5tm5vjm1eg
aMTGFI4hXAFAjm1jvO+gnPRS4q8UKpQqtNb9e7UThymLZoa4Ketgz8uIOlysNgM3
sl6+o4HU97HomqmCOVHntp3lFfC8KfxNpsHYGZRtWZbN23eQ7J/+gQuK2UEUcoiR
UuZ4aSYYp7tdQE8jdqaSuBKYsuUnzl96YNMug6zZBjpv6TJp+7y2tCnJ5xYX2RES
kZPoZBI6MT1eZfo11ua9UlrKYOzeQFLlnEeKiIhZ3gFFKRMjumYJ/1kikjWdQZha
hUZRVuFmEc2+I/J9g8cp09W/u3opN4ZTNa1A2jtkNB9YTTfhfkqzdDmMz0HyNQV0
0cnrNgD6aQcIWM5K6na7W9E/+OWAIMfBvxA5NGidrzroPkECy/x3Na/ILTBBrjLi
pqt0kXyUCceHb6MuOs1r1JO9MMtRMCTuN5iko3b+wMvCWc/agHoa4DiMMSKr/XJ2
kKDQjc49JukfltMKCy+NLQxKwOZaj4fhm+wErFeF1Ry/cyoTp86Sj9qmJN9KoHui
3ac1Sg3u19OXPnotEfKQPb0skKNjpiVRicspmTZ3EY1BCmL1Tk0NU4vQU6pIBV0e
zQsZcGZyH7NGGNQjb6vWYJamHXTloTdc64cCRYt43s1tT8MrZyKA/YFKdozZ5zXc
gqVGZ7VE2WQcPud8WuJ4akCZNTM5HUVUOIUzWFxYGEwHsK1WpApI6eR6cbpPmuZS
hcYXLv8+qXsqG+nRE8WCmRSmk8LiN17HufedSFF8RsyXvUlTF8nsQutxz01EA8PX
+CJaxEyXhC3KUuRYsF5u++UvaR2fwOKwqqN3+y0ze1zec1ph4/rVgOy8R2fSO1oL
+mvbOXp+9QjVb/qNWKdJlpLzo+r+SydJFU3gAHDE68SPuz6mC68fvwIQ6QWUa0xR
hF7oYVtCiikMNtcd2pNaH43wHivpVP9p12wtSiJugBCD6j7PlZ0mrn8HT0uIPmwr
xpOK7YSqu7XtOtuty07B3FdClqmzPGk+WYJcx1nwGfZmYuPW/ASzEbbwfuimyRVn
m4lMeqMOUwiB3tUefGsxcsU5P5+oNcLIkdKz9jtRb6ia7Qak2fpjPiWLP8G3YknX
EofuLyw5R+T+4zM5Bi3Il3RcRzjJnqBGtxcv9M7XoYvh5SknymMuz5YBHLP3wlkB
ZGxpIAavfxGd9wYkBNJiJ2WNiKqJHH7kZel0drN+rZ9XibPUXunEtUvsQ5vjaEXx
7idLP4y/vqzJlDBCWBYeADDMRNXCKYI/JyEH5XnpDleQqhPPFMWC2HZZkYwpgKv6
c5Q42RIniOpuk6zIalgx93NtwQZFuAzI4n0txeGyB3TEoOZ85JMTXpLR8ZHz+/7u
rH/FZSXR/VZ15N/sn/C7lw7+t/QQ9s9lcsHBlluTSkxQSrjUG1PdEfWPjBPEtT18
ZjwRZVKjJ9eQzS9fhnXDU/ohFYJZgSdXzy/UGZFspxOlDqaQt8CHAem3vxkbR1Yq
WZxU4RZ8bQx33ntw5t76HcEUNQMtOIBt2gW/mCvAB2tNuV3hbINLQXLJ8+wB34TX
i3ZXSHuOCBJb7jknZOXr8/NiWcrI0b0GF8b3JXIhd0J4Or28EmEvNVKVqyJieNm6
Eqt3yxwHAguwSMzN5whm/FFFfvBHL8/b/Bcg9Inv9Y0TCQCsiJLT6JzY1PnGGJC5
CSQJnitT1+y5/Q2dbCMqsiquwgiOl1OEw5Twfa0vmd1GHACk0VSy31M2tL/dky6R
Ri5OtehMKaZp4UapJNhRdz46UGgIaYlefsfUCsAdBkEefIrDHc0OO2OiTZcM0tQz
EgNNDm8lqi19uJQzQZeupKmsor+fkQHsJnYz5jN+MOCh3IvlsGDtIYyBbMtjTOE1
q2qnZKag31rs1RE32Sj+3OVAciD6os6MK7p0QvjvoaPEo/Wv23DuIQlo/YQAeonV
JXZoI4iyw3WRz3IEmJmIQqGbyu3YXJbcBFdtT/gfntmsQzvNeph9lBwsk8/JDtQd
GEBGZibd1TJOvJbPLfzilKoTH8Mi5o6W7GUgyQBXji03e60086rbklL4nNW+vLuX
4XqxxrKvVUAGoYFrahLxbw+Zu2c6CYtQ94XwltmurCih9aDEVTBARvmyFT3nBkAt
Cn3060qA5W5iOmCBfcX/VgVpWqJUaW7rJwo5cyx6dcWyjauPpWqVgAuznbUaeOjt
wZsJRStpeevtvLiHSjsqCFaKmtN6d6Otyx+k3b2crtvVD0SeDKJEX5bQsgVqHob+
al1GNqtJaE+6XRyJZPmIapRho0VzAtMAkikBtrAb6nLIp0A1HTEuytdTKo1Gg7eR
YBwomiAl1zTNLBc9eRomlo/+XV0dyRKFAP4XmuezydTFDn7Fvd84ssb1xX5TO/NW
Lnaz2pjI9Rikgz8n9zygl6tlRGFXfO6iRQDrB/92HHlu2oDd+ioG5eCvahv9ZV38
p5lBzcPODUHOSGoNA/ZPQBHBb8ZhpwUb0QrOtTRDYHSyJu7pmL5yR8lTe42r5xmI
Cy6nPgkWg6vt7zv4DOLbhE9LRwOCOq3cDZEaynz19bVtSKGMXphqD2oJVt82lUPn
KFRpVfqXIRT2vf7oepzUdpwdyaxZCGsyWPMjWVn0LfAwv2BuW6hxKQKezEB4cy/v
ftMMnEdP5T8VRE0NL05Ap8Q4EW8TjFGxmruySwPukPazid0/NudY3XHRhuGPnwf9
PepW9uwFQKbd03KJs2t3LqFav5/GQcDh2J1ZEL5XMMZbcVb5SbM1NuxxWqLbqxAH
D7GltGWk9BBSAyHDII+9B2cXioeV4/Za/j2aWL0BAhAxOGybUkVc1Vur2GdI8woG
Kzt2V+lKfYcBQaCr2EhJV3cqV0xv1E3UINw6QUPvKljCMnH0QwGasGdkYs5QFQe+
vytJBTXlOT7dKhP2fgSwcI+aAdiSOr90HGf5Lrf+6ReshCSELPkNJPYLqa3S+CRe
aSJ7Yh1r0qggj3xEmU8lqg0WrXEpABXKQ+JKP5g7zO9+otopZgGj+mrHHJDdJuy5
FsvNkdIS0kODQgvmp08nT1pHhTsFkCkqQ+LRR/rpLpOT0xcf37/MPxAyAzNivTX5
eLzcJ3LSgAODrQ9OU68Y0GlIIIhl/FqQrqk7KlRsQjMxLLxnESTxTF0QYp290mo1
a6bnWWoSXBURsC3LpCwsfAjz9HobT5uoALCzQVfN9+wynUESuMp1/EaSYxl27jh7
FqWEYMHGHos3M2y7B7X4f8D2yR9L4cGcUamXuYnDHAiMqJGMMiuKIOIdlpeI0GlL
Oj2Hfb4QZMg9Tat+nBC7xGlUybs+h0EMEnqR+DRnzybh0TUBqP7grIv83PZSpJ5v
PZ2dPGKlLWnkqEh9ADo8op3qXEuV/W9YV16i4zv0KVw/IgAUifR2DZZEU6mUyFlg
3J+WC3A/MCleVgD6t0qsZfFP0Mpl4O6NFk+E178V7nUKoZW4jR2vqGxEIlRbpXHo
pmmasPVRDaqrZJsjT3/6wjU7L/TuWMEazuNFuMUkOv5RLHPFE6H+7WVTvlb1DjxK
ez0ndCB+vuX+9SxzfJDjZk0azz2ko7xZ6maT01dRI/7hZ2Y22aznD2F0NJ02lrw7
/sXsRV3K1h/yLkqVBscIf4L0lKiIA0wDAxszCESDTxlCxqZQkA9qqSFZZ54yQzoK
d83Cgjt+1KlPBrACqnNvmdaJ89mOMxZ+AsWxkxa6Ez68EXmY6zt/dk27MhPwDKx9
9q+vnkOALo2rCWtTHznmoYMRU87fkigyz8GC1FqTjX2AJgbHxrqvGdfTsLxw4paf
YNu6tbs6sWlJ7zun4Z5MVZv/plBuex6DHy3AEBImPjv40hZfaBZbDRRADmZW8nKt
qGaOFUfRyiLcl5TLCW96PDB+9rBrEp8buaYLGFnlUqZTHDBhA8ejiue1V3DMeo4X
akmGREfUyyRlRu5853oeiqnlElH663okylWMsC4TzL3UeE3wISxZOZxMhwNsMNT1
ZVSPffUDXRt7OGGihJiJ9p603nmSo/3oFie1Cwr8OKnpPC2LdoGBiT9yuwlcLxO1
i3PNGw9sF2Eq/Qbc+6Iq0MFniBF2AFzhajeFUnBqNpusM9y5vcIXQgDN+GAU6jdB
2AJ0qk2f8JPtj1KT8U0PHq1ZfNO5/c1/qtOI9JHx13XKCCGwPVNxalkc3njXa+et
QQWe0cneRcXvvee3OJ9omN/++zUvVTJFkOMHyG9vOK4NBdh/R4KGUfvHWQzUX3vY
fvCY61bB8cSi30/cRN+j6zMmCGBGubub3bVDv0wez/fZVyFCK8qIENpFzpFKwGRg
UQE55YfM3sRBJHYV+29P8Kt7EeMOtxxB7uVs04gS51E7blvBhCvzVo2m+iLwsXWG
dwoQblw+rhi3+rlwwnhRG4UZS4nkvzJKEkqAflNr+TVIjMQCrebgYtAq+xq5XVa1
hXxV+fJZwysrvqiFuIOdGFcUT25fAgqNcMAsPQTL8qSO/zHQcErdczQqw0HAK2pk
8tsqy61pua8wW0x7X3ls6KJlubNO/EIa5xXvdWsxwTYQVQEEtSWM/dObSzYEtciI
Up5+3akcZ1Xq2MgHy1dNIcQ+nHyAzCPbOOU90TDbn0I=
`pragma protect end_protected
