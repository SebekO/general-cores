
module single_region (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
