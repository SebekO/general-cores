// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XPb3gRPNR+x5OP2Y/ISVwHvLNC0Sy63jQm7gL8mhz1LUuMa8hbLG/DtrE3ab3RIf
Bdxbx5SSv/WaOETMuGeVEmQ9ZTZUGVKx6AShrcxVDZA8XX9v4VWNfHVGH+UCXejM
ODGXeOoO9INxaioFAKD0mGgVSwWT3iUKBbfTVeurlOA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809904)
dMKl9tbbapv5DVDtUylYA4N56k1Yg9vmknWeRjI4deDdrNtk7uEKuwxa0ZDrLli6
gs5+5cWt9JkXNK9DUinOqzKKUwqe6JIKZ2t5kM1FXIfoTn/5bU2m9m4tIq+JW67F
oejKfv3JJtcAc/T7SSyI6ycX7WCc9AdNMY5wGzY/sUadCc+jGkaIbgn6myzczS1Y
/jkS/oDdongeglAi0D73HPskxinWdK9BxZDhLFBbhHJVOvlWlQmqutj4Jhaq85KK
Uj/HzGFRt7V9y0JEwdrvx3jUL645cMZisioJFDRFDZlaqWfgO2RV1uwxqtYaRWj0
VGsgg0vcOFxvKVFlWNOm/yB6XqSPIflC1/05E5phEoRctuVudlT1DTdryzISGdPi
5XHjb8Zn+Y5rtQcd3haoEzRVHro67YI+vDergl6YvVuE3H6ciHuH6lSjc1mEY/iD
OQg1BRM0CUuBjBXzdNX2DyCiSz4m/iQbcBr3ra7gbAb3uDbZXFjDAxYaYDLzx3A+
HFJeK3IyoE5YKvUcdymjZt5BonZ2jI0/uWZzyB8Pcyv1qgfIE0IWUjBmagluTGSe
rZrwp7jJ61KkZXzRHnua4DvZF1vjpYKpay2HL5dDQjE07+D2dwwnFkyet21dnopJ
utgk/jlSEOY2/oolbUaCOI1qzhAQEyUpfGZ5vOx4I0PuxrFyNTM4S7uE9YCjMTYR
8zx6s1/A9HpSuUnq7vmPz7YM9bSxQb9fBoxfyrFJ7HA56aXb+1YbqRcf/kOuhTTi
AaPaliAEap4h8+S4LfRdHHP2ZBjG3qOeY9JXW8tIMkd40VlI+TcA7/ODbE/xdrfn
yYcLNdSsuGarNCW8FtuHDsKxfjOQkGkLClQp8xqgh7jOWWI3osNAj9J6Yurhaa1R
yvfYHSQnmn1bpCgW58p619sn2vRkqsZsQZEdM5QbHRsA9XGy9mJsUqj6SFOEKrMc
aBUXT3zvytS8W8/7fxGtzEPJw9POvZrOmpDg1Jt97GHjMMQhpXtVqm6Shq26Gyzn
Y+W6J1wk8TcI9qVHxWCvolmUOxLWrLQma1LaK7iVxBvUtYRIf2wnSeyfF9F6zbhk
W8Pfz0+il6DYC+kNNxMpi1QEtY1EARv/cN59s/DcW0k9vvo9pfpbOZaoGSx7Kpax
w4k/OTlqOWgLovdDt0s9yp/9SMRzR/rmFKNG1FuAulG4AAe+w4QkbfzmF84EEcWm
XDPDhCL9bzE4VjKxs6uX+0hA8y1rKyuZq28x6M5XppaNcmFjfoZPVu1FRPNc9chg
efUaJ2FXAIyNpa4b11Wt6AHFn8t4PYa9VCS4RVmyNOWB0N8MBpXruLj3TPAG7zHb
4Qh/rTBNWK5GIp19RvBmwj87nKr9uBEajhfZdNXr9D2Ge//D6EEMj3/5ZXzNWD+W
DlSi0lOIw0IhOBJYd5PFeIpLYFI7Wnk3r8ycflHOmUc7C/gaF/fDaHMbCC4LtXis
LhNjCjhduRgVbUnq0PP2Tyd7FsZHLNnnAnsPB3X0euSyFEGrOP/l8IrJlArjEpld
rE+XuHdtPemBLIYb+Bb2JSpISz6LcLnh5q6TpH2K1zGphK37lliUWwuvmSk5cSs/
gZKAsfxGzXfYsUb1G7GB6PG1foYqZ2PidYB9AY5jLiK9mLS0EaqXVSetF4+Bh6va
ANR4MdM8P8PreYAaFMPqV16KgiNcYHJWl3nKEFskF5Y/xgMQpXaHV8AwBxNVFgdy
PMxCr/kE7beBnNE/uogkjVIpX4FToXXXu30VffV9v9l0p6bHx5mgd/nrLSTahaFr
wG6MjoGH2CqwKsaTY3UvO1ROoNJHSkUBveT0LdHxG2Ue6nW3MF/Zr9MaPDqGYZ8X
EUJYsdLOcMaPNq8IBVfm55u4rNDOFUaAi0c8FDmrFH968fE0IOLfKnH4fHQSixFU
0zZXQgGZO0eECEWfcrTOmy/Yr33oYyPBhXzjEt/y1BAfHWFOGmwmbxlqCc6KSl2X
IsNc8BC7w3Zk024k/KWNpQUzx1FeJb8lIkrDS4KFW9EvfTmXWzVG/IV+6oDQKRt/
PBfnIBqfXcWGFKhSbt3CbJLpfm7vC8/6KwaR8vJgDfGbuFt5uUeYN1bF7e8gxnss
+qlzckmLvugkJaTt2PCdrL1z9sUIXFIZy6C/rn6fOL/u3hrtDRpxaug4cInRc4vf
oFBJTPZVWVJ4wOemiZNVR3cKy+BVltNXhu7X1TMZnD9dwls1xGahXaSXhSmD5Fl4
+OuDfYHwbQVVYyP/E2i3xYB1Q5OC3czGng0r9iw+LrqlsLMJ/nAxf5HyhEAXkdJv
8cccNohDE2EFtl0MBspsd1Hn8xTMzEySGyskLXv0mTrkcShEiXtW+Teiw0X/L4Ln
wjzPoT25qu8RXiHWYVptGjhQrM/hPKwFX0e1Y9uaagRN2fjAt0SVNFzto8IMbvH+
0XmCI/3o6KVVu2AP4P7ezSiOEXkeUJ8eT8BMow0SkQhLuQ0Yu1Auw/kT/AzY4r7G
kBVEcs5n0H46iBPnhdPMV1f3cJ3JiO8+x3y1WZje18n/f/1hYZ7xj1odVKvAZQgd
3eyxsJnwAQANUMo/SaCi/e/I7/JbnemNe2gDspeFv/VRfSw3u29BKC7Asiw43AHJ
jXWa9Lq0P0ruv9RJDEq94oj50lKH2KYg+ufHfPwPSZ+lm8E2yhWJ0frMzoCt3I6m
WtX6SNGdb51OaENwlCHVlkxN4xLbepbp6+lj7bZ2Tsy545R/wWVcC9st0GpWmOsA
We2EYApE/qcKuPubYm2NVlL4GGx+7NqTZSZKuIS95tjyHuWedjtb2JJEG96XL6al
HlD0XuVQ+l0kDNyUPmSDysfCKLbwSD47o0VqaWwR94oTwnQKroYkdayhArzFxiRL
Q5sVSz4zB2KXh4Ftl1VISgS3k3Wm3klIimQn1WekY2doPPtwXsjrMVhhdvXzs1fq
46YKfynYxhYIrGI2X0l3Z8etiewyDKX4jNNm+e/xdvswRQxdhQwmNQzDzhLDboHZ
z04JiyykOf6hNcgTUlCm/11Iqo6sq5d5xgrzbSHJUZIEbyI5VYp3YShb2E7gDdOM
DUXGk2dlqL9E0y+QH8NtDT5W3TIGHeoeVRrUFOevA53zPqRrmCYDEAgJJZr+8NC8
3UFR+wPVaJ8qHzmRlpL7H5GgBGyoLZc3CnX5hDGlGtmiofzn48RurLB8P5ttErD/
Baq24hEBW2F/aK1Bs2JwgtR6d3O2JNS/7NRt2lcPdVHyNRSZ86IWdEKDhbTICDrv
MuEoUtAhs/3PZI/EJ5AZb19tCdZ5bSKX45/2Ii/NX/G61mswcrHO4+jrOd+52xA6
NXBw+sX4p7rbUNfTAqwj4+f2rZx0QMglCGopPT2IXHEF0k9xXhB5PBvG+kFBm2FR
y4zGEQ00zJY9GSyXIndEPuys3Rh2cPyaqYUGngkxFHEjbqVoUFyVf1xoI8nq8sQq
6zMK+SgRfAGSRSEQCP0++hdWkaaOWUwAv2/bKDFmBKBJt38D7K/fiDPx3Xd7pHql
ld9kVPXNBfZ1CCAbULCSqabW9+Vf5wGhduLfHGjQnEG2War4gDW7qh956TwKCYPE
D9M7V7wSLn0+k/useAjnf6/vEN6fqoO+iI+AOxMnwEqh/MrzggLk1DGdMXaZHSy+
4JT20xUsqHyRvTA/a5P/ct6NDL+W9ab75jrwngfDSF7oED6KZmvCdGhKIVe9sPIM
uwA6exQ/hOJh72aEybF4uDuXhKnjjnwa5eNcbbFC1CdcELsBZfwThnAPoxl6jxGM
8bAqTbQc5B3iYbG04meQQrwWaS5/1Ss2QPczWSvbnRE80lmiYB3D/mYanmw7FNxD
ldAjkSKKLjLnSoRjOXxEYasZP34kTQtZtdCvjnBgGe7QyTb7+D6s3/JpLr+0zZy6
LJKFRhyVvmsb22Brt6NdEFTFrDg8DP2E9oTY5gpQd/nCEjAvAiZICQ3+xWJPFTvS
norgPEm+L8Oj2ejQdAZ/p+d69t7MHnCjgW24tpKQeEa5oQEcdRMOpuAV07BS09p+
SmGDqqo6dQJSU+V14Cq8NA3ybo0nHiXSrxxrc5kSMyL5NmMXRN0sF/sP5jSHaoM+
P6C8fouC1AFGnuHOHdT9DCeJFPhy+H7llpa6Ihah34IKKmCV2BsJcm3mcB2BjEI+
dEgy4bPgMkJzdgHxAMxoWMLhzS+xW0/wAr0AAPTrDOrNrrGCTZJTj7RFLbWoFn6B
/nwxziMyMNi8cMQdCBrZezBXMfmDPTNCM99jB/Cs9Nn2rCnTbgpxONm0N5HEZ2in
RrAaHJ0Jc3JjT00xpjk1D02CHGz52qd3q4I2osvsBF/7Q8m2wOAibiU9Ok7yaAnK
YS6d57j7uoXTCdvwFRCBqe3aCBA2WGQrVvDig9Pnv6X1P6aheRYMGwtXsobxWGbF
nmLCWFPCIKrqTXFAiwsVvOx4EaczeqYnDnRA/2QceoI8x6DDvUpiUjrrsshmKeqi
jzg67xtUC+scpL/KYdqhHGY9I94USMrsqIqnjG6+jKeo7XBkcUockeRhoii+2fMn
NNuIxN+yvBASZHKlZBB0G91mYii7WDGHb0bqqzQztEzuDRZ/5rXy1cJXEKSiNHeM
GuxrJI5MBZWQHJX9rmdDMvdS6D/wAjecb5j2gipcs7DyjcXTH7AiyxTTiMigqfdV
3LXF95/kD4eFsgiFVGON05O4dZNiTZJe4za66ojJJVkcgzVacy9MW8rPOwp7ONN3
jWlQyqF0hyDup/eI1VabPd88nrqoK8UwCzMTZHxd6w97T/bYAV9skdcpXfVO2Bj9
p26KEmEX4M2047VmvgPB6RB9cQkUUytDeR/c8E9etchWz/ncOB8WpbyknvTWvGmh
s3+ToWjfB2Gh89CC0rvM8QL+2VZe2+sbW2kx1KdZc7Lrss7CxlHTJxYYSQFTL4Vj
s+6qwrfXrXz1aGsVk5HZEnsBkmtFX9qeeWvesKb/wOYPa4CTq+ML7XdP5KExrzXa
vN+1ZIT+fmw+h5vNp/3G4VKkbjrFnkeDMRsh0G2FTPFhdfBA3D8Vwg61+1RYD77I
PrDesmvskRZWNDKdC/v/iS+gxJKGbVOwIVZ7OXkfauxJXcIwdPmUKOI+jv3cfnAg
vjx/rRLK7ajGE1BhXJ8iqVXIJ6v94JQLj3oGzm8R421H31redWjyLFcxkTifiY0x
Y3z4lZDlcvmgihF7OK7UW6DA3RXeJXzOQq2VKYXYiVJDrpDBwJyo/HYxs47iiyMk
7m9/TW5leUU9UABISDnT1XJZJnllPwTci93RUQ8/FUxFgVCb2+avmm3eePBhC0ly
zcGYHy6vmwopVXttVQZJecSVZIJjnGZ5oOjeUAaT0Axz2WsB7KhSrARr3yr91NC1
KKSnsZY+XiCnj9pxFjdwKgWpuiauAfybqENQIGMR2p5RTfKShKoPsy7gVoaTAI6Q
Zuxuqb9QJBQR707IKAlTselo0v3AQvhUwtooA303nuGgz7/lhbRx7h1ag3K28smB
SaYplfwKzJhpeW5iriFsQzosC9hQ1omL+Q632twaOQ4UFdcsWOmM39T6mehLm8TC
1pBL4S12omM50UT7cJEho+dshgYhmjVB+0mAPMTy749gYn7yP89+TfCiALM70JXg
t5VsVCcG6Ito1/tv+Y3nAU9D+aujKzhKnoTcJ9ZGfzYzql/Y/WxMptOkdrN4lZF1
KQSZh10QdaX6QsLKPNw1iK0phUzCwwGL4vxdNCT8ZFNyTrLv69m5jzj+T+ssVnHB
lIRBLoaMmnsraVBtuWEw42XhTY6mttR1TtfCYv4tSNxRm4NKjxKAiTK4zBdNivpw
PEjDtaYxsxslW6yN/mfqIshu9zMTBv+7pe44GAOdu4I7du6qSk4lO1uFA2pC+IvR
xob9pCbzoAaI1iy2/DeaL2/gYf8mrESJ4uUu2SX38xYccvxGmqh+pD32c7GhR8gp
WyZyT6e3tYh2MH61qLIRGjTUGaJUkwwJkM49i3JdwXFdKQ4ravdIupmVB0JbEcJB
XfAZhzknOTWaXTaVLikAv4myLpvmtrcgNLhC8VAk3q082/hlkzOEdOwT58CpJY6V
VBchDOMPc+SGYW/baxxy2zwGVT7GKSpuXOnBbX6a1iwHrKDURMB1yQLpxTppUGj3
VeqnsARWRSrMO2s3bbqwOVKO9SIiTamar5+1g3TNKU0fAHIfpefmLdiosAYWHbJJ
p8wz/dOzZrJb1SlhQ44fGzJ+hJWeJERElx0bISe/c82MSsgWsvqweknLAeKRWBu5
KXKvITM81riq0qID7VWcpYDPEfSyv0/cc/R3IGycSR1GydDTDuznihhGPTey3zLE
y5l146+dNXpRDzgs0c/hLH2guOGzQKyqP80raTOAaYoQdtc91HI7iD/aN4caXv7F
RtfxUOZOTO0iqzL+SFw9Uy7R4nJJ0y5UskqxOVrsn3mr4SFtITPl4kEv/5bEfJuM
KGqV7nLj3rEHLT79Wy+JDsjIzj6yy0I6YAW2ykQhce96J9RVk61hOnThclO7g0ZM
7P4B98maujTfDnPK/Kv2gtdm1+0d2LmJkPh6KJUdiMvnQ8Wyd6tkP5OeohsMTh4b
4WM8LQJ0s3KiSZtTnLgbVuYZ86wT+pqc92PTk7PEtUu01s4Pyg8HH5X3FqNt9EHv
OM4HZfn6q6+OxtHHhhfPDqHwP02ki8ZI+lO+OJ7AVgmPkOn7NQ8QZDXDRvZmonWg
LhdGSspDGeMcP3T5DQ9PtPaeV+HqWPhXq173SQoAoH8865qCBF283fPe3haGuqH9
+SolQPxCQcD9ljTfFMvdAx8RdqtR7L+31IzAWHH7KXIK7/0464NrIEJCD46eQHeA
/OU1UL1VvQ1Qt3dfbpsw33gxeE6uh3QawtpdiOksYq/KeXoS17ATDNS7qnbJn8ei
zd9TpmVZ5RuIGw05qqlK9k/iqx42Q5jOHO5PD9GK0unlNo6KN1owHydAxk4vM/4/
2kQCkUfq/9LGqyEAaWQQ79jjvzTJmILJZ5vSgdfl6G73Puf2QRL6QkC6E9/PRDxK
kFSXxeVt9u1+zBPwblBAkjKh1Q4HDED3hT5Vz5NpbtuXMTfS1Jz096dHpc+fa/04
d+hiOvdIODwxEpR5pNoMDj6fPUUuxtAJLsohef8K9ZNO5z7J7V/MJ+/KeNIxJiaa
YaKpY+ePB6tWfvDjXCCvdyfhZGrJyznB7TXeD5jJPTK9kSsusZi27rP0RkmF6iQf
sUlkIUOu0Hp22zOHAVpHZ1SAfmYErk5lYTdwpaDCD6RE1evi1Xd1ehNVM3r9mys0
gLsr84VleqlNEjFSbL02vNHidSN3veHSFigDy7PVqHLmycNmm4SKdX1KvXvE3tGn
o9leddW/VZRfHMcaX/gRPfm0A9bEZ67sll5O+KNRX94nfzY99c4zYqzPQOIPaPE7
MLX2kWtJt94AEARIl9KSrSD5gI9wdbvp7KVUWsbhIlhIVx9Q8FN2CYD5WtRy/J4n
V4zuKwD5p/OXOB4lczrLp7FdcgBt3IQlRBpBTVUt6V/bylwKDrQgxOcnczk0d89A
qB8hC812/GQtz1Lh5+3Y4tRZ0Lsjc7QLbdBqbIIdLhVElXnAzQqrowUfu8cw67UW
QNAyD4qpN5Z9WFHGEqd/fYK+0lxSRMF/vrqcAInxVAVc2udExvy6zAT8QODoVoHy
6en+qFSD9qnK9R9WUq/YhIAoVZvGI/19Z/I1HVLcxgNchEMnSl21f7NqR80VvHXr
c7PX+Obc5nw4y5D4YKbAv1RfvOfmClwq20TnR7axJxU70diH1zg4KjfWpnbBJsX4
TxxT/fTxCJfH73NOL3KS5CvFcptNb3E9BuSoCICtjWUbrpsCWx3m0FWZH5HzVwOU
B7q/CVQy+/eNlAyRCu1nuPmpLd/jt3tttZ5Zv7FXXSgQKk7hh22/TxsynNqBL45A
zGZGqGSu3ZNVVTwkmGurp3KFQX1pl90JOEkrnRVbD++5r+ag90MrDZw/jfepGUHv
uYex7EVGsi5LeFqarOuceXfFZUtMGEMgTDTu+rnKJ46lnSeDNYDj67rHNNCJBAuw
LmwcgOH8SQyNJrhXsYBcMb4Zy9fZPtQIA9/PZnLe5sP8agv9B7fI/YpotPZkasdH
tPG4hmzTNCyo7AfRiK9FVfiTl2NBQLJg9qT1f/dSqH3SvrqDGpnS6GKrlJvOZQMV
7+yc78C6xHNmCA1oPOGaP3y3m7DYXDT0GtAexnDy0ZoX4YnHzqp3C3X/62XijYMB
xPIjHlgqZEUXwMPM2ZuN0bRd9T6NfPAT0UbYWXG/DNXJ+DgzjVRsUE/iHBDku3WN
xP/hct4TB4UUE6tj0MYlyNuraIF+L1viVywGGN0UMV8+OQ4AKtuKzdg4zdEl5ZJ3
Bf/n9oSVYWCVwrmhEFxKvq3MBJWSiSkJMjKqFhPn33LVssWz+UBdtRMyipm6SLM+
Pspxc6puJxLiaUjmqdJ++yWLHK5swDOnVrkTs7jZ7eQKTXXo0QIWDk/IlgxsHF6T
374rWyGoI+llBBR1Av512fH/VcKWMH/958n2a4+/pQELbg0KOE8jCVUikhATmh+O
gXMEd4ovaM1Sh2G34cSreerRsYB6+7Rm6ic22Ki760gk/hHFb6AV4Tg73z8zZ3ix
JsoiDi4xZx21LMsmx6cETUetEpX9HSDa4FZag9NfDbE/cpzBgiaCNp1TTk4mb5HD
SOsIp2gDd4TlZVOEFANr/SOV0whIXQSzYiqOpFAORDUj8uIJcSl5+QL0uv8/hDEW
9JqvaXevJTCFJmrxfcdq25KNSfsBrBPIPqs80+BVD2TgF6lTpH68vSymoatNcCnY
ByqdhOWputRX7Jd5TxWLOmSgH12+we5PIrhE+n9/MAdNewiDZ6Gg6KP54FRFTmRp
GODzM7zO2yc50z4m8NiwvmONRRNbJlLRrr2v935Gx4bD37lEakbpN7/qh4t+5f/b
9TMrS1F6WHZzUXyZ+248dqoAogwAqDvnAiBLVMu2INOc3V/0VQonZh9L4ME3TA75
da5r9ns+Q4immXoguNmDW05zHtVCVNG63m3haSPM1dTDzdwzy3qC3IdZUeHRdzTD
qqNKdaLc+yKNfha/cJ0Hpr8invn7Ur8HE723KLMx7MBn759FhHgaCcRMEZpBAPEh
jxUZ/XI9Zc3+Ywv/j2QAdCqmyqsW/ISl/jnnof542xRL6U25KiUV/+Iy8yXCPSfC
oaDL7Xda0jKJMATBHNHylPQBIJ9A2ZCtu6SxDrKs+CSnr9asM7F1oLjJtzKPu6oP
fyR1NYqcICQJoyTH4zS5+Oczlqg+v+o556DLjy+6wqhfg4nRJdC7w0TjuF3e8aaD
oBaU2pyeTh/Wr5giK3GHbq2IwDgl52bc9lgEwTJSr1bQ0KszKJl9jKB7IXDJowOw
hvgySC9VNZN3ym709524HFF078M81OxaFI6TqRNMsijVmIN22UGBvRwzcoP+5UrB
FYvD1NQAfgqBDM+YD3WAbWI+169t0uEvwa4DsXIIJHvCg//a6ijZxWGaLCkyxP0f
ZXG06npDF1Ymt4Mh4wMukeOdVQwSpDJ88CmQdqsPzB18wKu/obHJgzUlAue+F86y
RBCQ1g2EzWF5mW7DRGD0a2pLCbbx0gFgd9k/ch1mdj+6zFjL7TwcZY/uzB1Hbu+0
24G1sTJW+pK7gmokws15dTRXmDP0K14Ra6qgiD+SbCGhMUDCyGGouzEbva9yxVbk
UlRKtsgm/QOOro8x7H/ZeFgrEe4P1tXM3l6Aj/BeQvdbCyyXFgGDSjWATGheRMRQ
KpkLFlm3/DUck/mSK1eVyrNgG5beCjZSKQnrAqWKGMcxPLv4ae9+g3eDrBz3cnvD
wVPAq+e33bEgg5bZpIjTfLTZHbrfb39l1JoLk/3SdH48XYOT913WnEmDEf8ag8sZ
aHGEu42NrLQffvp8hQZ+gTY4X6/t12tcsJxSJOEjJdaYoIT/P43tfQFbDuTvjAax
LCbFjMXCrKdWkn6WUZFl1uZHotcH6jKwFagw345VwW3KsAj2Nf6toMmpNp8C4MDu
b+guPio5OqqRG9MSE4ZLB4UySDNKn+keN1oavBcSWOmfh/iT5iHHhynawbK8gxuH
xDH3Re23aRjaLUZQSi1Soj9WL27TyKuB3TOjFQuc0V5CkdwHM6ZzCaoZlQyGNWX9
uHR0MJcXEM0BPLsR4rkwayFl8rdGdjIFhX4WtVmiigg9NplfKBCudiFuPThOpqgv
KVUChrf6VWq4oFRDEi5aUIohRjmFEuyJtErirM0TNxsdmr9kBYreVOcX8LkXQf8e
GBVW3SyT4sEXlYLACpsfVQjAu5kaTHzAZ5PJvrM0242MYFJIM+HkCQLfM9apPwXT
SSCYdVN7/RFB+mEy3TeE1HuSih7UF01eOU6jMbhiCNpFiAALE8MZQCDRF0LAFJPu
UT+F5/BWk0luuOvgYUrDO04nZ1UbgrN2ltOazDUx27vEZnLmIRpTcM8Mb73pOaxu
Dk09FKdaggee1nc273XvG6bTbiuEHRB8Ne1Diqq0zJ8t34S+3r4NFL2ZardBErP/
macvnpx3smaSRCJaNu/KWQnHKa9wnm0tryZMKKJ6pHJ/AQ/rjz/OhceFuUp4Aw/8
b6VcAWMuj7HW2EP1tUa9DLqH5bZArboKij+hJcPm832TG8EZ2EgY9wrkTSbV5K8M
ZmHe+BFjXzFQdzO/MUyg8ctni3YBl3H+v7DHJ8T1MFrRfxfxqKJo4RYdwcc6OhHv
OZnkml/7GdFnZSXr0ONVNWJFBO3e4lXsQQZNpqvqF7yCF7R6QgA5JoIAvP6PQuYx
hM7N5MCKDhHu5h/LygOMwcJpRVLGkYlQ5klYU0EvVoinz4H8rOwhe67MFLUT3UAr
Y2FlG/HiRXlFsh9lp0cpadFqLDV4Dzp830LFcaGxWL1qNu/CYDjL5OCVeRMPlUrY
X/StFAPyZ8ek2J8wXX6rrCkGvR15ZVuS6arM6tAuSaz56V/n0SZtN4o6kyPf03UD
qz4+4T+ZUKMwvd0Ap3E1dVVXolaSuth3FBQEkg/H1InMUvQRfTJpMM1jBCWhZlSb
ni94eV1w/4mp5XqqDmG5XcpbsF3SYunLaZVt1j+MoO7Ik5a0UHOAsWiEHe1u2Y5V
lo9GZBdzHC0+uVsOQ/rn9b9T4tN+LzPwSPdD8LwljCCmGSkkStX6kngcNsM00xoB
ZCDMD6NrmqPvL0hWiSBTNffbWdbwK8yM7lbRD4hg4a13QVNEJmG8VwELFvkIBpDR
Fa7xYe8xmcvB1xHnokv1yrG9NSF8kTEZm+5Sb66lxiW/HM+8FaiyEXahiAXv702U
NtiJ+O5Y6Qfd8qSGqxOvPGy3uZLVwpNywo0E/88emy6LXYXRD5VbRPlyzamAnyfQ
rnP/Da4BRrvnmblTJ4BarmnuCFn5ern2pAItYZuur74xlcJCohkP7i2emVzAZ05V
nA91jnFMz756xaTc8VXYvvicsiO0JBlUCfs8hdLVeqrzLG9w9BDXD0kd4syrF0I3
BYRdI8BThDBDxQ+PKlcbJNR+Q/MApiKvu0gsa9WEJVzXFcbIn8aqRDIkXwP1ZEpO
PU3/9t3ydnvU1l4SbL4UfklqO+cydrHF62VWn55FmZiXLcYEX6mhQZSYUjqMF956
oOE0Z8hUsLPB61IUsf4RHzHA+FX/Qmx5BJPv94Pw+oK9v7Udw8vaCcLK+fBNhzmf
5kQRu1sI0AslnNILFsFiglyIz3POdvimsuqGh6dj/OLKTNV/bvXuEOypEnaI5kV0
+AqsiXBtkin4t1B259S2DcaUpyj8EFWqe7u5XZ5T9wbakn/PKOHzVqRU/hKTv3zj
1dEvAx1I+Tz4s3uMa+vwtwAI+ByGRBRb3Ks+m4Q8bgEst7sDCEXEeS1kkqaeJmpA
FtwX/nIav1ZmMPDqfeAOhjcRVoks+zYpa/LaoQaAO5u42MyRK5mXFZNSYyAN3Pto
4nGbDdoI9pDIqei+lPTFOiYvPAvIpvSRpvneVIM5Mtfu2k7I6OIiiZg1ZEg86ZTA
N+8ZZ04H1i19SLCZ4JP0nKGhVUSeC4Hcf6OOFixsEO+OmDhGwOx01eQ8PVl1EcLg
gM3piOfqJFNxhNzu2GDbwWC6MADcBIjm/dc1hpszE6vJLD0TYiyzZ3lVz+s2cUoF
WiCRW4OZdqRziEVjGwvmib0JDQIbqm87CWlVxP6cQx0Z26ejjovoMjfjERTbGpWC
tY+3jFq8tdvgAVUvvSGANXdcye5KyjGlx9Zky3f5tH3ywAzHFWvavfzVjvQu/eQ9
cDWJp+YwFiNAX6uXlhiEJmz3YGNAH9oD9ekUA3jPhOGF4H2s8FP0K61OtMZzL7bH
DfdqIHVc7mWVEeE7SNYq1L31HAoJ42mOep0loY4RLDhHujdJHFj8F4764CGPinsA
IB1AmmL8NPcfto6zpOvIaUx2W/aqc8ljS3jHt8iVQsxuzJQW/D6Y4wz7fHkv1zFG
vYS8qyiNBKhEhtir/VCJG/SijD2i8mgVdenUqyX7Jjw8z2lnXHt5ZxUlVh6166C1
Jmj1RVM7uaV3H41RfMO45JdH3eF8pxxxj3zUOzejdVyCVNtoR0CTAEjYZbb8OThq
C9uxLsjjtr2FCRTGc4Jat6BH1aiXpWSPjUja08kKR594aworaZJn1dlaKVKna7Fe
Q7NzJ15koCSStPS8iyWu2I3JBjxGp/Yr1SXuPcgaNhzNpz1lKJV2fYYEYJobUAi6
3gQ56r9PPC+5B1wc6gqyw4vSg9FgC3/jmro3uvtM5k4z3b1oiVL0SJ+Yqn7cHOlr
TnjYSk/xUIaS1XCYerIHZp7pHrU1ff02sLz7+gZg0hSZZZEfIDJIABFFVkOByISU
5fg4EdpVWIbYZEc9IVBoFAvAXYp83snhBuyFcrfN13adcxz4DW7Mk1nBuIAuqVrd
H2WHE9cy/sGmHR66qyT4z+k9voULtUKgSozdeR8GRZ2yyqTUp6dhi/hvA2ghdmRt
Mr1lRIqI062+SkE4TSHDc3IQn1TtmQUW19ejysVx/qpRaWtWNGfY4vGrTmvKG+XS
qdKuKe9CWnCk+H8oZqTvJPrFDXRqoG2sbgCy0P9JB+PVFVJ4FM6HZ8PSEKQ0P8EM
al+WMZGT6RDDXifMqywZA48+CAR7k2FAuWIgakwWSwsKc9ie1JtTtPJjdXUtGbS7
oGPZ34CjmEkuRZmgBOlz8AWVEyccI4YzBQzpZYT93C3ybgexi0SgICPbLWgUzb/v
3wQiLcYnZw6AOynAmRiMCiy4v1ZxMcTs4eZxMD26on3neCG8WLyFgtsK/261gGka
EJuzgTjVQ4OZ/Z0cQfwa3PpidJ1RqFrimcXZqJLK/ta/RPuoWn5OGrXN6zUHGA7j
+z9vV/UjHhRuxM5flsWRsOCIJRFtfaF3xw6WC50Vbl5sPiOWKNkgDBfNoWb8g6iP
jcr+eK7Fecjr2TrBJT625ev+3oQiENvfXQYJL0kv0hoafw08CO9HCZzg256+0F2z
jZXgyGR+D6yAz32lUH5uDWQ3tgbI+IKDglwC/e4wPf2XWqW9/VPLeRB3wZZ7tScn
o4dLvUjCSi9a4KrLruduSA/Nztd54OcCLfJPg1herqPtciieBrERHvXjXTrUhkne
Xpmj321w02aGjNk0Cf1nrYc4PSASGPaBuliHElbm9v0o5HsWjJCg6oUKU3VCpqIT
vCwHv1HgggeIbJQNX1o13xM+sD5oj3fS/5fFsOJEh8JgM1yOaavqgRTDDKgo6sYz
5c39iCx1y0fYmnN7eWudS9xwoNUObyqb0hvF28rqMPGWW/6MfFkMlANSMk/gKxej
PYJd5tPZQpWmWe27OJOUpq6LFfN90k/kGWP0JDtQB1ZDnKdwKKoGE6Qt1avP/mT+
mWyV8fsQwiJ8XlMW3BdhBv7Myvo+IyKSn6qEqn9VqkzBiir7KPXf85WWa7U/lF3V
eBObEuAytjUwjcFQAujUrlgtH5Ns0KJb/gShnZX6815+Zt/ki7DL6MkORIcKOl0i
A82yKDjAjv0vKs2aOMyalv6G199OmEFaV5+WVfNRvYiKzMpw+TeKIhSU7OAVUqQr
WXV2FDCnY27w3yvQ4MBFf3W5d/fkJ/K6w4lcx5hnKHH5HCxez0r9AcDn/XA3gJyW
nNn93tx9mxqnwIvyOOyd0KAj/jnsPr6uy9vncU3WLhBQ3EdOZ+Nzs4f+q6NerboT
WExSlTY40JcBuKgpVeD31yNpkUne1zJvl9SoFRaRt0X6IvHBNygmRuFpOvMOEOLd
b7K/O5jbOlQ8EwH4Ns97PK+I617p3dHDrv+jDAvISXpX1CIj/hzZchxGbQGxIPBl
dTu3JjlGYGfQ1xETFX9Ve+51VnrI6PlgbVXCYQ+i399ZTm8l+T4pXNuGRE/ySQMJ
JpMtXHt6SrB0O1klL9ugleqBxiDL+RRs41KnHqspFkdRNrWeciadXtNm/6dWrE5T
9iIsMcKoQbVID0mwHLEduxEw/ZBVfWJI2f7JUU0YNj1kc4FzaPo1uz8m9J/f1Pl6
ctyvj1R/8ersiUQ0JG/mWmCYt3k1kvrDMi0344BcqnelrTl3meEMWI/1NJWbfeqq
JCnYnZCMlQGL7TjMcbufY+eBKock+woO7m02kj/gyQKjkTIJrqkOhxmMbLiyssm0
io1e4WcDcVnfs8E2rtUeyMp1+blDoi5YNqK9bEHtcDJczqec44bgj3SXHvVuy51o
nhLK0V6kMdRecZ/eUJV89zKlsrTZzgEx3Jh9zwdYpjQ4TZp82PMAkg9jUgIdXII6
m8CGfvzdN6a5k5T5RcF2L1p0itb3cDWWVZDMfHdCubXXPK7gqKyKpQ6U7/fxdrHa
Q1qKYs7tdLXAvzQOcgKX32jXqCb+gYiDR2NtGW0WMbJwQlln0Idp2jT0OWHsHBtY
Q4aI3lXR5+0HB9CMyxwI7XxcR4xUrcyvMuGvdfemIdIIWSA7q0n+yFr0J/SJAZCv
XSe59sNZjKeqW+3Q6mUtH9WQKC9kJ0caeZomYgoUQOzGx8SnkuC/qcQ7Wa5OUYT6
v8TVkhEZ2PZmZdRvMsK1z4rGazife8Z8chg3jzc0mZHZ9f2mOS2n+zh4hunN2Ds3
3wh+/Y7imjiKsxhtf1sbEI1ZHQEMDiLZUYDs1D8QXvf6SQ9udUXTQcWMRxxPp5iO
cgnHWRDUz35if38EpZJXqYtgIS4DC7tyNXspkvbC6/pvQ5HSGUbu4Zp/h1SCalcu
1uvqc8vaID1s9Zu1Ut4A623fPkMZ5ZcHPhx04QEp1krZE7BlpPzqZvzvHZSLqCy2
QSO0dw2a4FzyzuFgOH528uzNJXKpN0HbknEwViOhe/LJSeBwgTXAzh2uWubBvo0h
zd9sJ4YUWQaGUo0G93mg8tr4mbUneHpBHcaaSlktM/bUSbgGph19W3RR4jhdaMTr
NNVcs58zxo/+UwNjKSoO243eyELx++pHCUqNRdQtapgy9InuI+N+Bwqh6MJcowb9
7vY26zyqmEIXb+v9jBrMUroxnk6IKsdH/fmupDTbgdpp29dcz7ru2tHy62BIWgGU
u52c4TOrJcK7TjoojRnIVT2Q33Hltfy+qqn0i2bF7EWtFVioZUcdXIzniXY0EJuz
nvdd213u4dHhyvcMccbKkBtqfsmat+P/95EDtYGKG2rHi+yhsAUba24RND0EUn3m
7K4TXVr4elI9/gtZT/FIP/feA8iyauCtqNI7T2ThbngjB+sIc+dcMSow2ttWF4cQ
ymwwvneMVhhjNF8/woyqnkqFOhI6z/qMFkFD6E40q64uqjSgEzmQ+0QmTkn4GvIM
blKv/j7xRkBU67snXTNnxowKDkFOnC5RbMVzWvbjzshphz2b4YTC60ksq/LtdPTj
51Wk2f3tzTFMl6ZtLsfV6hRoTZOysk8d0IPd6EAVVI5cpk5uBDEJphGwYqKTnvr7
vx+1s5I4CNka9Ly7gxQCUNzKkcj4nXdrQdVv/Qqz7cUvzUva5+5jNvVkpce/BETV
0j/Fh/3w4Oo5mEoG4xheIR8tAPyaiSD6GhUyOJvaZlJH0FppdmFlmlCZyFVSVJeX
eszwn7cQK1mbVy/HhloM1El+c1jBAVGn9+hPmzbaOopKeRfTTSZTMHfwzCyTrVQT
XTnX/1KdJ0lzPcbrBQkOdqbkL3XcSphfC1MvN6m9oreVSy2yn3342ezqTXtq0kJI
vO8ClQURgBavEoW+w3JZnNVgdVJUv9ocPWfpYKYEL+9sJ78RRl5Yw33pLPL7LbgU
I7O0pkeuAb18vanwWXm3a2upFnCZUwrBOpYqv+4etk0oJfQ2Y8GGTCF9zIL9rcrQ
ZdO6yQPAx7sXYg+tV9GlGbs49e86/vduA17CskQ4u4v4XSXY380B+9Xcx0lBknSV
J4/FSOB+8i0BpAkQn+QUqxLMzHQPo1cXHMwuAiZQomrkI08S4A30D/ew2xmERmOO
Kh1f3xrMEaPbwAzDMAwlXndE4sT9pEiqhX6qy3kNCn8ZeWNhMrvmu69mp/PBVcf0
UQf3ls8kU1L9Qa9f8cz2WnXLpmv8hng7CwlnGG72u1VQkDGDRvKstYYKaqDvSQiI
7RJwTBXLPuKv3mtjpxtwU2HAWOCXoK755VaR1Mue0lNrcKlP8FaI8C2f6/S71UwM
z6tR5eMLPjR/I4fwNnyNFfgcOWMWeCd/77sK+TI4v1RzJt9Z8YO46MfceRLjnLbv
vowwl6EaTPZjKKVGozQm7/9CfxwqtSoZrvjhBmf3KCxYDiSlyOuNSS2zrsezaoDM
0Wo23LKEc2vvCYA8mu36zSDpjcis6OhnmrTeGuIt6v00sXWMFnKlWJ0oS+mWYAep
zYU5aNxzfySq+mGisWD1TT80EvqJSPnJlPFv10kC1L6m+meTMTuPtNSp/WJCun0h
v1YgoIjcFN/CKYbBLf3lbLmFqWee+j3wW7iF5BoFj2Yk96roS7ClH1LS8kR5kxqu
584t74Av40C9jb5zo4mttqlA702gRqWldxTzQ7jTV0bmVYdIFk825OhH21O1zfka
I2l8aaXdctaX5QmhBZ1J1C2SFK4G936ZP7Jl69/70krgaFZe0pxbagtMVzqPxCbq
O6HdzHb2nNFNwxpBzwgmyRY3wclBaj/9GyhzyHCYLiZLBaok1G7ORUEZKTP6LAdK
bo1zmQ1auZuzE96BSMHkYEEVSnqVbzlAlc/pEQEecDo3BbdKLmZWPCwYxyAUJaGk
c3TOWpRByiEw66lSgetse/zTbX0ON7xQobq1LGmMiWl8IY/bhRVR3Ck1bkr52RPh
aLQKEGQ070KgWjS5tCqgP2PoqnJDbOUnZ3R9IdC3u/mGkPkRhMBDEf22QuFJnYw9
2mOS813HcoJifffoc6OALOqab7BI9/pMXFMV9JXYA92GaMi+1UjvkTYAjx09I90J
Oy1n88rd7NAcV5IUxBwGckX9xnAUv6yj8Mox2fRCqJxaDI2+bYBvJrQBuJw5QNSO
wJeVSC856CNiIdR4xTo0RtZa3GHbVCSAnHxQZ4EuVb+XRLcQCDkeW0yVVv5rTTR2
iWO6/ODw7YckGpyFl8jn68hxL3Svbkw7yBPjsNoR/JKYYOmB1VrkwYjXOmJmeysR
Bwluu+Z1lQrk61ohWud4A0yF3eloi0UgibxMm6+1wxlNpv2GVmPdFkDj1VknLTbK
jFlz7hJQvJlQQsDftu3rm6fWcR56/j1MPBKGAo7b8KCogFqF3jGAwah9vfGpVNoN
ZQcGAGCFoHVBLW2q/vm9gwNVC/qtGD3J+dLjAPEKM769O3jJZZ5VH0B5mN9NUu7z
KxlDS8Rt5XO2aYRzzlENSU4ky9s7xCv/p3JxFKMsiEin6lGWeTL08XacZLEmLd6b
okcDBjbWFQ9/MP9OnUMk8DdY9OF1DHH6ze0aBalKEoO5lDtGivjsEkQ2viWkpU31
9zi71wG7AIN9oKjxyGAbfK8oGo8nII3mQ5VfdishDqnSiwGEAxT/Jj6SyaWC+8+W
KN6OaaBisI+dOQkGKl6dpX2uL++99UVFjLEubRLGna8JuyJHO9DxpU97EBjtWpQx
wUXPYHerSPR1REGspaU4dFzKdJ9lxnfApL033mIrkenaBCV7WCCyu/t2SElyw1i7
pKVfrB/vc/s2IlMqqswPocsy5zrtv9ERBQT9JnrNBRW4aha9Sv3J0oJ3k3GQiwUQ
wllQRsTmHIni9B/iwoQTjJS2dz5Q+brkTaFu6BqreitRy3JDiq3FhAET3+8WCF6/
no3x1P1tWjNk8ThXb24z9YVfxa5XoC62NKxnKWSGTojsyTM5m/d951I96eBtiUgJ
sFYGFdXg07G/5FC6QjYK5j+EmGM42Oto1LN5Bupx+r2kWYiG9snGtFBykj/Ri40H
84psi5QEBcfXbIFwID3wsdiRF3teiD99IdybogvMk+KW/a+gkTf0Koj+8x9B/cLC
9qF1fYd5a5bY6rWQtbnH1d9ZX5/ntkBTWkjUDZMCk/64pN2mf7Taa/ur+vObaKC0
tVtGbHALnbVETezOLxAsL9cU67uCfZXFvVDRnBQggLhJ01a8hL/HBLr2XbQ+Mjl/
UnJyTHiBJ1YZX1E6xX+tAuuVXEO416B7RVMLoTXIwtF9yBjqOFfft/jL6yP1fvnh
222n5+HVVDHPhTOZqhYsglncmJiyUdW6jVuBBid0zAd9iFHS7Y8qDZ8E+cpmKywY
6gXyd6zYKLHG8a3qkgeWO+n7+6v4R+WWMBgNterAk4L1O4fBkaKHl4QimpE9A8tV
gQXFx+xC7Hk5VNmtYnGJ018Mnk2nr3+S3zmcXlC0CGCNKJM21JmqO11/0VdLxR8a
+6fzLEtwokGU/H8sDlGWdll+iE4ryE5WnRpdmGuiJDBtR4UKqN8cbjZHoKItzxrD
kP4FFciM7JV9qlAexhAPJloIKUcCzEFLJoWJqB36G2hrQKdDbMkesyUe1d6B65yv
lhBjbYHQxYcI7l8+IwAMeLkHE4bMgPMI/gbTwqoXRKADnsacXNrvjbIzf6eB3Lo1
tHDrayvCg0wV4lAUapyaKrjNjSYjloVe07PMF6cOyHEyW/bxqJwuRxqciUw0BRUX
tWng39qos7j8HrSc7wchuBUoH78gHtyxUfTYsqH4EpETTTrQwzKSoraOcxj/ADJm
O5MBDIttVWebssZwiOYMEUJ+8iaohakDGe/HwmuaiuWCCptrKajLXcRZFWLSs24N
ezGGoruxzbNWuFKRp0rTup6poJSl3UW18S4H9AyvP6Xg1wYViivDpyGUuqg31FHv
C8kuekkHSr88krurtTwGqdMMHwLqG7qKYytC1CGNPRFfG15rw/+yBchO6dMGMNmX
WZNzFhl4ZxZxsRwvETnhJQXyaIsISKZXiQQoOYBLoAgqJb7zUQ5lcHTtIqED42i3
gLrEDKcO/NehuxzACKt+cSOSDbAyir3YJ2B0p9OGRuHQ679ra6Jhylo3NJqou5xp
PM6aRV9dw5aX9PzGP2UYdCJAqzr/FBfB9SGD3h2avGjUBxOCOGHQAJB8GEPXRSYS
ittr7qizWnv/r5lNRxdi0f1dHAExbhKkmr4wWSZp/Yxq49VzCvksvck4lu4qPU3d
Pcl608tI17VqSGrmrNC5MmDaX6z0qPlDzTJThc+RsBhyuRQxdR70eJeHn9CamlMt
gWt0Rz0hqAuMqCSkgAiaI9J3Dwq3DQ1QMH+7Jr6rYrmbe9HUtLR0tyJ735Fsi6T0
CJOnlwvEgWaZuiF/K9HYBM/AMCvUww2TWHAGvVP/kUZYbNyoUna85jGsTme2Y72V
DpoyxqgazqQ7TKO6nqTjj6BVhCDAyDU+8y1thp6oiiNZbJBEW+VAtMKvDB3ztpp4
W+ogHMGbzn0Uc2z7/6bWo94g1uSlw+fwEyhou1J4BnILEI6eSBVryXbBrZjSpqW7
O+5Rryl7uScFetzwFYl31J8KGpjy+Cdy7kiHIYLssWoToXO9g3sMrcxuVUCMrWqs
72k4gmcBg3o94V6jNE5ILmviWkpto06LepljAltLnRpm3EZ2ulwaByxVwUeDlHoW
QVo0/qAH6gA90oAq6WYv+oz2eVePvnDzQtHbNhKWO2D3Uudalrmyfwaj9efImhRm
dC+mzwqB9035etBj3k7jgXPimxFtDWBtFCTP8W54sOKOz9zOVfnVjDA55z54AFGt
O/4fj2teDOUwKzOjC8+5E0oP/2mCJeaQJbgObsp/G/wXsN9rx/T8yYUb/TIvxIhI
VECEIwf3YySyQCzuHxe60n6l1FTigpR5EwYNBuiQvHd3bjZ3++2Bt37g54st023U
15GBGqk66pnq102azV28aLJsIRcoWPgJQByGJlF9hhlWj9sN01grQJ/aIbJeGxqX
OzGqGN7BvRwS09pK9xjKxMZdPSH0I4bBaRoGIBnw54Gxn191B1ez91f415ecGdv6
+Xbp/TZuBfzVTzs3FpUr4VVMCk9WPrnmL+O7CGKubVg6JgZZniegeJ2dnaJWbtx0
chegW9rKAxyXI1RDWz75PAM5+r2Q8iK5lMF2e7vEGtRI45zkkmWdsBEGLLygZCEv
e53JkRBi2nIyDwOW0vVJpuoDTUfAZyjxVbE7AmLZbIiAcT33K7z4GjcTLCxlaS/J
+AOy0FjmXJ+ozyfpFeebT85iPVcz5B/L6teTlJm3uRW/AQdnUa2I8MUbMaEnPBq7
zCwgN8I0ar4lLiU1a4oMG1RNDp2rKp55sLhc9iMCUkUoxeHQ6emsaHwu+VwtaNeZ
+Fm0reQ6O80N3wz/JpNkCOXdH15/eou0XdSlIa/KJwg3O0m5YWhXT+Cs8DS/PGus
lnOfuwYz2fiPnf/tDQJtcuCRP2of68HqAYtcFRVVgudVLuEH6fj8M0ho6TpDI68z
u5wdMyosofpuUwphOR4PGv00wwrCY5mpZEQjAmYK84nMYACNqDwilKs9+ZxvGoQQ
rdA0PGZ1U0f9BJHs5Vkwdeipl3TTphYkwIBx6X4ssjeRLPysYxx9osKdTTaTw84/
zVs3Qq54Lgbi3/n3AEhIEv3kiYECT73IzIJh8ZTZnNaFLaBVYAKzbgMTyVgqrd85
pV+pTXCMOd1c2fEPO4BdFp6PgOVm3t1QFADT2BgmUSU/71IJ6665u4LQXLTdTmTN
WHTCPbSuwZEChlvS+ZvDiaVnNTnQWyibIFZXxpsrkXsmeZdTHIFRka91MVuiiuVi
62wTf6zT28sm/kz6wnGOlxgYv8NepLtVMsVODQ+DUo8/gbrzGkAx7pO9D5iiJH5D
tjzywKO53AFzhTnss+yAZX0IqJiPt1XWo1/zsTbNW+zseWAQv+KvtGUCBfPJmnjE
1aTvgY0tL8hVuj4FDpXr7WU8YZxn5aaFlxpp+4/B3BF1DaF6AQs5jLHLQEmuW4ev
Qfje6k2WHfIQG8zqbxifW70v7A9kWKGtLV1RgkCC8CsbGwIMDP1BZFoTB+p0majf
xstJJS+1GAbbFECB+zW2v6/sU2J7NdWUil0TILwqzpbfWQnzvMbEEKYo3elsmQQg
AsaTXM5M9cothWE5OU8KmNp2iWAxE+WqMW4xq6pleURHpgZJvpR6pknjLH2j4MDZ
uDvtjOC9ea90btahq/iqo5PmMAP3XCeHQUt4irJHd4Kmgj1+GuGY6MUn5kYOxgRf
nf+CMy9YoWYCKPxJohcTTAJU+lZj1h1eKfI1LFb9N+IJs9fTexOsp7u4R8ibdkDE
k1IjcmkxTfNwOqwaZxOGuVXC/ob0CvtoK0P0GJlXBCjepACsLTpDR41zJ02NvVHx
eU9ttt9XywP29A9AUGWm/sZsV+AOAsk4iCKtNoflynICsJD/rc3FTj+oo/mdol04
VNI3QpRaYNyhc2hzS5AoQch/UrPJYYvLpvFxuEOys+4L4Z8salW+xWCs+eg7TrUr
pfRh01pQ5a0VPXW21Rx+SFmaw4fVSNOkY6RCktKhIGGdj/9dgZkZ6oA6B83tCStD
l5VQGn1XgaUpXUQ1ePK33dp7nDJYJJS4irz4hD+FkKJUXJ2Rq5fK0OVFDkx70TcS
sY8tRqY7OAVlABnayRst3wsX8i21N/xy5VZIDE9ir/9g0zJuwS1Du9Zs8rXoFgHx
UH5dv82nnIh/gOFTDUcjYAC+UQhjH9GniiAXqhrBLEfq8VNVjTK4QUYoLBAAgLrY
whhCB9kMW3i5cTGewStOZ4Wm/M/WoHgZPEosscRQ7IN4kqs6HcqwHPls6Qv6i8y+
u5S2kUvCJ6nZuwGQ5RpplyGZ6U2FiZJQLCAcLLJ+VY5u7sVZeSyq9X7EuwsBAojC
f9F4oPzNUctEN5QTlK7O/AiKMRUfrmP5fRz0sBXIOCYXHK2Z9rzTf7f2CGseAHoB
PmJMW/i6WkLGLJwMzwrw0QyGlX3N6uBAIjXHb4jo8DvzD7V3QsMTaELCdT2TDCX6
xaYmWTdb/RxMsyqm5kK6jvbxdXYfZsovIi91yCi6iJ90YNwzw61MThaCXlPu7jP9
O26dJViwK5UkQiMKlFdst+xR2DeAVnt0oCycHB5jpuPrnr5pziDMt5larcuHxMsM
etGPn9Kjk/O5wAsrfRdkTWByGmxOpN5pNR1T21MyUL9/b3hnXU0WJF6PBWrzqgvC
g1gtLBYSwFr2E571oKdIIFLLD8mn0N3htdNU3aKrV9h6SPWTplZMhbtZGSn+7bD7
SQmMemeOJfT92yLMirBXkcxgKNGsTAMwO5cy7iBIJHEGjigGBtHaApZv79vqq54T
vFLeMSVw3UctUC75MgBhcoaARp8qUK49wraicK0DBv7qIGD6Oeah4MwfdsqoYMkR
BC61uVim85hVxn292DjAw1xnkCiWA3X/pJQqK7KKoaltFYiIkZuHExUGZiWeqfqr
u50kkpvI3O01CkPesl0/coiEz/gwYQ09DH8H6+MmSCu60voqSQ4giLpJCwlVu2Aa
axivtUEmjLL5tBFBAFteReSPISbtTMy4eQNylEdZBlmWQFOEg3VQLpojE6VwR3ZJ
kkedVBxff8IWiG8KCkGMSDIpTrBUi1xt4qNtGfIlva2qvmVA654ANSoOtB/SJX/E
UPnIROAGjb8G3k2XXs6AT8XL1vWDmOxL5N4fH4OM2f62qNhzI+fBD4leRdJ9RZsA
BzUbDsn7Xfn18Ae/uxY5YhEHaG0QRk4q0LosoAqNJcFbRGOdX+dQapzY3livghOO
r53c7ROa5wbLgDN/nJYt+lUmvTr9UQ9pvDhNIqHTWXm8kOjwdiHN5efLFqqjSUOF
wQslxQQ7zQx7jBxiES5+6b9prBMIiuv1gf6MOoNGt7Hp3OH8xm36rOFL4L3qlYQi
obSm/VHOifFWsrAkowKqeUlCQzNGm6Q/fphHNjDq05742qAuxnCE4wghHxMqoiSK
UjXTP4b98ZWs84zxWfdfIRQhplcMPwSqszD8HqYXiNSC08xu9Z3zthiu6TZJ5qbv
Pyl1YaZVAuuImfe+KqOopCif/w9QtQi0W1QE+dVO2JJ4GzdlVSGf2c7tWT6ci+OU
ZGGp4tRpFFwkDuQaIvZV7p6TpnwDX+gWg/ZcC++IzHu5Q/tQwARvfr/HIXugHex+
gdtyBlbsliExcbN1TKNbHXlSNcFup/iqxEepgLcQ14EoCAJJf9flSSwjZnLxR8H+
bDuuk8gjkX+nzgrDWGsiESdka3omvPnSUW/lLMD3K7Jx+IdMeXtPf27ox36IlfCW
2qg6NrRhEy+h9IXGEI8F2EaGrG5HrA7TsIhRu0MZ5LsHMgVwD0kQDJzX8SPLHruu
O4GMKYKcGCGDQ7Wj5Ud54aMaZej07SFeV58ZxOOgv3sEK8p+xVp/JzGBf+xGqhT8
2As2/Y9uPF47XgaU8u5SBBPbtXnxbIBWZjWjcPYqf97DnoaAKy18r203N8OofO9q
ehBCvoVasaNekiniVFgxcGfEu5LlJ+IjCL/rPDcM8kt3yjwHuO0koLFoZsIgOXsM
mz8JxB8AOhc0DacvZ+jK9UgkUCtEwJ2kp4+DQkmJ9DiyH6jv1Mapl98L1n6BzhJO
u3dDX68NEfEul1HkONrTMk7Zj9/ExP7HSo7loH3XZ0n2wZalVRdWx3XKWDRpr8KJ
5aHUccEjoo9WXNl4aQurKVmhVhpuxaY/3ojc1HQVM4q7yX0JwDT5X/pDCOBgNY8V
i/3WpEbAIL7cnp2wgVjymJUHqE/IfrIdXinmJRSqE0dKWMlm9zApThuYFR3UWkMT
uy+KBYp/aHQNQ4nGo5kC8FkfmRiAvi7ypF8+T89XI4PyDdgXsBrRAw//tIlKPGI+
Ug/NErvR7pOmesSYobyxpFSbcRjEVR6TLWkOb7TVVICBc5BymrvNI5XWPhc4wAUL
AbCoIj4VJJ12HS2GM9eMde+1Xn9/d0V+EX2eHMp9ZkTXeotufqSgimzBNK3QHfyx
YbGGudyYm5cHrT5/Hs+viYCJx0NQAx0eOjJG77TGKdXn2JkmqMqROdI/iZSYGgUw
tBiV7cwg99rgKUmYJNCx+/LZ/ng0JqyW1Bz63hSlg5/U3MGFI0G4rtwFpQ0XP7tE
t1/otIFhTQHEXxr9RXSa7zV/2dX/K0YIb/vDdgC9UJBUU0gj894lOWMA+sOdDmWh
l+oS8nSlv1F/htZMdSiASJsnazXzd8EQomRMpqTdOQSgI5fj8NcdbNAHF0SxH/Q1
cyC9DhGY1YfNoLneGUUNMi9APzmFdeCokLwHftg5/7NVAkE3OztNbiQbgw2SXLRx
QeQhSnAB9YNaN/VtCnVOdawFMd+AZ7XkKcyILP89FBOXyzbO8vTgeirp745WudNI
azgNx/hvJKD/Hr2nFYfXAlji+RaZ9llGPk08gQAxZQDuxryhA0LhpNDjnZuJ+cn7
ROcCgbJLbp38RtoeryXpk/+YlAuaTcrt5g63QhSCHo+LGUGDsY3r2sj0iV7zc7BS
yxHPsw5ADxDns9Y8tvqXbI/vDei6rhpaei1MQkByqJYqkiDAaoreibuCYCfecO3t
QSISvl1NsOlOepv34+Oq84xS2cXplTgdXW1UWiRrnV9+xcZpBjTNtk5i3Mjhts/E
UgKm+7BAYj25XzzkTIfRRVHvB9P+fPRTYir8wOOqbnQ1fTuCm+AmccrWkjJzx0X6
8jI2ocNf9418vhvgvwdbo+4DQqXZb9mexxXvioLWtr/nbz9RaCPcmJ9f7pWgHNxR
jojDG3ceQX7Y+ltV721nH8E5XAiL1BbeYz1PqXJrbccDua+2tTKJM3+F26xJXiPB
yW9eTOQZ/JBCxMOJoKPICtlVRsmdISsFnIZH+kXParlVzAXGl0aqItZBo3absCeV
keMqPKUF4yxB/MB+vN/XWOga9lQcEeR3RZqjP4Qotv8OL2Vh+IbowOPHHxVrSnxZ
wtyJsESy6hBpDeJYVUjRJcqIF4P2eiYAVvl5Z496aYpEuRcBmYSYcmtzBrkec8Bf
i2ixbMXkhJBPbHCXG3NtxJ+Tlrz3mCPPH6/1fqriU0YMidmiBJZrPUnPjrK1x/Wk
lkAQz944GZQfhw4pPGnJrkrsXyTDZVQk0EMYlbxVgGAD6PELvXZ0ydxOsVDfGQgq
UA1vCXUvRvUHKzaczlvP8p1VRG19ftj4H6buLYj0qcxpGqmqEhUd2B2HRX0euivY
CVrmlQuqp69fDrCbMChZWG1kvyuvgvH9nQ3IW2qZpbGyHS+qzaq0ifjTst+VIzru
TKGXLHb18BZwR6vr6iw8dIS4f85Y4nym5yeLhHtPn+rp/1WJ9P7jfGqDrlkE39oe
2h3XAmOz3o0nM9+/LmQBfNnlBCagTtqqVLQZleX+lchyfBDyMzMqgUQs7d2InbjW
azVjrcNuzgl7jPOysaHnvtMKRlVtp2PSf6HZwILbf5Og1voMSViPosXpaG3DX+Rn
urrJLqm+cWornwhKIOjVTENzX3RNdhIlYX3bXG2qSQRjtCQdvkeeHB/6R4Ed2Cjr
u1U86W5i3RezAsGCrr7R4wGxVRC7luEqKMhXXA4/EoqXGzWjMvrEXMjyQ04R9UGV
IzIH8NFfjKWEU472z3VVV2cZ/A2hIrlNVhCsm1I8S/FsQN1IlednFwOVBjOQTXBW
+9jzXT2YvhYOmFq9WmRzmLy048V75sVPrruujkwNRhhfL8y5dzKMQYLLIhMkuN9W
7vC7i4NrXbqQDXD7QT/EK1EbcqlS/Vb90gf5clISXwEFhqInZBaPhHRZmEy10g7V
NETc1SdZysGzN5cJey/BwknWq/g+1rNgFLgovSYORHrXjzOVlpw+14SShS8wQVG7
72NPcp1zGgcen+QyzN2H3KmFaQH+40zL5ngqArOojZy2gTfZwUeap5W7F+OEGOiM
A2q5t6mRDZMBZ6cSUJiW12/nR1bqMcK4WNl/Si66MoTqVBmft8APXXSaVVvwV/ML
O586rO5uhcsr85NByY1auiIQ/AF12uXTTU3ARoAcbr4LcyV2pD5lR615rOtpgmse
eLtzVuq7i4inonF+OLvDp/o0Ttz7BFl+o6mOWpGvVk6f3WaFg+4F+JVyLUxwzIDi
ylnrugtSXylPjom+Qsoz1Rd1N2AeeTwO4xJfSvIYIQuwwt4qGJ4H6di9INAn7yry
qq5y9GHfXjOl4KJHjAstccLt1evgtcKI9R6CgwHaZ3KS4TBTaRu7LeHwkEKjbONO
PugktrIEBcHQqOj01yGvxHcj2lGxiQDPeV5fz9ZyR8uZy5Qi9MndXMKptnTGU87v
Nf1DFQU+40Nu5vpJ6UAxnkNC2ar+Ix1s/rI/PmQ51WXP+iPfwkum7T2+D12M3IZd
Qu24U+GXymNW7IDmPrwPWZO6MR6bLin1rjvOPjt+SHUE6UISm4HcNgvbBpxb7WBr
0hVecpu9D4yQTlLU65M2nx1gY2Ub/RgUyMZpYnYy9ETcLpHYrcwI2IXdHMN28D9j
E/HmJ2rzu5X35wT3pI2q1TsVgS489fFPzIdbnI0AqzKnP7EEN0XV3/VmlFpxWYZb
+cBuOx5J3pyw+ob9GRfFPf7IB9jeBRSl3QRe9w4U23jVVEUCfCPpHljw2U1H1S6+
Bz5C0a9sq0zzUeqOk2WqkKlOvhddREwsyaf1ZbVIFnsT6vKPI0ydWsyxDUszw3/I
pR+gUjYCQTADxE/K24TawI84PEbbBC74C0Jzji8rMxjkn8pyKq7uw7eyabXsaR52
eOdrLlDn5BvSvOtXmmkIxzgyUuuK76Pz61eXUHWmUKP9BnJM2VoCLvd5LmAG3hVx
rWZQHDN7bwi/Vx2Be6jYg4zTAxpLLz3l5WASivcn8Gj9+nRsXoTc0N3Bs4xXCuws
YHu5/BNNqSXGskyDn9s+bMuGoD0Dd1ZrcWE7NA61th1fToyUqA+rDQ//iQ4e4JKl
VNHTurotkqKw9RrVzmyh0XywZ89vfN2NaINqC5M3Wk1iSn9esHEDmKu3+Ow08YRn
4ndJ5DDj9WiiJI/AF8dS+9SJrWXjU/ty5NuR12oiJxOfuBmYG9kX+aL3oROOlhZn
I3pYg8W8vv9+ryZNzIbkOUPP67nAjWnr+0jWH2XHpSsDVf2ZBSCOqsqCuHm1XEDV
oor7wtOzclR4i9R+K71aVhumM2QUFxOBo0YzYkOstelFM8tcZumgd0X2DTYnVccb
WuRwnPfZ/wcOMbJmo6D6BYs0mZ7itPHvEVR38Xr9sf4c3+ejwyTUjjRmChQXZH6I
Toy0F+lLPNKBZUdD0WZ4FuQtX6aC/AD3fkfdHkxGZnG0cg4NFkiLf1fFOYin14Sc
e/B/Fredw7aqeR7AAmsDaduRWinY9JHPW6krbv1Lik0j3axAJyWRdBTmJnB35a0W
cOqyMZfXfd7FdS88xCtYPgvknYmnOnMWPDmY6ybKEEN1wihXCRNUXcrbDGRqdELb
dDdLtZUlogh4sObaD32/C8KMaA/88DgqR++Uyd487F5FXS21i5ex0gbbr6Gd9Qq4
62ZAkb+gcRSdRFPDN5FCe4WCQuURheFUd+0xOrDzUiRJVanTZtdIDwrVAFoEycpN
+N0MBeVscqKEJL50cFLH5m7F/NyY/yVCwfG96GXVCTFEXDR5Ny4JV90Az726p4cJ
1V+a3jCCYC+i+lL6ayRvPFrch6QLRdA/Rx07fEp7mPI7M2obct6+enevRUFXrxwy
r607ksVHBfQKJz1XfGBJrVbzMb6uF4PD/h8WzhR8vzaSOMi6LuZ59YqwAyOiNy8x
iWH29oDAIyMWXNkjUwE4Sjbufk7jytzZEb8XiYkogu9gQ8xnLKqnX8+l3O70ubio
0Dvq5l/YjptRkUHB770lrQEAl7Be9CuUu2yRzTIACVlsl2CnfxTsdrGinL2s0ETg
hSUaD+AcVjBxmC31KteoCXl2wGmb2zPgxK8gaalr87E/mNqGafn3C22RvzFcXwla
A4QYS4aIkTOsxwpSnY/klnwuHz+Ru0qCeFlRhUD0Lf8EfujpcQRDum7Zplxv68DY
TcezClu+sEBHxNjZwk8SUXHHizfd83snCtHsHC/z5aa721RbhT9OoNWndeiSZPTK
VC4Buvh80mWsrTkf3r4C9IKaUVwqkNO4TYlryQtU8Qo5byVB/tIUQfY8YLlqFOK1
iUSSJj7tDznQ1oduojdboiGOHQBnEwljdDLEDI7RbRj5XzbKChHCzBt7095jR306
tDau2yB/RaDO6UkkllnS5m8zvx9eJ+j1RxmzCKMI/or9Vz5d/8Atf8AOwFS9PgIx
qhmmUA/N3N2C/VariU8zGJCRR1fFrhPx40sYnMkNJE1X5ZD1H/vqMpdzLUgRq/VJ
79n5bFDWkyi5ATpyvftJorA0QuNJVX6T5S/0GNsYHjVZ21rHdOrJVS9sj59PQZXa
SgLoEnkU/IIVP98ZyB7nrHCfiRYgqppABME74UWLTR+TRy1Wso6NiVqlRoEOXsJi
u+jrOhPPZ3B2p/+1u2nyi1ss+IRWgJIhDXXfpOeTzOTTVQ3WLKUYTBucaHQBVsn6
7xd/Q5KLpNWK/zgtSCJos/35Iyzr/7/s+MCX5hW8sUcLf9y9oKjCk1W/Q5AbJ/zK
+WkA8G+qSIeJDMwgfMYEGfcl8VtCnxWYCO9yRLuLWZ6BuiKT1CgKK0cOy/sIuCu1
BsdXc14Fe/NBWNDO1iNdeNGBC96DTFV8RZkmgvUEtjJbek+tLbin1VV15x1xBepS
lQsQc3Z1ALAqI9XGcEVTpXBSIu7waGLJWtENYlJY2svv5Bd0QIPbp7KZjLtE0+FJ
COaZbpbGOpcSxxMfWQ5eMuriRG0m02vJzsqOO6F76HgQwpWeVApGpin6+mT4nuWj
P+s0oAg3yBJlj9tZWFHHajI5P2BdtAY7Chg1ZtcbkDfvqY2gpZFKocLzIiqhLUvK
wmnYX52mrdnk3gE4tRapWSCfzEU2N/5vrr97uFselcpA9clProh7c9QWZBgBYKTJ
sBIFL8xVtgRScZ6kpqJx9kboYCm6kibsR2XL2r4NKGv5mMz4vOIXdiIpkj/tJ9Gu
xWsVihbcrhLpkxZPC5+jPlvZrmiC14bBgP7RIpHwmK6w1LWiZwhBijbvVdtan278
2pbfy9flGBCUhQPeQpSOjp/if8rSf502Sy8xHcWym5Hv0f1U+cFMi/7aggO5q4Mp
KiYOyUpIMpMzql68lu10NpvvQiecXsQiMc+k9CXlO/NIRazQO+XrIbA/Y0hc6ph1
1ipdKqsouRiRT4eSxQb9LFdZgigcnqEKWlXCraUXxCP8PnoWOoUKeeEL5+gfAUwy
7p+XZOtmv56Mqyi+pGUPRxwIWG8oI3rKMgkmBP7oryLCUlkQJk9kT7tuBQ6dMN51
urPvv1382ukmoB/Qv96jI9vBfSnaPNIBfmAhkU1+BTolCRb/kCAzL8sIBIQxm+uE
lvSCiBqZtNdYdoPER2PZYeigPfTvur8f8/9x8YTYCqRMeOx3fPdL3nRpSp9NpxZJ
/qYnrStso6l2PLt0GlwXQKMb7cTUKnVNTYXLzeMrWUrJzXtF0yaBqOHALSsnehhE
e70WxFQkdiZun+DEcwIN9JcS464TheWsPvapxmyXB1oEgrWnuMeVX5fF4gYRE0XA
I05KrmXT1tQQO2IYuDjbjkVqSKvWoIEQ4mSyn0hRprVTHqPAnVO5goEi7YbvQhE6
Ji0nBgwOTGkqHlNtYmTA1tUd8OxtpbQH1s6y6htv7JVzGBJGA+0DOBEbFF70g4fT
5fKGvVvOx06neUsse+YP10NA2yMa+mvl+S0zuZJhp5Hg52nLOSFWekgV/upfnlSE
+547oLB+6VOC1JdeCAYiuV3IcpBz3Me/uTa0e+rPJ29tJUz5CsFtYHXl8B8rbC6U
holOrwSLs4DL1VMB6ENuSQR4yt+mGAG75mYWa2cwcBecFVMxTn9RbORhOkjDfoKF
IKKodnpi+wE0vMWekccVDU1v2/lKX7bw58U212XZy08tSyftUVrhIQH/FAxTZJ+q
XxL+AjTv6Ss2eCxRPZ6UpedFautV9xwl01bQ/ajIHVRfskCjj/p581B9X4PgXwrx
hxwAjzSo+yD4RLFcbCYb7NbitH8jjxdTlQT4arGSYGFU1h2whz/J2FdRjF406j6M
P+sO8VBBuwIK+Qy72A9Dz03l3c/RcilTI15a/ySEi5Mp/xbDbVmQkE1FmqbsbdyL
YMJZecnUvPGemfr8+UsrCsueRa/P82nzfaUj4GUkhQzgp3Brhb/PtXw32EbKqmbm
5pHAlV39fycDpPcSjHEEEl9NitnE8o5RfLLPNl24MppFBaVchZPVOhDx4zu3MuKI
/lBqRVNpURcAJS0lJ5z53EfS4mYcnvak46X4TBdkyisYOnW/5oT+EuTGkEkNExrn
7dsHu8L+sM6A241ReJJGP8OaTfpJMIsOppmDLzeyjg4eGRBOH7u06vt7pCLsttaW
7oA42PBXMtV7P38AmdsEl0i2DPV3WqOvreu81lXuERqmzW+7OB5O6B+2XfVRlgpZ
dWatzndasnM7GCDuvJdseiZzP+fJ7ShrB3ItNJEkG3uYnbKG/ubGak+MRzjwhWl+
mWsLX/qDC7OFLrGS1Jw0rYyW+uxxxyC1586+xgsyH4RX0eB2lxQtPDQO8mvP2nsI
zCy5TzDBLK/rwP5mplHCfAqo4I8rQeUE0ot6vOJVzGyyXElrBkR6i8NYIF6bG81k
yWNjH+Axy7foy74R6MyAJ/VPWQXJRe70nYkzczka/SCuXO8dEJsnudNBpxDZkIEC
d3jlfqFSuKeODkffkRruT6VsC48fjVqRPDU3xfcMIJE0jhDYMNxP62vL+tpzQJsf
2qN6vQdAMu++btFbkhFeboc2QOc0pQe7JBWpb4qCdvLM6kdAdPjhzNjB1HKO8D2N
QiYE1+OY8biIqH5v2MX/KLzsJ6Dc4pB6mbLe9r4hDVIHo7977+5lITw2XeSUtSzD
qoXyc677yrd503kyw/XsrCwWb+2/Qv6yvN7cv9L8CZBecr3zzo6XcmGi9gTHeygc
z8D41G7NAlH/OV7/aHdji8g/Ltta6/zaTgEhPYDqX9cMLqqgDWlQk74blUeuLW89
KmFY47slSwRr04/YUhw8lzd4I6T37PyzpC3xiUsesAyknkXpejU3pkI6dHEonjOv
3UXyycNPwrJHS+v8hEjn/pxG4b7FI11YgqDuOXjfVglpVo5vQvsKQN+PdXbUsCAH
1p5PImt/c8r9USwf2W9M6Xtas87KirlsRKbF23GAPmeZaUqbVYlxx5WCorUJExPV
L3Ds/plp2CgR40dMvs2bKGVBmVHcbLjsTbx4KGi1M9xqZcvwVy/ATdPm14QCDTP1
0Za8FU4l2kyVVDlfZTqbQEuGARqS//VsqvZy/SxEeXG+O66BliT8wSIiI/9AyNh4
kxsunu0d7MKMkXyOik7XOmj7td3MNUQRUoCkcGin45sDYdXS2KUlFXrPKtDU+jgT
MPAYNjemuT2BOf6E0TFxwol5SVaHdDTIuxIvDT5BRu/uWX68+wR1nHj8B0ccn8JV
4tpNmQfbbIXd25aBUOYNN0lx1Y3Pl1/+Mt4hSq4SqO4NfvZ05h68pIqcR7ZTapMY
x+ncV9j1oJ1CAXfCssNEIfhSjDjGxXp2GacDos9jcMuylXi4z+wsDAi1W8yZCATE
oasstMZrNaXuAHoucyNWx0Yhc8W17t00wU0pEDfSh/tTCHC2inWioh/GPRhslQ3S
blZ7L30MNdsUTVx1Citn2tzHJrrQyc/zHEbNER+qKmCPMnjO5f4EaGy0Pg9z1B/F
Ftm2OvfSuzltmtm7Q4EJhv/lbKRMwUD/kr2vX3EUQCiW5u4fLvvFWynnN0J7LiyN
5tnfOVIw/JDNzlfEj8REiG1A6EBJyuLb3br4EEgyfLdeprC3a9DG5v6uiqeiSgtk
UzM2eN2U5yCZXC5e2Q1ua8zMyeQugW3orXYMl+vX4OuE58m7xdoS1+ncEDHzQfrI
lugB925FCbVFRPfE9n4rxnFJjT3dCKtK/GEkRgQk3eqtvLqP7BopvBlEaNYmYxH/
caaZoRafxHSBDbF0eC3D0OjKJic/fUVKt/7o3BtEJVf2IbZJh6Ah6s1OVhLfPX2M
xQcrH9HAuEpBjyHS7lZ/qSSZQlt8CBETgrJ/SzvlqQ0v0NnHbAzFVmkmsASnf/E4
/yR9pDig+Jfudn66uVvE86nBJMq7uPaDs4FuG5uM39SM7Gi7ahCgkc/5ARFGEyJN
O5VsNlSogPlDkyGMWzbvmbvpKrQXHdBsPTn1eWZ8+WbZMidIUPVrw+DGRSQtVTAb
oXudIsPsTDbyMGr2Jh7EaelwsAkIjgwOGM1rlqnTym+idK/9BTRem13ZkPVJdSjc
sTTol19SliR0BYQ+Ag7zCZbOM1/jGiAxGd9Ha75H1lHwsLGJD72tdEZkq7hGrSly
ko40NaHTEkCpXcv0oxDZ9qdpJbGHmPce8weTyIMmUkprhF0ggDZl/FX3rPFO3Kl4
K5uNopgOwOpNP3Wo0HjFIfkJlSppnHxrzzI03Xk4xlksHDCg1qc8Gzq4piSAl02I
9ErizOSTHnUD+wRfRFuYakIokXAfYPT/MBFs19RhjnxctNilxhNaG8YA6LJOD524
v1UIhEq2xye1kWDN8QeIaetLNeCxyzGd2jk0ziB/Hup3YlttQwWWjKRUvad/rsNM
HHv8pjFmglukA7jWajjBuv3VF4GYywPG12z5/Nz1OMJgE0APsdwY6NlH63pXAVdQ
inMk44w1L1bfp2CNpM3B2RxGvReOS781xPCQKJBL1p6Lf7upsQ4eTF7AzicjldBH
0r012eXtYXSTXwh77/6c9IPToZPjoHYlTsSzMfhXb1HhteKa9m/RVkEl0+/cIJWg
7amJqRFnNXR6CUkwlv99ECGsWfGORl9OBSsYDeW4BpS0FzkPa5FqsiE0avEYOQ5O
m3VALwc1iJ1LKNR5Q1SzENTmnRoQbS7tzOA6b7l69OeRguBnCeB16+vVxMk1fhvV
ddHELU6knlNVPQ94Wu4im/wJOa/X30tPIP+su5Z1GXbY0C+7Q+W3dNYU7Reh7uxT
bmqpNQbYagFR6hZWrx6IO5Hh4UYYiD+OUHIdGgLvzwJr4hbNKs+Zg0+qPrKoh68x
AHSYkkuZy0Ht2pFt87g0uwMrDRBi7r1jaITOp/XrYSfmC4mhwV7IK8huQApmQ8Ef
ATyH1OMcZfoLAKTQFpateYRR+gXzyFP01sdoq5GhMOycHGycKqfx50ldMmlsr1fv
xkzXS66om/dKhEv1vodCr85QGb9d3d2TQ9V6cZFG+6GL+3locfIorKGgLDUoopn1
AaJpNnu1nSL8TU3D9GzN1S9hAtUAcQ33neEzsXmxjb3tjEyO7gZ2aqm/GcHVtIt1
xTopJZ1/VQLfmLnBw8woFWzkWcDvJ4yhohrkTZdQ3T6ZYviVOLLTa+BvOaNjTA0K
YJKJFp8TkUWwl/u5tETTTDCf8/j6V2S85w8m/zLmBW9cq7brMZpHRyC4t84X+Hfg
oW2idQgcvfXs/P5biCxdC7jE3+iHLWad/Mk8fWJUCi5ifH1nqMOdnup8q40n2oaN
HDgB5e7zbLCy/5XVgpIwRk20UtDdsUtpnL8ZcbZUFgZezmEMUm8eybSN/cPLIClg
pvMVRqPwobHA2DQeSMUdPIGfcxEKuPTrVddVfV1oa/pAX7Z8gzg2hIQpYVLZ9v12
V0ghswNaZvlAfMwvcP9jChv1WUQ+1hOYQrDXqjaM6xDx2CQkYANO5FFNU4xwT5kT
KFT4zlWOxy53XHFg3I5JMsbPRYgbi+ChbLddLndpLojdfm1MiCKcb3F3rMC6gnh+
fy3JDumLWpH4q/WunLiKFdaYAcyDAfhFqL4iEXYf8ir7ME40AHm0faEAnKIBu7ux
DCDT5+bccJD4HEoB5F1i093OwO/jBgZhPE2iiWqau6jkP3oPSKEgL9doJnQFX4Cj
A4SH92Zep9KecUbvLGuldfRpLCFqrjePxh3PY5kwSA01dHSwWnb5Xy92O0RckT0G
74rX+DIbphEhW5VGsNNyF5Kd4qy1ZtOODf1JmFH5SZpWymi42P6BbTmz042aapDN
Nkp2XEncT+qQf7gEsieDane85iEHsnI+iFuAtjLSqiMCyS3kLc+T5AXG6ypM5LUx
pbTP9dJiyPIlCAdys7HVqKft/TmUMPsDNBVhbSL+yV289igxWDRcGWjZFtWEW2K9
Na71cZjhmwEvjX6351N8sb1cJfhhZLMsUrclErnkLRuOOYV7kL3YiZlkjMiso7fS
WBsULEcm0lG1z2wuGTBBY4E2vy08Ot9XwgKYnWaDJirFLsBUqofSp3tSrObTIxB+
ACE1gHsvMM7EEg3S7Jw+FzPgflfOcWNcrYKbq6PVviqSRGyHt7fHBeDHyEtfIghq
ZRzidOG6XCBOpS5Spgobz7Keo0mYFEmjIE3K86MKbfbMd0XGl7+kOzy/hug3Wbpd
lnRkQ+suZFDIP/PQqtr2rUGpZcq77Xs180tigbTTg71hfYOWUKKAJrLmpQ0DrpC6
5jWFn/+rdq9AhA0abmGE9BXR0ze7ileSXuaCfsPtS1QqXRfOM8GEJGXslpDJT6Uq
YX4Of9j/cIQB+1dbTzmmhI+Z4R6w5/APIEOlYKQTN6VYSjNUwjE2UrWvKaK1RtXM
AxkZWAmjVJOkjdPBmL1QAC7iei0aYZ9C595IilMrH2O8p7/H0Ow2xOvI5VwHP5ub
AlsuZlbEs1/CHtodXsK9iG0PIS/XJws7qrYT+iRES7cKGnifPVRj3YI5BpQQ9ccQ
WS918cEa+Q9sBPpcFi5Ghzw0cp3KPmEFEeQE31Gz82NBMmm7FuEsZDF9AjJv26oB
N1fTAMdmD9REHLSnpKcVTOZoFc+stBigllfaWuZfYgGKsWD6B7y3LaUcfBOSjhbC
VvuhmHtfzXLO+krJ0id4XfXh2A5bI+X3yh39GkF9XL6IbQ+Ud/fWGrL77GDi5AbX
S7NG2DtLwdomVd0EMsV//IBblOOf6lxKZfG9oRT8G2zk8DIHrqhxdR50TLnsSTw2
IvzVGKxOOJvReXiuuu+C2nlycNzr5rRQayTTVD9iqN27mxGSu+AI3QxSbuBbKTcj
mcKdv+wMwGlqBJqM1RmPilyM0DbVcz8up6HTCA8jranCqOf4i0yxzi/m/fpbiEfr
lcEZhbnHmZVV0Cda4zvMUHlDhPtR4pGUtvu+W/a/MBGj88u+DrocaDPY1iPtKnGh
FuhIuO6/d852Bn86mn7+CD6AY+SWkqLw//GqGqVJ5J6jaGIZRQQgFFikHRtD6lLi
NtLNHB76Aj7MO7fQTgh495jb0Cci4ffCia9QBlRgBQZk5JYIMmWQRm2JGxFH9Cbx
yEllr8v4cDstWRxSXGPWew40v0QidZP33U8blC7WHGyPp55nc/sfnAKaVhnE1Bq3
pgoDsZtrw8t5axjj3vqElwJvGIQ520NouPKXrmS4fyxj6X93TdhOp+0Vlmy93UFo
9gKrXUw8/4NRstiTmdRf6T5DHVm+EiqM6HuohDoxu+GYLhKTG0w0ZkqzLbT3GjeU
AJsgazUNZeqdn4I+uMIojCnyE2HKPqUwpbeBw3NYt6AvHLi+z4ubC5IYEC0ANCGz
s9vpSKdQBBebzLT6epp9ZtLL6XvVlqLEShCtyy9+qX1PMljyzvN7M7aJ0LGJMJKS
ZY5V/RjOm9VInUZr4DedWkkQ1cDBKwNjxwM2fRyS+MWYDPtnWOFPS/i/joolfyZM
MNOzSA24wbuLqbmHKtatzQZmEeDl+krw94w25OXA5nZWO5/IvgLYWc+AwDrghsnW
jIy+l6JGksGk9cqVtcWBvm2O/FQoC/D6sh1zKyKCSsZUMICOcx13CsWbSoHCzBPc
iplm4Pzt9FDL8366eS6y3cyUK71XGtNPp/FMPor18EIhrY2oV7GaJmrlWYseAQaS
L8iYl0eMnWl2EQeeqZKelHj0RPte9xEAgl52B3ePYcofAn/z/yFdWdfPtobOjkw2
1LOdWz5vqNRi39X0gt8mtJCg+jrEFlBkbGBZSfWsw0BbkyQY7dHMOVTxn+A91Irg
GPb+J4GblGLuUSPSX1wcjLpMkbBHiK2yKvI3hP8Xx9EoGT1otyKG4wff7+Z7LvI1
8NWRWYLtt6MjGkVx54WMz7gniCM5njMDDZpLljmjcXWThaTpUiSbUnXi3GoVtwIM
o0FgQEl/SkPjpH8SU634b7l1r1xDQTWRAHZW7c5GHQ1ecAJ2UYCvLEL9kMZIVPLX
y81MJzj2rare/1HwRALxRcLhSJT1K1tFZCxJLPtluNYUJvleUM8ORWFtHauIr4r9
JoHC47Iab/tel6Uf0ctXZ7b0J7DSv4MdJcHKAHJfpdOTibkELAH+aJcB/gCsV1eD
dwU7LB+O4tOSr0oIj/Ekt978r4P5RUyYrINVx4/6rd/IfpR52tB7TRyo7cLWdn2R
j0cGwy1s6Het2+NyCDCao/ydwUZl2kBFuTtmDjN1FHvDGEKrl5e32TLyr4cHwvGn
tXEbC8LZjc4+sJzZR410MXiH/iRTNmXCNgzowCEaT24jrv+Myz9oZlF8Kd316pJt
DkBa7dz/joteOvpz3Ex1CChik9CIGUfoB8aZgx3GeFNFuOrZh1zN4DxpR4yqYa5/
1vMkFWWEXiDMyR8YgsQqa1aCy3bakJtH+4hP+HvazHCMF0edobt7igjBT8+puF6y
zDDZv23n8UHivUKIl0GV0PAJ1R2yj69opArXHvXPf5VBJRIjBFladKhgDKqo9smw
MKZeigTR2vxZfxymwXr1TLmUDVO+gDlUsmlcMELtnRkX45pu8NmRYL1EMwQqF9dc
u5/oMX03HaTRrdIuteeESgJGM3iGT/GcFwpDmwdNHrr/sxpg2ceuU7X5FSayyapb
CumRzJaNgl4JfEkjyNrI6XqxGB6gnbTbgFYuqPaTqX2ex0RiMzBFuGMXrgrhj6NH
VRAqDrh15u5o38jMAUehi5hGgsEVQQcGK7VkvWL09MGz/3ZOxRL8GQd7fAKRmpLf
tKNq4Za679a3fD7LP7gOQTIV6ug2oxJNIPAogDotwGzdV71QEsltvykhzZjTIYXy
saOxE09KF1RMvgtb5R/1PBtRx9UEaApeXyc/PtdezsSx2WW0tApBKcRweJIyz8yt
NKhTBOPiBmrQ0wSrs2yQOeEBo+Slk0L0sgiG8zfJAcauzb/omVw8MrbQi/Fvya4S
WBCOAI9HD7R8rtfi/zh2FF7LPGqqx9ProG52MZzXtb5obYFfkuQoauuIHfP/2tMS
ri2WwSosPSRGhkKEmBJIcaU+tXBArgwRBTFp+GKmIGw9PrXyus4Ui4+mH/ZZjXwS
JNjMSo8kqvHJINv6mN8ITBVcvdm8NYvfQB5iNO4DzCeAZWUoJx4/9YGRDv6zd1+q
rDgLCeh2PYCkwnAJ6CFY6oOdhEABNtjMmKK1SYUo2jP6YVwMGYN17PaVpzo9ulRI
yo0fR5vOwbj5hkmd5IqgUvHqcfKPkpHoVkadui7MTmNWPo8WweGzud8PaPsU9W4g
8maiD2A+UJ1v/71g/SmAjy/iNWzj0zMgDJHDA2V8JOXaFzj63zzk2avcvqIrWMs6
hnMoryXGlHhn6AJ+eWq0lz1Le8lUONICB6QpzVbq3MElye5fE+XkTJzN69l7RLrw
xd5e3wYoRyA2IifmFnGvqtYPbFpLO+gbrzMnN8pK2vYNZd4z+6KLjMw22smZYlPI
g7n19Z7TCJEAngJL6XJyZIcxHFQcxQpR4Vj2MvgTT1UPpXzKpj8jqHWiwATjxRJA
GDDTsSkYE1tI6Y+9ZPDrVR6iBlhECjGoknqGAbkwgOzbNIkOF54mnXELJMU7igQV
wCJUJMfHLnMJtHiYRLTxxPpWxNZsZZRckVM9fJlrVWEc37ipD3e0SZC7kFavh4ES
pprGk7ohWNcupOv4zz+gxJfI8uu3zu+SOUZ5K9UnarRWD4SAfRWDdfYyXRFteneQ
R5ej4QZWKQH9Bjtqyl6g6OngZw3LZjtfptdoRItX1ImwFM3T63VWiuNwovdaDQx2
tIJMkIWwRK5A2NEBIh4gyMSCOmIKH/YxrXFZ5itGpY3OX8SmpC+Knp5UY7D5Uupp
c7POjcWbdSasDIbMZMjsHlhbEbtFBmo0xKMZqrSPVNurMbdnory2/SRmdhqKw0WK
v4BYFZEiyXZBkRmoskxSyyCxAEB2aYpVyfQaek4jx1YOHvBnkhT8Vcp3vmcARls7
nzQzr7KiPu69hvZ3ZIdYPMaIbDm6DtvwZf9TO0+9Nf8ygHifiTDruhNclqinytAG
McYS3wMp5q/lDy04R4FUQd7qM006SbfLLm/rC3//bfITvOHRGtZ9D2hKmb/puHMJ
a1cjw530LOh2Yz7NtsptLZZWl1K3Y01fW6H51LLRSPzQT6Q2hEBfhM56JSLmefsH
1KM5Sb20QXJdCKrKIs2ZR5oemANUMV3++oavLQNX0CCEyRvE2Xy5u9uSN2CUubuk
PYT9CIiuSw4W6E2aCdo+3scrs9nZHXI8zE/OcqcXkqqizwtfoC6r2M9OriGL2dU4
P5PhKYCK5e8nUgRRt1+zqICeLsIYEclXIA8kNgfAjZYX+IWUfbal90JAFpwuTUi5
PHi86QII1g4m/DmTNCg0MXYmSiULfxQuAZ1KNk/cvXWeFVJh/1np2RCGwtATUb/M
KacnNHx6TLw8TbtMTiBe/AiThr/0aBXLjSrYlbd0/yAvWCgNjOJqMYhPH2ZN3i1u
JKi7du+znHNo550qaPXUkD+qUERvWLgG7B0ooDI4Jlxgpjo15b/9rZPpr7rQt0P1
fIgwwH7gUVENabNy4jq9toA4LrzbE7SSYw+1wUhC3wr36399yhwvQZCL8z/zo+Tv
sxNW4bDSatRWnUi13gRzoR4fLP4zKNwXIRZ7Pf6RJv/r39e1o7CbUQR7VnPFrDBW
qm92cjHJ1iR7HyN89YrlR99XX7E5LybmnM73u3N71Q5+Nm3cLB11uQnpCPGoUhyX
KdvDbjck7yt/OLnWIz9aLrLnrdagFBktlY3m/CCr9pVr2HDvgJ+/JnmpQJZ5WMGS
guPJWMFn+JmdZEbSHAqpUQhWozQNyNC5z32eIZ30SsMnrt+XcpWPjl7Aer4N0vOa
4O3cjIYQxZPbAAxCo41hfKFsuaaPaXDpN2MaxQJEXaVrg/2HmtfGTysdqNB5FaoV
LdFNAO0HLOTUQAAWOgyg2zBAptrNZo2psVkSV3EucfrK8jl7QSHYTD2ysr5Wc/Ki
ruJ2nAzmaZUdsr3APTYfQiiK7IwRWFK4bYHYbAcYsAvct8PNBmaJnm2wB2Phikx9
VDsm1MEUsua8peHkcSGl8C7mUXysIa2iBm7xXuW9wmccVwkyCrf8GaEcUsr+UlzV
aGfVjdDbQ8e3hoqkSVm06o1PiqRypI0Z9hqMe1KZdzJr1c3RXqgt08X6r/RP9kUr
FhjEi1zC2mZ/g4riXZSYSEJTZscf2pKZH9TTCGBuAna1TGun/k42KdVxKuXc3i37
AREKs4w5OyGj8l2KMq7HXcghI6dSmnycGvA7PQddnlkaxgEJXLkszgHpHtPhD7c/
ls1aafZwys6r8Ai2CUa8766KwgIahJj+MPwlbrSpha2lWL1an4IVZXCRMbTTOXQx
XRZ+0up5IfGQPBGzyaDNDtM6AQiDF0x1KUdgDZpFaPr8tb19xfZ2CMJsWlMh/gxg
MUVibbXHpaoM4D7k+roCElCP3Ih9T3EwQVWT2UUQIh5Qj+hosutQFDTWe9RekOT4
kNXzMS6zWz3dBOUVEgeUFf3Ygt19bwizLhPG1fOuH5k6+zP5O3ZEHyoLS+THjtOy
S6eyKA0BiwwvNL0z3oWdhVLeNsJpkP/pIcL+iRVuGDcLczTWeGQ2svBwB0TmFOqw
yeuDBYqQdnkUGPHnlHMMQ+OIZyfuzQNh6N873zXhQT5dOVjFUOLjk6PA2itE0wGs
Msx8KosT4k9U7J0gA7ITnrspgpZOEYMvsVxT2ZPELsnudhkL8FxySKpHOHKssJfH
OJ5rofGUl8jP13NWPlIc+DmAuZCquPjygOqVQcwpH7JkrejLq5yNilliBsIIoVK4
0ORWlBy4UtSpcdKntK9cECfgBiYLsnadn66LRB28tPhsvnnMG/SqMDn7WAG2Z8U0
z/suv6AdICnjv3SDuw/QC846FZUWezJQUOhq4vnZHmfSBeLO0anbH3yZ5yoX3wNJ
q4CdFwArOe9OgOPPlVPe9w9PDGAa6iaLNFn8pzDbziWK6GGCiAQlNlGMxzVVhJBN
mSgvOGAeIambq9e+4D090F1r1VBFy2hWYmRg4INp3vNb+3l8iIrL386CyjfPGw8P
L0Y7OQSNtJO9hSwLUN9lkDLEodQmtqZnvjXZK5rM7A6509PHJH+m9N2cA27RpD84
6lB4GXlSmtf1zykr5CrQMS42FN7AfCCND5gK71UUWXp1BjfXnyGn4VkCcwb6upsn
tB4PkyO4MY8kr0JpfMRR1yRV5Y9hpWq1Kryp9OY7luHH7zhNzVROZhZuifFWHyxE
PWc7qulgqT0KeSY0UO25V4fhJ3Cj71W7jHbl8OWVGuJvZaddheG+Tn/dOTTvVvyK
/crA5J14v2xUDFxecviPMOrbl4HxDbK8nSIrxGu4+K/8YSmLvrWok8D9GMwinR0t
Q/Cif165kuio4b19F1zZZR0MsjBRvlfokgk8GejFCZFR6AU8QKrlZhinS9Ij0ow5
6bm72PgXU7gBVB/g6UY4QEU8y09yTk1lj9zkjoo6lYc+8teXonNTl4MXXdN/kYmE
yHFnK9vGdHufc6sIa9S4IJMKhbAedZFgLHANkuNZ7DpwoP+EFc1s9Xd6OitD/Lr0
ePVaVrp0qdTCLjlZMlZTg1QlTW+k8xX1Ydf2bnaLCAWNup/SnJgBif8s8z/jbFYz
CinQ/N7PVh79hQUOsc9rJ25CjQZkxlo4RWHWq/AxW7nQafXGdnBwuuHxKotkV+bN
Aq4ZenaGqyFHRP7ok2xSD1xmyfxWG8DL1kI2ugKHUYB5RkTK8J9gDUVIGtF6qRWv
VajwcsSABeOWlzyPlpjeXEoek2Cb0Iq8qVl9bQbjYcsRqyxfT9tgeah3bg1/IdYU
Sicl5lTbFbHcnJvDVpt9XJfVZSU1hX+3ulx2aQ1OSaP8YQf//T+Lc0F+x0mxxzay
V0PK7sV2ZJ8ZsPQ6JlhTptaK6ZEr1CH/CmNt0f7zRSk2TViLLKGMTCjnLCAKvEf6
hIPXZVyNm94mJyfWtZMnou6IqfI/j4hMjWDzHBKub0eqFMb09Rem63blw0nFRtHh
D8wKWsdT1flo9SZAfYh4/LZVmtDqAT80C2YDgVYqF71y5edfH0ISJ1ppNb9YhQ+D
zxyOhWQkLu+b3BxfpPaM5kIRtaa6S5HermHQ5IWkWYzyy6In6p0Kar7VR6RFd7GT
fkK0uVX92gzQgmt3NCL4w323IBrGGbcch0HJxode1pu+i8XAG1WDQdG47KXoeWeH
+Qo6Rf4LQcqb5q3dwho1vdmick1cLtvrqCBYcuswNbE9pl6Cf4yoCBb1apGC9YEj
TwZJtmjMAa1pv8pOkzM1jBASYJ9HvO1AYd7dZuswGQxvLQvIUfxd6oFkYjBziTBs
kJaVj7GpRZPfz3hFm9Eiyr/l3Si2ckgtKWf3mL2BKlfsN4cADgAXKPC1F5yRBNlS
heEEuYwtsG5fzfGV/cNr8I5RKKNlMlZg8eJuTTrDk/nvGq1giJNguPBelqYMR8d7
EBKOEQllDGwqLK27OqoUUzQmoT1Ylq9nOZlUhUBOmbUt4SdlPOC1gHU/kp03ZF+Y
lRZjyrZBU9iV55zP92ChttiPy5pfmAjD+UlSjd04PwEqWyFiFFEOXemqMeHsC2SP
qtJb1eSkfdImIK1NzR3fGdc1ZLkuAkfc48GxqMohtZROsErm+DMD4zU+mP9lz2oV
HL49mqT20+dW68W3n5aYPmQ+czoHqd82lOkOVWUAoLHxrB/JnyrWHpN1Lxep4VkO
yEWgx99oMkKJJwoHBYkQkDBo+bpLQWqbegWAdlJPIBac0qY0vcMaUb7A6JGinXcB
ZCZKuHafq+uSWxHCqeOr2/RnGqz1DrB1zX3HQf/i060zYb3g9bzEmVzD8DhlLq9C
VApvMAWcngN3Q0V9rNlCFkl1pWT0csiPB1zhir5V2mjG+oZZfLBMbQJLAycw85yb
u3BEJBIinp2qxvW7KWIukAuMAht2iuCLBiC/u2xyKoGjVX6StQ7FmpIe0vz5oyHj
RzezZc62G7NramZSVvHNK4vLu/wWZGGQUyGFQw5wBJwN7t9QD9qMXwZYn0nM1OhT
rfSG8YU1vjfgw3KU9DS261Y7uTNC0N2DniGZxUZW9tatZuVxEvTlSGh2EXjBaNe0
gSk6H0spJxl7B3ft2t3PX4hqCG/LcT4Gvopz0idOS6XiKRCuLfSNbL3DCAXEBy8n
e8t6eq8IWXRRVqM3R3Z3/I/Vn5B2jyuFKDI2JieEr7K38xjfKrV6no9hbJY40i+X
tBQojddizhROEsqMSImKXkh85Gni1QmGr1DcELSeTaZml1Njf5RuxNuxK4G2X6dc
O1mU6msrH6cVTIJeZOS+LxoqI/UJpYblGJ3yPde14Qk+fVIbx2AS2n5X/3MaghxD
6yXyn+7f3PNf9Wa48Twuu0DGYnIIZcGpdC3yU/zNNd9FNdUkbUbFwthAN+7VGDbc
C1lYj9IvIoTImcHoBL+gMZipMLEs55ToIUrq+DiP/dprRgUUPdDZUgHB84SrVuN0
0ZqvTgRU0a2CgEZMJHs4cV+oB/wgkzd+5b+4FvtmUWwFYu9iK/Od9a8WpmGpKpMl
5ZMy6A5haaBV1EgQxLhVtAxGadzxoPI/mAeYLHqXjDvOkhwDRMrLtlDZEE893g4V
lk/O0lRudWKJ2T+04CtEGReR63Rbd1auEfyRWv7X9qc81RC1ccLTD3bHtGNvJW4/
jyVmd3drFpqxmKxh/GE0PswBENTJp08oED+Q6tEEi3Fl6pNIdPU7xf04SdyqARx6
wqSctHsfjQVV5rSoR+r7Y8L+pXjwsRnDzSy+NdYpJMkQSRepYOu/bMLTdo8s11gu
2cB6N6hxEgcc0wlyNRriKWq2MvY4NLpenh8IS78soEDiuZFcyA7eiRfTuJmCRM5A
/mUuzJ+idGS0WA30Va7+Yrq36jyAlQ5QGzrOGQHKCB0XlcH/Oc5c86Ku1Tt8D+sZ
imJoZFZHvIOCbAh81/qgqzACj3ltEyfHCQnb4Rr5IPtIdhka2yW2izYzcpRPbq86
kCxY+DgU4kt3HH79JZ7opPjPWcGy+NrUjDGjMet4wZZRI1IUz1DOxRZ8yKaDE6S7
PqUY489hLahlGoZX5gSmbL18b6vGSjv/iahjxjfTyV1u81400pTFl4MFQ37ibYWg
CzFR3iRgDxv9/6SOowy27LKHKbQmdBJzxx5mT6tyYo+n7e+n3kwrtUr77XEhyABk
jRTXkv7rrRVR6wpPd0H1SwfFyznMwLoUpnILEbBezh4HP+5DeymBr+UKKEtyEG7v
anJM9ZuSzsSzQn7Z1k84txs39jV5OG1Zhz8/Jy/GGOo2xahN5Iao34Ukuy6kytAr
ZoXDz6LgEVUq8/bItGyS7foz82fFUEmD72isVCaESNr4bqN19JeuP/ImzDgN7EmX
nRiA1Pj5SDX6piM8HQ94R56vjj9ZXphgn5UTSZwK+Mw2CLvFia1oozzlF4VD1tw6
fdcL7qe0C3PuSGe77n76mIUCHz9zHzP+Gh/1j0KwitVU3zHY26FFd3LjvrZt3qw0
hfNjuAYZS9sh37aKUMq+XFg2DLBz9bCSA9mmYndrUvFoOxhHUICxcQ3x6Cp3gUoo
d4L48eI1ukfg4EAOhfIjpruRoWlex85H2S3LbSpQjtrS3NfIqH6f71YFpEqGEkYd
2rcoJJFzTh8y4Xmb6tkPhEGk412MalJiBftb9HRMbM/J//euHSh0HfIHg8UzySIA
PewZe4pPOv28sqFzXVv9jsBoXaayXohSsgSIaIeS9mYzNm9oyFWikPcZgfEdIDbu
Z6m5b/DsF0ZOvLne7mcS62Fx5YYfoVLGbKBfUXgq4rfUbxn+ZWWxbi5WxtbVP1uk
RRQDbww5RyxbSQsB5ue3xgB4pqIfTM78vRsvvLttWFtRHX972HEbJ9t9sEujgQIO
pRg74q5TgCbu6d2PqFxkhmYG73NXSqKwp+cU13xZK3w/C8Q/na+yHfufWKTf0zKG
PEdPeBBme447NvuPbsL6nH/4dnkql2fEoe1HiQz0EdVoND0SZTfQto9y9V6fDSR7
/TVuCdvLRI3H2J7d2W8ijKB9//zSoMsVgbz8imkqZV+ckrzWe42jPVELdQxS7ns1
mNqwPvJnnQ0z430ketUezqMI0KBOCOl7qkv5ioj+OsAhd6xuEC3PBtEWh6W2kVcM
nki1pfQY3AUKLlQK6yQOp5xUJpbS/TtdHASKqeJRdBCX4DJUzcZNLNzn28Nb7OGT
mH21dCp+LFHcUFF4CCRRdtXqS2JxXkIFRD5K+OHElKto40viVmHOJyF8wvzqynqR
75u/9DYGZxCVbz3MANdQsWVZpMr5UfYpymNg55QGenAw/Iz9w5zEkwmNhAL9MSHb
hq47PaCR3wCLCq0UytOo7+YaqEf3rDjMz0O1DsKIYTWyM3Id6PVr0Mi+UPlTgvGp
gC9cq6ULMoFLBKIvv8JZHPb1EngASbt38L9bWoEAK77uP97iKLr2JdDFqe0j/R4P
bEOeUlAt21/24/fY5KEmjy3U5TEA2C0WZbAEeyf0TH1WJg67F6/4fhZgSXxLm12D
twh3rLaSe863nFxfCHcn8obEZfptkXUHQD6FkC1pEobz5wPnGWQ45VH5EqHGBoaV
9A6stbJdPixhwTrk3mtYovB8tWqq2f1b1h8yRpkrZ6ju9AVQgZEtY3Bns3FeYCB3
W2kIVJ4oIFUTkxUh3HdPh9u7aPJbpYu5O5B00oPHxRHA7E7Fr/exrPfvxWv1lF+T
ZMF33SPUBAAGNw+8A6ag5sBprUaNHfk36S7kqn4+Ygn2gODjWE96pLLmmQvIFLTF
4/tcatEnsJ3shkVBBtTzItf/YnqODvPZB3bjXWJwbvf75H1Ypl2JP/u1PWiZo8Ro
kwdm4SXnyYWYBYx9c6OKSocY2MvISp7xaDvUs3ONoagEZKMsq4ZuvWBXyh7Xx7gf
+/O1H5PM6uYdN00TXy5JlAxolxkWttV/y1JPZHgksMt5/Zu+PsAjYNq07tNbH6Qh
Us0nto6SQz30HOp0/Es1CSs1/pIRUxg7fFuX1UKPS3PoTrIO9cIVW+qQenK7OTdd
njHz8syymrgKIg0yeNr+vtCNFxt4ogOt88yJ+FxbX6hxjgMdQ1XxG2QBwyB7K/jN
iXSM2DtrYMC3tg1563EePi6LpW0FdFVttbHkXNY0HeMOJpxtZclqMdV+SCtINtxR
oMAWm1OimwX6Ot3MDAgB7j66Ac5AT8nGD2/YTmbjR3q71BKai9E/gUSJUxwPRTCn
PQpm5t6ImfOInHfl9DKWoJE8Nrc8R60vfC738bpdkXETQ5s4HM0iRzF3AGLI9To5
ACThxjOzVeOFDj4c4ImapGeBOCCJHret2roogaqvI0BfCVxW79YzdjG0R2mIzdBH
4uyAyXinDeu8jgYblBYa/terKKvofOvPk9/0z2KbJQ0mdlfe1qFgRBM/Z46f481y
XPWelTawpY4O8n04TiaBsiU6X9O/ruk9Ax+9/uvTFj4Mpp3fYvWYNe3gWkhahsbi
2ISaFzsNZjDboR0feM9uUn0yho/MrFsQ7YyeWtxZWMfQqpdp2AEo2cW1pCjPvAzz
CX4aiRaJSVBOwGvjCmBSGSxQcKwJbWs0EIyV0YUIymBnRy9fbiaD+dOeXl5ejrQP
2uLdYRtd8ccXfu9fRy0kgSXjFiSylh8nD1c6j6YFrD8yZGMhqkMcbyx0lDriwXCW
FmDh7WDHZzQGJCdFWuT0NjWxQan8IG0ORhrxTbrECwx3fnF1BATMmtQKHHzjxbyQ
DgGdBkXpAZhmdmTiXqJTDBKQL0wtVLKnObY6PDwZnT9/VR4BbwqIy1RlezoO56WO
3xSFqOUl7SaswI7LdwkorIu0WZCaM+FcpEbRrNY7RDVNtMGkOioIMo/xBBiAyrAL
YJfDN+AQOdjL2xipP463JFYEBpVB+wLGdbyGCjyPHOleGbiz3dXAi9VPaKcnczUE
UFHzRHcAU5SE+gBBMvF4d156OTLFxSNuRTtf1+morQuVYRDRX6t9mGOySGXtaQa0
dOu+zAe0RyP/IkPEhDklApzHrzZautDxGX8PB11lY2r0FuqjAk4PisYm8L1Cgvw6
/N0Bf0iQU/CgB0lp5DvHxbP2N8N30RTSCNR+ghkARnbgnuVGLk+2lI7+IcmEGUYD
UQ8wYoOikG6kvr3cqlND/XSi+PxaAmLfiGyA7eb18IsWsYDQ5gxH0v70vZgArK9y
XSU5jIRfrdKllvFQpEyi9Aqx0EHstwLGRu7SFKMzBWfc7vWvIKff4PRd70vJ1xvT
SCsoaWY9hjbXUhwUxW1eeWeIffUNAcaxBzfzA7hPWTJmq92ZMmycjXIQS0rRv3Ia
1k6Y+cXhytopnf20Gf3rTsxMrwrGrRrCDeqEWJ9vvW5vAS18DD7BaxeRcOYbI744
8CDdmqE4euE36NzIMPLXIzg3a/6AwF/Mnup7l5zwFq2kdSceYBJpPeR9x+AYlPTY
aq/Aw3TLSE+sERatmiygJ8FMaTE2gRaM00KzF8iFjXPcE6pju33svlC9oANT+tNN
AaV8hPg+mFTyHl+X6C3mHpfHeuRYvrxFP+/+Sb0nEhE9sc5890EwuOyQka8a1KhT
a6zkyMPa+ea5jJtKT1OaOBgvoJldNrMkcprWvRb4eoIpz1QSNwQ6e40i0psbKWlC
+AionEWOc4U9T67s8d8nBdBrfO3e6gXaWmSeX5kPkvCjjlx45wWFdCCxwIJ2xNS6
dX4w619Qj2am/ez9Fw7RLJUsvyVgXjvmOymMcbCcB01dkAtJVyIMTsUR2Y7IJ5OH
v1I0SHvrF+NqUJAgWO7etUuuBSSfFC3ZLcuqqU1Q1b01dnNukKNJ1QOtRfUSdt/k
njGCytahxgk9pJoi0uf4YHQh63DNrA9TeGynlynNgZTnszVXUMoDhC/zpwTcMhQr
coVTrHI39Qoo2NrgjOOvernidaP6eLY3TiTVUhRgsEiGsxxJ+uiujhbFCXuLyPSj
WXbacjagLRAAyQ2b9wpKCR6I2MJqSbqTMZSebb1zUTjcrDooCyH2nKowQ6YIw5uy
YnlbAMAmQ/AWC4SuFEc2ISbAu7FkmlBbzneL0Qe4mMHUJh+aLpFZkRO0YsDX+nIG
TILdl3NZCtWE8w5cZfjdfUa/fHGoyDsV/npeWVLIKOwqgrDDsyAMsC+OeAwXpaYq
NhyqUOzwBCa7kT3pBiH+IPTWl3ToYnDUR2rmz/XyawWJc/OWAPhxXHVl2520ennW
kVOISbNRt87xrEpyJdj1qrOsAbBjag8JaFcEZ16hDLMYHEtKgJYmy9Yh2xQa0YDT
nDdTdq49+YjU4r5YiTFdJ9NV47RbiMAqRRuDYBrupGe+Y6ls05uRMZKPljOIVhBY
2Pb08kiI0jv99zlgHokyAL2JmxdZrZmp4IckJEjH7S/Itq/eUzS74vRq4EdTUU1z
5ch/38J0gJiD+Blyi8FVH5ZUvKIGYwWCdvJ44XZ7p0fMYOhq20p390jgBsMboHfq
Ku3BWep2Kr7WI2wPapdfrXD//ygUoJpCTrk+GYWDllUcXIPsSOP3r1/F7jSzMiG/
bQPhoQICN1PZgItr2eql1vKPtTHXwJojK+zRM/78m5iep09DXw/JhAYl2bDP1YgZ
yrg+zSstOV1qU6uILj4mDPjUKtZEBIdR8M0ppuEYS0vm+H36uTTj0qNMukC2JSkE
+YdP1pe7j7X/rGea6JxyD/wjJxDy/SpnpTEcROd6Jc3YMz67KwULbdORELb4HMdc
Dan6cxRbiPYm3F4LnAJN3h4YEdHEMdp3pZUZijN7WvBOpTsEvTk6coH5idnpxuDs
7ErT4dpzDM0t0aIpEUIQBEaCztjmFcKJaq/MnziNih1gXuphAKnMCTJtGgi09KT7
mG6OpUDGkeW14F2aOjJwaI5Gh5GfO0rdlm1rSkK7JdNimcrLxq4WmF7Xu1aM4+DH
QUkwDkE8RMml1WVe9uIVUa0id8BM4j8UxHx3CGpRI83/sVVN72yJX92rYo72jR0U
nTNfVh8x3yz3mWbd8lGKoHnpgiOjhKn2PD9oFlD3VOxzZbwGpGwie40fhdEUDvmU
dyxge1YQbQXr30DtKNk8OWsU0M97XMCiIuABjjxpCWRL9v/weysuwkIcolpZF9DH
QpZdfu5LOk3DLijBh3m503ogbR+EKnMcj7QST9NbC34CZVJGH63pyEZlyLjhMYnU
iqIbS5CPOnj74TpBx7GW2DgdVFIuLzCT7eHabB6p5yg+UNxc7IlwRhvWMs/6UwT7
hmw9nemlB0bMh9pzg/iB2LGwdykHRv63l5/yw3AuRLqRmTnaBKqy7HubS20siOFq
0sA0K6K4FU3XldnTO9xxNPRhzZVfGvybbgW47zFzGJfuhZQfspiM8nkBXy7m/lnV
/LUiboD5DpCwQ7p3MbL+/U33HZlzzZgov7Tc/yTKsgaKopSWT8rVUNwMiEizI7cK
2jOLfWAXRcrGDZPaxHvbHfe/n/KToPo9ibacFmC3D+fnwvvZ0xlyq6Olrd4+ZLtI
ow0SkL5Yd7qB4q/zTMcyMktWstNAuMKY6TI1Vnf72e0C1v8DP+qLfH5JTLhwi29w
Ca7Kg74pDAWfl7oiFjT25IGbk6znTTEvktKie9BsI4aBb3U/PqYGXqnHdPVBhsOv
jeNTAjOLvQul82gL5NIQa4dPeGy6PbkSiERCes2UdK3Cts+U/gJ5EoW5bY/7Cn/s
lFvyZ61RPwerByFam0HCVUCKVDp0ZiSpu/JvjGUSGQPaoS+rWDhgIKdGZAzQ1tvy
otawrSbJXERmx7VCsXk2mF+UNdpKivPbTJAX80X927uxTV70LAGbaCDT9mzELgvw
/DJMs2U8drpUckJfZgLrPZHC7Pp9kM8iA6m4mBKF1Ymyga6zhnXzWytMrE53k+x8
mUv772L7TOjZVE9VcFQA2CXRX99UMQEUBIjzRYpV86sQYzaFz3VnDzq3P2C65At2
PHMU5HgNh60UQnzj0OA4uw8OGkjuGg/yYE/MsFqF12HCCGz2dIlk9ESHSmR4hISi
decDQ1tC/pNSAiygEMbiKidTmkL0vPH3sz0fkvwRR/RK/gFnLFrH+ALBZds7dMoE
Ps/xcTiF0iWerA7jL3LG31zU45Ep4Y38fnqhivsDxWxMvOhJTf+/BqPnIkFv1YH+
96WY+NeBo2swDsMq3pl0nfEmd/GAu626F25lzzOA97KQGBHan72QErMKCBki1mB3
nXzi4LlUSXx9sS+4y3LUPRlYskVbHR+ZcId9rBdBZqwDDOB34B8AskgDiY2woa8N
WVgk9X0R96LhFu0VqpbKtAp4px3ThRXMbhE6Mj1F/TVBl1f50uuUXKKjtTKETGFY
+rPPxInMIkc/YeUgJj/dyR4uuiYq3zB0lKh0yA61G3R0Yx3xgl3ZoWRYhTOEx0hC
A5M7zpfQPy+cvt8WYRi7AdEW9zvTQyTZHw57zqx2TZ7OQ2/RfsT8mR+L7EWdy8x8
kWktD036wDbHpV/aI1GQlDY56Xu7gAtyhtaezcdZDNSg/rIHlCDv09c9UQ36x7qd
iWqO4iA1fxz6FH3l1dQmwHOtC7fXkgt1cIT2hUsLFxqJ8bQ98xB6sI26Tl0JHJcD
/6ByKzxRfg1OsnrDKrOrBOW5C2trEsi+2XNmsVmMvv+bauyNPwT9iUiH3HPcxN9+
ososVxSam0mJTqGhBSqSdwCpQ9JppA2qZWdJ081k8ItxxErSFCjKWWtPgeeCbP5o
Pv9fMGrlf5MzuPS2vLVicRHzWqL/thmz66q6jfOF91l207+FaK7OlIkuer0cLLh/
M/JNB/Fr6XaiKCCBV7Ko2jx0OVceZELbt2OIxLwsGE0w96yu+NdtKFqnL488I2oK
qSxNROhvwSR0PkrNkyv+7TyyhYEaSB2OGcRlkiywCAGzdmXNBrBrayPejs2UDy/p
SPSx2lRR56pWY7EQ6qQs6tspjopZckcsNVa50EpWS2jkypa4nNa/dEMpbcGq8UTr
0PykN7BrOsHPCQ7upHw2Ktn82u9GKK3JBSfR+xO6YeY9dBywrWOBeUzFd6Fd55tB
wplRd4cE0b7GkqvydT6mjbqjajYDtHxIhfU13fK+oTw66FxEvjAuPEZsWxO5u3uq
A3gEJsMfVcj0B1z+WL5Gtxnp6tOzdg8gtkSSk1oP25/cuaCVjG9Dc3udtqTdQq5J
Qz9CcDBgLCk3O0ggZ1HIL7DqLT4rccl7GrLV+5tmJmkYczo89S0r9beS3GQY6MUl
QizyiccXf7xUdv6ga0i5035epSj72ERRkf/q2NlJKk6/yE7QZvZy5sEfwAX9hz0+
ExkiBxZh+fcvqbrql89L+NVBfI+bKXwTELekfr/rh0HBOKDVMoU5AF/qdn5x5uK6
54XsYh+wc4BhqAA+mXRlf6TLKJH6KXD+g93JoU8UKfR6j+HYAJaNKMQsJUF2+Mab
geArWBqtE9D6zuZPrXWtMf5VIrCIhY8oaJIV7z6UjyE7nrzg0VkvJETP6mr4MrLr
/QpgHMujrjqWMTwbpi6HC7vkzEh3cCnuy2eioy7dkIe+wVOCfitTc0pNdkwiHqU+
/RamfNh39lQ4AAL2UzLKI74Ivtujbk4B/mINvW2mc7A9iOqgdyllaIVS34jjjOx2
gXhy9n17l67t94WW/bz2MRF4nuxIaEtwHnjFSdTBQOvpU5ZreGbREjlURQv3uoXf
W7jdBJs3h1wnWr+v/5hrcd5Fs7vMY0z26E/BEVCKrjBNhQTpgOPg/QjB8y1O765m
hic+fLs3Sz4/zrbpNyr0e0OLVScSRY45MvYY1hww71DdGBxvQTOkqVqJfKV9u9N3
udvxpDh0+14JokdpDJc8deru+u3cLWWUpOCrJWE/oB0yEqJOxiMd/hQqxtfCN5fA
cmpNtJaSuVUb1miX3zAcp0earVqC6pPQ3Z3PE85i0k9z+jc5ys0iG/A8KFktWDBc
p/OWCPJUhzke9rrL9++h4T5w4+sguOb5g/a2jmqBtZN/D8UYP+W6wrOji055ld1u
b5w/yL6wtiy2Oqmp2Eal87VhgVW5v9Fc0d0PLML5Fg76CSD/jAOFMXVrbkAGFIQ3
VtUCbd8TSUA5rc26+PQ4h/BJbrfoRb+g5mCjMV4D7Uvs42FPxNlDlC12V1uavDam
ULPyeAon9Dh85/SUbZLW6Ifa3LnJhO+X+tjqSEV8XxStSLG4heuZV2jZmlaRAH8x
OlzfaG6MuZa355pgIyaYWa75CJXmZ8GUF0qsihtnbUhq2JzUkZTCLwxsmQPiqnOF
BYh/hIMTb4M9UWR0vd1cS63PoPCUY0SBdz8U+Hsiz7j+12y2tZp4BObGNGQTHxLZ
xEwrhQjWmX0pj0B+XqX0N5HP77FdLsJe9Bn6CWFSQeTpBVU0/VmjaDpzfB/upc6n
bnSD8wLYGxQC3qzdPgs+RfRQLHEc5RxiNBpBGLMPYnCYNCN+blMoUEeDedrMhydX
Ic7kWqTfacRq4AohrqKVHJ+hdqjJuXpmaBZLmrD6X+r54fTf5gDZ2UP5VCfjvWRM
5toHqTacf45qf5W00PYYrudRRR/08dbB42tjdCu04gTyDIF8LNFafJFHvZOaMxgX
ccvmFaOUx67fuaX8f3BRAxADb+mCyUOx7YfaWDgM4px6rpO7gwR9p8Ob5Yau8MIy
ShuuY2ZzCC6DbVvJku6GZ/lB6JTA7aTJV3yIH+pWobiWjVjiU8fFL6xMZM4i2RcD
gd2U2xIGaiC/kZ++wtDl4wvUfoVW20b38rhOILmONOP8ta7NNZa1HVHTYdjRdodS
yv4ZfWiMDSV/S4ihR9qIebN1nccF6Q4QL2R8szQxwj8eLQ4TyI6iL3M/KmMmt0KA
D6lWygYGCR4txlHrIbVGFP/blX7LC2CPtUumPS91/L5Vz2uliP7FaQnAPYoO1Sk/
Pj8hNcImzS9JGruejVmqT3oIv9hCjV3BXMVCcveFcb/XsJJsUI9gpJKJSNwksYsQ
hkJC3qx6xYxvrZsQ0hNsouYj/PYVMT7H5xjb9S0DrA2Xl9JOx8WP5iQGsU8gjkLP
N52EyJg2pMtcP2NaUbyF8GaCj67LUpI/d9QT4kyRDLp9yxDRO4IdZP/96OULd4rL
vYd2tLygZ0lN9oC/lhe9YTujFMxSYH2hBerg6HpohtMlbOluyeMJVM/vBUNBnVMT
1IEIaaMI4/gtfKDGxTRld/1j3+EX/S1xdipTN2rCPft3IyaqEyWfHlt6WdFJ1LoG
8TQLECjlkgVF680iPd/Wyh9ECgforfkOVktb6HFgR+FeHiytz0P12nTxWBccrggn
+4OpU2Cv2OJcmBT3OmU7DvZ7OSiRAn5rrQWCtHgVBKIU8fEB41YC9jC7Z3AtI0Jr
ToUB0xXQXdH2VCLeDm546CRUR4KqmcaKu5kcN3j1BGH1OFo1tRYwipSghQiLKoiH
HlhowpugyBm61q5g/rtVxbzE4J0l9/LOCZt7Gu9Yftx/MYP6OBJS0ClIurGyMsdQ
JGooWBwSbl37MXRzJkmptg+40pPxZ16HkPx6JzYyLTWeBcTZnMsnSsZ9GHi3eti+
cKqWI6XxW49oc5iTuQAhaoJpJp4AtlxURALkIE4Ox6x0P7T6SYNl0bHiay8Qq6b0
leHJraexjTuFyVKqyAm8fud4InMXSAVfIdQcrVcMqT5llJuSSVwQdnR8KsRN638z
XqJYH2dCVSVgLAimOnDQs5he5qQAxuxjcHuoqEsUuMabIWK2Kb9P4Paw0G5iD8Fy
JAWq3DeiuNJ/F/9+M8Ys3q/ZcPEwrB28Xv13JlH3mtEhSiasGZx7asDlH+HAHdgO
+a7mZlX4Z8ZGi1aumddOWh5+LDy1h7Z/+yTsMKFQInyQwqmcVdfhz5A1bQ1FNDG3
uj3q4KTgKOvCwa346E6KCqMtKFKJbIDrGx7IZTIuGvWxydkGl/oY41z/mF2bqZVB
pnucmTW7ILboiEproLUdgzA5mUkBEerZ3dPO5tPqquzugZJgkpIjV9t68N5VjsmM
qWmOJRRJukBH0KhvWpNKc8yXdM6NyszR0Lq9a1cjUE8T4v7vXoaRwDkisrBm0EPb
ecW0ICr+nC8Vol4ecIfC6UC4hbtxSO41NMWOqNl/u9Cl0gr2ouJWPVdmprAXjhEz
zXqV00Seg9G01/rN8dfmRRNp1PbeJsQs62zypy1KALEzKjbKof8M7aq/B79tSxeW
yjoozpGoezJAo4Wk05zq2iYkkIEAb2kIglmxPIIGnj9JrJw3Ci39xGWeaiVzV8o7
Hrj5iORLXuwkMkmcacqbsoNXqUVXv9jz9gPJnQEX3AzhoKFEh3TcR9rtr/Y6oQ7k
jgMViy4UCTOOHKY2K8xoNBedF3fDB7rIbdQbinmIYui4pA/Rf3haGiQlGiRi5+8i
XYOFriw/oHpQayCYDDxMaZcxJeVgZv2VgVjByNXm6GT4/j90XnP1AO6bg9HBx4LJ
3kgbAeO9P818/E9Lvp+KulzNQS9/Nt4CXmE7wPv15xswUZoYzGuaGcNxdDhQBuAi
wSzzSvtNAaRQDUNKX0j8Rj0F4Y3/NZAWTfqqhZNHRkPi331D4xSaXcLAdbD5kO3Y
KdNsgFEN6tcyf8Qv2lW1ZXQdg/uR2XpLJxHSSxS41Ou538hP6ctnRbU4iRKAhSZU
neSUGMQWrpZFRaZw+MULj9mruKQDDOUfLwUBFmjtJEU9I97LmFkKXalExCrYxqXx
R9edvArpFRbqiE+Dimbwho3YO1MkK0EgZHspsY8ishsd5rIhBD0i09RoKGJuJIsm
4f6Vk7kvHS2ENLoX7ZC2rB5K/g9nRi5641BRRbjwsH4m6uNfafrH/bIs2MHAm1y7
YovbGJoFYeiMqaABZEHSYzkoNdjhxK+sxCqd4tRwrove+aRWx09Vmc7z86VCvn+Y
qOs6BraAQrgytuRu3lnLKPFj29LkLMqEPEW0cFYMFFQqI/Em3LPhXJOAmuRm9EQ0
tb6xUrvuTyIUfhDpvNa5to1QEZbf3Syoqs8Di/mfC880X/QVHqTMeevpiipduavN
mx2Nfq/sFa5LVsmaBiRLSJPcqB3Aueop8NSpLs+78TpjB6cosn6dMjp56x4QfTxp
mYgV/k2EZavrsblQpseiw422hNd6KLIN2fJ05Rsbu/s4JUwtwh3/yFdHfEU4rcNP
jW1ze7c4evoWaELHlGUk9p/W1FUOflLxYGrpuZRPDA3oRTcBRzMZy46XDp7YQGbR
ejI1ghQgLWofFu3PMaaVZKuuFLIuaA2ByS+z3AzHsOgGI1aIN8j/5exUcjRIdCeC
x9JYt48yxkJBDmTN+K4ZrqU2otdwc70jKFCot/Pw/Zk3V4r3pHfz9sRC18LRT+c4
IplOEJIuf0K05b026yBjHjXftclhAYf5xEEC55h3WGrsoERJjEqg5EI1PS86ubRW
QttaDZ+91Hk4hEYT/TupVa0aSrEe1Pl+9U9O/1dT5ugmZ15iIOQhV/MlpDDtbiJh
VS8ZvOWm4Pkyk2sUHoN0tf1Vx7a01CLewNHaHit3Qer0pZIfMSvPbG4JOTyd2Gmw
bkrHjEuMbyhyHvIT2X2UfKRm6eu/2jTpMxv+Q8J1SRzKiWhi0eWnHXkCNpfSfI5A
P3f22aQ3hZffZPLLDdVFDhtxnmP0jBuGwDr4EFJpwI6nYbbYFSPRKHNdOXXHL6fR
bccBYeVq5eoURL6+CqJdQLZmr/tc8E/AGRsppRQyYEaFNwgt0DW1kwTsQpdyZECV
JGIVEJ0LUC/2UaPUKsL92kIXiyVrDH8keRwLy4iMCMfOneD69F4lbizk41SXEzzU
P2vKVmxiHmI7wirXqLcyGmL7AIcmKqzQn3mRGYR+CsVKgRZuLbGmI2MF13l3IW3Q
1LippHJaRjijuXoXTz8T4c4JrVFbdOs1u5zWSR3ScTQADbgUgwx6pa1y2002X1B2
PAOFVvVGcbskn1KB9RW/UPqJpcOJ85OHD8ZrdFPz+6FWiDiUcmKKk30d5t7MEpzn
Hqt3n/l38+0soAGnpCBfA5qeFgHDfo3wsKFNLY5FYCYLY8Eu79iy2mXIid67XqkH
Rle1nkUzLjwsZ3ybQuMSeN6Wk2VxqzRcaXR7yVUrYg3HQKS7K/VTKFLSntvp7CUf
xfwZc6wJhP2Ud+fqtAa0PEP8Zl8UUXzfKxbKlwD6j3Z21fw/lD451R//rvyZnIBC
KNjW7bbo2fZ+tlOp6WpQgjBYw07FyrH7so8wiODCwGZvdxu0iKPXw/Rn4dHpWgk1
zAG51MrCL1DTRpbEOcnbLi0URWGtObFigQALChe0/AaCrqpMSQv0KQ79I/0fPDIW
js7QGk/r1dbrRGs+ZdsaoK6Np0FznM/G/CJtMyU0tMr+kx/qIOIXNZ0DiNSI2kHo
v/BiZwDpM0Mtgv7zv8yIE2K//bKz7Kdsgfdd5JpOqJGHmHzmr7WzHSz3/0PztrJP
Cua59zxiTvHHYAMChfuKOW0vzQObTGR9EMp5Xlx9+fePAsrEH+xb3eL9bTTKbNpi
ttm7bVH54csTFCF3JNEnbXh02A0FMNXhgyqEG6kQfps+Frcugib72WUBBUJkZGfg
Kgvg9NDR9CifHSiWDmGzwr+eZHauvLb4XvenDUBEEd+zMYTxe0wQh2iAj1Z4P2st
PmCMGkRCpfwsI5kHDc061lxebP8NW+AOxZRacVZBbhQt6ShYBrpJ0sT2KzT181wp
xgwZowzn1y/wM0QLf5GliXlaxHhngLSpPaG2PVuGgDMU3qr4JWDI1c/XIV0D430i
o9G+XnDF1aSpADUDZYlIb0VmS85ms13fJJzZ/xrapWh8STV4wHOjz5eGi9c8MXvl
MFnX5cfF3NUYSqOXxZv7VZ7s2xNtIpg4W20PrY85cUdqx8NwM4BDzGPHYY/LFxyO
nqjpZT5wc3kXtu0Vp/acWeEbKAnipfHf99QysQbpy2IgHxgXwx6tkj9EShYQhc2B
e9KE+7hwiPsBCHOSqYrK9zFzjswmYtgvdo3ESGKubsKIgRjJjLAnU071YlbNYa0C
4IJNoBAAPLFzbPNFychV1f1h3dif7fSj9CKWgi0zjai67oNjEYR+IkRGol39CYrU
Y+6aRC7YCDupV1w1BREaVS3krJz9HxukKD9hKZmDgP/d+DhLD7BVLNqAKolD3/zi
DvHzGiN32riRfSaLLSvYZJCge3EScewnIRbo7FhkhygimTvsPjLoY2HP2j7VUr4a
JQs6tZKiRYOJTDFW/nHTja3V8GUt0CxcY8BLlTKpbYKZCgnCUBti9vnX8uLRiQmv
W/vbshy2OJM5OB72kc6SN9ESa/mHUVro09jy0e8XMwpL+KUQQNUHB/LVOCEXI+el
+wDP8udQRKFtBX2susENDmrwlAsOuNDT/7d+mgBUWC0zRa/bGkx1FDD6aaAvKh0t
hHMbTDLf2Yg+iOfiVugk3ustxMYijvqr1gkTze1CfSeWeDtsmZ40qpC/DAEm3r4A
g8PEejtrfhi5qLZZgkR/C8nWCOHEo95do7QqT+avBDAErp0nMo59/wnvKSr7YUur
xjy28RUBFzPoim36iOA1QFkr5Pr51A5KP7cRtNidPASZYoMMzTLLN5VyjEgSQ4EO
yYTNlSuX/8JpU2nckRupyRKyyuuGOtZiQMhjVlTlb3I6FME2aXrxO529nz3MVxyS
4jQ8luM3Bi4LhpdJ9G9EKUiZk95RcKTzQHX9k539Eq8mDrOpnrJT1HECpZfngBMA
VO41G4pDFGal+D2uDKyd38k40JHvH7kjzMa50bzzeq/Dj1gqt/O9BvIvBA9x18PD
98VMT1LU4O7zzdz3CR5UcL+e7VMXNtjY0vYCiB7wZY2DKFue4wdBZL2/f+SkM8y9
/ApYKGjUnD2BKC/HO7oUAI5kaOO88qrAVSRWEFxU73EwiBbcrg2zx9UlKiZaFWLS
nTF+Y1iJ3JXgMY5QzLIW0gVS70yL2hGyPP6ZxFOMaHGtgEmcpdscSssj7ADpv737
BvdHh68fGQY5/ZGzVl1tcwt2tEYiaX+hXPJdiDnmwBEmLxXIeQupi9FXzrEXWxTr
HkLhc8Fo1dXkqbr+Ij6YtWA4xMdUpBxcg21V5WrqzunwH6Jy4xVXnwt7csanB36h
fDY1GKPZLtzgE7IoyI0PyjXVFw9xRgT2F7Rn8cZD92wZRoUEIGCJF2ABXyLrCS08
TpQNWLSMF8yIAKNukdL0Y/HYQQKZ+KMtAbF445sjrgWcO0WxIcYZYQpy/zACNAD+
mq6uh0czI/maFEsEgUREVbFMNDkwnA0cEPsh54wrl091qEFGyiBW5gacdsT2glTC
0FKNaUgys64iFEK0R/RBs1uwMuT853vmKEUA6hQ7bCiyfZCtNF0+25WX4jIlwqO7
G1vTrPKtxVXKdiwIcQIQQjPEcSnhdVaxAt5Bz+iMhEGnbVgK8ipucsDS5/Gf41SZ
L6/VquIZ+z8waqpdvclTo7KOTbdKuf6syzcuCRxg7/hh58nBjOtl4QZBeTLRY3Ox
Xv60j+cH26q6lairhIzN98woSJ7lRPa8ghfl60yYGVIhzXc86MpuBKyEp8HjnGG1
6JyQe8EcBFoqUBqLewtLsDoFxxR23EL6J/s/iTnEJvb8CfkLyHtfVi8wlOw4RZTV
sxmCfAOzlDySWr0hHMu3nGF8heeDZGkmNNfzYKrrTJlQjatzlyNFI8kXumLojgja
sPbupUnlZQAFT0J+yxX0R45+HX7RPKbUaXRqXDFrmpnXyKHnW15GJXNaaskJhH5h
vE+TJmEJi39nHF8Kq23Iqndvo6UZWOz54ZoDgFjzcoOLckdh0LPQ1RTKSRfNGK5D
34AxO70mBIeBm66c6idC2a8UmWKxOMDFgdFjnK3LVR/OU+tkRM6xSf66NqFnrF7f
Hr54WqyFx1UazmkVaUJ/whyPoZksi9KXA8vCCEMlJYsAhGJU8qj244FdvXzkHzjc
6IXK8wYeIVHGMlTw4cHSvdMGdPPlWEzkXLmrAOLNk04CtQdXsVYoCtgm4DYYwyRd
l8c24l60ITKW0SpKZOpvemqmpVU1bac93Y4C83flW5sUZPufKSa7iP4asNUy9Yew
itX5IGF7XU/f/q6Y9oErtf1DeWnAzjOght/wDqYo7RwBNeFbh7Ol+8/LB4uE38Gm
NM03Sot7/fDQOyyj/qGzbL/MNkO5aNpax58xgwmBJRsgLwO26rJyV/MYz0Ba9Pvm
ZUzprrcLMM5yNWN3iHlp7dsJpVYSclQqKmTvf6x2cpLG+qmQb5/ZuYwkvSKZoXQv
WEvSLJr3+1ZulGDCw1nMivTC9/IVMZxAwnpdbDU9iDfWv3CpPatbj4cwbwx0bz20
0KCGUxHjN9BO6wUHUPQcCuuU6320Vie7S/Ns7+BIwkt62P8fKX/GZuPqEvL/wCV8
yAUSIaoa0PTcZdgskaZCIe60bBvfk/+EJR5k/6DezWRAqkT62JJAQQUDht5tnLfz
Om9OpqFSHuBGQyDOdakq4k6fQDgLHz85KON7d/lw7YYUlQO23AvWgFjiePAUPth1
LEw3LL9kWePQxPksCaAxOGPLWPzf+kuCF2fXXy5CHN7euj5T2SBj+yA7DTiw6UhC
+NZ0dCv773j0F3nHXekiFcIl8RfpMcYZ7kxJ0WUbWCFRy7i52iJ2RBtFXK+6fZfU
Ohxv0cWEdz6mOViMD3NxdQCzgXRnufN1VIDajpvQ8ZJdSY/6vzVdNGmRvvCGdDd0
m16CGdvMMA11ZAbNVfoHcDLpCv52vemP9Ouecv0vxAalUvcOUU8RjtJ22+8cdIRR
w++EWyqdI9dcrOudSAfEWXQotRZIUZWkBOSy6x4x/8MnWQ7Nm7l6S1nqcCPOpwcO
8N1DWseWLew+ojnQzDIp9Pe2OmazIeW18hFeww2WCBDRxdsJ4DY3C2KdE+toKDVT
86GhhWfPc8kLnOOguXewcffCrtQBeFA1QEEKyMVJunyQuD/P2w3zx2zHKPFGKsWf
5499HBg0obm+SSasS5NlZOhPe+OETShh8M+evF/y/r05tRjsQjg5OSsZD3zrLAKK
jJG5+VQbTicUo3vlii0Iuy1F1/Uqxgw+fXBOrJF99s2raBc8ULAJSpSldh/ajWN5
1UAg04DbKCQJb8RVWLw/IHm33G8Sj4YuXsBfmM1e/dGr5bzRKW3Koy+lF6RW12Wn
PuoZNCZZKHRC6S4txCojv/LrsL4ASuD+xlKsmfdNoJ9x7Pnn/YkHs1lFMwDELOqA
WXgIhQdNNzvitfUpU+UPjKLJIcZQivLM5qP4hDebtrx/P2VfhwCZLhsYwTR3cf1z
2tlPR9sGd4oHC31KtJHlpqo+6eWI6k4Rl+jlmU6TRbC7NZ4QnZYNNUVvuw2hlWLN
Ulz5vnnHZLxmxPpyqdc278CBrDXl//tjASZHLIAwiN+ncfAyuI1BQVXA/bsNzrxQ
cjJn6UugGZo2Ek6fEQ6Z3LxIeqDLHKfZ7QZkXfDXAL+yVEb29CWXDjB8lItSGRDK
/rFcYDB692z9kj4AXhQWpc88xNDvnDM4M+/D8CTuYCg1bdbKORCdrVe8fXx32dwh
MQcGL8XFdub/qFpGStMs+Od3Z4WDm75MgnQ8xwhO9RZkcC39Y4wOTEU195dcd0gf
N534d5p24C7/bqhMw5bg3ULGlay27ev2//BhxYNU9cSpD37fKA/XocaG/GwyxE0s
6d3PLJhknd5bHyCHpCERVRXbrMEx4xe/Df76AluR4YGx4mT32XvyGDfaPKJ8a3Ut
rWXLL23bLx0jJ1c9wGzRXU1yxQuUjLZ5vh5hzPrKgrfO4CFNz0lFF4HVgtDE01zF
fnDPjCwGV1Y9+Bp3qeN5wt1kL2Xapk+RTxtRWbilhzv6frbsRFr+f9G5vo1myB07
Jd0GiALHsQvFpus8pkjT0JsNNAIsgbLM+7oKRuHqb+5TA17r0wcC2OmfB/WRpzi8
LvpG/PWyunUcUFfibV3EPZ1e9V6vpm8XqstHeIggZTslNq0We//86+0KIQN0CEWD
ixBHp+WfZ+IkxeRyJ97LoJwaHUy3QcpucZjA16D44zm+YB26yT1WUlCVs2BjBd27
9iatFboQ1X/pN+2XScFuexQ10yxl43APE1dLIN39lf3sKb8QHgDQAIgxyDkRNV29
RRXy+yT5xicgp92x2TAlXyZrSN4DnjQ3uo33TqajpAMiCtbewV2ak1s3V+u8utUA
l2YgZVvric87N00UzkMpUr1Ds1/f7y4Kze1L3fLqjzNUxKP2LVSfqDMSsuTXGIwb
D/QkQQAdxTfcqj8jB2mHeBKg4GJ545WDMkYlWb53XMT/ZdOKjASXLCj2N0iFbr9Z
rS5kkTQORqUpdDGEIwShdn6O1maMjBHQnJP3A+a7s41tHroqkywfIUWmPofQ70Yn
ooqg/gUp7sxrRL4gP8um/4kQv1TcRoAJAK52vJiiXudpGnfAX6jUcZu6JRDhYuVB
/1tJMvbvC9lDv4KS+dIAKyVWjL7iUolShi/funuNHbkfzHhYpx2xNAjz6fjcw3Zv
lcmbmlJYCjCOGdArL+xtSTYusltPmCM50Yu2p9m4DScah6DsJ+i4sY8tgLlaVdU/
mx7nVPjLTMEcKazyAgRNE6LqHiX2oDH2jZyY+9fCD5hWbaWWQaLSBIm4QPlnGOpc
w6Kk2UR0+iiKfv/HxJ9vVFxfhYDc4XjXTML+do3VU0Pd1UHcKou4ieeRBl546UwQ
cZ6oo9bJu92F6NmzHR50HUyRCORBxX81yMknSBigqBlLV8fhLil0DuWmOLuBYYu2
+o23sncLNWNynbJCoRPPsoSQAKMytKenPs2p45d0jDeApFCFVv0Q0rAffQdKSeFj
XlufiEcbVmBjbzZZ9/s31+mbVRuChBtCh/PrIqGZNYOA7qxLmCimj2G6oP7GHcjT
iosvMYFH5f4l6F+6baiudkuDAyIWSP9SGZth6s55IKE1ljubGleLkw2Wr57x1ZA8
epNxpkXaAx1ulWrtY0EeHQQWpsF1ppK5XvYbTOvt3FOQG9fI+q95xpNip2Jw4G3t
38eMH++K9rh+N9SjD1YKrL7OiyI7osdAsFu+jqFCduRxyrwiwydLLo3ZK6+hsMul
GhXiIIXdzXxgDoCIr2JSPKl810+b7+uYA6uW0VWmKJ0Wqo/ca2giRGDd9b/y/TOL
l5U4Q5EFjBbZAl3QzMuvXULawfrQKegeUlx3ttuHSc9C2gESXupMcIe4tt5EVV3c
rxI+XeNkZdJGPjNlJtjVmRvdFDU1JGX4cFDb6gCJcApY+4SopZln2CrpuK8q4m5N
9YJcd/5mTLtnu9RdytJoa3r9zcYSfiCXg0mQ3xDEMnTmiO0d3CNaXD37h23BPChw
kd+rHcaDFkB/BA42mKZnsuxy5Rx/mJGN3EsEIcjvuJNDgDDR14dSJubnsueuUAvk
cgV+zIw9NSAZsIP35zW8cYxh7SvyFTBBxHwTBcuVIL7prb+LE5SBLJ3uJbUOOO5S
TXOq13c+/AMTP0lK46kB9ba1Z3nCGRVu7+4UORJLBJFjRa1z0YHx3VwsG7EyGlnQ
uvew8cLGD6cDx/zEa+4LPZaFciyu36ZJH51+5qffy4y5JMq4P9dmWSXZFm0gZqTT
mIFhBIjYI6fj+H8t+q3VD25mMMD2bHIYghRf3ARFH6lKHGv2N5aKGqK3vYg6C1SI
EXhK3pOz8A+ETlZf4qbR08XAXzOxZVk+CiwVDR2wd0amdBeDy/XQCnxl6SuYtVuF
XGfxKMUWEdjbVWKY4efBSD8CCMHK9pJX32ApszeJ8fp2kVdTPHBWscSYD+ujiX+9
Eik8hrEF5OwfgJfiwIuzM+EPC5NPb/lqJzJ01YnfShIak/zjUeObWRN21j1Ohx8q
+QiDK2i5lXhIgiLQ9bqkWsBWKzbyGcgmv9Qepj7goj/TsidMLdoy1xBYncrLyaHH
bnJt9fksSKd+JFC7GfW33c7IF+YQG6i6PoBSlwOHzlD0w3IBGuyAc3mn4TKZxJpJ
sOq0k+juuuaLUEDYG6LGUK1WxPn3frcUZUzn+FMip86Ydy/ZdzVr78r9UCr+aq2E
KkoaiiFrcLoWk+fF3YtNLWFejV1AARcG2iwsFp4fyoF4DYHQzrWSA/kKwQIR5Kqt
9TNzi9+FgGFU2V3+iQkHUMcQOgjhDNEgRPR4ErWsJISRScRaiefqliBQlWn60p3y
ltZndLztKfNuSnkTqWHOe5HonGdBjn6gO3SP0W7DlUoGy2XHPM1MEuJq0IrpmXCm
dsv8mtn7cg34M6zku+PwAsiHr+TY2WIsLxsz/cMg0G+M0xUSkH9gHipnl7gyjHup
BP1WkeubyeZG3+TJpbGeE30FmkmgEySS+fWHmIKu0kAzASeDOJWndbBSUt5rpl+d
Q9CKjnYYgut7moeR4Kf9cgYPJyeXZSg5hZ2VrMRTgOfjPVd4gkzwMdn5axTfBMZX
flheoj5FhSJmG22MtOC5Ys0SnodgJqzsaTvFWVKN8GzeTLNIzQKrH9Rg4sAqss5a
B5RtLKzNTphX8Ip8vLZbbivIWFmeNqKvolhxnfjCf8/gN088Au1+5nZnOc3kR1Hq
AI8mNaDoanektgKvZVnwPFNu79e7mgqb+H//9A5IlxHQSyvDND+O8x4A07Izw4JV
ito3jgzYXYOjAGUVz201TrBmunhsIaz2+avXbH4XQkfSCXMDnzgWY0U4P1WXCxtk
6EflF+s3xfWE8EcilY4cDNPOoFDMJHkXhKQTVX3NKBJF7CPL5oXh0CrTcv6b6tAD
apFl7PhiEnfwebABoBY+ykZgrRtufkGijbAFkF7WtUX7sRHS0Mb+WFw08TAlEZFW
iqj6bDLcNsCJZ9lm/tGkAjj1eUvt3O6ft8b7WVWm5eL+atWg9vWRrIJFiwpPO0ul
waYFsEjwuwbQ82SBl528gGtbR5TBSpo2XL6XaZSvcBLBfGJbDnrKrMr9BT/73XRa
sQQgEHU23unwYNWzSMxDfu6ZV1zjQKouMQHSNC8pB6fhEh7LknhytCKcnzfBQVee
0t3A53qXfuzvLW3/R7L2pPz8wXTUTvuckPwMaB1VjEZ26miDnvVCV1RD/fCKHjgP
7wqpPx9ffRzWsmeLSgxeSCASBEcTmkVBR9VRsasYle7uY38yvmTfGIqJeBi5tiJA
KEXlQ8gNAwCqOx9yX7mI1cd3JTJf+MgdqSS+ZnM7CbS5TpLZXspQ2UlRhQ9EgXE7
z6xvtRDXW6+jQoLkQqQXSOgSS4euywRqjPnU6d2CMvfoX2GT30JqBTAPCloFROMm
GLBeIoygollQaP34L9LyDEm0+px81VjLf9jdqaEZGzXx/Q+ldrKpruNSMSI0TfOP
ff8et2tvbF45d6d9AAPJO9IRWuqehPHw8ODV9W1WldS7VJ/1BmzGDuz0CZePGqGQ
1CnR/9AjZcfteIFNcRiXs/mssJL+6Q5HVWgINAPg22w/SK14wLo6jCE+EOz/dbAd
L5S4239748f2xFIhgqqRmuFU1DcJr1n1WiODg1DK2Z+YA5JyUJhshekUEl4zHy22
BtXOsDCAV5B7oR40vkYIoVZUrNSsbC8yXnxiH2DFXH0fax1tA8L18EThGSHnQzdq
ra4O7RxeICWX2Obw72IaCEUs+m8mXtKTHiU/emoagA2eIxgCCDGNQxgSTUW+1rdE
g26chXbSq+lvzSjJyy2/B792T/GKoPF5OoBy+NvCRxUzOzmRf5eA/p8B8Jjn7Ure
CrifucABlExb5Wti8V0hhY1/5rMBVdvnZi0qfOkTTF+IZ49tFDILr7JxYHOXwEi/
+HFVX8fGgKcR7QtyyEz+6SP9rq/ip/bGbHTb6c6A5gG5JkXiHD9dbfGHEY7LgWXZ
chciySRZQEqTc4ynhesvMv+p4KWDPNlsp8A6jGzoPCZRKZ7ADS5Pcwuu8dHSM9td
g3Uz0faX+me6IJ6ViitwNjTWfwMQoVdwfytQvPEkA9iYTBJdE8W1zEmotpsTiEwC
CVlmhgDcl0ypcMNfBSjUej5FRp8/8r8wKlPxYE6oaJlhu452qdaRLF6c99mGqi65
9B4AES6NpzxPgf5hhZSsoxqWg37zAi0sVqEVBNXH1EVSCgDqncMskHz1D4oAgarm
8Rns1cZPaUzw1bMJvHoouGSgG9d+ZU0fr9xILKV7a2WZgNNI4zPa6qFP9A8GomrZ
NjDn+KxN8jzqBX0OUBqDAvY4odi8l/GCqmKi1rtEM/F/bQ6d9Rn0/nsTdEDi3hW6
SVeF+5TrUHYrqOvN56Qx4x3upc7Rn7hL8Oy9dl1KW9a+vwtvEhCY0M1QHz3zhdpl
fQN4YKSHHXY5mSqD9Eg2UcTTJXgwPmR0/dBKjtWKox4ud5Z4+AYvjRX1XEfMSNrl
4eMUR9HIVp7ECFWs3sV5RWaBH2LaUf2UtQcfmejHmo6dN4li2nbGbUD4Hg4ll7/r
Ba50NorpGcHyXdM7Krb794qOXJ1moc5M/gZoXmWvTdf95dKOZtrMejjD0YfSSaN8
+9VqgrkgXvpuxtu1DPx+eDUOTBfkF1Jrocc8PukP1+tHnipQETQJRfFRtT3kZmhg
bZNZJH2yw54z2K3GJn6RGUGaDc8Ucbvm3TKORFiYa6EBY/JIjKFtTPzx72nyTjbO
8fTT7WwHotTOqIsUZW7MqryMZ12zN5tF5p7/KrS+G2nWT0nHZ1aeq5ZFDJm3RGKV
h/+RYk+Zwhi5qNz4wMxJq9qUM+Fa8g0i48RIta0OM9v0xpURRAaA1n6/SbhOUNgO
qZZd9bxiYcXvLAlig7zBa5LeGmsv8gMgzHX63OfIB3t7iYVM+8q+N1zPoEDsICdY
qUWJJ9uDw4juAvC8uAg+w44VtM7+886K3raxOq1FLpKIw4i7t9QSA14fSI9ttsGm
AHCYvrNYS4+9TiuQ+ZtwbKtJ1tSuGbs9ElG7fBkJbEtxOjjYGHhEFundD+BeJAgr
6Q2/ZCDdzzUiTPz8NPOqwbWwNvHtPhZ4WdE3g2yXiT4ePSK0BzyHWca++7fJ95/S
SSYtM2aFuERjJ1lDTWq4gdzZk5DcfxevCLP2N/9gYNRWsXEdolZCLT+tTtDag6a1
WMoJ1nY/GY3MEXNQjaDk+CTkXAmSeYKWb5Qs2aZmKTUerqgtNCvtfxHa9EC8bFAJ
uuwvWGyJUK6pXeEnDh7zI6QMWNLX65ljFQPfTd7uNkuX8GFkDAZQZtZCTTRQdkNM
XKkE2JzPImIWQfUAi9nB+o8YWay3O4o3Rvg3yWrOxtw/iAWt/l7AywQ9cLl1/wY5
hBVMYOY9d6VftC6DvnfR0NDhYs6EoWC5b/iM1LmQ2r/X+PVRYsjJzLByBfdZkATv
Og+QAOFnFZrOwiISv6tmcTCKfV3hr1FbdWmWS7vpb/L8kB3vEQDYbCCKB7qaXz5E
E7o4ZcBr3NE+OT6gYvIf2QhW7HcgrU3dTpTXOaqGBAD6PaaObrc8aKKlnW7TUwcc
TKZ31EY65eHFHoa+vgWo8AOl0RwkRv9dgQ3osl+Z+v6UuBzoWoQXLtfeR52SWljt
lnHSnTyeC2ltdTrfcE1iZV0yRWt5HO68t2PAavQBWSOAtCHwiVH4yipahs3Cz7tU
JxBqjQuqco8NPSW32YpVI7L8UTnFLeiu1360LRNlMzkhVc4N7aYf5mMFN78wTNGH
wEOTeE6IsAn90GlgilUyENrDbBsPDcHiXRZMk3NpN+d9HnnwqAWczKZwNISVLfDZ
oN76FYl59CPtFu/4wzPH+RxBSf3zQTmf26QSQgSK+3SvxO9gXnnpik6rtodEBhNa
rknhpxvrtGXL/hf6L/PnQ48bg1DtFQxnX5sNBFfX44/xOphiJwqJUguOd98WtNzB
vX+1c+L7yswEr1jwEx1wAbtjw1TJ3LJ4Nv80oTGlJUvHzuXcw3YJjbVUlsET0kPT
lyIbRP8kVeqLtbW1Ldszm5G1j0IgxVAP3qdMJfGQ8Ho4GE7wzXjpg7vYZbBHALHm
jNnObMhnDtyxUEpJJE3iWJz1BR+QthGgs+0OR7UEZLhgUSGhqBkjXJHcqxK72NKx
VvtKUbi4+RMOM49apJWAPZaiHEyr2J4ah4kRXP5k8YHq3/W3dZXXOqjJCHJ5yDUC
aPTuVZtnehj7iXirBZC9c6wuypIF9wa8gxN+3eeqDKkn7/3JkKWkJGY7miVasLTu
SLEttkXfT/ur1mJe/SaBPswUFL0BEvIfQ4nUitSh2EXgZrbHNAcpw3LlFqQ4DeKA
a83D212GB5OQYBbE3pXRA7q22VuMtP8rYV5pogPNzwxnMGG2SzvjSgLYOqRlcLOE
IJZBagUSIcRr6PTcvSsTgHutFatPgn4FAI0aEkFLLVgA2nxsC7bVKJ0ho0fKeJcd
eMNyQadoma2vNAzKBOGRDZ+gILYl0nPbZhbEjxItdEU5UVDhV6oDM740yBsHUcSP
E7Qi5dGXRe9KgpzH0GAtERTgq2oUUwD9m6KSIC7RfSPzLO3x7jOU/gQWdowKT+y2
DHiijA2aJwJjWoMijNa/D5qt+CWyIzPZUInJcJ8tj+3uL6A9v90zKaZyR/b1Rnsb
XZ/8FeNkxYjNUBEfqM56LdoCoaTAw8jhnB4hV662ezsm7z2zeLmaCmXmoFwyVjuW
nbePacioMZ2tFyjPVMT6G3sOM+T6WVvzY+t8zYfjRNuZRQCjuVMfOn3UH8nU3u8T
nJWQ6gXYYrR6DAsZX3ytiSLALj7ssh7zW7MhJ8/yRnKR0pkF9VavL70x2pbb/Fp7
glpl2JDeyD+tlSP3l8gB1lDxE/WjbSFQRSaxPloJNDY8lmPnocjFT4ZZx5azFStG
2UCKbetrxa+6SNxsqWMPfPh7L2NrZuoIdHN+L4rZ3X7uDkFj9A2wvONQfl1/+yvo
LbqYnzKoNIKhQmEOnA9cV7Nxj+KYXlTTy4jxkkPoc64rejdcbbTl9lEnY09ZvJY0
n4W5++GsljyLRmU+I86W6dKFztGrAcfTNXIKpR9gLKfObLgTt3Y/E4SmXb5MEZOX
se+RAWfDvlp4gA5mn07M2QXa0B/N9GpgAW9Hngq31y9sb/PQ0OULB/Wd+dn7Vhjs
1GUQPMhQcU5Hqr0Otfnm9CU2/nE6wkJBq8QLYepNqkq5OwrPrqRP2Z1qEUMbZYWF
Z8lb+Cxp/5M+Fswb/l6ZrufGnZ18eIClkR+mWscDxU95yq+CkMpPpcEqzPF3qhvX
tkkqaa4Jm93tKXYkYsvWCm9K91EMwD0cNvZPOSPZe465fs+EJYLuERA3WJ/MMn4f
6Nl0ZGNXjl5VnhHOm3DgQqsg4ccolJTFEq4P+8DnFsegJQPMjhoN2igvSukjCmPJ
8D5Th0QUiqe0wVICGxdyTakyW5nOzSa+y741SVzKsGkgebHX3tkjDiAhNau0hh6H
2Bj+MPlz8gDPsyXwL1ihFyEOO/ujsSss0RyMGTEwOSpZnXHu9TXeYzG+mWDFdMHO
3thM4sRRddlZz28m4y4vwPQiQFbFly0WSUrntF75xQ+YcWYUi73GQsceU1Z9ngpE
sabfbNMGWSZi49lyUkxnpw/wEoADQofBNuJbgk0uJNexMXivNdhQftTk+bf/IP/J
dQbKK2beJ/RfRRr4OVIzoYV/Wa7ZbuXJyEyBugPgfNUkgZQkhILbnBOaB1SlBSGR
lilEf1JPISv01ddBhalIKzAPnBoxOH/uMV2VIPTMB5DneJy6/wtwQxI6uPJfzgEH
5AR04ghqeoAl0L3AYt75onDcs66k+HG7Bi/k6d6X9HHs0/LoIGyDQ/2wk8gyYC4e
roDjx6PdgTffnaa2XXjXtXEs7AOYPt8hALk4flMckBfDnJLDKbik+KlK3aXMm2BR
4GxgAw8rYS7Q5BFJMbDxXET+LrJkiPPgJ3BJn5FOUvtojXwur4g+zKwN1mlaNQc5
OL9V/YRJNTFu7xwBdwTX43f4a//eA0F151T7hEEZ24oNQ4f+27P3FRWKsAOMkkOx
Z5t3e5YiqFV+RZ6BTknPjdgwPDcAOb6OdCVD/PvIsiSLeYeFBIyIFUAty5gMQ2r4
Huqeu8zbh+Lh/nRSlyOOLeunNJRPGDX09f5apmUiPDXIBOTYa4AD4bSUOFhGyYT8
kD6DbisAFdVJ4AK2xSRo3yyaOEecUvW3XBG9WLmFzfDM3pdSYN5A8Wu3OlBpysHm
ZQt3et/FYCTqoqhGHPOKRg5CzXpZalkjiOK5Z1uN8yBpsxuFwqcVlojUL7kH9qXu
HmBG7YlICVKKDn33NBtBKOmTqrklHx+hmeJPbjCvxmbQQ+bPd/SynGQaqfhNxzer
LqjnKQQJd5qsjbH0acJEFQMIxVBI5MXfXzqeo10/qQ0Ge5r9shktO7mBQbDYeP+M
FSbXLalwtYmgKgGFwxu3heJ56Z9MfJMyY6kV+R4Df0haLCYgKGAlkqEtW+EfK+7w
k1VNGL4YDa5piXYyJEB64wDUDV9MSAFROzxy+bPQ7GmTFs67RhEz2qT5V9AXIOCB
zdbHpoejA11tnxUBVfuvQ8jnQCe+yvN+F/vj3v2rTqvB6+Of0sjbcJEq885B/nwK
nIiZETLQhQ4uti2q0/Uc+38n5UPTgpD5VTpH3vdh8OTOTQ40dtWWqHL0+e70gJ/+
Qt308vjUQyG68k3g4cXP3zopHa+/abtWCl5JYBeyFGeHnqBexqhM4L10Zw3V71Ps
94n+cfmm336WgfvFz/p1yk6vEi5HtxjCd+fuPIPu4stieNQpPXc1yLM3AXB8sdJ1
aW6ekLqkWVhrnOYfthIUBv+jLtLPVxis5fqjBvuuFSR3NMMvN9j7EG6ZIO2jVe7n
z/6HZZFcEu/E2edVYoz2Bn1dms/jxFazmDeUVZ348Cumji9nIPkQETpb0XsuZH4i
vUgK4G/h84u9dyz02dZu0+WMCaWCOOI9/9gzgGn3uiDARA1AlhOMRbv2WZzfjAf6
cUw1CNLtVMT995mumNNSQLa3gJnZnavrCG456EDGdQxRmx1lBdSaK2P4JMG0IBg5
RO2cuSqnv7ZQNgeb6cDCPUcl+Y1bBaH3iH87yl3UQ8m612i0/2BbvVCgIVu/GTGi
wm+K7NuC5ZnLf0MuscP9LbhSitE65FpDprtylUTJ1g5PCpsEA6vd0SXGurw5SXcJ
wNoOxCVM1lP8hgDERtKhKuN6ETw3O75T8QKJQDbsxjSuoBobH3lZjr+a8rI4h0bt
zAuf/CDO0k0cOVCZoCY9voxm0Vrml7Feztau7ey2bo0ORPng68iMF+auHyinrY5x
cTiMaDtEQ90kevUf5QlzRJHbN31zM3noEOvXBN4a5OPEC6n6kgveX9O9/W6tZxEk
T7Q47Fvx1UEBB2uh5mjdLjs4xE2IwqFdNhMeTes1/2nhRmJp5tH/8NdFBc9xdsYy
/8rsS+TVQIiaBVmlJ6WgpEKWnn7oC5mqjm1TZxBENPpv4POztRp41sFtYDcjgoIe
3TH5RSPWVmyh1a0PvaTrvEdgkESM1C8b1+sCGke6znTAsZQpV5CDU3zhdP2QAEyS
E0ODKQN6HLsmMqtqg1y9rRZF3l1z8xlgLyCFU5qau8TwWIlGAxjx6XchQWX4g5aR
4XW1D+7YvB8Fd9/xMirzEXjvIJjvR7/o8xJ/w913K7lTjawvDCkjSNo/eLqYgRGo
1yENbjUu5OrR1fHW25d/C3U/AX0h+xx2Op7Tq3DeEeLMaZkqHX35DhLquC7iVkJl
lty8HSJpdFLu8mk7d0oUh7g7glqCn9pDHxI+QKS2YlmMrYtXoAItyUI2PxgwHEP8
es5fI6fKZZLUosXo/rDED1HeO1RhVByXSinoNMcaskVR7XWlGiQ1IsrHlPvFwLbW
rVu5L8cDb/Sk8S4k/mVvS7qEgoiTWmOjTuimWQEmqnP3xgTxL0vmHHyXJtXERYRr
Sp8Q8IKSzrYebGEjQ//wtLAB/jyLcotCGlqeKpBXBDrgj5L9leuh+8c1VczLFkZL
YY1cBgUBC46GXG+ynaBbAlrUaE4wJe6GUJn91QheNG2ZCexCNO0PToa6oovmR/Rq
blDR5gFqtFt+HP3eUeDSX+NWNf9EWZZlfIMM3ImaJIbsBqTlwrAtIBLlnwewaHyq
oq0Rboj8Rks4d4ParL+Fk6rbeZvCR8pLCddb0ExkMWRcUQdeUSAApUZTFccISyDb
BlQ65i6ybiAyXqKY4fgKsBDTB4ayz5iJ1nWo1AAnKLFasNrhE6fsKEbHyz2lvRft
rdKHuv3RvTppvTh40SVmztIXiIwiJgJSv0CMVcXZ1IG8aSHTrNYa2ybTgX6Va0rW
PMZzmrVESO88vv2BX+Rf1/0nwld40BksYX8pRnHBv6fd5GtmCnzxnxyphZcwvrpp
kbxN1YgkNTzwoTGDYKNJwCLQOZIevpU/QfZbz180YnslHFPACA6Om3LEhPNfP8bE
RBDQL1skMv+WB+iYz4oGZb5sgPe7w/UfZx+80Y69rs0Zx72hBKJikM8SDBgE+Z7m
0edj7Ixh/M2DHd3NW3rXfysCTEKxx9/fi7uFsvLDzXaH5oe4Fh2SVJ0wKzB9F556
6bl8Sm8wfQ4++YJeg3+4o1miULHP2j3bSnyvXJDxhfzdDSeIudBqtL7bBzOfKY7g
UX6h/kNZlYXmnwVzs4f4tPXtvBM8eUfNuUpIg0OcBNwpEmKGqpx5m+phvf7xrsoL
8g/4qcotE7PMbYLN3OzZwTxHrccY5MS6EYQ7zllgY0h1BcwTIZ9FYStT78/2v3zC
IoFKgVbFQbBB7mxD0cotJmfG0vGEV0sAjZbQO7UkhCfSCPWfo1+Yh5uDfejKs/xt
FZWAwQMBoCyUddzGoMW77+pby93rJQ5jwO7iMgT4O5fufHY3eDjKYK4HX34VbNA6
A1IfpsDiq9N2C3iGLlA8gICv93t7j2AStTJeo7G5dJisUiaCb0YVpELpdfDpdBdO
h+ZcYSTEEl9noBhayarmujHKxggckEvgdYvxKLu/EtF8wwrp8BR9+asDQikQaFyZ
a2LVm32Ekc5mulgsmv0vNEZQ3ytWPZe1Hdm3TMM5mr19AicoWGWBG/f8AZdnJWkD
UnVDjRuquMnfdYvmmgW7QNnoW8cZT838DFCII72qNdCKwsaa4ScKrGwBGEF0IH6D
oBhIjBIOdf5ciX/wineW5lDjMQ2kvOSd0me7+ofYzZsmhUM3j+8tQWHvXXpFEbwK
a0AGP07BvL09stNrRYEIXD+VREs/tk4MUW7bNnNYD7b51LeZkU+TQ5/nowOJFUur
76biyg95l+GdIvP4NcR7CqjXrR/dZp50CijW1IU5Il0w0YlxO1wxInUtlrVd7itj
81jwj2CXWyEz/7sos5NeHmCTvOzxQfZmoGsK59Gwh2UCog7BsYPn1DqQ3SwPjFdB
qhFByeBXeH8jxoiYj0BXfRUebaC5ZAXEQvCcGZ9t5rrfFhVvx6SrWGTvt+fJ5v1z
7ogphESedmGEuyM1Y9/KNAauNkOX5TUDpMV5uGm05fsCnzFp459sx7Z5INngB55x
RtzkAvobBp+BCsFvMDt86dUHxgZJCqP9R2FH8y5ihY3D06dSKaI/GXqgJi6TFQjj
LuU1nJdj84/MwTZXVUAT6U/Z1+FOdz3/FHzZCI9MNK6Vs4lGyvSNGiiE27+Gcwf9
DVHnBiQAEqo8k+jhd0b6DUlETs4/abTaAFOAvxClHqKvsnscWa2cuZjAFl9b6eUp
NOKlg6FdtDzHBoxFvDWpTx6oTm0aeIjtxvDocvsWCdaYMoH6bQp4m0iXxaRY7Mbv
87jg3DZnYVM0EgHHTyx7sdHYwTMD10zaPV9LYgRdB5WcQyCcPOtKYlGKP04TpUKA
p93zXjtOFL+Dnwas+PIiAvBJrpu/tCDufIyQLI3xkTgSPhrLpWogA4fBRDBScGIZ
vFznPd4SoUEBmIqejnYnhMDu8tmh71kME4MDyU9o9VJOEqQRC0ldKdVQcWZGaMef
CPqHdUxDXRXV9t0nRHwPLRf+zb3cdR3a+z6ap4OXWginltj07FyWcQXmEm8Ol6LT
w39npCnAfGl3md+9hmYqzRSt7kNzhFlA1nN+Am0vYeXECS6AEHhigNLvdVwP0W1S
lfKb/SIDsZIq9fLMufdO+EUw0vAWeRRDi54UFIfjIwond1ds5ka2Gdbj5gy/Qaj6
PYPVvDFm5Wkbcfru4Y95+nou/2I70jj6A9rfFSOc4cpqieGUqpyEGqyf3O6CvMAI
85XssiEsaQmKgXcSVCD6kD6DNEwr91z2q9Z7tGXADUSg9HdGUkCe7/tG1w8egf9e
Iazqy4qQEKySXuU0xP2m33EJUT3M//iXRWJ0hT6xdVJv0Mzpwq/+44bX1j5+jkT/
Rh8uSX4km0v8Mf4BV1dqt0UAwEQ0crF4MILTWgfrvWpOHhX6B5wpnLd1mzyzgZXc
h+/B7eAt7160gdblv+AedU2LA0esh4xTU+JJMpEjWHgdaN6uX69/4MFX3k8KzPGZ
ndWgdSVgBHOnPYiqVJ9cAf1lcNoPPBEWORxIkkXRV1kDdC7WZwhctBPw1nCSRuvN
4Jjg6yB5gU0GNO46O8fZ5S0evCsG2voJhA516ONNMJFfi1YeV9y1uAYBvLXZvimD
VbgbsK7rICiVaFGrnT0macE5Wic6e5NsADEzm5t1RefpisXftI4kq03JJtQrA4Qa
vy1blFj+zle0Vd3c3KVOILQfA+zf78o6/T4NxEpQO6OqSYVJ+ce7VV2b6LXrmFvb
zqFSEXbH1kb4d/eiNzevsnCJd/CjawlfM9qiVXlBgWqTz951snAo0Y85WoYxWv+3
OUf0Hxt4ZGsm5vQzMVb6nJhXEb1mRyYZpYGi6qyg13Hvh0O8tYR/P1z3zSQU9jK8
vxV+L25b3ucFssc87beOYAdfte/Gvy4QTErCyX3g2/VStgujtp85lwR46LdaTNIS
DNyH2RSCLPcZ6fQvQzM7nWbgG5D6tk0uwws9xVuIbaVmxe3ObDiu4cMEZF6Ew65w
lDiKMbLeOy3ixcBo8k0OvAsiuGZsggysQrXRRxYJfqbMDGmvJ1nBldueXkUmyE8C
KaRjpk+zDWgIFBX84M+/IOl/mKBRlQhKg9BgpuKwaGz4zV0e8kTNtEiBxmK1zw/f
WtNK/GuTAZkJlxD/QKLK3vYQPje6TP/DhHyKt1jLuoZriQyEngsRhKBpVYpBemmQ
H94myPmxGAYSgpuY5UCELWleAK8C59elKtJpiGByQss0qsWeoEiN1fQSoBQt4QHw
HXrJw0LJiU9wX7qz8TIW4Ffe0bPfyjqkns9G7hoqOQSvb8gLu70lRNl7aRkFKkLD
Tx36UJi+d5AMnm6vVe4pwlF1g4GYT207kiHJvmynfeVAChZyN4uj8Z+1NjsPI0KM
8FWt3tPS2sIc5ZUAxKOVSp+E6liaP+mfwfbjmDQQpdHprYSl2q7slFpvzQpdyKqs
q2kIjUSzquqAmaoYw/3RAZOJpK7gXzkdlf8K6e5OIopBiQf3waXGj6nvWwT83nz1
SOGZo+uXfewjXAtfhSIJwKxJKKgTTPyWmpdGSjTKMvtrPdzs33b3HL4gDCSN4Hv9
Bs9ZTgXVmuBSI3BQ7WW2WCE25w1chm/ZZdSRCvNqLOoWnAx4fPbnQRwNQRgoOsNJ
kDeqZZTAno7QxjOZBECwaXf8GLDW7ci+Szm7MtIOZeHS/+OUzbpkjTqUaIFqgkUA
WztVooK1Yk04abRffVLV4624FsZeFHdbJFcU6MftKy+58rNhPX8eV841owGslJ+W
4tSVlqtD3lAQBYNZULlNT2dne+MWvINvCJuVJkg3eP2Fp90R4xUYitO7/m9WKkvf
jGW0N+o1gorYrjyEG2qBvhVbKPINnnIMzMoWu1+UQr79zviTHjWp497QAMctLYP9
ZA8EWVX778xNMOOmMr6t5V3TddHUxvXBA0Czr0FkIPH2liaC3DCPo/bFRaJYCHfx
0/TG633PUYN4Zoo2saJK5vn/+2/mfYe/S0PokCIVW/WB69a+oKiu4iIuOlF3LYD0
H4rQG2QkcEjq+wsw8+lAiDMl1rthMDxVuU1ztEYQvK2hIaq0Z3oMA/yvfpNScLbo
diCRZmjTMLER8WoO6yE/et0zfL8xm6Z8BIYnPUaDAEfZCqRItsRWD/BapsOHrWJX
+AYPQTncpD24LP0GyLrbPnMmIz3ei5ILOaV8BG+ukde1v14ICQP0zlMzpAbij3pz
CjIxNPDssJaOWL1fCkrC9Kn+ehPb/KjvxX+H7/oEmKUQ2Ns+zIo9GGcSwPdXUTO8
kxynBWAMwrOaS+MSO7ZcqlOV66d7fQD1iyKuUgsVFQ75419ZJlwl30RYT9a4Jwy+
n/0m2GreY2UU6ChRnJh/LP4hTDjKRshr5/9R/g47EQYuGtGiTXmLduSYM4aQLq3u
t9A4lyK0xhcd9Mz50A5v54IPRgUa1AhHBs17mrVa6xJC/x3E/qz4ViVNGhUwm1Ow
ROD30VP4kNtrNPdRELEedl/qYQ3fGgOedKZYHWv2bgylI8e14tCO6TU+NwlYaKT6
olwjXNAaFNmi/xvMPOiAbaBEtNzooVpRMBnMv3Wp6xjVqFNSkpbEFMsySxBy1wi4
PvDgSHyRJsPKSoxzImwHTGPEtscJeFUDYoV3g6JEEIExwFVBnFXREbykxGzNB5ZY
5AjU7QKBErFw64eK19RWmmgeByGveMzfPiMPaip1Pgnc84IVQ9YSaaNHyYL6viXk
e5K7rNmmGK6oxKcZ3KsoUL0X3xtVcEt9d42fzgO6MfbMzxfRM917zBlGJNtMNcBr
B1ZYj+efrY94fJvCi3HVotMolcwr1+MM4nnVrTviRr9kaI83aEPIDO2vGI2OLDV/
J4hcjwMk97KuzPpvYV39mfPnCPKPRjMkxVmwYKQcuPyRDFeONUiZ61MziRZMWzvf
qsdBB7JoR2zIdNUOd+EEpWnM9Wnnvx9UpLvblpnabi4VCRkhFbbbC1DCN9jWLr43
a23r+nMptwfDABULEUir2RPL2Qy5clH/Jjw2bP7zqsv4amZY+ZnaRMYnSJ8EGhq4
Bz3IXnazbbc17MjvjPszhmgROoG5xaxiHaLa4z8ABEXp3iXFRmnBkckjnbLFLrAH
NVQxtgE1S5XqpP0CcOKIzo2aE/srr4rmoTP+K9RZ1t7++xwnuDn+0yEjQPh58svM
irq6WntIP6y0fWL587lgd8yek6ynG8L/fSyXGr5HXlpZoT2Xfw4E2a3bTevdMTX5
GLqv3TUnlGvNglRZ5uqpdB4tGkIPtrs6KnZTm91GF9oa/8OQNopxORTHYNhaskOF
3g6dme/kP9ldZR2CWSjQFj6T7kVRS3vHRzYQsQZo3IdzHzZMGvoxMiYao3i6ySjF
GpyVsnV1JrItNjWkWRV+Y2FXO1Zcf0VGvsNHbJIAYLPqoUewdzyxyfVUiFJjaAIS
mFFWUFCb+UXkaqYWG2I4E6EQDBfOy0Z9K2iWh/Zo8e7UDzHBcEQ9bq2W2nzjQgb6
hUm4EZuqhxGh+W20idaRLG9vWRPE1op1LOE0/tsBmXJ28491fqSz7oAgJU0fszdZ
LdulaRqSpakq47/yKxxfechKoKgXS99gd4Vjj6zZruGQR22gVeMeEAarR3tkRcTO
KK0fnDju+IJ7Q8TmW22NMKcadLA45eNVDQGYyTjbtloY8OOe4cblqJBHszomoR24
DDiRe2J6q/EWQtBpW8ZXXJFRZP/LF0sYwZFEocFkL7FoAqd5xhUqq1nvN+tE0OdO
xFQTeN+51/SYC7MN8ihAbd159g4j2Yrrd0sVRLrFY/wZfurtnbWBI+1e8LmJfD+y
C9qWLSYwYsUAQXAuAbgWUdWRlTDRDyOClDstVs4IXHpASymSr8h2MehXaN75Rmy+
7nar8kaLb2XmJBRXNc7N24b+kYdZHn3iEUyDpAVRlCyQD0wywf/kVeP7CNeBBKb7
HMJHeo2/jTXZSzGWaCL8xkHTnNSsG79yCOn9HblmydBiM9M//NibkrfDY01evIhU
nO4u2mKldQ4wiMKFbtquOVR1JgEwJULox+VNFGkVl/wjQMXGpTM6IxRfIME6TqWu
BeX5M6W453LA5j0VsmkNELUVIN05ERTPFoICuq+sgUYQ/4zR8WHAXmiV+PIhqrxe
Cp8XbfAOwC9Xl6qqcBVWnBgWTJFz/atfRB4t3t9ftKVXEq/rVKen2hswjE1QSe+Y
yRFDb/wqYymjis1L6Q607vJEiJUPIa7BprbIrVm9O3zRAQ5osh134BSbBgajy7Qv
LTqKLSADLmpju/7aYq5vs9RNuPMcKDOWzYv4O8pUR6GWv57WXWZ0++CHAysXkCMa
jals42JRDNV4VdydQLv2EkKtanoBNkurLpBeDaQ3gv18zuGIMZgzCD6Nb9mi8fjH
8Mjh4BXYeGnWmxdvEJ++9lvGAHxyiYKH/wm6qduYGjG1pDa9C3i7vLojvMKcmtgC
aHKtq4xBrlmGcDftOL9ByvZY/79GgIbkg3+rGx/s+kEeyiaBjYy97Rdi7d349+VR
gBJ0PqGJhyenly51YwqF0Q+Cy7H0yWM6Ca/t7szXZoVGsGPaQrSRYfrOLrQyR8UL
D6msC42X98nHEZuftzSBvb/G0FS+/RT5D2d2fYS1D0/m1SLAmqk03YHOyYmzroeK
TzjzJF3id4kE4QLcLuWnmleNxgCFB84FkUoUYeLiSGrEbkLUGlNwCpk/z92cAIt9
7SnfwVmIFojZVohjIlzaEyoAqvVB7QtlbBy2DpGgd69bGnwtmXKZNw3baqYVYkDK
GVVQ4KuUOWU7zzbYEjnij2CR3g96mNHeVHoum4gnb2+0ZLVEvY8kHO9O6TkpOHOl
ajf5T4K5RodvClqx4E7dhXJTzlhC7xr7wk2ngpUF3/CFZUL3XzqsEHo//u/coGpQ
+vp1UCc84UWfX3/m/2DdI5XOYIF+pzja6s3jbann1jK7mHIxjY6D/H9NOdtAXhjX
Rm+nJBrFLicR4cx9RjESuj2FLDbEV/RcqGBFyWzOalCS6noUqiZg8hEfixT+ZJnt
HCD70Veecb7b9NK2FZ9yZeKRptKaqV8Iatqntd5zbUy3SJPUow/1upo/ETz7PEvD
dUYMNhbny8KiwBA/AotBboYVsNjxZ+5MX3bIDX3orZbNwSdwAhjJ/h3VzirvKfHP
JwDsFJcT1IK9PWEOpdeSXjpsC0AeFguIw/jpRS/NGm8G+KpF1+OJGtc+JvYIwENF
uppnJbBYjf3g33BPh9P5Msbf8sUOz6CC+M5m3qqwW+56WBlg+HsDSqHpwTXlOriC
8WGbL6/dAKNJZXifTLIJvmRAxo4BPWSnUQFcV+dZmtoGid6QuDYuKMlUMOOlghtM
XSahoHe6FewNI9zWiYaKYh9m4KAzOtFVc04Q0y8zeHhRcaL29sYS8ucNv1EFTJ/4
qrPqUITF7xAn+yDyNfESJJt7qK4TwZr+V629TK+bXv4lT4nnbcqMFoFvqPmkhlRh
tDyh9V4WBnFHb/azH7JIGaO9mPAQiR8QeWfsbkquenxkL1jyo3Exls/NlG5B1g+p
7IfCFiMcLV+mH+bYb3i6MBbV7AGvIHRaMAv4IiZI3hrOrUkJ/rmHb567S/KjDTJo
0nZR7uPKWLSA6e5M5FDfy7noUkpwiUt+lgzE01rhim2rb4Jgu3iKCq+5gBxvYBTu
utfuACUgLFhpIcUdqciq8fEsRAkt2TV4W3gTsvrTYePkT08wqIYbY11tR04KPANq
HcWpbWyC1gGilmnvfAzqlgvCdui9bWK4JuSGKairrHi3zL0C3PIhq2Wqmf75wD/7
MAf8ezKLBZUeU1lj3BzGMob7Znko3Z5SLGagNQqey7b+Kpba8Utxp8C6t014/2zq
gq15oHmM+Kzek+WH9dCfpcGoyLJYAAuTUTU8ESjpvYs/ggJlPm69GfaBkh2aFN8q
JIUbq5G8OpTFJRetYOTZ7Cmalm0r4flriAtxAgQenqUiUUCsnqIrtB7bSxXn1i7r
61EVZ1BpcCE9UFqwFtecGH6YRG8kZgZDEs+5Nq+EArX4nQxneds9eDzm1YuO1802
6u5HIeW/KvvnrOBFQHd5Fbzejmw6+8tizzNpczd6NOnr1z2t7NIjBLamwMfoCkP6
Sljvg4g9zUCvPMdf0nRt0/dJhDfVav4Q+dMjZbV//wnExxroR6oQNKiaEaLwOdz5
8+SqbETjIYHTxfTTrwiO/BOA+GVo/eHUny3jy9d2uTkspyvmwbAKWEAtaVDhOzLc
7hwAvgIuCiWTLD389By0GEsGNz+jBQkO5aMjKn6//+xMxbCzNYHFbSRVZid/DolS
QO37d99U0R30yAoBKO4UhJsgVPSCHdY9A5FotEAP7cQzUv3LbIdfiATlN51YNx3D
b9gAJqeatdlU1upptWiibOz10yBrstolaBbaWNvNLSuHZgHFAN0VjhBKY+o27vdL
1RfY/cC4tcgzTImkTYl19jolGaG8s9b4e7aeVn+5a54l+D7VaxPPJ82UU5HxjRNc
1HecOGH2fH5sO/tTZFt8ftW2UIuOEAQoDfFRx7zZW+3Y0YvYqiKS/2Up+6FQfB24
Qnz3MX6eka7vlMF+NGOUEUsP9iXnNhxjPukineYI6Ehsxsb9foTAeXrqfPFDCQ3Y
34tTt5GDp7tmp7WO9Qaafk7nrktAupx1CssoHP42yuHTPNbjjCMfHOCRg7ZCAJMi
jPO964zBQV2GPi2wBcEzBPJYjUghMKz5fUe7MuDtg7KCQSHcYWgg3Zohg8EIOxiS
m11PxqJIsI/h3YFxY6RikuGZOhrFpr28qd1S6uePeGAQoAjgJW9PGm6tI0KiwiC1
8uV1gqfAyWDotK1rY/bdoJhfwlwjvT7ipsZWyHTMhFxTFnj72GHKTfEf+mojJrUG
QEa2lreLF6Wo3Ni/WjEvGIfakxO9EikUoNygiy9vOeRZiyEQ8hnR7yO9FuHtQW7J
RpJLOFGBb+OOPM/aBNcLDfJAM9plARAsAyNCYzUowqPJtID60I79JlNE2rLAJpH3
KltCJZ2aL5ALqmwZaNwHeRat6TituGFTRryfPD9FjVY+ahUsbFys5IWaxbZanEzs
1uTCsYsybDgyC1LAW7cE4/HDY7/ZQ6wzrK6q2a/ZyW/cAeBTJjnqW9+5MkZFcroO
538rZZUKwR/HgPjyCVkB0NOfPcqELlnbUeFM0YxNhKCIyBCBm5+ri6+tIT6DYZXR
E7uYG/b9RUMB+m3QvM4OGi+FOrV3VYKhqf3XAL6lsCAHEbUv7cE3TtyNIRKAtrIf
meb7A6uAIz83X8DRCCbnCUqFfJCxGqNGp+ktve/J3Eowl7HFN/cDlxdVOxkS3dk1
TGsZJq0mGvksbNZhN8sQLfj3Fre4ls5hzCLfU3M7tO7bi9TCgOdUMhxDfHCC1uzv
W30+Z/bby6nvOM6kgPkFmgZpZhkfEltlsYf2BWHCkw0+8ZCyPyZUelPuQDg0QASF
Q6qE+Xl4nzMi5kdM/vLCTUhMnR7khb7xz44UKXPbsxs7ZbzQiP9LWdcNoF3itK31
KIh1u7yFUmCOcyCNiy6E9VBnv6Aoq+iJ/9CKbAJm7tz6d5EY5faXOFEVMPmtPcES
SRdrjOV+tUYUkcB5cMvEqeWFXGhGlrw5whj9H1p1bzavDHLjfSh0dLTZ5GZLm0lA
aaraxLksFmaykvwMDyGulFzIHuZ9ne/uRkr5qooc6nOk31s+lxH93Gv1mKYkVhTA
hVSYgApMgqNtdu5a1+k42qb40HA75rXxfBzDSisX8qphqWcsF8dCbCKsNvkbjNWW
ji+BJhzqFWvBurZ+ffNOJ/+7TI+4K01j9QybOtlKdSAf36GXiYteqPV526Ga5KHJ
d07YwX8iK5nGOS16iHugyw6cqDGf+/aR3QLk6YGqoioaDwuX04g4NczUnh9IfyTJ
goisT7H00ypVcwD5q1ENVKxeiiATFbbhZaNnZ8mWTnHONbKauJ78PH+MHC7bxoe2
i4POxVACYcMBGTrBskwNKHMvyV12La9rDbbaA63K6mPK1KMW+zs9B9ywUQqMHdcy
pkys/Iek6sF8Oar0pB/b1Pf0MNVjRXbgpGdbAKL/1BKFRWXqw9GCp3me+7Sn3P6o
bUmv3J6J7k3TftH8sidswEuYsbV3ElLnZLbYUeVWUcJ32OIUdGxYRr3YjPb+YZnS
hV6pFBWtu8oHDNMhRc1H8sPyK7SsjJxiAWOPCtD3EUnRTYM3qho2rDrj7bI0Evi7
ehhSpdloiONv77+geSK+QwCY129kjGHq4KGGYeHHqt2OXemJiqMNoa4wLZPGRPLP
sPRGkDJ6A1dO+xmSahERlq9eresZGtCi9Cd7ANCV4AnLKBqxK6APmSHQYKAXc5eO
+3MG9F/VBv+kFi3HhH31it++7SgIpoyYbu2xk+n/cm/Lys+Ax+DuFFI+zFf8x4l1
FH6JZPOfVqdhE5InV9yKuZQKXlxLfY6AGl5XPwfeONb1Ydcab6BcN3NdgVVvzbVA
H/76OaVmukA9+4ncZdFIp6uYFgKJcCrlTkp5J1SoY/rvlmquxJ22X9+Gij9H+jiQ
0rHHmcwWvlM+O+H56WawkOJzKbwluatztep3IruMdgVYZOc9GHKKAawsgcCtIXw+
MfRdmauD+vU+uRHox8TQNOThfcUJENszmQGNDUAwLpSvJNmeRuvSASaqJxm8/qN1
kV2UGKjdvZKcIFAIye4Yui4avhjeKOSp151IyQkgM+7h+yRrEzDjfNbdM3aEG213
zeHfZMVnH/6Rcut7aDncKU+72gWnHmQjoTmZgVfVQ89+xaqeu+GZjMjxYDFkA+mb
Sot236tzGuC3l9RCkmpYiE0FExG/ZniAxHoEcAgQ56P9THMpMtW4cavFUlOY+LQL
PfjLrhUqgVG3aKIM9PQXPQiO9FxCiyGQDQa7dGOmkCWOWD6ombEOE9cgZXQo0YWu
Ol8PtCngzyW2Pg+7VUQySgL76wq766Rqy65GwJ04mvAKW+1zzXXUeEY6PAmjl6cM
sz8DU4b9zUGzfbWdtxhJb9q3D7xORZ40s74p+CiBj8iqIEkB4aTkOztLamhYhHHk
dvsbWFdFQIb+/c1aWtIsRHs4fCl3Q87MHL9o5cQRV9wnNad/NVmwEFiUGsUCsLc5
KbyJTggCy3XxeXkpHBIpNuXyRDx0z/LlohZc12fP7GiRb+EmSLyWeAnVWI1tJVf7
jyyOLVFnuWUCd2Fm821H5kzvK26Sas+wNeSfiRHOWHV+WK59MAkp70L3xS3McsRF
hlBUo2spMnngxmSp1W4D0txa6sZj4jv7nYhOualYqtCfdVyK04WZZzlMXa2005Qs
X+2lQxSbMFzseRvA//qS4tqNqmeX+Bc9Tcbf2iJlLKNSY6ujBE0TRzQAdZcv3Mry
xDddxQD+8O/mJlV5s4ZD+iVDrJyOVY39Ppnbzov53U92mSH2Iup38X0FWljYDrHi
5xJwCcwCfoPq0aZZKnEd9kBPyS5u8AXH+XUu+kIZsNMMde124mlDkRBXoQtl4DJF
6pTTL+nVPFXU2GiZ/A2KV/afGtESg6xA5rGohQtKanl5PeQY21m+HvybHz6zLgYO
RF4oTQlPyfD02mHIvpu2VdDQzg7abhJed/+x0v45kd086MexYXkUMGegRqQOHvjF
kTKWleuzMcoHFEFIHUMwaaXY6HdYPihiadJGCKNCfROjpKPOA0G7MnXbRC3BPu90
EaoXaAGh9gqNjtieT+9mufeNdXGjh//2Tt7B/rgmkac3cgc/dpjTjutoi7cjVVxd
nF8Jkb4dmruB44z+o5kzkXzP+vGID8JT8mT9EHO2EHU80UlfUnn5JfHV4LscUzqk
J4Gm7DoaEsziqvOKjUG4LjEDlkWtlbur0fUbcq1MFpeD6uPKfRNvjKsDijmFI0sL
7rYrxI8UZG3ceHM+OBt9CV2KMe5ZiyJeMvXrd8GaDh6rVHDUTtltbCKyhgcABtPD
oth13+rHqNlpeiRWZwlrvdjt+OMUXZk+ZYqG4+vOfn/CBPnesEE1V470y6QUPc16
D10LNQGnBKB8LIvHfAzt28a7JMcWn9FzFtotZQOIQPiQcTplFCeXWU3Cmzzb+9Uk
1iZhpiFksuCqOoMAm0f4HRJ4zT9a7grED1M1Y3KmHV9BjMxVct0tN+pw1wtcsdIO
D3aG1i5unvg3bKwWhC+CqJc1IWCo98UukSIDeMzTuhDQapajSU6tZGlgRjJe4CQA
lXlr1KgWgJ46FCIg1W9ODid/ShgX7j/AvMJ0QMJvzScXW7Y5tO6+Y4yKr5TE+CmM
DbaEPSgdpFS8CA8A/3UqNrKObIuQvEYw6YO6dXDr/x3KHd5jXONfFUr5Q0InEhh7
QQRBFLn1MF8ybYxhHZi2M5Q4gpGRLRJ+uHlBx67rc6ztH4UPv60JOKmkclyM0vuP
Nj3KWf6taGsBzlPvqWRv2Eva3Xgat/HsZVkmTfx2Op6UJkqf2QWmFPnTFJkBCjk/
aNsQv85kdCtgMPVeEph9uzHD/XNW5YnNiWys3ckTN9i/jW0BsQi3PpmQcl7SBz4U
M3YZYKADxwi4Uf8h84J6TZTax/eNA1aw3buADlLnyM9e1whWzRerYsHnDqq0Ufuv
3rNT1W2Z1bpCm4fJcTgmXLWW4reOQ3WUrbmcynA9oD6X8hIEkLh5tQLuSBA/u8ZH
shE5jRTdl6mASVshpe+O6AXrkrHsEH7/0qpETDzs1HK95sUsKah567h33hlTnIU0
D2nqtUe4ZNrJj2ikm4npnfG0bEa6JCS8/zyb6e2qVq3jUSADUphm4GCaO/m4ReGg
zeEvI+1ZTS0TOtHyShiNUwGV9aa7JiQIRLpZLoqZCToGPR/RHwOXhfgbvfnDgDyC
QnPLrijCFRdN7xsfNVCFdguOsWFYaWElAB0bmIabg9NEOjjx8N1E8F0LCike0yZO
+dPwbX++dOzgQZ+XedkBg475LJbHjzXrMhe0caCHVeGRZie0TFOYW/6RZSRk95Ku
pQZy1FzOEhmEsTWFh034sYlIj5ORgJ6F5GaBcUIkpfLsQY41grr4LREOV8/5l3nJ
5iePFNNbuiLgmeEHS6Bh/CubxXU6SKYKs0bFum/kgdLdzC3MSCFfk0pjSknepI6q
YGG3JBycKGyZqkBp4ET7PWoxRGAOSlW3JH/9XBgN6NzfDmQ9H+FjXjZlNbqbSsiv
LDWxs9zqMaxtTgb6QMjcYNxmRzPDH5SZjAYED7R+u8MrAlurELT5zDxe0Q8KwFLO
Slf9Jo64TTHzEQ92fYFUM0UUnPFnn/SPdBc9tpz95bTKEb6K7LxkW84vmYieEVR3
0NTscgXkxIYmJERL1JudBuMjI7Xo85caKgDSXt/vSjbQQvOrJSFqYHLQQGMqBSRK
Q3Sorq0cQ1lkzKOGObvxJuC/z0PULmI/OKiRjFMQw4Feeeyv1e1waDBZx0ZPc0Ye
1rslsM+/ITycvXTluxqrad5b1E3hO6V+Vl2RI1ow2aU6udCcNlcPnoIcbfs1V2Of
oioPqAlK3e8bRLxN5LoQ5SvMyKeueGLWrRD/iCbd/4UWNethWkG675DpBy9FmN4J
SAMjuAg3rzuXdbxQQrLTgAW5diXzUxgZ7vvs7d+K03J2lzRcCs0GvqXi75gMsyGy
E7x3o1cD+7TFc3i0/yNRwmSSr3uJVnjMH2+W0AvsxTsmssmfDY1g2u0f6LS8QduX
2GLjn3ehTOlWT5ujP9TO1q9R5DgwAtxux8Cbh/A+hnx1dvZs3l/wxzrPjFCXw7lf
+DAkEA5tl9XRZQl/BqajhYGel0KlS/y1wI8tRlQvFJcK/kN1quwTtE8ImmKxxn8c
wlB7Xaa5VkM8O14J2/1HEBeqbNGRC2ToKU16zIwwT0m0NgHsm6nRqVRLEZD19G7D
dgfp5rvo2kSZhNqRWrxtdpypaSm3JTsz3/uAcuT4Rtb9rjbJgsW9X9V+3Cmwv/S1
PN9Gd6gcS6hRw5Oq4FrchoPOX97kKLFqQ8Wh+m31oXXQBsSkVDYkjFIz+MwegMYw
hb9bImhfBvVldU7P63PH/19llpAj7s1nF7Lqmu56wsGNb93EzixHi9mLst4wbWi6
xLT58adNqQCkovb87WnDNn22eghjA9Kpzm8iBam64YNQZHXxPOL2FaPRk0uloOA9
8NG1D76hmlVwxYCAe2cCWZk5Y63Rh7Mh7kHnm9aonULBDurboebjSSHesJwzFB+5
p+6dOwLbqta7TyL2S0qkZN9dGa308NlzukPdZHqYC5K9YohxUmTcSUAQLYxE1rqO
6j41fb3PssNLYibCXuzLkCpw3vffaqOwRsL0T02t33zFiVhjoGmI/30yqmYpRPMH
OdrNPnH93mXSHfoPt66b7O3TU84gdYJAUpPgsk30gMz9oAgJ3eROsZ5amc8ht8fw
LMi667cFEIwG7VLubBEb5PvfnuHXjCY8E0AcT9nxPOu/SmQZ6SgGoq/PoTwOdRm8
KmJa36l1XHwkPiBs3CUaim8x0ajB3kMZ+623sec2izCiSjA2Tg86L9yaS53/G+CO
y4BwCJGgfbCgF+se4tVkZsrhENrDNKjEz53upZjrkfGay+N+d7jPiUAmmvRAaiuf
CEq2y+akZFavFzZJz880u9BhWTqiBBHI8158sRzXxM10jqoBxDrwEJAdZU454VNr
F4YNFrXbVbWznFdtDpAdM0UJtYZiMvvgbcZe1yuBzpCbFsdWq/WOjGdyIerHoodR
evobkQ6XWqFEMgTt/T7a165+UE4g815jMOT7ZjFk38hXcGS2kD/Yw6bW/G7BlqhR
yfpzGYKphTF2zhElvWJZvg03hTxyRSQLOm7mcJN/psBs4HK9Oa5W6hO4EZ1z+5hh
xDYTEPd/e1v8b7zO/s0bVkq4UesaAIemb9t5qw/TILwQN5f0M2KiO4Q8XF0TYpIw
0KK+3xU8OrribAkZzTIWA9nj58i+dyu9csFv2qUr0phkdy/xVtqdKr3w/B6Qx6Xt
P/4HS49sxi83hGRLNX94L3vfkjxaD/UV5o5+IJqp6rWp+LbL0nbnvXivaSBHsLTo
QOk8ZIaRiExwgSoQuPphVLBSltjF5kkuVkDnylR2MK5bC/nC0s7FnBlqb+W0qArA
fttIjGS1zdjAK3g+pysH5EvNflyKgLi15dIX96s8TfoLIDFDA3DZJXGKYZE9ic6D
2q+NkvFF8L5fB8uRBkravtxs/MfFgtwMr5YPqYcBNmvh553Sf31qSBIS7022zT0P
vPvS+MSTNGXnVta8EcgoykT90Vs+E5xxXONU3QK1tj4zZP7MQmwTPCY6Dlyl8N61
LjYyJ6CoSud0rvRvULicjpLZiM9YuNaRQW+N8dtR5qwGpzyy5pGMQzVN32gMwa9A
0Vu1xol0ozaZBk837YuH9MLVnIiFue2xJ38LY4FC4YKbsjeGeNH0j1ESwCCurHAC
1JF9HPq/T4ZG451whvqKS9odw2K5FuB3JXudE6lej/62gUhZiJ+Pyu6o+IUX17S3
T+syhu+BZYV5r+coPRjqLo4VXcluIzpwDyV6FwBiyemT4yKIErDSNEzTQPAnMYJf
9mglC3Nc6Mu8lQjVM/wCDfl93BYhUAmHP9XYbAURM/xKviXjWl/oQI1ESc66oqgU
MMSseKYuj3lgck4QSQ+WPGQBde5czJqlD1W7lnPtDhvkoNcBWqp5jPZmngV4Ta11
QcxsiQvM4gHlYIMa42hC8JQE+vAcjtmwoLwcXbB9VQmCV52XtvbpOAfvtu8mZQEL
xL36O+DPNPwRrNxk3DLdJcF2sfIRodW5Lk9Lhh3Hzif4YciX2+ovpRXwuCrEye1t
ZEqXjlpU5WumOuk01tbzO+PqJNf71nmeTr2QBXEjm0KMCWwtgvbSUmz0O6ZUsAvs
1iMH04lrE1hgYQI3n2QIiiMmSut7pp8cyk+AHMBWcDZvdZbFH6zLG7iSX6Efxi55
ct2Cn7HFRQC6GikdIhNCdp1AzRvrczsTZKPFWUypOBS6mtKs3REdLq+n86R+o+l2
q3byqn0nWbc8ptLdNT/FrMipks6TseXJm7waIlY7G3+OX+V0gR2DDC/bi0eU8f6s
jnHj3DiwjhGxphqVxnYGxdWhYSURPDttkb+BiTIqxXOlqjcRs6R5N5F505zxspn0
YCIQdnyVIi+Cx70cE6ToYNlxTHHNoRIdzUVSeAlAgHiNXhpUyIK6mg4aMgf5qMqa
o4JL/Zkn/K76rAsNdJMOzvi5KycAgICV+EE8YwBaR6pYCsOPY9QqGGW5HF3Z84yB
u8U9k4EOqMAzAHxroUtno6HV2Y4Pj756dXExL5qdshHwvOHzvVEn4a70dS/9uMRL
mKUKSWM5FhTCRRFWnyB5idIqBl/q2DEADcRay3sbnY3c3UGcb8ZsnyZbesLYqLhW
qSlqRh+IdU0C+J8xajJ1dww3VV59MkZySQvGTUTdm5TMhbMigO9ACDjZFRMOSkcn
KDg4wHRRdXv9KItnrlqKW0thfc2wg9uVR5wW/+5QLRVL5qTqh1Fs7qkqgYlqvKA1
MK+t2M4ZNTqNg1yKoNEdr16cgbNMxPe2cqIwbMdU3oXSAmJ2Ol3FjOm/T+BLPsPK
35srPv6AvQKD0gYH1ITplqNawyliuJFiKb2EZzoWPvy2wo5LTCMvJdVfwRYn3+er
ELzNrUBh+7eQS4kr0zlvYjOrGjZ513l22UPFILCel42PubE12IstJS5GlZmaxgwr
4Gapa9X3lmzIrJJmpqfwggYdBQnS45wgKa99x5rS1xSs7q/BYAQ6h1YgA7TzxL8V
2nz0RGsIE5iTc/JA6jT23ILekVf5AGsIc0si1HCW4k3NWKZOSD+tNS4fw/RVLkmK
V7f/aAcctdv9ZSuz7w8oPvNGzgteY7lndUSIQFOpxuCt6Nqkt5p2Rmhwdf438k9Q
NQVEgCrayb0zGkbovNZnQ77vIDi4grGdzEN36yBd6zT5iQ8crHfrga1mskwDzCVy
MJbWRobyIeMpX/M+GgwuIOqlOh82lZXa2uyU7JsYQhns6bWjaTTRg7tq/qUp0fkG
jg3FQ41n/qxsjcuZ39IDiSTbAmsaH+l04bFZBHEyjnAHAUFQBlqyTgCsq28fZlSc
bo5UTKomczQnfCAdFoVH2JkzpPx9Pi9X1TrJqB9ZjEete1h6Fs0wPht9EEHTB/E2
0SXpn24fAurIJAB1PU+MWvUoPVsTEcCdiOI0EjR6RQb3P++jPDhamVG6hyk3Y2TW
glq8mdBAtJMB0My1yKcta9R6lC0XwUNv/v7qnAY6wBKmiB8kw3PvcsZiD6zdybAm
pj6cnUNmxH/obCXV2RzjU7nUdcwwe0Wp9cgxYLieK7ll9ga4p5OKh2lcQZYTbKUV
xNQoNnA0TYDtk42E5QGuukmgnxAC3YpgNUtm+hA5eO7olozkY+6+pVI8arCUFWVw
pBP8kabUjyxntUtp7O+YkCslyBWec+Z7ldr2Njb+8YTyShydlK2/J2XR+Acc/JK8
J+1kv4m3owhR0ATPlT9O9oCh3pH+iiICSuifTilqslzDkISQfJv3jsQ2M1fw0Sf8
gx9H/UP+iVd5vYYTC5DYlOTbsBZAxOj7AivTycCzOMloTMMK0yA+ruPYja9oDsmd
ysMsfcHmQUmURphAdowggyP6aHUU0o/8BHen9SrQIuIPr8GWg5n/B3Q9EV+arsJ0
wTsHRyWvoLD0IxmsRuDGJ8LxXdncaXRq1Ud/LBeac11eGjN+RKAxeHPsTjlo1nGy
1mlmz855RO1tvjn8blUdj0o/mFTwAq9OfcUyMrDwJZsZzoGqcH36bmILcxsvICVU
MqBf7pRGQFIQ4bSgpk/KP4n3Gg8W7UqwuwNmNy740Zm8LJR5yjVLXThcfYId4YkG
U653a3OzOvv9yYq1URlBRzsv20yWybeILfF7XWx9XSnX2p57FduNJUVNQLQvOpQQ
k/Wu4OesBp0UBMCa3dnIKtq36Xu1LcBPK1fZRmYs2i0JYXzDcTsx5SORCqo0ak/y
fzB4i5wUW2LfMB2n+IMWS4dQDPfBOvJXS6De35e6N2vCmTxvx+1XWP9T3PopYafE
F32AJ47WROOd1kibt0CNalQJeIA5Nb8whYJ/rKyF9DL7LMqNSliTpYUdgF0qyRln
hY0s6Av3YsbhUlMCJdTeOvEbNfMxScDCtQFgSMKeK/QK2GfvzAD98yslKHDClhYx
KwHMzNlgHUrLB+IzdOEOa1snxzy7GuPcm2HisGAPSYhsNxQyfrrTNVq8TszkyJFc
tbAt+eJ6xskxU2qTaYrrlQkoLp+jIBu0K6ESN8y5Ju6Ne7MyLg96xBunA10VPjZS
JNdo805kf1htnz1w5ZJ5deRM31cymIPUcWV7e0ZOStrVj0COhga+pk3w23J3wEMN
SkZl/Xj2pIuWSIiZdl/20OI6VVLy7D5LomOc3PuZ8O59vahVbDVxRli9ALz+5tlQ
1PpznaIwH9OigAAqTWsk5DvwxJVWQrOA/wUnsRrQ6/zEG0Uy3T4E2syv+hYwpiIK
eWXlNRFqn9kooLTmBO6ugzIovZQEgFmveHpbWU0+UkVMWujpZD/NY4eZyyXYE6Vi
244irKBJFUZILhTI3XxQ6bHruYQmfI9NLz87sLnEBv5WMPgmLnrfkz3Opc2NOZxc
g0UKWBh1g+GdLWxeRsoo7tAlgVPKbhEs274WsPlnHUlfijFM+pgrDbVjCXrXms/u
4cOvxr0h0O8lwIWAUws5R7Ed4Jk2+Iw82jwDT5Sezh1MKDL7Oy/LR3Re10IF+yUq
SFwThsMN+liC3UY1XO4jcXJuGkS355p163U26LJVEYnWFMbr8gPvwm3xuzPuxcGy
RLI6bctIA1paytFUJwE0GnYDJJQ3VvsLwDkaTDs9UaXccJ9VO4UgM3R69DotDs71
l8sZNT/8XvjQkWcCgWhfNMg7H5y+MN6VTcFVWpEFpm0ulbtdQSvBOqJeUeB0cjOn
VeRZDCXHC44WzyCaUOPTOpR30ZkuFF0pDbbCpXq3xSJoWWo8eov78OfuZMbVU9Sp
wNuwM2e0btNH7UrlSTJqahWlQsMgL3sn1gyFAVgK+8h9JLUDtlnyojJD02ssQd/e
7oIMZWsSFVr8zQ2ShD4Lr9KJ8zYF3I007AHV1QipzUMyYF1KOrMLkMQgx1mvherB
PXrrIX+c8LpTTUTsXSs1orgIKeve32eFuuXSLLg+4tFgu/JtF6jOWKCgD2C7dR71
Q6Cr69KBTReoSTSpF09Zg7H+cpvjgA820aoFXTWHzhx4Zb4nMTwDANomk0aTxwPP
NOMfh4VZ4RZn8mpc/7bWaQtNNb3JBRuvU26DqwSkjF/9GqWvax6JieVQAZsf2PQK
Nqug54M/RIX9a2QOPEf4nv478BPydTCSS98CV9JLjjFiHE4Z7gwgQtYw+dml/3CY
XpTtt9rnEungFpCqTx9azL5rM6Qet1S/oDFfpWDPvNGhu1mgrGvPDiy+FJGmd+j2
1CnxmB9EfZI+VFiyXMGVcSPDc67fObApL31agnr8KFSty62VFEcH0r+tuq8WdG5O
la2z35IIj2FMLEOOQV0jAQHhQzI/JNwnXFuoLl8qZ12cHCbBGARsOZrRkh385VT1
JvyDXye3wmOgh7XqzRabXyIx1v9lb9Q8p5hqlX3/eaZBg3Z/jSEDnw1S3I7O8BOM
gPPfxkoNmZL/AVmf3eDfeVj9r5T7LgLDidKbLvYpDUAoiED66YPdQJUpSAvVuaA2
7JMlF1hDbt45crbYaMTYSl4a4NNv7VHRbivsOE/y4TTy1qYaBRuPmrfJb1TRynpD
PJ0zjV44vqdoqiMxddgsIR22v6uX0yXjKzM2imWTrVBi+lc0UZuCUFqS4/PxDTep
2fp2HyrIOUNsJp3X8ISYrzV0kpybCzeNG0mwZFr7KdK38ERelq5JuaMECd8BO0eA
rcXDcNhs2NTiZWjC/87Qq+LisYtImp2m6yxnVO0ZaJwdB7pZExdVdGTpNapDFQ6/
mYY+4TJ0zGvPiQ8HCgoXqadGM4jaYbocTCRfm3af1Zsd41XmRykAnty5ZCAKrV41
cD6K31UZJ656HHcuMfwddoxllQbICbKAK3z26xcBHoWMRTyh4KwWYHIRAJGsYQJU
hSTy+MikJts4WUFsYIocle68Lu00fahHK74QAIrcOczofeQGxzA87rW6SZbrf7bA
N6TvDfCIy9SDbxNudxCM+6kgEP56lYOn6flQ3ZWec3rJAt0ST/V8BugqT2EEM5jT
a1PSHJf1a4dXNi4Tic/NF5Le+yj6CQTPftnhcR72u3vFCsCKMwFUP/PKvMxa/hzU
8L0boxZ2JE9sHmywTleO14rGqYUOeQYnbio1guHG1ZqvXhdlyC8KOTyGa0a/2lGR
kVwWx321PBhsqAxJ3C2ExPgZ7tsImsmM/ipbCHbMaAV48zUqIap24fwvRtrrHqD4
4dPhV4ka6xWoNZEW6n45fyr0wFh175KaCLM0iwqS5H1cnFRrWgW7XmbS3VgGMbxW
Rub43UHdvLMg9HfQXMBJAbLy3EOGvlb6eFVq150tlygnR3aE6fF9dht+4iGChuix
MH71mB2evhKtnRxQucBL1SXmWomMEJ2Ybjv0+gZNuehCMoIpkoQ/QexIgHZG18oN
VfSIRgI9jaNmw1vHkWI5vK+iDaYIli1M0f7a9VB1NubXxICkdbzgqLOuYYKfLYOg
udR0ir0ZPlzRtyBzg28RA2j4PIq9+c5tnBYIGvcI/bvjLVEqXG4vutUZfDPMHRG1
OKUMLL419EbsxrhhiKXXBfD95fJoGNdc2NrNjh3y5g+cI3V64c0tmSvFL1CrDj0a
K5cbgWr6iJcMQcJHc5hz5QTLaRDBIpGLGe/ZgyPZ4Qs2pyS/2HPVVr50WkBZmjiH
wL9GL/YplEvN+PUI9U8amrAdgMef8jn5qwCp+cCwFKMgE+KuGOuyzZBIMpI/aYUX
ErjtMOodWe6otHhXuOORZnNc3F0m0+EkREJDfSNCHyor2mRtwx1RipEXKIKSvNjx
MHoKNdCP4ifyjKtzJV2e0xrM7GngJSnDmoczoNQAWEjPlwbxzNHxFvMEehR7aofI
usujkjGUS3dblQBZs3DZh/K1nheVZ5DX8A/12GECfxNfXgUq+fpbfU7C3C7+7YvT
KVhE8WZmwWGXHPeW48NA1H+9L0fTk+ut0Fg/QzFdUltGtMfz2W+oehofhIWPNyUI
iD87KtvlUi4EkQF4q6aNJRltNo29Ii4sDiwIyrEXEcBYEg280E1vakoQ51O8+t3Y
H1/uB2//gOLCrOpBIzkqhrGSlwz1VLTMmFAfnhk8DlIJtQiOB1kC2O09Jz23qEup
P9rrLhSw0XMNKPeKrJbgOOQZIoGwza3Tn7mvGH7wcEivQuvX/Sh38Ta10c2sVci1
1O5T4Pt6a8Lmp1EIUGGUPv1VzfePiuW0B1VBYjRI1boAkAzcMZmWN4mmbnB0txE5
foplcrdUt+q7lTbODo7QCZD88utRM8+H3qND7pM5LIe5/tYN6RbYea9bdh3ZxycQ
LJiIvdQfvZw8jik1srQvxX8sCla7WC+nRH1MxYJkMift1Jsb3kYkx4k76oa1ESfp
FgUb2hDSmrnJQwFIwteRUkhnVCZ/YOo3+3+tp0XiGKhnbcK89J6uOTUnSSWTL6vs
KOspNReFpdgKPhcNkYvS4ZltAMfQ5qtExIlPNL/HpwHESTPJiAZg+h/rfRFABM+7
z+Uyqa93OY7V3bv3bFviK4ph3q2ChbhjOSSPDpTVYu4JQeguSZ9TyB1szM+8A4t8
oCckuDVK9t3TY9xZcAxdfrCjUR0UXboTonIRGEm0VZl2QApxm1S1iMH0wqz8MnB3
kYkhf2s0qtZ+JoibWvLZwE8zw6VHMzJsaLWjpHHA3i7uzjUwz5k2MUA8SVwdOhlk
ujRy2TVRl0oUf1zwIMArbFXhd/hhDmJw7N0XjJ/2UMt0D+Nal5UzHT4KsGp0wjnC
yawtkKvpkSP1j1RHiceE40eloqzw8YIPz3FdB1esRabefwUqFHnKTYrggTKhLRpy
i4AIeTx7gwN4jrBPdj2Xq+uXJxiMvepd/mYK85zo6CDtVJyAu1vJH1z7opM4YBNN
tgWYeHOhZaaIZzAkrW8LkKmsqltISel6eQ0mEXeV9f33JIfJHD4/SiI9zv0QIEpQ
PWMunrWEvKn6s4im2LeIdlMOwr1J9GSfiyTURHBpyy5mR0VBoYb1qvu2LoKM5N3R
PJ97p79cb7/S1zNz75nmyPMdT1E2Lg9LHQFWeHhHUOfV9MqNSqW39OJW7v0p7sLK
VcQ353l82DbHpppt6vsE57QYQuqWG1Nhb8/9RTUb5B+5b+tExxbbhugexydIkuFy
YR5elaPK04lKsjPuE30Kct0jGm+3kVDd2cIEQ5Z+cI7HNw+QJMV8ccq7tnhVpDAB
6V6Nnee4/7C7+7rBts9lZ7oLz94qsCHg5wIrJh5sB+C4PPtv9nrj4m6S0HvFNNXF
sKBBteiFSyv8cFvIDDk6aQHo4hC5GE80VHD07A6iP6LRtvHJ3ASu4vRbStZRccnU
p2WkT7x6N0FP3BVINeMklB11cU/Ob8GD7DJr6VV66d0oIyyz2twKmFaJIkNeMiZd
a0Q3GXZwsjSat3E6b3mSFYHgWAUWbzV0yIYCVnwys3trh/jvOrGNh1WZ7A093An1
l6jno3gUoA1IshxRf5V5dmw1V/MjMlEacfxNGZ7z7vNmfnGHkikQF0qEvT2z40sX
sPMG23YiQzk/w56De1wV7j+FVmTm2Z4O9jFFC9PvZl8MJoSvcGb9+8LHQVOilCbw
7ebuXoAswIgOqr5CuZcI1jd4aLgkpiVe9eS10TDNwSMdxGxaUGq+kA7VXHLgrnH8
cMqf/0rv+6jPCLnuK/rFXPrIqwXxLqGyAczfQXj3hvjfgFIRIUWdYI9ggiBHW222
BxO0hhSwqYXc5yOS8SQJrL5aerW8Gae738HeIQlekyQ11MquwKWkU6gbcK/c9cLp
TnnM3Jwpj6h4kjM6bZI607Gn98QZt+fZn3e8PfhWQqGkmTAoJxEqCmPF5gq+Zu49
Z6CEVet4kyB7gvl+sC+oYqBTMair5KTWHl1qugqW3A8M8LInKWBjDIxDXT1jlqqj
pY3ZubChhc8ajFhM/t6JkKBrAJ3HJuoz3eHT0586V2pNgtBhwHsX5XDyVbFdbB8u
GdPVBKlhtsWSepKij6dLBPiVnjcY7hnoVdxRLqWLc5ULErTuo4I+TGP8+EOyul9s
bYGhyLqMkHroVVf4WsOPT6bXL9EyWG9z8fed+7Q0USqTHWbx5A+TsD/Gfj1RNFKE
NvMpEvKO2U6pFEEWtQDWTh6xx0SN4Oebiza5TVj8rbOQgapu55/GPc/TKpE/Sk85
hLTCAv762rDv+ULf1/aIEqOyFFtirXJjZB93DafWVSIyEX/Z8QdSbBtiknhpfrPS
eFHy291lEZajCvwuHyf6WLZvkOWuwGNV9cJ+nBmbzBSOR/f1laMNG5P9NxsJwoDI
yw90oO4KkUC8DUBEz2qjMrMVnTE8f43mcjRsZfYGtbf7gjNOou9xiW6eFaVRLgrg
m93vqGCSY1WAdzj2H1R8Xfwz7RkoigAbftDeIufJuvFTk2SYhwkdQMRsK/PKSbxs
4DVgTOMtszupkWCUVC+ueVmNJ30GEPQo8vaFRej/4b62cmCDWfXDdgWotwZxYrSy
DFwkNmYImGCLrZQtYXWxjNFfIkKCf/HaCKkUMc4qRt5MRDOs3H7GuZ2RGHLb4HQK
RFqRUBulYNXsjORCLWf0jun3tYGX0tSt13As0SYZ4B+ZhaFfssVj7/DuirorqMe5
Zz9DTkd1X+5uMGNMqc5NKKoHOEIu9hHCmTWcUyrBtSjZzr/YcdrrBd/ur24Nemdi
87cdBydmXiP2Lf5fR0PJ/iNat/vUh8Z+4e+db/J8iP5bdy/3pxUmZNk/A5+d5rjB
X1KDNjxVgl4zoqpN8uC35DJcf4cnFToQVZ+FIlrF/N4RnJA9bKw0mKUNZs6SrU+u
lKX0W7pq3p/rtlb0eN69GBIzPzjNicbmXwMPIYePVtyc2o1x0lPNvOQpeeymUje3
ItAt4s4uq+r5K1uWftZnsLn8dohZUDx5tfv6Dw3Wnhf50Q0GJBwIpNWvxYpYQzxM
5ze29fsbF/Z16f4Z+n7X5FMvzHM9G6+IezjceyUkrL0PYrtWj6RpfhjkZMW1n4wy
wRyASNDMcVjPTmExoNGuIz6Dei517wjEpwOfTSAlyr5dydV4hLhviqaYRjqmUBlP
00EdfWQyyLqN9KnIW2ukIK3Fxw5EXrGqaVzGMSieQKQWrzUQb6fs4T8IO+mRCqhX
DtWByxGMdJuqwR8FVGSQzk3Smxuc+r/qsza/tivyyQ87DDY28RArUZWVTahOL1+0
S6rWVJpSJMqvj697whpSr24INJrUC83hpUHeCI8hmIK7NsWzIWZxa+HsJn+9f+oj
TB8RG2gg/ciDAlpdR5V1eksZbACGhAbqU/fQatHOrPdPMlMY5gFYtWCY5fOWVVcy
E3xzm+EYwil/kwNAK82V5xidgn8Z/y+rZAg7ZSEilQFJL7glIeWLfsZvGRbv2fAc
kfMTo7gDvJG/yzILjw2nWGAeJsKTE71nNwmbHeV0rUerGBYU88k0S174AMRaPwVQ
ZXDbJ8x6x/s54YHf4QZ4wR/Qm592RUg6437aBRc6TqEh85lDfJ8wm5P3bto81op+
qwF1HuZmoQ+ldhCam2uoGEPoVSx1R3tpF8DgVaKnoPuUUd94oMcGbisWZxc/S2sX
DUbNGG/memEEpmDrjZGzYwwvyCGRjjEHvGtbOpoyMraDO1Kzfep4s3eyNz0I2+k8
Gu31xCg3RlSZ2nVod6+eSxU/V5wN6VcciUB6GqhscNzwBbFYOgSbIY87m/RSVP9g
om+2SD7j1ns4zbYxe8oFJ2JFCXoGPUw3oQLB0PxJoxJbpUqG8HDreT7NQpprOl8s
iaZuj4fnhI+CbFVw2Aaunm+5DoOum7756xD78qCJ9yK9MQSKWb4dJn+pkG2/ektn
Be3mC1+Qvkk9l1cVSAaGxd8XsiS678V50CLpKVhN8Ud3siJn6qu8eIlt6oH9uzVg
QoZ2MI2pYEaC0IZs+D4gen9tBrI5Ox3hV0czKn97M+eCNyWYCsagWquQAQcHgwb7
M5dv9mg6uH3iu8Ax8tWHiJn3llykoH1pir9z99s+VoFWqz7TfdXv3PcS731LL9QB
8NyGIwhqDrnEgt5jwf/j4cjlFMGfDkPIkrf3MyXvjqeSsd4y0piCCTmHfBQpr/j2
DndJrZxQ+KxYa0gLzmGT9BkBEZ8aJwvJ0borf8YZBVqlsGcof7HXoZOQt+//YpJB
TTLb4e1gkytz+0vYmo1Y43yKMaBwfz2Q8Lnrteb3cvDyTPE7LneZ9CdE7Xeef5zd
/JQm9lrnqmUyCr3VssWanl2HhHJbf+t+PbFX25A8aC4zM7Osx2A+ao+IJkS8RBA+
aJIBG2quvTjEYov/i6JXp9NwuE5lLZmLJrMw6s2MbBjB/B2oYYL+soSCXLQiNRa4
UHYHhtRMIl0gkB1oUg5nlFLyVf20vwmFf9/K1nvNwn646taSz/YzC+TgALqbh3AO
Q9mmoItQPxFSH5s4AB00ToXrYARjcbnVqaoOf78jA4Ob13+/cbp1ofVa/1QsKO+D
bkEraINxJS7Ea5dwglLlT229+mcnqJK2FHtnr5j3TdT7XxlODXe2tP8QqN12K4+L
wJHMmfZ05Jh40HoiL3KGOUZ+88MJeKfHuP7iAxbgzbxJB74Kj8W+MTWR2CYWAuZt
nUlQ22/a3uKSwrdc8OgXypm+jJ5VZJGwzx2SX6cGAg0OWtVc65ifXnzkg6/5j0P0
KDK1j5kfa5AxTXm7j6FOdMSzgyn5v198w9jknHENxr1W6AH7X1PW0zOYKt+h/Dnv
2zByPF+Rf/gB/bL2rvUeOQIicWB2uNYk1BM15i2fQ6dOLGh9T2PgaWRuIxD0rSeU
Ji1XiluDyZp1Hw8/3vr5KJXFy/X3r9ZARaieGNpFbTf1FExy3WVNi8RbTheq44IM
R/19f9gATbhLO2yfEY/3xaF04W0DUncXGOODqs5o6PkfdqdPmPVJkTuzwpmCt4+N
142recrWyRom0k4udB2LwgNsR91LZyI+0w2P91ZHsPZQdeLOJSfhrWXNOMweU2ft
Oc3zYlQInu7w7uNNQ2z81rAB6VmbRwePuPOrX70ktGDBcCF//W1EVLkeg57GfSOm
TeviZ6iV+30baZChkgy2uBBUK1pI1+N6OXmN4lFtvES0L/wdyRKy3fvc/g7DHlr8
/GdKmVld+UTUhLwYEHgvO04xh+ptxctgQh96mAlSpwYGMKrORi9XGCW887p8fD7D
JSGGFs74Ce5w0QgEFuT490yQZaBmCOPdKBMqtr3MZvkUynfw+00BI7y9jBjdFE54
1kzwmu1dyICsh2TviSBLjvY2FmaZgZ1+w3XQ/9vIYcdA4ZJqslSIQeqjMhLIjAfw
d8aXfqROf9hFPmUVrLh3iNcBv+lO1jZEqD0r8AYaqfC3vU2LI66PcJSruibrukvw
bqVNfDDh9xhCibUeN+vHNook0g3IUVhDAjqs9GJhIwKWkKWpChtNRGAbkAd53CHB
o1XrC1Bnrqbyn6s18Z0/j3DNhdtPgivbRJK4TBunlQomw3CDsU2w7SbeZZPMWgtB
Kc7ERufw9EwKHjXbZzN2HRIofcI9LNkofyjxVAJO0p1qY8ro8EjNg7CQ+NNfVEJX
m/f8BFeeWl5Hc0/ymlPllDoiH7BfHXBdrJXx2qeE27+D7mDdwTNbLMz40g/+mpZY
EFvPyx4zhK6iJh15yn4wtqSACz7s9OvRafBAqyawSA+eoyZuxoK1aT5J4X8nE9bG
5/nQ6Z2gr5UzM/nhwkH97e+zMyzAmBljy+8Ud90l+62uHeXfaHLhwhs1gwHE0b72
EErCjpxx1BdFBXrzwnHHXJg3R52lbnYPBHh40g3dpPPxbQ7Non53ha8vt/M5A+hs
yaeidiO3FXjtylenhgcveGYcIlrwyZQhYYmtU3CgWzWRTn5pWxnVbrysQr5aLWTc
7Udpfg3bU9w2+Qv0uSKnk4umCY6Ocf1lv0ppdWpoDUxfLeFahEXmfv8xw0y9Kemq
Ady8KZZLTgyajij3cuy7mbtI7jThRuuT8evTYAYkVums2XrqYObhzwrjblBoNOyX
OmMYmkNXdQvyAYinv88yC0V03vKvGhGlma26mLzgovv6dU71UZAH/geFkmWeIpDN
1OF4mlpEu1Xz7TWBKZ8JR4IGty5waeszpXkJtKTZdUvNkAv3aPnH/u9hTLnZXciD
a5w0cRq4VZQL9TjDfZvQD76DLNpWJscC8OyrnSOzo+NdF/mz9V9bVf8WF3XUZ9/x
6KuJx8NohxSMn/daxZu/MlnLbRlylxD4u+VoJjST7GE+7qRPPe6pTSCG88PILE7F
EdcpL9jEHxmodTbf7Ex+tYzr1WhQGBptLII7M7uBrrCJc+vJMguU5l2wl2zqjdbh
hQbvivwyxmP7rZdaXdUDPv188qAXFXACGmseQlpWT94S26xBib8bOzcnBKkqtV2o
NvMAWNIRGrD8O6m0Isnyla0VwFF5F9QAz1Go/Qp0W4E51r8VtmCrKHX6k9asR+xr
DxaNGWCd2BJM97fh3S+pLzJSQb+LMJDX2u1jx9DdwQfrsnoOBaGkyRwcUAl2Q0zi
dGhT9Rq7lyGQyJLcQ9SkScF07y2xx9uPDqktTNPxmqBMEnItY/VQ56cxzJ+y9BMW
1pFL1tfWz9bgWgf+LZKTY1FWRmezA70j7Sc5pgWFYc9bHs85YOwKvWobqKGmEYfy
dfeoOi8ry6BGx/AA0g66ahUwk07eFFb+hjFVTgiK5K+90BQPnJQ9/Ne545Q7T7NX
EXvOV5rN+vftOE1fY6EHQzzPs+LNe/xciCf17nK8DhBhVLMTxj1ndURyT5mpOwcH
bUXSIfmYK6epH6DSYSoNZA5oFChNLMVRUPuPxgBvHxEhe0F/NUl3zfR13LfXJN6C
A6R8Rqi5x9ogR8iECmFfCPq1Y5rpg5A90yr8DO+3M2UXEpH58rC4f+a7NXU72AU0
u26Jl6DTq958XbaZjhcCbzpPmk/ilddlnYwt/fHtOSGsjdEL4f/CrrWuHqem+Yay
bHsfbhBLrz4ySkiti9VesrEvW4VHOlEvuw2zvbjV+OMSieSyX406ItIBtd6tLZG4
9N1LpvEaqLh/U2qLtCAOPinD/2dha8qQAZgiY+UB88oNN1KnALKyZMu+esnYFxlj
Ch/e3yv/AB8i8CUEbLU90p4Z7T5eIYwQ4DuG3g4QJOnNH7sqkR1837+LNWwFXnse
PoD9A0rEjqllU37/ZWZwLczhOO4KM3O7LIroeeESQYomhNV+U32rNBnrArFKH9En
LzQGBTYF0GSaq52YgVnPv+zNNj3TaKcP3TRve5Fkk8eylxAana5y/o9THP130EKo
0Ur2jmF0XB0BvOrEdc/37WuM04liH5IsUY5hF/LtzAjzy++6FbQ6AoC3xU2p1UbN
oD7DO0gbbZy2JTLOpT/B+CEoGq/U0CdYKwFbVf65b9Rq3mqufFZ2OfhDvS6ENX8E
dKVvv1TW3mTVAITqk0x0PtYb7g7k08bbSFVNUuR/qa7e0rWrYxuCNZY2AUEuQ/bt
wIgbH4l/ZaCXTdbxo/EEZ7qYl58M4vGQ8/jIrJNnpqltJlzSv4VgqzoaP7QV9Xnf
XDYx2in2Gj4qfjlq+3Ax5ejwuh0fpgxTd4sYrFGgR+UJ20fFB9/HlfPIehyX7r0Y
QiRbJyzm1mC0NE/OJmKB3SVX25LvHCSgieetv3elYQcvG5IHFNaxoNVGDyDypUTF
woMLYhAEnpfc1oGZvUrC8ztbSxiDuRGbGvPetelRnKvXlrz76gkOjq3oAu0JBFh6
wDmsQLSqC72f9Lp50JrwcpNpPAmGSP+FhVGYunU6ZWyHn60OOwJi6yLAoxI/2O1H
GuDHZ+CLyY51YMpnWWe6muFkaywHB5nj9lQ7Ss8qWXY/M5YJsJUGvRW/nPmgai/E
4f2Kefe+4F56MRxdCj1hdBSHFWzeQRyr2IET7JiY3yDOR74EwLpJFQxRdUukiFqb
vATmHDVMfm2nosADgP+xCi/eM8nTyWqxJgpPwn6F8gOHBAUs/qS6Sv1A148ch8pD
/IMsXwI7f5Nse1s4WzA5b92zlvJjIc/QrwMDM9z9L9QohCLFb3HbndFAmCz0CuBK
JRaIiYAk3m8bjX/f/rgyT9HfvLU6zmWRGFKEiUE47/5dT+SfqYCVB4hJ76Hvu9ol
1eQKcGNPElpODmpsc04KjRgitbKHYXujrm2hC1K5/NZCeYyZFs+SoTmUzhhZCKsf
qqzHAexADALUocXganOcs/HIvUG32JPqXoSjO3TYodmcVirCQL+tS4CNIW3p/v1v
h85txdBYqLvwDjKOU2yIqb3cops6FOK4VCJUAaX0QYzmRLXvK6ZRLoIPqiU8ixIA
zECWB/ef2E+/R8nMiABzjVq6U3ny119T/XKuGtzS3kuqhs7+pC7vwfURWlNmsRob
jKqHSLK7Oh26mIDDXzt+KzZ1k+kCzl4B8K9eYOpzlsBwXDP/IBwpfHrvF0/UHwJs
PPfanHmJ/UVin7UKCAui/FgbBWgU4GAeZ/tS+esGaxMN3ztrUb8jQHZMU2QhVUJD
IxLmQdokLAsK5q9K1abr601NWo1s5edmGmYcnMGVsB9xF/pjFZPyvqI1Q/N/9/4s
GSKvPQp5utW1Jr+SiHZVrOtqoLQ+cAfXDv4LrwK3KWnnN7/JB59jVminI3k4ivDi
B9vdEdVNj4mMyEiYKFzqaf/TkNSvFxGZYzCtWXhLu6hzC/XziU7sME2cqLGxp+vS
ncQGxUr9edTh1T7zCiYjbn3lT1vNPNZi8RqH+H5Q5d1Fxo6+wwsjsFBCsjCsgoLh
WE8D51u8KvxwoZYPcDkz5wfV84O/drFb82mTdEJjf07RtAsR+5Nhd4wEIZnVgJOR
6tACmr/EWZyAml3xwM3kXLYabDr997Lm6KH1rgiO3Mp6uAiFhDBusiMB8mP475TH
DG/LASJTYWDS5JQt7mFsMl08n1G1UplStICyISsl4qv3xY6pjHcvRzdIkvnwwow/
Nm+zC7BdX1h0LabgTtrXrLbDD0EKiEElf3mW6VM0kp3JXUG8ppqjkqdlGS6KnAYd
8CTzU0KWNvJFjKBg3kZoe8dYOxXRBWIXd5LvyFDK31wvLTZ2kshBprNt6EnBhZXK
6CN64mLIT+NrDsuNIxgpwxfvLwVI0imQJlTj0cnzIFbZqFXURySoeAfZ/7DVq/FI
YjfBdgsyPyJGoRo/9I7dDIKKY349vEBFOt609oYthyXFYbwqOdMadE3oaVnxyBGU
05Z+c/i5qk8EmIYYPuVY/XhDzm16YMuS+5olR8vpTNk/qhXrHXp74DZW/ryQ74GE
MCH6zkw1XUMy8hKGWt6/wdegNVFzA1efk89d+LR40F+Xc232mnDWGI6Mr2Gp4CnV
NCiO51GAXSIJ/kZtvueR3qWKVrGQDOcpQboSvpwvYVxwsfEJJndAGI+z6L5oGFPN
4ZC8758+GGqjEAllXjgJ7Kuyv/5Z6whHILkHAf7pxEFWDWVPl+n44fKfobgZRQXK
rkq6b1mdyAAuI4e3aMrAu03sDEEEPYMWcqEgUz/B1A8n9nsxPPib0p6GOHoFVy6j
iJsH8BKMYNsNXLeK/x9bNX2W4zp9xRzJ3TolfL5HuLR4+ugQY8zdoilDoSXlXAQE
bOGPcl+bYEHWZC05CqHKmLZeZdz0TlKjAKl8PsedE/yBF1ShC3Wkk5aCjXiP+EE4
VtyaiLifXS/fJj20YcKqt4VmIFTbrcpYqo1YkRHXQ4Y+PsIVflzz2xoswoG32seG
XKEpD6qI0c8oLYj1rdcCM1atIdjKpcmkim0edyTGhBgZw3B/Nlj4MO2P4QfERiNd
LjA4P6a9BNsargVzDnl3pmuc18V0B4PpjFuFwZ9Y61v2QRnSUcu6QdzP/kDPvIey
nOqKtmhdzhNXcc4zd8FbRRgia7RzlH0ItJBSPpzFJccijJFaZvvT3EBve7wZe4u9
Yn291B/6Jgmtg+ZqAM5E2l1M/BljrfUNWtGk/A/jhXNXWH9yVd/4sPqEDQD2HY5C
gNJFcs5gnqSIkUDchm7fV0bntTIV+btDzq/sRy/pH6b+fayjqk8/rxbAkrBNb76P
WaNEefrW3NQFLRYNPCJEmloj+ICnjBOfigruV6Clr3GbitmEiUzODJPJhlQI09pe
wgY49/qNc2VtFiqhwoP8z6FnzzNuiw0hlxLapOxQUbFmlv6QTFPUyJfuSxIyzWNR
vNDYM6cBWOLgQnlcPfl5/vWsPvadkivs6pLcDJEgLuiIT147oBgeQUv0O8n3yYRb
rBaxpy6HWtLPGtHzifQ35K/I+yHi23x0erPimDfNOR7bOB76sGA7L2M8PbsVsBgT
QIhIARkl9K124w1cK6G40s0n4BgGK2BeGzkKbE981dBuqLAMFaowyaUW9AT+kdEb
g1IggYdicBUJQ07T/ScOgjE69rr5cUAl9iD6FRAiUNYayxTd3q24vFY2K8y5av0i
tVtKeapHE7l3+CTjV8wJ3mxQ18UMUGsGWwESPMbDSq/O4rsShDODUAQDtu8dMCdq
jaI/3K1X08ZHY2LZgdoG80/QlbtwtadATh1s0jgtW3madcjFPXofgVSfR1Rl2P+h
sjEt5gVWSrMGgdwRg1LnYuOG4afeD9nqJZQ3jH3BHU9cWXtPd9eZtBnAuk1tYt9Z
wphuFyvKr81jcIBSrMnBG/iiNMZIjcJv8eec6J51ZBvfFp9cOK1eqN1Cd6Gw3aYU
RZDJUa49UBMPYftYrrrzeOLv++IB23LtjFz5ExOpzFHPNsV92LX7u6C/gUXX5HVL
COK4WurUDPns2Z169k4K3gsxH1xzIPSt2xGxMASewDDZdouUa9tSlaQshNN2Fu00
l+sx80eu/nyxVOajFfZXjkBTXn6Y4Y0beCcwHdBFX9kuEQPe9GM2ApbxFJcbYE6X
kMIQrDZZ4Q9Ft2W7Z+C8loToE1WyENDcTptrx92WRCKeJXq+Th0ZHA0wJSIuhIbv
SVPGvWtWqrqqneYc+0TG8r7u2V+s1XYMgaI75L1zf33A7vYr6MmIxvqo/AmgJRwr
Hcnw4s5NjT6X4PMH4Uq6QThfVOxsDrx/VVJjYDlfPble7VeC95nj6q78Cz6XroMi
VUN26UR8RMBAUEo0ClIzSRu35ijAkSdwMPLdCNUgDgDMU3FseZSe3Fcm4Zr5IIay
7M3hhIL/jHkt4QJ7Bl673CKXy/DR8sVYjk+DavndCc/F3RlSzl+zePassjULMnGJ
lH/3RhCGV3sZH0yTUMjpMWibuXfWQ83GQSsBIzPd5PGTHjmiK/STc1a4ZktZtLMn
n71oiutXGMzDXiKgrjvo3SXyHTzP/CtXSvLEhqZI+IGbqJ0NWQ7LNrsY0GTLPE2b
5+LufCEFA7xG7XvSExZwb8t1SlVuBHxA+vjAbyGrqcjvzqzBh6SlgeoR2gZ+0/lR
deGrfjYlFw3L9I5LyLJfgQFoP9kbmhPOuiAzpttHF1PRE+r6HQWsc2yW9LEtOsCz
ew5xnycvIm3k0ksVnm/gtMggwVv9dgRD/W4OzT+YPYaj1c0NGFlK1zM2Y79LrvOh
IrnfF3ITrgHutPoIuhvW6r6NLzKdNY15zMCp3cubOHpqgawNddv+vbgauz0g/xYd
omkypKjMa4dVPSzNbNcTT36Hw21TF8NzYrGs7djj2gB13FSLeuJadFDojWE5i6hi
51df2KULjfJow0yMGjHG5qEjDonqxAJ1XS6vbOmhdgEeGTXhhMo+fdAtfq08WBZ7
7g4LOAQkh/Eej3cVOFoEL5JWrfhIYyF+hV66+ofq3H/mHjdB7AlauCviD/KE4fvE
cA8ZoWi1tfhRqRdwKauIESOlTL0EcoWLuRuqZH3G86Vc3oxLAGPaHIFO9nfHPdBE
bfVCKt+nnqshGxigMAQImhoUP4IaSVvCLydHIHqJBqTHZ023pk8PXNGCEcQPsWDo
UhpJO07lfAFqJIivxPh2/x6PdQHzu6w3l7X/TakucAJLhu7/8LjVb6KEzox9FPhi
DfKxMU+fq5tW3EXtiG9B6o5zVBRMI46NwIVAr1w/Z1ix4+Xx2biRpcoag6mhVGZU
ZThWi1xxvSOKkYcLn0Z7IiZDKjKJf3n/hpcSl044GReCIeIGuqqip8ihVvHjp9dc
37gQuBTso14/ePGSdxLr5AztyoJ731+H4IutsuG9i0kZKiJpCYKmTptkevueEQoX
W4yOx4hURxZGbR54s28AieIuqfGcqYQQ5rUI58Gsl+y6n24RHeQR1aGIT0PwQk3g
7wCmMmUHhDGrvNVpWzMSzQoiun9hKhxmOOOXyWAmBiyX684pAjEoJa+JA2K4VeCw
dAanBnDfpfwcNNy2UytBKU+jRNasTuoe0enzhClGTGav5VZXPcEYJZCXm2BgLait
zBbPsxDP/9snHz3eOeE8p2AgJ7nesqktFgHVYa6mMCxHX7PtJ+lsAIWW5Zudz38I
noytJUP/KYuNAp2bVJqJKtXT2dqABkDfKkIXQ+gMCS9wEVMa8SQZGJ/+c4bZP08U
Ka5pUKqDlGrmAh46cl1HgoDkTopJCjoj9thXPDyk4WSE6Mg/1C4dlwCcQ1t6XDP5
bsUOoH/SblZmVgRsfmDpmy19xubmgURWPQJDK48LZpN9gG7aDWZiYNjIGuOaA9wd
p4JCPpsR/UNF3JHoEJWNgnsnm5QJdotMgsFyUkvT6ARJHZRbsvKfEGFeQR8q2gmy
eIYcIGyZ8Jw8CWkOfFN5xrhRp4rIXebJoHihZGhpDz4ch44f4w6jGM8pEfFdHXc1
6PkOwMWSsB4GxzYUlt9wDthNs0lc6fSVESpnxzatRCwZBDdKe/DChVe+v+6iVDmV
QYUN9gXfeItR7k4ldpICtgrCkh2jxqxS+Dd1Bt5aW62HVjAnJSA9ppTJ8pdGdz8x
hK13n7eLVfYDD0H1nNX0Jn9OL38tolEnBtYOtxr6KX596jdMLfmoDfLqMdU4kCAj
h171pkPCfZV/vJnnKgG5zzWu2Yg/wdSv9lrKmlJfK4HSn+gjXHUcehSUke1NRpgu
eqkaRJXCpE6ObIcWsHvz35PHLCtG+Aa9Hf+PQDIbm2cbaPE6ZWgJ7A9fsybmCiS6
yXjASPnzwQxRLARyFPF34siV69N6eWEsJiDnjwKB4DQwyxvMzb3t1jQveZP4pR96
lEgkz0KQPFrkDtLFOWOEsC3gFsKPaxPRRxQvuveHQ3g74M6mStPe6yPVmYcBzZOh
WsXmjUs02kT+FWVo1OclKXfUVyEvL3xeXt7YX7C9FxepQs9D8BWp/oKTJxR4Z5cp
VyTaV1jPj28h+CpB+Jhtm4HSWc8I2r0fZfbxUox/6CgvZd9ccQIZSjA7yMx1UPLz
s+gcCas4tQIvnzkZFcn9x1ZvrHCHDF1ozohWG0oOXiu+9/tSM3GmPudadXUtnWju
VrPJ/bbsS4MiRuH29aZ0gho6Kbwgc+P1aAwbal/0ge/Vfkyv/t3KkDRY/51ztRm2
LTJsHKKPu0tleuFNau9F78L3+JgstDUKtFY2nryTZCw+kaceXmkbWLfgtqL7IJzv
BvYLjAhdG1G7ITQqzVzQIX/2W44uB40aLjnyfDBPRcQZObg9zqR977R2AdGt/Lv1
4jT5FHZjEk1/BGcXluEVAvSCy7fNsy/WoKPsj+BD6R6vXQHtcv9O1oGBWpbMVeYj
1T8kMeRmc2pvhVsmPwndf14vpZzyNmvjORUeAGkEmTtiino8LMEdyPJ21UCVjPz3
WlPX3jAdf2J9oDFKIzXT1Dn1nnDXHb317Pz8JTqzX0eTPMeUYuAIp5MakZIt6IQO
Ow0XTns2LLS6kKaXlw4wpz+u3Uje/C66DwEHwcu2nktyRWSFjTP0w5N7LQlBYrWO
Zx/6rky6DxOCM9UAt1uLhxIqzOpbSJ4PcdJYbcqgHWzWF+7n+ilJadgmoPxVF8Vb
PjHnWBqToH38PN6t+R59o7oG7Wl5KRtkxcRFPqdOOEkxfy7Q9MtThOJBx5BunXaq
zu3U4uHtm5d8lcRvHkR1WpAbwtqQLl2+d+obJgvDc0sZhEVTWJZ6YGgS80mVTuCo
BR/5L4Cp/XLXPGsYK8eEMCiTdPsMvogoJ2+GMpcXEfj2+BQqkDK3at0XKwTeS3kw
C/kmbr2E2R05UVgfAEYz1bcc9FD+W0XpUEG3tajuC5cbHIeQDc62LILPKsOIWU3H
tgiuIlOdDK3F5pPLtWMobNH/k39IhuSa/YEpKwGSelxOLhNpvsoFg4fJfmhhdYGa
KcyniV7qE9/0EMpWIBYYVzdhYzXrHX0h0GV7C3EbXoTFLQJWcbB7FO3mrYLSshp/
huR+z207qzdR1gfJ7xPt2M0qkIj/tx4sS1FS3q+PJPZEPkiuytfv40I1fh70jby3
yo3n+cc8Y82N1W93oqHGA6pKPMJB1kFHeVY7rNjH5gboAxzOFoC+8K9hxHUEg+6q
FlTru0gZPTU/dx5exPo28NytyNJj6j8K3ir/VGgI9kBCb1jQdKy1c6uRNSiY3Au0
4VbtttcvpCXyBlOpou9Nni9n//A3mFS1lXkhWtJUGIjvxN8XSuHQRDaozgKAxEG2
iwYHORrkvSmu2CoL4U8XsaMBCtHshEmm/X2dIVUTGAsC4Ze+iHZe9tAFjwJVrlKW
AzqSe5OvePhSeXidBmX5utlOZbIRJf3pcNHDm61/dxrPCTFAi/DVP1gNRsYM4xjs
8npnPPqw2qpWDvz7CgQ0J9BkZpIRtK1sE4vYiFS7LJX2Zj5Fk+Z4GTpkG9Jd2oBw
Go31njyrFj5emzkX5HnAW0YHfU70QoFue3sa3DWtpiLEC6BnwHfzhUtgG5MUrJQW
MgpUkBjKjV+x9daWunhjW2VMvELxhI3PKr32HKHM9dfLgem5M4isKlqryJibwJ9f
OQQip1ELv5OepzyqzEgvO83RCDJnmoDqGVVNuIjzRDYDQMf4tN/lTL31VGOSZ0tD
L3HE8h4XSwC2MgMt7Yef7GwSUUL1G+2CZO0cw/KBLABLsez2ESZtyZL2SiGlq3c9
/L4ru4De6cou4wiZgOJYQ5GhSPlw7XkdLInQ0Wt7jIi7a8rLJiQrBaoePoKmgyhC
0AWPZme4M5tP3xc0fr1alcAfPYqT29ofd0JEraXPr4Sz04lVCrptQcHvfhVqPZ1F
lK1G3KFoSQ9ctvriWrLfp31lRKZzz0VN5eJSFmP8FiKscjIgqVo4uFFP7llNu+h1
Ew9j0Duyb94Qjy8F6tevuj7Y+PmEZxpmidKbNqxoOmKriQ+SXCQWYdQS1Q6c1RTX
RKBAaNnff7Gp2QUH6rKZKNjAdKYloykvPQn7YeVD8If/P9RohJkkgteb4y911Fxr
8aEkFQ7UwRQsgp0+fnVMkvuliJzNiOICPV96pFGFN6jpp8jZani1SphkdI1Fy88K
z6/0y3HLxuTcJIqXvoR3a4mCGQUZa84pKq12KFMSrfDhsHnUsGHJqFQnkuy1ymB9
J1QU7Xa5DKHnoNqy/VAFhEJiY2XllXwJRmGzk1kwNDWUFuTouv70BpO06zwzVqyM
ctKfhrRpcTGK6LGRA6Wi3MIQ0JaOVYwKDCVtRYFBFkk8rG2kXWn4EAeoFCMkbWD+
8a/DtH0NZZFaj9m9VAyifga6xXsHL3bE9WOZm4zZaL83mCD8j0XTzWNP5FScYnmX
clDMT5OgHTfBxNYj/l6dg8VvLy0c4IqA1dUzWhuFCwf931/WlFlJiM9Yv7Dh+mDh
dwpv7IHEGEd8Bo5xwiAo5BDLpOyCWzoFu/GpJu/oWDva33cQ5k7KGagVmwMiM2yQ
DWxDC0YvbZDZkLUDmwwzXRAEcSumPQVRtvA/51M5bbeKmAWHwcojgq2KXDqJKx8C
LjDUHRbeZw2v07C7Cr8ii4CT0fu++tk84B/WmYqMrl2HZ4OKMsgu5W9OPEnaKMvv
Ps1xFDLbJuXhrrUden/JFAsv3tWkl3Df0ZnWdtAy32Ui7n1o4BAwXJ5mSiddNBly
RSdby4MOvCKlhnNAp+O6Of0etDLUcviqH5BDvLiGpGkZ1uo2VkjbgBWjl2Q5PJIn
s9dVe+Rf67uRpZXFkZY8QuT/ScHMRNqPIRbwCGw+zpmWmyY+T9Swy08mxEfWDda3
9DrTfZINWx8EkbujU2NNnXNuJzXLhrOFIUcChoqtoWN4EM+2LHt/3a6GZjU4DeBk
/5sFC4N1Wf3c56pPXctlBkvmq2CS+eVrCtquyj1sgfVxPNABKCCT487/Vs5tNf0K
0VpYlKgKbVkAU3/udDREjnNlcjwvRcTcZ6gdIM7Nd6yOnFw6lZbS68rtlgqUNqM0
xBajl5d3rgYSpUjynnqVCAmmJ2rXZu8+GtjrJ8N5D98+PFjwAic/nXf3QQ2LFYMM
y27igOzn+QqvxPe/FvPTN5jvlA/1KT12tIDoaVy5PPCbdMO3K2iyLxHB/LOaRQvj
lXsFhi4+wsrvDDXOXcU2MgfDikCRTr0JHa2pctF/6BQ688tnvu7CJApnc37wH+lX
Sc5MS1LSao3Yap107gtapATErCKTK8fp1NU1cIEOWL6IK96+DV77VFyOpMFOusRK
k1zSzo9fb8xBBW1h3MvhhaDB0riG2rE6U82GEGfx3u0Pv6yhbZpFfXhgW6di1L9N
8BpngLf+vxOg8jyqbgVb1YB2jeQt90IqeHHN3PKOby4dESr4pJgpfaX61vQEEqY9
1N9aZW+gfX3mV8utijkKGGOCRMZg2Yp+KxTkGJy+fkSPP7Y7l7iXVqPhB1S1sqhR
FTOk7hyAs165yuAsjfxd+2L7azQmVgmnqqUt4p4wIJhIh6CIWfHpH+1OSFY5jW8v
WVoQIIIJeipKxslUgK1UuQ6Fbfe2O4rQyBQl7m6pTcd6XdE4+shzS0OTWBkZgfsf
WAgx6pJT9Bw4tQ9C5e3GxJN/oSADlzKNstLcZBACnlxcNwhYpfxUGYxTmtTJkI51
V0WfUcj/exXOz7X0/OXdqNrCVHUy9IWjznC2hHhoaMHPez0DFMy3pep3FaBsZFwW
9cfT0mDWYEQz2Jn1kAWg/FhlLaFOEwpJ2b492749q/72rgb9kGKBiiIXDyV3MG8K
8Zs5eWbTRFlwaL7z2u5je/bYfQUGQvG7GQ/Mnbxu7vaCJJO0KNXSFVRX36jVRt63
iHtEyjsrJaJSCQQ9JSe0DSRpIILFXhN0aysedVs60e+KPyWV6VTCL4CDzszz3zcB
uflHz8N+SPWT4Ydqe7pH6QFUL2BIwM/fTF1zdJnkoLhkETUOuQlGRSCyG+0biZ0I
rLcyeClPBrXmZDpXSQ3A0hpkzYyZMB8mkGLigczOh/Rfh3SpxoTHg6Q6pu1EXjKQ
EhvDNMap7YkPJxA8Y/mHLEF/a5QcJHdQ3SL7ANvpexq7ApAK0jPdnGBfrh1VA5rt
VPdbnMTRMQl9aReMgkQHkSwCYwXibR3VLvRZNuq91h2ujZYABJeQp+7xDCsapWIh
+/6vWVxSwcAaZsmUznO+RrxZwXg5NYuQ9CQjf3mzSNwsoZbFJXpI6bfjpDOLtrx1
9q/vEaYqJa5tUs7O374ixxZsmoh3yNW+ZcABdhGjDBuDlbo79bWIoT/z43fVn/nS
4LJrcCkYffs8DmOUXII7qyewj+Ow9FlAfrgTwSXWePHg3st0/f+d7HFCDBBXfuBv
PKwu7Q6BOB+mA/Nr5yKYJJoZcoe+mivSXxQJh43bcDYlp2FOxM6s4PQP0kRXRdYe
HMcje0PAZyR5SHHraaObLqkb4uYX8quQZk7fcOL2Xsc+ub6tgYjE/kceu7mtBB39
LeQbn4TRnsHR7rP8mJZ1igf0cexEZkKeeaAceMtnEAxB/maPk+03XCQ+umAOkuG5
jIhv8IPHXYpFdPxTNRJqivXPSHCJOqRLKWh1aloU15unKSTDF2x4aRKs7DoqpSCJ
SLEzBXpWIxICN6lPqUzShQ4pOrP2xVGJuwdWj0nLG5D66OmzoseVHzMnX4PHvUpp
RdNvhw35iM8xpH+rk7CWvMcdUKajr+EZvaFVJJxdnTeBhNiJGOnyLTQrBj/wNza+
GP3e2Gw/8hcfbzQHzBifNsT7wLYhPP1piYihmR69CuWBSZvK94T4ocUnu6z1YhVr
F70QIn3lUzJQ7itCAXd5C90bbPJWxjyT9QIBHuTsmvTxvNQdgbkxFkFnZa/7lRRL
CruVfpV3jny5Crn3trajPL+i6MFuUaUgOY3iIcLbTVkQ0vhs0IMyQGV6TdKcVeWB
y7qvxDrngR/tEVFwRAE1omAEwrs4Xj7VKEC7Rzn7ChmhJ0On+XNaQU0UWcl7PS41
swKB6fFEa33yNxdG0fbma/pAl04AVnfqdxMmrzn9kEPMaVAjiDfBn/e7SYrXrh9m
hXfPOL0gaBKGRR8v1M3Agi6YNyQa5VexRN2iPX8K4F+1wEaTMdHLop9GlE+T7cF3
fJBC/VZYew7FvqEZ+kPwEkyDZcxQuGWV0B1rJfCyHgd9yzbmCGMqYbjOIGGg6Ovy
SvZtEytizqASGcN2qnlwDGtAr5hqYX/j8osaggxJXr4v5kZ7uOmvRViraln++Wiw
+I1Xs7YZUfRiyc2vW6wvjB96drK7x7AGLm43aMCdWaLyUgXn01k+YHyvB2lLkkE2
NtXL7H6O+tIIvUPTAj6/FOhT3jVVCKXku7WHaMETzucfqjF1n+EIOgQzBBwAf+Fi
/E+w7y66+TsrfzI+uq7KMJdNw2/bw9bCgpcR4JZ1oFWngsvoxT4lF68ieFD7uuX0
YtDJ71Z4c1VofhvKH2C3vU7B9/I34siIt1uyzTScjkA6ggXP3Mu/DnNO2sXIiE7U
vEG7g5aNaEuNxL/VSEwh4CcTRV0ak8qfi75lCmMkrwrf10TKnQNK5b8zblKVzUQ/
1gPFQ6cp48N7Y1Jd0LpcyFDVdq307Q3IZY4B1aPNc5leV6PeJ8IYcrgVhCkfxaKl
0SpgqbP6DdT9kF+G/WDBHzj2bK8QMA+qmoQoeAs0VCD4fIFcVbTOft2h7aXl0zPu
1bSb8hKe47gSvwnIwjQc3AdqMH7v2kU+bFceS34SLmoYsK0TVHkbS4E2hCRXcLYN
9YJ4dBJxY99flFQsXERWatX+juLzlCegxRyNnpYUbB8AdRjhdYnvIAdzu79ojsz+
hhazL5jrGiUsvv40+6XNk5kOTURpt+aiJObKf/7kyKgqOaa2TIikye7dLiIZRAGo
nOZfF3Vfn1cHmLghq90ocXzTpCI3ZMlnj5B0By41+oga8MT7XjlHVunrCwV13wVS
52L1EDkd+ddRH+yaYcqs8k/AnbCW6KJvKfkLywW1J46H+/D16Hw/G7/lLnfk8mKU
Rk0Csm8+88gFHPDVtPTXPsfd9HCX6lATq1qiM9+g1xv3LnRRuDlNxqT7VtK0DFuj
s1HZTjRCLqVrFxcL4M5MOMFTR6I4Z1nRVKEmLVWuxNeFhYpAgOlh97f8MbN4eil/
SJ9h1dy5HNRcOW9KeuB1xG0l4o4k+KabrzJgoEMRzhqOiY7fTBLD/PHddnR2t76U
/cEe6ZakQ1HbOBSCvTMUUlVDcrF/pj9mny1iQz8Qo8eWAJMNXEGwjkecQGnMrpJd
kFsxVyvjLJ5frHDQXD7tbwOB+GFHpCYTmNStJSzf09foCqbTLnSCIs01fqZT/oBD
lHZR8FPGZx4aIS/U49jUt7sb6H7rPdT/YAAEalC089mOHgg9J2YKmBpxiSeHIUQA
iKTNBI8giT60KPDFxblI+vca8N/5oPxpTNd2s8aT5fcKUyGXizDLuzgOE1jh/bLe
bqisAjWDkb0lwQFFIc9xQT7ErlbnYTuvQYxVXHvfGARlPJR+1jYpSTR9uNA7DHf7
8QWE4q1q6w2lXMF2UmjOEx0EN0ay7ab8FJmPwBQiMfk0Kweb+ktfuQb8bF9nfQEF
5NJETs+HVF8GArqqr52n/dIxJQxAIgzFR0+kisz0/FiKCHsnwLlbDiC5NfbnpNAH
ZN2y9Nea1ikuMlTWWKW0dx5un+gtz0U6npxAQdNWYUsJy1ZEZceJmJ4ZB9mTYcTS
99og+0tWtGdpnBObfP2CRboagOC7nDFiFeluieogqcTMKSEp8MifGIoXMJ1OkYcA
jP31WLg+rRXV0G4h80/SmIe+bZV4rpxCZR0ftVcBnxeNU4AzTZKuqWuRSZ0pr1+F
FE85UpVxqNcOJwmQEv25bA3xhPin1wODdiOGMppMHJcklneMSk0+F/UCXVVCMo1v
g4gzrlwVFzbbfLyR3iW+AUPsXv4xXzoS4CxRAJtgYkTWMAasNpSq3CzRpGLYfbY9
iqaKgT42u4xoaq8fzoVeACmh9Zqx1UPhNklGzY1zfGx4lLLFZlwSmFIxRtv5Uw4b
epf8jQ5s5rcpI3BLFwUn0QNPgHRuXT4VrO/g7+pIAv55B2aRIAS7vyELAfBkRv7F
xFIo43O22TFXwSyqM3pp10UXzsffInjCULRZ+QztHdfxWcAw4c3W2j693PG+kGsl
003ZAJRRWbNcE2iGEKaoyErQFIAAdQHH+mZgiv7ifHJJUrqXr1gneURySL/+UVz/
xrlc7YhPu6UdUJMYB3/Zm7Rr3PzDDoi+oIYzppyRXmXXw7jCFNT/dKvea9+DbvCX
RwDm1yN0pirw+tsj7OURdRuAMyZCBgFRbkzuR3U0FN4/wmCUmBv3cWHCJMBVDaHC
pEK0otQL47OVBJWoviBx95tJC30YUQjtG5sLi7C0vWPhlStOk8KOulOW6gkikylS
F6pUKdgmxKhb3ICP7rc/p0+/Zw3EQCEPc+lCRO1TibKXfl2vNO0RjAE2nuGHn2Om
4Agrs6mXH3YwZcFZzNhahtgYy4bmHK7PPKiy9i5678cL+5wm+gQGjAzP9k3obR1I
GqeUFjQHCGb94XcaEqeQiU+D7gpHGlaaVH0WmMq+9pK7cMYpTuJoXhlTooTKujCH
tRfLup417FSyoPw1kScDTmzeH0gqsv9Ts53jiXNOy9MbV6JmjlSu7zi2vGGM2h7g
/UjGH+iRyM3duhEnRnc2VSVVFjaYyrjhZbZxpE+q2URKBNN6f2DWcZR4AxANvMm+
31/7A/EVZLjQYv71HRPKU6WRdtg1gBTeQnby+iJaGJZJHh7iKaZyKbymTAVPCG7o
xMfZXpp6P3TgrKaTjK27/vyUBXOW2e8NiBKSDk+fn5X8v9pQ9+5YqKHmy//Rm/0f
uZvwgUHBiD6ysDpJLdfj9GXdFzmg8CHrj5Prw25/R0VESTIawjHlLqGF7YvANPXV
aVlcu800UsZtwdwX9t1m6wSMqhIku6lsdFVIjts9B4hIg/xMjhd6r8btYUsBTKRR
HGz3X4BBt4EciI/VI03csELADfVDqHevwgDSmyU8RW/fxiP8DtTRRl5Cyvo2mfpJ
QZWa6CdzuRtvPx31xCSQ2EOobzlIlrTiuSDh8pluhLVrT5vJaq9RxsTkX/Im9Lkp
ifZKBXaMlA+RijBClxcpuZExwrMcoX7+5oCCoHiVVBNkXiY6VcqDnfSlc3HEmwRj
nhoMqEKRLa0i7x2xrvEbcCDP6Qi0ihw6DU4ZACfzp39y31HQkGDDzGPqYRdHLMKN
fDCKXnR2NscVXRk3P5TA/c/yjM1j0DGeyr2AFIJcQ2WV2MBMGctr4IhqCrlLp0R8
IkPHk9pdNLx7ftHH7T/yByZTlmtcEYDMnEBS919eJ/Colc92xEHgGe12V4hy/VFO
AZ1UkFe1gkeGwB8d3AbKgORThWejwHW/29yHCgsbNJOB2C74Fes8F4fhMruqQ3j3
QZFNXh/xZiP5qcjk1PFU3SxHqvimkB9Jvwo057yjnDwLY4cJYaezZXjzB0ycpUv5
aJWfg4shDCWRI2Z33nDrnA+aJaVMx0tSVa8WJns4XVOohDQtAFIWZjoBb8Dufdev
TyIVUJOhCiWjmKBSCdhpWlubumQundEMbwFfb1lw+7GrDn/EBv07urZ0fZUZQrlC
Dnugu1LIkYQiDIs9RVnfwWxuAADDRcgHSgZNFhFHfnQayKmodf9siDBDRaelo0cI
sA5fmmAdep7JLC9/jIaIqiwt5Fqe66I2VvAVwyVZ68zXEUs767RU1JPzOjqBCS+w
ieXpPYsQf9qEHTZneRhzucCUTwqJ4jTj73est5lcw69+z2ygPeSKewNemHQBpTEZ
e9JxOs+xRzr9rHhe72LFfvBcqxoDLtzPWxpG5o0HEgJJnGRSL5JuSmLAAaGgWXIN
o7KoB4TFyg+2SbE2BbBjQQwbjnn4AUBKwo6w+wj0sCPLs2C3yFNEhiK9ep/mREHL
n/QnJxNaL8WmxVlZuA5QrBEIEu2CS4MHP6wYZknNvW2qR7AWT/HuCZ0sm2X0unQS
wmm+q9qnFculGei1lpbJQBSulUMl5pYrnMQxzc9gDmYfT0niUI+HidR0QR8UJ9XC
zNgH6hZonJ2ZuAwu4QQopYWAIskTHxM7dT6JM/k0yxIoG4ioQYL1WxDbIuSngUDD
Cqs3DjMq9Z80+7IjB1Qm6rWQdGwvTPi83CX5PmyhbMIWZEMF4mZo54twwoCf8bC/
X+qsLav9ZoRUseEbThSrhrrMm37V9+dYuKgkO1ExQlHBz4SEK9GIvxiVlkUp6DnP
wDE3h8NzIGtvv6Iy1tVEpYjzwXa249InerdjpeElU0Omf0zFqEpSUIudgxTRM1hb
YX2jiq5Cc3jjiuumYq9ixDZyzlal2UCZQLubLe7nGBIn8roSlnj9eTt1Wi6b/0op
HD2b9TQGEqiqEaOWrw1c/wGxd+0NgpgttrrXN/RY8CjAUZkKE++TSIaXpSgtNIn/
b9tmj8NbuIcWM0upnUvDmYcAJpMyzmQgDVQ3RX822nc2NU6zXuo0hdqvuAy0uZKj
r8s0DS5SgmNTrgLbcqxlUL1wbb8IWPeh8BlC/LuaZLlxr8/fQZvO7DLnI+Sn2CcZ
q6BUyRW2U2nRo+4FzgcV04mUunGDvwAleyaERsRnFoi73LGFGFruzok+Rq0cjWc/
Qr4tt0omzvGV80sAI419xWFTQqaQdYxCqAXEIZA8oJPd9/wNi520x5NoviwBV7TK
Sm893rosF8GsUwhmshFXHYfBE/RI2vqYlKl9RYWzQAOHUBWBJsb8eMK1KYL2cECU
FbeNtD7+3wwrgGiagTturFeX3mR70C5xgHok5tTTJlledHkI3sFJ3N/mkpnc3oHZ
91u8nbJAIkUoSEhRYWFexB96LO/MpEqjDKW/BKdI4RhsDe6leJ00XJth1KqxjbX2
bkGws5CRun7qWTzpRCGUz9UltvCaiWpp8hoyCMJH3n9JeQgKVspE/2rpj9kW9tgj
WdvVlk8IsPrp4Fskhrvq9YyXKVMQouvs7QLkxyCcuy8T7V4RD7CeSBtCFKO7z4zP
SUc1/yoPvr2SieiRXWvHJn2F4POjVz91mgdKjIHusjaZbQi39XfkQmSapxsoEoZv
x++WxdsQXpRG5DSr/L+k+dFepUMUknAk1KuCH7gw6bKPbz+Xq5znVF5fLw9gOcl2
GEeE25bUZa9OqRznF/6v3dILY5aBHFFXDiCxZuKmqiCN1Pd4Lz20jOZuy0SKgmLn
7NUwVrpQBt2P7vvBdG1SdcSzLUhrJ/PDXzVq6k4FPviSiVy/xgZSp/nujXKHO0kw
ZmIaADONsLORDASJCQ5KFEQOtu4Y2oxWsf3CyWAdIMlw2ZbqDtGTSCcfHCk0bW5h
9JVQei2z0UsOPC64kYLZgcasElVhAbp/E/seIKW+LNL6ozIFqepu5t+2voG6DYhR
21m3VwCT5o/9YqlsCiMBLij16Zcrv6M5iCgAeieks6TE2S/PbwNGq1hxULpD1lFO
XVYhYfEndVwaXe2bnmdd8r0hg9J/wxW7tycNvi+rSMnx8uyfxeVAfb3LkYYpBKKq
pOXjQF+A/aMNCknojceSNXDyygl+efb/JChRvsmA5AmhnkOjKysx/kLFC/ms9G+W
tV6TH4nBSMd6pynCDhUeQgo3DdWHGtvuGHxQNNbZ4NOHN5ar1M9xEWm6eDPRkNeM
HbvhY+jt49bhRVSZCqIORmpHuj0cx/oRjGNP7lF8mdIijehubTDDpT+Wk6Xv9r99
LFabie/6PdPf/sFM2VNBt3mAdKL3YUGW2GLQ+U1vr62wWG7FKsB7vK6OWYsIJe+6
OgkFaY6CMCrFYAlGauodSfUenCBKq08zYCiO8O4guwUELMIsnPkFFUJDSTA1pFy1
WcL4w1oT/UGK2uMBv6jUT2QPGtryrwI6klsuy3DGhfvUDEGN87M+2g988ahDefH+
23BkpOFgLkL4GMYjTJqU9awrTcNAvSgNhO61KkcebDe9bXDIbzWQa8d/faZG6LDf
G0Wwa1gvqE3GTifgeQ4vgZa5JtzKtfADlrYkPNO3P5un8zXvACcX6mFmfh0LmNzI
QXSssYMIBylsTJvntPqZ2JdNW9g60G4DmW9jhboNSyisLkVdsTP6fSAP05wnGEaU
WEUuMDa3x0sO7hNVasT1GChr4428kkiL7Iv/X5AD1ncNB0UPSZ4Z5JCWD1QceAY3
CFGta+6+MB2iyJHx2KqaXo/Cgjv6YLNLUACueaL/Fp761krBZwFUg5us0WlbQaOJ
NvA5AqZI3jUyfMM7821xhylbPhnCXEbKOqH+CRDgip+9Dec1QOQS01NU2qNuaODh
TlpLD+HMCfJ0RL8MIDFbMACKqnBYx8A5JB+bDlhnd2HE4qq8cgyhiDZ+0agDZ1HP
WDwtyqWGS8YtddBT088OT4jMXgjWAqUhIePVbu0oRBOtYm72a6iOw8XvJDrvlvIf
KGVg18QWo7itBXjX0ezCxQqg10XPakRwZEPVRanJUCiOwPkd7Ysq04IhUlh2zlYU
hwfPSQYoTP1u/2hFrz0cxkipXizqKmEUBg+BHPKckm3yiXHeHxnZRFIdSvaUNwpB
WBNtEJ/14Umd0Kh90NHQGiL0yeMUlkW5GJNQxNr1d95Pf9iYuR0BoDget68PWRdn
K0gakdSGzzd1/H7DI/Iy68vcX1udrUCPcGcQ8Gf/AwIEMZ37aIBKuNuWK6Z9t/+v
QbNUh5gwrmXPf5tAjorJpA1CCHOB0Eg5HYOhtZS1F74URmHuVmETCf2PYQ83cQcB
NcG/hMaUnG+sPVSImcRDcHLati00voMDxoRHXM6Y20JqrAETcHyjH6ueJlg7QHMw
bk/hk4m3IzeXXcJP6M8JX+Zvr7+UXDSFGN1fhexBTxixbDH324TnPWsxOlMgjSrB
H4gJVk362/XuHsEcPBHiB+jQbYJN3ANcl/xZ8HG3/v9NO4gPhKl41tv2/Xcu08c0
wdK9a+S4iMuBSzAsCl/v27QLeEasOs5dPnhCUcGNHEABjJooxhKGPQyYckMcKyCq
I+VS31sqeJ7oj8/HPWEdSKUi9ucfcpXBhy5d+Bww/bSZ7FrdBgeF9XPC4JH0rBLV
XEvNN/AhMvQ9vZtiwqyESk6x4XBIfu3nbEOAhGDcVw5OMhMVK9iaaafhJuuNzvX5
cIhD9MOzfucNLq98urxHlazyJjtjaoq7nbIkxyZYCaxZ0dayvHpAgoRjGktQ4mnE
FFgcYgLdp8gUmeSH4dVq8TRIx6oLgpayLOajfmpvoSlJAD3+nE05WegG4z6vW5AS
xPLJkI3EeePVWR21Se37BO233pVgVXcBty/AWOVNnlRecMRkbWe1LZWH1v6A94RQ
1M+t+IFQuIttBq8FmO8h7duWPlBGVsdYxA92zuSIEv25UH4xXRu/tE2QkD8ezkXq
2a5B4Wb4Q1VBO/aeFrESeeRj775DU3TzKvOA0q6604GYLd5YahmT5s37kghP/pTx
8vwNyLNqbt5OJVfSk+y8jEbyDsDJtDhu6R9yFcwjm97PsviyVKAv9QricgVj4hb2
RuuMKpi06nL1YVnO0ElyGf5rr67jALUl8LhJ1hSIYrfHkNeTgc7GHp2ax9JnDDtO
BSxtGVK8Wopn8z7jwz9/kM0lqfuE4B+PktmAGchZmslai/8UBHEiFZ7ptkavBCeD
LwX9DdLgEQqRJ7o1TpT+jfueEI/PPXUcUQTTUXAXf+aUYcZiK0eN4M92b9zqwCZ0
Ael4hufg1IyQdJQjdqPnQoEVi3tTciSrCXKInE06s63CKnrSnHboPgGp9Zp4SzH7
aNPP07su404h37lHGIfoul75z5FrXumzcgnn3Gvfvki/3IMnTU3e4XHQq+PVRGb1
YvORfNeQY/QwG26EjGaiMXvJLmyRfMfiuvS1bJul29jj3Bdm2emyUedmlay6Ifze
braCEBotD4HHjOQAj8OvhOdquRJGM0obDfDSWSuWTQ6uMDKEcTU2YtvWuyR5Fnhz
sz2ZEFgCH0xO1NS4WtuHVO+hwuWKMrO+i6K4TubjiWPFomBfNhCIzCVy4LaC+fmh
odgIdgHvx/8IYHTP3zTYTS0EvODQNe+NfhJf0ArONIPMoo8E6MvoDbOGEM7wBmz4
nQsVP0Dv1TXHNvJsout4Cy1gTbf7d5NwNQKEdhWhGYrKEEBWuhcYna/3Rw8Jb51o
ValjCpAt5u+eD+ghvN6EgudmESljj8WyDbj49JYFRlvMgEvWFy2AGftXgL2YRp4x
DJhXFICFpmEsRiOQFDJK18X5Qtuy0WX6Iny7ZKp1g9lKltpWI2TtQdbyj4RD0leo
Rb5i8XEZOIYhhQEkXc3PBTYnAn0SMzpd8rJDLIohWUlgqsjwFJ0wjVFcwIUETgnS
tdgVUDs+b19jMI7FWF8lWTXbH5SG8muXUSBCvnMnuZcm8cxIhj4zcddg4tzhIx7i
cOa71M1GV4EBEK62Bwltl2Uu7PaaAuGCc2XSVlsvGZDpDODkV9latOaL+CnmsDmu
Zle+gP1z02kBXpeEly9cC1DG8w3mhaBUF8IZ4ET+qTDKmAMdmdnN7wYfZHSqetMA
3HYE0erjFwGUiWAWYu7+x2TzLFAA+ej9oTpygWqrsrs9R1YRPaXll75iV/INofzU
KWTpxGb2XUHSfWJXiYchkdiygO5Zc2CsI/3plw17a4Vc18C0BpBrNaSE66gderBd
U7hvVKhLN7wd7MWnNva8Rptq3XQYyBDv7SmIsixu+GMItFDY3Kn+cFDVhNAGhrfT
nPj2Bzx9KEHtd684pnLn/sLiDAsE47LS9/XoGrPOO4sQZ8G/Abs2E9gZ0Blfo3Sv
ZhWGlh4gR0U3BArMxvqkTNEO4F0nhkFcCl4AJLOQH0uZwdUs05H95xvv2VfoiwI2
7knHXfQ5+qYH8kufS0GVu6/DSDvxisW5B8cfVONykV9uQo/HSzFbGMRYbwPYnpY6
xsy7aUnp5vqd36dDqSYtGrMkXtvOPLEfd2USgD9cqpVQL+GgpwXY307yFGgnknwj
AeDElk31yYic5dzlsWaRqTw1YJ+SLp+pPnbArq48WhwXQsMPNvfRp5w/zTK6ROHM
POmW9HI2gAW3WYIN1HCMJv+bPrKa5cpK5iRQnEL8u+XI96cw74AIQn+u81OXuYEZ
mJ5leEu14v+0qvjX0B9Q+HxT3XK0/qD/R85jMa5hM0C8V04j0CJROKt293vgHjXO
UC7pctzhyVyENNjVWikWBM9plT7cWHNSh5GmcmNJhrmWFsKF2IAzXFbByYYuzXmY
JGDMc2XB+uWbAK0155d17YL1d04tubaxHWo8nNqPhbXBucCmUjAhycDGpRHcuTNq
j+gwkoBpisGxfFcy9HZ515i5FUFlIwEH6LGozcYXM6BtThK2GI5lFIfkDPjzaeZe
eGVWvDEqldhDfScHHEWQJNq2E9NOqmKhaNPJwwXl+srHEjeVOrd2mvU5Oq4FVYvh
u3Ixmc6Bsyn3cAE63eV4dZIbooFSo1EJWKmmiwtqfPe8gfpJGiz6p5PkIClEHg3K
Z0h76I19Wh1CqLGR9ulYt5mz4e60E0WX16gGHYQhgkoIrtzzuU/2LTbXh7lYOVa0
QWBWFSMxKYNO6ez039Q70s2uTlbY/vsgtaYHya1M4dkf+ln8aEpWdk2ymHUD7aXD
TdhgWfIVIlugJ4s0+F6rh2OzEgKyAM3qgNqe32AuzHOKJTrCXGy7qMMbOGfpi4/o
15au/Fmvq0l3J/yBpht+0pXSL2SFZob9B7yIIb9AUmkdEIoJNs+un4uMVb40l5Q5
jipYYe066vfPlHUzhmpbRq1BOm2l4EfHkA9Wmhv6TzB/A12p97RiGVMWkqsT89Rl
JKsGE6sOecrCpahu9POgBV9GSUoLFFmPn4DmocIimHqYByyy8DhOOjTNp9mDskoa
sTS6vNlv4rMq6g/giBcDk0FMydRHA8y5cmvXclUn7/NpXWvZ4ls7JoudRehUYPpz
vkTGK1CkouWHbIsi+GENlBhqDpBqGHclgr1fjT1v4iA2iaCWq2P2WEeqDNpefFEb
23rGnDSwTKD0yUNPXRaBJy0MqlBRJQ7Z5vHjUaMBDwFl+fqFqMXtH/5RuTxNSvjM
rtBviK6cbPkyhDoHpcMpKIDLIgq6ktX5cXOpsx2DCCFWp43kaCQ6KWPr7YWQ0YIq
HrzJ59gPT2ku3mo9SWS3DV8pI5wttqcZPnv4pU3SLHrRrX3btUSgnluNO5y7ZcDU
vqcbzItHhsQqmoj5II9+KXI/r+k5TwKxxqco2SRX8bwMRJRJW/jIq9L3eRWqnP89
4IdkrnUQdU3qqE3xJoH3r7q2cYRSiQKZRjGj6ip/QQPAOf1iAi4LnXdzjRdLmYo0
WoAytvs9Vugi0Uw2UhLQuSiImyaGpGh21q4RqoSSUblzlo6P3o4kaYQlys3av0ww
GYPLeL9RxnyppkvqgSnqOkyzdBWyP2/8WhvT9Png1XyOiigljvfHuU2nNamcEm/b
bjRw865sMPhcRZEL2o0POjwzMhhMPFYTGvRkvaw/vvye1YSmZShb4uFQjy5ujwHq
DipU1dzFz5VbNqzlEmi35g1I3j64BAFArJlb1jPKjtYLLBVMpTh5f7HC9TcUUlQt
F7MMuzN+khKwl+YdzH3aOXrf2edPcK3vGoWNfZ2Fj0pCOSriETIKDZ3tcCORlpyk
ugApDNtIZzLetopfaAptuH57Tq6mx5MTaEIeGxzmyg7RRxhcThymt8QTOfwM9RjB
3kaccIqkfJaHHFpM0exvd5eZzU9PtAqz3QSpik1QzH9eaCTRqKfkFe6rtQ0SUFjW
Ks6qnzhoL7ZUeS67f8aj80u4VmSvucShl3k+Tz90cFecv/D5udnN5f+/79vu5NCv
FYksRAIzmn0/K+afuFdbCGq5vkPHn96/em+TVmjqwfHB+sYOfvzUKrakczyavS88
0ec6tsB8h08hu295VPc66sVs3J/ti2Ut1oATrQbQ//tTz6Ov1GCGijVlYO5cwv20
Rk79mQwJOvPFPGysk0gdXGyZ2mNWpdkB7Pn+5/zfEi6LDknskSC3onmiyiBhQfqc
EhLEtM5cq3oKoSmHGGGKJFmTYME2yZ9MmXBAxJLBUKDVjZR8ekI4o/zm9IfOPV5C
nLgEWu6oga5AEG2r2lRk5hrWVbBuQd7LPzwu3AM0bEjRRWem78fgY4JLw8F4MteM
IF7SmMpqsbgHkrEBof1RePTE2a8JDbRBm43TxUFTyXhABZXj7GIixEBRDGssdM/z
PVonbS4MRmXl024oAzSsG9XqdBHe8oAEewQgai5Tdw2ngv98MpNR0AUppcrJG72e
DatnEg/0eI6PPLAZpi6zILfzDXkDXchD4wciEGZufH/qthcppW0NpNJMYRtHLOSN
MHHPSgCkjOThpHmDn0iDT4+DA47Og66q7vJtq1Q8ZX1vB6lIcyvqiXPxDdid8ju/
B2kDqYnOmuFXw60MjoO12IyJmbpSdoy2YKVLykYGLpFeqQWyoTMGKix421DQGIWQ
//d2yjB+j+M1aYAQVEbVy4oV4l2+JticJU7nnfVyJ+zA2zEbmcgNO7khZne3bS2Q
tLEmfsw+2KhO2JyoZAy7SHW5v0nG4YoybmHPjmDp3el6ARujF4wI82V/79ibGMbn
fU/djLHs1T9vepzfPZJEIVt5nIyk9XG+hQ3oCbttHuDhU2qfxRxO1gm6wt99Uf57
6TPa1z9iH5Ym3zzUKQPxvhc6reHANDwQCy0W5STuoOtO+OVfESiUU9HZ+8u5WxrO
dIcb7BoUjxmpefv7Wt0ewRr4RMlGbeMsbKdYKmAsynnO9nDumsEmhrTiuVQavyJ/
0QzrLwTTNCYEpENpS1TFwrT+eKwfdnYn3gWgwQpp+u1cWQ+dhZCHgxFMtOfxnlHm
4AXBjZwJ7Ia8AUybFnxBRrJwRmNDbBFNIqQEum3wu7UMmH1bZVf1Hd9oDadkX4yW
NniOoOXz5vXeN7iuXFsu3tBu5vQQN+h6z4HrwYxUIBgTh7Po80T8phCm9/klQIVc
Ekc206ljXWJfCvLfUdjmJdqbbs74/suQdMwFaGShM2Xh0BEtP+3KJGN/sUMnjUxf
1jOuJrnZmJVk/yJhPu7nTjbt/wUrZ8G46JgS2aY04rtx7b8e//vWC/r6dtlji6gR
RTYsiDcoteURDtjTuUGQlzHWRDBXZ4BLI2Ly43WQy8mvsHZoFUfrLZYByWjeOiUo
stGeMS1THSGFpY+t4AfNzY4wUMZdE9g8fNyWwJu4uczgaaV5R1nd8qKIPMcMbuMB
wHgV9KByiMdODvhgrYQ1RWQhXcDcbWBxUg/PYpE9NTPD2gM7//rlxRlO1ImBHQyU
Vr5g2pVrHCJWPL4r4cV+kPYOOlaXc2oJDWgOZHt4K5hwntAkmCH1VHSP4Jbs1ztu
XZNWETIsus3+/W0xcOZtA9myeUAa9CenxICa9ZpNc+yV9J4VKSIBI4mx63TX+yxp
s3nEM63bPmASZos9wrOiVyaqB+VuWj9KW9QMzkDt1P0eL5+hy2sEVdudoXE1sI9o
D6NmoGaq0xqojCQieGXwideWBkZhYthGD8c01hC7Ub8HHa6q9EULitm3x2t5XxDU
1dG6mw8NwW36bGl1GYDoTbPYG9ut+uEa1U7mTgWtbXLJhADe7hk/BG67hyTtp/Xj
TdAKztyHwo6BK6kzd4MX819sUnel49E52y6aJJJN9jOmX9oRYA6LG2XHi5Ko+zz5
67P1fI7a1urLYeSWvTSo0ZDdxAnOiXyDnhzEgZJmUkcRI7KJO1pkwtzsZjVlKMNY
7mJHf0evSvk+bDUnw/bohgEE/jYSvPQUg/mwHLHBB3f1kS/5+Klfg/ShfNAUENB7
jQWJy2Lk8oJVckDSPPWVJwMK5YLwfM5DjhytRkh7atirg/E/Ba2SksibzMNaMcKN
/e/Np/d9WV+d8UX6/sUUeOxvEicQtBk2ZjStFKdLmkYAPiVG+hYHN2DLolTnD+sk
JxFJpx3F38SEPhLNs5MtWeniLSLVhtp5PffR/Vh0JvQ3zgn79DWXP3ONfLTgaKTZ
OnxpFv5s1YFAxpz6rcHAt9d00QSZ5waZFx4lXsNIfzS6rps62CnkDStIEQVhKVZo
1txn3251YjWsn0tARpgXGeweXA9UQTOXnUGmzxd9OJJlw2BN7U7Tg8IRNyFN59ao
J67y77SuoePO1Rxp51GBCfbGOWARbavDLGX/BoLsShJHYaJRz1FLFfpaLXdxyosX
tfOdJ6AixcmTsRT86UOfv8egty1KjC5YLQExY8PvPChSQa4ihIRfN0B5X53R5WDN
KWqEOqhiHm0szSqUr9aC1Ud72xsg4D3GYj/gOFMCiKJ4PSQgoZbzgkuyv87SOAMY
5tGqLargS71HQ9TXV/KmhgrkW69VBmTbFGgVyG0P044X3FCMjgURx/9b51t5+/M5
OWQjI/HkLnbS+Tnwp5Ty6tRt/HUIceRysVPEVGHZAGMvHLC6ZLwCw2QO+p0Nh11s
azOZ/WbrucygKxy2P7DeIW6aJN7We+tCkKkx0pdh7rSbUmzlhuBq0L018AV6dVrG
AG7/uXmo0MHXcFIjtuO3laTj2evxiEjIP/jP1lMKsQYLtOCMwaBPW8a2Pap+JAn9
eGQDH/XFFWxkqRAdwDogfJoaiIYx9lhnhAATU1SusQ1nsoO4akpxKqf3gWGVJOHB
UdGKK9ukPMuX506lKLdlQ1UGnriWjys3SrXbLo/2yICO9ARY9JPmAbqEmZZCPy3c
LYbnJihD/Gfut6iua1bX27kR9mdkQN9ld3oeOZ8Em0w9tEo82UyDeao421MKO1HE
DeItJfl+PH65ozYKzPdFNtJrXkhBBAgmF9s+tMzol3qwv4Bkc7MxMhZ3izNXXjgG
Wg6dLZrtzk7XAjWAXZm5hfhSKX8Zmmuc9x3jAmNmkwq0083uZRB7XcOnRBwPuY1T
jw6l/c7PEvk7dzgVWRPFxrMjZP0q78vqofBs13quRtFDRKtpcTWbc978zB2VDp82
1RZw2iUGxo1YeQ8opLM+/XeOtUxoJWXnaGHao9mpb4Qy0Jz4hLLfByvSmRgs65vT
j2HuoEiuGsRMcti5Lnsgmj0+xgqgGJ2PtvArmzy4tlT4rWF/0shWbq58kCP8EKJJ
4HDBR7YvcySz2zNjPT56K9LA8gPFivuMhD0o2CskeRGTHNdISBIpltPascAJdmPL
NRFy0hhmDTPpi/Y3UQ9El0CzcPCvAkqrvJwbJ5SbyPEXfeRRTappNo7PaPr+64VK
/1q3kuyib0tpZ5Kl8Ty1ENKiAL4Xfm4q8UwmuzHQT3SdfWeJD+D8acpNnn/64G+d
OtY7gY/pStAO1i0oxuTcyP8ROEhFMbUNRzX4yH3zCMTFBD66CyhCr2t448AsvnOP
cDJl+M8bXPzRir4Ty/n07uPHABFpB81z7YfNdndNysIHaStOLqu+EJXaY7bkzE4b
ZedlJ533eKa58fDTB2yMr6Oxybe9OIx4VhTqemVw29PvQTX96FxB+P5B9VOCT8OY
6Ogpqcx0oVJNY3e8K0drncOaxdOianixtcrL3k0KMQpF4YGqUy4X+DBE9KUC9C5X
xDfFkwznGKX3/ZXWPBylTaKG5Ji4LF1v6sD4N9JAqqEcGoQehRzjbD3Ciq65pomE
gWyHi3IPUjJBQDj9kgE6VylbUDZVGLWzHetvHwN40sgE2oVsl5nSKT0X8t2UkLl4
nDeLvycVQ2Lmm3q7P65enG6lvhcaGb2blfZIpVyERBcmXHIgHMoSUxfzBH6oqbWJ
lNDFvRdgr/fy6exqU62SLQchY1nohk9+h2cJ7vdXZ9A8ZiYx84FpjMUWJ604VxfY
H+0UNw7Li7BhSdDm2TJgCADXRKy+LdeUWYfGiZNloYXliVJ11hUPPANw/m/oXyGU
hwdYlXcQc+NYHChPu4FnPg873SKAcsqoYh3gD528KoIwwiBqgIBdiFnbXshLrOED
WWB6pkg4ONdtLDLsL6f7m7lQElV1ZTP0ZNAXexh2Cb7Qg627yOJVcqiDENAkHKJg
rRiN0aVyZGvLPQ+DSBO0/ggRD+J0VAAk9l2BYI2PM9qyOMG+a3yv++oP0cDk8lbI
GmrUEyctQdlsj6MIPw6mCckguZJx85jYby4TQjx4JbRpJGoLc8X4SVnVjAmz/Nir
RxDUO6AGf1KO4IiMAkLPmevGrgiNdzhUhcIoh1gYjpH2C7vI64hpQjQA7EyXdGtQ
Us3trqAZyBqfKIq9VU4lNuzkn6D9r+40KNU06w7MvwHqZCgI5asxPpLwgJDw4XH9
N/GLwlPN10HKMqvcnE8sgAJGn7j0PGtkUIBAd1R0pGRctQc8YeSUojbY7Z/UPHNu
j1dJYrjwE6YTxC1FpGM03hQvKk7sogEQxTYlBcXB93Yq9QCcgR3iZKYc48aG/q6W
XHl6Sy4KkWmxIE0xc/9Q/mmV2YwLdi0wl85tENbS9p6qMR6EdZe6PoBYDuVEi8lc
qdCOaSklABZhO+N6YzXFW1aXf76Tbe3WUdoHVtSYbSU8yDlemPF2jMeABYw1V+zr
HHmGFIzMhOPTMRovbzqCOWsbXVMDF0BBSLbr0zcfNKnlSn8hmFfPs3g0hUO/1G0b
lT5EhJFHZuRbLgVdNQJQYBCnMK0r+JNRA4BLpXoevjXxiQ1y51SdnXrAstth26jo
valmFFN4qJQNeQA1+I+DVV/rHZN26+O+qvNbuIdIPKami2RvqXhLvBpCu2lsofQl
lUnWpC771Dx+rR23j4dtYs5jRO+35d7AVcGOq0bOxlDDXhCzlKlt/Otk7scojyZF
MP28nVHCgNu7uBx8M01R1/h6O0iXcWlLKHHv+BW/Q5eRqCaAF0bh6KIH01pGLybn
gBlHEU0fTuA3CTgbq5wkxP1q5tFjbqGjDOnga2b5WMpys44X4iAzTRQIOo7ndgLW
+BJX015er2ybiMbfpH6NvpggEnEq3AFnxpZfMQVVfinQMZklteXId+HrnKHQXYK9
ZyCrygwwzy425nsWbNCUWyaFN5tDfco36Uv0jG5DEbdt01l0oSpH5GEDPM1wqlnX
aF4vcUD1TEslDkHp+MxMtT+NWLCOJ+YDqHgHgDf3jeHAizXgISGaTYyv6lIEAxr4
/N+23qA6OJ03R723aHwiXrs//yKpSe4+iapY4muVUc1Z7mRw8IEx2yhMoaYeo6p7
Ut4wIn4/RUWwRqLfVRfwI1xBSX5BaVPSnhmZMrQby9Hm0xpr6hn3cKzaFr0z2e/j
2oYBcclVaPxKYwtQHvdsTmjSusBC5uWsJia3DVT7bZ8MASxDFak/egV1UgSPJmE9
Z2KhTTVJEL9m7J5+aDOelQbKrKQnGwkcES53IfpJwCjuUCSN5LnsTd9w6/OZt+df
oeiD2MPPy3wB6J6h4uM9etz1ZKBxegwdipIilLVvQQ7MruRkkYMQqm175yNrt2gr
L6EHOGcozsHiSrUfdzkvn9PiOmWSjYHWePlBzwxjmpJa7mwOl96bp/aJ94bSWBYU
0Sf0LKIfHajEbZHjIenFmx70HloXuDZmKCdZqoPsu5+uFhyFe1HPc+jei/iOQIzn
4ByxfA6StJF3Dth8cRsGBBi/oxgCzQIRr5jYEB3I3ZXhtNfQ3K9PMd9EsWVqDMts
z2XHR1DeuvnDFI27wBcsl5KMqmx6aBbquybRcNhkwsbZA//G+JPapPDYXiaBEXP8
1uexNW1h5jMAaf2woQN8q94cIOunT72oMUXFd+9j9Yt1eQ8k1VIWQTzir3/8YHND
yhn5mJ3oZ8qZoRWQsy5udaoQqaYT4rJW7M/wv044n1rKeI5m22nGkVZ2HKFwRBok
quEEXVIS0bzEErQI2EbuH5o+4soGFnzwrkKWOTd9HE9h78sOTQ/Qyd3U6ekQYlLi
FCe0wpk3x2PR6WvyaJ0W6JNfacg4fJdWJthFebAfcteabQ8kzupexom9vz1vzaoP
eRWq6RDYtRoqkIy79rth1fGoFbcwLV9t4Mk3fwuyHYB7LmpbioptZB2fN4F4SAKo
v3JeAZq8856WYZZuWVdZE/Xi4DsNWs/086W6krZ21N8sUgTmChSlO1uv96+VEF8e
+c8xIS98T++iU/3hSEcs98mlOG/f7tByIexLhnE8Ue2y73joVJIXP0oNrZL9Z469
o8ZDzBdeAPi5SgvUxLq+b3qvu5VuEc2ti7JVlBWFirfvYTo6ZYUdU//4/AKAeQsb
DyzvJ52p5xSwyWs+a1lQOGjzGVH2g8lsEfrpeQZK2SPLbrRJo0PILsCXViFBh/Se
RWobFz7EshnEhy3++Ds4r4JtmSeL4nI9Ie6UFvX3eZnWqXNIlWaflon6U3p+sF5X
cFj4CBStPxuryEeVj0g3GdvLqutijblNYVr8+eE0924h5dQ9TQ54Mvpyw3vRVHCC
vsHt1R4pKlAW5K5zSAjyCLPbqRxkFF06N46rfjhmEstzqlUoK4UUC099F61+AGZN
d+cMODMMEMUZLB/7kOxuX9iMJpgx/2YygUYrQODQ0ld/Cs/jc0PBDX9FBahOasqD
ZTg6k5TIUuYtHSySd0s8GGjE8e55uRQ5p3j0I6LGaKgohXua9kcXVxgRLmb9IjDb
cNFyzbJICN4bPecnxLcxN0L7dyXU+77mJTs0zJIufDYL6/vXhx+YmuYL++HTM8en
RXT+PbM5HLZYxjgeOPZFVZDkLDWkuHKlGm3L7TprfFpd5vpo+KLO3Yd6xMNcQH6S
hBlb/7TLUXvgUXh/GSKN/UUyreWAPVSviPyBgjiuWDWny0Lz2ZHP77Wl5QqVVZ/6
NkXMl8+fkpiZwRrPw4I2CIIT3D4qZb4btLyA1Yk6HCSo0NbEDoOKv8gAFez72nAG
ofN5CxACLdTUXqNUjkBvTrviRCBW7H/PEBEViMFN3xeTVTMaxKcsfm3IzrVD4uWs
nOgGl47sTrpFXtklYjoN5LFkuyUSC5uLQOvb7YteXXscSYBoYFpOEkJytZxu+LVE
CKnO+S2oTVjEfzx8JtbvkkjTDMfHgbtTluFJ8aBOVwOYWxQu2y0N69zjeUMTmXVs
o7fSS7EWp4lo1Wii1WjxdsuXBvHu2NJG/X6Ka3PtbQLHXOSaDbUOucLZx+z540IY
vGR0HAD8+X0V/0Ma3DCGuLbnbAkd2eHgVWUlVPcWaNK38c0blvoP2ZKjYNdqlzYp
cwZDujB4hVLMwTSCMY720tdoEmz/iYpbTuA465YYC8KjS6gZZHwDHi2ol0asW2X2
8T0as0KhdMR2YZPIXJBwNFUS9rwgvObLqoo+V56jzGkXzZDzvuQGziAn2EPOEFIp
FKXMLefzudONAjAGatB0dZLIjXzSjdIUKyyLYxDe8lyAFKSPNfwt1ges+aeuxWYu
4uW6ZmsVW4rXr7FBM5OrZN+4mC3+HpXzgdhzB3/OGAaw4WOverKOnTxewgpbjdBm
ux8nJCV1Zf0yRa9knLAfOsHZARdl7v1n2A0MzRnx2Oaii/pRX5O4irAygySBrqLB
dPcA2pUXdoFUsC5dWgHeWecP2Tw12mXlFH9u6VhmtZnj/27jiGMnwWGdns9TpeX5
aFWs+EFjWFFRtjUrg4pmByGxe5r0ObpCnUy0akFOs0SZB6EVnh06k0HfHwD3v8GI
KZlM94AlVSzNQ/g+JI62dPxGwTSbVkYndPUBZsQxXHQT0M91jKbFgZRIyxPEa9Et
Ji+zdXH0Z+qP7PIh617HJkrpaYfC4WWYDcfaKOk5ViMFedIGgxyLBiFXjfgJGZ6W
0HImbEbE02+Yk0GQUFaIN+BBT2GqOmQ/DQEnZvyquJrOJX0eserA5vrnoiSCI6o+
XgJVGz+8RAWO9rt2tWmjaDox3YdOLWA3bxq58LonkHiL+ADWEC6PyykKtpp8golW
n51qMsOxztZyiTCDcOAEin6NaIrWnrobMPGzuhNMtWFikpe+XBaT6pa2Q84rK2QB
uXYQ+NJ8GL/jwfuHr1XXlYPot0mlUtxOGwkTLNd8cTmoKQsi2ClcX7kX9KJICGXL
+S26M4BabpzMdf7MUE9gpjGKv37dEXifuu0w1yuIc8TaBN5ydCB6CNmvQ6ZpMgn6
k/8UMHFXYg+5mfZWwwDLC95ldT8Ddn57AXJFiZGkT1mqzB+14miRJ56Wa3/hLitu
OthVC0A4CZSHUsnte3OC6K1eq0MmpdPiOyRmC3iB/BMMK1Evlgc48b2zE45vQzxn
wRXjvQPj77i+yub2Ny5KPhLq6sMSYDlG5x7dZOHOVsOF+Fp5jryTG9Mqon9w/L3H
H/Oisk50QarFAjZgx9EySoIt7bY48QuoHNZbvgL6b3FgN+17hEWv8RvIzNlRAWvg
FY4gDMHGaef/SQsER3PyimTxJywOXHqU+l50TUAuS5hCuto04mlIepEvcaEz3NuZ
QypD0KTFB+st4M1eWCzDWAHdmSoQ3fHaXhywpRYo3cRfc7Uc3M5PtT1Sy0cDZIEL
79zTKDKqzhJwt/kMyYJL0M3hIlBQn7yVBctw5lkl8It1WtCcD3OBdv/bP5Fz+0ha
xHrRWFMi5CZsRb10Ma6iYoW4tGXsZRawD8h6APWhW9Uh0sugxzEjpDVa4kvPUd4m
OYGvb2IGjsQnl22m++aDQ6Y7QU9S5pXZoZTj3yzsjb/vntr6yKr6qU8a5Ywxesfp
a/wzZuB8aj9Imd0abMFufPUeaUwnDAWltYda43meYVcoZPEARbfp/TiDMzNKLGSR
6oOY6usa6w54i8D3QB25ascMyCy9Czlue1EgxqvI3CufAjaSMfCU9K+QP9MtwkJq
VEjcn8QkwRSZ6NkqKQwOgZ59i5Hyw26GobiDI0CyA33fKoxEqC9T1TQLeBdsvFm6
t8edta+PF2moKw/CsM+NEFgLztyEFvkg+a4asuhcwAQ8QPbBb2/1A3SeN/I2egM9
t+pEENg+DGez84/z9ePvqtNK1SwyO3sRpXB091/l4csOyz8R8cY4jj1Ir+QDGe6B
10nKT9Sjqn0St//vutGunqsbXaVYqpSuNtzkMStfIzEaP6sei7wKJNcha51XKRWT
lbvEEoaFUk+FsLLnZ/3xxd+w1B5/qvdD6KLGRFtLzgycS5EcCOuCK/OOVbZ1LBgC
oEOAu3cMx7Rb4nprmFBtG1h3Y+hVCLEnlSS77UUFSP86e9M1LYCpwYOrLCaVa4YF
+Hxk+fKMbbdJ/eBsRwUfv2yPLygt8sMWVyhMyP58Dli6N3NjcgCfxcFe5+nQ0yIa
L4FTmQRDiypdDyw+ceJ96sMCKxB9MkRGeGPDsz6tPtgqviJaAnea3eUnid6kY2Gt
2IIhGEyMdv6EHIDHtu4jRgxqf2/bclpxITRtw/ViaUblo+YMSx8UomBGy8BIyg5g
R+eYXAoU/7FuXAU6fyVL+hA1cL5n8AI3AE/eaKusb/9vYRcm2MQxOvESWaXrreVG
HTRDxzuSmLsi5gf/XAJGx+ZY3mmiSCX5RlXQmkMC8iZkEUXwrx0VfqxFYi4u2f0h
bCeYkVKmv2WqV5yHt2D/EsZyzeNNmKB31yc/tZOhqUCJvRzbLFOh3R5SCOdAT68j
vfDJOcDQ2gTQrOjzVNaPB+ciHP+czO0ORc1BD1IN3ZmNPrtT4sxTorlxWTiyk3hY
+1o3nq8DmUi6qR5gY/nXqQmYb2SvKrt4S7xH/n2avBHI68A4Z6jTzRPgSSNCsAtf
DkmKd1FY7W0lIJ62jAm1PDuUg50+og6RdxNBJSCfHEWSGqnoqyY8ZLKg32aJjOYQ
WZMlCxI3x0bIq4t0g5y3ORiguZ978ssR9aHKlANmnj1erkndZdqkjT2OCRwmDCpg
H28L/ZyIheqrcpkr+enuenuLq1DFpNeQh77wTOZDqn4sxwlpOo5SbKIb/M1V0z0Q
xc14YRxrj6M/4EYtoFDNHqIj1l3Q3ui2oAdASVzZZwIRzQFY7Uuexzef2kwdqRlx
lU/T3H+aeAp0PLQXFPYTGU9paE8qCpgp+b6M5uDzGdx9e/VXZm7ESoqCoTZsOTRy
Srb14BH+UfIrflJ859ZfQVLogs+ezXD5MF1XqKe+wkART08hhTDYAYyqB+zpP5vW
7MWEIyFqHA//FSPy998D84pAXkW1wjE+aINKn3JqBhf8QShXLtjwewuvDGt4ze9k
gEBTDS6yn7jf45DvXcI3It60QFlc0cTCd8dVOIHw1cjeTIMEZMY8fYH6xDgqiAwQ
7F2U+0AllSpLuS8JmT51BJvsuq11cSOh2V+vo6du7jBn5VB+YQfnRVdf+n2s5/0x
uqPKNx/vgXUu7AE/vTP5zEy0dVz5iUQG1Dyi1debUX29ddkm6KDs9Roo2wEvaRzj
6ZrjUWE1tBb5+FquqSx/Yf/3TstaDRfePhFrdw2k0UURn1ZwnSyaORDX3o+TFNs3
zxRi1dKy7Zze5ORamG3UHzLAwIpjJO7PqpblTXk7WWv22qbavFHJiOLVwdNAwmsn
339+MvG+aM913MxVcMpJllvUiwKB9nWrUIG/3KmJv+h6hkRis4+OjL1Zs6iMPGsX
mIEc3FaFqpbJJW7U2atmM4rKY0UTqtV33SAmDyxaOl04mw7hokI/2aluH4rEhQlF
rN0GtseKkiulXzJRXzIahoVHsVu1bIlEy6ybNVREg9pNIfaBOTnEjXVzQCWYGp/R
3MX1+s18Af/gPFMNFFE29TmUF7LHCBmBxu+AaN7/NDr0Mddcsf1M2gFEhqRcvB3c
dxrDJSqotD5DRUXtvv57+GmMEhrBAuBksrjsEIJo9SXGuYvQwK0TpdNSqNIGj0jc
dPvODxvRz6aekQPvYGxwufzo15uRH/DxUB/CWIDKtCABYS9OgcQsUeh5YJBKsPas
K2tdJoaWzBj36s0tyv0Qip7UOHKXBodCL/JSA5VTvy9/HGimkZ1qoUpVyr5OeC6p
WWSV4HExpBSVn3HdKnKC4DiyXWrhap0TaI6FrwA4C8LFWYXBjGl09CC7ixJZmdxl
k/sDO2y79anuq6G0qgbIpVSja48oyF8889fqKyoWys3HvnluOBWO/1ZhWUEKUyb6
hjI9daOjvDD2GsNeIn5H813WiHlICgGisi+3XcCVvqVJG5bFg9vacINtrL3rWpJF
t8im+DkJob8DP8usObo2SJlLBouPV7BtsNT73hg8t/t2TGpMAHLc6A0EQoqlGy5T
ov57uwSS7uX1VudTWkUzgONNqAeuimv8P7jSgONN5GVOWoDjseDlR6aKMbxfH8+S
TDgGGPckAFNvaeGCE15SvTTJtpSco70TilGfqbBkxNlDSJX8k1l09NG5ObIix/rQ
NxrMlbSuMGHJAHEb2G7QbDPcucuOp8/NF73aGyNuCZaAf/bUZEbL6+9EcJ/WybLa
+mwCDmXAM6h3BdwyYn1Ol2kO2Tp7G4Va/F7ANmcHtUa1+uYydVkj68ZKh45NcbWF
5hPUa7ec5eWCv2LR6Bd8ZdMCK9a310zY+EsZE6Cs/9Vn4WtpOYJW+i+AaBO+qgEx
BgBovvy4MJ6B5lXigtaWL47dQU2gSuctjgj6P/IKgom9CaBf+/D2d03TpdbPeM03
5TPP0eSUwbl0Q2V2PIMJ6MluK6DxrByPT0iacBfOmz7VEl8tGzRk89X6wG8Nr1Vk
RVuma49p8vfUKR1v9BsNBvxK1rDcyGx8K52QnMeWLMP6CLp/pU+YUt9e5QQYUF2V
0nWY2iymIPtm+HwubPwyo0mqpi3wFyS8baEbkWNUnce0VUn2SHRqxYAWnfQ635HT
NYtMoLRL6pP3I5exIyAnsxcO6+2DlgIPE1FBM/8EQOVf1GBMI6XhPcd0o+Is47mZ
ggJAEg43MdT4nbKrZiYNG3BVpMP5A0el6LO5+3vAxhivDCmqDfs1OFM1tb8R4psK
2t0a/WPHWTk0xl0gdeR9Zo7ZKzmUFNc9a2eMGkOZNsv6+dyc44QVDw8hu6IU2RHo
1luxgETVMIdzDfnkFMo2hN6TTCb7LRsLkKsaBF2b0lJR19Ye4R8oxJnuLQhFf3H0
HTi/THzN1k+gbgjsqIbUzMAjvm6dbp+KhqUlv5EX6SHRms8+hmXHbj3AC2pF4gy3
tcg+JlkAQvlfZBWm1lgDwPqhKHNePHDmzBob3Unou8GVEJpnXF/fIs1H/yA3iXkb
+WTvm7TNkFePvOv1LbjiBSTeYNAMju8SH2NRvpCGg17P7l3/7ZKtMKXq2Mj02S3V
biPEGSJ5fG/Pk27Y9ZlNG31AOou55M/iFShQZBk3cHy2bYZMHpd7QReZfB3Yk4so
CpQsKn88qEEblpdxjvZc653Ggxg2wHZStqO7Zxh8HlWQyxwrn11tbXM0MsVn1MXC
dQ5PgJ4kFnsgiZ3ELQKtie40GdGP81UDPv8Jp5MjFb/oygzWdxkyWuc8OPuhSwg3
XruQnnfNkMGYW3WY6EMhNRwAmcyE+C2g77p4HmbAO/vQ9VbFiXwJOdlKPHq5ZnzX
e1oG8J99o13ubuvchL1DJPuC90ekrfcGfVDX2UmFiVhH06DIyOaH9HiVzt5FfLQg
HQyKB9yYt0T+Zfj5Qrxdl7BHwger7omOKNZUVZy10hpwgveW0YReUd2GonZSQUt4
VxFYZqdc+Kqrz84L4HDuWRz0oAVu4nbv0BkW0MfUYA3oY4A7V+WcveaFQ+/fuT8C
PVujQCE4VvVAzdIrVs2/U0VmdbuQWBfUMxaNAwlHT0uLWY3HsXy52Mg/5fw/8N6C
WjkVqx2aC8uUI4XhfOEMTgy0bm3prdBFLnmcpnMD5wgGefyWbb4hEhNzp28mc/dq
qxFfyEGYHiYAHvIhmr+qt2vpvcQt4pZU89bMRNNOBJAzPYKNjbLL/CEtHKAZ+RH8
zBRrZsJv+rFaKdjVgBNaqCB8HwRc8btcD55i8Wsv4MLhB1svDJvXO8UTVqs2zCbv
hmrhs156IvC0nouiU4vcHFSjtXqGTKy7vKi6Nr00bdhtBBzrudwjZ0O92pKl9mOh
6GPOmyKaP84Hiu29xtiEIP9y8RWyM1E8/sAP5onulNAweTcl4AXwmfmTHkQOeXcx
nQTPibzceKZNgOVDXvfQDTyi/yYZlzRmHw7R6FZwdI4bkMorHBhnE2BgbFbmcxhw
4OL6EUeL54LXixvszfzCdbUnbBKAkSb/fBL3uDILIIQWSlOwoUKYPsfPMWkWXnuy
Ww6C2bg3SCOtrYEk3uw753U5MjpXT9u4kh8YDEmmtpzM6ErHyK7Qbeix0n8qN/QR
r+JkmEfq5+rpbjexwG3ixtLu49gBLEba8Ze07L/LI5sbJQLfPIwze2lcEpW6dqGB
MTiMY/8B1TTa6mCMQZ7xWF/ej5ZGcBeJnlFLNwH/DuKLH8x7eAlpiF8/0KkvHz+2
q6FexuyqATzKHhP4joCMOU0g3+eozQGJDWll5iJel9w13/hefMeWMIlGmi9593Ui
fwZa5A/8f9T6V7bCYc+krxbuha0QAxok89qnE25eG3pJBvU+M8XSQo1XhKhV80Pn
WvT+bVbsYiJl1zopS/2vS4OK3JSrhJ44eUHGmLtCIIadgDN91ajpteaUV0W5wIJE
5YHl5hvIeNJqBHFEWVO1oJ0J6S51fAa77KHIZxAKB/K4kBjaZ3qRD+29gUoNV+O+
CCLt5RmFU1MNXsfbgMT6VfDDjSwMFJUdfZrLgiQNZpa2UKlOTCPMODXyiae9/lg1
AaZSq65mFmuMMbYYA6U7wLSln6KVY52rk88girTlyQnWNyzik8q2/Yri+0Vcq4MP
9cnz0wLIU1ldGYdy5MwDQcgcijeX4fFMi0kc3bSohCswxroRZURzxAtl6vqM9/vi
ikCb/en1fZkKncERzCT/x/Idm10PY44wV+WK1iWiP/vtMB6waqJ2iQ3bFRnKUsH3
cGXW7WfhfOr1BL8Kc5cLoZ6+uMzduR0/nwqDNaVBLHpN8FjB1Lqym18snKrWIqlV
3UWN5NSdr89CS8eIfZb/ogPXvGTUOccyGr3OeoAGCrhpJs474w6JyxZacJUMG8Vp
wxtdcq17yPMnIHVvcySJIQirCDXwj0fC7M5GricfBdP0VCE1OURRLe1WAUPyVSGr
tmWevosWffkS8FKdlFBJu9I5XjeraZILYFfmQA2ahVqxdQsOxxOQyoFfaoPg0RVF
K1nYK/3HriBnezNYcwpH7dwyQxJDYbKkvdQ7ukm0GWjBSANRdwAC+jDmmSMpe3q3
DLh0fjr0GohFmcWbYYR7AmJbHFff9S2JPTGVSoxpZxxdhWh+HOWRd7TFjiNHc5h7
qJhdktEvoGd2NvB/8v57De0A8hxjiZGBpIopagfpKjrq2Z1/tONv/oznrTp2gCI0
fycHztMehjtQWd+LidRrAX7wa3G8oD6OyOLiu/SnJMKKLhFuDiNiHLRWU1KjvJEV
bmdeFSJt9Ut9QCohfjLR7oSkiuS8H6vN/5su7K/bmdZgVeKrTK4obpi3l8io1AUl
TkEC0fgDh9mCAK1jFswKsRpkMprVgMusMaXZE9xo2G8PepfhGnApTgNzonWqDWxA
BkwXWuMSUi4TFu7yVCvkxPbR6LhJRSB70bOQU9CyVZSZ26bQYXI/xWHIUTrhZEW7
jO2enCgM76JX2WTjK4WXoKhWKUavQajM9QthZVYuTzRyYGvqtzXIy179azOnY9oH
ffrfFQVcE6OONWlU945zEQCxMxh0GdUAfXHGxZC8fq1JYcewHU3ExEkjMpScfC8Q
l75ioNckL6cU48Rb0KARCVer9SoACbZpOrT7Rbvn7P08+7KrgXHezbJ/Tsbc8KsG
Xodq767SGAiW7TudB/A5hHYn8zvqE6B9h3r7S5f9cPlBYXwB8T2zfzOb58gGSRom
OUOgvUplJXkX2VNCe/FAQ2O/uvdeOQieApHDL1kqg635MSv/B6+Fv1QhHlDilTWY
M3GQ2pW3u1T1SOeu6pqjSBpvLkysS/SGllBS9J8JvKlP381/5oNsRy5GLK03DJjt
S0hTcT17DeJIIv9VFj5sTDljiNC6drLFPep7AphDWfHkjhndG5X+39ya8dGEVvyF
QAPmyXxtQRIKapI/36ZtkTcXlcoiBrnP5n/I1VibaeykeQ+VBDjshS+haI+5fq/W
HUT2VBsQ0C2hkn2A9Es3iAfUVMtZlK2KVugR536It/NjMUd23rh/94QYhUHm4weW
MK1m8QiPCDfSOgY9qrSrJEz/wp7II9d4kR4+7ZdXweWzXE0IvW9tzOycW/4xfSPN
Nt/CmKXSSIXtFciUd/mBuo6n89RK3zwAvhRnaLec6MDwov7TyexntipDUs9mNZur
IES4/oVK743ZgdASjIJoAE2RtBmx/u2QaCEvWcljAaGXutey3p0v6Io3ePZRd6Lt
ZcNMYQCsRpSq90IP6Sth9bqXKRNnvEhMvIQ+vDKZkAqtcG/6AOnu+yx+yTMcTSRG
wt+/1WlF31cz0teXkiG52ANUOlskgiv7ayXbMO5kA4tVaqcLwX4dMyc5axnLapTK
eqQyvB04e3KAE5UEouze6Jwm2IcO4QFZ/H6fdsNNVH/NeLV9xitrqAAKXv8DgECh
NUNe4pKF9dbpOuX4SOuRWkl7EXPjoDZoFTiuSk+mHu9k8TQhgHxiH7l9WkhLjy4X
F8LW3D/YsA0ZYK3zVxZzYidaduNF1SCVAYi9R6kPzxtckaJU3m/DQHh/dMiZK8q4
0xT9CTTdQXIraL/TRyziJviAxY7y2o64SVQ53UuOHaGwr4ga8wlA4mvhxoytvf8N
1GmnCUWepilYFGxOUZe9MxdHCXXyDj4gVxC82iD+lJyL5ISAYR9KXCuepKVn/oE0
eUptywUTIXr5fC5U55Ubp0Ebl8ZM3zb7cPUSZQlhrQ527Zw8Ao0lLUyIl1czdONG
U/cV5HByI0/ZUa/PxF20pvVK9IASO0EV/1BO9+tT2RXUFPn2HVrw+HQiBy2TXZzc
miBa+9tmVrirmFzNkvWVmZTyqiNKS6MrCnArPsuQrh1vijwsiOZYyDvK1UOX84w+
HZmjc9ofHFZN1utNJaCdI1yEuiMuUDPTZ+4+CMUR8kFEadJGyAtvzfL6xk38Ve0R
OGwFunp+VtEMODMVB05NeVsMR11wzWc5Aigjd2oaXv8J8x89Pq+czfH5pFmSBW6L
NRf65dMDHn/EgZ+bJ/sX4HbMUnxAJgPOoktZpND4zdsqNXAEaZlvDsX9YAGAojLF
JewZ0TJ56gm3hkTASm5rUpjIQeOzRsfSByt8z15BETDnKVxfnDD20tdSCpA0kUcu
09fFqTmbSmO7u5j3DCjjTWfcenJZ9PypCLOnYVN+qtoMr30+WlZurkzz2kMrlp5R
6qrroRuYgO8h/Mf1rZmqVo4JI3HUDfxPrxVNNj5cF8eG3UxMzh5JeCo1ikw6mrwN
frfWgYDV07cRhIgsYpqQU+PuJF0fqlbb920G6WP5kLXYBDCadTPV8y3wr5i+nugN
oxlVEX9tPOsXHVjbgAimAv3Pyt5acpiVdBgSI9ucnPVeky3AgWU3A+ML77gDIDlN
4KqoQ4pVA/yr9LnnbNHXR+c6UJ5TGiWw6BSnblS5N+6YkMmAArNkYt4e2lFlq3Ad
X9vwivuzi2TIqgo7lrqBGiOqGWW1YhoGIkA6JKMmQtqXQ7vyLjs2oI9P1QxlnMOb
tPAqDXwNZLTHqa7sx3Jrwm1tVlAybgUbYgXd/+f8Z3vrL5UeqPoay69X3cjLJdME
hF5l7ZmiX4qwm42VKb/qydw+7Iwrk1bgCgiURqgxAzv9QCWCyAxEAUiW2t3LwOn7
Vo7EddfzS9KXunT0lfl8dhKlUWOLkh0LgR5QCxQj+WydFSvbU+4VXpf4K7cjLOo+
VLbIAcnVINaYU8yrjJRL6Wa1FCatDPRRiUu7pAZcFLvcmjltNItCu1f/W5G7uiA6
E+Jw0oWGMs/77+tFdriPXHBrHvIjf/hiA21bJxFpsWx3QVTZiumXq7wXx5kgqFQn
RoWEgLQW3IALYXsmBmZ2mTgUZ/qjIWNFGgDfD6NDIHmuWPa9/IhrI34v1/TmelDB
yjoiIP1NVs2LAFfo20LhNaU4Mgd/QP5ugCEAsXaIwUPG/Aj6r2a8jifvqpNnolLi
D4q8BHs97+IWEtD/uA+xj9Hq3r5/S0GbVZWLFrmXbbeD73iRroO7vEE9ydp4PkcR
vY7dUUMIa5cvXI9i/YBjfCiql4Ty3eCQbTEDznJINjCtjUCaI+Z2sd+iqJSPba/v
9ADH4n1vWTAQUtR0yCEsH9AIvQjvIu6Kz4DVmwGZy6c7sE1nYwGcK7IylqWzg7An
H2KQW2CthgQL3CWZrezhHjomJ6h2mkoguFIL/aB8RaSnfgKOu5NuKAYn5g9R3nyQ
5O4/hbZqxCvrZxKcMcivjbc8IPRnuf+qYLFrh3s4lfeHsNB0KN2CUDztM3cF7Pjq
yTxIwdOWMxZGI903QXfyQW2l3TdZxenAEH3j+494S3wYe69248bzpXGVye1traps
duHnJZqvLwMVKC6i2Jdmyj7jF04ms/fmygZUjAl/p764TNgu2bfH8iQ1jZ/AynvP
2bkg2roh+sKricoQ/WM903c8eaBeE82Q+RMlHzhn0k8AkU9nNnUm0mwhrK7lP8Hs
yRDcUctcy2cSerOkKeucrgPgmpHTaP0usJlSUgQF6A/RcKTxmO7GztAi6qj2aWw4
yqym0ChtW5c0K1TU2HhmpHLJbS9u1mr5/E3DZ+EZQzEPJqseKk21OViHYHVeMzzo
ZNzx7RePNRs9OL17QGZuvNC1xzCdBmD8RcWN7tWW0sIP9+k3EMqzOH0fzKHzJFt9
H+eAz8/W5eH4BSnCFqVH/0ZmXRzavq/XhH5yp+8zR4BR6GZU9o3XoK+d50iofQql
soZfB2EBKO0TkElhK3TsCrNThe232m+GTbgQVjcF7FPFRJV7bm3T484EcsaWAn5u
iNcvMN1eCHk+/gD5RhLgV+MN/WQWxF7uE+uqVzMEX2zFbRVuSvOqBORfxUGOlffr
CLFeyRck9QZc6pFeV/rNxFpxWAZ+Yox02v+D4Ha605WAIXgIgaCwChPricRD2FxU
/n5zXNUtnorU+dE8mqafEUb0MS/o6sc3YU0ZewWaEyw8Y/l8XY9+KbjVEjQalr/W
bgoTeQTOD5LK7Sc60bYWpxpbSsgXqMJnP6a+tKfYBcFCfMt14W2Uvq35Seoy+p+L
wYLcghWg7QbqUFCld1DR77/sQCD1dEYJX09g4AMGewvkq4yrDI1WxD4CTeY29Z7S
52btCNPpla5P5eUomcQ9W1UZrJbzlShQaKcSpVaQHoIW+rP0tdJF1AYvrpxHVPQ4
qKVbd4egakt5uBi3zm1ChQVL1+cfu88ZmthNkE6A/GycQkpMFDwQluCmytfKCd1h
XwLyfuINRInq46GOJhf8M/NFgTNH+/YrOZtRiTkLfAbO+fKnjCxWwb9NQ6bFCUHq
Nq1fccxYiYvqxMaMIkEY3pA0DMn4g4A7ejXXqgKsOAv/UT/HMt8rIVd+v/I+HYN3
r5jR1H2yQVE/NXclvaLzSUOZh65Fhc1z1lLKZla7Y2ZQZqI/kD/7179OXd87Qu7A
c8zRf0gO5ES00X3BgpyH8XPAevF+04SFSWYv44DJESpnV33b0LKqNLvXfVAHgNSN
jpAmAyFJisCOmc2dLQ9gZJXzbwqAskN37HLyAtHuxsjq8W5me9T2d2wHWnEbbdnq
cmdWSpWjkvllis8yOmPVPN+CMhv5klZAp75z/QLfvLQRJTqah666RPqdZyjp1+o7
yaaRxlEjkn4qShqjFiEgrUICNppuzJ3gVQXsN+9Wp0zExHERe3ISozr3uEC15E0T
+UMwxFN5otG2+Qz7Xom5zr+wV2zqnCBRlkVL4Jmt2qaJIap+pBG1rC/mpSRthovl
6f143QYMH2msin1VNxWgVmveEdALzD2e1JurQpmHgzG8sZRfgve5bA9YqItLWJQZ
IWwAhDIhHk0tN2mo2hL5nz8QVHG4wiNTH8eBS3Tj3Bt7PXex29zQX7KWgBM0176x
7Cm20x0whBGVV/cxMj/peXxSL5Dz4KXhdOWwBzGNfh/I5KVLFmyMfFbIsSj0Ivyh
FNMA2PHaX1sypI8RqwDHfYsFC9HueSwayYSykzGyxoJ/FfPlfcQyTmgsFDiExlhV
PkaTwq4d699WwuIMbFWyaEQl7eewQ42doa4ZkDU5X/+PFzF8Tpb3zbxXcB1bBkmQ
Dse0xj7JxlvbGXAsmFf6QXicfmJoTjr6ZXV1XtkF6Nk4L8xLFfnXIcS7Q6ethZ97
oawn/gV3lTXY/Etpw5Cegi8hw1D6pYiL1ZKEca47HSKR0deJGOCjyPd03UoV8ZOf
pJoacWNUEcO569PlLLvZcJAG9eb/nqdUj+VJfLnl41sz1vF7UOgC4o/cGABAtOhc
Inu5/vxcoVa9jsapIgl/WCxmzMeGfCYJpQMSEU+syAepn148rJfNMb/94mVc+Mz3
vTy1CvyGO8RjPZXexB/dPzwbMISRbUIZR8/W37WnN6OnYCaeyRnp6CObZzlgA2Yy
4lHZo8e/6R2yRkqhwten+gJc0jpWP//urBprgpZp/k5xwPnZhxvKG/KWqyq1dpSv
OSmnWGQuoLX0zesEqk77v5+X10WL0vcEpdumxzZItu5tlCX5Y3awH3kWM8RzyiBL
0adhm8oInRutRNUdjmWH96VPthJ0TGJHFgaU4cxpdNrzvOiEfJppg60NLkGMgsUx
1DDLTEJweSVjWqxkwrdse/lvIckSVsbYUuSd32+hwN3BArcignEef8HPVsH7+K3f
6vkgEqHVmsOdN8aGY44od1vjm/AXQkELNKFbYeHatma9vMaqj9dQOnEZo1Q6YBFQ
XmcKyEEQ+QcmtuyEQwWBH33sPLW9jtlIk0J+YbnjXbqQkze7IOo6iz9rXS7+C+P9
FL2m9S3c3ArCjH/hEnBlLA0FR+PsK7d9kvDZSb5Zot3HgXcLUrPuHD3zeMpIQg+O
bD6jHEqomAMDMgQO6ii3bWCKHzuP21LLBj2IG39JfFysgHsxVoxj+tDRKqEwWC3j
O5Eu0wULtE5MwIHosKely6bfOH5xXM4BpIeuB3kgBt4d2Kc1mTqrjD8Coyq/PWHi
Glj8XxgPBqytssHh5HP6kNpV6282wSxtcFO9E3U37lgJbvKyjNnjXrQamBlrPTp9
3jJyAIoWDe333wZfGkKutOvla6fJAxJxYny6sRTkT/5ckEC79HTKV92hnFnGO7Ts
mYCcamgZazr9J5ndkWlWkMmCaVkWpU/jbksa40bG2/47JXDbn2dLnEdH330TfJPi
pFesHYZS+P9CLlDBhRL6GlRt4ZS4nFCyX8QDCeDq7Av3eozSuvYVPcZjZgaEu1XK
a3nFvFnrScb6U679Q4Rcaz1L69PVrje21GFHmlxGtRwbKsYa/JR4butwylJ9zYYP
cNBM5nvRtyT4iV5wBepq/OjFBI+HXQwlVRoTzZfg4yI4qyNLnm8cBJme/1FVkLLu
KiRYMCxeOhIe+pWFefGY3s6G+9fzGYSSPJE4F2B8K+X482UhOV3UzKk6FHMSe7LJ
HKyad44WiG0BYKCL/nv9ClaCMiNn9fWbQ4nJSpBLgnHNyOS2tgtkOOOm7mNMe7yN
Q23df/YhuVBYlTOOBg/8vl8aGOJkrTtETIS7mVAyVapHGEckZntt+4KyW37jvf36
tFWZXEFbfi+d+5tgLYo9+a7XdKg+i2ooXqpnUH9eMjDGdpziHkU9/MSU8ASTQLN2
PLB6AAUC76ZRvfjOFbqPIfrZ4btax5ae6HwRdWryfHXdQdw4oQlVIyUJ7+kyh0eb
V/744HSlptLlr+aSd0ouxBEXP7K2UxmOD94euznrY9NYun2wZicWNfOKS+ZyLBWX
qjhtfj/fbT7td2nX6tVOnGnhz/jVneLizbOVFGyOJu01aLf/d/8U63mYRFpv0D93
1LH5UCfgKuCgltnTzCasxgpGtRNML9C+1prTG2MyLoF52wITYJxhTcDX4CiUa4XZ
BlAN30WXTSNLjc1Wr7qDs/umfLMedfyj/+hCN167/kt2HxcNFTWcU50CMS4nvcqO
7eM6V2X6E803cGS/z0xa1Uj8BRxEMrNcjn5NtHy56fCUrvAXZJqNGS6P19GlgmEi
ZM1yQqAMY5eGs+wdqrVH8iPKFSWFikrc1D3IwlGKCCPct0LjScCLTc7IL669uqnr
74FEJuVwp2qf+AB7Vu7mAsEyCIBDsj8SNdqgvqxr89uG6a+iMxZhcXgPwPUCowpP
aQFcBAHDmaOFiBLqx7kYIGcEJF6l09+EJ+9xtUdjOcJhJv0fe/e3uVfdobVdTB55
TbZKdra0Rw2v4t/XA4cUBV5MJBQuy94mDgZi4yEF43QcQHcH7P0OkeBHYIiUij1G
NG12wza9smV3mbS2KNFcEXHjUT/YlP0NqySG1G/gp9ID586uYCJ/xebhdcC21mP9
Q3rE1LB4kbd9EQOjy2HBYJxeoO15FTUIctX2SX7BBTJBrKtzPCxF/J2xDZ7S008h
GpROhrKjkFv04JbNcg+hR5kHAlkuqH+qq50jkDf8NVULyASxls8Qh2cB1eIRVpCW
OIW4xVpKJMOVKhBOYdLRL2wIb9+ubX4/LWF6MMP1o9Zqf4DgCNfZbBfmzp/I4UVP
sC7zA4xqbxZk004qnx9FWaseNxp6RSs+6xpdyh5HKnbR7adaRW9tUOAFLuHCivx0
HpA71XvYi73wVQuVSuQ7RVm74Laf2Gs3tkChxEnFX6aeOedzL00ac/mEPHgPEEbb
yzCsFxUg/Ksc8UHMhuE+0tzz/b7wGRJ88uO0ToFqZASu32UiEFquv6vdAsYd5qbJ
jkN2s05sJeI5P8QZ0O26CpsGvgSlDnbEQMIXy5L8yfVnLbkZ/TOrfQ1RJrMgytCm
NknSXeNPvTq8+tPogwpDA/9S/PUHG5QWvGJCBuwDm2gc+GSgC8WOUwjuefqgjEO6
sohD6YczxJIphN4Bmdm56uKRR4RedxWsxpZh635csA8KczR14tEGB+gbxSQY47s7
xZzhDEEPxhZvo63vyBmt/fF87xR/YIY8myBXqFYyHooqYrJW6bJ0VnRn0zqaCTUi
kGMbChFbYcx0xDs6Vl8RLAPXZR9vlciEuyZs7OuEeXySKZ89lL3bFN/RPBhuuUtf
zWXlmusKKRqAWXXcfN0EU59nVhaM3GBcNPKRD67Qgykk3NmlLfuzMuBQHfcn8TYt
tZkh9DwzxkIvWJVkswdwF/BNwdnorBAgHruEMKJ1B9Y362bf3i0tVIO1HVVmBbgY
kGWFiYJeP1/9n+qljdDIcrQsQD6iyehHh+qhi3zGMlCeVXJy1KXx5KqOrHzvsS6j
yCdv+9l+CVAkFcjC/pk5mxvtQXVeQgon3znNzEioUt/DPKTWW4KWWnuHaLp1Ye1i
nLZTEqYr3HdiqxW3KQ4nLSPNRQIDJedSa3S6uAbklehj7WAiuRlv8N7rUusuPuF9
gIm419ZwHNukdi3vrqDHAsTqwDMUWbHzeQbqtRgTHgYMYySIeiTjTFayU/3FXfND
wtPe4RBM8PFEO3gdgN8W2eGgXRWHYzdPamu5gxTwG3yPRENRZw2YcvGdGW2Jl9ys
6tR92AB2Ia1ckUC9fKo3UzXZqfoCnDrybAO0X1ciJjw7LEXrfTzz5AfrvCpSLYJz
srYDp0JP8Z1DOLmPvSYtXq+QYrgBSggHnGYw5xNrVCowb0bh0ZPvc7BZTA8xqFJX
cSU/oNZ40dWO/XEf9qz4f1oACzHrsukpy6Wfq/X//keeqVSTNdm6elnT1MNcp8JT
+9syg9EApZePVhp2fyTI6rEM95XFFKVMWbO88H2MRHDHRFpawf2qtmN51Q8V7N/5
WAtP8faH+5ttYoxIHj+CPoZdWuf/VOgosLa/I+IZa/iXZOaruHpWQcxB2is356Yo
ZHauInBoi1LvwysotOlDTakKxT25Tu/8Lf99TQGRcCCbU6ouI5Lx76thjVPoA8Ol
FeXwBD0pWF8tIOrwjKUFaVqByknAzGK2kEgGFE+a4IqcbZuf2xUd3p7gjwoCzRBo
YpgKDnIrKS2wJ7d3mTHxkR3+BGKpKkOl05UVVnGgALCNv1B8DBNCExzAL6/Melj3
tio4Z6PuyfBcstZC/iglRIAzcIto+QdISneRaOGqIrnOYg5IqExppr17waLtJ2eF
EbZ3md7wj+KnYVuNfyCY0pw8ZFBopcQX2jJny/2b2mSyjOvhemO1oYO6JZ0WDE3V
0ivfgeN9zEW7kq+QZfydHKKJJDWb40PTgmyoYR/EbQEPpL9xOMtNdCzBNa5tJYiQ
pvKx2A1bOuSoYOVBtKBR9f/Y+7dNmZPhZpvRHoBFYyDOt4FKqO/7egnl12e6o7/O
uERE9SAA1BI/QiTtXLfUCxrIbGldZDGEN2g7Gh0aHT0m+8ArsWA/EI+Ayx6KcDPO
wqGDqG9KV9+UnvmZkVYj2mHKM+avBpCNSANxuVX1begnP0OhsAukzs5ahKOF6pH9
Qbd6geN9aHRcXIombXUoLadZ9a7ba8fsrnkwSfW4PBL0HHI67ULHH+9cCHfVhSGk
3eX3WLlqzjzHnAoLX9et/5lNz0Iog22IlmSygJcBXt1dp7oW1eh15fnzMVKxbFfk
Tk0sMKvL1aAQtPkJEY93nUe+QY11kPhss1v7Mwg2HIvFLNW6qyezhnbFPBPsh/ap
9xvUnvELvrSj7hNi9t3mdQhi70lFhFa22R7Qmwn+minfYjSpAaVKjw4G7X89PFrV
Jw5ahWnFs7KlLFFMy2fImV6Izpyf4ivFuREdRz1zFNT0qeFCwflZFp9dHPqFAIGD
usJ8AHIVyRJMSNQnBLafQQwSopmzdonVManfX3ZQUoZYvEvhcxT5w8y2Tm1tL2IF
ZVtuS4YJnbjA02JodQ/poCJFpKGuJNBAkxiH61+pOD5Xao26ZyEzET9GSbA3fEw2
i9/VrE6Yv8PVppskcnamChUGgHT6CvGYo/9w/g+idkMjrtI10qqYYZ9pdzjXKKZJ
d4+04LqbcI/FjVu91pe9MXu0Stujs4mU5Yq15A24vK62+FoKQ0ThOs+sBjs7E+6u
K8NAB6TynUV1+Kfk66D2VtfnwuVSDKXNJoBKlZhtjXVOYBfMi+3LPZroJ0PGzggd
ArU/yN77pvY/Tghc4Kxe/kmyxe3SMFWOks3Mxc+5vMMqQc4kywgBXAm4LJpFj5qQ
7hdjFeLeSKLW5EZpftubtxWvxmkAdTO7matPlcxY1rrA86oo4DTvibCAvLc8LRW3
IgVJWk9VeJgzscSS2f1euJrS3de98JH1QcmmgyeVPjg1B87LjfWlpH2M0xHzFtnq
ZWsWNU0lT3iu00hDhmjUbjUeeFHjCaUe6AELHN0rgQTyMMJbibmaM9AkCWWre9Xo
JQask4gC9ceU+KZV/AnJeYwTD9oRIJl5537L0zmZskgYFNfVL+j4Mz2KAhRUUtzo
q3wY8Dy7MSTkV1nvOC6hxRbaTV4sP1sTayP6V4Yy9ascemIxmbNT4RR0KmMAhVP2
bT7FJCNlbVkD19lZudBWDzAE6vI8svdVf3PnrxZNEcgjXwjauyxBIDJ8Ftbx3wCi
zW7GCr8ImFt9DNIlwwD+jbHvZ3KR+ybVuyLNSs0jET8DPRQV8KAf3J7i9NcZnyEb
cTQhZuNDzWAdAqGLgb+54SIQAt4ePZ3YZlQMOocI1xFk3vhDmXhLfPfwBjgMsvas
M8Szk2PQ4LWoYCyuyC1xbbuPLgELbEzWZQH/7MW+HKSJYKJqwm5PzC2BBcwywDSK
b8dt0KkqQ3J8MqHLNY8qU58LDQSDkkHS77klp+gPg1RH82G/VgZL3l/vKRlujxHT
CUA1RKqhWvelPl7thKlPzYW5UF55MMkv3iwxggG3ffK99AVEo25kaW+MJGWhWNZg
k0tkY5RX41thW1BFf/IErC1XOZBlPxlN2dNeQkJv3K/W7WTMCEg8Bq2wFT5VaWly
2GCRDgwP7dbQXkSJ1yxz7FsYc2U2dqx1alGVzB1DwyUWSqa3Ggl+EZmQ1IHaMBXj
NhMitwf7W4Oc7CEla489OU4VZj4/thSEY3yLxXn4rsuDSsEylDbmiTv721AsFsor
YvE9YpDOgYY3oPG9Yq65/Pbq4uEd4moHyIDMwYcsncxBXtMjUt9KgTLxehzQzvCA
ZL27On79jhVMUqboj35Ag7CWai5qwxEPMURIF6/tUVmyL8hQea40SVOAwJ8LwBNN
zYuWH9Hg8eqXUTkKrAdRO5HBaVN7SkNklAHdMCTM8VOFuavzNc2ZJhQVkO+SOQHa
lv4R2AZVS3yRzqVlNN46n5eVBor/PLNZq1YBonthh1qkhA2SNx6Ntzk09ui25USW
KFYxw3oUYClkHQJpuD8D/NnZQe/9zDQgqfFNB/vy3csTiSpM/SwGsPcGud4XwtgY
+UociePdwx9tqHwhtkrwMU+PVFcfOSmR970WkAY3GD3aVn7yL7QXQthyKEm/b2CH
1EykTg/wSwOHp7akmhCG9vpK4hHvPm6lFvEgV7qrY8NZwT4LNYoBDCdbeprH45Ry
Lmg2CQG+gc8c6sboD9AI9e+BWdQ/MUENDjbiL0A60QTk16uJ0e96ibwAezjH2ouH
TG5OJDfWOk64GbKGHWDRZMtQ0UjB0lMn+taDXNVgtYVhQTd7qZoqvY0dgdChBlBa
1OwIMw3MB5FtJ78WK+NvJkja992+LVKOGKXvKge0KYolW4qAO9PeWpAOeb4sdR5J
dYO96kxp6SiaoRoqWFxqdIy1eW51IZMJhDG6k0xp4geDPyk7NZxJ//MJKDM/yCZ8
eQ2yz0EOF1s8zTKtxn09hWLbatxvwVQ911fw7rxlbdWQokph63+79npNSSZJzSpT
WkZv3vetQsd+vAJN7jU7mi3az+7P/je0iIyLV/Ci5hQ1A3USD0h6QalGqSCSWTtb
+UgMmg6A5ZIpqWpPGoHnTzHykebYqxHvwQFWZdEURZbnwouGUFplDv2Vq+1AGtUi
rt4lHWgYpL9ZDQvvASXIqlZDAt/ZX0Wu0kwtBolB2y/oG6x9d8jFItVAqwTibgqV
ps+dMmQfwl/HMCq3/2Wl3868FdSMPv5IJRv60wt80vpNqkD4poC56BaL0PkpIxTj
L45ThXZoRyjSPb0TlPL2Nbw5YvdW7LhGlYHydLOGmsDT9lr5arwbjUcD7kSdaTAV
CjBRoYPgCbm7cxuzJpNduymxQC94n8kom/UkLlWjdaHspuC4A7foOZyiIrkOdXQn
FywtVUqX2l8GB1iLtPbcQ71GaE87C8N+YejGHtiUhDUanMOEeF1JpahXLbD74voa
4QLM699L/1804iPDbak2xN9pi7D2DSHCeMBb+5I6/jy99gaof0z2wZZpEzAaVIQ3
1QrnWFC8m6kcQu6CjcX2zVpttoavHIbSPOqq3CQonTyLfVMFGaHI+65xiVZg4Tq0
KFkpnkkiGrfvtbW9UTw/m3v/V6nq7C56ZZAwEGN2HoFteyx3RC9afamfiuDwMyI0
NDsaz5rfFvaKjTDq/PDNUSiTM5xXjMwxSfjTbYPR0iG8EtU5axpziY5bMLMdMVUQ
WFbrIte/ogasP+7GHfUmePJLJRXiG3Yu3L/vK1ChT2GHLIrNES/zriFgao8eDpZT
BFcT5sqG0M8RsHFbrgVIaxrLPpBiyXLP1Dz+MftZOnqQHaNE81KFf8fZk1+RdNFP
ob4+f/+SXBmnnaZzTIrSYaPcRyg8bHqrAUP+Hz0yxC6fXfvJXgKIm9y73Jdx/VTR
UPbYFBhApKSXe3kJ6nXZwbz/pAjHTrznujSQpN9lTXh1lfNIjONlBKN/SAX4TqBo
GE+paU5XDt2G8GSdoTfTTzirn09IB9zRGcJgCxF5/9gWh1yWnx7d4m6OyhHAN/uP
OQurxScsBflWMIZ2RVmY9ClhM/yRDVUDAItY6W7vCSr2+ujv7XvH8N4+UkmcyiLx
uMrIwyY8IkOWW+Rc9KnIuv0FJC7XkcApwxwduXSYdkSwGVKKUa0yWMTxNZmb8hZS
/BWTQFNqDKDVMpFPBt3apNSl4bsOLdK+2Tnektq/JSQXfeYxGU8C4+zlNLQdo9ap
7KRZrx5/0ieNbyCT129Kk6S/+eIaKstEu6/yyCy5Ct33TpxR870f4jtZPurgDi2T
YOx8L4919DPND9q2ipQIA4H+ZJZ/jZ+nvuUnfk3m9Xzhj+M96US/fVy0OZcnKRnr
8/DEk9NLhq82Hn4jNKAuVO80yaTLkxtHCWGKYrxc2jmSFs12+W7xe2dsfgGWIsE6
i4eKd4g9lunb3VPYmmweaERPwIFoYb0/4m9S26POapAh8xApUWD69vjUvSukk464
J1FIxAZ/w6XhBdHZAsi8j1DLZysGPuwagAWS8IVAE0/gLziDyAOC0vTIOYUOmVlr
OA4Ri86t2lX1HhTWjAFz8oGzseyuDFWNE8jpHi7ZBD3uLC0/OqBwascXoOKglZ5M
OA/T27MvPvZSZlIblrUBW4uHrV+6fSeqS40waqZVni7gWPogsLYKLWtC0pLikvwS
F+RtWViIIF8U8Gc20Lr2hxDqkDjAsnlKPONUj9cB1Ff6bar8tLbwqHgSHwvVjTIq
9mHDxkvdPu7ks38PESyui1Mf00miTtFOOSK8M7v2UNnjvfPtu6krrdxnlIf38WPs
TYfvVEy3mwuIp7ooTWBp/j9jxwPdH+CuKofF1zUecB36g7PJI8jahZ4DC1b9zRYU
r2ANzeH6t2X9ADzfNvjj0OaelaQo1U5Ty8otgESqNpgoKDw8w/OLrmeZ6bZUKtGN
wdzAvYB/nMvcyffu3q7LNL8penGPIbl38fttUHgXBIb+Zq0/t2g+YQn7s+KQMIWD
tYVk6yzvWJPsX2QbrEVRHJqsrshEwc0NvZQSvGAoThAgHOHmCPkJ7ftc0rhrbozH
+lyYXaVJ2x1bBUmfnWcxOgrsjidpNIyhfFOV0P4Mvw5fXwD9OjkmHNggKSum2Ozb
zb/ZibF/Sbe0++4pUk3U6xeKwuCIovxiQ5iFlnjHaZg+s0sjWCM/AEa9SRRqpOqy
VTNnTbTCS3vhOu5DndDO3WaR/0JtNnNGEFNfKGfjem7vJ3dvTUd/f8zHjWL596y4
ht1IBONCSGCqCq5XzupeifTeYUzGPnapHEPyurmGMC3OpUggM75NeoulvM7z/su0
yOUx93LP8FahIpkNmNvxmcI4f5ChfQcjEc9C3lSocwu4QKgS4cqtU1D8V5Nr7BP3
zcW7IuvTfrtIeaRCWgD54tlGJMhc5xMPdErcmnGBNuGV+zQhzY+nM7KcYBF1JTpE
29SaCVnzily5zjEq930r7UkiENEIrjxbNg1IglMpxZ22q1EavAyQGeDHVGaC4rtk
8JyED14TVorOmMWpuOYZJ05joSmuJWfFBGuotTUuw4LLp3uX1hfjm2TAjoIh57LN
FZduDLkMgPm1QU1jJFRk6wGCDk+x5yKUQNhDVnS1dhEC/trcr+6bEYFday96MgXl
MN9fLauVEeVxXrFkRXbLaL1979sg690Lek15g4AOQPN19wRtERvODo7NzpaJzbkj
mSGnbhdZNEkHutWx7xQZB1JkiF9uDBFoQB2JKv5LkpVUtp4frCV2nokvdzFlq9th
BnAf4nUvJrYgbOdstQo6hkt3E/L74qFFjAmX4Z57SswYzmLxtJqxtyHcWg6PQEmw
OFm/sboH7UvL631tr+H4tttDVfKD5WYE9yqgu53KMBlnkI5ewtw6hutKfzDRNzJ2
h7edr2YEAjtEbdXZlrHKRQ7qdQqSrtCuXCv1TynMvJI+lJeYI35SpGwZk93zJM8p
kdESyhm77Rfy+NggLGTje86wkN2J8cllN+q7nzLPMGbr3RZoUFe1MM3LRL4zPw2X
6OMSzU3bPRP2e5WNSEWtDO+I0p1E2X4YoiQmNSPZEmYZzGejtW+RVXMDa7Bc51EO
h3vOVtZVNlM8BKhnLGm4B7DQyZJeELvgqcNa1QckxFVD/69v9aM7ZHgHanEEegOM
gMdG/nF1ic2h+bW9JTmVvMboRpXQzKfru3tgkYi9JIbRW9kOrkTsKlJ190MpU7oV
RyFZ8C7loyy+ys1ROq4FrZ63TKCVkh8XVx9fAQdPl12SMNBtcJa0SQDXPtYjyd54
QcQcDqP4Dme7Q2N2erNmOR4YiZ6dwrnJjmaO33mjF140P4Gw90njozPgPDVixMOu
VjZIsgRxdKwmb1P35IMYx7qOV9G3etSqN6T9MgSUxbfw0NSiqDae4NUYjxNGdDoP
1KFD/CIPTPMTEXaJY03+B6upsjUvrueFWTc+iYmoO0cPoL9nnlqOQrhPWPYkQfh+
ZJL0JadfPXn32av+drzqTKi8MaDHAZ/OROl/vv+jDBFR1igve53a8e9jCVoopABZ
0RB31NHHQ/eIL/4ViD0LFKdgB4PcwAoN2k6YtIiXewut0PMWxrQE9PIvTcnH6xzO
+QA6oMFphRAwKzfPvZJvuUtnE+WH1D+STZk3Giu1/jLPuqp1IWDpezS47COvQUxP
w0vlOKr6pImrBghowjXg65Ifl8MSMUWl8ex69XGhtcsFtQBbjo3GM6ETK+WGinWc
LgLKUcgqSR5hPRCwCEHPMlRPytWZUE6kI5TSs1eOZP7z5Tj1Mtu206jDVN6ZLAos
H0lNDgQDOWlp0r1LAmRrZL6GirlfN6WULzS0xKqenxCqYkGyf43G6avX5kzCsASO
B5Cl6I1jIL+dHUui1i8AxkZZb50WLz3gcqCDIr5T4lgyxenp0RMpaZD6lLY/O3DX
9wAMBeRs1fvR2d5ycl8IIXz1Ks+6jJML1c/YVgpkT9nxDX7Q2SOlqNzH1l+vKfCy
Hlhi0GIwjz54lCj7wgMJCtZ4vW7yIjO7HP9R7nVgd/6GljsdXNLxpj88ee/14IRd
+Z/dJGI4qKqSGx88+QEMIYxR+YWEKGRelsqFteR/Jxk8diCL4CBJvLJxWmrOEf6e
4kalmc+1lZY1zGHO1QlRBOawM4KhG+8sCpEf0snBNCL56BDYMnSrk9Nu7JVTz7hS
Wxyyjor9mdI9CQfLvmxJpYYa0tm3t9uJqxvXRn7MsxDvQHE4mNk3kFTMFr80UsFv
xsASWXGi9vCUoTFFujQj46Gsdwm7WyaaSfelkaHXQoa/2CmO8irZEQwI28AVj33i
HKo+5TN60fCjDtrHhhbrOfFiAPXwHIddZ/SSeX/i1TC3qsL5fyL4DiI5xD7OTJLW
9v8p8a9mo/Ihq0xQ839tKboKYvlOSK3h6UMfTqbPY5ScsiiurCU0KHn6mLYAG2m0
6k3+1yElKAA6M/1h+IVMtJfRZSvIOha1L/fT5xsqLhQA4XvHQ6TqXQa1aPqEh43D
E/Ml09TgYXULWuWLdDcvoQvA6DlKEgtQT7KDK/AygGniXWwPvuGPy5RMXQOLRN6c
zTouIFpIRHKgI3fL3g9OsAEzLr862HV2gRov0lxkmNowRTyw3inq93L3VTFIZDvJ
RqI59Jd955+OVko51qGIxxwsvKuVByv3WdgkaUx/ggEkYbQTyMtp0Igli+GNgMlj
Bc986dmq6hPvwWofnEXQ5WjUlupwuzhPGR3OlO70mpIlsDaUMuD8uwfhy/SH6RL5
VpYX5LPyo1n+0vcUev9Njw6fHnLu9KlRziogm9B+QVELYPyJfSmV0U4Wjnp7wjNc
klhWFW4t2HLqokM257gjQ9jcSOh/eeT2FKU3UKIh4DbKxMKi/3EzdeWWM93CkzpU
5yjx35J6I1J9r5OM9AdRbaP3tLmkQDGDqAjsUf7OSq+F4GsLcFJmTvs+DPAgaBfR
2lzAJkGjaeCZbjLsj5WrSujesDhXQLUzYaWlheaKDN6ZfsJvB8HDJHBUEumJmPhc
NIeuItASmYh4jmOEVjdQAn4a7rdUMKoi+UdNb1HUrCwrbeHpQOTm8+oWpJmyIqzC
jTDYMBLaAeO7d7HodACCJgv/YoEbYHg8uQ59W6lMfUccqxde7sGLRs5chZF4c1YK
770zYO5CHXI+U5aTxam8HhPzFY5TnPDPzv7oNEszlbvHRVCVcNHoZJdiI5xURApm
s1glNRqa4pD0bd399YY9XKEUP/RXoYikxX/FdjZ1/s6l6vib/kxDfBgoblMmHEuX
HDOPFoNrh34qV73iI49DRxn/f8mwl5r/xNYPqpBmnyNOndpQEM9Wb39zviYEZNJJ
Y55CyBEbzWcnnRsUXFIt7yXJGJ819sHkHUUBhbCTIT1a/IUOvhoQGk8DO2zgKQYN
AUSPFup9AI/711daptS8rgy0hr3TJzXjsOy/9xqr6tHAzCcD0MQbp/WxniUMUkE1
1MLCroCjYuchswekBJiffDEppkTgb/FXz7lcOiukGjvu8Vz2X0YlC2IyqRqWbPT+
lPyVNaoFatwym3l1QarOXgadggrxoIbZ0Pmpe2qj8GRW42PwvC6+hql4WehS7eS/
RXYOqFMBbu7sug0Tr6CnTgs3XS3IOILFQiSfpj2Y1DBa35h3su5FRot/OXQ0US/O
gqh+zQ7s0GAGW37ojd3xzCTjcLsZCJF7/z8yuZXtvPDLTB2grQiI2lxKzI2360Nr
IlFXZCgsgPBdWQwamTdGtQuSq3jYTjTSeZjorgVVw5nVqUCPhrCD+GN9QZ9oL2he
WRBbbmTWBkauZvu76n41vL6g4QQUvucVDJVZno+Uqq3wUhqfFi+55M5t1ZLm5brG
hTQfXCWr+AZiFa3vGGCYQjXtYaPzvIrORYdHqs7HzgQWBNWNs0cNSdfUcXqDfoXO
YxbSZSUVqFANvfz7RxPJmGGfBQZWzvMgXgJgW+/WnGAk8VrWmwRszZCV0Y7rLBKh
gj/X/6lMXR9zWbqQnz/zg8Ai8Imj+CdTwMYZOr3yb854cIwttFot2NFdNwfY4Tur
FngGs3eEhIOcRVSTKZ9iSrtsCIlAGB45JL/tW5poyy6BOE3+/UU7BJakUTZako83
V6B2psBqu972zesMhDsyuVuGHolRb8fz8KKIK0tTajLW6RO8ell1BvJpazFP5XCq
HFh7odanqfrm7SwF13kThtqx2S8gOSU84pLX7ldsot8/ugedVrBfvu6SY5JysuSJ
5pnT4g3W2+WPCGlGPQGEl96ZgiY/jwqX8t2NH1aYE1tGMv/ZwdAdVkfyBI4uoenZ
2ZDZJ1GvmqVWj0z3znEt0h5iQrH+6cooJDOcByCR8vkArffyafsCy76ZHn3eGGP7
hT3hTObD/fNeyzMyw0vwhGP3CtJb5JKhRGXMCMaTryZrsuVn8uZqyrxwFLAVNJoz
SAN8VLW6Ftg9WZ7s51pyQVGcm+pft1Gk7of9ESxQdMMWC+D3wXJUkcBY5WcmpuCm
6haSnF73ud89RXido3Gmb3YiAyrITu5Hd0rULVav3PqgK2EdoSx+RYQIYnkWetb6
37KrUwxgFiE1+BEVAGLu6DRf5c86I9nb11+WR4QQZMeN7MqsTLzp3WwqPfp+sZaV
mq0hVVApgifI885fyl5EdYY+0DhkTFxiKgIb2vtTeacEgX3UlNMJpTRw65JMk2YA
zBtK482POfzGQDrIEB9WpyS9U4NtC7Z5U8iMWM5802bYRw8VEu9uEELAlsQBlsUC
65MMZD6JSMyW6K92gX3PU/2jjLvnFuo66uMBrD942jq3jaGQ65EIKjUJexTsrrDm
sItTykdV5S9emRjwLpCpMCA883AP46soHlHSI/5njyywva2xGqeixTR25O+jL0FV
z7g4Gpz9xfPEdjklXKWez7Z2h+S2Ku3cQisDozTr5iOlB5Emc1xtmjgUectehq5K
mexRUjELHISrUpzQU1lAReJ6j0d1wcegx9suLS/yy5xitoG+vBAtQzVr+CwwOY3X
Nl6zz0NxNSRJoXrwp5+RP+/G1bjS18ocDkFKy41okhXyggAbJinqh7ZuJU9ymJFj
jzJpf7XNV7U6Z67p+CaJDaPHOXKHhxe4HktuTmlvhOdKiUNWAzd7yXG67rA0j3YY
jS4DrGSsAlQcVJx4OLzrhR8vw74XxCbV5Oleu1zvEMvYenkRWexQQMG/udU3r0JL
qGY/5PHZdr8vO/h3WJEOzzO3MJ42t2O7YxaXoXu4+z5nO+nKPJoG6+U/PtwCqYHU
mzTdQViiWR2Yu3w/r//MmQB+H0i6t3arp4/MaFhBZ+GvqShRYWUOND/TuUBSKoHu
g36V04StCX64yaB+wLEx3zZiMjQqvCYLmlQNQtqDUhpujRrwZzDsygbBMNQ95huM
VZ/08FQ/8KKsvfQ0upL1FvR9/srm5afbav3S19OMI8DrOlx1jvBtihPv3fPHFRNY
qqs8DNEMObKS+w8u8mVaGoCMgtnafhosV3o7DZu1vtA/pUYpQ0fDmnHGNFawLrfy
JC9dIYhhl9Cdm3sv52Pf9XrDAg8h+UbTvYT8FfPMvS9I/1jmgsvqnGBS6XzPFNDI
hfr3lkldB9o0uVMojKTJKkq/qsjNLOhRyIolg6iduAgGw8oriA1bm3tf6Lb9yNQ+
tCTUlacmboBo88fKo4PrrYPvCgd7j0h3VdXgxGRQ6YKbPaSwTyEkHMfIyLRn6LeA
XoDtTNqUq6cc0A1IJx9glkjlV5aBKtSWZuYJu4ffn66saWZtOWg4nToqzOMMIHTl
4ScK+9wXXY4xrflOnqxJCkPYICSs+VMpXcUU/Qr+pZFEUxIpx/7XoKvN9Ukzg1+l
qf9j8MZ+wbSGdVftPi+VkIAgBSj9TVfj9S2UKUEuU53f4bdREa963H4MrNNQy9Qi
d0Nd1K/o8b4W/nHyBFOLglLKxzFvY9RVXWAq/9PZGRTyU/bM8id4DX7GdFy9FADk
2baSsBl1avXo/SSzZ5Hj63tcyvAlom+6KyMYCE0BMeZzi2YTzUk1CYP/QAgnMBVD
7R9YIAqNzFUDGFg7JmHqep7EVKMPCR54fEiSuvXLcZJk6HuZWJSL4JzheqMqdSU8
uBF/UqZKju9G0N4ab02AsWfUZ2SPaPBd0Y2Tv3w6tjv5KChFOn7f4WJgmQTtMusR
gEZwI3AJlc7kq06YfGMiAZfOoalT0bokIGtrqtMgtHOZhic8/l9LQhxcC7ykc0bU
PTouMONgZboByoPBO8sx3wsPiG4/5QhGdGZ2hjuShQQy+vxEGM0aSm/jJTNVybuT
An5vKdvet92bu/Q0pMmkI+5GkRb1KosvPtNJQGi0aWvQFz1rUyUDfQ2jjMtNcgLk
oWdJq/GIeVSKr++EBEIw/bn9AqM+64cYBTpmOeiNfxyhTYuciSj0naBTqMHkqGBf
wSROs0Z1hwyD7HEcXXY3HnXa2VHGmts+2sNMAOAxkGOq23wnZppqcITt/ef/jdlC
QayKv46HyuTd5VwEDOZXkwK7p4f2tTFWzJyqPU3Mk1bULdjo4pdyfFlXg/oy3FbY
gkcKWGG/zq2Hl5DXGFNygBaChbPnGML9K8eSqefkHdDpH9/KvOVyNJP4BfUwlBXT
dVWb1pal9Pk+0v6qNtdxYFvD73ovE9pYkr3vngyHeZ67spHCIa+N6j/Xez+SaZA8
kIXejyx3MuP2tsw+GsP7vD3XoZydeoxW1ko+np2bjZU/TLqnrrcHFcpIPQKx0k36
8/87EZVTleZ39CoyUCYfrfHrQB1+riDftxtrvX2cx8h4Ceu5XHte2sQ3ykC9B1Vq
W2B1St+vT5Ftu+JavP9O+abhVowG2rLANte4M6BzMBdV5nPJj4RNiCzVI4KIooXg
KaTGmSfkDL4KinFZM35PNRbVrkPOhoBpWJdOuXSyGlKX2VAN0bVUrHIch3oiTIzt
4syPo1TjhFdKzeCC9+p6XNqf8H2ZMr9RMzHX04ywQWoEhhq/J4/bRhuhVZtUk1dj
x5rAphhByO2GKdEdDT7MCNPt+1LWAXNFUBvysXSyNHDP44nH/O8qF94c0g3lJh/L
rc6C4aBOwFObPi1PaHQA5ZiW5OhWloCC0ezX7z6CuMI45nCzrDkxO+pZQ+hulB/l
Uy0JqraV7z2mvr/FuSsoskh2EGBP5nNwMN18yYAdaKPk51cQnazekanp5e411kIM
mOaI4OPBAHODZm2pTgzwtq0Ii7IO85vFueKaHXeLyxTS/xUq/ckEx5UYs80q3PWn
P/DTCLu2wDUd2oTul2yKW4zvtcF1+BOEySCukduVHnHpSnKhV+Ib9axBu5/H63FO
RXozyE85oTZUT2Ru+lnWUTgjzG5oQrrTNpYIt6FddFPCLb6hsnXE9gwGsb4ZK2fF
+9EvxU+mw+Wp+zQUT2hLeIwHqDdKnRJETNOHlwdBozGZInsVVO0oXXzM90aLtTtp
DZtGMaVAXihpwZ/vDPjgQlqvMWDc/S1ObEvVEUUL7lX+ezr/hIZRF5102NKXl8Kf
pyK+rvgoHqkLPvO/3SKJ9mtWnEYxBnRB4gqhJXwxwDbw6pzhcRIoLjRTq/Mq3TLe
tStWNm1DAdJNZURf8EZOZ+vLx1MW8UjhUVMqJsVeHGzDHDrZUOnHWxvHguTUbh9m
G2lQt6DOuZdI6mKRHSpcM+GGGckavNOPV58x/bDHX4OopOTgE22oj14PtCds+VFy
jZ+x+XFBHCZkt0aXSQssuoSiWu4qTqcPDyHpNObIl0Hh1kimF00XLK0LNpmx0cuF
/fwxKYNCZiaoKmJKU9fZKVl5kLcZS0quxUzmcjprx9gfR1FClPvUbrXJo0p0QGyj
LFWDsfKRY0oiG92sE47Hwm4sP5fxWGgQkmvqyyD/9ZxkByo0DZUADV//f6lAM7kW
1imenSoCEOgWFLDZNTuDOLb/vyt9bJMPVDhLJuuyTC3Ffu3nAVYtkShgmWqwAgiM
pmrImfPMGLtbLDnX4xIRWdI/GGCpCMnC7N1q2XzX8unrzTIjUtHXAvJdhoatyIEH
HFmpFzWG3VwGvBgmPPb28gBBP6v6tz0p+V11fwn3v8qru5QLypDb2M8PkG0xWLxa
1J7p7tVOwflI7CpwYATukIuiFtUugPV0KgyRkIwsW8aKo58czvQ60KXh1ppX3ApQ
HyGOMAcftVmrcbw8AmsOjN9LDoRIStswAhSNbog6SeU9SZ9R6uX1nHTHI4zDIrL0
ysUUj7efKp8245ddhyeJhuTS6fWI87go1TDUTpLWBw9Ycrf8NCZzK6p4Pvh9rMgB
Fj+HofiRuijuB3l7FWdVBmyzJNvpNqonI0ceuAmOH923vhlXDAVlTle27WIgCHUr
9T3zFZx7TLh3y5rX0P4yrsbAEjEc3yT9i8PqQ4aW+yO8yrMiqfkxONAaeyZwZDK1
5hErR5OA8Cy+k4kgTCbU/jYOTv69dZ1YHXlFABYbDwINdydIGm75yvqFfUzWC+Nx
L1I3x8gCP2GaBqQny8YiDEzKZKKJ74AwnBdt0kXdSAjgtta5qpXl2IeV/0DW5qf9
z+rK6yxmPoBHgXu0+YpPTixGnVT+wgSPjrLjd0ATxQULibzbrJw+/bJctdTQXkLF
Vf/cl4gBxu3ZqZR39xyvW87/eSQFybFdoHvkF7dg3aiguMOLU7eNbuFE2vU3nifZ
wY8DVBisWx3frOF+HO0GhW29nNBrqwZl5DoU4MX6eR2Ax7qf1n4EhlefI9PSvtvV
roEMaBsk+YOhlUbzunio37XCOL/ACry9embYNj0R4Ad8Pz7iPIsTg8qOKsDFXflV
dn81uH1XmzbK5OijkcDFabpwRUbVxWpfW90Yx/JORN1d8yw76yYc9QH1z6KTiN3L
sKXh0ZnFLCJPgGNTN2pFXnSndlOZbeUY6SjlYMAK4/nv52SWKRALmZ0i0hWALFQB
gS5l5ziAn7/87SirJxNST7Z0tbgbVvIJ4hSxedn5EU+zqNC4oM8dMSfQxEiqG2zF
pltCg2abnd3kXCOh51dWSvIXl8/vEi4udfxcbL3GixEKl7zcAdeYfnMdXuzRVjEO
l67vKdxohvu7ldWT61Qs6ClW78R3eyeupZ2QpZc3XJ5XCd8liYfhv59Rni6ghZLk
xD8Rp1z9Y3fWoQF+a27W5L5sZzAoqlwIl+J7RUPfzpr/qJY+NnOLK6qKbViTZbD7
BsdCmElghvhG75bv3C4hGi7tI58NgKYvYOalomkh3n7uPyMGwFRe7MKt+g1X+mDg
A8mm7BSIIJdq5hxAEcuk2DwnyTxNdhwA8tizr26Qzk0OVoR4lYEo7G7X+pyZKLx0
9Mnb6gYrHrK49jqYERSqCL2gPlEdlYRspHwUSpawgG75C3HSYAxnqSvIq7IpqiRD
lRE1TIjiuOwkwZQS9n9DV5IbpxZbkkcUSOY1oJLkxOFsfWvKSyVjxMikPjE+iNQu
XDBil24VjUQ+/BJrEtO1mtSBR6o+G13AqRvbUBzgSx/VtHip4bckzqkyqvAWim5y
LZjU4hCb6UVhriLoDLcFJQPcUJXc2rRhQUtTIWtIhIGE1vMxhcsB8d6TMpqAMOK6
AfiymFjfXxN/02RCKYPBV8loP7sRFR7OJVuTwKrckLDZOKn0t0t6AvnB3sueSfdg
pUeq4b+ECKOc8KJ3i5M8/XeW44BUEJuyrxLht2g9zfUU808VLOZ/JihpWADzohBX
bSSKGUPXahOmPmb8+3sQu4fCCtF1gwRfbC/xLgGOUe5Pubfl/8uUvrV3xdz0/D34
X27fb4FQlRa0y7R9FVIA2931x/Sm3YHvXb0WA0SJMss6GOA+cERBQFXyzuxMdECB
rADZLhZEgqLuCBhDQjRfvpEVsxDGQ5NKOMJIMy8iGq5MkquKwJsBRadp+jqqTVHK
NGZZDZlFzOrdDr2OypcWi0+xUrBfKrcvyHSs3TbemT654hONJvvtdu/vFCJWEXHf
S9WTHuKXH5VQKC31S1E4Qp6Z8jxeut/QXepKMtReZ+E2vXS5vYFyU8GBTvAOo+Rh
XtvKep/hjGEXaryOgdAEwCTPIiWYlIrxgpiW3/eWDHRTnR/7WzJef21QoGu2L0gt
s8c/yR4HTWyYx4mIeVLg7UnhaBO6dclZzVrkCrx/ymjegaWaeojcZsYEC93TchzI
MnptRCrsn56mPZe5+f6mMeK0RcwX4pJgLgF4S6JeyGEZKB9qgtWJKKYT9rEVf85+
WOlNoS28kZtqwinPJ1ZvXIrceaquFfb+NTZ1weAvcPHdxLoaRKaohlHZLOFepx04
8zU8bjH7Eea1pQels9DavDF47Ogkc2Xh3aWgjaydTJoiD7qo8E6RlLfJMVZmtDG1
DaCuUW82tja2Vh5bRceG6Fwz/BpnaBrHj6P4WjHkIwDQ69L29ma/jMfHFWoGD1B5
ua7ESPalAEU90TAtzJVQOQRJO4iLeits29tXZNr/OFUF7UGDL00S0kByoEh4FyIo
d7b8Nwr26Sn0HW7cpgwdEs7IRWR/LaFNCdXWSaB+K0nV/Qu2A2jmkxBL3MptFT6x
eDJBP9OpD3NmwxSTCM7LcXdkeeHlmK+uARFbhVmi9NdJYEtNPodepgZ9tXilPQk8
y2VclMvtRIsly93t9s7nndieTnx96gnSe9Frxn/q0+aAOC8pIi4t+ynncgCZuHGj
bZtu82oEodCvXR79qdvDDMkW2g7jUW+CRdMJmSUyoiB3x8/tBkG58vBtq554TVi/
LMohuo0Eyy7NzuGItlmBJQb2q1F8lHYja6kZ/lWvetRiKTeDiqyYsWHI1BWUB2uU
qLTU7nlJOmpmw9zgG0ho1Iffp0UzUAqaz/HGCXSwmICKXNMCu3It+94/tGSheTgL
aj9b9+UMHcUYGiAYVnEU/Jk4EQY76zLW3IZuwp+NsMEebWX+1ni+TeubKkTY54Yh
Jq0uV+QBt12mRXplnNAghlbLDqpWCyR0BAzh75j32ERFJ5zWGqesi56XLVD/oamn
RFqyIY13r5IH4Q2IZnUWAQUqTfDv9lC57VDUQkejB7K9KwMxSd+N3/16s76dfEon
XBUe7qxWT6kafRHT10I/hmqplYEYLTdlUzM1FYh7KYARH18nih0SrEADR8NpiQiM
zEkvnWok7RqlY2/pDElT/dLTQEhmU3l27kCU2aH656fXmW51yM6Am00bQjyIcdEj
nlvonfaYBsDUGR1HFwpzOY/GtixwM9gYRKpmJIUPL2YSM2Y7SHhtBdXxpDSiubHy
zkSz+9calUQL02veCQjYdc1F+f+CCrMKSrT0UjrG+SRs+yatsJpNWwb7QJgWLmPx
NVPfWUnQ7ljHiUtWeZHcqkZJyWzDP8jHlTb1hZNKJI1aNe/hS41JNvDSy1ce+ufZ
JjNQx7Bb3ROIydcaiWil/5b+evS8Jt5Qqd+Y35eLw38LSaXaJFTS9HbG3X30b99w
Mg2fp+FWRp4J8l81+kkKarktpY0gZMRJHUTdrgdwRq4AYKAdMZ7YRizLYAV+2Kgs
xCoWyEO1cjdFY3Zsn9WI6rSCTE/VX9vgnPNuZTs9HBqCG/6snp7mW+wxZAx3nmSk
mr8FLFakxHYzoMBsEagpf6JiHiltsFAmS5b9DckRB7IdP5vEazfcqDqMjM0xUHoM
UsjPcdvov2cZmZCPBJeqEicKaFmXUC+ge7HnGRV1hWfxzDOW06tKRPstVTy4o8wE
wpwJOU3jZ1pbt5ToDJIbtQb+g9rhP48ahxVoyk/TwAZNaC03z+XmqKDFLwUiASg7
8hc3Z2+hlh6u4l2HAWeiGObmbe/KS/JXCmwxb8y0I9sSNhW8v2394HzM2zuBu0xY
NsK5WDAkpLZ59c1L0ovobxd67wf7qvABrCkGT43f9sSF6jJ7bXwcWC1z/K7S+dSB
aYTvnmln4VxBx5AaFRA1G3T2pdlTk4zho7xVubEwU3C2nD4Lnqu7Ph54SdQRo9J4
a5pQ/SejZoFlkHOZquO5O0dskmZaxn+5RZpY8JVJNUER5cUUyIb5iLB+Vrwd6xnn
8w9oDFjlNQrKY7nDE3ysnzja07tTZmi9lZZgFeqn+OV2/TvnbAC5YWpC/GDDUtTj
sQutiI4vEPNrfSWKxxRaQYbSj1AqXwrne+SL5zYRwhiwUykFWrfH6Rh8pOd4e2nx
UYU1WsBU5MxNuNzAu5A4Gy/Xm36DrSKrEChnE9SEaPsBZQvJYgS794Vl0ryJofL/
SYdUzmuH95NOTq7yDee6ToxLeHzoDxQY56zq9JKlMLWEgnWfVWYRpIKtv4OSSZP5
6XUE92fR2EtlIQ6CrzJ3KRnx1zqwV0/lsUwP/p+XymrMUmXgmLowcatOyFqrRjBj
W+iur4PZ8dy9L0E2w1KEJFWnkT1WGxIIwXJFKrxxydf4jKlnSHcOpaRHwq3Sfb2j
684j5pbbGc9GKIhw1gIs1p5abo2hNVKtNcxovTcvTwBcDXqYxuRZZt88DYZVNnG8
hmygkWW/Sbdr1/vrXrEZoyl1hz1M5HJ5pBIARJCVMrBNP0tBE48AGz4/l8ImX9et
+z3jcwVsiU2qrsEB1d0jHzJKMaOIgfvyj5vVRwRcuSDEU7O0+CopkjAYXEjxRTdW
lSpPd377f12KDVdVwdgPfrKxoQrtYOIHlkcFEfpRenb8O4GS53VywhH1r141Qt8+
lc40reNKtJBCTa8ZUotLKGboqQpXpb4+TCk+8JFwRN+Vq8xm9q9u/Q4eLhR9IVz2
zR2Oyq6jd+HMpSJM18Tfw7C/Wver84hYWjMZV+zZSve+aX9LQg1oqgwRGZyp+YaA
7goQuZVUuqlXOWHCLAM2MpyXG3mFo9Zh333z0d1uTX+ABGo76DB/TrQQsfrcVDGh
ohPmpjPy708balAing/Fl2NX7jx9YHF8zmIK1IagOJO+1y3FVUao8/9ykyo4G/Au
ESUl33Hh0u0V9+lxdCktkfeLcCagTVjso67hznIq7HTrSOBkbCLhZD8coS7DXVHG
eGyEJ6q+2t/HCbcczdOXoZZW7AJ8G+Qdmc6PUJLFMY70oDti0IvqwnlpS05mvkwm
wusFXUPN82WvtlzsUse9S6iEJQzE5SSoB38mKZdkzyQe0eEIEFrEw1mNTTjMLt3c
LfNzSBsPtn9rDFjqB0zrGmY9z7Opif1NIzyV1XPR5lz7dinrxchMgtnKrShLhByH
DkV5pumi9foM03SXccDha9bX4HaYXRwC0vjBdfjLB6Pf8n9YTMrk+Lvo5wRd6FeI
xaSseLqc65FAXKvVg2FDlQtvQCnSS/S8msaOHNyeH4AnNPNeosnvJrxoDqtHS3p+
HZ+Az4Y8rvc8n4puZXgCJVIhiEPWVm9HpiBndzMA9N0E3p0vGPMZNh6sQQ5Ii9Mw
U3BQ+/gSo2IO0vxdZ4fJfJE7BCWRuCedTTCodiXUH1lNn/xNaoqBMWo3Nn62+RwL
IRGYJXVEelmcTUlkQP3uJJPXobN1DLVWcIgouHBJepSj2S7G/uFH4jqi9S7pYVtm
eVKRdCel7O7pkZi41J5vcoIQ5/EsvbPfrYrbyTt4N6au+b2xmwVxIa0bkLqGQiyG
Zv28moR+eKnfSl101ZY+Up8IAfQ4o9f1MmiBG8Z5TrWt9gi4yVzkPkZYC9kVhIeq
4OzLXaSUE4DNB7yyKeGdpXLWF8etspU3xyD54WWs5mOB8bozH6AgUiKZlS3TBIJw
YgHQh6Ya7bUOVNDGJ0YpROsuGGV9LH9mv7NqJ0Hwnw7pLjZlBn+3SSMVr+10frRZ
W4KnOY/1TykPh7wHMdqq/cSVBZRcwRE4d1oha/uRnkgc3wkX3HxDKCLV1CFt24A7
KW4Rdl/dhfdRoO5gd4iCCO/CQq4I3hRU7asCoYQsQ8jPZzLJaX30MMVUbp7JiIfi
PF/LQKilrmjbsmcWCT4TYdzzqV5040sXnDbH9gLoDGhegUdwmDlnDWxTMfn/ySOW
qAEdbAgtP0s9IsKaUCL5hjDcH+TaJZqPvE6rM/pB0XWuZuwkUthYCxLTucwqLFHP
Eu5ih5xOIMfe6MzOfZl96p45nrtlHQda571w9xpjGz6e2P3JOIlwp68K+J0scV8J
jZNNCXp9SC+ap5qsfWN+yGljhlfwL8Hm7dqwuh55GNsiu5nvtIjPitH94U+3+Wzj
AKO27P3fLS+VnIMTV/orQsuUaaq20EGR3wBuYRqSRtRGPBvb9gN/MoHeHUKkBTb3
SFVP8CmdUILQlqEE6zCv/qFvZwTCBgU8iAXCfqVCn4D2KBkZ7hZNmFzPCGcjdNRU
rT0xUeD3ko1ViJsh0b6TkPc2D9+FnLucdfXnqv1ZiuN3cfJJVmwqpw5BBrbFRdIN
9ZYUVLW6NAeeEQOCIwtAgx1bswLCvRoW734uwJ0CJCtCvwiS87erBmnoA40zb9CI
pwS/X48T8JS0GN5W5gu+Mum2xVxU0aC1xsBvRzvW2Lfg0MWTgJKrC7BofhBojXO1
vPE5QMki3ceZ3tGWjDxBhgS3SACgt1zvJJYAn0AIJFaG/UG1/+VLp6hkjPPvbkl2
oRTWHYYRgrJnJ1f9IjYh6FmMzbJbkC5NmFJW6XM8KdsURFw6slBlYlvTz6wGphjb
vVFa3OEaorxKyicJVzkNM5tGBlxqAlq3bDIsRB6TlHU/USxCcSOHj5kXbnuM0dp6
J26onmoREA3ZZkX8yqeVXPGjzAk3AvBTGEqBVkwFKaCwC/4E5AEO+JOLCxQRk+kU
2DQ6vfgI1iHIGO3NPerAKJ+G5gVjnH0n24MFZfLIRGWjhDmRm+s79jA15KXXre2a
pwYJEZxIT09SVJ+auUbkFUnXqelrcY0qdLyrxcgu7ypmCIwso2sx9bTxsSI80MSa
d4QcZuRrvvyZMUjEqQGWKIqMQg1OumZ6aaHsFt9Ct6OIAk+co3D2hcfJM5X1Eeg2
pGMrB+suyGBLyhwo7rIpSHHUZhYgV8i89YNvLxeZDrwWehn7QcNt0HA/BS0/BezS
tadeGZImaqj2N9odiz4WjediDxMdzvxhIpRLekG0+WTzo1/2t1KyW+CaXu/0IPLF
wvrgKdbKK9gX6B30yvrkk1S/OQ8C4/9MqX+2eAOHAbWgRpZOYdv+ABWWWfY6BZOu
1XFfDzFOfacqJJTmX5LpgV1Y6T42KBlpJAQrF27kQyJz3GTRj2hxCZIUOlVpWLlE
V1PINIzuP3LVbiP9F5M2WzY/qVQ24MkPMgxc3lYbvYN3LMnzP2lVVQbnNLQZa8Wf
LnR46/Ne5yVWt1fFQJAcptuGxLTHyTWjO2wGcqsi9uOQJ8ER8wTChfnh60SqF0oN
rbDC2XCk4vAME3J/x1XUUNKH9Kvn7VW1DJFRMvZpQc10uyK5aprbFOCtDV19ohFD
MjNJNc9ogtSeq4dqKHiKvnE+UmEdANfcxf7gGt8GrTXHMzHvfvNDgNEnqfCZXsfk
/sghST4Kvpae0cAcVk9is1c+T9wZpKUTEUl3Be49/ety7KrIRAhiffamiMbyexPz
vxVRKQxN+/8ZVxhyUXd9wd4IWdwmwSDDbzX79KBBGlR6MFXQlPtSDt8WGATCXjrj
1rFoarcGqY5mCLrqn16ULgD5NNB0SGAyYwzUNgekRvK3TIDTBtwg0TWwXlsaDA5O
dRIeS2u4sKDhqCOi+PkRRKW6ihIn4yqe1OYIaqCWp75A2ihpreScJoDVGy5C36wB
0f99IfJ5b9odnKXb7v5WhoUwuInp+c652BJpIBxBVOgTrldszyqQytG5AzelAPsC
KcEICehgGD1EJBCJUE03pM9q4KYWJKo8D0a4ITzL+4Xaj6su9X7s8ga9+wvCy94w
jMy8r+ndAbkwd/f40l8uWUthrzjjvSCKyT/JrvgfuozdcfnPCQe1pzXjJfr8XVOR
hIxs7L8NTFso704aVbtF/dn7y/ps0sM8W6bF1xLOByolyVJooFm9m6HiBE/wj3w/
Yx4aXJHbNP3K1A8szLzQifjAYrH+i/Tztfxu1Ps+TN+aMwQrXqBE62g/U2xiq0Fg
5msXAXYzmqA6lNYUr83xdB2Rg1HtB1iXxZAnIBgn27J8KnP9haeUXxadoOBIc2m1
IcOXSujPvJYsFR0EtZ38cxwZGIWJlip0XMpT8AlWEM8OSV9wNLX9k4R76RtTVtYo
gizdwiwnsfL2+Hw+wedLh149vTdQSMQ71gUySMDRqknPXjlY7iXhIFPk9bmuwIeh
ExFufCqcRNU0lM2ke7FlifndABCLD50v7yeC59XXV15SHd2/E3IGe7J/ZyviarGt
uIqHWmklGUHEAtvYXPDEDogSKPwtsvIX9dndvhQ1eGWSEjcJ6kEU2fsbFz2+Cz85
je6L9Q1AesoyTk3HxPansmE4epAxLFXLUYJD233EqJhc6PvlxwW7Yh+9HVTS6+Ic
ZF/aU6FuQ0QnOy9dXR12HdRSrah4q/juAXtKfrs7FsqPnF7UfNjWAZwB7Eq1LKhd
H0rAEu7rUkaZXVmfm/90Fc9jWxjeKw8Coo9wpLnFxAjQwjTi75ZQKuDZqy8GgJNR
sz5BubsdPFZnYMHiWIfFVg+dwqAKmoUke9ZQm+EuSYRqvclt4ytGYPTjvo4xHjcI
rjB3d/RyYH1YgZHngA+SOfCtismZ1X3r3YVrOv5gDQyTzXPwhzBRz3nm0678Dhsl
QhoETwr4esKv0kQOOUXGMF9Y18OSOBa/lxlIP09SxMyyu1+5WeJahaLt8IkB4iki
SlXNHx0Umsdy2Edsjbi4WOYQPhEUD/yaPLQALR4q/a2r4aWpL1s32G+UahKB2DMd
zxGfcHrZXKnr00ALyvN7OumkYakQOn0WfAP0gCwa23oLrCGbDE93+aCZlhzkfocY
3He0ugUWywg8gwBA26nM7flcsNUSv6YuKB+yGVpiV+dxKt4ye0SjJSXXjouvxn9H
K8nLSqKcqiGFTPduTi9UUhMMZihUEXaQXoCS6K6qCe9Y/51EOBQAEVihsfblYEbj
YyjLs8ho2uyt6UDUf++WnxArcJF5y8XfpttYuP8iK4vGTA0RiFoGL/FwuBbC66Iv
inqgI2cwS0mzNCq619Iz22s4UMF4ZXK1R3U10lf+CZ16DZWrer0ejtg15XsWXChW
8FsM80xPT2GOABOkXxA3pT1Ku2ncu1g0cmSbVwHPJN1rvG6pGOHm5q//rQoRQzyv
CS5ZQjxumvgA4//0x/fGmPm4jZuXwLI1na5JTJC257MDY4dqzqSsmljJtQbBKJCu
OqdRFlPqKt262LaBsGtyohykj/CzgcMy+63WRpNo5hAp2PyJQYQdYiMAA4yfLm7N
yJbu5OvQBAP6T8q7XYOME0RFHG1byVhmPVgldXGtoyp7B6g0hKPMqkJc/1CFYW/t
flEIR/KrmgplyjtV7Egvw398fkpS8N06P5raVZbFRlIRAVb3dwBom/Rm3POE6P8u
KT1TfnZ3T6IJ4EIwrwOxh5h+Z8G4sgtxuTW1nfjxOAHaAQVO30h0TQWMzuOnLN0c
GJMZjenU+VO3+BSBaqkeZwHOCDVuVgJuGzQokTL1RX/QjVAubjQZ33C54cYp9xkD
LEOY1X3OXJu8uTYcSnOAvO5JQwzzWWntk9G6c7of0Ock/cQQFqTGMG7c6Bk+ROrC
sT3QOLz5v+LE3j0CRLCP+futeOer754tp89Tf/Wrl/zzYIPRdEE3F1YS9LCeadl+
lOP5cF0DJCVrlaN/d91xFSN9SkbnxLmzjsvSEK+D1PF1AJwj22plj2HDDuef8Npp
8uqyRaP7mFXQIniIAUaptiVa7saDDjv23stWzI4grCw18zIMehT1E284iiyHFyn+
h6aMZRtQdbrBbVW6teNFKoVtQHl0b26yhlGEiNzdMzH40JjMbcRv89csYGkCjVD4
H6SapbP482F3kRpL6QcnGlQGfqIqFsI3qHb+Wp+L6eLLytOM0NdgrbLTLKRue8eZ
xUaMtPjVIgrJIgSTLlHrVRQWZwnRKvC21cjeDLHkp4qcnuLilQrupScBvE5MzNUt
eo4dxrBDpqqssX2bZogJj8wpAElBde3kNTUEr5tPCD4HITt5rkpcCQAZ5Zti8Blt
NodhrygdTBq1IgFwBZJUvaBFYOIW7PboZMKDyuM46Ch0dwweu4thYCW/CzKvacFr
+OiAK3GmV+l0Pb3dVRIX3b72HaIpS5/+LDR5T9bFpTG5wMiHaK/yG1INVqzRDDZg
VRBYoreTJShYtUap92s95ZbaRFVX/lrfV4BZoqxhL1YM4Uj2UkEoVWZBz6l9wd1Z
iuxl7mSF26g0IQSbwRMwYV0lkm5F0RbpBeCQBtGEpwUYDEPoL0JD559NykNyYtrS
LiBR82vKoB59VQuMw0h/ho/ud2t23cAuHSjRZ/0C+tdiYnqyHY8Jjpb4w7XyiJiM
n5SMNZFpLw9nobuZrtBDbWNsKPPLVVUnnBrf0sGo19UsOgaq6cPAr0/GL81H8Njv
vUz7Pv90ocO9K2yemxiIG39kWyc1vGvelkFMpzYUoF0BWAjnFSkSVicEjrymlZK2
/CjNIA5tF9vq3/lSNB7diMiFzH6Nwn1zJIWf030gv4343wK/etq5taapR7AEEpfa
yr9gKfS1KrNYSomBC6IEc90K3Qg1EtVudUoynb0U9twvOsY4djPWr/5Uz6Fnazmv
En6k3oy8pbwq5tnmIGHhA5RoD6tnEmb1d670cDIaI0O1TNeP3d46fmoOjBniVGyS
f7T0PBi4akxUPzVpVRr9SGxjT/kYjzInhelSJ199Fv56jrPsP0NPKBNk8NCOrZEd
omb8+dnuri6DEx6CD72AH2ff/UcS0z0Wnw8+WVBkN8yKNQpsL49EGmsdrZFQNim8
32RV3x7c36pjb6G/Hm+7QFovoDCOI6QLAG+G5eTxKWgFFo2ovklHh27nHZ2/NSIF
KvhKzlqU5gzDsrgCjR+LNLst7GUCTEoMSNZlKCSd02UlTUhxM4Ms8+Yr3EWD8GvG
aHqi49fRihZwWv7DOxQBpON70dBHKyLXyiS0X5wO1yXeYYSayCJlEPZXJi5X2stt
u8mSEAo7aOBUAXSSRuCkClOG2JK+JtIjaH2Q3n0yx5Bk8Fg5TJqDfClYPYwNGmqT
XbtFrGBSnEK4V3hJJ4+VQkJ9XvzHI9GJywiFEsgRI4V3mA4hT1ZO3+s+7+vnPy0k
Nzbeg9s+W9moaDKviU+MGoAMJzECIhXVSVYgqF02gD8d6+FDVqeDXYazvEnUOai8
ZOC0d9mFXut2oJUaeP78d5poXlNL1d9gafuU8eBw8lOvCHvmhmnazihUpx25X53q
hciJRD0bwT5LfC1jCcuE2l6HLL0sk1dqAbpUPGI6ETYCPUdR5nK0uK1jTdxWRIl4
PBlPoWBqJjJTUx48ZdXfE1ddM6QmRLnoQkHiUl6I81pag8bl/KU26BytyWI0P0Hg
Bvfx88tD0hTjzBOJWDNbT/mn/68zztI2fbDe6OaalS3SalyQMCqpK50bLtVXYVB/
/9nCwIMTZ15KzbfI1b2/NH7/+G/DnqKhPdCPz3TK3IVYpW7l0QsBylLqK8TiH5En
DDK+BcLdn5++s/Pp+d37nu2GO5C92V14SP3jKXA3bCbbZZUelK+mjBPjUjFjiET4
HkjnBBfzd3qZhK25OfaOZKwHkyMeHeUYAygvj+9ha2hurn/fbfJMAyzfz432qbMG
04t/We3z8ibEqMhG0hZLFpwaLpEqU1Flnv9O1K1Gom8c3LeDrVEKPVCxITnij5ze
CYnIhQQ7gEdLF5E3dm/btleN46+w/QIEy1NWdv4AelHaoB+bFfu2fQIyTgtT1Ewr
gm0B8BQ2Yl7lq28UC3kTzcgSK9wfFJl73sHaYLz8SQ8cyS4JidhyxoL9oiybbBMd
r4fk7CepFll0b8J7vrG7PwZYbGuKVFYicRJE0ueUj4h3Dqbo+9mVR63ZNpmG2K3v
0AsWI8iu6eShmeNUGVWscAR/tTkvnF7mfmGJIMdiGMktqu0Cwbk2FnM0RCCQXRJI
eTIIXgjjOO1gLKom6xJfUoRd4hIq96XE8F1W8ClNWRfHlVCSMgpCKDzWGZLnkT8M
I2KM8DFtS0sIo83mL6VPOnzGeKqieynBtnL3+JYHW96GgLWhQzAABzBZeLudJaiK
MG3zEzRgNGGIHTdEo188QMs623Kn2nYMVS0oPT9shwLDjgYQzFOlG0vLLjRnuEIf
oAMIAkKwx/5gsSQd6KiriLeL3UIM8C9qa3tgCnydfvHc4AVGbdlQ2Bn6XzvpuoXR
eN4TEhl97zk9/YWMBvc35r7Zkn+38cHs0IhC9gd11KgTnzfvkyCbLFiDkpBmkobD
aqark678/EqR9TaNlSwp5yTEk1DEmrA7U10RNDJ5bytasu/za5cxut2xBQQBM1bN
Ij3xeUB/N1isoCt2v1AZH+3CunPvXiFm7iWugVU6HlFSsjXkuC1LcuqBRIjKP/xz
cg+FI9nJX2X1ChKn3adlFt8DC45uiu6yhQnAB28GF8oH8atVczYavCVOshzasVrE
0MTyso8YdoEyP4WjfDEernhBWay1oGrINOUDodLjnYwWwT1nkTH1//VN9duVeNML
+zms9b32CCGY3lcc81eefcC8D2Yw+V9YD9oep4j2PtuyJiEr/VlRiFZsrrHoTUEL
fyuL8kSy2Yj95H8t72xWgyJoaLBq03c2+1XvXkAy3CDtkgA9GS4bRsf3bCxDiYxH
QqHmBdX1odASx6HE62+V1vLLvg8GL5t/LAOEL+GEJ8UUyjUIbia/s2doxc1XF9Bh
Y/A67LvrL0GcSJbWb6kv+Ng3v7PZSilmDp31RnOx+wJGQcQf/Vof1Hesop8aNiiH
sZV1qhsHldhye9Uj48/nlnzBedIBtBff/a8KYwSoxJDxerQm49b5SJWBREU6rurZ
zSUg9EQKqsPQB4EpIGBFsxi1/aEY3YPU7TproTjcBzHJXGth9W9Bbvl3oo0+YH/X
6rK5pRn4hLg3OZU4XP3+FN3WBTHxGH3cZ7tIvx4wvFbQ6OT1iXBqsQay0foj3LLu
TmAkb9+TphFODJZTEn7PqWGxmEbYYJxOwK81pM1KNcmoMlt2xnlMXZBHwEoTW/vL
ko3u1NS+HzlnTpvxtPnXCgMxZ9aLgoAxO98CPGjtRg58KlmWqEKKGpasScpsYCIY
kXRk9/WAJ+AJ/qkQ6yFtAiGrKfxGL+LIEso2nRw3UTvQWY3fcHBIrY+C6zd4gdcS
r7qCM4fJ/P/YP8kqmnYwgZDH886ESdYAKOSOkJsYIEnUZBH6PPhs6XWI7IL8mV8N
yGBvpNaWtFUm0/EqDFbnPzDvLpzWPWzeJFcv6XN2rHS8cnyAoMTgk09XMIai0FHc
BikQcunLn55ASnHq+Sq5Pae4KKgs1xXemqU6M1618oLlfgzUUcwy/A9bTEUpHTkZ
cmuxQRUQRaEabnJ7dUVEKWmiyfaSDiIfEp6JqL+4BFULp6svUZxpKcCv67CBX5Bq
E5YDy++HQf131Y8DQa5lz7jeVtWU9B3qNgLRVf8dD94+LSW4d1YTMOFB+lQuwYQH
oIoSsYOb0XA6aDkayVbrYVJQXjGPHAHRyFF9uGdXIZhIObk1SQX+AseppV46HcUL
mHVmf+pWuC+qLZoyG/RoCTyBKto3BieL/816HeGyUvQkGqka1sEMrWxtF0al2UPa
BnX1S01dp++spYqxkFgks3ix5OUngxtiV3nflctWFZ95zIuASuh+SU9TmpX/+QSr
D0ttHhbnOyQrpX91tjCyM6TaEEEx0S4L+Fn+w8+Ye21wvrAA2DTAxXxuBhnXVtIj
7camteLzanq5R2AGw2ki+HRFRTpaIBmKxIA753cCERC25H9aFWQKjZgxQjV0S4xp
5TFTQxuN7gX0tpjYLBzD7gsL1X9iOSYYwW6pFHDF2OgirrQ9fO0iAkLubmC6b+nT
ig58EqptnWxPIFDeRCl1wOXySYM7cnEYwWGg3wvj7rONNRrKWpCs/Qq4h3YdEXVU
h/J/92ULWQzQ6kRP3UazxKCqOKoqb/sugUkDvxt0eKgiStjvUngW9pA8tjOlPhTl
PUx/K4o9lWZxR2OYsyiQ1RBQxvXtIm67qPdHRNRPCmxRKbUSyfBL2s62ShG16W1G
/hiiiQ16f1p+Jnqj2QRen5tgNxrg1HMCBwwHR8YQR7GolrswXv2D380Br7KY/r3y
0OeuXZalgL8/B6dw8gIZJwZ3C5jTlM8SU8hTTZg34OEoku3Bw8BNIY6JF4xhyVNT
RIatxskX+a8is+t2SIyitIC0SJ0PMIW6sR+yHJzc4CCuNrp1zyf90xhM49HiGYpt
iziimoTmBpEmQi2OfznjFt+gPMJd9Ax52W9/G1WLgGydEX2PLgSlvGzahwJ8Bis8
F7gZ9oh66MuhBY8r7SlIWp4kPAKcBaRZj4kUytw9hi4Ee3yUBEKtBDIrz3O5KBfH
U4NSqPZsRE7o6kPmiFN/U1yNbhO2QYMH3RMakRydaqtBk1wVY6Vi7f5HFt9MSArh
DiL4MeUVWQgfQJQlWwlhb3zuwkOn4qW1UcoFdnxCgmm8cUpVwcWkCcao76zD/5Mt
LEiSddPaSrYWgxsPRo2Emwm6Z0cVT8Cstx72gJSjt7/O6u+SAPN4Oj+gpyFsqP8Y
3oElv4OkgepyWbBq4aucgoc24WWn0yztA5GjdZAwADqaJn2um4LcdYbZNkK0lMKo
eyJquA6VQbverr/p+bqq6FHkh6w/CRuEXGhTetboVBIhtPOT8EKIOovdpdyPjuMn
j3LJihMosyYVd1LJXVmdkbzwbngrmwmK5dy2BMuOlwsQJU9klbKxMtl1a6LgFsFn
XSYc7PYpKG2OoMtINGDFHIBPstVP4IWaQz6oPRr1RXZQyRxOPZGDrayKz8eo7Yss
vQMn7CxfaFutOsFDmRBON1ZGvEfNbh3vEWjxM1h7VSQT3DWqXsbj0y8gWNjXQbt3
H4s/fpabZEPxjnsL+MyDUCt5rEmKSmygcz3FbYNauCibsbz+adbqZzcEZfTGFxNl
7CLyUE2CoI8hOOitp3Xxz2M6lPQymTNvaT7Sen7A2V7do9s0NOZhcrFtdE/pcy82
ewAFJkx+n6ZqAxybmObsV9FQbioYO1wysHTUAeGE4nG6xMrYaa8Iw5CVoBka1moC
hO+dheYibcwYxDYVOkD9FvYun5CW2EgE5eWw7LINYVSUWBzIZOXEGufeuwP7fg6w
/+K+GOtoA5iOn7Z2bYkiXuoC5YHkUQuL0qQiHhulvnmN4/nwUkAsI2kWZPE7vZ3Y
AYkOxAKKrxKc+FVCBlXcHBi8sKAURSMA7EWFUCDpSJJJn48ilwFV/UjL15eH9zhK
giwJfc21194vaIXjZ/qgg9X2q2LPpLHt9QbGPFTVx+RMazTIbc279t2bOMHXoKxJ
KxpF3TJO/VqZoRVGuZzXMKqUHmfqKexiJF7ZORB8H4dRQCeT+SqGzkwtoOq0N5jF
dzVYNMFMoDO3xvHNkbiAM1xcnYOpL0ayhVKBGlQe5ifVMgAjy4dCDiHjdAWl0wrK
dvfO8WZ1YiiGMtZ7B5KFPRlZPYjAX3LgUKhqgF+sA/duZjC0EUnGI1OFx2k7k7aQ
egRStr1C54WTMY85OP/bhkEDQdOM4IUl6IIhgjGi7mNuIb9Pgnu+XiyWOg0J/uLx
XJCKvRIyQ60ixeFq+EiYSNlZ2O/VbXv3AeSBOV7z9Eeo124KMIwkGHsbweO4AG7Z
iaEWk9uP9Edv7YbOF/r13j/twmaRnEtnsal3VpgWG2rCzSng2R5gLnFRDMdXJht/
5CeFJwYwly+ujY1KfGbZy0NYCzQ7iH0qGps6I3f3ldlkYb1oEPOapSfzfmNvupvL
lWQTIxJKcMUcCbMiypswSI6YIoMdflBjDsVeC3LXO1BAXOFotThFZR/mwuijuo+h
lP4aHWfQeLD/nIkzwLohk9ymmWCBHIbUfO76/Fem+FVWM9HfQEj5aUAjU5xW2+z2
yOMd1E5SBShEeygIhsVI2Drk1cS6ZhGql9evU2O/hx5LcPNj4E2fp3cL5iXC5JUH
90eSmL/J2LgBMCBr2PHqX9C0ZgTvfsRBZirWd4jF4DVRoUzY6lPSxZN5291hmEA5
xOkFSHmygpvVYvyH02XKE99b32P1t8dGvFi4IodVGKB5DSx1PpEatlllR57XB+gH
2POuIFJBwukyXL2QwmJXb4V2uMzFsH67OdzywSSN+FUzrIhg4UcPT6Su+DDRKE4f
V+xyeN35Ju/UOefTA0ycayiBoNyADwayUxUmqYREhyIziVhG8cHcPhxFVO6sIAnb
xqVVFGbSYe71PO9+PIUcrg5W0oHJTFL2CPQ3cybiHEi1XZcZYDD87ouUo2j9UZcP
vRrIv/LIzVTdsvc5Wf90+o/YMDZrdnadTBpYbDvyoHAnEv+yKlnkHATtHM0t9rCx
LkKSFNIsToaXMkdyJUAf65Hpwd4hyQFAq5tyHuw8ZWwl9aDSxBQ+ifnLvxr1TNEf
c0WQF/BHGd/dCBwfnCxwlqIRJxxa914kR7nM4COpwax5SHZ7vpl29opQTlZBbAZP
+IA9dCAROGRcaJ5F+RK+AGmzVbIKORfOrYrPLDptCHVy/f/Nm6kavAbDvUOhO58e
s+QYkSFIWQXqW3jfADxUaqi4kaGTZuapx7h1zn1n5XOfRlZ8A8uc8qICXNMSgfQL
fczWHpSGV7QvKZ379WDMGHLELTjPOXclRQ9XrIhisDFtEbHqG2tEXBucN9R/DHET
OcioIDIbQ7Z3sc4TAl2ml13jpSIFlBilpycQAwVXc7aLuZevWpOCEEKnoNWvf7qK
FRLInVBewgPZHqSdkrK6B+G4I8xDc/aGKkzPHdjKLo588Bk6ZvWvRxbJGJYt/DLY
7IatJQ6etqQrYJH9m45h57UK6+F4DZCDY1iC80iiqG95DV6PZte8izcCutzFJJzE
EhXAK0T3ePn3tl0/TEZVtQTVPeucf3+2BiwL/r5V3Fe43k0U9o4j+DH4CdCl40A3
bqtfGZxqX8+QsQ+38L1aBeVSB17yJ7u3L+hyR5jlBMoRYb+jut802sZc/ZIbLIwN
kQ7D7MzZVgFBPFJXeSKfhmn1AgygRMp/nXtlAve5oebZVqGAqv+qSJe7w+TnpXDw
nV26tNMB5N8Jig9vRjsQ9PGWgQ/tG8CwZSeVKMgXRYrwlq5hegfgPMNrJ7ketbpS
GjvLJahU7xTNFY+24atG89W46DNXZh7F1XT8BTB1oSa1Ggt1PIAxt1Txhb5XdyfE
VaxbD36Gpymx3hyAYpwz6CKfE5jWulZTYnugZUQvMiaDzI1BcJ90mNUmIxL6HwaZ
EInNF4WLid4dqOivtLRj8ok1DGmgfXiHiWUy7GcrSrhVNCCNV9cFT1beZG0PiRWJ
41L7VH1Zv9ruZTu9zRPopq5qpK0iXb5cT1hNqAJFmmF/NgYMHb0+VDxEE79Wec/i
WR65d/b5zt1/p3Cv31nyXGEIdHGgw85PrkcZadZlxLSuxt0W0SvP+iAV7JBif9Lo
YZd3lVV9EA97Eqct42CDQxs51EswcmxhJdTajOnhQI5UC1NaHHUH9OY761gd/oe9
bokR2C7idh7Pj7924iLqN2/RtRt97iiyLhkLwW2VFf06OyQp6XBHabPBU2P1c56y
vDm3s1TE6yMu6orbRSA33C45/xAdLOPS3vbDow855FfJdAzWrOzYhtej9YH0p7mM
RmbOImWKwKvkRW5M3fNeimfrK9+nnv7s7U0WQmlabQbRzydWTpANGAcosnTYc1Ur
QYy5REhokbEQDwSHzloBAecv4XUXa/jgwaJkG/OShSJSZ8+FEr3BI0KC/P1xcpTa
FTSzZqxCb0+XBHuAATBgfT3I1slwvSpgjrx6Ow3OXPtqW8lB0nKblNgAarhVRtWa
JeB8NUP6LjX05TZDNHJ6rWbU8gHsb4yv92IxESjbStXZHBkrBgFAYSDbbESl1I2+
3aoZtXJttNj/prST+PM4Xytst1TkA9XcJHagj1F6yLuNqIRsEQaGTTfr70wsgkfb
Y9PrvOjEkl/Xf3Hua2C05tC0WhK7fX1Dc2YANpXemAagntrr94iAhfhzFw2fg4o1
+vKvspFypw0Udx4undsiWy73cCmVxY7E82aL+IAYR0bCS4JMH+7pItG9LGGivJro
dveAb/KJTunZUH/VZMb2Qh+832rCuqfQaexagw9fusjMw6Sej0iX+JGPg6INmrfZ
fsCt39VpXHpxV3Gj/4ileIOicrqVKnwqmjClpaijpby+vbD4U/o8NSQiobEC6FeX
iCD6XL2kol6xVhvBLHZT1ekvjmCI61shoUUc4wG+nYAt1BhLHTvV3oRI+TIVOQM5
8avPsh68KD+wcB+esYSi9kQHvfSQk6mU9wOSG3zTEUyn974ImttzRm7umNkAYTw4
aTUc3j5l5dNrYhTpzsZxyOGBgDAB3r5BlADEPgsyCIHxiXZ6y9T6AyEJrJGQW8aA
+Nj1Wwih8TXwyDqqZFVnrwz+2GvReJ72uvpTFjirY1Es3yHW3qZKYPkdFlCsgr7o
pjJa59//W2PFr5wmasKNBmxUmZVwPaX6FPHSaZJ8vWk+awFiun8wt0bqS9GSEhLj
5oZK4WuLy8nOxASt1xQoRiYY2DE46vNZz2cW5Fsc/J8KrlJZREs+e/hPIbIDEJLt
0RWeZrMa0yUo6ZWmJyySCNb+s5PzD7WKOzA8HGwL9FryV/MomYbeYrsjPfk4rq0A
Xpm9urEJaqxoRJuk3fcyFmELqnjsr30aODAJIkVSnSAm2tLkT/WEdOusV2q/wWK8
PfOeD+yCpmp9xa/KwfvgZKO+ihXCLezWLf0WXNGVt9k8ZcRRjR2DU0eAh8ePuxSb
Cl/Guy6EmkXvarb1kkuIFj0nLS2nHJ4YBhpvPde1W/LVBAc1rJdKOvoDXOKRlWxe
To67cfR5UGQ0nG1yytVM8I6sGHnI5wUDfFrXjnz0t54m4NyWelZ6JwSW7O5EUPyo
6HLQyUjfW2EE0Ka8/BuPnQvAb4SdyL+LjYZBP8LoqTQ6oLR0Xq4ZmCEocqBkLJQk
lfk10IIqeVyrnsU/5Pp+2g8abtdVrFsk+NZKdggpSBkcdNDnpC4yt/73XGw0HvNK
iW62wR1+pCKABjK0ST6F8aH/MkB+HV5c5zdIrs7F7zJGgm0RfM2n3CRC17uMscpl
KDPwUKuHWvprLio8GCRIASo+/3iXmXat8PQgxol0kL3ytGdjfb1lvCou78iZlL1i
BVvUyEeq4W2xJzIBueavCXeFxW9JKUtM91vr3Wz15iqDo2lWXh/bZFYRJRvCpMRr
TjdGs31qUS/xGc/D9uyMg+hGHek5SnkyiuHzC+ewzos3pRt8CcSGEbD6wkqLh4/O
uB06e28DKoy64CRCmoXSFCo5YlmU9O2zm7cvzqlOokYpok4D3XxictaLxd61PfDA
jnOk6WpJ5QKf6XDZGmoTmRfkqfOGa6mYIWPTdKklwn10NmQhPw0i6ck5OrLYsjhs
PjlT0/TgHe4JohcS/cVyDcO1RKFlmnKf3N8TgzFXV//aj73SF+OLw7pXBDT4h5Xu
8nQ5QUvRbL80ViKo9WSyKN8IeYz+yiqT9iqqUrldVUzpzqA+d7SaofY5lEwo5g2n
1n13GJU4gCGv1gz665zDRnUTkcS1VcRyNiMRetgM5XQlRwBuoY1jxb0vvFJ5LRfH
9LaGbXWSoTDUx6f+t70IuxZ1tUK3BaGqpo+3pV5eSyqDnZ4rDAE1uNciU/tBpa5F
OceWoTLP7ysGekUbl4J3tSrIUmPvrrPHy5+8PT8snSTqckDMR70jfz84hfxr2Jsk
IvdcLklIUWjFj6W3Ys5mGv8UThbiZhrJnaxd5J0PMC/IFLw5yHdBb37U1OvywoW2
ZemxahUxtzGUbY5nbieY96oyq/a1L5ANS5YP66BqpErYtW4nZXxUgx+3t9hbbLgt
DWLdFjk0OotYn/HBAv+w/w4tTjRhDoLU6UrR4gmOGe+RtCokddfMN4n9hX+jaxQj
97ReEg0qFGcAyVTGJgaJKRmf/lFxvhy4uieMf75kYxRyfdMYjjmY3STnlU+2wmNp
ANjckph3De03hBAdGRqNC01ASfAjGMIrn3889i8sUW97UOCwFiuDaxNnuNfNRenn
kPSZttgAa6m8TW3DSHrrOtvU8QKp3zx9TRiNsgXBkOCSvmwSNpZL5Ms0qkvcRCyS
M540iBuSUqZ/257ZkHHyOn6T9AhoR581dkSxk2qFPcY74Xu0bTa5TJ1zlKjBDGY6
0GUZ4x2w+uEfi86cOP9vSYawqG8cM4yARSEo1++6V4ZSFnuxPDails3tqitDXdec
jkisTqtbCw+Xw2Czc8gcYoPi0/+8D49SMsunfnaHpEPdcYxHePyA/tXICZgbTRYZ
mZjYDLKUcfRP92n/I6GceosEPvwFTIGw6dKMkAFiOquOCzsSar3VZ5dvZRsCQXol
MVQaPgRglXy964vk6YuBv2p97QAcjApKM6ipxfAFX0qDwXI441HWNWFGUq6aOsUb
1LTT5rvGjVH534khw/vT+zOC+tCn9jKwXe0RtmF704V37PeFKZQbIz00VFtmaBpR
Mi//nceY3GktaI0rOUS5EJvvg3AEntGJczE3Urzerf3zqAKf2OuCNDdsFSKOGOEk
dYFS4wzYTnjsk3jxTdOf7G9YnSG4VJy8y2QpHsmrhMqTvVZO3Bixq/X/xFidIvuc
SQ+nFl1NFsAyWbNbm+/ypU0csTBrCqUGmhIIb71RgCDNtCF1IAITNNfCKTeJ2Bpg
GHC3elpJS7FFB4L0CbvEYPDHz2+8xLA0v+ldFNfPmOXau2TexLijJcQfTeGSoK0u
ujDpAst27c2S0BHaP6m+NvWFwgJmB3+sByWONSfe5IQc8b9jOMfOmGbidGDKjusx
AGXGcRf92pu0/1c9iE4cXy3PlZRkM4Huky2n6o/ppVbaMuliMHfJsRTwtjFzfrOd
ykjIRcDbJYz8+hTo1ujym9GzScH+GVTb7cXfe24knPqn5felWYbxc5OX5FiU8YXj
qxoW35wMn4/u7FABKsJAvhppwmmtcv0p+AgmayYCrJn6l3HNB8RmSHXhqTxA+TSw
E51ic8ojRp+s06efHqPz0xxdIigxzswa20OWPrXEvnSg/YAmPPofe5Tm9AfSURQJ
41GU1OumjdaN4zB9iRxZvphC73Ls0aa8hpg+esch+Zk8mUQwEckpPDnpRWs4T4f9
j4YrXLx+ZJ2L7Iy3fPoK9Hi8Z8UZ/2miXQYJ/bMYLHRFwZjGXyN4LnXfblstJhRa
bp0pBb2cB+M2qwoJgWmClKmCUeqX7OUE5MlpUDJ6XDFFlUyr/EQe0+8Q3Kg6rBAt
MS21AL676l+lQw2vUZNUavL+ePTqJOi3fqTYEtASDPJgx4dh8IPiQUSqI765uPzY
2d0Zxsj6dcnpG3SPEWj1JG0eakO5Y8aAK5zniMcFe68YqMtP8RAkcpXvNf2z9vg9
ZU6QTZzoL2DFrMUGkI+NwelMe09yZAOaFQ+1zMGtRekr1Li7olrh402x2cmbSeqg
rJxcdDrycfD8RperKGRtqBBx1LKaSh+DZY/k16La6B0+zx+GRsr2FgfJvUM1u6KG
N5cuoUGgqGhv7fb4vUt9Hae+p8SRAXWrHFpvP4KezZ2z7DfpixDb+nnQstwearyu
IBOjINZHSYjPvg3ohJOUPIzoNdh/lAPLv2cnonas9YsJDFTL+QQCfszsdAk0e3oC
83UhVUu+pTMZVCt/RNDcaTvkpxkSaoQv8Wo002FlDnBu4voZjRK1uzATmcPDmeAW
Ro3otTvmen16dxVo34YEvv3/P55spUtKlrD+tlgtdIJY4RUSYsgmZhCNRU9cWC24
rs93gwK0RYw9GkjlVTfaDCREkH3tPc3Ne4jy5c7o23NwHods0LBL0PoTe8xYZpKm
T8f9eNo+xZyAn0GFpQVApaY+1N8K/VmJbFKvtCSIT67Ecr5yVTdxvZsiBMRXFmnx
SzA0FqdkETIH4L1/EO8qnv1HaYqogSmyX/NVUFYdaodX4DPUGGNmf/kJCPDgRgym
Ijvp2Z7ME2i53WNa6fIIcVJX8IRbgrhd0xvXWmIYdnFRN38hEMfwLLv60ywqUcd3
RBFdA3xXo5cpbqhnFbW/OyniWkfS54V36kt5gj7PnZ67mM9HBPAQ8PEPTkKd/sMR
VYsTeAa+FeHQrtyqndKrQ7r+l3GH9Szr4JkQbUf7wSBuRDvSG0RM7PLmiihDtalP
k9u0/lzmxR31+aJSuzmBYu++pV+GoDhOIr5A5KFKR/bAKXLqNI6DO5j6jaCsUDLJ
8/nItrNTNcGZ7tv8zqX/4SVXUhIywQYW6jVEG/dbMVs8yHy8E8RiS5ZqAA9nxbA0
KAhErcbwYG0Kqs9H868umhEMXsRVw2liqF3KoIzJeh+MAKebFvMvBi+2IEZaDOsG
62kki/WeX2ZEc4XuNQJOmzzv9NylhrtEX2rUNrJMJxIA9rRokE/sgK4sp+NcUpwL
isIVyFmULQylWfebm0lj6BAD2pBNWcK4S6PWaFbHeQTS7wU1FVwv1u63zz84nLdb
WuojFp7FkFPEUOlR3iTNGNVvP56IDgLmNra3iW4wiXzeXVVUGNQHLI/meoGPmpfu
8sAe7+NEDTUm0xV9exLbWUoq7njHXJY21Vrz98myHKsScv1PhCIy/YoUayB0rB7V
i9O/FKQiVi1N+Ny9Heqd+ntTk2jQK8/K3GwJv3F6t8zJV21xGKvUxSW6h9L7vtY4
FecCe9AK3yPbZ35rLrRHvgEwD1mnTmSzo9nk7dRLDAUdg6Nli23v84zcu+u3WCb1
rd8Iy+xQ5XsIp0kWv5BDt6+zvsaVlnzd5GG0eD16uK/7v5XfPQ6WmJlpUqCqrR6I
wxcP8/AVBYUGk30Q8uqcVNgH1NA78ZjQic4RnbabQ6JpflOiUr7tRj/0jt58E+47
X8NlR+2miF89coFyj4LGBMJItjWtGqii8kI5bMMMk/Pg5VsQwMZGB0DLTLum5zOb
DNBgh+19+xQ7IkMP89fG9ElbjxUtJ2aHeImMAQQkivEJSyGo+FKEf43Es6+c+ema
eAuIiILFiXvOUvKGUV6Ffa4YFsQbQRnDoydwnIo1I/570pJB5ITj8tsH2rmulLBm
uMLY+7WLSQf+tau22QpVwcKYNaj9cx5F/vkdRxSm2WRKonAPC/g/9+LUXKoXMdMi
eVHJbQAaNIW84rQ2+BquY3ZLrFX8WJ3dVKkNtLryLL36WlrEMNJFi5i0RpEaH5Wr
vkwwBAuBdRVkoreQnP8kOSBZtr6TDqucXRrnYDu659otjV88hauBLN8TOKT46E5+
y296Or6gn7z+NnWVIXjET1rweY8D5GGHbdByOsHr6xywugd0ft/py/J1v/S6CRel
kotvNKebpjinA/etaMby+icX6/zbSkS3mL1YcMPHeqBA0cnsL9zFzFhpgxAGHwF+
6D8XHasP1DshXtK4yQEJKc5bsD1f8iq+zOlCbfkuvDu4cOxhuLZn92xEVKaIx2fe
wrwdXNpjsCJpjRRJe4mm4gB1p12uq/AOXj6MIfi92sL4SUmYrry48BsuRGR5JzxF
Nndd7Wvk2PTA+3ZvM/amT9SnPan6d+G3teS3Pr+35HAViNAot/tNSIYp4DTiuk+7
1wSQBmhqu5lAYratBpJpQgYIbXvIYM2mfcctNH9rGOe5bFPqDufr8Ht8GoFdvGPD
Kx4Zfw+dvFGBtP4KbE25NPX2RjFdqkUCgNcoMORoHtuheTyrzStpllbc/wl9HwBO
9Hz3AP3PoO8pF/CxSc+aTByBdwUYjInHY9S5l+MtxsMIEqae4fc84EZg+OmAJJkG
gKevulbdW2kHUe8wX+jf1O59OfqNSJgVW7hEv3XE/aw+42prCr88Gfn/ZvhpQbt1
wmpRZmdsiyfmMHnGcWZVUva/fFkfVNlO0KhjLf6hZDj5Q+5dtPMsBxHWVIrGkq81
V+ZiACwBv877zZSRmhd/zYAhjgRiE/EzG9DMSPtdMFFoUbapQbXpWXhSwHF6ghTy
8UASPN9qpHWgNUyJ0mG+DwUe7hIbADW6DltYA/8CE4yiOJxTmP+eS7oeuy2yvLq/
95lUkibOpfNsk+AgJxTh9qenamZwSFvBhf4+cmpSXNpfjJ+TI3xFyccfORyXYGpZ
0KSyL5ByJ7EWfUfpWe4oZWGBozmvTfeqcpinkJ0hK+SxLgWhACoti2K1hLt3O+7b
rxgGuE5NOZcZK0odweeenk4N/R/MI46wCwcwArEiu/Gq1K6uFf2of/pvu2ZKnCdk
gRYWtGreZ02thu6n2l4yeck22OCSDdwwpKZ6lDAkdVvoX9mNevgKyi9u8mGCmFaf
9GUjVUGI3Ro1aFlHpis3mbDRdHLM2vph+IleWwIebYWLPqLBUU0YLI/YFoBRsyxs
yPUMWZID95S+qGZUtHLSfKG8P70UuTZ6SAv3tv7IdH6rKUmh1pLejodx1X8i+tjQ
ibxUn+T+Vf60Llz0jiu8MrI6IxMDg5TGjvQALf/8J0r7fpWeZBKyE2lss1HIIX80
3WZ0JhSaXHahyginnNNHsCA1C/DmTz38R850VZVSGj7lTuHFDJh9+jZXcqVjMr6Q
c5qf+tUgxG9Vp8gK8/cTe7IFLgI7g9wpZjFx4cJn9aT+Vc0cBhMQziRoxsLtP0cK
BOIH/RvGlSZhOdlMcguUxFYfMOGpf4WTAq2VB6T5iqdSIfOE7ESsLuVYQY3cx44I
9O2Jz+Ie9cncH2re9XFddm5n2NvBMHSJKAt5vWfDYO3ksirlKW/cFLbcralfM2ZC
OzVprYNTtRdtSzQmwCDdsR8zW9wR3pfqPF1t6Kpbn/RolU23yNRmBYU2xemc6e3T
rOHezk99wNyGUYvB/8NWdSt41o+yO1E0J9UEc3g4Q81vs7/E6FpkeLb9DmxDINpU
MMpEY8YBX8CkZAW7GMwuZO8EgJYa448Ao23UXK8ch+V2/1QYYGgFHW4NJBk5tBZK
mkTciQzM2nCLf+A2+CwM7pJ0WjmZBhwsGDq2tXv8uNIa0lBwHm/JrTI2pg+o3OpJ
qkFLS8WFlnVl+8zWGGTTcvM/w0odScrAprFNCu3FmYcNgfvEk2hw9RA8rFInY7lq
i8whbqtC1DXs8yXq9EwM9HbYEnN2qrWsDfz8R0Yz/pxOMOw56ghJao8rj6kOikDA
qvQ/jdJSisH6ifMaAxgNl3peOFD3k3CFkJi6CYYDFVLOiKfW6dxHMVwQ+2X5ygNI
jWr8pinw1VkRQ4SekxJR2449a4Ew11OnOOfFyPZgaUzI7bbwQaH3Y7cKA5VhTgAV
LL6AbqXIYijFWOGoU/qV2EwOELJ7523VesFgMZe9BQhGHMhwJvw1Gaglh4AHG8NR
M+FRUyfwDAtM93TcecHZCkBBKN0UxVLQjX9ZZT/anOqVF8qo6toetV7p5g0511QQ
PsVsOrsOoGv3KLDTSl/reIvUsBALc8QkmOPtedGonXTuxHms9OjyY/qTzqJZIGk1
XA6AEmUeUIkgGJsOh6NqSHINoFmXrtHHhCn+eTLlFfhSvXWOKOptVfmwox9XIhLt
z5bHNs2QxFWiSeXRbohIZOvXgan3XvPQ9zGwIOqdqTYC9dvO1mpTI1VkRC6XVPA9
7MgqZ2N9I6RDw/tvcMEfKfD10dBGG3BUhFas3Z6f+/dgFGMoJ9AuooAuhtZR2FZl
1L0c2rR8LsyDytr8F1NGZXO4VKWduH2nGkSmNFnBZxbUc+Y9fF5fv/QkGn30kYfn
q6xr26iggT2SVq0mbsXHADtweOobIyjKQ8vwEtbllbUNekpQ8DQ5MqSuYh++p7At
i/yis6PF4RkK/Y5kbmu1fnhZUxyh0UzZQnM1pGguTvf5fUm2F0cCukpigKwJX+9K
ipVLy+3QkJF68oZ5R13J5Kf52XiBoWcLD8tNCi+9XJBBk5zddqr1i+/Gzplvfje4
t/YIxPGJv6L3TZafe5H5+otv6mpnliXbZseAVmM8VQAz1DLqSOQkU6dPXpoX4pnA
uijs9tiFtPocu4+aGCa2NZ686EfTOmEu5AtrrxfKGgaGC63m0igh0lnD8DFxDBd/
faaWdRPwdJ+yX0V0RCkatcJN49OAfe8ZSrKc8tBmFo7RrQGkLGmvCCBiUPJZeNvo
w+LVTNrwG3YmPG+LmP6K22CqGet2jbyohslj3L1/5MUUuymsG4ds7jSPwhzCDKnj
vNzhdiaQG6s9MZw9vTPq/+lIy5ZOHtROa1VfLwm0eNZkzyg2pBNlgSde++th2yax
CTcEs7zih3lA40ifywNBJgZTjYcXv3ylwZZTVdtCY7p/uofD0fxtnSRIGSaNRckl
So4RlFQ7Ym2GMqCoYNFksqa0YWPQ9qxcYVmhV6qOQsdqjL1Fc9TTlZVd/8OnaPMN
YVgsRQkpJpHmB1E0aKH/4xiX76x6/yhexJhHOLA4FDnjkUfyGmBv9BEsVs+hYUdU
ky99VHQpKTsIkeYCcoztnwj3XazDtiklwGqWU03c1WZ8W+mTSiPW8iAUWfLzZyLE
WWxPQLVwjOpVeripYfkU8oVA/iY98cxmXrxPCnXNNRK6g3lCDkTsmW10m1f7Iof7
rSY9hP7PU/rNo0HdmoV/EydPKQ3/4lLh9VTcAF/vGm7+UJH8O56yNc6X460vCIGc
SPPTa1L4jqfrRe/tv5vfF0F46kfvxq/6yOpcFYxcxIC/2ja23Q/XoTpJcm5iKZED
Lkj2nPaxHPzmO98tSZA4uMKgOUgVETR+PD/T9lB+pQ0lMDET8nUQk4TDqUFqvTXH
c0ww0DLqjcHrfeo2CQUo/gqt2nW7uhywIW5NKne5v4+f1f+d5BAGW/bULqqeHCBF
zuaYZ57Khw0n4qO9VaKNnTl7HrTnt6enORXxQ5E3VKPYke0w4UovOgilt7Lkpyzb
FCX0B5/G4WlZm+DQ1VARWlHQBYsFKjT8dlLcERxw5NyevrHbphnSwpI+J8Pugl88
ux81R1e4Ltd/aoFYg3azLBQWoqNp7Kdz+P4ZVcmE/wqfyvF0mPbYGoGNGlNeixBH
p1t4TlhKiOVmxld98leGljNTIZLmVpHGH3F4e4Ru452HpRTvcBsYxZRclBMchaOb
P9Qdl5zhVF+zyw5AcGR3iTQ4Sw8UlFDtaro0aI5HD1yRUe03DnG+aBsgDS/84Na0
V+xhUCrI9wPffeySOrv/sqLDRODJcC9clKt6VaUsem/fL2yvuFvwO9tO+RVeSrWP
hn/OoITxDMgokqwdbqTcCveHzaXPNMnuxH/QFXJAvPJj+DontqYS/zcE9tbeA6YZ
VUj+MeWiNkvSN4uu37C8laHXjsB2qpcqk9TLAfOGcK0he9im+diOxz2jmxA0WRWJ
OdmOG6swWxVZf1vswiWp9xt5wRYg7EzXd49o0kgPU/gAKP7jLS6h+bVBoB9FtT4A
zjwkK0DmEtaxzVbwmgbBRC4JRs+ZpTnLMcchjmS+Fr1qsSBI1Zs2rukGlkXG3edv
//UzmqbpqQXNipsU3QQgHLu577woZzhAZpeO7/DRQSGCiGsGec9lq65atOApwX4O
0PHpNkx7KmAn4dvks4byfDsmjGJNBHH8WKusT7EvgwnOnM3dk03ElE0pMMgH1WLo
6c4EvL5P1RHRXeL6gteMz2qc67UYgxfwj/Cqb2JsPmUnIfDRyHdxJE0H2assZFIX
SpRUg6Uv30k0YAw1IO088HgubkofaT9Gdzfvf8odSjTffCf25Rs7YbYR6DANVcCZ
NVobXMXjZvSh1/fB4Wh0QM6C5ZHuJiiDt/6jLirdp1ghPuAoUTmQ95zviUwpjhM4
PHBQBAtZkglGAd5vMP0/4TAsGSpTOTv0YWvfRtIvBW6ms6Y9Rx0Pmd1LnEQkPLzv
Rg+HmBJMdBVulrl/Aav9X/gBukbxcmuG4l28PWwID+5FUE6wxd3eS9l/4CXH98sZ
oiIchcVWQ4pzZ4gvmVCcZg5tfKj772Gnx4nS43uPsN53KrkZWcCR9ZahO77QXrlb
oTMDXJT5XQBApBPgHd+CCVgKUa53AdApDkHr3dAIwahHPCYNMlX1xFGiblGpX9dU
htl0xjfNgVj3eXlYc1CmyTX76FMCnJHPa5Bwa5rAvcCZhwwgMDHCdB9A2j8BsW2P
xYsH7yfPgTIcwB05iP/+6ZMCYLE876UzpJ/in2ZLKoFPOgCKdMYoO6GHgE9RpB+u
CoeqaNsgOF6X08l2BLi4lmNy24ezxQtpJiK1Y9WCBzD6H9BDy58DhRYKj3UXp+1x
wPOPzYbqSIfPED84s1X+Wzw6XtaStt6IWydfAwQ39lYjwX9pThTjjlUNSmAKfBl/
NmoTmhW1puWEsjNxWUpgpmN2ngpMdsfvkh4CWAk8THnM1s8hGqEMF3eS4vPAnPlP
BmoISqwjyLDHhYC5SnpPdrvXN2C6vZAc83TeVEC4CimNzcVqO5kZw0tQBm22/aJ4
DRUYWxspMgzyEheYGMB1ZX9kZQcnPz09bfyJyMd4lxCEkTDPqsSTKzi4qlSS981p
a7gtRtwbddtIxXWSKJ8kTfgRgBpxgdGPPBZjsb1dRi6QYr+iGTQ5+Zdq+G6AXoN/
x+AKvF4IV73Tu9mqJMI/zIpWjYu2NXmb9q40oiRfH46l+PtCmOsPDxKhx2FHoCGa
dWLZvSQg7UH/JgfonxNaQOoXKFy2Lxk0wdxgXlEA+yRoQ2uCJtdg++5Ag+U8QPQ2
X5vrS785Pt1lCDwctGCAWBFor+MnKGOjSvyy/VmH+4DW+k1Dm95nDIsYXmSqPlmz
1sYykEAzj0cK++Cd3prqKb9uLpZZvEqNNIGi2JDwtErv3JIWDvmild9RtORoxxkq
zAvp3IqLDvhRLnuSgCn3i4pwx94fi549korQkrlddh09q0N+bw48QaIYDcf1DQOw
JAqziHUBBdnlzCkIuryT7afchIb0Bp7HBV3MdNFHwveacp1oS0Tb12JoI6niFoeE
9GLtgEwwtgGXXW/NG4Z3nVwRwg4mENCQOwkJGaZeI3deaaJCqGV5Jh0qGgE48v2Y
/uzRrhrQfklybpHauAqJgIn4ANzdDQIUSYJn65qP8yas0dYafQ8WtZolO47P/fGU
dE0dx0krzspsLsRyDeKyUoSYQheB46YMReoRQ9ORim31mshij++ZTekkNNBGdrb7
huGMap4WFpIrhpvYi1fJ88m3BWQCyTKqLpu3Yt8kbNZjp3e0F1LlDnhKTCWIk0Vg
oGOTzN4qwbFism0BbPQMBskv4U72cqc9i8pOGIXegu6paYzWzgVMeZ3+npC3XY0Q
3F8ZWKiL0oXqdQGtOvUNEbCcs2KWoPnCv4GLLHQGXatm8YV4focB3quEjKt4QsBP
+HnwA/FTm4ptNsdCizfK1FSx5ZtIwS6fE/dTWwap7OS8ZNgvJYQKoaJNJvzkpfYv
r+1Zfpx44UmHHR0oKxxIAjb997F58eVDb2XcykxmadMQof70I52Af9BujbAClOL7
TQzwks23b7MM4VoXM/PqeOh4BpF4ltcqbTgMNf3LeAKsYcykPJlT0zKyLm51Ws7F
kOK5Nm9LMC/JAYD/UQG9wylHf3n9eMfVSVB6/rOqIIjikgMeFgZ/jnlpsB+Mb023
wBvtSRDRMf7j5mHuLPvWGm9Sm7rrKq6nqjAe31H11AIfXOWFhPD47CA4zjqnnEoj
WS/IjJFnQoyYII8J0ZFvXgQCfGsdP3YHmPsksYjpgFbFqMMHANGIL40zCo+aQ0Fn
riy0TWn3T2fTogsvC0Rnk1yjx+mcsuha98lCu+JawWZnWc+usO3oTIaXVeZOJVPM
GlFXzAF7oZ24xg3nP7FiCER9Db7n+aX4KAMrhfDlTZXlUNwt4Qk9DiSCK/3hQAri
3LNsnZ+BDkF/z/fDHQFyxivmNc6oK8h0Pz8bkXz+hfNCj9NToMmOy/XWJ9KWw/oA
2UgZBNTjC2JBSL5e/MfUwEHZVRl88EOZRzAqpDhqsWARucm0aOa9ZFv0RbHiFt6u
hBx2QuKmYjuMYV4SZdFnzArXjqarfneQAVnGzqEOUMjHf5eCmcYNGwftHw7tAtPC
CAFYhyWrTbB75O7OL7cuzMAp6t1nS+nMf2eWHvSre/Kg3p1+wT8eh0UKby2y/fzK
gI1xamRgTfTccTEMb5BBlbVI4LUmGxzdWaH9+qexmq5tIoA6sgFyOGhjcNC+Ef6h
jLFK5EPu3UAyYBFOd+MJUbNbr0nzgxhkN3Ihp/hoF+6q8+kkRWnWZsJbPJ1ozBqK
LiQPNHQiRLrAx356/XvocvqrFXp2S17TFIrlv+dYmLN/dqkqQdQs6md5NmZHq5U7
XHEs3AM6uRuYuFzk3ToVsp+lGyjjUCWA//hVnRa+cvDE8JFPPVWHph5vZbmONpOA
SUGfUY3Pd/q9SQfAGlfQPFpeWLnszrSBJFNhYt0BNccGC/yiT+/enqIc+Rkw3CLr
BtkA0ZJXNypSmzZXsIhFCO8mqsLDgtZ8yPHENcidMUFin0Av8tbokzD8dpVznQr7
y7Y1D2YruZw8VLTW8u7gTZNzXckbzMuBj81sYPegY+5IAKnfMPRGQeCy4+CCCHNM
olYLELu6YRyPvExDGQmXaFRBKZEEQcEh6SFgm5RXGrXkz+/34AdsuRozyAYOKMR2
0jSxx1FjKfwPgedk0BaYHjiodaTfFXFJL2Welr/m4ho+H79ANI77Eza0QjCxSW4O
9Hk5hXJKhBps2K5jG+gDSroRe6XQrgrJWC1MaUA7C14UVYlzDaR89V7PwlRdhYJv
U/NsqttvRnokVuvIrKDHIvPM958RWLv5uPWvF1NCcc60tRF0tPpce8Uz7ELHkNly
/AS+6Py6MzwC7E/Tcu1nvBfgTsddxKu7BGYUpvz4uJsvHiOVi3iU7fdUBm97HBHh
jxNjRrHAwcOvJBB0Ox4dLfivY6W6QjpcroQoKj1MYB88gnHYf/WFE1HXGrszJyXi
HgznL1eYMo0jLd4nvTFR7/2eDOhl4DXY77SGc8minU0vPwJVwyJ+kE5nYHKO3Nyh
3w4MksJDW3lflxY4BYU5g2NLrZKnS5uITufJ1g3SVcEjdpwkNDRovOvBxRDD2HCC
KvlxoOK8t1JmdQeu5JxMEC0tbVmFg9UzrLMuLtPSsVx8/59OLTAEVwQITeS1HTWp
6BpWoyvMh7x+KuGlj0bdrVrgch3iZthF74S6enrikMWW+J/Y9qMt9DJLV7hNSFhd
NzYRN6/KbUZV+OHsqWy1BMdfrggxmJs9BlINZPzV6H2BxMDiu2wJXfaNl+fq8ahy
ynvC6MG4/APPRjmz9XhbiTf4bOTM/9pao6Q6bKWN6loTuUA6m5e6wypfaLVLZ99H
NaaAZxDBGssHsHgemSmqdCxb0hdLaIvyA4+s8Rp4NDs+NDwpktxl2fsoPUAy0bEa
03ga8Tb1CSlXBadUf5o3vluScHVVoUF7W3sCUO2hdmtlS+wkxaXvtoqu5abp0u37
5DhYXlh0TdSKpzs2b48r3XfnGxq5fOlUN1FTsT0H8oBVkPIHSsSTk0Qr3XYxFM+A
gwtLYl+e3k01XWUlxw0amO900owNAdm5KjGxqECewNjmm2vErTB5IH73rvb5aHUo
uBhxBtZW1qHGfsecebCGK0/jeJDHTjg91RfVNIO1Rs43tpoj6rhxNDMUxummGgqy
It6GUN5NBzvsedoWzvTSpNFcZC2iFH0bUKX02THvyjcxIdI8t2YwWszWxFEZXbGi
tphp7YwdZ4CN+d3Gofkd2kzkV9YB/Bk56hFiAfpMANnC6GX9gd8HulO6xBA/rS6Z
tc59B0cSKfWMkOIIopUeSKOdn8OJWjjbXikFxwKX7KvcIJY//wz6RmRjmYdwhyEi
Hw1IRMoLh0hF3/k7LbPvNBO4NwcrQpe06kA9WWAb41O7aoAjJSyc6Y4GUvfoxgse
RYxwDIAkl7dccY0pYVQWCXH0dd+3jslkl3MhBJQca6HMldSwHsGIpsZxRr9hIGzQ
GvgWGn5e7bMr0OHn+kS9BIDDKhfft2mUkIgnwPgmY0lL9WEYYz99wah4k9NTg938
sMY6XQiIxG15DF2LMixhPygyy3Y0Fsv+xW0KNtxn3dRdACcd1/BQNnYb0KnPNHLz
uO1ftgwHietbDim30kYQ/SXj4Mmqb/PlJfojPddp4Sgjz601lBwerXa8DXWhUGBj
Hib6Fv7BCPWWE5chbtA7K4evartZogeEPBHBejsXC1xdZSYvYoo6vdv5zfbJiQi7
Ss9iTgAz7+4wF00V3snoBuSNjDzQ3DR/dFSwNhRzdvsHsgqYKXjTklU/9KqcN0C1
ouYSaBq0t/DnD/9WajShwdoEu1NN2MvVZjXqFh1mnf12OIGpOl94khniwtWgqq43
9b6LCeF0R5aUIvnMXeR8sQK3wlAoX4MkR9IrBBwiN+wAaCMYQIhX3SS9rs3uJwKd
Kx6K22Z/SDPSde6RLWqCuS0eUVJDzKzymiDg6iOM6h13iDsSWZK69FGFYzzw0JWl
F4MYh9NXC7yiNgin9Cieb0pG0V5A5OcRgKIwFkhwlN0tKpQjxG7GSihDB6FibqB9
pNgRR3o8jUW4txfOsw7JGXeEmcADrB4z8NbioewVCScWdQaOioYR6YQZJYwCj8nw
Ok5+1EfbouIqSk4S8h4o/bK/C7kDf6fBYAtTJB35oBiMj0AmsCNoRhmM4EA14ytA
k8vwu/BmEAUtMNvsxFziJO7T3Y+t8b3AfiNsoP0pVQVQhgLJkfrRPNwvGqoXpHSq
NNfw7l+ZT5S9R8HkssJgWgPHaJNPsgQR9um3li5uk5YK4O1xZMc4eJyxwNuCMV57
sky7NbvGacmqkc+6IwOWeKPbDb+Euo/qIgReh0+TIaO/E2vhYlScDV03iH5UQENH
MhF2VFPpYpBz821LhW/pU0KzI+2HtuGUVh8qefaP5kBbK2jFgHRVS0TdrEOlJs39
cdShkizBmOCsZWJvMIkwdKpdgNLJEVLQkDunHPzJ7BIAuGrbgdnKnHX+eCHxTTO+
Qy6bzmIXX5ak/dtfpCFswCY7EHbW8Q49OsMpx6+0b6B1Xkr1M8tay1+Za49k4u6T
ScMfYwDPob0oQoLg2gC0A3M2qBClf8QKPwMxh0e7V/Qsf5EQxGlbKDcHwT3GbS9x
I8pdT0091ZyvG73r/FNDooXiafWYLClUd94xeRaAznbmvST3H0SOL0tMqAb7bo4e
vJhYYzTMQOVSUoq+nurTVVYY8461Dw/b1rRQjv9gxOe9CARMJmDkuVKOzD3TKpvu
TB2abFDBhEknfemwPGZX8KqO9K3WU+/VYchn5n/p9/f118cYnh/VHUHH6DxvpLe8
J60eR1sX933YNr9itknDiFEB+emOfNHT3xyLm4KJDFIDS6uHazm97ZZLzlg6sEfb
+lTlBSjPXw4k3lEvFq8MMnPb/HL3HulIGJeT5VwNzm9cn4HiumTLSLHKbrjwS3ej
hIIWj0uE40vWCD5atgTX1XAffD7hWJ+5mMFEHy0NtoUfmzzRK8CivO+DrKNKsa8s
enpdnZd19oa5Mx9XZghJCiWO4+w8y1fmL5S/QDxaOykdZ9twJ1Qta/o0yjeVY3Yy
mPy0wjz33iHM4z2TLFnK4OBI4uM6lr+1C7UwkRnb7SvPS3yTMAQ1O7OjjuDPW5Km
zCIcOU8ywEs4vvVDmoyBEh/EgMhNpX6lac5GBAuPjT1suCSPGvw4JpMg/1pWNzGu
mCaCMDEI9UVTloljj8XLeqXd1HCZLfDJFcCPjGaRplv948Id9tzLg5ecg1jD59SS
2uaYe8IeV69ZGjaoeVaLf14tNIrMJ8crahP5pfAXWVldzVdXg8DorxOKNZoAYT4v
yCc700hJ4XlMe5vEUF8HxGxTQRY89GBuV4RUkCfzF1PLH2q1yT57rGvVighulzFc
fIxHwoMOgMg5CGrAZY/tHDigI2cZ1H+KeJ6SF9LY8rWiCpjIf6eqUgrY2DhHfVs5
9vnGoPeYIxa7EzOFmiBOVT4L/29T/Qj3F/VoiPcTyLAnt8Kv0cj9ZK2yPjFmrdVr
N/jYis8PYqEgFD0vXT6j511C9hJZnYGEKAbA0hhl+ggK2dWwht55Zn5X7o+KLzyo
MB7QqbiaLeb9UxyG9WWAYZAdLh1s4rrp+oOFqkGv419sTUPGivF1Iqy3fTr/+bmS
sVheUccuxx5xpO4lnf8/+tq7kVPUoGrstaIQnXli85/7sFkuyiZUrdbNN2Xag9yc
TBMXpniQQujfJt/b6nIeIHEGkO6cOcRNClTNSfZEPBiRyhXIylQLqK83snfkCLHL
QpXESICGcekdnCHuY6HRaUZEieexm9+GPDrO/LYGyM2EaXs7j1aVCCCHFjrCfADz
yzzPHziyVz1BV8buUTdycvDkWGsZJde6uBfnpJRQ3mIhU9IB6d2FQu6pIyxPr1i1
fiyJdKek0X6GC20AjUzNnfuP4DUWs8E/UuGZYJA844DqCamrCnomRQQq2wrPKhm9
CitsmuMOaLY/rIxw/wDdWCMgarp+ZW81+LMfGem5936L4ZNE2Pa3c4+xyYaN+vRs
1S+UoeEZ8JQKmTxWmkSxUVKQvPKtcFR4kfFmZxsbJ/QCG2vxsKJwwpeAaELGJbmq
z1RPWNYET5UwiL4RiJbu1wj83MXHVAambTEtBIVntaD5zrx/HOOX6lK6rfywGixQ
iKRYdRKAEVyo6UX4cAAfFTJHczYVfghpiU45+MTyo81PN5AcMLBpu8xaPL73x8/5
l9Ue90p3iP8zRn+8IbGHku2wDpuOVoQs5iKusyJHbhMzYK9ZeA4wGt4Z2Ajx6ad6
atSyu1Tzup8GSwJ+JYI2q+6P/K4Q2e2AUDzPkIgWVfvTWhdN7p777jW6BtVZIk/t
IQ4KThYVa6gbDnPdUSp1uyLZl5dLh2+pt15EU5ztFDNGvEubG8R7pYoxDR59iSzp
4C1xkwaIntucSxh8KRtPug46zzsZE3drSFjPp+LDnWiOiUFRZPbB4BTGm8Yc8Hmu
S+BneXjzkZYL3V8JY+Q3unzlZ/gB2IepfcG6H6ufl0J2PGIdga//7JB+yXn3pLIH
UEoV/6ufoKXkqxLZXCj4RZ6OmAKhp4p6tiEF/d54l85kll8oc9dGQzdI3HLQQ/N7
GsTeMBLUW2We+sj9jL4N2Rc+DXSR4ArFtLTNbCnf131EQPTxMxE+0genCMboo0um
GgmwswUWJo/iPRhwiXFtlK4VVin2et8W6vsvVZ63Fox23ZB4/+oPyb2J71pzlwnC
1b1ANb8V75bgaiDOJEsVX7WWcQcYerslLUqGJNvYPBKMzyyuEIusTzygga4zGpis
cDaKmkxIUzGOyMetxd1BEXl2dGTQcSYzoZ3ePqTuU5KBx6flRuERuvwXdXHzCjdO
YS8zmk8KuUMzoCWtEB83NLbngNx1sRpu8/F9bgxaLlxf0tMKffvsLHgCNtyMyidG
pbUrWtq5Qu8xw2/rx/q9DK2Z5Hgf1OwLL8tVIK0JM9BIMpar9SFg3rjcSPkHqJKO
7m1kYMOzmmrrwWx2EShO69FLkSt4WigeDyD+IU9/otA8zNcYbzwJ8a9DXd4SH+5D
3W0sH4sDtMk8YXvnoC/QytxXeuLX4r8Re8nJFpbHyuyrlGiuvwy/oyWEJjNFEaIE
mh3Tus72fHP2BPS+8bUADsnyFgO3/46u4RDDSYI86q40/ZuOlDyFFHcNTakkJV4F
Q/scmNHj4EZZ9IeV3+oq5KBOouzHlsQtB/ZzKod+ktWhEaFmJUPvI3c8ZRX0PniC
KGdnyLNt4lTPDKqdww36lFWE4fKPwmpIT826JSvZb+4pblcKGfp4mhe6r0ZugJMV
V12CM2urE0L2QNMdAjN4awSjAVBT7FdNjqtFqDD15aI7toXVv80Rdyo79yCMPgaY
BgKTezkGSNcgucRbevsXzhKOBnKuCafTGo8+2Eae2KsX62UmP/U0is78PrykWHhQ
ua8VDyVyS2+DFzSRpy9MUwjjbGskPKqN6iq455/kLTh657OhE2FOGP3vLkn0fRig
sQ0rzzzjufryIm6MepqPqz7+ZBHXWV1K6OtYwIBv3r3O9BOljc1EZt6HwrKvVDJr
zc96JlgM06TikINjlVsF2TLqxtOKFJqzv29AdF3SqEyt8kxlIyZKVtqZOepBjRvZ
y+oI4bA11+MRcpmBxRVQ3NyQD1r7GTvNwfchmTdZv968A0n85m7JsFNudFgVQmMI
pBuoaKgtKXLLEi4MWq/GqCMKvkqZXP0Hp5lz+5IH6iHIbAozXVfAcf2ATsi/r6DU
9+C+h5OKtzYfMe+HWc+B/V5hWsvTUKXop9+bjWLTl0kMgN42/HATZXbr+WmYX+Hq
r2p8d74T55ucGddXMBEph+owkHX1h8I9J3MLiqZNVOF6qv7XN9A7uLd3aR8Gm6NL
rcw2cQj6MNCUuAOL7ZKX4zECtIH5paASm0mZgnVGhQBzlqAyRnOINdNScIqCiUnE
szEzqpyfydcbE/iQPbSWuF5EZAfIb79n9gT2MjVPmNWLgNU4fAWMS2Efpy3wQLuD
rh2UXAubg4uN9dFzwI2Yg7S98jykyb5mxErv7adZQSx008wikJ1j4ggrR76AcLVk
ZIjacWekY3BjKZcFzbcMqF3g/pAt1WxKpFipj4FDVCVNqlLFDYlhOf0Cy9XseRFP
RkdL1K6ufSr7EZo3h0Eonij59IRodosLMgUItGKx3epc2D+b+ztZCVhdg9qBnc/0
FnYDIpaXRzVS4b1964ZB6uVz+3j6eNnLAbIyD7eEzOU5YVXz7oo07Ef9CeeZhOs9
F1qbw1bEZaytCS/ly0zKe30eg/FJ7725vVDpPbdhwmToAApBhoVAXWPqKqypNyXP
qXkogsMpzlxYP9KyYGcwfS1INQ1gucV5f2cf28QDOjy7o/mNTajI7clYywW7Zu9i
UFwmJ5yIUWnYOOg0wwLVwjd09fmMjq8yXXbHp992+dOr5giOUiUEpqCvvu0TKHBx
dUhq1OEe5Xjs9Rnbm31PTAi6H0q50lyzWyocT8SSDV4YWYlGpUsAEDObqV/4/+dz
aeCuA7efsoopgfFj4iAFdgvRt/Zdtp3XC4QIPX6hgvP025iZVUGaYTJUYlW0dT5Q
yr/ubzli30Kr0+XcRkvu3XQpEZ/XJAxliPDcHAMzDFPXaWi3gD4GO2fxy6WWinOn
n9+JR3axLxnYIP6VzFQENYRW37tpzXbK/qsmMjPEOjmwq3741CIr4AC/vDLxNWf6
MSrVR0AWGl0B9txmoRo+dtkWVouYlHRP+Ecj2NG7atgMfQWjiEpnhPYElqltubvo
oX57ydAERf6JJjnh2pJEkb0hOaAgvc+ZV/Sv15pGT19XA67dmm4sgaDnwk1rKoL2
GDQwV9tgDEU/uC9PxpPBg+PT/ZH3FGaHNOP4kIYCOrxaGzfOWQtlqdc6dWc49TVG
PMwzls+x7S0JC7SIyXROEzv/KONptn6pJnEIyNijsV3aqp9g7A04rwi3R6C/DTk7
mup3VkzvxZApLZXx7PUIaVOQuXIUQJWttIp4hlQw75o+B2KnUKZ4Z6/q6jRrBgfu
9PeHNbIIX0OG6cBZ1Z3XnS9zTl+UleymEBSncbkMsgt0BAdaG45ZycuXHtHU1xyD
U3Qotq4cXgYDAbfngE+tLNnNVP0mcf2l5dbo1Cl1bwAupaxdJA3f0NzR/oGnndLM
M64dhaDoRrfOO3njYMCOS1OCVNvzut339l7wi2IrC6or0QJx4ypwbRSc9ZY8EJix
A1mF6mdsnky0+5sTb+9Z8y3iKMIN4nWycJVEpro5vwZ5HjSE3nrFWAmqW3Falq7+
mZWvQDvSbn2KvAAHf1Dtto4xGxsVMthXj/itsNWYaSdvvQY1DWEGg9H/jWU2K6FA
yfulqLvqBJrAvSZ/ftaU75Z1iOuxaBk9wbPySy7ihFhHmAVXR7zie5xQTxJMefpp
7r6f2+KTi1XOg3O+gSZAV4QCp6rWTNdYrc+Wl3wbBLluqjAMYkz+b2d5dfyrtBT6
VedPaYVCgsqf+Zh3naeU83sfMQKNBZwR/ySW1mLdpHBbxUjJR3A4exiTE41Zqcxm
mL5l/37VEBLpEKHkv33nMxdMCT6R2d1PAkmT965kg8N01x/NHY1jnR4mJ3eap018
krZ1Lk8jlEWl5JddwahtEmxGTLsCvd6ZKA0JHbRYC69+EOMN4zV1RovGYKLdAaQa
MV0FvVZ1mlAFrukr1Stq6jGxKCMgjmd8aNWjaW6g8wkfK4E77gqMpOgJS+EZ15AG
D2CAbelZVRYsaD2xi7QQmEkA+eRP56UotfCc9C92hJlHj2MaOCnSHOSE0xleyydv
7PPkvLTtMurNeuwh76bwOHWJusu3vpeaLNafVbcoVkZN5bhAGDMVgJVBI943A7pd
i/grIB2YqM2vvCFuAwpVHKdkzkWNLPw6rskfMwDnG2C6QZgZrMDQ84W7YMg4AyIa
Ig3lMElfvpSFRXdLBw7wYqWqf5zdSyG6gkigLQ8kzQwoEs1TB11MFVZHVcHOCwc9
5qCM+tHa5ceBxm7LMZGWLD5Xnr7EaQovvzYNuuMOLeOT99AV+C91fGH7t/yA0aM2
k1TWhh5KMZtd5aDDDOw6juif/6dThdkaB7sm7St5uS/eCHE0MIwFLsO1poXZ9ebw
LXiwngsgSYrYqRxPdTBzoj7M0e6fIKC/lVze5ZHJFmB3eDNBRtZs46Hm5i0OCwbg
duO3+rlbiKDCsx84guTjZ3Sq9C7BMzZh/GAOdOmfxns05HjXF4u9+ygNu++zndyO
JN7ydFWtPNtDrk42KegD+ry1y+BxKkRASrsvPalWQILbG4TrjhUihvsTvgYSttXy
KIhT3HywtrGXtCJ/F721drUiP+qjJoh0y8aB+GqxnaU7BHhDC/tehmAgy0/WhpWC
afsHPYdD42GLnX7lUxThAa6OqPUU5XkfcCRCnm1aiYXZ3n/1FmE6vExH8dNwjP0V
GP3iWVdOLuEe1zq/XWiGInWO2QDfFr1ilpFNrM5VAH8JMl92at7UPF2LuexQInWo
dAtzdl+iI8qRHb4y1hdy9Ze14nx3bl80ir3a8OorTUwJoaF46+l9ExnoZXPLTe0H
NRE875K/TH7MMjO6bpDQXQ3ozxwzgQemSlsk9xbS7LwTDxjExwc5Eioolyr7zbYQ
d+UcvylYuFapvTzYdK7MqRaxEa9ZM/RqeDX5hXe1PK12dCfK2XOYYCIBGBL/B1D+
UT25DMt9Sz3fplB0HMDw33N9wXfvpsxj43XXp5svEFd32aE+VNHT8/dOrfo9pIGU
4t6iEFOnBO1vaLLe+HDdG8BXHDCEOgPRTk1OfAlNHBX8vjfAYP5lN43ZvrsGuqpo
bZusCaPLVgd4Bpi479SuAz1mT4VvmGsEOLZXI3kH3xh/drSzAaS2HHM6GsSqHaJa
tHzNkPbQ/kWXJ0NJLFBgtFFU69/Y3bEYAOs2W2aePYbkf+DzePGSSPBqwoSdif7u
ZvO1qujTDuASX8mUPDLbtiNH3UJumISZyj4yAt0oTsj2YsS5tFvYqSKDmT2PTamT
4Jmn6OHqbEUMSVmYWKYT4RisgGlW+yYWC9mpqg/79UFgsVde0G/PK/zCuBj60ajC
BAaYmL1dhhVhEZl9Y/kZ8Se1Rq/Jrhvrgi25NBFPn4LyH3kZIVZpianSv1GUeIZe
F7xqim6bLrzl+qCQ7AovBbfOLAnxLOzcNQpHYFs9tlgfyq93lhd8nlLjGvn8Rz7x
kuWhVNkrmzicznyaOCIJYY6lOUxRJ73c0D+ZvuMIh0YKaSE0sRqNxC8L7pe1Hn1O
wXoqR7Ogpb+IdS/RD61ejvIInzKj8dmNDAvAp2+BYVRJz/HXb/chxnoe5L/hS6jW
kDPRvRWD1yDyysBQDdKJEc+/Xs+YDipKyX6J9D3PGjMQ7eYqmu9u9ecExdBA6u1V
RCdOh3DzzeiWrFHkEAmkdcPy29q3dRz+w3DglaS+TCRKvjZH27bFFmZXA9Kp2v68
qZ984R0l8xw6n9GNhaYUDvMwRWpyBflQy1/7j7omoMYP3+urgOpslKpROOhxnfS2
QdvULXD4IAuZMI3YnqQEgzWHWqipOekqy18pmTVezEenrdRBjIda7CdrGb3GGYEJ
3Gf2O8sczWPWeOxFrTClQtYqw+WrwOC/fCWaS9lCMx46z7lr+453dvtJjG+jiCAJ
jcmLSWBfhSCdb68Ot9tnuvP4CGNq35ebb3o2BZ/+EmBISAoO+wtBYCMIB33eQTIb
qYElJBGHI7LeyJMFXGXGrVrl4bcAi8Y2SH9Bx3EPKFfH+7in0WU5djqzRNRAHpj7
+SQeszP9ySwL4VrAQsV8gQf+jgUrea6eIRGKRZdY1jA6d2F7JkdlIsjJhHXQoaN9
/iz0qN9TpxjW9A4CD28qps1pu37wWyv0Z9kjoZFStPSv0XfSDWOALctMjKyXPM6I
yhJEbsCoMHx/lCUF6IX4WzQYbtYiAGBZMRDeyEpEJkc2W/goo7rh4+wXTdRzx0lV
TbwPgftZ6+TIS7nCrL3kHP2JhMGQJx8buAlykV/J9GbkzMBmnmA/uMxudsBeyKWW
/7m94f5XQXg3Qb5gmGstPeRNHXuB73I96YgLC0n8l/sW5MbvWycnugElbJIK9/AG
rGRb++e1Q5HgZ+h8aJSk9xMfQ+AW9cLZ0qk8YXwTguEf/bcoPraNYolNPpdjH+cE
gP8lXe8yKVbZThkVm9GyKA2R+mZzaJc5yAvMwZIUUWO0DXsZVCSuxqX3pvwEiYVG
+TxgtYxVB3s3nDmnEz0FIF73pC+ao7nyNBF/Gd5Nk62+dA7YeamMzMA5x6a/Tl2/
/8RS1kxCwplWUzzx/AezyKIsEmDcpUDJd2I3OyQyvZd0SI/+SNvwzM4VLg24Yog5
OTvs2XqYSsp2YCcUmotMQCOoU+yrTCnJkEbhkZZt9eE7E+ZhFeO5/STlArPUm50R
ro+k3IvpOTmRexQbddj+Fepok2F6IurB57jMLA6TaqIbCoJoCEhMPKI9Pe7CdE3f
hhBsV/V9KplO/YjO6//Z/18bwW8Qg2t2qjYQ+PCfrdpcWgQ9sCBG0oOxyNPCZxmC
Nq8wotqYJdMllX1TaYJgByPrKlUFnBqVYY2nJB7u0lT2zkVqqrDKsJg4XuuJBBs8
WcV3WCq8aD+SRm2ZUszX5RSFbzSZZAf2VEsdOxC5BanwBE7u1zWV4bIGDqL6i+W+
xFzjq+/DWDPyG/vkQrdvVqofQSN3DUmzAO+izKjuJ/yHeS6Eq2wMDs3UgRokvQrb
LDnLWHSOyh8PQwrrDwXSTrdGzTaBp+4/Af7e8G/rLFKG5/S6ptOR/2LS5ahKBfta
ovfnAFzVuGvQ1Yg2I6+kRcVr26H8ig4kENYMqRG/oWWiw4FgVE8lV/38K2WtiQ8Y
QftUc8nNRIYBDEUdvRhuU2xPeY4EUK8yMTgDk43z2W5oULG9sUOzoLdi7dHkZ6Vf
fvBOLEO21JsCnHQ7RHNRz456d88z4MTpm1K1Ll5qaBlcYLuAg58f9Vk8Yn3g/h0X
+VYLyysJgq3x7eeZ2gcc+qGvHojm1fkNTKN4dVGP+rPCLx0ZdT5P3o9iiJQq5tXX
jlcmq1YkSXH/nXmBofk72jsozWH0O7pzi6Er+GQ1gaYDbj16H0q9Wowgcdr41JXE
MdtQ+FPCdO00idq+ieXOvLfnU/zdGNo2nx0R6Oup3f34NqVxI9C59JOFJNCgDjX8
tAV7puzhAZCj91tPDWhY6CvwNtCdrqXQdoQ2AX+D6H0TSNFNM9IbI2qjMg0d+FFS
EeZBjMqUcVYvifJUJAUgIhgA9yH+USuaXoVEQHt0MMTSF0EkcH6Rn1DqpVNgmakR
4q/RxTeDIUkQ+Yp1wh1IkL1QJ+ZtBf4PFJZO90TQmquSXiPwNiK4LMVFqyRrfLoD
TlwlunCrZ+R3RS5Ql0i9o3OPjxL6IySU4ORG++QMqEtSiwngm+3UaqtNDGh9jrBo
IYd98gD2R8imXyw+VnjNvrVrmZOygjMYboePwvrMMJmq6j2siKdJAGTaPka13SFW
gMEk/R8dd5BPpDppfgCQVbcX+sy4gMPle1svs2CQvZo0hiGIrN7+5SLlPW5mZSK8
4L25ofD7sC6Mxxqaunlh+PuvfJOrEA1+d/qz9btLEcdlXbqyXtvPbe/WK+29Awoy
udQo5X+c7BY0Uy9lA/2bgEC1cBZ/xc12Pmy7H6ia6M7sPgajiN1uc4kqPAK6IBxl
LQt2bz9uFi5THXporTvMLieAAizE0RTe3PeR0w4WOf/ictXrXlASVh6Pb0ISWIoa
yEfiAROY7O7Ga62/EFl7aNggR9F8gtRWgyVweOJwK2cPz2BOcRkRrQ8edY/Z3zEw
fbCT7R3VeQUl7QVD0etCwFXUoi+k9bWsfBfVnjjBeOaH7OGzEYqqMpphMpPWbaLe
3ZM7VvvOAxW6gDZQatcHHHIPdihLm6csNz6IdOmGuwDhW6FTlchIciqrUtZzLWXc
7U2fpODv75kVrZUsSjtoNYLZsxNeLFVYpv6mLC3GRftkfmY/eDLDsDaPQtMNCykE
61InsozfrXdRVbxR4dkq8PKeYKPxBJlb/4ulFmULeslfPr5uT8z/Dc+r1fRA0P86
B4ObgZxYCiYha2YptOrVWVDbbMc8LB7MCv55ezkwz0CSDXE89sl2aUgMLORI2ms9
MnIwW1uxegvqx4dxUP6sCV/fg+KqROyUMW5L3rY6UNCMSzrE/NO+VcAUtyesDVKA
AQ8VM4cxvV0tDwl9CZdMtSFMx8M2cftodW9hRnxU6adpK6qlnWksPsHMZ8WZDbc5
m9l0SWWuZHn7m89Vj4cB9GBtfFMNgvIOcdUXNNhzmStayB8pe9/vA3eP/IdIbgaw
SEZqOEhWinsHIB7b7HI1afZErp1ZCbOz/Cgq2EF75DKjLQkrtZ+J/WmLyEOLe2vz
1nvJu3HQrIUVmhOwCU+/GgGShPi48rs0T1aCbbRdQtA78dPBAF45fKvcHeKYcAbc
cSsG4YoPwGNCEE+a/COCAbzIopOGaA9JLULz+tSis0t8cV1STFYL01K/z9dj9vBP
sKdn8QSKexsvmQRO1U9QPk1Y51Wxnq/uwJU0tvsRZ5BNT2lm6mFUVRPoq3jqdKJd
qdbopyhhF0x9HRxjQcOKeW7YBX7ghrGIRUitx9eQiHDmkOXry/xuVjGBgl3aa9lt
acWlQ2TtPBK43ikIX87zNSKLO00jyxm3e1aMZ/TwSk/PTN6ygVs1GbrSg3B1odny
C904LG5BIT4WwVdQvTt7WnxcbzC9f8QSMl23WUa2WvfnuoobSvWPheKkUbtEN5MY
WpNv1bIkMjoVcg+k+DZqpkAeHmV43zU7XZqx+HnmUQtj6P27PqfNUHltmVWiXi21
tLKHo7RUPjeTeP10CL0beQWXQaon128res+bOLxf9wtL+KlexDgAse3S7FygrmJv
5HVAQko/iEEVsFIO2IiqaIjb6myzMTsdvpixltKL1x3LKF/G5tQimXKN8q6/HPYn
TuvcCNqbxY7ooSfXbDwxTAhkf8RO5+RdhuDLxPcGDEClJfBaQ225hrSSwGmdD0SC
xXD/g9w3kU4bFLvzXTepiaIAl6rfwQatX7hIugaYjmHhWR75DARCEWNVSlBgSE4s
tCr4Bkgn53sAnlVswwi7Xboa1xRaHs4WIDwzSHPv3SmCcFfw+DZllGEe+LRLhtfX
U0vim1LrFQ/WHJ8AzhCc2TS0uQT0xvx/c/1dNb5shLLS7RwO6Y9IJVXcoMF5Iw3g
TEf8yqSkjlrR7tHM55ZWX5F77WLjS9/vxUsKbhEWehKVpatklNSlUXcLHYJBwuhy
x1K+T9HR5PyjO8Zkg8S5iknEOgtqX2dAxCWcY834cnDFbWBsdmyicHS3bqrj8BxX
5xFSVentFsOjoDP7ohPt4n/qRiyr5AV7Io9W81uK066oLUkUJ7kqDLvMfxIWq/N2
nc/oVq696ggTpefrhCMeReN29yoLdu+E2Y5D7BtejipzcDSyUXb+PdZYwxvhzTP+
1SnvGTxNuVwtlpMOtGKpVvyCO1ja7TRSZmptYA1fXuIp0TBDZTneW5ngb8PH7xqk
lJ5vYJcB8jsmZrIl3srOQk7mBN3xUzbWXIkmAg3iQWSwIOtKrFDQbfzazG1kvL8p
wHs9Sfr2O8UPmTgopXPztQKfaB/tiEOZ8Koi54v98+7CphlftPHc/dbjo2BO9EG6
F61eWXxAuULLwr0wrr4gIWu7LEfoxeoKIcKMKq6o3j9AmWhFc4iG0C1VQS5l3PZf
ia/2dfH9yh3SC1/+GOPF8lw7sV6QLnh3jgy1ahpRdLv+OWm9vF94IyHNjUJbeHDI
UVj0+FzetTlGsvxZtKrnxyaUKfkZtkhQ3bi65rrTuzXBSUHKKU+wZWxdIPfurSXI
exTsA5ZpdmoOUT6r8whCV9Y4yNXF64zp0jNzXClMLMJCrLPeyRuu6DjFFGwqyDZH
O/zcaDeJYoAP+5c9nhYkezm8URdPaLPoijKAr5In4WanmsZNDCz2InHV+340rl1E
bSDttOkuZTLgYJRSz4lTn31ZtBzORGExYCJa05VyNFAwDf6uFIhhuMUeXLxfabOh
cVrSemAEgOtJ4yO5ocSxmN4dSeVzDpnJaoZQz5M2A+dZLMGgMorPyek0Qt0GvJJZ
ayf73qOd2+6yshEVOVIFADJ3aI9VAL3vAIYJ+ZoyDY1JvUWvrPUUgh5tvDOmhTQ5
f09e89v9bzYb3qWjcC+Q3tl1dueh0VsHTKWZB9P4ycIgLnWGZEGE1IM9jpv2VGQ4
TRI+IX0bv5G+iRG09N+fEipZVdFvqdVQNgbhCsiMMdYeV7Gjvxvr77VHl/BrYSPV
XYMnKErgq49GOXCPR2KlpzEoU3tANS0SfTsdaUFyHG0FUwD2muAUq249WldnIu5T
1mDI1KBNeuGlbmwuUEBAAyG9WWcyK8c9p9hg+SixiuxzYeiDzL1tofw+lkQQXHba
bRlc7ZIDcVxMBkAnRR3yLEv+fBNyuKnlc8Xz//My0BNqiCZ5QWBgDGKm53cRt9Kh
z0MnvYYBNtb4m/nksRkXZzzgpDbq9zTYIqjNlUQU/T3hBzckCU04XOu8+p2VJLiE
CzFdEwiSX/iMXIE9x6XVat/4kVTMS/XffVQHtc4hAdhV+v7v/ULcC4i5Bvh5k6Ho
cPLZdivwEKA7a3qdBBf48DzvztR6RLtK+2qVbNk/vx181xCyjVFNmEELVlgvFGLs
I6DAKZwuGeIAuQlY+5HGpQCJV5D/TU+MK2c/HPFgNPreFbrX5pAWpt9AExoAP6rO
Lvm2Z3/CRUyVdshw77BFmCRgkKbgeDYupgIcvk2q1h1Pj5z+j2mTzdyKaZoNYoSr
l5t68Sw6h2umrQlU/b4nwcpwxFRa1vaLpHcQDMywQwP4RYBrXXqof9D77gQ/kgjA
1GAqDqqF4X8d2r8Xb26gN6dave6fBpmVkopElsnUNDokw/Jgg7cgj8ZOUeYWf9JK
HQFNdS40zEf1X/06Y/psRfNWh4he9L0yOV9+DDxY0KdBrM7q5VUIvbLY2GoLwR+e
vf+pHclVlo64r95TI26ms5eFye12X1etaZM2YwmJHu3clPLmdpVWRM104f5Z8G/A
zD9w5SEs1RvtyRngAL5e0Pk2yVNOv9amv5C8b2m1uBnysp01b5b6UD6CFTvqI7nK
CYUzvda8yXgHAqi0tuq7miKVuf0eXfO0Nbgybzw9LwctZdUxfwMwpGK9KOe3KU1J
BmtRTsc1yxAJYNtk6y1laP5BKk6Khb+7CVgaVDY3nQzernytze1ieqDx/WHl/X8v
qPR7NOOsOUfREGex8blAsFV2/iueUgHQRl56BOqgDCgsRkiTc0QYU5TkwtBfqtON
h4ViXgLaYAdDf0xfICRVzZAxHmZ6Bh9SghHJZ5fw4Z3x4L2pfZgYx2vVG9u9Ny+h
+r8/XkWaNMV27cveuf8Fzpkq+HfN4TNwZtxxFfpBrzCbmSMHJCQAoxFrKiFxyCyq
avjtiBkLxIcVF04hpeXB+CSkCuSTVXxCQUoIKl/ph3snrlMeAZpA3mRnSphWYVn4
q73ryalPdJjRLErtv/PVn66vjtMBQHMu3KwNe1Zmk2wvKnsWNaRd7tYYA+w5sCE2
OvT/lvhwZk0+91zcSS4iGakRPrbdgYwCBcOfc/bbuLJSofjiBe6wkZm+ovHWqqyP
gDUudtFyMS4MxVnC5moxGxbEPAvwhS8j68QhFvho9pyeAu0CwcmLbdl4Xqkd9q3e
3X+SNqfavd6stjaB0ggr5HoG0LYHZXgy/ll/hx9VlZrbqAr15NphfAOEA3Y8D59g
5RsrB6usikDOLXyNkovpaBTKvAhm1ZbAzAQUHUmMt8hlrF6UWnVB/Y8KqRoSYwTO
FQsfEzzAc+LAjczP6lnVdq2ryQIBqpb/BpbyNcNEsGj9qPMX9zsDBF5DLmMchO7s
WOVyng9JmrWduU+geFjLh22a+Xc2MGovbF7jUps7u2MNm1Heh3vwk2ItjSRGHfgz
wW8sCgn9qAmaDAtaEz+iVa9OUElRa4+rGuZYCRN9u1+zCGvu3yyjqGwv04NOQGel
Jmc2E5XFIrxUa47Pxpm8rqGu23saQgHtY5vB3s2mxOepFh+GcGzPUj7sueS/eYcD
ys4SoaQ8GRDDcTMZCh6GXMAThcTUw7z0QKHdVCLjAWFYXekpSBKarmUQNYzfkvXc
j26DMubZV6nyFG5vAim4aKw2HqMDvlY7RrwhTdjVQHQ77+tShMrRzmAvnIsFBHwg
2YsY1H4oJMxWfDPJoaWi04iuknmWaiIPFZIrfeWoY8poldYOjqdvwlmNUDQSM2nn
ico1D3c8SF2A2Ac9DyKDuAlQ4O4DmETO+Rrq3hgJfheTIAOuWaZ9YGKZolMrk72C
pRGKzo8MjT3Zk5lG3BhcagKtYJn3RToQrhsQSEJGhSEstMP34fil59VCO0dHxRfR
h/ra3UmzDfiveRf92X5PpWTwSBja5M3E/Q07/PYOCEhpR51h8TLJnacS7EDW8cMy
etTpufxVFBWhpfiHyfcmMOK2gohRJd60snPRO/u+Se2FdVc2+j5ztT69UI9fbgWI
mzWrKJljlz8QyCF4jlAiDdLNse/V1UKo8pWPAiF5aPv1CPJlLNt33UVQVm3uaE4d
JSjTrlHm3henQUvIqY8oT1lUwQwCUARukZj3Q0JFHY8yhpieWbBxZLLiYRuTSbqm
gZ6Kt1KsLb+EZUh7R7KdLTFIK52cDx1BuGV+zEiAyTLBe2EQbCWG5RiO2tRlRhx0
mqhH5D0LjmZ4H5OgwPYmGyzvnD5FdfybH5fcZIf8BBqupxlFBueyIpcQjezG0x1S
uSXAQagYUOGjE75XiHgLgJM6G1ngtp/EmTNIVoWLHukp1tsg1u/U7FJJ0j77ER0R
oGy4jEYrMNLjFTURN/C51jMxmdg+5zHWrObPitpqMMze142sdeKGfJvjSX3vEVh6
ChLi896n/UiKm/wS10IKSXRAWt+NF00TVtow7ABEW1e8fCgltTtV7ISuQE5cSipo
hbBIOkzQwTD9Mz0j1rSOvzJZhV7Rn1INLMtLQMx0Rhyh0LSref4COYfF3IJOL/YC
eojxjZ4bJZgawDgAyIEKo5hGYbDuUiSWs8C4b9oigA+Q9ej62pRPPg5NUruEnGdq
B57JD+ykJZ3ts4sH8ftBEGpiEntGnO6fpK+BDtOeHe3pSKIGFk3FyL5napg3bmNC
+OsApQ6+6iCiYHynWVdvYy/rHFlMTrizf2aPgFeoSH1Dmv+jO1ZhcnQc0cnWbAXi
rRqpeT/5Y9WURlqOuNmXVLrIUrvfV71XnO6Mgmff/mDOtlJjfEUf/Kpcxy4C6E6V
ags+ntNdNL0oimvCgWxhytD3tQFQH6kjt+5eSMT+N2nALhr9HFc7yc/+u0bu4YFA
oidjuyOo+tpWRtAggAbJsHNzsGGr+dmZuuNHZUekhGk4v5wzZfZE4IXe2NeBIdQT
EizRazkvjpDrKnRBMiTEdqn/sVvdYM5CV/yaRQ51g9mYnDzi5YCZmO3bwKsAN9zY
JTdqdn5eHQDm4SgB1Ja1wb/S2sSavCTYKfmJLcKCtmqsI5N5GNELwyiHxJVvAZof
nOB0c7cVCs9Wp9PQQgOYDIsCvi1PtEdh4i5PDhcJC5NXouCiTtE0PWnsbmzhyj/x
o62ZqOWJbbXf7e0J3N+s83UJTY/t8xwG+KFOgHXcRQ7K6jH+P+2qsADR2T5OPQi9
39Xh3VaHlFzomIUH0YRjssHiFC6wlVCNCRMEJmQTxdV3RxQ+1DnQ8F3TM628+TUj
/DTn7JAHoj4DVr0PC7AbwAG5hNkqGqhQgzmG5E+WxHKhXN39k8fRzqzhuo3YpVXc
hXsOKFNl+3N3hoQs80ujDSUuwguLZhyi2+4uIqnEvsEglfO46zWsXWhxiBIObR5d
4EI1Av8Qhs30v8aFtUh5zYnhf/KSEC9EOWDmfR8XhBbzSOfFP4v9OeF1KTp0bhjj
TNYS9715p3ibejRR+jUd7A6mT75ZSuGBmQ+0Jn0JTJHTGaE25vEH/iGdhgeNpDyi
uBvDcbeYQg918juI0VJIUDcI+OCLUIJYzL+gmZRDOtX20X55O+r+8hAM44Zrs1o7
JkOkHp+kgGp7gVV/4MKW9cwT1lX6+gY5YumbSb3xI7JJjklkDb9jqQU0j6TasK5x
SDNlmZ0SXABAd69z5DzZtYVvk6IwK7zUoXes5uZ8nbQm72BvL3kmb2UB5ATxIk84
GFbziPrmwDFDks4G73+3+WwxHmoVYgpvwt49A8h9Bv2UjQcTadfq/m0MkNnnXn7N
1g2qZUEEvkooJs8yiZQ/qy413HHc41hRCESitX9odsye8bhADApp4+zVCVP8kOKG
f3wR5TIirOCv89GhWAOp42/fsyXqEcMZ0GqJTQY+G2ZNWhminQ9hR0HFcvpLe8nL
DDnfiyr7O4ERbjm/GEPAGaNkehMrBQ3BOvJJjy0OFWpm12LFuYuhO6q3qx5mewVO
W5zlakpimOHVqJR/VkZXqTS2sPReb8h9DtQDw1VPJlOy1r7APMrKUM2aPS68qJ7i
Q5YpP00joUfhgef445Raof0w+4A1+PbnwybukAXxrqHePrvNacgnHGYDVbW2yDBT
+ZK51NTXn12/kxhpuPPNQ0LfFZvE4Ay0w+XeJHFPCP/4BpbJLsdDqj+OaPe0px5G
9akb+GpgYAHJdCvoVOyjoO87c/3334ZuI/nIT5PXwpKcOuuwunEpBZ7u+bMJaHKL
MI0f6rOF5rrmn1E3eXKmGqxiaZrjZk3dQ1hLuDSye+g8oaaa/cgT988tYl6Jr6Zd
DzE5gpRFvn5ZsPoOa5rVbsKNjWRlefbB5gL/iN0DKKB7BT7U+D0XJnsK9KR7JZqG
VEfpUhmhSWzDPeUQJUGdOE3nUw168L+BOEWA4NymObgPiepg9u+ewtStoED66STI
Pc/MVt/+1Y+e4YhMPRklAqfEyBIhGHXZNoco91JdwzA8ZF+WmO+ZQOAyMVj6R54k
jXnK99zJBTU/uxqa9r/lyCmW5fwHW7W3FX24KAKU5X3QmS28/Gm0cNS4lWbOv4S2
UmfwPfksPBdgcsOQ9/7bjsZUjGKcdXmoMLg1Oomvi2zInAMNAdPoP1kEQcmJtw8w
3t+Rv/GqvtfENn3Ir0zOfPwaiSy4JVys9za05c4fkYtQIacz8MTLod9juxgxI6YK
aDpyC1oXY/w8VkBv/GDrfh9XvTX2UuMS59dAPpr/BIZSAEYCdUtsH4yCGzDQtUMK
eXmhM7xiajhPtLOP6tWU9Jl1T/7rT/DUe9w7zK7WACZKTr1KGi5XTKcRkzrwuCaZ
v/yBi4GKbmebCCfM2wC6/BZ6XRfSdSsRCa0pwW83YOPJnfZVz+l+bO7erDZHCnU/
OPfklRG7uNp0A7xH8CZvR3NeOHZSmz6c705rBqX6hJO5RmdlSri2Yc+hC8DsjIIA
nmqYIwRworqOABtj/QmMWAChCcpYyQn9E0hpvWUky3KOlCwzag7wJ3kF8jD7Rnb7
3/y7cvsvMh0cR7y5zt413yibgzMUG1RXvtLYi/U/i1LXSfRMVNb/UExG4OMm0PDK
qxey/+BL9XWLZlT9llV2qY/8wO0HZ68EDqq5JtpR/VSxub3ULlhWDIiDHM3kQa9K
li/0rr3dHkIppEVj1cpwc6xInoX1qBYembWHxs38jmZm/lLaer5Vyk9X0fBwkWV/
5SXcExfh9ZhBPALpU8qlaGB4EIvgp542U+Sf3pyfL9t9VbuFvi0dTTEUby+Cw5ds
gb5Bujz+oyzBtFk7NVzjFW0laG9+4qXDdDH6TFM8uU0IJYwE+shS17Glhww3D8kX
gmTa1BQm5mV6G90TJJ+2V0hkMzsBFIPW8Yrt7GY33qv5xY590/DUYaJLyMNpts8l
JpwDTXpQpeBWyDcSXzLZkQ/osG2ksqpqC+wJUZK5+r+QOQkOqFGepRZ7s32vRno2
Zk/uU3h01UxQt1DwdpTAqpU0chtDWmH1ubkyAi7LReD9oqtKVo8XlTu5b4I7XXpj
0b6zM1fmM4wUCMGk16MbkAt9QYBaCvTKlnHfkmhtTStLlcYzdwiL6EASSLrO/x/4
l4ztJT1LQngjUJBVQ+fBGiTzBK+ZmhY5X9fzBj6TbLLpGnNLXtPiu1EjF48HHHph
bLVBh3Z0URIMJABcNPPbm0o3SqtnyojNC8Fd3JHznvCTm4vuKONXaKnWWzbk0xNi
5YaeIdAOAR3vGhYUTl098L151oyRoDxW+xtS5P1meFiHetFARL8sRjOB4RcwicLa
Q+yZWdYHGIYmZ8XPYXPc+RaFN3kV35qQDuLBh8tDJ8GzYkrlysdOFBQuK9SkKnX6
E7gBeDo0J0lQwTxftHFKVozJ9inBnirhvNycuLaATy0YYJD2CU0G/h5teCvR1/Ok
UZsGPzktRrW45uj5Zz49bDQHlx3APwu1JrOx3yi1Q42m6gFHcS7HB4GlL4+w2Lgm
WeG6freDcEmZxMscHt1PS5ZS8NVUOF5+4ofF5FmI/JTNm7iQqUmc63QMv8I2ExfM
PuQDCAwDwUWpnO77JnJahkh6OSgiXy0UohGeBnGV2nVWJLMSFFBAmSYxN7XjpP9p
WLWW5ilIDlJ4Xopp5ORant67ZdL8bBm4E3Hmo6YsNqGtSsq2fAZBowVENGFANOyz
iJZ9KlPkafh/OkibjZB2dtg6bPGiVax25d3iC+2XiwgC4gBAlThMgYRyMKV0RqMZ
0bCsPB1HfMV/94uxD/66Vdtp/iqMLoCwsMStfnBHLZtW+yRZygwh7mPdbwHDaecR
DM6MfScfTKV2n4bnUrz0jbHvxSre8qyDxSvLo+WW0v+TuwmQlYFPTDOg+s6GvXd1
71RFKNRB9eX2uVAPcV3NAQ+vw8UsAEXlpmBXuoJD+I0Zn6kTzKsusFYYXcxB490c
RDrLYOJYFzjTyFKWWes19k1RTKfbSzugY/4B7vfW6NkiabXWUeqXX0GNYG22cS2w
aJKEz0FVOp7RdSB6p+CX6v1BqcTMXiSsEwpDcPxpec4jLjNI/pKZfwmBbtpnwGCK
h4iZy1ytCGVOFZrthWLfvxt7PBLchU4LXY/2q5VuYY50+HKBpssSVd6G334LYA/Q
666njkjYlO9R3fbHTnxvnq5GbD6NHNN4FRDg1oD0FK7qnavUAqtHH260+dVVXuSh
bA2Gwn4ZnqCEME6PN5Eg0CqcWxkIEGjLi6xpNLxWItMbeCufe4+VmfxwHbzwlXe9
SSvC4yS7xzMkwu8IbzITQTOqJF8kyXqDA+qD9wOf2r4PrxhrC2Syr/KBGbTcEeYR
xhJklrzhla+V97vF2z0j5enk6gzcBnrhpAqIs2QkL3CgFxSX5eHZ0f28xxpB2oRI
izrL+NW6BgMTOjNJ797WdXP9+EovhUI3PsEB37iSkLOc3P6wcNj4vjfGVV2IEIkA
xICJoqiiuRbCFu9+GUaTrO4BxFxn9JfM77zfhn+mMO97KcSCGxlqI77j3yBPQHIm
WbWu/Wk1KPu//3AdHC3I0DY0d4Jes+4Ej0jGJEhtxBNVQZMIltT/gQZiGmGrpndR
UaClBIu6rh2V52RSLVGKcY53yRDRbAESzOTLtdQb1VxafRHUWUjAxUFShmPZIJ7x
yQVcPHfCQUcan2cuRf9/ql5WzN/bPafR/ssw8mIRE4/ir88zjxhiZ/2kzepBpXFC
nTjujrZdzl/37yX+iB6nPnazEC92np/mIeXmk1zcr44d/RL0Xbs8cqHspg62QVPY
GR4lSA7GuhkouYEmbmYEcLW+QQUF6eiQQm6sFKuNHLJ6HcDsv7sQVyOr8xblqwZV
kQzBE82KQlaebI0AroLXfJNAkrLhvqu15JIxp+KPfXTznFxtsOoDsqQeyrALcHnj
X1sWwtENMpA/WXbfkNl0/tjmZDQil2vvn8Zn0nRfFvDZrvWe7p5mk6L++0DK23Xk
oYtFrpb9y739+93XjqQeVvxS+tjlXIdrQIMOUP5HSuqcUDaRCQHDVOAvtJqgNxZ1
wLBomayvDOscGewo/VBoDOxeF1bsRtSSFHE1seCewTWqGBFgojNUAIkgIifCDq67
TH1GenOC8H3KXhh/wDUnVnbl72qRkaRNfzIh3wsMg2XtE2DDuiEO3NFqxmAKS6KB
5GmTB0TZ9VAyVqo7u85bYHjZvthR/8npvG28MvdyNd717FUkDfJgiy/UzuOxyust
eLDCDBrRFPTq4sAx2fsAwFY9ks4Q+Gta1sCTpix9dthD7OmFIHmwDYyhsSmymSOB
kg09/FW/+KSbKJ97Z1gkGbGWf5MnC/KAJoMPgzjunNnDlYGhKazwb85FYwqOosAZ
qia2sQoMMMMY/qmxUOUFlaDB86N/ycSXTKLCBgn/DAYQ994uJXd3hwzrv1BheE2s
f/K0uxdG46qABtds+ShWbb42FvUp8STFPxX5KnEQRYC537oNlHdAZNQMbioQvPSo
qkBCGoKFJtGC59eELOhl6WMvlx2Io59m2afa8isDELnjuULeCQ8QUJK8p3oqYT9L
oykk6vC4YLd6cqHvuyTiMCsZT0Cr9f3hnss7+TBUAjAvBN1clVRe+p9/fgEw1P1C
p2SYfkCX4oy2VvmfgreCf8ont9hjFyxm7pbgpx+q6UIRXvp1pWkMKsqvSAoaz8RZ
9ZJSNWub8a6HOFKPRawm9q9rf04hRtusn/aDPVyY7Q7VjavprUQcpv1eqIl6tAsL
3hER8ZqQrwApXVPH/fqIr+DvLRQ2m7Ov1h2mwrGSf+lx/xryH+mvkUdrilvDamzK
K1wN7ChwNeVx3ghX7Qhcz5FT0HhKMaB+znwyvuCTNGi41MGUtnwudejt+tPD+YBy
a6jAYNCEE5ZluLKp0e8DWrkpxR3wY1FL7SYdfmJHxFCLLfCWRbWSdlIOXufVE5ll
9IgOhH15NlQfXM3nMxZ+fj92VrY2tUM3xTVj59hSBdSxB+2ZnZMN3/HjoknwYD3w
YF65Yo2st0s/3GA0YMq0JEK7ktN28Lh/kUlLoh5RoNtc0cW1v+xIQreBXBKp+dZW
mtcgAdbvarTp8yGLIfinW6dQWfzZJF12/7/YYOrPVeENiXZ5asfee1dS2/9hp/Dr
/nvhd8fD+d92BH/+W8do5VCSINPL6V8bk23p1xRKI43BrBiMzzL7oPffJdow/4m0
CNSwmypkJfT5xqD1OrPwhY++CvGh8bbRQ/yIYbCuG5YUYkDGIRxqXXETZ8Bquw3p
DfccgkvWrm7Jr+aRw+nxP20cZEK5jqEfEra0zKpo2Cy0GYEwpODmaL+wiJ18EwIu
z/BaVTkvSJhvKYfKBEtdo4QvNdFmSGE2X24fqaxUkRQvNBkVKob8k073iexJK7Hm
1ws1l2YApSSg7uAn+jGJ9v/cu4ZVLXSsL9eIzcHLcV8jgF3RldKpazIzplzhc0Mr
LgbUss7E6cQKeM7LWdGMDHAbFxQUJCfzihnwxtu2cfwDS5vOlPM5msooESmJXERK
zM8pWve5QEQ/e7nY8+MqkR9K9ZndT8r1HsYr+tXHT9lnbf6nm/+fzBQh6vqEiHHh
MiMNrGJXmX9leTr389hhhtIpU5bpzB/O3n7YAy44HRk6MBRKijSXsWyolNP9EPmx
3zCTc16LbkybUCC4oT9ZtljuRnOSPpTiZ4ylKgaRjMaMxz0Gow86hL1e3o5Z/Wx/
gD4wswECfW24dmzqG1JP0zBEmuEZzL9utAWN/HxeZwDbftZamLX3tHUU+mSoGP6a
kSJGwrWopQrAp2Nk0zaLhqERifH/OpR35CALvewIya2x/1QMQ95aycv5xKeN+jM/
+2frb+dugLeDC4Ph3g+EubjDWzDsohFRaW2cC8NDr200Lcwy3qXJHTgqKl2kqJK1
a4LYiUwVMqBQYOjFAIp3+IRLK0bAVauVuhEsTokQTrK6Ry3rRRUVRvYxlGmOKQPw
9wqBBTMI3l2U1r2ERi/Ja6ooCV8qnqAB/+VMuINVXT7rcCYZK3Sw6CkHzUe4+yuM
HlcMmRJBz7uA0Xu1PCgdkPXYYI3qmBTQL049NOAMocSdktySq5iXMOknVNlY7YvO
hEFnnK7FZlSh+FuErP0GNGMpbNXleYqclO5icwqI7l8U8Q3hHpWKmTK7g4OnBWUn
roMNsoJOnuTdCVZaPhCRpkSJVv9G/5vClCHCjqU1DYT/Jz37nO2xBR1U44zCM3KF
EMvEI4C5xg6BPltq4crSS15bxCjBTzgKUkuFmuOIgdH0aL638sWcMyNH+YIS26MR
U1oyBfNw5Q2g5rufPYTA+hdORiEETOOqraVf0TwGbwj/uo3aebwAWZGvqc0RjgxI
3fjXcSopXOClhRzsZUC5jW7pST28TNRbGLGHEi9B4w3YDod2tJhE4snku7c+7Q2t
7BAcUsB1nfIpvO6knohCbSw8pinSJy1av53j+0MKWO1rZcJ+6W6cO2i7oUm3qvyT
UFUO4osBJp8LB1T0XgueWoGP7BLSZSbnPYL5jTSOVDmLOD1GV4tIe+74DOpKcbS0
/KHts6vzMFx8CekxeFMjfqTf3wf3JPcdWfl6P1qzvRClO1JFNQ0ItnWOebOIzRud
vFdAl1h55Bj+JrDRHMCuUiGZ69ddAH6djqFWnylZIpwtlAJyY4uKA+IyM2x6qTcD
qGROXTjC6q7U3gI/TIMIBtR650+gZaWSWNxKEQuOvJpB7cfG4dz5yFddqGDf4s6d
Q+BEWHEZGp9VE0x50Ck5B+THw3LsDP+NkZ5LqcqIQTJhlcG1GVlicMfY3BgjKyke
fCmLGxIqU4ll6r4Gq00vKx9+2XosPjgeiw4jFs/LYufKJJ/G5vNjyQjSMYH9jB9b
8dKWwuMx5Fs7GyyZQTQUs2cBqUkQ4rMbqjsEYqjJ/fTDoG4cwSDEcfiFfs9EfND0
uAxUfvwYFV/GSdLr0ydA6QkTq1c/eoOQgnltuoGlDYA543A2+kNsK4lh06brjtif
HE7r1CKKycCwKq61N1Z1Q0YDoPqGSo5t3hHTDmFA0DVVOYlk+AFf5Q7W4Nw90x5v
TXvn+fv5kqTZpAEGCduM2hLTMtMNWGPR6oyuPu8hA4ghG+2CkVToFlcanlpLZFQ3
qgczYcJgc+5mlIbkXNTU6VZQsyGJ0R//rEogYot20eoX6RMpw3AidT4kUI2mgEJ6
CULXAS3wNQgNQeWwWtgnEnCoBAh9X07KXximxp/37nskNSPpBkdbwMjLJjxMGSuy
MYHfZAFq+GghFZC0pbkDD4hnqjX4UHt8G+9UGqJecru0FbMvcUE3hah4eQ+k6jkX
b5OkRtawVcQjNzfZb2Aipp60hzPH6ZEGL1OjFlgLa+GF9ovV1qhrwGNbrfpGVww/
FjuQFfUtR3H8GmwdXrgWzk9cfdeNq9wj1/7iwe1Qdu7z2e+eUVqr/IPtAjV4sIlJ
o+nRcQBZoYvR2zUaaA6mnqirFflShvZEr30Rh/1Lef9PYmqNQb8IyT9S8IIKoqVA
teu2LDVLOnvDy1UvlKS9vSjBJxtwhXMVLqpLONbIv/+KTt1KormRXM8wxncLHSYK
I3vWXFUGzpv5MN2OyJA+cvoHOzWm4ujfiGlLKUJtKkQ7B9ppO2gOuIpwd43ZJK3y
ceL2tiNhwHQUQBixmAfgEU04IMvd2g0+lAhu4hSZl54xLpX+xk8v7Oc97/bHt4vv
3HHKMlxSXkdCCi1TDGQ4dSP3Gg/hiJ4Dw8doxvw3i9ZCYgQZuKgwQwSZZgBig9oA
31Hj2Jwnc7i41DqCMWm4fKsUdpdGsLhvihW0WXm1HAChmfmW7PdpGFp8IxImgkn3
RhDK8ezHsY/NqDap8HRGYtf2SSdbf1LX6CFyMfVS/dwsUH5tKGLsFWnTov8t85pm
l3pWfOE6B1ScbSgQFKAnb1LkAgE8CTEdeiDaBq52nZ4CZAvyFTLRT+lcK2gq2aIK
+e0xOL/FgDD5ZWXvw6QK4sV2qye4uSR/K3cUxV51+AIK/FQ79kgl+jolRgdlnTbb
5IAdqWhJyvBkukZ/mOjdNUMNbC9RMNAhvsHzTzfqwb77UsUVnYCClpru44UBS3np
h7vu24y3rUh+lIXq2juwa6PyW7mFgC6WAafBqDItJ+aRRoKCK57i6VuQ93K62gWl
QFyXegmjg6OE5DlVecA9crpB/s+Re4z4iyPnoRnMgN/wFgbtLY+h6ba2+/n3XNzJ
184weCn5RggV6q8CfFCQl5uRFAn4OfnaU8ynOu+DUtrwW/UW9RVf/spk/GUhbISZ
0hG7uzl4Bl1OrvQ3vojvf+FlCdQZyA6/8zTaIuVI++vYybazJVmcJPN3N+fj2eXd
B5nbMxDAoXFcyBccBANqj/1b4hoRP05SABdxXct/ID0wHORf2iqOvWvo+7yuIQoX
eBg5m4nEreSz9c4ASFgEqUq7hLd+jjXL3cYY9HbWG1N2eKIjK2F1QIl/Z3FfCRIh
FCvpGDzbe7w0FgX3Gfpmhi0AZ4M+6Aoi9/qdd9KojwGVI5ZiD62k5z44+QX7+AvP
SHA5GflfM1QdE1J810ZK7cA+0ykUguATxnatByxvd99Q2LwRhWDUNsu6eBwFPh/b
BZtPMvo5dR4L0oIvpqPzyHwsU5z5ae90CQigG/vaR/12wxSRgT+yFj/oiqZCcWVS
IRCm8r0oWdu3r6qsW7o4G1yR9BWXKFG52rVrfRFED0CRwtllVymQGpK7BJpTRoOU
C4wBlGnOdFpXXVt7dbdUI6icjNiuuOCANnfmg1IEfXRx3iUSzRRR0/zBMempSAfT
Emp8YJ36BWQALdMUHcnMkEhNYnzfTerpjEEUAZ7Z3VmqMN30flDZbT/1EBQjvWml
uEKZkhfuydTpWIhXb/GtiOFRNfzEAZyGE5Gb/1YQl0CsWMbGMBimJtB4BT1GLQXc
4EMkam2KXvjVg7FEAgdQFboja7JZXifFhGACuzQnfiwCKQc54+6EhFC7fp27XcTB
tbOvOiBMi4noHEaNwrdc2rt7Zn8xqSDbxpm19xg1BZwTuzzBlQz0X3bRwglaWWeT
wlYPGnr4IReSLYBPKoBMTGqGNpfyM5pOn8M81YC0ydLJ+SAiFJeE5cc8hewHXIY3
UcKAtW0fMrcoF6M7GflAcTKFPe/xEh9hFEC9WCCq81AX5Uw8hIH7zfSC+xiq2NIy
iDs84pxLmeFxJUgORzP7vYUfHigOHMH9ykFczylIdBGt4u7/EGEiH0aAi050cpVb
J4GTqOPkCtDQo3skVC5PNNiTpN75bvyE0V8To0Bs6iZ6830D47iulwFUTqK8GSCj
sebuNafvmGD6fDKK9txCbd/fhLYkudAeMe8aidVbBKds/armDyP/kz1KIgqGoPVF
kJ/QFvdJ1ML4wjYuBuEzSPpBtWEQ/ztiJBSnGmghDTabnbebK6CSGG3cG3WMT5Du
jl2AhBJsFvwNlytMtG006nNJ6QD5fXG38VSZojiMPUeAB/P4jkjE7GYQsbXkiy7s
Lv3r1VoZ21NrD0ozjPQFltk8DlZgjYCD8e8O9GXgBUIcr9L3MmJYglAJb1Oqx8A2
52Hg2s3hTpnXGjqRoD3ArcWYuBnDUEMa+6oSiBmEsntzYdWN00tKDHnvUfBR1/xt
01TgOV0ZsvHCy48hd/NLtj4WEGgqHc2d2eLEw/QUqilGwEcz/UrmS+WQbejgjc+6
Z9XCk4M/vnnYLkk5kTT/7vBUsCN1h9GAwT1tLRtUAM27+J166O8dGQ/wAE8Q6zBB
h/iwhIl++ByNyssvg/ampCqcnVzZqo5jtIZkoulu5eOwI/QIvQWbdmenQw0mSFYK
ftC3Mzg9C3RVCNh68k1WmQzkks2fTjn5lq4HMxzdc35oQSdWS1kyoBqldR6vGQWh
UqLoBTVjFuzJxVpXLXqe26W6lO9kAYHyfskJ3mscbk6XOf8UAF8l583/D5LUta+z
xjrRzE17+5gWCTtEHEaXMcKuBdkql3LjIl5MkaLexqfS4Y8ykpbOTKRzeFsyuXhH
zOK9cZ34CGOvfomYAG4OdqSMO35EIGRqPQWndpa2EgDi9lCiO50MHLbj+d9G9nxK
5gKjyz1hpuUwTt0vC6x9ONuqiEDFNIYvcjGLobVxPHEY71jGIQZObR5e/TFZ1dRz
6H2tBoVLwiTmGeVjPcT9mDsM0FMkDhxcysvibM3zfz6y9bdRkO+pBV3bqw4SH+BA
OW1KGNC+5EdtPqZeo2sphQy1g4yxLWGpk9ze9+y05JDRzxRfiuin5exsAQKbOAqO
0c6RU2beLvtGEjTw7VwZ4pCZixAMiydODgldkbqhzFaP1twMPVxApqJO7DIskPwz
yyA91OixSi0qUReOPa6pOKU+QqlNQVk7Qr00f6P9qZEfBl3CeWb5JsUNuIF7LSrZ
OkwEGcgUxjM5ehrPhc+stHCYhnPx9am+tlBnfi8r3XhEMY2dMKpH3ju+l33EFxmk
glYFSQpc0vpsEOoqexkK4EPoA1n4Mr0DruFSsjdqa6N6PaYcj1hMPZrrYkdGwKbZ
9SILnh71Ck46M04eLzq5wRkSr8BpsOXIPdCdLYYmf12KUmh7qX4hSgvZf/MBu3QP
1cUi/UQCk4gE0YBFVaPquXn19wYIVK/dAmb2fmNojX/nRQI3vgSUML+K183Buk7j
56MGWOSIchRTtxj+83RgjGcvwZyyi9KMv01Sj9rnCRWSHL2xPNqlaPyF8/RNWX+Q
yNguSMS5RBwgaulLiPbP8GqqsMy46+1OeLu3zdFI7rxurZYrzoJR3FeV6ofbNUL2
A/WibLqzcJiZPafiibBDUDI7GUAdpi1vjOV9uZB0Sd5MtuQXmnUqZneHAvlYvLrf
akhdiM45QfbbqoO3evINAjxctj2xVC8wYcSbwliRBfPsYg56FBPuLrjZ5ga20dFV
66+hFyNehnnGy4twmUBFr1VkkiAKPZTSAmEOoUSvIlhjrIcGyssL1ZED5UanDzCu
H1LMlnQuGTrFO7r0verVBt9k4b1Y2P0EArVslgqypI3JZmXIzeQ7AlplJfZ3f1iV
50S0hUAG9me+BIyjXzCq6nCTkrGtuvzybXeVqQ1FUsVRTl2vnWRUH5LQzmYXBwls
JAqNnctaE/Ux+qhc22OMO5aePLFH+EM8n/kimsCAosVuKqa2CYfavWPX8Egre5bS
gj3MMdT7dLmnPcqVqBETjqLnBfYAoQUeAHZ5b6QchWa8usYHUiWPpxiXVKm/+wdT
6Dl9JArMh1v+lOL3qKGYkUvrUMXSi6p/jbcpzg4Oc9BgRnMjoT2gckBkwS0od1P1
Jfpm3pYlAMjN/wmOKNa0DvHicFwTXGnLC2UwOIN5xndRTeuumLrVjK9ztUGXvQnW
D3CDqmJSbNFRttDp2NEH5Ca+8ZbLTnyG25KzK6KTaJf93zl18Aki1Ken4/qU7ZpI
6erFhi1+w3PlrC8JsISaBapJMjSN2LpirCxTbjvu1Pk3JD6q7VNgzXNO+S5kO41y
41S9g6LosAKjNV0uj61o4r2xte0l40r9INrRJ4NjZal5pGBe6VW8SwqUyri2dJ/4
tRBt3XcSUzyZp6W4y9DQ1+3j3fy68sNQiqSupcXhMjQnNDYVVDvR1rM1KOoiasyD
o4KERNUBWRRdsWa4U46ikspVqH/C7g2Q8tb5XumvBxIs4iLNHrJMTU6I1OhlQHA1
snHLAxvcYxD0jpq5kfTwzL1XMkoQdkpAAGkW49IL42AE8jH099lfzlyvE6vnTN8+
M7HrCyQav0Or8g7QrSxuZxViQBP6gElm4WPKkB3tzcWSPbjP4OohSBAKy9t8vTdE
zUB/ymnOd8m/xwpj9NZgk6gfq+aUfKoSd+kqixcbQttmtr5MkdepFGn5OsBjzsKR
KCs5OFp5Z6Vye8/Ui6LQMMkJi3QDLNx670o5JOqT28+kKqL3/AAnCVrZEDQKoqYe
/AZ+InTAggg7NaczYw4h+dFUv25O4jsKNHLkOl85sI2udwC3BR4k6XGfRCzjUEo9
Nnme6Gn8pa39V/6qRdoE/F1lpZff1sghbwJXnxWBbCBQEetasTufKpvtdMuVk67N
Em0Q0+6z5PNLD4VUxyi0ELc/G9StQJmtxUvKKl4ArgfLSXVzalD8ji/X4Zf7jlmZ
QmiipStT9z/FP1o31tvQGlmfCO8v5fnEC4PR4OSFHKehU4s+99LO6fvmiVD1Us7C
NP5CsqEgVaYS0qhNhRCHEb/3Ts0i1m/Wmckc868lmPBuI6oFrAKieDDsXYl/p/JX
9YH6OixzVj8LKCI+9k0T8Lg2EF/UFzHCIkLJBsT34Cvjhyyn1pd7AJMKdW8tUAd4
qB390wHeNCQ0uggZRk7Ra1R2iSVkHjwgY8hqlnkJQsY4BmXHFLj/SzOhBNT3Or4x
oXRwnGlobKKumlQ83bc+Mz6Ymw+3jwV8ubxvJ7xFGz9qtqn8Tkc+KNg476uGVC7r
V0C34cAV4NGQCHyLPNCNDmjhLpWZ6sl6kKx29nxCvRADEWZwAxQFzD/CduN+WdwH
4IMAbSyaOKJ9kEfh5obLOyE/APh026x1wNLgBoZqzplho0dyDhbRYLVV6gI5yOti
pwszOaEqMlCMrxY0NRXC0gM2a0gOoHyLEzCO8CvDVWFsAZpvYF30YOguxqB3YZB8
K5sbsE7X5QPmMrkc12guOYi1atXwHWS6+IcetZTQrg6SNb0XtJuFsboqi/brWfXI
z9ZjEirXsJtlxVW6ziddnQt25Rm2plrAG7RPCEFeZEYTQEsAyah3fzHF8ILapIy1
nL0fE6Fl3wNl0QxR6QzZvOvxjg1QQYzD4JtJ2cp4LZm3mVrKB5x2nRMDpnBkcDpQ
n+OU0r0qi5gbCKV3EniDI0t4l3cIK/8I6TR/kPeCHRIxhVTFbc6HHz5jLa+2uwjT
Iz1oykmdrkZU1LRRcWeUsOkD/8JHs1CEVw9aDK924dB43dG/qh0b0zoQ5P/FEwwV
pp+5mTfIgyfCmxypC+sYVS2fmA1Tqjylsjf8b2p67jthS3GyTFRNuC4fAv8JF61Z
gvsJ4YuSDIQ02E6BvfyRIiN/PvP9n4AUPNMNYg2w4Y2Y/CYNoJtqS1JS02dM37SP
SDBL5zc8rfOF7rEMHP3czLRiTKj1xh4Bv8YfzSOrBrvW6vVI6abSV+cFKmi5ODbp
2ymH0VVlpgCp1ov1T65iTSB7ok/6y8L7YBtaCM3lrZq9d32CWTxJyvSUmihxLuS2
H4WGTfd5YFDOYMJsUz6VgL14LhQ5VqHHuDA5/Akh+UEvYDUw2TIh3/c6sZocTeAs
GEQ0vVgNe2eTuzYS3APiIXXOUAGjXU8e4Om1oqqghc81MbDrBEamzY05rGW9iIUW
SwKc4mkzc9TQA3AVBSAir0Lq6jEg6DB06EWqGR7HXXInVL/jIuHI8GuoyfEjERFa
hakfx7gMKn44S39FFom904JNOavKUHryNa8eTkUO+kT3fvZ8YoS7kXylmN7TicvB
/gJFLaBOV3WR55QZKCF7Zic9iOFK5Q3Bqs/65FrTCqrRdKSoxK+Mx/RXL4hWW4Qy
zxb98W5YdkYY/RXJ99sMDRX/JwhbpXqk8mSZl3MCQlFTN+we/cew2xSP3hyxTSNp
Hk4oPk5enm6zcxJzTVSYvbAM9yJSjJ4p2P5uTTWG2Q+I5c5fA1JzDRhZ3JOCX6b8
yLi3A56oSTExPxtYWkaMfvwv3M4wyQJ2HKqk10DxpYWTQco5xkP+ZfHTAAtm1u/r
1uKldqoZa24rLUH4e4bdbnjJgFnKT18uXutS+D9uOnbIRaNq3+XETlJMUv1KHjRu
rCOAf4Jyai9b/QUFnrxE0wV0tS32C1nxijC37S/7rZz8ToHr4OKHmcWUDatgPAG7
9+pCV5WBtMQgaaJJkQhikyYqQaOt9ZZcuJW1fXJOB0OkFPdkTkUKo1aShUkvxpo5
yT8trZrMkjXGarpQIl6fFxX5SBald9Pl+cr7787MzknaCcFmqo8UhS5Ds/QwLnR1
kNTl34r8EiP++EH6795j9HP4MCpYQsDN8j0hhMj7uRD5nhu0JIzLk/0MP4CtNP++
Ff7xJNZrCeA7sjZIBTuXMsRsNlpMCmcknSwB5jpLygqkFCZQ/DC9V/75L5TkAh1M
Z0z4nLdCxXhRigMW/Tc8ZPZBnhTim0psY73d2USVfAeKKulURyuMKnfpc8FOm0IX
Y93K0nDKCDIQyvrXerlOJNOXIT9dUckwIdjYkvOcUifLESqZTJmk7+Fj8z0iA4IV
qDvu2h2R97Co5orl9X5pAUZAxPzVnnINVJr7xYnvsTSezFj33LXegTBqGAJxYQdL
vZdmFYy0/R0Wx+sD3ljoAx17vWG0IAtWqPJG9ohN6foq8ugDhjMxFCJQepNRuyYE
e23NCFZUbL9mQOec+cKBUajg9rBm8taP1xxNSvu7MkjrRIW8sBRyLx4tJTXgRPyg
FqntgLHARZYEMuurHDnxTESRqtJV2YHnX1EHP1InlsBsmUavjHuq1h7pMbkpKwpU
skuSmyySbbod5/439qOHB8zbYEPRwJCFMeAZKa3kV1cea76U/loW4uzsoJPyb41n
06TYP7WFYn25+NWxiZuYm6+7VCeIx60pDmHObUrHGmWups70OAuK4uQcu5RIDR03
kgvHqsROZFdg1++krZiZHH4TPnMFnOAFmmFhbHolk2/vY90gvaNXJ4E/1MUXHNj+
t2HcRB5CHXyAI+PNxebfSs2W0oWiQkg64+B9tNVXjiODGzoIdtdTj37GdfRsRwzU
ZZLtUrobUNH95Q9M9crysh2n9+ydu5cWtxlzmPKib45LyglDIUlVqpNxns4cwaIW
ycCbrpB+JFzfcJimhIWuL6MGtnypoDcgWamhXLWe+VuCwQv6SilfQRc/Pb3HnrRq
R43k8V16adpekHGretm3qG6960phmddngFtpzSKH0acHxzTHnkc6RczeP9m/tNR0
P0oSDxOup9GmvMVNpk3fynXTMAoY2IlUIOtB6/lSbRpwO+9hif4+wO1LQiVPiuVB
hhtuzI79PML4QN8k11iH/Ox5+sDiUM/6RDkUzZ6SO5vdnHGyWZq/tOIhgC/awua5
3Lk5dBfumgA+fWJypKMBpp2Ddrv///g091XVRUEnV6VzRsWJBM7DJ2IksXgH4qmd
f7nFJzX0CtgHAnJTCL06dsl0TSFCa0RWCtDiimF5SDBQeA/BVWk8W0+cGtoNt3Wk
iuE1Jdj1KjsAdy55XUQz6ftBjqj+jO0ze8C9hJqOs3lPsDngEj5p5hNmroQoZOr7
NnBKhmy7OHZNTDehlrs7yml4egP+nsFqF2/PuWZRwEOv9VN/iSJpFn0xojUAUYiZ
zn6Xo+kj59+yaU+DAEV34ejyis0HhN4olg1AWOFSzx6NZPuAJiMmbu1c0TwsZ+Se
fOqrBfeyfub3BBl+T+yR+HLGsS8vbPfKozpX2Av+gkCsaa5asdkpjxUD9QX2gB1M
u4uqPYA+uHlRVlsarfZ3jnftKPhnWslHdgBpebvn8frHr7PtUjBd/fzrUXF6bmEH
DZ0QuZoIKAIGW9uur+CEBnuQAjVScMJxkb7d5yGRYm0pxoQEJBqRSwqT7ymO7yBR
kafUeA9NWrWNWJRCiIaND3845P12Yz11EJSIs+lNsuyFCCjCzhr0gsnMmW+qrOpo
QSNMmO8eZFdhIKP+2EqEVpSChg9Nifr30hociKPAiiSR+EIRbQFHTmu9gKzo8IgT
umwDc7InkPGZem0rXNlKcOwLkU4u4lU3FzG8oW4wcU/+1CWOpUogofIRzEihXP3Z
s5LuoOd7OCdEKEUJJ7ASI0ZAGBj+FBXrZIvV9dEfMF9q2FD+l6/HULlVtqa6wqYI
Oz/QPE42SrkQV6rI8FL1oPE1bxZvrFQaPYMgIgGHjJlxSPZJ8EpIrp+9MyYNcM6v
rxe1WBE82jSi8d8OfM7n0k3ACU9hb+YFulf+Jq7fg18RKJIe84Xugk88q/eN9DJP
e+F/Cp2Fx/l0rr0zx7WFG7FR0KgHlwLWA0s16Aqbi/W3WQh591IpeXSWPq0+RbAn
Uv310pCjKuexgvkdZWy+Cf/M73YztP1kA629HrBkMgEadQqB16SWhMDbFoGuPOWD
UQedkWwUF48se7j/yqDNi4VFeB6KBlRKtQVXWQwAv0z2yf8RRTo1atTWwHhkREbZ
Ylz1jz7YtL6qvS34OnUAa519XBqMYvG1ZK/22c3HzzNI1CLTmZyJbPnKDMKd4vcw
JigiUEuJZ0KUB0khx8XmK9xvdIVSZau5CVOStQfzI0WI4xsMha9g1Er4EPxSlrHw
Sgd5A3Vg+OP4rBSvIHp/VpdcKweHg8BPXGDcErGtfIyPZoFb5E7wHpd29m5aJUlR
ADRweTA0vOTKFA86vuUDyHlhNoiCnZoptKrWVGJqWjfO2q6NyNLpvdU7rYPwaUgZ
cR/8xpMWO/Z/5oVsl5AJWfW1L/iYOtw+pFgWa7yiid0jnv+R1xExwaUdZDcJXGfo
ad7ovacpA7pPhmdoYFzUN6nNs+VG71uX42iPoKL2/e4lbO35Vv484INCHaig1qiR
zXsq3yJ9hZWqXg91PGTZ/eXtNIWSOXKfra/wf948HoL5XbMR2KnUGKr2JMnu0ABT
yomv1n7/isXGUrzqifTTz327tSk7QE/S3HNvr4lJBKi2EKa/71YwBpJ0SGD/5La+
6pINgIAjgF4AZBvst7+0joUCtNU3buC2ZuvwPwcD1Wqvf5SnCbh5/h24bihyzE/C
/5w8DO08J9hdd4f7ql9R4+cbWYjhuOYXenaFBr0jijIsmD5MUntjPZAd0F4/GAGq
09DLdk7G83d+BLbH0IYklADnnjRX+zVxTPhNjnBNq43a4UFKJQ6xA0VzIC5lJWDi
pseVop06bWa37dk54lLwDYbIyCgUtW1qGZ9KRcQFSTq/EL8jwkzSFVkITzISgzvy
KUN6Ms7VgSeoD7yG69vhkp95fIwYNlgxhcJ8OLlLXWaRKeUfOSzdwpou3jODiv7e
Oap5YFwX7tkUegfB/Afe8/ECjQjKsTGLoCRnpLOiN6pTOtNkMPE8N4r26k2aRjzb
kNhYZWbr7VWE27w9OK74mn5aant2Xw6t/gDgtuhUvb7U+fHXjxImCzmICCI9rIQv
gWjuY21QxiFl6yKwgela77ZMbp3/pfjdAKdAH0z2ZMsIw0a+nD91nl7v9n/ogThH
NpI0pW7gO6dHPJqeqrCtNmhLf2AM6Bj4qDxmCnyMla+GnAFFMALOgGanZLKYDuc3
lKYYerlvOdfDCGVmRA1JYF1UQF8G64BC8QhdjWcoxETC7dbnMC8rGn03MhQ+a6I1
NFjPDx3qrF2Qc5f11dUoT/OEsKzNAZFx4L9SvD5BzUMFnBQvvdZyogYz0pIb9+qo
rg42YUVLuVsJMDoe4Y3rG7Jk5BlsMJAO6dYOSBeKMV/QxwH4qX2cGAhGM6s3axoH
U9SrU5cCodbdwxM2sAs8LPO1B5gZZts8kkQ4wIZkwlxgNvSFc4zK1/tWb5JnU2OV
90cAukue72rFYlSHQoulibzJm2soQ924REWByYa9MHJBUnj6wT0VVrosXIAnC/bZ
caH9XoABvKTZ+YNdOePPWRDQOyeJiyQv5E06SpVjrIgIriyoG3cREumjeWTBEyNj
AkDIfCeUaXPw6RcEGUB7QypCM/vwTLEEKq4jQXCUB+9GUTCF8SkBkJ1YILk/+y0n
RxHUWFs4Tyvn6+u+8if58NbDCHKqWj7jHdq7rhLOTR+XoT1GHQ4rfo1qg8VMe2Ei
aBEQdeVzxMGK+IEe1gO/reUROlmh3chtM3W8bV19obBTHf92Q7U1AjDHxZVzyKtS
naKUrgUJkjEZ3dMUQabQHH6AM1oWeeADF3mvhC5fke+DG0qySiL/O5EeYqmF58gN
mrdOwCcYH0iyRrtXBx1ibhQb6W8fikDSGCo4wMaoMgcLFY+XmDqhtYfEV6bqhUsN
CHuRTH6kQWTdawwMd63ruVPohCTT5XmEZSydyGVkccDJKeP/B/UXqwJdc262luUc
sxQNffDBjsiRg/z3bfGemMNmKRiTVE9f4K/Tl0T3PC+OwrXjsGpNNYg0MxOrczos
NGY5D70lWhUsELv0xzJsVeJRu5IAwNGiL9/JNayNjuPpau5qNSIs4RM3NqEiEPhz
hup0TffYgicp3Z7TEHI3wKxf6Le4BHr7zXkW1hlXm+mH4EB+EM1TFH9Bti3SOgu3
G49oGqA6EzMitDc0r27TsTF7XHfCXbG2MFRcIwHQEZeDqdP3juod4fAAKfMAmFR+
cI4rwBO9NXIrNn7smGA93s9p4n02d7FN/TTskBX0ryFQHUdyh5Iqo92d4CuaQjSz
E3ZjP/e3grYU0XkoCfNVYh54VboYb0jd1AE35INqClFfPO7YEEv4XvPX0kN0CaRd
CXtOtMphADWDVr/yePpDPPuaPfCUG2Kjxh9eH0T8TdBmmT5NBl+6PDLujYTvh18s
narlLQKUbT0P5nJ3itFcSzcTi2UwfWuSxDGE7q/SCbSiN7IQLb+eIQMZOLuz0aDg
YE18dcXwDUU65NtHE1lk4tQjlTk2d5/FO7j19ssVEt5tHWK+lfpyYhLRYiq+gGxF
7n4bsAKT6lQ44wXlJv0iUZNBpxaWMNocQ1DHi6GLJIBWGSy1WTsHAfpbjVxN6wWE
9+Z4OT3ZmT4qHJaLXU3Ut+/edTyucS/vpXXUO1h5v+vbv9aXr/AVOTHTraC/BPHY
fXq0glm9wliyQ+6W9SYLVzmtnQKcg4kA28kPPygNlY7Pi9qkEh3MRD4bLs7jZ3+D
QWngIHHddPJEF7CwtQUjmkBMTnX8qs5ddof+BFTF0Ppu+QzeHFathHnenYalu4Nf
hwRZ3xogjsiHV4/aBjWu1EJq/CyxzhoBioZs0mS0OvU1NkynzvPv5nGi27A9TuzM
mKx9DfhTJLnT3Ck40V+ff+Ynst9C09k27WLq/hn/naLz1E/p8TzLuPo2j8kwVQlu
pq0g4DSKngXEHWPir3nGOVz5DScVVkGBvg4xJTvc1ouBovKWnw9AhtEH2rYHZ/05
bx9Ee197lisioyg+8dCboJmI3IeUod+YiHji2YFStzMtknpJlVPDqnu5AjAx60S5
2JWLz4A88DXSA6sk6rA8i9AIsts5vy96IZr9Z23ZD5iUKz9UreX9Td16vqCh7Sq2
wXBehSJz+yKD0EFlnbGqU81ALJSMZQCOodm10kAVozaTowgGmDbu6j1sELJWMn8s
qeLIb0YMT2hzroTW2280UOshXz7f2SnhW4Vl+i2n1nE+SM9fX7vYmVgapEZxcIGd
ttIjIky/BW8vV/wmbzQztBNtOMnyRsZ7gML5tTz76BkeiD+WkEFJXKACLskEypXY
Sn/1aIAzZB9rwa9W56Qb70TB3o6LDIqNIxCde+31MfxgVo1jK1D2nmIl75vz6QxU
Ysg/ZnojlM56FXeJU5ovaVI98jP12JXgN7aWOD6mnhLeW0lFFtCZmh23a1qDcvGh
EqrlWIM93Fjb1fPotoOiO7WGPRdgM7BtHqLkPNi74SGgQov7O4e4CxWRIVhMV7Ul
MdYp/SwZzN95Ge/OOWXb7vjd36nmfjUFVSH17D/RFFzxp9FaIvd+qkEurmaLqbyO
QLrQVefEzp+SLnH1/tEwNVhX6d4a3TU9Gd/u4x6y8EJXLjAp02iEnLNgEa31U2jq
rAWgJMnJOKUaUJy806plkmPNU5ArLN6+AWqMGuW7gfw1I7tQEw2gELnpSZ3JEkvQ
6CEM/qi00bBV11HG4r/46O0ITQhi7SmDqVIOvp6NRNaCtdqpTaX+3sSShMYLHs1e
Kppc4uXVjpF74e/L34G4EEoHk8hffW+Qb//GNwkCC0G7Lra4c0Eylkv+upHTMLmg
VKw4S3leVFa5kWfBfmE/BIqr/lTHT9ILVepqOZbz20cIzeII+RkTpBJfjOwi+Lu7
SVF17Tc48eZpDWLQwZxb3TItdQRVeQs0TmbUgcH9NPDC5zwq1ZaBA5j88Nis5Ua7
K/1JL+B3b5XqRVCG6d9tj4ZMrArbyF7EFkwP2roaMRoix2+1xOr4N3ZAV/zZAwlW
pDhTLjw/oN1oeTFHYgSV6h4WfAJeno4yTHQ308cr7JNti2MuGIQ0svmYEpJSxO0g
UcKX+UMocT8iIiM7l4hem/8hPE+CO7WfI+BNDUcl3jJuVtf1NLf9Be/tRIiNUamU
deJJIrOOSuHZhv1UkymUEmqZ9orKyZvix9oCJh1PMMrnnRoby9LgsUkXJbpwseWf
4QsXJXS3ECOkl6GMbkiNglMoW7wUGkMcARa/Iqh3ydBimizdG1tNW1NUyh4bUIjE
KxoeTxAI8iCicvqe/9bm1kGt7coGsFn9DYld44hGU1xhtRBSX0C4FLnZv4WENZqz
tnVv2qZWgzFgwzc4tuu2TzAkEDhS044j8yaeVPIE/D8oc9U5bw57+Ebe0Oaqw+h0
1l3V8cUvHZN1BPP8BZMom9kH2Oeq6/m4h3ZcGQzdpvAoC3qpeFFxepeRrLJZv1XB
WX8VrugLsRamcsL02+Djcn1HdLJuYCoXY59lNQzxZFspBRsA+d0tMXIoNKcFi6V8
AS/0QijnlnbpPpy/dZ28UJzDRG1cegxiLaSTQz5TyUi5MSnQ7/eG9xG1/XelA2NM
1Xgg+bodXkUTvLt7yepby7rQez7Em1AyTJqt2j5csRVHDEud+Q6lgwRPOISwY7SD
EzGx1XoY8eUs2AtkOcPbocO7+YWlP8Mv+tE4PejPvaNaSPSqLNc7Jwyxxffho1qz
ajVwN3+K3Sg0UgVd7GGq5JiFHqJQZ4mCiWbVYL6zBw2V4QocGpE7vovFX+YVIlL0
gRUBBLU56hck540aJ85sLUYPz2ftKHmXTohnZEOqTr/w8QICH0CieaJkltLxTPh+
/SBkIOMv2HNEBzKkvdXjLZV9Cso9wDJ9aH912Pc9ktQWG/Jg2tW9BH+1Rtn+DmNO
CZisT/HedEd5JVYxr0EvnJY/z9wHGsbbC24EIyCRRIfJ4W9gys1zP8Y8bacSxNSh
/xhq8kHau5YsQHVB0LbMDdU9c7todJmf7jJUcHQxVRUzPJkXSO8+ibtJiDsUG1C+
ztBgIvvEw2S4A14yDp7+cEWtmmZ/AlR4dF/6Slp9nMzTkmV9W6RF1q4/tn4fKaQ4
QWzG5WpF3EKybTT22G/I9J4hberZZxKyqGr/otRdjTexnDBL52FVzG2EeEkTYEhE
C9mav8WVJeNauhRQoxc2bnSZqrZ4fykmRruhJc7om3Y6G5Vmw4brbmlgCcbdOyDn
umMM03DyBzy9DLwlmrG+5I/sPHB7Vl4z2UbXE7P2S/m6Zg+w8RQLWfHQYYsvmUty
LjOTePaF1GkCQ0r1XchxAOOhcKL6cGKytMeTw3Sx3hMnTjwGgu85u9kDwckEPWpl
hKyuA3v11o+Q5XOTaJO/US5BSPB2BVsXHfyJu2taXrBAZFCNuJzBXD7uZBjUHJFJ
+nDcDBjROXIGizVf3u3Rmfy8M02/41K3621CJMv+SKsYic2MWcBnkt2ar8Pyw4NT
k6NbMSa90gKTlUoVX2Q57b8wg8Vc+JUCxga7RkWnG6Gv4C51rfyzK1xldOtEU8tQ
PlTJ3uUYkfe4jTBt3hbhF9qjnODyZagIeQ51DI0bBD/wIy8PiABdwqsuAEdwhcr9
QXgZAaHKDXq6up9TAl1wmlGDNerUCWoo/DSPwzmlvaVvexVEV8IYkOu7bUNH0tlu
gh4MeQtRyzkku8qw9v+YaA10CNDnUw/yMmrBpezQPcEldVFWLZBQQfaf6n5crdt2
/DgskqfstRRFe9DkzhIwKxhobo9kYvLh+ccT0qN1kUXLVxI3F6ouGGssWhUzSVFe
gE7eBX1q32xwf4eZtBISU838+g0BCaurVJgzc/DMhK3E/Krb7ubB1D2F5mW52wl4
9GHzlqqa/02VqNF+OFevhztcRHI7vxFSTz5YRsYxukxc/SqhQJ6oM3qAI2EEH4Bb
ZtAwgUaOuu6hob1eW50U1piMZ4HDyGwPSfIuOYgEFcdSoxNIUGsazkEUgz8E0MlI
jaKrE49+WeKKtJzPU3Cpzs1BFF3r55LeT2X7TBODHeufFsSpSYPVmgU+3C+8giZA
ZRrtrDJOqKl9h1c1oN65JSc5pTshDogM5yaLC98kjz4mUudjr1zsMViC7hGCE4PW
7Oj5Luj/WU6jmoKX+h+9kk8F2bIjnt42K4pqxeNdll87A9H4pobFWXVj2WyqVI53
gqEtjxmQQWgG7VcL144sS8XrKOf2cgXg3n5ZGGtN/D/E4+h5P8cQvWBCA7f6ypw7
8nQhHkxxiPEkxhgGDoaYIxjfOrm3u5sJxMmNfMVlSjwo8PZLJfKw1z97oRKs6P1b
Au3CrGFRvOO6L6QNozWqlYnCUNmoL6MfVdgv0na87m3yx41eGbxDUyGwOeR8Vsbe
rSP8l2j6lthl5glhEb3knYjcj8NDeFaWbA9wLy2nNYWpv/z/iqcUX+WZMmxoA+8u
RfkEnqbhQ9Xayk1og54/D47Rd7wxClVBvRBUFjko7kh48m6T0TOW20mT8Uf7+bIS
JRyf8R53343f1ixPFbc4+ZVXvcoLJ4J0l61CvWy6cd9aoe2lW7RgrPaul04XXRi0
ptRf4zXq8QCdkGTQiND/SqSwbVI2GYDtZ0EyAaVsqE6Bxac5h7wjc9XKqJSVe4+N
Bp/AQeWFIC0PpevvieAhwkL2mA8d9bhC1idnU3rjcFR/QBJof9hDmuU8gsUMH/Yb
kgGvAPQnHkYZVDsFmObgQvmwO+A3E/YyYRD5i8uCPiZwmJNMywi6UIpRq7THoSRC
0pM2C4aKmQTcKsU3vbWiyyy+omBNYSkI9GA9wBRaA3LR9ZSXenwlOH+ifBzaG4W0
I3lEtamCXMxZgjHeFf1JjN9V+uJ2wQKvxmb07rWhy/K2QntIWEYASsSavjJRjrat
reH8FvnwOm2dUmUcOVzZ159oDkQeTYWEgYHCC0FW/LEk3aVb83w7M6CA8/roQ/fv
yAUmK49K7l3I/l9PwhQ4Itws6NChdI4u2mPnOJic8Tx3fGaBivOjRJvg4DoYo1Wu
IExxdIig+sUH8IteG7VscYWBig2bi8DrAZG9xsohad/e5fotMZaswnUU4YWRPNXf
taEfNyEOLmmg30a8/vFGD7WAgqgH1lcDDISSvIBzTyVVWUYNnfC+bSrux4eYHUcL
kT+Uvjmr/dcu98o8ON3/CbbuA+2mIIMUNcececifOiKhObsAvTPkLLH45u7M2Bi4
pjrW5wfhNK9i8uo1+do7PuyWdX3kqF2R94bx/EjBfCDEnJB66V+YvhpYmYq40MlZ
dGMdHRodosfOTl5EGooy11kZ+HpJcjEjpHTVXWMCs8BMg1TIamn7Vgx1V4xjStkN
aL4xVJEMuE8yPbscSb4V2QEe1zyqLv6S/GHqvuuIulP69SrQbdtztjgFocXubyNt
yAUE2wINqdj6iglgEhhbGmuDJB6X4GVC+B/bJ+WI7BWPRsj+PSAYHX8pAZ9vl4Gb
RYMdgNmVEBMmlmgWb2T/DFb1PefVCacct5Fn4n5knj90P7mbHKgxn2zRNPD6CQxf
P7OtHAnC40gQL0/8Wv91RlURsTtJzgBTrhVXiJ5X6apso/9J/LDlikJR9MJwqvHt
e8N2JYWTBCR2tRRFF/bvk5r9QLdFn0nro2ieWbNbh7/eBup+c1LsknetsJLxm4GN
2z0oOCs9l+Qnarnn4DFXubDs0skoXnZvDZ+HZ6MzzoS9HOVSdthQr3DE9AZbKsHu
E3r2v81LdfjJJg/91eBfCjWJgZ5BWed0ARLznZmZ8SHdAidi3Py92OLZnoU35eKP
N8VO7pkR4+nylubGq80kqeCN0yMO+Tt0gc+S9xyBGvJYTo5VWOfGNEIhuR/QOU8A
XvrvcZr+3K2H8PhsYte2LZAps5H77lFYrz2LwhaA7PYEOCaac+OfG+HGIR7bTE87
IX3xgoxg0336bhrU/suwLWrni5bAopn8I04R7CoJLMKlNU2kPwd6krJv8T52tMg4
rKopdfVGBW0dQYgNa1XsKuxzTsh8z6K5/qu2OF3PSLFe7Ga8LqR6Nm9LMIFQSs5L
i+7oUwabinEylpodIwKUjC9BpAkGooufi4EdY15MuLeludSMAIBoH2Uj9/7Qh8Yj
PGBG1hiq8j2M+yEpCQ6jXTLKovrllgPHAqvx1eyzrDfT3+rUupzxEJ1uLHkQSlmf
pcTcUNydKUhs1SNRYNY8fsaFQDw7KbIdSKrXN+uEMy8AE4JmZgvAAlihetxWeRxW
3sGUh8K3HRXlqqi/2Q8V/JAN/JkrRwSHXlm1Wlly7E62HYhjQZMgAt8946RNumig
nQ6DmyuvOEIYRM0ODYgbVzVG78ZdulFOKWbolVdnd6A/kIYxWzU6zn6C5hUPqDRz
qAM/qZuHK0Pc1Ii00zW6Jka7SylqrT33H01i6T3nzNxGmyXpNMahqHIir6335ffP
tIl+bYhqlGQct/n/2A9XPAJVf8kHS/BA9w9InygRMJsI4QXqRo4L1+L4em3aR0zm
g/+4B8nhHNGoNNy6xzGARELMNzn4njn1Wu+8HfoYCoeypZxv8x/VRQOfL81IFPA0
4Vkr5b/KVe48PNeMjKTjNZsCqMnE8qybUpOM7vygGSwjyoSdo7uEQwuwaPsRlx56
FuJ8nYCVe/arICPRK1ZLEuL8aip6tXFroKqn2Br+SE8+Kt9Dr2WHgZw2OeT07YbT
k4lNACt5jnlIkhsq/6/cObB5PSyvfQ8rCNekOxR9cRYuylXuC5nF6jsxI48FkbfS
6Qufs3qEkHnmPc3mb1bZqlqCRpXdCnq7T2ynSihu5QiMi/gbMNTrZVKj4ykYIi3d
WR1ac1C5eZDP8ki4HDjkHVO39ZngOwYWrMzVyjSlBUh+Udu2SsnO0y0cfOOW112U
6Asyji5koZqvucE2SXRFV6JgMlCddRakblLb/810mztoO7MRj8g3bEFg/xPsxban
Sp++2dIja06BBgzM7xhWfnRQ60wWYHYeIWsH586WBpGOhP8GaHBkr4tvXGzQDPQZ
rxg3Zl/Skrdpt4t9PzN0i0q6OMAE29RKXNH+HwxoXcx5k3xDgNls4o9w/mcXK0ba
OPV/x+z48eiSLh3D+pkVN5UT4SFQ3dHXhEsz52dDhnzztxeW8YJUbhPNJKUaatgq
1XmYxr8MfTPI9ECCOEoTDC95moxY1qwxsCb7Ifm68vHh20q1w/nY7zXLhtg/Yj7v
tA+cZjfxn4fFpcS11Vnic1zzsZYiQSGN4RIo1n9kEq+LosXi9n95bVcCSE5c6AHi
3ojnwgnVzbSWZ9bJgJarY4Bdxz1nRYTGNbjP4j3dMBKwOr1g7t+zbBbQdEoThdMS
jlZkQP2nns9w/s8w07zCNg6ttd2ir9VHcwTZeh8xoJyy1cCYDMgQESOjcZHYRgBW
yKSvmPEeTRs+6EyVBk6WusS/UmxTy1wx6+ca8khcbMq7PttgAXAg9f9Du49SjU5B
S4eRPtGcDwh6yrJZ10iy+F2nEflyin3P/PWn6pgdVgVQsfM2K9VQEtorymCE52+l
kVt/+x/LUe83cYM04cdwznqtdNh285jsR33aT7wHOPa6+pJEcJZiB8V6L+dEVtWD
UBNWnLQM90cOCzyGcCcy77W41kntaRHTXkMnZKlWD5bKHj+DS53p10HCZG+oxd/f
rG48+t6PRKKiCqjRhs6HotmPFcpO7USkF56KAEEDKU26SgQK8yugux+bSfYDPj5N
CBHNYNHBWzSgFt32Id8HA7HdZXir/jG6L7LA0zuLrnVdKnkzRwJcvBy/1s9ae8+2
4THPjUG91f4Bf2lXQ4TjYbl9mlYvKS1BqOuHwusKtny+ImDgNyi7XBPojGkThbdu
Vn1M5oKrrgJbqKWs3OptP+kKYI4l4mwrSAJziHo5OgJ2JUnMjI9PBWZqq+BfYcIG
q0OyUv03bc9148vSW6RwIJ2fhp3GBbZ8ouQPlfeUXI/CDKShOwKSCPwAjhw9m9fm
UOl2lpXrzKBMvxBO3T+ARjUeF/NcHKWuLQ77pmNMsPBXotDyeVyRctJaRmAbRkLg
IuGOaUGVyGdi3+9y9QVRmPoktegav0yBraXNRPnkk08EaSJ1d/7M1nXc9KD0qGcK
ZltEQ8hqsj409rTw545QlW1yWJw09aciLlqHQ0lc1iqjRDlHzI4JJ+VHL9/d187y
BUZDE7cDZFpYaF7yti/X2NGyfK2EqNW72BKRri8HHWBRq604jgmGZBCHudZFcJ8Z
tasmY+iWnEsiaLjM8rrzlWrdn5cyuJXPlddoUnI94boVlC1Rbk3uJq4RtQyuEYpG
ezw79fynJgrZ6MKVh0gHwWT7eiVr3FW6Ph2gyvdAzhJFEG8ykJKC1EZJJ8U01Wwf
N06u796P9icci3QZF1+Epxtw2rYO3IlnX7ANyJzoJ76UC0hNbj8ZMbwD7Q9CTC8q
KEVGqOgivA6Es1+OGlJk51XEXcUqp1Bp7AldK2x+K/3i/RlDnaIqB+hvpFOYxiXj
uugmE6XlRr2Kze8R91kzzlMrkJwxAzZHMDXxdWXY1v9Zjnf7c/kQMiO3Z8wvkale
nKhOUY8DxMUo1uscykfrz4phw02vPvBRuYRaBdZGbXQSYvNQY8diPB+52RRD5i7s
3wTh0okhnFH6QSulEH7Slegk+pO/1axR8P6a3czqj9I6dFCh27z4QeCp5HsqRAxy
M/ei7UQvpjzx9isA8uT3zfJN89631LQyvsLeF5b64Yu2lVD6Ez9GNIRyjFXhIuuO
GcAhyI03Gda2OmJy/akursFlth/YgUqNWCVIoy4NEEf1o7XvPGgiis6cnDvmp7xp
jTjCJ8yKommpRC+x3GqkJ3fTOh7vyZGL53uSIfQzUNcpmK3WXpvwLF1qnmY9iLeO
qDfzZeBINZug0KXlbY9SzN+BpV/mZxp8wuq221eLg74Mq0G26sQba0yDVrmtWcJx
7znoVYoM3QW2y6wDUn9PeFNQaulz1lsbreqNHg07vS+++qjxaNA4ibm99ONudqvb
H7m3ywi44WCLnFyzcGddk05tgHe5wPnc8o+/QWgdVvWVyQh4Z5TIl7mvZRsebCZr
kjBj7XKG16ULSe2CIvvwKFkUYuBsqPGccnyx3yrNUhedXZeHoc+RnVCR+8vTUEld
zBvhQlj6zBXinTwCqEKHJ6cFyXN7HylSJnBS7EuB+veaXqcisZcSWp4N8M8Fz+9f
daZR2Cn4d805rf2juRK+eiO47g5+9cbBEKnK07PZ2xZWhP4k4zMx9ALBBRXRBGBp
A4UBbbsUtEXsU+hfMdxWNFG4XmyFNjq8FrAQr8kqUKMilu7UDXs3Ka+CjQng10sD
F3JKwE46EteV2Su1SA4zIo9QTSlkqVbX9OcXFqVzLhlgDdSmx7LQn0uA7zuuNFsP
IYqx1AfexedAiane+APXm9HHuk4D5DYiWVYZUOnU/CHOidTwrxzPNlt8YnLRBOZe
VQC3WRxQDyQ4lNpag9bDeeVhXLRvBu5V0l6XbJrZq6+xZ5DQh7j4MHtG2lxWDCUR
4aQiv1hki1Nb+hULZh9BLlVPcaQWH9ygPGSDhRneX7qSVZ+MSVRbYhWS8r029B/1
na5EbsSO7O7tD41btDtceILYSBrqO59CyUDOhyQ/cy9fUIiEDRIUB4gZXaST5w87
Z7DUHkuMaioIm4g7ngldt/HTTLwtPxZVewnHZ0dmcTZhJzSS2z4C4Ptw5IAoMVj0
pNUii2Ch04umCz2kUIafJAUsnO+BY9wKxp7vCqaWS/j/zgTIX5E2ngPSZkzdAMxh
SMHrNQN5qOwp/1EUv/5vHSxcaGqOCf3YzBgLPSK0i9BgKRdHTK6wQ+J8xnLgqFkm
UzMSHFC4V981acB/HhGtPmJ0RnheVJhx4jCj6nCSviQbo0NWsPPa97haUseblPKx
A13w1PkQ+xMUPCRLLuvtCs7uM+IMM84wX4ltpbTmSIsq37UTrhuPONRtyY4xiHhT
cS0u7e7Wz0iI9vEwzO/LTNpRDYdRXSydlzpZCHqHWls6gbJFjt7nBtBtUCOjSUZB
T+EghGG3asMS+voxxZR2k8bfXTW8zvMVUnH9g3dEDWeBqh2wcWly7d96wWMqpppY
tY43ao8S+pVR0ysoFRP3UhqV0KCjpWjAkl06r2yh8DVmy5Q1/yWhk+8hPq8PfM7/
A7U9e3umV2nOY4uitLTV4RvgY/xH6ORi8G124HiQLBUZXW7k+a2E2qkWw2dGCEa3
1fI0OJ5nEuO4HRxn7wHoiDzz2PJCEpleAm7If/cKMBvGWJIObviUZptWWYVZT++x
wofuJB1owip0u2Lg6/cX0NeIW0kQHvf2Cp9xh0SI6EL8w54orLCoGnfyBxEa69Zx
B8Wx6Q3sLa1QfRD3Y7fPk0NFdDGx3tDi2pgwW+9FTifDVTKm+Uz+BWE8/P/cPk/D
DZuiclB60a3EPpX6hSzNB4crcvlZbz7bv86Y5sDIAxckcRar/KneYs89SRgw2jeb
DUeQQldlSbAuZM+TvR10DTfYkLqmlDOJDWOtu8Cs0BPI7S67OvBTe1bWPzODchwy
N+tuOl8UcTJ/KtpKSVq3e3CEPcOb8Hg5yrs4HLWuNArMvadcr6q7CmSVjj+NOnk2
CC2jJV02Uf/ScckhiPrKlwanmfGjjMl83PkteKZH+6iH67sFBzPHvSC3e9+nSduK
TneOB5TpXp4aax1wouKkZI4PrTjWK3thew0+u7zQLqHukVU8BFeYSFsw3DgppVGh
kHIRoryDrVkOy17pTafFFvIq5Y+4VWayIBYkfukXTg8fhNTSGtTEwx/oQJCrKiFk
3k1dss6M7Dt+FvH4ut8JWi/AULz3wWA23Y7osawqda9XRtem+KJ2UciP+3CPkwUh
5hEqjsC3TqTsW24X2TEHSLtUZ9keH7fJIucM9zDXt8dFB63N+7uuh5BPuew4tFcM
PgvijhWv6ymquvdvvzGaF98oRgn7mZitDTkcxI03QBI8tBNzt5JdXe612LJqMMLz
CNANqkRDFAAiV8QIJoXxYJ0ut9zV9gq/G8YJKBkK0PtsRZDm0hqfXvADDOnncoca
g1mUXrYnCUN3hMrjClGjbjWWFR0kp9xyU/q+yNj/Rua/3J0w4TrewCmAH2tBEEYx
xkiSZaRatkJU656CZTqal4LgCsvJVVKsPa1kXpwdM9TtFal1J71t+4Gxi7bttjrZ
a0vpxu1kF3aczd8VHsqkyHIBkvx6Dk2A5p6k8vHXD4kek5TD2eD/r+4Rbt5V9RkU
OYUElFMCxMRyTlcUCgu+27b+0hM+EVBmVv6XTPAUS392QIev+qIoXjP+F86okGMc
/tO33cye1V3TmVO8F7fbDnW8prN8G4n2oA5U4yoPbE4GcgAATUGSMoaeNpewoiCs
fuDDD5+relO8A0rAL5fexS8NKtkSRZiNrjlU62ogL7qhjF3mLjH8SQK39iY53dvu
XgPxFh3+37yC6iGiL5qAV+OlxRIxZGNlmzuHvh1bmQjr5cN8lSJ/BIdN3MvRvFOK
X4JI7KRsfpzreJc2iO3kfDkvDipTSNm4ldoiBwl8/vk7V8n4zSgzwoB5VGTz+q+H
g+xjkcIzuWYag5CUOxuMvzqrChmcX1UtkdVz4eNz7TJja8ypyjaeu/xVrvkljkzs
A+l86jLCTn68vPhQT4EgH2Pr9GTN0dRS2l+C7zvs6624cipe9OV/8rPZj2huFwJ/
mfQp4uu7Ke0oD+zfRuAq5Kaas/DHnPbxlyC5fxzxnQGsYjm72BqKHcYIFnWNWNsp
3ILDewyTt8X32+kowPr1iWJSAx8r5M9VnhESSAAM7YFQZ4GHXMNfIH2yx9kPRgDC
jhhfOlcQKGzSgnvH2G2OAoNOElZfWQ/h50vIouaILcd+w0xeYa/lvU70f3/ybbsC
/76luAbYpiXWF0X0vVi+zJ5DP1OxHpqb+p3ctOxmWaGAFhZVjprjSYMJSO87+HTy
6YMvqd/9OJeJlf66mYePlyDI1EoJ5q+wmMEnEH8IiR5uu8m3epX0hc9qxv9r+5Np
HRx21seklqmlkBQBBg+tABEqfa6aJbG+mjRSc1jbAueK6h4+okoB76thSBD4Z5qG
XX09ribMoeOrX2QgD6oT/a552g0hpWlVgFAjs08pvNfcT5ErWdfe2+mFQSG3DYbE
UQ1CnygScpRwIkd8K82bvFK2YP5MfA7VqyaVK0bJ3ZFK+UGkk55baiIhz0K4dILc
KIOGgZfFSqZi+HXd70RDcMo3EjZ+ZR8ChS71Q/7Jy6iXoL5o/4RRhJWOoM6zVIj1
d4yQoQV/nWBqaxnqRvr7znPvwFJkUmAKcbwbUnu8hfoH8eV2sm2byq28uCovrJ49
qqgE3e7HuBcU5E3lqE7VfpYz3Y9wgMi1J02hRH24jtP63rxd7yfJIBJWjWdtvFny
Hy0LMtLi3GZ44jVV0OtMuP5EfzyZMvEnIo78mKZ65w1vAWInloDXpsVqJiuk4Zd4
bthyureYuzKAjP+MovUyoZPuveBPXihYFlHw4/zFJi1stDXjWSBIeEevp+XalChX
tZ8Ig3Gx97z3+jO+DG0xOrmRPA5+RizoZC52EyRhFmmPjm6vQ7Ljb2Wf7B4XXDh1
Y25vYkWyjRi5+V06QZAPg7KA6Ew2LeWU7Np4czeGhjyjy6BWCvvWCneTO3BpTT59
EZedQQHTu+52kmxS0suHJDfcAcqJ+o29atuV5/bYJ8deJzxnRwmlCv8j9Z5jixy5
txcAGgVKRb2FzvW1etg2gokHl+VWT/0UCIQx84Q4+Dv8VCrZR6D9R+TiljWdGWGc
VaI+LZZoY05/LJu6NOyjNU8rXtrBIHw5mMUpJqrPxgdWtvCyd3M6kUz4FR1ROvW+
/0f2FcR0SQl9Hl+z7CxblfKYKyVZPsuJhkZATN4pQ8xvz8NcZippi+j+ktyqirNh
Q4FUBbfravOlv65iiwK9Jt1OUy57fswwJTLhAIcxXNGu1fOXpvyHyooXGFg7Hb7E
17JiKS2CuTZEcZ3VkATIZqhkPEiari46Cbr4IAzaVMb5NySL3g0b4P+nexL142ut
/sXrl8zomLLNlAPhCsT5BP4IVTFD1+LuDNZinn5/j/zIj9s1LFi93HjFLAVK3mD7
A1+frWsQC83ynoOSDvjQ6yCeqdBkOtLevpZyzx/MraYK+G7yNleb+KMoxA1BD7Et
3wZEdOhs3s1JcRYsluBPQxoNLPNDUYlYQbSx7xG0VPfwe0140PXxjc5TYOtetamE
Ml3qFtUZothuJ+KxiaZ0fvDT6KoXdgcyrHkf8DyCJiJMhTEI0amwWg8hkGQ7WBdg
hH5K9ZP4KqjfTnjV09LYW+8ZjKU6K4gF98lPiIdXeA5eZKdyYgRjnpnU1se/cxW+
GtuQPOG9kEZzoeZZMAzRmCGKrqzYpwJ86Z7aXYvABf9yUw2k+5jGJR6/TDQd5wkN
Q3EIyAplrFU8hst41RNPrdwxI6w3DISdZwZ+4o6vEqqTEAz3l1mL/tMTJENpbjvg
n2EOVIMZuzbaLFzP3vpy84ozMO33hPL/XdgszFQuAq6DOY1VC/uTMvQOWsLhT39R
KfwuAhmtKbBqd2uIykOtThBbHHXpG483buYyj8PhJxucm5Mi5SgDq9orXMLhu7vF
Uq/1WIjD+n5jNGKQI38x9D6DIcsL6SdW25+c0gzFEpCRP101QjxV36pdM7hceMeZ
39o/bvjN8VnhOTraNioD8i3mc+c3MBcGnpmpsms8Y88F8lBKRN+DX+Vhbp2fEeDI
rddnfdrrJz8E6kNcIHiXnlgTRufabCrvIOli0QvX2emgoq+GDHLiEVaDZSD6bSm1
KHcu456mMKfYqqgjfxCB3fI/34y9H1Y0oxMINeByp3AJtIfLXTzEHmd2kFevfhry
7f3U/Z6dU+eSQSTA2MYt9OiCipowgHdHQ9V4AKkbBWImyTO5C5CouIi5qY7CK7Hv
1J/QMm6Rr/DtSWS4fIYTT5mnJ29qH5napyziienk+hOSpNRJSBFXQFTC/V6h2ip4
FnCc/Pmp47ugs/5THIX7Ma5hpbL2JMYB1gaH3BhJwg2nL9qMvXszy4JMYJHbPIVo
Q1mZOp/ttBoC/uTHVNCyZDSwehU0ZKEvzXM6b0KTCbMmcKnBIdYno5DFgyzeHwUO
uy1DeX92WhQ4uORKJrPVa2Rs5cFDBQcbe9JtbXU5MbwOa5VFwu+ulU+8STC2JNdD
zzXvQPZILrI4+jxiJCnNFnO/WYprf+J2nN/ojhInePGQi+tXvUwseNi5HG5xGNiC
s6BFcODB8Sz9+MvrRAJMDcDhR5e7P0vckbaKPqCBmCuQZYnJOAi4dROMGBMXpxdg
EB5JTCew+N9ORlOMRQoeQ1rCEXEwjzn9tQFJGLAtf4mg0B0YZzzE4q8UlQ5qLA/i
+WCNhdPeOQZOmrl8oxR7iFVuEOTp9b8Pm8R3YL18O/H5R+s7ytsOBT7+CCox+7Sg
j1jDIOUsBVQkqzpNhDlQmmAWZjKq14wFtvlIHY4aQT9nS4TL+RuAiUzS3+3Kv+n1
FS6em5QiPLJLeP6+jdsUhBtV2uBoDl+00OaMdfgXApxbNyb8DclgwBNHbTJyisga
Ym8Hs90djm+vd1MkdyHorq0teR7sktZgSw7y2FJyavjoRpJCscjYja5+3wd6Kih/
RtTOFglYAfLxoyWNepwbK99Yre4Dhafnk2AmxOSCsvWMAsymMte9pkbcW2TC6yyM
DTskZjQMaLWfEGVzokxIxedyxJOLZtWm33JqrnqfXRLWZfafldSdYvgUnAnOOy6s
S4UA301BkoF+tk/DKxf+0hfdHttJy9LkvRns8sVsJJcxDJ8bpD+TkzEzuRBJEDdf
x3xqlDYltWRMX0EBUQyUud78QdONuiSlceI6IucOkAGFiP6wFF0MNUNdUY/knBh1
QoYjd65UlRCrz9WGFtUkcEth2gw/t5LOMU/o9RVaGYASE4hqFJzHUa+MdYV4dnBf
DqL5NRE9hhp7I98l1Mz5u7s8/+SFyjJzBOX9Q9xaMpMPj3qGazMb1j/rgoCqc+pA
2Io9750qDEDcfiAnn2kAbZ4qeNky1U47tS32IY5OnOVVAahZUCs9GblQ40oJl/jW
DB+vH7rTP6OG4XLTVsb+FRh1a6SBbwOVtEASSyHppo7+dErmxOEAc5C60RSMTtYy
mO1nhN+Fdn50PBvH1unTBL+YjZC6WUde8xKkNrMCR83/qM8Pz2BJCy3Mituuybh7
QGti6/gk1gGi0iUdPNd3ueeRoOL1Vm/zQxqWApzUjtZDRUEuDXBMkqN1+W2v/HEm
AJc9+EKz+sJLXa6Rh31sAUvkwTYhZrijReiQuMW9mMbwRUySYRetFKR5INYV2+7V
6oi20IBo89n+uwnsxqVhpmCBU6Pi3XgP8LylRDtK+CLNUpK8662WfhlPWy2REaQj
xpSRszL8zpXYW9aS7a0lbUtz4kTpVxn+UpY2P08PuBl4jLmHK4FXTwNT7G8XdCq7
wCWj9yd5pnTUlwlsecTbFdoLpCP818dta8eEHK/sqZdC4vKC6xgkSId+IRuUXE0B
w56Bm6WjwWyyNq0sFYiEurc8qhgnOx0gFvLRdhdFVxTCMuXxz3BVDVoJuhpa/RIc
EHtdhG6W3/rTlgnU91FJFTPsKk402otY3ybbIZKg/C0xDYq0M0Yr0fObhBIsLe7R
NGo9Mk2a7c4GMRjso1NsxWZ+tSLhYq5wxnl4LVznzKxMLDlZ9Sh70YYeF2WxFatw
YrqZKl2fM8qZuAjDIQlXZJ8b/QbgFvDEIbbooRBRumUxQXJ5iwj3Rxz+8zDqU3cU
q6nR9u4NW+12JryPFh3KVEvXFVCPDX2nxQ1h+iwxUhTIwK4aZGmW6Ms11+JMU6Wm
eQu80ZB/GEl50Bm2FkRKz2bC8f9ZKv4l8LDSBCMKFHM9FLwcJ00uX0Xk/zUNTDhD
pFf7wwkZAme0kdB2zcT+Ovg85CotW6edtmYxp2OucCNAT3K0Kc+3BviXp8LIqRMv
KhHzf2gMuHNUn3jJ6dbJ/BvWqVcdMs7z3k5lxQmbzynrlBHMwXkdVeL4nhmj1ufv
GeqFnOXNCm5Q4fw6j6DiRLl20YIKdoxOisBiVztivuuVb4TyvYwMBIiqXoiE+2hn
jNtvj2CvrRUUhrXRAdwzNenG+1J4+xOIQL+NUhqU1NezPaxFGgjF/jCnMkYO5/+P
F3ryGG8Da/OUG0vvRQbraspsH7yjbag4B+05tIIkVo+48WkdeOHoD8G9JwecE7/0
+1aXnSqy8uFpkMzBa34IVEwzs19wp82bOs+Lkzf4kRgzLcf/1i6Bt0M4K4aQVPMA
29z4VXpraRJNTol5Ko6q00QrSjLd0ZonQ5jJx4yySMmTpVZN+bA2u8JzYs+MA9g6
muLp8zF6WXF2ulCOBXjPNlF6VvJ3UBxXmGzExlfLGUZig15XkyO/aGzdVEsjvEK4
Mrv69KRnefmlAWN8sGhiCo7ivUhbUlmooKx/mA/whRQEkWWdGGldb87W2VRaAWsH
Za1mJAQVoNFzGb0YutF3+sJJ/Y2+JYGajcRLYG2ddkOmfq9VXozL1Dmv8uy/ZmBs
eXFZMFpRfWit34cmyHXAieKAEKeP9D7Jg4M0FxttDxaoOe5kGScKgN1iG4zE/+L4
lb7OjnCcAQgo+AasxsVOY5/7fDAd3srDd+QyHjiaaoyn8AOvjMiINpFu5OnSu99y
SnNoTzRQcBsErq7/g/z6YqTmyAC1aqTb4Fy0Mfl1hhyZFg7RkuZQMw6F8Tj7Ha1+
cAJk4DsNT1gsUz64O0q8eXJHSmT0BrUnnr6aLsxZX9MUwPgfZgSvvLDPEJatLsjQ
A1lNzd9LCHxgrTjt4NcMrijESFeWLLagLdN0MDn6Hak/tgB9GMdlPgkqzyYF6RF4
eIPyfuuz72LwgRQrFzTKzy9ADWM4tZG5Wis3+6HIanxK7K8yDjiMh2rGVIdmAGaN
XcIt4kzqL6UHrs8udow9yefrAbQV1tVwacUnS43Miz8cW+n2/c5uRCN4SUX1e4Fg
9X7bOEsUccV7s9eQG+1U+QrRTnAhDACLhTcTghcVlCs7vfY+G730DJdZYN8P5mej
1RRdILuknnd22HlbyL6QUbp3hxg7RM5YnOzRLrrqQnbAA37C45prDwY0+oD+ap/I
wX2z+9rZ5c2I8RiwxGylggc9lrbLPnXWmr89YOE2HI+npSIm5TXbI6G4SmhGPmqG
eb5XxQwAQKH4HWjW98bWqptwYS7LbgMyu3dkBEnlHD/iTV5q242LmHvGWKYzgKfo
6dawK/e6jJZEItRRfXMPwwTQ8rFBnVrmRD1NSehXssqf49OLQo61eaKVknxROpg/
2yji/nwKXfoCZ21SuVhQ5C+tCesPxUSUsrTGTQQAU+fxKRidqiJ+xcni0InExTWc
uC4Ojy3MlGX2ggE6+aQrRIJRKNzCBzOwy59f40cpOGY8CBjlyXCbYxT4EmwFEM+8
8ykyIakey/rtoHoldDZ0sSy8+B8CRgCpcEhD/QqZC4Kewo8gIGbB2Q7Fk9001zGM
t/0l7MHGbfE5PAsjmYV9L6oVEUurXIhmqyj53W8tpqgfIh3I2UTa6p4f6TUgwipG
lXr+clVtlqK9cLnwSd5m5gQdh7LwmTFupevsnmiX48qdID2J/ODzSjVWANRfew35
VMwGZOXlsIY407gIUpGxBfSKZ9GnrQnzYeW32Ma+L+wi6GnSERbS1WawwuDFPw4q
C74wOMhzR83zlK8VdaNaCp/gN0RRIikn9OBxemNj825kfcH+B2gsBTsR+aD6YkrH
raJ/q5R3xUg7sINtQgTq1/z7SAzhSa3YTlQU9OqfgeXr2Iqdmz9qRfOI82+vnn4y
4S3jUqmZq2k+nr83bywC/FWbtnzNcvgaEAv79RpgqMgQVXNlVVYYESLGE6SvKs3o
ebAgTYXIySyAw2vA8gcPlDinqkwcqEuOfZowYbU+95UQU7uKj38CRhAklrMBzGhi
2zgd48nQ6bpAQc5vjsLB4U/IgfH4uHO3NdBtEvxSyPkAImJw5KxQvPfPCfN04W3q
nbnXfCIDp1HXkXpsIaSKjrP3JckP1/I1FeNrxvbgTSCa9bZ8sv9FXW7bCRScMHb1
BB1+XRpTIU7mnKNkgbf02wlK8ZxnHTH2ZtoJST1BPrEVUkxSwWh9Ba4ovL0KqI8D
b1lOjAUxieFUdAWHSda+hhou6WIhUUO2zetv18/FXsm8Hz5TU1xu33AzMSXDlLC7
WgOLV2JPf3JuJ33LS5Lw92h6cibobgHRwv81FPaAeOzm/FwbfGhP9zB929c/71eL
8Zuhn3kxpFvtcosbQpGNNnOwasy7k32aiXQKWvsyLkMUirMK4Cs0NBcdm00HvJFm
3Hn9ddhkKAd7xc6vpczbFDLDOBqWUzA+tcPu1jpWRybhD0P7VVIvbOGFzGQP0r3G
zUj6MGa6QYHPr7Avvcg9w1KaH/O3WFIV6lGt9FLxleb7KoNTxQm2HgekkC7HZ/aI
eXrUBa+R6Mp5IcB0gqxoWTVzi3YSk4SGSXgSo4vKM+laq+Prdrrjcl1+Le1AJAfI
RU8f0muNrY3dPf8DcvErV47WpAMI40n3XeHvQdXO/4WkypKvAdeU4CfzKCB9zUOv
Jei7ug48qJ6blZ48cVAuWnhWJhBEk8gWKb2A0/vHs1K9QCkhIl2eX9C3+XP1znsa
44bGJkQvC95T2yw5K+QnbUKITCyzVogInUMA8LgACUeUEJjR3GhHRBRCwCUakMOB
Qx+npdGlExIE21Mkuv9efLb6y6VR2ofIGlWP83WKKQZg664jsJyuYjLdSRke7TJt
Yf3uzfR4tpQsZU4S5bRsoSQgfMYR+6IBRMROrOwaCmWYonlNRbi2Dl6XNNLvHbjx
uYMUTVwRV3OjMm1VOP/VTigBc9E9ECDoaftue3uIv6yjg1WW9BU0wZM1sp2twYnB
QYugZmhTFQkD4fpdwI7e9bzfDZak19VvPgSX51i556A6F2iTQ/CyFi775EZSpbuY
Bb9kmBSBmQZoJlUsTAD7idVqkALWOkH3YEn1iRBXJ94f9IR3V9FXU35KQfw1EKH0
Bry3pJPb3Gafbiocv5neHt8Gd6KWuve+KsLTARJECgWHV9Y30bYPLFHmKb+cJGFJ
tMovB/XBpd2JHsBPe9pqpjt96A8qqXnPZ638MmLrDEsAieh9Bq9YyxjTgpllIXeb
FkQK3tePkwOi2mOInhgVbW8NiYbcDMs24Lu2PD5ZYTEnKLxisglLL95/pd/WlRH1
67w+5UFBmpBUkFH4MYoEKM94Zqc7wHc8xGLZEYO/Vj/cw4gc70uNSDrjIJq0ekzk
ZY2umIBEUBm6SLdOxmwCEQZzQ0ol9PO0WKz/ksF+eIRCAgECImPDAAGxzFSg2Txv
BcXnOSEICaxC97Rg+pLpiEXl9XF3sWKm0IJkxoQvJ0u6aS5/p2t4BAVQ98iQIPR0
iCVicHdXNqih+2tSyX2WR31w4lGcjMMQE7rhMHV7gDLHBzFNox4J+xySChBS86KE
X2Vx+00dowGPIMn815lmpbaN43gm0Z7HQGiIUBf4Ik7uZPoquMFRTr1+6Xg6M+b7
IyvSwPkPQlEAkZ/8aMYpZoQvb8yfN/NHsP72ayuswCoJxq2kFTdePLzbBPvUc7dE
llNzR1/C3yA46BDfq5mdir+IFF5NyXmcW7mQb3WVh8kCQV6RrS8XLuKC28kY0FMS
K+moZ/AmsYodFsn/zrTjRwNNamfgfSuic1feIboOmiYRZO9wVrRt38cP2H3b8KeQ
E4bPUsA12NVBuf8dQ8Rq1qn5oYPRJuCKuPyqNJAV/BPF53C/ZbSGEToAblWTQw0f
InXDD3DGWnCZL5883ECqUJRC6XTVa9PIlJyMjud+XKStIsXsj4pCDinGaghTFg84
bfZloGUjsDk0RE7NhPGqahcRct01EHZYeFtPj+hauauSKfbtUadslGwM8IYgAL38
O0SRqStxFwgaXv62PU8B9fnd4XQA9EVXBAhZYm8ZcRnOl37J5EHwTg2g1Fa9W2oD
cm1EtUxZPr18n59ZdL1ysKsq1TyITAVyiSNv+Vchz91QDS9CPFrgknuVgPQb+A2/
zr27GYGe5sCbQlWYkO/ckpGHehP25ZWfWmjknV4BxsX3ezPpbCkslfXZYv0HR5Gz
dtlPkZAIdED7nHmMC661I1/dwJvOf/OHpLEwTLYLu8HBszQuObmO7iDl9c3Yx2Zt
YmpI7+xXywG6FVjWwrFydf21ynTWrFtyRxPiqUdLMGk9dAGRO7HkNppFssWM6iAq
9cGRAauq7yFSDHs1mZFYW0Ob/AcgA42XPV/r09USX+v+27Ym+fHD87kzDqPuG5Fh
ecfmBawYzVThlcZhDZJ+oNNdGWKw38AatPtom8fHsI1FxmjB3DYTTkCxjyOrQq2p
MFwqHgDAZalA2ezi1N6ppmuLBV7K/Z+uNOp9G1/nQsg4fGA76yvi4qTle6Ba3+Df
OxbhZb7csLl3ba8cY+4VNqHJe6sN/p5gs41Y7lp6/Crho9naGqdlF+j41Y14GLd/
3F/baKem0Y+Y1ptWtMUp5N0IE7YOdo/lty4TvKSTDDKxMrF5v/8mUZhOsdO3cIzl
y1ywsifjuFqmKYJiXRLhMv0LNzSL3TJv4ne7oKFrMRFsyiFv1yWixMRYcc6/9xFY
AX+psDmG0/iZQ9BLU4VsvSVmkGzILMo+Q+2dO6nDOyN1PZhznnX8d3A53fjUiC3h
8qk5kwvNvq6btL/ZtrcooAeqPemq5jnSXC7zlyFyUofnksoUlb+usUb4XJMgiJMx
PzbAwB+Ycqd74l1bRRDlJyqC8iMM/q0pvf3qJqp6YuJGI6izLzeO7wYSe6XR9mrQ
fTybMXYLt4yx5Uir5f05NhB05elNLqsUB8Y/fb3wMghNLgp5/VBc5h3vhTSeHhs6
mvYkc4PDQ0F47zVpr2u/Q0cHPeSZiJXhNArgvj+eKqHT3ns+gpDq8pPZM27TYb4W
Nngr3oxqLLCtGjM/IN7iBgRkLYt3FELG8myaoArTKi/uzYVESOvNmiESnjI1nQ7Y
i/T0ScsFoYYxiLS+N6pma9+GcEYxyRNa1ZLF4mj6w0+AI1lUDfuXcnECe6ayDoFn
pQYyVZMYx5mecVK5AjYDjWyy4o4BgAZT5hLHo11IkrEeApvduJwfUz8Js0sQwquE
L7WYgrZ7rjLTAMBx0hGjZDE7bRHQnyPo/POyQd/X4YvUvyrZVFzz4cFMjNKq6uDn
n/0ezLS1db7qEKYfPb11sRJ9XDRSszI5TpHAhYLQrUbGb9RtePplVbryeZInUDvi
dbLsJ3PaJmiyxaoqwKTQLt4J9OFKDK3fZDOrvjzSCKLWC0a2AYjVMT7N7bsgDWIo
LZMbaqFoJjMQ2r28ESmQVjdX29FIw6aGYPd/uJkCXPpV3Al/rzt68dfsyEVndQi7
0M/5v1qM+V8AltXV56Z3X2x8Z4DlUINtHUfmv920aJGjhEfSJu5DcXENefy25xTI
7SXvoLTNcIXRAU+LeL8kc2Uku4QaGtZ3joQUZ5qYg+g2y+BdddMSe9PunTMrkqga
QvK833FjArsVCrKbGRCO6SGs5y4nYhzVMBhQO8iAiPhFSe+1m6HgpY8DZc5uVpum
VBGJPQExDvvS3OWDXK03Msl5tPBct2LpZOszXC7F5HCbEcJGPOx3Rwj7ImgOMwzE
zV+Pyh87RmQUQ6xcLXJNG6UH+L/q2X8sl2jt0Dl8S0RrgNjO0PycOQMMhuYTyma9
m+GXkJxbEOg6icj4DrVk590jpr5xNPHX7lYjJFm3WngFJ/ndq4wNndAMl4nYo9W4
gRREkv1eEXmRGtBTAnqLY524A7waf3gyR/JgTikj6v5oAyLcyFsnvDoadzw7Dhk0
MArSpO32wSmkE6G8S5eEH+tf387VS1mr6iy8Wu9+gRZQ+qt+peyODO6M/AJuHwbm
KZcKNO+k++3i+DYsAPHHbD02to9G9dkBksxvbPj9TV7KDn27qlPGVxfhzc/eurpm
/0oH8rlw5TOSns5pKpP5nRCKbV8sFR33uFAhsvYTTNAKI7sGcmsfAsFk3F+ioeAw
aWtuUyRrTusA68kEBbHXjZoz1bGUR2JiiPpCI6/UNVa16fqMPi0BYqcoej0SDyFO
HvwtX2rS39KzFmsjgdA+3zZHy2Z2HnLRu37ybeFUxg+ZjkC/21oHqDFw1JJqQexa
SE1GIvccR2+pVztA/UQJstOIVepHYWHFp6JMH170VPi4sMkIboxj1+nZc42/sROd
+OO/pz396A76DfLcA/r/y04Hgndr4ZpgVk2UaNi/ITuUSwfpoC/aseKT7y/KLigB
7uIW+JN0TX5AFFRmSjrcBmPPAjy4vl+IzNhGeFKTbAEB0mLXTNbNKPyhIN6g+GdC
bvdk+kk2FswMkfQklP59N3mfRhDuepkgdJC94VU4EVMXXKcaiv7KgMBM6sauPi+n
XAf3qOh2f2PqCayIzghTu/x7vBLr5MX2pZM72CxJikf73a6OVwa34GkvbwguVsVY
y8wz7YrU+zIavngTqbILgv4kM5o1P4xFKxOYfZJ/xgCIeHZCU3Qy1sZv4/I8aEvo
cEbxZXtpWJDZbjBl00tSyepqmhKncQhKqwvTv2v5PMcYUBtVaCt9BUBbgIwaWltI
XYz7naUZTUsj0O7371lBW24Bq3aFpObLIfCxjK5zCxsvuly1Kc+qwVDCLS3GH5v9
mAHnqAts8dL46Y67LAVVtZewLmq8QT3zvDG47La7Tj8Fvv+xHzJEeSYgyQ42pLI0
wQDhyIA+N4LzqbcO11IFQ21tB27F7zkjc4IwFJ+D6O8Jzzu/LhRA60vG/4I9Tqha
SOKA6++EzjB1N6Sw5KH6+qpLGSYdu+WusRazTJ28rOyEKgLXPMhF4xMMkqvs8Q0E
QTAVhHdZbNeI0E4d71rRoL1EdXQgQ4fboMpdeSSzj4iE4EGNz1i3xeS+l7y7v2q5
ICb4R5/I+n1U/T+ynSubGZzNVJ6wQci9TANxq+kRD3COuiaalY2CE3E052Ke5XkH
A6psgMFhKnsMhn59Ixf4gi/UPA3KqdjBmOfP5ZXW1lZJI3yKO5uEkhm4GcXtiB8c
PrF1dpckZQUj00hzfcZHxtNeThCMy7tQxHcMGRLqyU422Cyf1CBOj551ARUYlnKj
SfVmYf1qT7zaJKimsUOlJtBB2KHctHFDQxmNoIii/6ETaG9/AOsgAiz6lbj7D3cS
N3FU4oQbT3vbu9AVurt1di29/vfmIgqxhAZnULDcsQF4dhgAeNtUIFsm/2zjLCIq
/BkSQfQL3fkeapUNH/mXkzwr0c+iUiqF66tqZxz3GauSgmSGJDd8sO1Z+PEI0DcE
BC16XBgvD/uij3mIFN4tXMsgO2SaTVerox/OlstJLRCp7vInyJ5Hujv5jaSUVb3D
ltz+kXRiKY4xj4UMksIBdclqc6f4fqbWsUTk8DpXPTrM/DzZYzOSSk0zomGT5jRa
QvtcZluUuL+Q0Pz3YoCaojsMoTYIT/+EqrGeUOQvXpX/T80JjEHV73cKGw4Cb8C2
/H5dxg6OovDTZGY2PSrBD9Q4wX7rWb1KXmt8FLeqFMpj09n+Op71aSuAo1HRVA2j
GYtS4RXcY0Hk/MZwGTYgfqjktDVM19C6SxPrpKA/44dyDQt1HWaRJchNrYmHwwgu
mKSQJmvLb7JWS1K5B6swnyPak734ldkQunjyFvXF0B76avwOOIxjKCpazjZqHQF4
7jTm3D9ZfED/vcGAfPF1m9ZNQZ6kGNchA0XaDKYZJTxQNvC4JuD25Cmi8rt0xFK6
U3WDMwRKnbz3TOZx3Y2wNy6+unnyo0qA94rUpLj2PeovRsDzVRTKupiHFwYCuQqB
vXp7R/mKCgvci8U5BeM9fofnZsrp2y5mlZqM8vCGp3j7fJPjWg1JTWEhlqyHNXVD
eVX2oaCQNzEC+g46VTuyaPMGkuBkI5uVS86cAhbXHWI3KaF8cl0Gp8bm21kP/U5f
eN89NgWKNF441tpAIvKsuqM3OktBCwK568qridVjGVePlsQS0P+nu1mO1fJE9nrr
NbXx+hi9hxXQ0QC2Xv+dOIpLJLaxVBqFX5pUTBS9aWZhTOD9BGVH1qY8k7WGK7zZ
qw/60S0qYQjVAMXfISJ95aKcEqOwW8OPyC99Bo5zQjr83oQNtGGHcP9juAD2/SiN
XlAeJW9fbkHHklnzfv2iVlur3A6es1uRtr0fL+bTWmlUE7V8+YArw+/wM8eePFsi
aA0/zkNWi1HFm9oUY9AUGv3apsNHrWuAmZMbqRB+bw0bmGx47TjXg6Nv7dIcRD5q
PmFs+uMGwG5CX54jAp1Ol+EH7NoXJH9DoTqnzuS2b4c7Q5BN79srK/OG4ulcr8dl
wmOluK7PkQ1IDrORG6n0qWuIJr3NNCc5zHevF9v3xuIXHuH20BUJvVfV7APLm6K/
IXG/p2Agme8hPM4lTUK52A4Qn1jW5aRDaYzv/LCwz3onHF35N7SRd6VXpd1Bv11G
hreu0M1FQZAyvPuZn7ODy9BU2CHn+YKu2TuDAmJ4yCU2FEa9fjfZsmw2sg3c65Di
dMUhK2RZj1avkd2T/rmJU51KkpC2SjduBSINxHrgC3R7lNGz/YQkYAyzlYcZ4nLj
S6Hl3iAp5ECFF+8Afras0Ve0X1umRJ36dVHQ6YCzDu9F7YHbdDSjlrvchBF4jSYa
izURw9NOlQOtUHYllB57b+Md2I0a/76w4hjVuwq0ckDQScn9TKNiSqzmKwAT89uq
0fiQBcJ5+48kB8IbHpikeo/4xlTUia8+VNg/JRaXuZrXLczkyIqAvWT+UYdHad6U
RWj4konkKigBTbSu66g/VZc7THo1DEVwqJJxO741MsZQJAoPFigrJw2HRaq/Nynu
5vS5SyBEXyzzlYKJq99AP7zyYtecuSEzIDi/v/dZ5o+eEGYewtKk9/iOTKKxh+cb
qKpFOsIpqP1+N3yaPq1VdAsx5eIDhDXjtjPwEFWKx3iA1Awvy22RHLll2Fx22MUW
DHc2rvkOjQzq+d73FGk+CyfOlJcA14m7fAqEWw5CxNctPNI0VmxI8A4JiNR9Zx3y
DhqhaW4dGHomnmbV6kjHznTFpZlEPA9R/YC7MJtbXjEuCHot2DKnGuYwXQCcwoZp
IUCzmhQsLovcEyD/p29my/UaM6ndwaCl0UO/B7Ma56fujvAKXvu1ghKOzPF8jI9l
3sESgI5ew4DYV3GB/e2Zt7n5AU1AqLQj2okKEIsxngit1TAhM80gPpFxMbThWp5K
W2IaF228jIuju9mU8if7TxZjjYSfn0RVjxXKTEaTpppSNdxbS4VWiFnsxka3X9t/
Ru7t8QE/CkPk7XgdxYzJ55Te8suTsbKToe6619u+JMOMa2Ouh91G/jpx3JgJx8gw
aLa58rxqPr76diVfHbctu1Jj++gHyDhq4WzAFtWQU574HiPAH3b7Y4+pEMJOIVNC
YHiK4+YLcbFva+yShsB7VHXFCUhVjZ/V9upN9HPWOBkfvzLpHRhNg0ADUzJa9htp
s+0e+BUlHD27ak4d6RM6KjXH/Khopn5cUzsvBavyHBXWqc1Ke9ohH1+/Kjk2m9fU
KCxCTnANlZ1F/nAmuq7HRnR3jdh0vcXaAsidGeH5nNoopV2N7bMzeshdt73czCAL
bVMT3EiTIO2YNM0qNu3xOS9a9fRq1peP+yOiTmMRftGq69DOCjl9vngFpXxz5oBD
8Plgj/hUgloamu75hemfFGPaBV9RJ6hdfj1fu1tILg/Z3sR0L5xp92k5zHuFzLsF
9a+v5QJ1dWheZxxrzvrEzX0bGbmPeVpOb6Jd1FcP2x7ZTOsBHeK2s5iVFWP9Mjy/
yZjN3LCdmI1DD0aIxIykFGOj2XPNh6KJ3XNOBJT0TvM0JBLFAeoOjNxRjXqdmB2r
nBgohvOchC+oxcBqwroLkvnp885NUM9HihkUPHOjrmLQGWo4iMZYJtGIuWSYrISD
+NTdXim8CGTvicqQqg3x+MnftUYnERMGtNE3pW0y0EUSa8FNzmqvC/qYr4g1gWPU
p4oZBrT6ssdxN7lnDiOfGIuzc7pU27R+1trSdAdUMRaV4KEn17hDMaPhz35NRYOY
jo7MDNK4XV2C8GSnthtWlRxxq6roX3ZaUAZPnmRLNn+jvaKsNPERqffsIMOO5Oxg
jL5qHkYzL0eTqIFJhKYBLamVEP9z2ZsQ+tprm+DYHIsDzpiPFfqOWSlZE1mleRCB
/IESmPpDbyRKktyoPxFswlx99lyGmm6H2Mm36g/w94oaGFiO+v0Kp9tNG2fnrFJI
gOP7X0CNVomTC1hnR7cm4qUqhTwmal3GQZ0V4T++wIOQKSXMsaDai+jYPCu6y+Yl
UhfzjzLRhxFAMif7AJair6ISdSYVZd8tmig/ymv00Tmdj/9SEsGsDt+azPJnLnyH
L5KJz/s5wImkUBhhndM9p9AYcFNbNkN5eLalJy+QgF9VEdpN+iHtMnbDFb/J3Kjx
s41K/MCGL2AcxouKSF/BZ7ZnblxzTt4fk0/pGxToH/cwWnU0jyHBlxyf3CnBRcQe
PW3Mbjdt3fUEB+l0Yg2X1NQ0WiwzS/yaPDUT+h8z/CP2DUthMAZlENZ+SrIonTXi
tW6wbf33d2jZgGgnZDdkyM9cV/DwNphaMBaEH6ukWIi16b1egMZnx1eluauOTED3
1r8gQI/syT4Byp25/0cpZyYYP5RDfhlxC98wrYqLuZARWZNWi+rs4r/kbCP0b1+B
m1GQ4DGvs/j1RjKijrypxxRN05GjtNt9/mAB6vx9Q/2b1IfdqLUOJ1AtEKWGXRd/
f1YrBdRnsizOeT8vRwftR0uei+UpXYmTQ5CNH8mXzvJAZbgZaM7PvuA0doShzIps
/8DEWnFXXqi3IhvEOVhhInLc079njA5r26wxGvWPklEL4dGilMk79cMt8kku4ae3
nt4nvgxlYhy24lfng/6Wrym6M1b+DquWnQGaUbo1GkdQxyFvL2LinZ+mplBhK7lN
xNoAyqgLNQ2arytTpnSRHI+Mrb49aQ2DcANtwR+Ni5fJSCPCbbVJ8bqyXGNxrutJ
nTlwy7ug1hOSO90ynbOWhmMKdyw8tJCnNyf5sAruEQRnztUpKMrhDjMiwmtfyJ5K
5RQikiIYDB45OEITDF7dvzYAfqQymIwCrr5FLXa03XbaqXkHLOj9T5qXTw+REloi
TQolbj2aXk2vFnZSCcOQLAO/vP5lJkcDZsfj9zsgv8BFWcskF688IMQ7uiEKwxqr
INZS/thWxd0RAQSOBQMg5LI858yPaefC1F+Gjl/vN2LOUsB8N4NERCbHhRMtedWT
mb3NFXnNM4AuRY0yRh44O7ece5809jARy9prvZCQICoIfEI86gnuOactEklvKP/k
qXyuW9rimyE0EVuT38Bx4Zy0OPtzbRCK5S5MP3kWnyGJxPueTzIcsTKn20oGRiuk
7+y3A3uE7KGxoHIlHEwX6b+ZpXeqCh7uK4GtUvw7/pI77VXsEz3uvWgDV5LeTlDm
RFONB3AHDYjAq0fyyLr2tgELQIw+xvIIg8pb3G3oVfmKBZJ9Ue3d9g9Zq9l7QckE
1wEZTC0YuOLHXir9YMmRTEij33K12VeYfa4TmLLIG8iosMyxZfLsRF5ocsvkPAnD
hTWeUo4dJghYWF88s1vblcbeWecLtgfOuT815vKzxi/xJVyb8pxFNQ6xnwE1kdVS
7CYHbB4YU/roTUmuVg2Mevh0/LkDrdrTNj0/+q4IGOzBkd9n2oe2OykodYigLlRP
dZdtsHjrbPbzKgh8LwsTVL2Gb216ZVbNxthwgBchkxaMV6x31PQOT0L8qRp0zeok
X/09RH6qTl6vVv+eC54QA8VHykwsbxxObSiK029eEHiPkv6DVeRKIztltsMgADJK
SKxFpZhdPe10FdgZiROyig0hKPxn6EG1PqNzXNM61hHC7VYc/V8mvmGDyo7UL8+J
HhQACTOgJU6lThvWX7vOuxX1rvpWOtJP8j2UNVnxDBSVBY+A4lvyU/uVkw+qxWme
JVBhGYCjmHLQEjV8Jugq+kuZ1k1mexaAwhF6AtH3NtQQ1es0lZhpHSIFEOzu/Dar
OYIEyXPOOYvx6YvrY5J+N+h9Fn5ggTNkqjBjvPAE6KBMBNcDGpx3w6UM3e0s5Ih3
YFgufvGVclx8Aur3M+e0ogEcvIH0OAO4o0uGl+5lJcvY7OaczMnzxCSOf0kaWsUM
bn4av3czVdknt+AFioGJZl5TMIjCmK6dRpWVDxFOZdBaMO0XdjQWxyWFAlKK34AW
tVwY1eNPdx9Kxeg6NFTRg0MAlWQgcw50eNevdU81UzreJntSC3f8yOnbzvDC//sL
cF7uLPX7Ff02wh6hQ+zIfryoGm31a0uKQ2AJN3PYnR9Sw4rkVkn8djsNozs7jHLm
tu6hwKpsn5OyizgInNrG8WMr7hN00emLoceBR+HfeG95TL5NjBkqU2aX5gKDRZAs
zlV1nFG2vX+KFsf87l6/M1p8woD4mtUjaN0FCj8FZLVobqpUEAkMUbfyW0KqwqJm
RmcCaNkW9I1Cc6VGYeeF//+RIAePjuRp6o0ZUj+Trqi1mX8r6RVcUrhdycE+hpYs
207s/98wBVeM4166tA8/pP8vqswf5HKHGaWJmX9qCaxoCZqFOWapLO1Epdwd8wJC
2j/vQIpGgJz/0mkCPUGlTu12rmTxgoZdXGaE0S/B8Y2ktkPFq4jKkQa1yoqSd6c+
nBzkAbreGlXTCMoQtUqFY1XIPHFdRlKkoTsBVqaSFYYroYJZNz4FT5UsbOo5rPa6
nYk5AtkeVakb8xxb6BOdtoCZ28D7uuawcndIWeecZevl2QPGD/5nNikVk11egt1n
WqFTpaA59E/OUX5Azf3PRR95cEl/uYhfyNeQnURWjQ/eTTkQu5LBsI7A9hpJ6OJJ
W83x18p2suWs/tOrT+S++MlYbLdSiA/PE3DLQj0zYkOrK/oM/flLHPXFpWLu1dea
Q6Rro3voZ2qPXSHZRagIK1OBPV/JPiy+eW/b5yrfYMDePzjQTfgcGSDJZ2iudCae
m5HK07nPwEILU+9pz5Tn730A7K8sxQCC+YvE/R05II4J1aMNU2oKtgmax7xNr26Q
SfV97f+xSV+uXrdiJvgDOip7K9daxBXQtTaC4ySHd/4Vqjfvlmsn7IQVFovu4RMe
21rWqIRXfciLt7JOelr3N/wQ7+H6DIcwgvT9MXWprPR18a92D8hy98K0Zh314jml
C1s7hooLAw0zAAkETriTJRKqr5j94yFPQTM4cWAVsR69V629xIvYLEFtedZA95ey
s5K1CWZ8jByjW6D74MiUGsdEIai1s2SBG40VyL+zgAyW+vdfChSIeIkDFkTm7Glp
nsrlNZDCykNZ58Eov0E3PwyjCubt2P1pmp9qbsTRdwKmG7+ysg4hIHMvIRsdHA4r
ke8DQGEKbRPOKfZrWrz+GzbYo/9/L1DPtk2aGhGV4ovE1PwS7G3Grh+JTFkOuufx
0MLkVSRAi7bo/VregH0eDfFIXYL+WNmUE0fcZ5aNIftq5YETzxy2nNmzEYO6BmpV
Czawzu+phHx5ZGCSTrD7/iWjth0NLwfDDK4Gnn2vkSVMdPEQ8pD9HpTqXXyYcxTO
rCN6sHlnSIZcLynFb1l3Amc1rAMesgvbM9eXZmuW9GMN+e4W7T7iznL2KoGBiQEh
fra5tz0U9WfWbOiWKHdXuIu3Is/Pz+/mnZt2qPNQCRqLaOAv6t2+7jM+SE4FvsdT
ZelHT+LCcW186RzLm9A6p8qZ9Z+NTuxLaTHCSHujxAtSh7UQCq4uGr1crdIxki1h
xnjmL4SFEWUb6GeqAIhzczIyk1j0ASvWAkmTNUcy0ZIHQLxLCCwO2QtBflIf79iX
anhwwwcaeH4KbgJKsQLGdooo0f2y0HxxVXgYnwWVMTFYsxYwn3W49hnGC/PaMiSM
OqZ8P2wokDAP7pOO5mRivoXP6int0bJQvIkU1/Icgortg+vAKjHfzh06vVyVvvs1
xTPRlAt+k+eM33156zaXEcF3yTEF7XY3qrMuUKF1kgw+9FtRzeh47FDF/9qK8IQG
KrWhSsPS54Lw+VHBf65BbZOyvn3H+HC8NjBeUXn7pRyWOhDHlp5HlQYkWI2ww8+d
wVdGdl60eLzbh0IACOfA9fcdUkspI4+HNZa42VZ2hb2hrSxXabBpC/EFX96coraY
7InM2AxHFY9Rs5AqHvlS13PQ0Ur7ZqTyQ0D7E6WFWaPyWGr39vL5wZVyxKrvnTD7
Lh8KF86EKkYjOGyscrtcGras97giKr58kQVlXkx+ewgup6TrJ61/ZODJduW8xWTM
SVal0+AXqjd8eGBY2gaWNmW7WRUpWqGxBnl9sjI6kzaUzmOxLhJxGH8I0NjBjwI0
W8ODy4jcjTl1kaSmx1x0qSyQ27JD0/C4qH+o7gbHWIx/2UWKYOJWdpvYhuhtYU4r
F0vhemeh7pcPSbgICx5MgvxSSOo+wssBOcQD3aQVXFpwph7GYl3HvwaiKox9ugHq
yQGxbFClakrYluSgysmZ7n5dr5UNmKyueH1dX9YfPXOLlpWcsgxT7hCw1mjznfZP
JZ5teGxIK4R2Ik627RhhIK1mb6PfqPf8vEMpYX3MGgDuXj0WhNpbINLWgqBnLRD0
OzGmXvh+2LgIQSZS5o5Gd0H6jQZseJ7o17qIkk0rUAma2nCWB4hJvxy4iZbAGixK
hKtwM6rpE72Fymg6qzkNChyo5gGd0ozG9dIzFUdxjlFd4Y0+EZJq0VpXheCqGG8t
BRf/kJcKVj8KUxjbg6qqf0Br7vsrvEA27dq4VT3rS5PSYg2IgSAr/8xtSJEIsv8T
rUrv6f4F1R+jLPmxHDSqZg1OVXFeql43jzJWM8Nc7ovU/mJT7W6N6U8ICS5o3Olp
w930PVpHV88lcgxJXN78ng1swFrizVa6HO2cdF/Ri/EHC7nS9VQxQDxMT4lMK00d
7OZ12a500KxYG+07LNtCpDHv4AaPOQk9O8q7aa+oJvFBk8O4s4hOo1ieRi2ytnmV
Lw6LzAWuTZq0XnDJ7blLWkFkpN+LMDnrk9jgnDE3D6D105OcZjDZ4aLTBpLBvmfT
MnBO8v8pDiqm9nD+kFZsGtllpuJ+5gKoj3Y0LiYRyu874RTga8joG/1fcwn2e/ai
fxSNxjCehXoMw8RH8R/0xBJpLpvj+InUED8JlC7hGN3M0sJEL2+Wy2vnpeVzRv0V
7MSpCPAnoDs+jzdSm8IbFD4nHFHs0yToc9TYpGivlMubujJPk5URkfd4cswywU7F
tMF+62kzV/ees9Gp2I43XAvbbVY1+t6IWbBgL/ySZj4DjCHU04+b1+nWmml7qu2+
hrWvuoHCm5vuS0TnmPbwja4yAxUh3kg+JoUZ87y5JeLgZxjQlnNyBaH5J9LMuO9a
G+wkDe5MvDIz04udRRMst2RZ5XBxpeUNnhhn24DiKYdAUuPB29ZcWeXzonWWgBBV
JSG0BBJQ/+TyJOOX2XLF6koOxHJFg3RkIFICZb72OXvnVV7KC16EofChZypYUBgJ
kHZ4RJToDMjB8YMamoCYT+iBHKm1Rca82C/0GIphJ3X2JmADLlqJrhYoKY5MGrgh
7JtJ3idBHgO7nR2fFniqZZFyGGW7/tOwbrVrcgzH1p8nwmPbdKdBoZMo9zq+Hdjv
YwZvZwDAUOVkzxcSMYOD8jUu4dpu3Og+K6vFTIQs9Qu+ZhjgfeKIeLA/hzXkiDxj
ehAF74VMRUq4B0XgZWidU2+m2bLkUTxtqhgqzJ4h7HMqNi7NmEM15l2p0xY8bkmO
CVoZF9/f76b8g2zL5CCDPyZwkbSAe0FhD+f7yUUx7jhT6lmXQ+ECgNAfA1BTQT1i
UIYsTS2xXHBGDPm5oQlOcCs2rh0nefUk+fXBmwArsmQC/8/rmQzk+VVeJOiuU/dl
y67tlIrZ018K8fEIAQ12AiR0EHkssY44NG9jnxYfwosPnSSGq/AuHRF3j88Yhi6Z
qfOnZ3c+GufUFt7fXC/Eo+v9L/uMNgww8UBK22OFbUK6ODXXmVXXbX2VCFbVLbHu
Xb1tILvElZ9owVyNin95IO4apx56XmenzaUIGTOMjtKCLK5obBh0IHtjARDasePS
xWCvmgCETMb5U7cvKcROzM53LyBbrRXipD3r2qabVehMGCwMcjQj+KnzNZTveIoP
SsnxKrICiNi3lNaVZA9QmU0u3QHWyBgRiUU6TlZ5dgf+w5FlLaqS41kcDflm0TJo
xx59OLw57GBT/fVy/MZdWU6n2ZlUzz5tywPh/OAchQH5yAyiGRS7PJT54ATAAUC2
bVQMdj5hNtmunrXy3epB5sWji+aFM9X0c6pC/j3myJe6Y9QSzsV2GBVtu9U49s0Q
qi0eVKTGKDETat/euhQLBJ5UHG43sfKkALwZnFmoK4LW+zqyV/JGWJ4tNnqygg6G
/4lZsRPg8RFx2viy2tw4P/L0eKembcn4HyR6b6A9DeuP498mAZJiESz0kqWVWm7R
CZG2McjKtYrLgKK7OQs7xG0/zRt18aC7qgLBdks+qKiRblSi1L/aq4IL1iKzwuoh
LQf6XuvYlZ+CipqydbL2YPrNCJCOR1U1/9aRgd6kNl8DJka5bRw7KYo00Y4PVGw6
Xiw4iEDWqERwjIBeqQ4ISdmPNttOn9w1hhEIuA4QaedE0HazfFhpD8jnKnTu/qUm
//XOw8kcojxZ+hGN8LDJ8fcaEff5dsIBQP++cW5fIsw0wDf828f7LC+HsdUuqxXm
0jzYQyVhUHTew7oIRkcDHi+AMlaVm318rFf7H4PzcM6CMVrtIbT+gdI3ozrohrTS
zI/rcPkrsxqxyZkRsDhfFKBPYRA2FrZ80Uhd9I4NYN/KWdnZY7EepuVrMpzUlO1l
cUhOwWoxMa4o5XJRFFAUto7MVfVsbBHZSgyEUaxOiEANmXQnoAZ0JRQ8MSphSsNW
EYG/2PPfCM66rX6aH0KG5yVnTlfiBN95ojVb1E8r0dk+GfM2fOTsIFiITEKLBrb0
viBHlSo8sCWytpcxrmQu95d7GVTXg0bFWk0x6bjHhSRUlSJ7PZlSCoEP0Tfvdu0y
jHmshaUVMP3RmnCRxc1RJ4myOdhb//zZnsRzczfrTETapHHEg/q7HR+vuYfWM0KB
2PeEs6pny8pWHgt9BkSsWkg9qCzOHcEi0NyTOkSr2dKIaTLniXwgPSSeDJ9GzdgN
R7fqO9CEQeS+odIgVe9MnRSLj1UNwH40oEEkz6TNbGG3J7aWT/x0cw/RHd4TLbif
Six6gudH4gRtyR+THjc4aPm6Gngl86etd6gsgJt/h4AEOms+NOTnR4hfCKDZJc6a
h4tjkzgyKimYdwRMQ4TFbOV+8yBQixwrY/3Sqx6vLwtq2MO8Y+DLmwSu7HLomJ4J
BePazxiqMsOFZdhQYXqPG2AI3+c8B/ePeMw2AR+zcyKv6dHxIuC6pbUW75qixfh1
aJAmuixtTAlDROhC5i9iStdUiM+E3q1/bTA9kZaWTpPr5NJHJSs0+VOms/OXVV5M
sF6QGQecMDYqDyTkNPiAORMEVsNx6aMee69H+vSWDfYvzNNef0bljPGn3YeKnU6q
exT4Nq6yNzVpE/tH09RsTX9AoQ3/4uiKshxvjdQ2oXg72OtGfCBabFrvxWDEHnjU
UfyVevj8f8kRJk/lYZiJeyIjF7SISi6aAArhDHIZXjtP77QGqRSfugM2idVGH7PR
8FFqpWjIDn705qw2R+h0t7Ym62/48ukU3fk1NZmLoWqraHb4mibyVWug590EMiNO
GTYQSPI9OrJiB/CW1xJsM3CBRaO4ti4PcbUxcmM+1ulUCikIrB2DE8SWjDWnreQW
8xjWODBJ27PijYDgy6+vmajSLy4YeZTdcrYbyQJ3tU0sivddf6bBd1Jzy/m+HVya
T8Fnya+5JpSQFEccm86n7uZZRlRKgaezymqyR67qq101t0oDn7+hLHHyJ9gpD5b+
B2WjKHYTUj9uBNqUf2h/XH4bbvd+NFcD+Pd78Z8bo2DLrOTpAXtewS5w6c1GQffz
pTjihdJBDzslmY+7IIBzbgoN52ouNeaHCvmjq3pCSz7+z+SML74K4Qvbmf7+OWlu
3BRgScs4IO/5H7fwHOwef1nZoYyOVmS4Z2cWEDrhQo7YV5v0+xre4Ua3D3eLErK4
L6UwA9YzAdDZByd8T02Yw0DVtxhh39YagTt57Q8HsyrMd6Kuff1jQSBqDcYv9MAX
GeW7qnnOT1keGBUHHH4tdNBE3W8v3Gf0F1lxTDE3gORbyzBqFONyPYAR/iTcQlBX
pfuM4MkUFWaIrVFVMNveeKEeryQlPtanwg6og9kCTgsG+vkGYPNuVjEA6k2dEUXl
mSHfNb75HosFa33Ab8pocuyutDflSf4v5/d5GxkcPLneCVaZ9IYYRVU5gP1KdAWt
Er+4boYdoEtD2It8ct18UI/CjHisnFLHXwbkL7vCi/hKqOd3M1g7qSKSciklSiBh
psyCV45zy2ObdzbyLngO/9AxT/sxH8YX3W/9EGKX9eSopZB8IZ4aUZBRtrYqjPw7
PxPFMGHaQxdAf2c8g1f3FGwTlpuaP0oWUFhBWQXtg1S2h1Ha0Egj0PtNHAul+icQ
ZXfrdwT0UgW7TjKFvdai4afJLwYnEzaa9zQd7ZRzbFMh16+GQ8Gna4gylK28d6hA
6DTY+cSCIsajVoRKYbAXTtd3kUbFc7zBm/Lrk6vqicnIPFUo08fs6cWvE1ckN0dc
5Ro+U+j7mKfFIymZpsD4T1zzzB7/EwVdGbraVf7Gynbm3a7yg6jV1cHKLPrmKAbS
yXksdMOO/5inK4c0Rw8RdQhZmc8SyiGaxHHyg4PCa3FSpzGcvM11zRHob+4z+psZ
Vya9eqtsbPGYBI7GX5i00opSFGH1yQFMPMC4GXmVHanRw1/96S+iKE3A30k5HJJ8
PSYYvOuN1dY+ypgwGZZ5OMpBTzX3bUB47mcurKPzMFmVA6FmI9AChoRUEM732w6B
ME8tHiq8UD1OcZHmWmmQUoyfdk1eWVNurwy3BqyyaOAa0Kfk2OlH0D3/VDLjtGxt
xNpjQaSGdDy0kOj2mi/07aS+LDq23LTRh8LCBafVy18x2F814/O/Ly8V1KbN4mWC
6HMPYCj3y3OF16WpAofSrzrlKnyHR9fcfuosYwQ+xKXgrN7fRc3e6qKGrBT17npK
7VItF34dp1T/X1TN9pYiI3oXlImLB64uOJytOVeKrk+dvPTdksOqrdQIY3MNf3vh
mO2hGJIKuEX/sTd+xFK7suTVdTq9O7Rr9Zx/G9/WcZcXKnvUVqorUfgfGIeY0NDZ
cmvKFitHD6iyvOMO10OIXVnmd7E4tNS9biZiBJfe+dpfUDUBKnog3nQ89ERHlxJF
86zdxdV10btSM7kcW0iE8tIsSuqsBB+vNkw+iHp4Ygff9xPD0vUeAD7OoqQf1fO6
aE/SIvkfMGh3YSHPNLA0xGqSFjv12EvmcJcAaq/qsgHRbnq9D0J56TPB9HuSU6/M
UA9BtbKzKM4fbIHB9hZgHxNUzlTXvn1iMPpUqCZOWVC0uBHR73QMUz3czVbpWrTI
Op53zeO4hiHVc5oiSU9xxSmfK85gLVhAv0DFX8+ABhgZWEItCE+3EWsonaxAlR11
Vw1HehFbKfwbjSa4Zu+qLWECTbu07Lc1UoRoZSvABfXyLu0s6K4o8nwnVGOboJal
Z00A1iYxCKCGStLWjZBwdC9bj2VUi3pAiP6JPSrT4aNs5MQKwJeIfubSR0aC+6ah
hw0DHyFbM+3yHIJmIMdDuW3DOtSwPUrgS9/7KgLWbnwZHblXMZkjwuXiDj932GoD
yI8yOIOphcNuiTFi2uKh/91upZffemYViLcz+6eNXLVk3x3AbE5Lz59tMTEWuIu7
bobtigi5MZ4lzhOIcqT34eEuGg2F04URR7XpP+O535L86Ars3hZG9XDd4Iqu5CzV
9lsnG6FYC424MOz6Tv1O6BGc+//BnfpENFmrtZGGVk7U8CeD31zWmMojlJKuKucH
R84i9QPFyznMKCeZeyhDbt/dtNSfOSx2fNta/igJVjSe7VpHQHffgXwbVukPeqoK
m9nkX7MnswVU/47c1sz05YF9kF3t2AKV3PcE8Weur+u5DehVuMex4mPPdjHc2ha+
6f4PeMRU8DG02g/y3zTUj6oJnWbQIEkdS+OrzPN47iqUt6WlX8IJKYFbgFzgUzyY
5LKjLRHADcVVJ4+aBbiXePW6TeQyddIOmcIh3csaZB7NKogQGaHiMJTTEAQhVB5T
NSqpmKqaKJR310BgQLrIq8J28xDRRJvsVTVnCDL9bt4wbGCmCJe4k99kHS1/aBPR
TNw2j3qHnZxDBqi543nUh5nJ+GR7IGLHIbRgVxwTrPHgbcT57ciTBtUnU0nQQtfu
wXdZaI5xoMkoDezinynq3BC7neQQy6qIMiavFSMNO7maZqRPtN9baxlI/F1U2PK5
bnFBddh6ThtFvhA3/btdKKj6AbQVMTrozjddtjleEtyYPjbuxfd20vvRyf9nKHqA
jNROk9Y2+epBh/UtDKsd9LUkg4NuMRY5v8Bh2ZAGt2ujv7+NX6xp63pKpZUy/3tN
c+ghHjylrjORO956cEYS5gPVSt5EbIBtvUEHie0XmTkKoj/qV8hlAoLgroO0YiDG
/HIp4v+eioppITXG9XkN1ChHubNfaUXH6A6QGnce1SgkE/PF3+AxF4J6seO/qein
b/A+raIakCu6NQ+KeR8PD+OrG6M4LBN89GGcLFrTcqrVfEp5TL1JpIOQ6bm5LqMV
XFsx/kZwjsoqCj6l2OSw8VhF2LgCTUI1tgmgLOVm2D9qg4hdPaYz3ezlohRdZg5H
TeEHIsj8Ti/m9ikWSeUK5imCR2E9Mrgj45wzdzgb+k7eXgBQ3Gld/NLr57kmCVS6
Dhr5PDFY8beN9JNjHUMv5S4yl5P5EDR/iT+pvUYid7llfx+ErPuCJ9Yltge1pK7N
UnRUejCOE9fvJuBBp1F+preOrOvoTFVGeFtinBKRttWMQeKLCYmeuo7oZcr7nJfw
1hYPOgXoyAOm8T+vns5g6h/en/+55H4xXR0RKctWNaegxWC4IoH8W2IRhZgXsxCY
l+zvYdvHj966QTVd7hRjN8+tF3cSngh3M1zcnRFZMcnq8mpQ0yAPUd9+8eOpojIU
oYLTDpne43ngxU1EgN5QWjwolLRxVR3374oO/5s2pFq7AvYDKFNNHjCpXBzgp5FD
jK4XcEgpCX3tZNpBd1gx7gyFvGhJrcXrcKx7qRFrZR7ERMrmwaGCnjhWkC+JSSTy
tJ2jxZp+9pluq0pQ1jsJSF4cbq3VrZWx2rjHrUpRzRy4tHNokfdC0/dHEW0TaQtL
ZU/R8e5s3bjgt2rNMR058XZKKd4sONvvL3yKp9ECEGqDNl/pcFxSUAwYtuCd6GVx
nthmwUoGvQyXIwxpKte3oDYcqCdks5RsQcM3SKNz89b6TIQdY9MCifpIgQC5BGJa
+aEnFckvRGY0Wzi4p/KhIVrheQsl2RDGvJYNGI6wUZm14203qrntS8ARWrucjSKz
oRg9HdWcXkVb+lNbXZwSofefhP34A22n1U/bt1xdvY1dV2LzHysTpvZz2TKOLzif
o+W60KSpokosMJTOJNyBXB9vupdrK9FqfVJuPprSJRjbp9vP+aH4qYqc7FUwYrww
gR2KaTGIuW5I2Noj2aOck5QKyt93d1XTqEbJaJginS1K1vnXhHtW5MZxCgliu/8e
otLsSVFKC3x+h2vCASkcQEouBJgxte8EYF8un00arLD89iARlj16GF48kbPxxkyH
h08/95OOhvdGUEZXUnYiXT7HPQOzec5dPlpA6nMSI2wr9tIelZ3b0MmpOFbR5MSa
4sUXz7+uRBFRDuutbBEAv2Dzf+XNKshjcxGdqnjhq4YzrT5Ss0lUcNK5fpLanL6h
V1p1qjogCyucEkV8iPvFVy3OJRQ66eELaW/41MQMt/CmxIxWKylHa7B/6r5vZ3li
k/HmG6bhjNsEsuusPUijRTVOXiCqXEMidLSCddoDlo0vzNaV9+8RXlMk9PC5Z0WN
K9TfNUYF70lDHyZBmqD9tfCEgSRr4/2q4MKd6tHz1/3VNSS2vhOhf5eqHwvtC83/
jARCq9yPXRlluq5gmyKV8CJfiDtl5w8D8zlJmAilrI8lTRfBALmh32qAfbFPrLRP
WlppaCSGFLiZs0/BRfZetnX0Ew0sYowNsaZjhQp0TBqjzPos3RFMBM5zGxy4O1d0
a7uBRj181rBmTUZWmk79amqOUbpm+9TFFVNOAvjIfknTcKxMTINR4eOWVCOmF7YM
ihjeTCJ7BNdvyWvV0g5/CAqoUd9TTDi6z2VGl/9aWvXVnWjrEy3/7eM7s9ck8ya0
s9N+7/LbznBSvA3yGL4qsdd972EbpBzvgD/iWu1LMArx8rrF0Ff4NFTFEeBu7wag
TpJIT3cl3unOPUGIHi54IdPEf/RISXH+pVtunbMD9iTVJJO754CkeBZldDuu64bK
AxHtDBqNQ7nMWugBJb3YjTVdJPzxj8/b5okuZaIkZo1/4KuQNpwrFvGfO7wRW1fu
H9PUOdh2wDq8P0KZdGPk/g2sgIOPUHFxBFGtoeR3P8bpQoS+iqWo9J18KV/CJ4jo
CS38ALAwmRqXnWeFk9lHph6fcjvXJOfQYjS43F+n1i8GD7CKscUCLJuh5dj0ZE+B
uZhaGIhhFBFIBliAL+UbYN+gIcIITgDeCHYTImF7+STuYiVqqO7jbGnsifYsX+D8
Msexem3J3hH5/gbt+5OxtG/Fll4hDJR9O6JIRSUdVdRED6JMb0SdEWubgd6r2WPD
20VbfaY2z9m3oFVgxGWwGOWpNlCvwdSILU0MV/U+dDYIskazQYzvWCbFNJ/SsaHH
+PM8c/q5bYXUox7FJkcBsoNcMQg394oc6lbpMNKaankL3U9vCOJMG56Lx7kqfN3F
fpmQCO7GwWDzgJX8p1IdTt4V5wUeezgWUU4jCmEdGby2gpZ8Wp5fGu7mt8q0PAv3
I/uiWccW2F0gHJzsfN9UbBsD6n+x6Kw3Ov8444koZEEkKlEoLFGPYCUAoqT63I+V
GfUiIKWN+866RA104dH644O0A07509JjTWtBMD717oBHzPE5wk2u9gLI4T5LVUm+
JoWh9Rzk63j5HPPxG706szZSeWoi/fY7mJCmSdonH/DcLXstm60RI6xfjJrmEujo
kO/fWbPRqMX1tqvxiPgvOUJgyDy5xkUKhXnxj/CQAJL9aFnGQR/STjfIuPHtTONJ
4q00TLe7gLs/zsN3/IqjaO/5DvGwBv3diSi4aKVJSCof5XfFhRoA79lORJQ+XXat
gUK/zoKai+S9v6aREVcCpjQt/sFHYi1Vpk6OmfYNlzYgYB8npxdbysHh7+ui9VNo
+nsyz5Ifnpx4SUbNHEGMU6CchGz9G2JVBHF7xHfwPlzsLJEAltGYdV+UnOmSGyqy
Yvz7HWV+H9WcO1ZUPKIOyFYj4AQptNe3SNNnETLGacqwVdxE7PyteQR3taGMLp9s
X6TlkJygUVLmlyD7QsOOgxgKxvHU7k/YMuoRonEPyew1V5t+wvt2/rvBPbQqyggV
q23/OisLHwemkw0kXYN2cjSV7Gxh8LDtLmWRAujQslD8Pv95zoie8YNA5n4XcFpT
gl/ORuNpAQMBdrRg8GQxtnYe2/eMMasPICsheFOUFXqsJIzxMjSf5n9R5rFlkhNA
lEzl80F19oOL2jTOMnRi4qB3B60tl7k0RSst4fTrtPWiUjKpdLEo17q7ZPLSihLi
+dHksjBtyhDADdVDm4JarY3bXgkoeajwDLmUYn7j4clkfIr1O2GKOt3QGXdyO5ou
h2m+eGaUsSDMtHf81N3YxQTpqqpxc3rwBodxMKDeoVPsDK05baVMT90f2gCkMdHu
trjjpYfxOOrY/mwQM8mruxS8avybJAg1Ea21cqCbCltPYGn7PomFCBprFR9KP5I6
jZmXNLGZGYjwACkwygvJfGLaIoSBIFFWJZEx50T+uPAZ9QtEFiHar3oPLSYLDXyn
lOzsHO4+U0juEyrkLSKxY79Nos671XA38zHbNIN2+/mVH2kPv76njGl782m4/u4Q
Tfhr8KxvZQQN42kr92RMWsZ4wreQjahg+JJfe7Kd5m2aNADwvPGPlwPQgsu7iwFR
OrA4P2C6U0EksuorOwZaRKyFSju1FHXQB5R/RlT1imLmNUQCcud3EzhNcrar9BuW
r2kFq6hi3oHm9t29VhaXbTL3qmnCslZL02KoJHLHLEJtGr7JPCgn6DNHfsRXcg03
0TusipQtdbzamZuUDuV3COvbspUXbCvgeAmkit0PASWiSFbWAUKq8oRlUSXOfdCN
6NNjrg/FgK3YPGIfqGLgLSlAmaxkQRCPGTJj2VXmKiV2xmRdAzt5DijufTg2cYAt
gEiUEbxGVDsd4fZVj8C+pLlRxgeljKh9W/EexocYoK9hktygnfskX1iALNPcMC/A
mHUEHjgj6AB0ZTmQ8X7h77T7NYn7+nDmAmoeKvx1XKwOcwUBiIofETe+y0OAgTOH
q1dY8HxFV15ABHa8SdTWfhBw5M3xZGnHx5vjJ6AGBdUf4YhcbfYrkNNvVSdkCXHh
kgA/bH0FvF7VeTQMuAk00s0nZmEhWxqt3A9hQWNx1tsNNW8FGFmDTWCtNwMP6VRK
6C+Q6oC4M/20sPDjQcrTMKWm4IiBVCKpQP+1ERNJ7JlSfHH4ifCGj/4+z+JiuSEb
HkVlp6JTLXhxkbAj5nmNx/1mEqrwWDpa5GI9PXL1AU3a9PvLFWm2/62DvMLT35zZ
e7Ku/9thfUjMA0i3EfMuLubA/Yy4Ug+XbvxLt4H1/tEvfd8+as52PrDJPZW0tWuY
ilrlmAu0LbwnXkKl4v/koNUYZKu8yoEPFsvFyfysyZEVmXQCPytz0Ng6G9g0Ea0R
Jjl15sKT8VPHrxbED+eRBAkq8sdmFOY9a25tPrp8cpRFhZdakkW2f5/ioV1zIuKJ
fJRxAwwUHBkhChOnYe1BbopAKlcB5MEGlW4FzDCe8oUhdlrYBrItwVSvrVjtOtec
DNF41tEeuddfr5z9UG44w5f92QE5pRG+rGl5lrJUFdj7cJ/Fkvwl56zNLb///Ch+
xKnyc1ZR3/EBvV8Cs0X/UCB03zQDNC7AkacmqDyN2+XuLurF3G9MM9sOkuXAIzIf
sJjU5BkdqD7/F8vFxOUqkio1duQ7ZZW+XBuml8Z5XiCBDdD+YyZK9wWkwwKi0rPu
eNbe7PdscwloTmfpgCm6sZ6CZxiCTbMY30Uk73Mu/IS2NJqb10hMY+OGoiq0VqdJ
MgvwFMRnzNusIxEfUylh0Vl2+Q39jfq0FschRjhMQ26V9p0M/plGPCtdh94JCfFc
pRZTkt8uhF39K2+R4HbBE0fpLxs+6l4FW+FweB3ofKWMHkrDmi3aKF8kLuTlujFn
wq/5izdfGJfmF3CH+oE6IYo9I0FY0SpqdGf642hYRsr/+BhXxk9kzH7ouYZ8unfl
B4qAzVJwvBLM9wmtDM3V3o7SbIdUK4OIHglfdtkcY/7wOGwMgI+IYaOKGBZnJ1RB
FePYLaRc0zYkg4MMV+y9hMhTXEKRpWoEB/b8UDl4ZqorZCyQXRshiMdcdem0Isxj
pnqVnDrVIuXZnqcaR9wpOUoWXJTTUzbXS/jKdHroD/OUTwCtPhx1k8zDidzRCMd6
8m3OBwLw0aPQY5JU32LPXmgSI4whRqF2WRxQgaQCIRwZegW7A4o9ILcoz9WlQs7A
6LATYDgwTev9qltjAxQ1MjjA8uCckpAtYXKflptGRQSQgpcYcv9y3Tcx0Rm2+DyC
nMpEhfq+qVlKQkVFliLA4uDeq+p5uyW/0RA2v6Ck88vqwSU8Rg/PS8QsnebdUKNC
gGJyoB64hXE+PvbOMIw6a5lAY2UjIPBTVLAsbJJHt9WSK5FXaTBfYh8C5teKeuxP
BwUZsxzRe6496XPsjiZnHnsFd8wtZJnHRyCjBvIX/xg4IPvxP8ljTGGmnUybENNP
ivURcRg1tCutHWC8bcrW01jE16/8s18civ/lFbcqDu57XtRNJvQF2cWaPm3hNc8/
r0/TbJCr9KJCQUr0fVV7SVL0pEF4PJlA/blroK7hWqS1KfF70ePdof39mTma4/XC
XMYRI1qzUSrH1Lea0VU2N6anBP31r2sdSNk5jr9QQ/IcK7H6DumvFeRPKtGs9Eu7
80C4qpoqiFk0KjjviRZUuvnjGIffYl7orRTaRkahLAFjcV5yIxnNMbTQmlbkBIDY
sHtItPtuOoHDyf6PGDVD/fzcA1TjqmnvdzjIiVvWeDE04XybAFLbkHBnkDbYVHDs
fId87XnlOCZ5o+8c/8rHyqVr5RPexXJ08jx5P0VwQE32/m1NGBVigWD77BhEUtwD
nCSUqQixOSOVgTqrH7+R5Nmoacl52zuwt/Plfocf2Qo6uwBtk4rp7b0iTJjavxcP
rvvZZR0PZRD+aJweqgPOfa050aJgYaMiRMEMZJNzSIDB3lqphEiSo3r8bzg/H3LY
CuaV/+1+rbO2afDKt0+RJCmIp2BI5HuPCbgaoUCS0wOOShgyol76Fau1GW8WOsux
n4n1SvisLJFz4dPiFNEuoURfWoFRqKFkY8o7GhUUEjQW0/ydAKZ91p2q3HcYI+wF
pThatxkPaIrsluKXxdF+c42+nUwogSOhLlOvcbhTyT8axOWurY3Kiiw+DSKEp5jM
zcH3Y7Qd3VPK+SlVHt2eQTKElWZ4OflhYe0k51nOcRWxF8sqJGV0P2I2DNsUqPFt
waQ+FdoOkLJ8CthSqfEA623pQf9Mnlyjg+oAQtv9fWR6oJ3nN0MxOdRvi4n/VEaQ
6I6J/ol1xZDEUdFTwMFTnk68IT30QGIYJT6Lq1Wv15fV51z6vtyaxtSvgBjVg4ZC
6A2tx2Oeg7mX9F023t8YVnYdH5ebufJ5IQypzEQUri5hV2OAwt8XdpKPsla9mVdJ
mbMJlQudmAwaJjbLMNDmPAV079DDdUOb87zfH8XMTtjjdmLocmDwe4TI1VbQmLft
1ytEPyZBZ4uXhwKqDS0FDuDPgmjfBcEgGvE5n1o/8WHEjCUZjKu1NvtMqfTgqzDy
W9NOl3cNgOF4KGn1hNKsu9g90m0quHpz0Qns5yKYMLDf4rbDhkIJFmWuByvtxx17
eX8hFAEx3LfSphKMDXua/Bgaw2SzyC750p3TzX5KTphFhrah3yO9k4quoBxGTMQk
j2jwTiDfxAW4Me9LXuHN6Y+vgpYkffqj/478bKGh+TXRfvprxBrGBUJp5x0BHOdA
K0JPWMcNhnPP+PJz/ulK+agM3VLlkwXdk3qUROaH3QbLzhlk2qnvaEvNf8SQDNS2
t51xBTCe88UXV4hYBrFAsGK3ikfDYA2NmEj+0y1ix08sWUIP4esRUGV4yGQwwo3S
HQmul8kX9E+q23Pw0gZ/fUYarM8y7NCI+gpJfmVH1pOtHbs8ySvX9QK3x/kP/dB2
GIV8ftnyDcEsLtmUNOjw6u4jt/tltDeAgGa8uCnjVPundepgwPp8idkqRUuuCDIG
Q1Gs5YEgVE5GWfu7P2qdfO9KLJC/thjb9JdWJxW/HXmwvL/r8VaYZZDyE8WvHBZA
9s6JJgYW25JAapGEO010T2V5a/MZJYaWqzm9eEEPmeQd5rYdwJ3mr6qpABAHdmib
/Tg0RIEU9fZxD05GEqyP9pq1u+J2hmdftSzqKvCsu8nUj8z7xLcgIAOdlf1bE4Ru
1JV8oI48czYDGv/QCHLTD9za0sy3qbLunOqR3H9I1+3yGnJG9ZySUWI+x4lAO6Mt
TNjh90XqqsBN/+v8jtWFg6sXdao6cgeeM7cbA+umkysvdyv5qPFqU5T3t7XXLMFw
7pxo0gnyed86XKoeC3g+GauYjHCeDsycfKcSH/7vjv8m06+zDcs2i0f1HfI+ZFG2
xGAJ2s5C4BKkTkNDARXbacYQfPl7RTaWuCmvN0QxRvl+x8mnC2ywptEVM1ccJZaK
rWujcJxb5MVmQJIC31KVOBok3zGchPmUL2IlYs/2Tj6RRWSTgadpP7ll9l27Tp3U
ijNiVHT8mtHsnPSlW7SLfyQ8eINoTn1a1gEemC329TtkZaYyYmCM8E1F+nEMoW3R
2ZtSmSJoPClFvGy404N6Rc/UeBntckduKLHfhV1O7QqacXmOIBSFUc8CS+UY6ijt
M6zyalWBsf960BrpI+vlUxLBi03vyAyvYMqF96Xx8DAb/R9j7q1/TDXkErqjV15C
d1TwCH4ZJWcKYyk2ibp7lUlQ+rWUbVX2nphyJTp5ERDu0ZLVr2ea9bOQmVZjaTTQ
tGb25xzjcmOmTNnJl0RFzD0pPRs0joFaGnY/UMXfT6kcNx4WPaU5mskvDrEmYRJW
fFk2EdBGDIINnUHQFF10tNveWJPSEwrknufrqLGsV8MnM3/mMRcE3tSdKi7uhy0N
fW4Y82Pbbr6JrkNZTxBqGbSsTK+5fXIh02sQZmPxXee4mOK75Qi5SIuTI7jhWwu+
BQD4G1gdHDTkZGEbrxPJK/v4O99PCZtfqxJ8YkbIJ3T2a439HpnOi2xxcHaYbS2P
paPtHfNamR+lK1PbH8k0Px5iqWV9C2PlmoCQSpVoD9CvJGvDdOp1k/kPAOi7v7I5
yorINkHl0cKSt3mrycHC/G/FBcEeQIxxkgXNAI1arUQxpa9dMxHCeMt9ncRwPEEP
mjGEQVRyg/NQnQuoWOjiftoRNlksEtEkr/gBMdc2YcCQ4sSwlrFwv6JfxyFnRUFW
9105AqZJjxP2eRtY9KVzxauFbz6zeuUVv3yqELWpZQlZePaysY3/7ucCxQY5yXGb
qvdMGNf/E7k/xr/LLVIcFwmcrclZdVDKFEHaoPOeMrvM9F10UBh6m+YxgyIs/FTw
pAqrqeGzteGcDuVF1Swaz3gAEh2fNJ9IXuoxbZSO/NfYTv4r2KRkhQF4dHU5ANUX
bD21w+hiSQzF6mffmHsFqerqXtxSNq6YSFFO27GfikKpoLiUbx1dNn8ONbJW2S3I
6nXhuhULoF687tv6Bf7C6ahq0k+ODUdFflsrcV8dlYTP7PlrPqNvJplIbQlM1EOd
XHKe1j4dmRNwJwK9UGBuJ1ASmatyRFFg7C4pKKePEUvd8pq9kwjKLk1uHKar6BX1
r5U/nuFrlDu3QEjkyRYK4Jcricf8sBwTxDtNlcXPs4W/6crcC7aoVLHV9a3j3SYX
xMf//bpVUojXtWF6QgeEzZbq8wdqwTigUofg+XUeD5TgUgJcnSW4B55csxowb/Zv
JnS79TD7DNvfWNqW+38kbyiFvjqtz+0YCH/LMVu/4oi+WUnJlUWERCp655O/56hO
GoOlochF+fLiH8wEOiUFaw0rBtLSpm5Ql6YHreq2bpi1h3kpUbJfrAMF4tGW4DAl
Rq8oCH3rLHuEWYWx8HRFm5CIl+Xlg1I8qeTtXzGjT9DePrdRxnqmDtwcfw0Gcd7C
uqpX1Au/KFhrYwMb6aHAOH/Aprqp4FSo/KOVaFZMPAnQeht6hFPAVHBiV3bV0WtH
v9BtRtoqX18rNO5mveKn4C6bSvIUFU9qB5ITgC2o/O8vfzUDa7qcVKJ8RHZCTF7R
OLJqbqcsXgxia5oKp0RkirzntzGvX9hK7xLP/xjCbakjRoDVqx7kI11ywPzRjG8h
ZeigWQhUhVdotSpASHMhtT7FLSWvOJJID9mriyDkScUNLb7q7VYRZLmd3F9319kz
4bBGYKNeKJEW8Gwwh3dMc47RxbHmyEqJ2tze+iYmH+jbey+ChX307kiBeUF8rqbS
o7JMI7HuiBLkzM3c/ipKbyWGQfcIEpMzpD5xvv707cdOZM4YmWALKvrH4yvZdMl+
J5WsYyzGJiYx5RB66BHeCMg0QOAN+1Stc83zPXSk3Unadi7Wu+dmW7Y/YHllUIwR
xtfDnb7eG2BSKE/dyKFwjKvzzEBrhL4vP089xqa+Ee/fqTVfQ8iH0CBvsrbP3pe5
Ypt3r7mBvOsJfpCL3poMqOCfMCfJ7n2bsHEPhkDppUEVMvn0l5x7NfUMzZvHV2Lf
2mRrv2MqTsZvoLDd6vI63CCoWd3La7gNbq7FjG8TTE0qmtGFFqTh4Nl87yMz9Tsk
GkEHp/8LvLDslTOrGiDEpXtJI8oqL5FRIueBGT3U5PCtUPO1IFgPxIPOrtrTUpq2
fe8VVKjJx3EUnOQ2du5APgc4ihMhfg8N+NdXfk6N+voJWTyvxw3QGdLpjB4z2O6S
5cKB/Aef0CTFtEL8bAoqaPjAs+rpO2V0orgif+1BxZjEiC8IhWWWPzdzAO9dlAvN
+uN6UPWFTVSwot2a7nD8p27/cpzISm6Q90OtjRO8fM20TwQkfMBlq7Q1Dnflcny0
qt7xjZjeQKd4ugecEe3pgoE+q+CMmkk2xj6acd6/hsfuhNawFewPvGlKInr/P5LC
QmBHvRx+pW9PITaVfNKoCpuz6E6aMkIFNT61sSpa3j/UTD+0mkx3KiBfoYt755Uj
ARzHdlmqXBtMZxfjVW8dKkI5h++iNKLsUeopsNkYugcoDLKjmckF9VO0hFhUwwsB
AjXx29yHIzLOZp0HZhCPJppCzVPntK8SJPUpwD4b9jzmmN4aysYEGk5KwGrMVLZV
H7U/NWj8EctrG0/ayXEE4AIiE+PQT5xnkMd+e60ijo6puS8yHYSrJ8l+510HdnQQ
Vs59yAvmDMAzEbKcnYf9ihpb7qPw3EuwdkuY5tepYRIiV9BKnJd8WjNZ1olfkmTW
yJNfXCcDWpyC38Bv+uxZLqjvmJQBEMCJFdZQSnlzHlnFOUJQPUZHIBSTTsgBVVcz
QoVe/nz2ag1QSQF0eIlKIixrrL412Cs+N2KmR6pZbltYAOrAuGej2sPSVEdm/mD/
VVAMp5Hwm5xpBLIEXbZWYNqfFNfPWdTgWzszs6QOhmTsXErUTkLBcuHE0IuWuHr/
8ALmGFjIBNU7Ck/+Wn8AOniD+V/D2oKwJNvtOmdJCt965UW02QYGG/Xh5cBYtrLP
qBhVed18WgStEmm/vBFTCH9eeMvCarl8z+5YaV6AaLjhbowt5tyQMqXblIz/vQxB
AcsTBhw5dK1Rv/uKmT83vlEHsaMFCjRI2NfyYH6PNgQ9uW1eVmk+AqPTaQKdEwX7
/u5ME4l1mMmo2Q1hTAKB1nGnG9R6Vh8UyyTJPyk7Obv87aZQQK9ToIm/PLF0iRyd
ADpqPoKvay+GfO1dp3z74Gctou0uHDIkmuqDsM6ucKX+Ay2GW5fkp8U3drig3uKu
n6gUXfGRlFbi9uP8/4YRqkKlSKxcMyJdacPUB94jXHKyP1JfxOI0hwhqAYaOql/h
/N2DF2x3SeZvNb/ILhKkRcL/3+KP8eQe7FiNF30X3La2kPzpbeQ/uBGMMCz443ha
b4a4hexGXaac0nljwdTxgDDmGHzJTAI/qMSPtznVucD65yympcUhTERNqaPjkxIE
ONbTee781LuCEv0dyDcw6xi0ISao41OtWaRYzlAfnS92PajggjlKP2DeHCnG5iZc
ERcN7bSy64CEzWVCGBRkbAfMyVeCwfDJ5wvcBssE4pJIM+/yhq2Obs2QsCFwLunG
WU10i46aMfHH1Nf76KCu5nixj4l278Rk7f3dLFpR7ur9KJ5A18KxCHsuWkwZJPlU
E4LuMxk0r4BSxVJF2q3ZiFrYIigzUkboEDqqqhJAUZ76aJ+CpNWfdL3PQPLxxI/y
lDEKicavfWGErHfZ1fHTuGDXzb+bsn1CRCGDfne9wwi58Uh2ZpWrnUsGJQ2g2Eja
0jmFxwncAjmSKXm4M0VQlFA/bt9L20hcACWn2wpBLoqq8WTGN4OO/jLaQNKb/YNc
KtnFbxRkcAGGKhwyIpjQTRrhp0zxQ9yRQ77L0ldVTiVWzGi0BwmNpzkP53jtxGKC
KNp+qRt0GpqLv0BxPr7pu5bhOB2axks7QN2y5NhwdDmVGldH7xrmATyoaFkvrATm
b964aXhR02vxg1jvP4pNjzBckkl3MY8ZYfmJLvCpsJPk04FiE9qOViewHRcFivR0
v9Phtl4z1717xKdrpAxUUnHM91xFRD29g7WJTxD39OL5SXSEi6H7HcPMLFDT4e7Q
B5hBrbdyYA7u8+PpRg0MHB9DaQHkM163GhjYz/F7gStecYHozWIZZv6Gr4+Oh4T2
btbZq6OWju/IuLKjuUxentVu4xJPQbSURq2zft/VVK260tJVfMx4+l+vCGATRhA0
9cQhXHhnNkn2z3Fjxd7umPfKT70gApzpDjbUBtoOpryGJuk+5fZJ/Q6Pf6n82JJh
Bt6ShqCBegIHsSBf72cfFX78OXEfPzsHIV1VaVnivM99RNFNUaC8Nf0XeVxUkhNz
iDDKe79DoGlDKTB/fcnDXBoGJh9+N9LYKaeYXcjy8Lneq/bSkQajQe9VHOOPWJib
RQhrXtjRiQuyQ+mvnXGH/bzJdgQ7tMLpCzfXXmZ6gdRy0cBfonmODTS5ZXxTZY8a
094o/yiMsiuPz8hoKMnjptYUW5a0qovv1JT9eeQlirbsqT92OrOUXicTMVjcAlx3
CALXATHG9rjNNnR3N6u9kO6eiLwrrxiTywBuoVir8+J+u5cY7FmGUbS/08rtjOT2
SA7zUlC6RL3EmnMQwUxY44QHBz28+l++p1LayV1cCjV7py/01V83sCRA32/QcvhO
cAlbwVlHojd2PSmRUzj+77HtyP52aqE05srnQDcNiDyWegfNZV/iw1B2IReLWNnp
096RPMBjjswqpeuZKYaYeNAu8GaPNNiWLqEF8+vX2+6VQckJm9Z52dNtozRBDkXy
Eal8+uLI1P5Okaj7u/jeIm7diY+CS1gwm8ECOLiqzskiwKAfth8KGdrnOrQ5R7kK
+8MoXOGp8rEFG6pcG4AXr2+F5xreLCUtLIhTU+JIXxsAzr5w2l6dy33pHHgMC1XS
3BC/yvP+iNm3aTm9DfWgKhWJ9vlDXgNUxknNSRZu0pBrna0kNCJr8nt//bhWt23N
hSqIz8KsZDWoiE0tTgVAK8KXP2IP7s2Ak+7YC6ngXN/2u34+wKwlkoZX3uGN+mIq
UcbW+5njz/0UUSVayMfG8S63XJdfkGZiZsZZXZGfYj7+BKVzL3vQcOvjHpLdVsg3
hB/97HyOXmvNCVbVzDLgBHvd4c7mKRfA8lTpa40q3PoyltlH/rkbe4CnZfmWRT1N
WLJtsF8eRI3zTwQgOOud0OmqCFXr3P1F+P9vmUY6vBer4vhXQIknV6zs6offVwek
/o8U1SSuxiXuQTbeCJ6GwK+LSKBsiR71pDSqEEfRJOqVJV0YiBGKQwPH/fwheFxK
gs21Ckgl3QQELyEAuBhhRCOF20mnuQd2lBTEYSdvesMIeJCVFfHhHRSCoJEEB+33
jKkZ0/NkbOuqbunBagx/4h8/TZIK99sbOeFr1XPHPgRMI7zFx3S4qlbOSBY/uPuV
+gw4qYMIc7Z3OuSh17LBfmL7hx0U12KwQIU57kZy02NCIiPRk8kTMRXv4RTsbrA3
Ihpivkw+rvNSmckqjgqOft8oqpnQIhxtXgGjAts0SUVAckBqP3LWdaSPmw02BHcw
08hguZsZtbta6zzx+3fesyBSwQjiFE/SjJvTaHrg5+nXd6PklWlX10TubiIiWpM3
NIZGBipGJQoOqmwrm4wqOLOBs6Ri5eGLDwkeU7QzfXwrpUZhai0U0BQBFZ+lyTV2
v9VSAGNGWdD+eIjtiYoXu80e4GuyJALobQPLYw+YPm1HPOVc0FUN/OGJijv9Gtf3
OkTN6q6mOt1M/H5OV3u+eMtmCXXIuoKKwl8GyunYBSSZ9nySoA6wbSQi2JOWoyyP
zwxqAmBkYQaUv5XtoY4065F8jUX27H3ASgt44xLQT06T9IHcQBgVbxCkLbAQPKdq
SAAxbAJs2oSjPHfz3jGLwHxrJC20jK6soJ8CCLhH77sMk/zes34YgSR9rYmcqcnZ
3FXPzUd/PTTUTVURB/R01iebPiTZ29dWIUFYoDGuGfRUJP48Dhhy6I0EN512hY1a
AEIUmRbobPYvskwoACuplFP+AJFL4i/Duat4oz/Y4b77WlFNf8S2JI99boUA5qGn
0tmsYwVJL29vJ28sMJmI6kG6nCVFQuAkmiNMdJWF9u1H9PZsNLI/pJUne2DCoOd8
clQGZ+xRHbliY6DVb4oFBpXXRdZwApjEBUfO6P3A0QIPXwJMZExN1q5MGSHBiaLf
QeHPjBWbKQ7s+3NSwX+ZM98Ny1Zv015O/FtqcCO3+EwoPKFlBPpZU/VHvW5bJZjn
QBHNXj19ElnfPpVQDqigD7AX1wPnia4DBcVy9LIKVv/BCHpx1vDkus7bCSkkQUfv
QVyjTvX2PVIYVSghWjdHIwo9+UTAkFIGf4c3ZVCSohpp0VGg5N3ZYPPZdRMToi0T
XUrCjNVDMUAHTp5Sp2p6OoectaRayA+Hx0elIR1m5Yt6zvjNmX17rv3Odp+zt4Bw
kM7tmmJSZt6gsJVDjPyOcgs8ofLePVQlczZNckagoZi8PdOSmRTBqGV0pTvDnoQg
Jkqm2K4nyVi2sW5Qx39py+P2rLgEfvsS47PQRIRPk3YC3lkL98n27QHQuTDc8qcU
7/zPm+MENnGy3fasAJ4khoNj0og7UhwXQMFTToPOHrTYDzWlgdJiDtB0Ebbr3Ok1
I17/Te8pPHPhpmysRIv+vg9KY5T0Ugm2SyOgiYIKFA7z6nOHimK0p52oRq+DSdGp
bGUNk02imfGj/49amI7pNp52C2E0rUQFRR8EnBy8RXHs/geQjit0WoV60jsIWxoY
jt1TeSYmoJj7P4zfvdU3i0/AXJgm0msgQDSnJrZm+gc7BYhIsOAeX8B7Tw/bzP59
TtS5VaL3S2lKGrNTTcQV4h65SoIzn1Cn0Fb1TfMdZNqszkh36zz7c9a/wyUAvJt/
9gUojKqqAHvMZfw2a6LpvzcE/gN/FxzPvBHtl5v6obDSUtd2IPNoaA8o0SnpI5DN
5e9dxFSY6KbSruAYXT4ZMGgFNkxUQa39K3h6WkcyKGx/DtQq2MXyPYwxa4GDPsvR
CxgXsDmkGcfWlEo+bYnMSO5hitJHYX2+Co0KxzoKpCrKkInWtkC6eRxaGq6MIP0J
e4lQyyYVuVjFE9bdWNRuzWr+4mTxb6ZRP5FAHe4O/PuYGf+cSidqkyLrlf0WueXT
YtW+0UmuJPl0B4o+hBH1JK3qu60MDRsK51dwgTZ/+Z0PZb0yJzws21WLyyH2h7I8
fj28HuL3nYnEBOwjqOBqtEIlv9Dqf4z1zkQtfzPSVj+ilJMQUbE0jlL5p1eIPlJI
e26vLozp2+QDC1BlrG6oQkDKB7DeE63ecUnVnkbSgrTDBoOcjK1hTVlM9LALLNwd
Ntg6sNUZZfknAh8FICoZMNHKVaXRPZLiSGqjGV8FRkEboyIGoGDwlnDT2SWaS8dC
ZTPOvkp7J1FpFahCH1Rnud4tXkiorQLQNjqus8ASlIpdApFrVckEV2R+osC7Y819
vDpAxK0BEjauMgifyhK7HTV5onKHD/vSwgNC2kQHgEbbbIZBtqfjTn7Awzf/HeZ3
rgq/6V535vFrlNW9oD5NZFeNq+MhqGUC+II+0Lu6x/0JvUXSK34PBcroLEmZglCa
2+q7RESlH9cFwaj9LmLEy6DcQFGs7oprdMiBHhXZTZ27I5gqNYBMsHkwMFC8kk4O
Uq09P2DDX+OCGApQg1oU+ALggVIeJLeaFLmFsm5rwLQJTbASUUp9rfGzYc6VjCDg
yd3EkCmv/Psy3RJVt87THeUMV8IfnhM71JifRjWyTtpM37c4fdf1bFMkw7c7z4V2
ShEj63G5hv7UyJjav+Rlb4/IMCIu8yM3kuC6yPV3of2SmdixrRCx1JGalGQ/Prv4
v9StkWhr6g9mqQrVLQWdHdx6N6swvWz8RgA7ceJ4dzrNn69b+pnYEq2h4c3AVRaA
HzQ3RBWEmj7IrDkKDniW2C5ITTWhclU/6PKTqN/YcB316y904Y83qzuFJo5cUkSG
IBNgpcoZMYjqLNgpAsnyfrkUg38RCBIdbfl6alwtmWqm64m4eL7Zg+F92DsRhsLq
+UpbutsJsV8CxujcgJ9SaptJFPPHpZXMnrfxaS6giTzWW+2QUB25apCfHz6SXvoQ
mJqPjNxl2QFY8yV/J6nyVKhF6/wGvdHBDYMUWlujSm3qS0tXu2HHIs6oBdJep3RD
VLoqNs2GVwnZ8f6EDGLefY/4karuo2R+fcC//RGeG71KfOS9fjQnPKAKCN+fUN9i
n0udXI7YwFO2Mwa2WBKU6lImJko4e/GVXFPCNKyXgJI+bnEpdb/ki+K0O3I3OL+j
GVuud6YgV+9C9HhNXN11SBYncxbrL2bKSN6/W7K0u4eFLBqLKwbcQzi0ucrXBeJA
OdT4mk0CW2iDY0aDO8syR3EQZn+ExgrRRKlGehE7XIqBWJHovC77u/Vw4WpXybEX
YLchFR7krIkTdJViog1mAdZ/6W2v1EHIHi5pGiuzudWWFVb0kbas5p18L2xPJjq4
imlzQIZqPZMzSKnGb1+RBwC4GRygtv+IoKwWl1B/UpUsJVGHMDkBRPP4deBe4kgU
5WekXJoIEbg26nAzjT/lFtS08IrX8r1VOlV+shBxbhvjKQ2gp+uAqDNizVznpxwi
urLh7h+++MtXuGbbzXJevBXoIGtwyYHpI8iYrT9HEqUQbURqQzdYCtXzp6VAWv74
gZuH6Bv2gRKyDhEtuOjgv+1hHoyRjFfsLXs0fbbfhPmHddSPz8xuI5imzoR/e5vL
wzjE9rfWt+H/U1s7oKCG9l1j1n+mFkaXOqZnj5kMKgiq/Vv5RgSd6lCrK9tagOJt
waTaxwoqLg0brz/SESlISkHPXeTkSL1Q1Bb9VVDcnyS7NycW7Qrn3brT0uP2tXLV
kO2++sF1td8ByhfBp51pwGNVIOPsGZCWfgDAlMOBLnDvVc0Halyj2BWIXV+4QZ0A
Ojp0n4a29pCBsoAioQAwqiANepRGsxRv0+Teossa7gTqzZZrZWuxKaMK8cZ7BKDv
ZgxBXVOF87JZHS5SdDX9h5E7BiK0egQ46R7RREHF/2hE8hHl2WI64Y+QXlrzXoKY
WRKAfZqvD+NIHxklbo0HYNwqK8OtJbpruKnRoHoChiAkHPfA2DxOmX3nGa1yqv+x
XMnDBUizFb98pFm7NlC96BtKfSY7hhJ4sk/5CJvlmam8PUBnXgY5dZIxTjKM8E4W
QOT9KUbiDvAa6pY2dAO/7RSNRfRmlon14ymLfulWnhWbFD7f5OqVRJRsO8TXg7E0
2DGOSr7limvdqj/l705fAxYDe/9ETBFJ9GnAK/6KsKWOQC97Xxlm5/g+wdtXRp2w
8vbBDkRA0gTDDCO4wF9+AXOTWu8iiwrZVxP1n5kpMGRZVWAjLo0UvIOKVq+RHtXd
aNKhmVNv3WffJtPlHpVFahOiG9hRjpjyzfaAe9RMFYBqQb2pXhVI4Dq3AJRsSQI1
YL+kwht6WSipX1ohlGrH5vrKs/OW+BgMg5nCZTefdUiW01tWXwMWAGJlKKTrMnFg
E89egSF6B6C6uu9rumHj+xXUFoVrhtu1C1AZ/G+RFM1kKl0ZanQVm2WYMFXSJT+A
T1him+wmlNEYE43BkwtxkbDZW4Ob4bzv3LhrhSinLaLjKVPITwWUG36qHGetVmTM
6zzSeTPfNjhYWQDTNPWcvkPdXlYypzQmi8w6ZFqFjD9i7mBvDqFlhknfgtVhV5eK
Ba7s4bKxxoXj/3qUCbUof8sCf1LdwCLKLE41c3elG49pLl3tm035LuDjzlXrmlj8
ipT1QqYtTD9yidiH+iPhnKvu+uOFm+A31WXUYyg+Ks57uLn7AQ6F/ep4ZfQOBPtc
xAPo+t0JxdcD61w2Hx/6JYn8UmCVUUJ+HvCeSCnK41dZz3pXGm0qQWfxgevJGEGC
XFUZmkcNxC0evF/zW51iS6Ub1rEnrxhTnQnHZY4YO0Tnh+M/TX+XcLK+B/RcO5h7
5oUx0TbpRbXaB6GE9qkQe3+cKkM9aAzqIALxKfAQJeL/kU/EH3HeMhhIJEXVKIce
T9dg8C9J3EKFXbW82/e4O4RBqf3Ej6oVRUuU7kM6NY7V0M59SbRFuOuOfWw1JSut
O1TLjYeCx0Ix84hbNwUCjIfoRA8nb9QBx75bxYelTAAymqp2CeoeXwcyhXzB0dGW
p6Kb7L/+UezlCilwK1VETCnhpOJZt9C3kZMpKbvwODmxk0kwilzxoFDiPZGe6E3e
NnDHkXWuNRVV9mQmwUBTwEAhDYzmVxYyC8KqUPl9fBWQ56FlotzNOYqmGOxG/AZK
dWMCt0Rx4H0/FfASwWrdpQw6IeUQcW6eiS0nn3G/qJSn7f/L0PmERmB+SmB+bMVz
qTXdzLiY1vNwexwps6LdZFNn+WMKxcpNgS9MP6U9VNyIwxSbvyntCosW7d7qpkVK
OfXB1lYBH0K2m4tc90gfHXGgnv8TWqabzliGYEj68cFcrHIalCb56rPKDLfYS5Fm
g/fWdFLj1kuu03Xkzg7jq1vxv4zemoBvybdNh1k5XrCaVtFHOEjTdjI/WkE7Csjd
4b1bYQhz0k7aRmKEpwIpS76ELCq9os6PnHCSw4noEKTAdaIYPQLuDDu5UYc3AyCw
ZtRlLuI55fXiO1qggu76rROb3dDvDZms5VY4VG88B54ymNP4wZwIx+598EKUOk2o
AA7RLYUc1uNt23lSGQthvs9HjvoQxWGQWWo5DREsBkG9DFvywAeKcbbT/7PR3vqv
VZIdxufqTBB5aHZacXg6G1RSkjYnJIocMjq8CF+Oz8vLJiG4WkT8XmTp5YqtFwlG
S6UZundHk6EKh5VyzS9egECU6oW+aFw8NGJXfz1GsGhSFY5Ur5NST93LtP6EaoQa
o0BfEW1Qx61siC/jM/i3JXC5PbmyhiFyTGfBUChHOAi27EOxYADjsFs79D7QBcKs
sOeDe3Xq0kYKO1Ll2qn1FQO/gX9I6Ho+fjxC+mI8SJqbDUhSNaeByfj8fmy+UnnZ
59tMAS9vESBdIYMMnn8+6ieybCwRBlkcLXW7fI1JqkGVsnT/gBYsMVUwjevjgT5g
4KSvBVVxFuXbO1EDVoKylEQg+1NHX8U8F+c5IOySBJFd72ryXGx3pvt4LwBETpmr
a+LYrY7xUFTbL0Po+4tTZWJ0op50njFDscSB9QY9P7j0ij0aOKNECPBFVurkoHnJ
wK00gFbU93ulFIK5BSCmjRySz9RKbBYxQHPuCW7I4151uey6/zXrK5vVX4UYlzZS
qap5+nCdYW/jpCTyZQU6Dt8ZFV3VwcY/HTtL4MtQ67s1YlGTsEQSuOfIfj/At6SH
enRh5LViEc0wLhNbjMq6u/YGLci6FEjT4ahMR+Vvdktt9AdDDdu2MXp9/DhrmAT4
xywBIgOFRa0tfxGILF047ExkzQrH3WGsISNT6UWBEFnqV7HclHsB0u8zd6wH/Kcb
XHKn3fodpvGdiZ3Q/1vW5Io/DGKRgQAwo7UwM6EyOtB2KqHIx3N0T1QDP9o9DV3Y
PO2P/L0/hamX6px3HJ+zleO+kME27LY+HeDRMd/IXZVBMX51VgcIKePdgshNvfTJ
btKVC98Fm5f8R5ffjJkYkG98JEztUJ1/oYEfRSZPSVrbKuhfzWo/mKdaFvShu00I
wmLZ8tqXUL5jiit8OB8rKMntNFvO61Iiq2780KgBArRhPyZWmZRZwbEVYyWTnMmK
Tvi9NjfJ9WUGy8/6HDloFvXVVM37bCkEvPzzF6fHV5v/15eoCnlJ8lq4ZH6qZAhU
TH+oX1+T8hzbmDE6o0zdHxzZ6J1y/LLIAm1QjREDi8XwqVw5pGPqTkb/bdgsvhDW
wFJlazIDavmYNY3I9RoHbeZNgnKKNIdVC/1jJ1KfX4PqOoCkorVPRlt9rEmapdSy
qz9FqeRGM/SapLARamHAtoIMGd0VntEZAoBhyaaQJT+Y3rcTgZY1F2+gsE2TP6yk
ut9YJahum8sfeiF6YrInQ5z/phBTix7qZC/XaTzvOSo6MqvOkJHJ8smG8ldTY+ty
Si0EF7lR0K99KVD3UFVix+ieI0LLQoe+TQYZBx4oNpHC/bTDavlX87MUWxCIkAno
Q5eNcM/wvlu9NoAgbU67gupe8g5f0UqYUQoZxYUIpWOi1uwzuxkXEhjxR8iEdqfj
Usi/vNgAMvWvIz1lmIsvo2/YqVKutlSeVS0U6E+42UFL0SIPBNUVWZus2d7sd3hp
kC1iWsTTwEtRfN8YJFJP/36mSrJ9aV3EuzLElqm7GfGodhPOWZXEFvfmGA2iz7T+
JLdxajKafn0+CfZqrcYOVZzLRrXLEueuWVDRyTo6nzf4gOS9czjDoIIGzx9Ln80D
NrbYLDloR/afsCB06wUEBvpAGptzt+8KAxb6HAsYTYM+oIk502t395CvbQFmdSID
HRYEgNOPjehhRIdkzxKCYAANNfHjCBMjpVRX7b8GtAmxEabXBbOHoGnRla4E/SSX
nyfp01soinZ6hoyPmoFKT+dhVCj5gs4BWwTkTwXI5+nGX4loBz7sKAYLnQV/g/up
rD0muKeahSS56bZioe1pXajfZ5aKu+rIY8CecEpO+EpCfRUaXgCnOp3chpvQuZOq
gybfBly+a6a++D7gTihrEi8tPWvFV+C1ZEEFWn4zXAvNpZuWvzQbNScjucIoNNKg
Z8d8lEkvmM3qRLLAwWNTonnkeIBoBBK94uDPLBZf92GpeBWZyUiDK1o6ZDe24xss
wU7yZHAOc9SG/pGTnotmoXfJdmo7c1wAxf11g2oybs5afLukwM4on2AVyoTOKoAG
f82O/3rO48IwoaNcrVn9yQsGjk6Iv5tlNPDFVhDOQRHOrEK67Cp42NPlw6SBKhKE
CNWS9Gne2rWoWCmzzwJgRJPmoYAqPvRx6XHyN5QPnLNApq2wmMTx+nxXlHYwZPvq
6iCMYcxaBkd5/PxlMcesw0m1o8WTwNaekkKW+zxrrjxPzfpGoOI31JPEhZmTRp4Z
8l8vuOBVsOkPCqhKXTc6CqMoX8sqXJRph78voLXrAY2ljLSlrDYWgxqVjRbifdaH
Jgtu8oMfp3qBhC6WqqRPEGLr59WY0BPT+ARebfDUGBE7a4n4v7HHKJMTPVYMaf2S
bj5/4dYXFfCvz9leoeypuD3kXHT+7SH735nvNQESz4erz+5URF/qdD00O6M+D7i3
ZY2lGA1TDNOMrz4P80UUufu5j9tkgsK23U+ZQsTNqJtb2HwI3FyYbT01T+cwFklV
7yKE1+MaNAA0PWe56/dkgB3SAg1oamOoHbLBOELOE4tupK/9HzbKJmd7mp/f6glD
kk1Hj9mCSj39NeIYXBbnSneuwMITBF+5ZywFy8W4A8bWBZgNb/H8D17Mox+nNgUc
SjLXulVLxTmOh+4mfpajfMYH9rzKW75SfoZwdSGNvFl2U1qRYWUsdRYxyBydyO/I
lfX8WJPXOkvO5+jNX2yPr+L7eLFHVsHmO6mAKC71irFxKRP/iZEjEUAfzHbfl/8x
+G5aYHSfxgSQag8LDLFql26sR9mC0rK8tHMUBTO4H6za9d+pExH9+oxnsLYbgYGH
c/z0E8DgkHdRjjP4xAfCicKdjAve/04T2Bl1acEO7wuwJGdjiIvj61OFNYOEhekR
6BRLw+/59++FwoUwxE7AWwwknP0m5vntKCHdej65oI5bk/RXYzX4ljrCOf7Tzowg
FI7D5pXYthgEjvCWbtp2nqdC8vvWfNEWSxJdSpHuhinrWbA3tIkpjm4mv/vfGU4z
XF9f8MIaNZrclIGyv1wyoU3fGKDaFcFqaiMN1TtiAtasVtTBeTaWOvYZEg1ONLGu
fEBWTV3ui9e9bf2TyYL01NLn/V7y6SYTtsneM3i5EgLi+w1g/PD3AfSFD9TkoUoL
/8lH9QdP/dpogxJVXbggCIS2kxn8YoKcxRJw6gPUqEpuZ5yaUvCLHDPaALBhuRRD
euUA0q9DKJ/Qzl1OdCWjjaiQw1Cbww98pA+QAJ1j/6skN+ZgOCainHmq2Mv5lhKv
3Ncg4NkxGBlVjTvNvnOcfxx9AUsyPh8hwj/+ydwKk1fSd8CzgGL6VONkDhNRTj6H
GlVkLURVV0rLd1Y/WoTkeJZ4Fk9X141uniZleddDebaqHnkC1Bol7Arsdur7TLWo
KYxFUhoBJ9skVnpmvDrGB78qK7H5jiMU47ff1hwQpuU0qonv5HaqQHTdP6mgTRgN
PJNFUW0i5XMwrsWYZqMYmTOYpj1vfiyyR3N7GmUT5qRZZXvmU8k8azS5bdzy7OCZ
Rt9/NXnleysZdC7ggT6rHCaIJI0VTcqDmPImQEJtuk98ZdXQwXxahH6ZY+H4yX42
m8s8Gm2+hrP0I+Xmb8DHBqpTnT6/8bS/bB3fHOXYrdwLDpn2toUMyJSbTFw91pkx
06URqf7gpo/O5JwwgmnUdlK+Tc4AGAdT76QuHxMnpOWlbqDkwCYn+tF3Y9vBDVlf
A7tbKE4nm4jqr3mzZHPAxCG863rwo3JCAGafbPoydsUzerNoI1Dw81fCKGHui2zw
eyjO5hHhUKHP/U0bI9ONPthawlxrxnomBYKq8wSa/kAJDTbXB9ogHsXNNiwW4XaL
lL2DbMBVe3OGFt97RAJhNxEJZsW1Rpbe7kAZ/b3DOU0na55p/HzbzrM2dxotmpbh
7+ZoBpMAL98aKaayvWje70P6AnMB41eY7nmngp/gTa/f8oD/OOmtrtUdh+66EexI
qNLfxfPIHlehNVd544ecsb8xA8+y+9SQXpHgD1j3CC09q/jDB2NPZG3+QJS+bRW8
P58DQHrjhvI15ctv15mMeK1HUYOIUhvMjRxB5aT1YyA1qbn1Vhma4rpXYsF0Yyd1
v1K+fZsvs8WgXKkD6Dtj/szw8q/YQxT6WsIYLSbk93YB2SLhs06tW4m/9Fj6GvvW
ut3HCCMVl5ukFikWdI27wL4jCnxKGYWCNv/ClJ9yBi1MYpjfzErzXk9soJuYxMtV
vdHPF30INKWH9aPyeXzYytt468NHxy959p2kF360GLz/PuFiB4PCsGT4XoctDxrs
iaRgRHx7CqaSVQMi7O29gpgNkqqGIfufnKaBuR+PR3fdj+ehAvH86Q1sh1S5JgS2
1Lz7oK4FyCGkfdM7rQynW/uobjAhxjUMMRqzcbhjkIf3FOn8NleECARJr5wdNRcN
RUOF6A3pACjJhlRDUmJqoa/f4pEzLtA0eqfW/xzLooVe3SfWMkiwQvNiNiAYZRIu
UqHSXtbCoP6Yz11vpcJKtk8xvOe9xS8vs3pFfyTwIlhwmRZlvwsbwMwF183cD/Dd
m18f6hcUN92lrJY+3/jflNWuphu3xdtYkC7GgHcIb8zKr1QIyjF/tMPokvWYBDU7
aI3Lru72DRDYcuLWbtfJ/iBImCssDu0Ad6OcO5PaGXaXVr/Biohjox3kVO0+mzfa
6gGk4B3GksSoIRG6Ezk7YnfqTo1ut9odA90cBvGyyPqydkWHfn17DK2rSzLVm4Wc
PJumeVqDc2kGnjtjk9TX571a1IF8hBAJf0aK6WeZj34Cb7MQGFrvpJDxTXFJdqbg
JhJID3OmNpXaERwWD6v2/3CArnC2nnTuS32ne6pzBFsZdxE7pSjfbHPu6D3u6T8D
oTk3T5oULAF8iNs36XvvOcVn5Nn5cFSAmBeO2asTlMW+4EjQYZE6JPPDVmcwfntA
4AnEirIDdBlQRUwT+Q4HMZ9tqK9w/3kxyhsOGnKSpN24D3m2aJuu1QkFkIirllxm
/jks8je0/GpV3aCrVJf3Ou7cM3XQwGjW/6V4xHMGSnev6Cvs6FuJ406evKjPr2Of
lt9kQir0gU+788KernTbQbl+k5ksksgzzYTaS0xJjIH+GeY6npEGEXrSa+BUMh8X
4/bAYNVsH82/WZ6tkRrSkPklYXXe7SsN8l+ojKSGh3KsARhZPQ5dzcXapo/oXvOX
uMI1XZHTpIKGZBLrxaMdesqeypWhuajLbYJvHgWwEkQyUQ1U9EQUz6+7IeUZhwjk
dIBvAcozAj2gAXIKgpDL+clw1xUsQO82R2ZQ2dT5iRraOjxHRrac241Nmm0YOJ+b
CabsosZZMr6ZfPz2zcp+lf9rwGDqNJiNVOTXWEqsBoYibfiVs+Cgnfe7AO6ixO5s
yUojvaR55KC6TmXztk22MDWKRQsNfoHzkCHYm6aOTzi/scNFe30Ui7jGwsJpVRb+
ACOvOsjZtF/y+xAe3RtqPUC5sk64rTyoCsnvT09JCOUUWIcstH+9kmm6JjdUpbot
2CslKUdDje6wjgyr15YvAxNqrszQwyY7HSfDfsDazgGfTK8gvzVz0BRqjz84680M
21PLxf3tWVjcwi5i59jpMtIQdf4vNaHTIDRQGGwcO7k4wBbDk5xlxUEvu40DOz3l
vYY6d7GaivMdV0f8x3sVKmcdD1AGaD73SC8p+PFL6hPNDjFjpym8+Bfi3NW8Rf/u
KlneEaluxUQ3eTUM1fgNNzjRZ24TZOt01Ua8c6fv+N/Reta5yQhs2PYZPXBQMUTy
HUC8f+EaMnBTESeLgqQU+hKTA+0bftaYLi7EX3KJ24iijt7RPCK33yEn7dv5/+FH
Pio3t9NrXBDdmurPHX3jhx0MCDXatNQYE7HKteV7QkfbOG7/hzXW/Wr1DCgDp0Az
GbSOd2zWevNM18NX7Da4GvPCZJjBZZBipA0pkpPEVsG0rX8hUwljmD06RIzGHhW0
AOjTdGQlymX8uGEibdhDSTRz9zsNakDSbr6U2Qr1cMwwAa5Gdthno/zzbgOwRDWc
GyQfykNUSQ8o/HVSNrR6fm29pk9Lo3j1wPtgh9w5f1bv8Eq1ibJG9CmRK0RXXWzy
ArsryhntHs7qyIzyQ94KGmHvZ0roMsjFXohJoIuAVnSA0aygbNq4UdoZ6RA8LZLM
h9+FwA1dm6VCrc2AUwKz6k4QMBHCuigFcK+vGTwJWXPQfyJTnUcBwXD0gL4NqxJB
bos8FJDuBCGhAW1fDXyoQ34OPtdAP570hnSTkyGHdae5jTRi5WBLx4NUsJIgwePb
WoysYCMbLoX/NFz2Qrr8XQq4lpen8tRO1QFOSZnM96t7G6Q+t5SRtgMyxCY1b+Vh
dkiLh90w7B8Xa/pUqMuo9RUY81AP9Na3yLb0XXQ78EmYENVgQyzgxYDdkJVcrMPn
3lZWPM+Cj5T6WXIKyZMFtzErppJeJL+vANqVTy5NB6mOzb3FhvqgLRYa5KDR75Xz
MSoP5buZxlYBSVO7Q4YjFSi/oY/akspk15iv8UElsHo5p3nrazE//xZJBbdNWzGU
CG8iENnLr6LfEK2M2xGshru7i1ZsuOu6sZCbVrlb/wtcGjnybxhLCfSDSH4VJ9k6
Ro3N0vwffyCgxnhhW9sWvdph/BgRGbHdkdMmp8UC6X4VU1ziFTX6GrFF2CvhMrwr
dznIlbsr4WtpEKGE+cyWOYKENMD63ATiwmnku00cHK458FcP/tN1Wd3TN5iWTPFS
NcTeJk2sgpAy996KpkE/BFZnmy4vzPONgoVcqG3NYWUNKHAO0NPXi5F8syl0mzKw
muGXNyrG8YmByHiC6W/W2JMkxtVQ++reUxzPIdqDU0RaSRvdWlvHwzdSXoa1sSJ/
o1MK9hJAH/2Fe7430qmJbb8bnHlFbokUSBgaWnRLw8f312snqK3qx7MwULwX+RYO
lUK/zSWK4rOuJu2IIg3fZD0RVAyiEvE9u5WdoDj9PVXxCwxSq0aki6hbmo1h85Tf
ELVvIiOj7sWYhn/ELno572V/ExlgtGIEgnX0B/2u/fGrZptRyTPR0p242ltPMSQt
CUPtZ/3LMK3bRffC6ML+Kebdb4Xf8+fLw5P0cZaFPDOTR479oh4xRYYYjES0PyPv
h+Wc6uH8jbZQwURvyDWdBYJ5IsWIwXUbVv3V8AIvOssuNPMvFcHBr8lQ77NgGY3E
+wy24roCSViE/XhGMRpmQG1QFd96FzkL6BI36gYgAvpwWYN3OGyZDIM1VhfhsXxy
78ACIisrZQwe4//ZzPy0urZvSLp/Y3m9VxSAiMIdyPs3Y5adydAqqGqHg9rNjyHZ
CIOmpfsuWlvrS4xJ0LEMPJrfNRiQQjZWWMO72Iv/O5erlesx5KD2aF0gk4J/chW2
GHkAVktrLmknyxuf3XhA8XtzdYFTFZfwE8EmdWdUK9W8eegYGEBCEO52xEL8qV/O
vIb4vEutyhTiQphyH/UfWWfddOePgNZXMFNtt/KuOjUrvKUqVmVBn1biaabRyLt5
dTeqz7w2o/G6sSHNa8wrDVvU63dcz3ZuUF7T0z7odd8+NXvP8EN/VAZmTi/oU/3U
xOFXl0+WuQWj225FqG4oPq4HlFqTp9nlFoEzW7Lqp7Q7NLfOdg7kHynvuDU00VK0
iqAXCIu1A7hh2eRimr0aSw692SlSLl0GMg9U1kzZyhS9c8tEw8CmfZHV+ImXt6Y6
BctYibpX8sHZjHz6Pkj3F+8QdBsyoGHHDEl5FYf3TYcN7asSBMwPc1yQ9vzi3FqI
lpBsKzlo25XayVpJku8VmNrjXCJ5q3xqZkwD6tsTXwkUFymlSUmaNvq09k1e3oe8
VqmluqMqQ7z7pZIjNMa1MsPaf1a4Tn/cenJEpTvJdwitV5ykaeCsUqU9UoVXS4Rq
7b2HEEVGnQyeMTbKr530bKhGUB2fqoCn2gd0EPr1Wv5aYIvNgCoGctO8WxKEzRPT
lpxhv1t0yneCf+dNLQW0cSZtl17GqxE1NE+hJGBHZZrc768QyFRtbJFYeopdbaJ7
KL66c4rfBeV1ewykfy1RsAbSKkMYtHz2fRkONV1TKq5qjMuIhqVX6bdcx8q9Z9tp
RS7p+2O5p/jHn5Mj3nWUL5uWwW24mb2ovR9jWyrHb+kPGKG35kmFKfo6npxwl/dl
XYqgr2WCSCKsfUTIfdooTzNoZTk70SxeeyTzUTBafos4x/cmAEe1Es4XymPPDd+q
MOOU2eCzrbUkNnVU17gU7dhmDl4JbZza6ssdjFXggX6RzQDRHUH7XEeKu199BC6q
OPdiKIg3qyHV6Yv3IWXGvtFsYLQeQumtJj9KariowbL97Ar42BMRVKpbxy/QqAaK
y4pyYTdSCOecKLNAu804zL2z0v0h5V1fn1vlL6M8slmGQp0Mtmos6UmdudUT9ZiR
EJd3uT375uVFCsVs7m0ja2wClvcTUi/cV6+aZFEB0WtC5WceiM28XaNircFIHxLX
9/yYFZ9e7xMduPL0iRLY5s5Mx5waPe41b9u5oF6MGMuGwhc7JWVE5FZuHHU7Mf/0
VKZWMdSgui4XWxaEkKB+AmfqcqWiKbmzgpmjRDEtiorPRcqy1TmzSVjiYmT7WDj/
H0cx4jRVkFm2Dgoc6FBJ0OsDXiJJz7ERAtpRIYe9/nrJTat318YPVQVvrGHykBNc
46kFZ6VGvTr+f7hWSdXnznmejl8Tk8ZgeHQvmxz0qhdPQg1KyLJRW5E7SXwldEFb
U2C3ZeK84JbXJk5hMPaxmJYJn8pFBz2FdJoOvxqYenfhQipIGc2DvBDnmES6NJui
yiPMcVL5ZLcJfBnmAlIByou+LkhGMX3zuOeIMObMHdyj8mnHXMzXCIowsQQ8HhQC
vzWbcnf7YJgWt8iVpDEkqG4FlAmJYyG97YIa8XHvG2ciUANd1tgSpbTTSDJCKjci
OG1JAtPwHM+j2qjEclsl75G3BjPTeP/Cwbw53i7Rul/DivcafOxHEguaweTb+Wu1
nE/2pecdAurggzR8LBGIQFUTNc824eny07FtdaSptTzvpnYVSaOq0nrssdX9mSXK
W2rHg/xeNwlTZbt3+sOjaS6Sr9OuuYJhz0sIACfN//hBAjTICE8S/O6kRid7Z73i
jEz8TOWVwudYf5bCT49jfrx3iWG8BVHWwFYVVSQtH8qvKUHKB7si5b3umUqSUtwJ
rt9Ai8IITPTEy5Nld/aLuYlQNk8dBiaF6sy6vrORloaRY1L3vbNiWULlIV8PYsv6
/Yx/wOpJjLZTUiVlBT/N+YAXiRBGrh2XndynrYtSEyA3/XWNGCCUVlONwrbd6VSB
d3IyjMjdmpLssXvOAgRrJ80IKwsdvzBdHtmL0ae5dIJEJTqME9uD1I1y8Im0LYPB
K3x6xxLjI7W3Hu5S43y4xzm0T9ad5sI+2cJDg5/G1nimXfgK0X3Wgc1go1cG8jWm
0Y62lVV4aT6MsJltuk7gu2uVHkKz7sbBvbH/9H4DjuXm6LFAw/GEs7x4sYst9DNX
WKnvbU97EE2dp1+N9mO4QI7PZt0fDj5oAGLEPGOSLvDymcZ23JuYOTKZpW+MwZIA
EQpSK4l+ewj6yJr6skltGFkqgGof6llxMyPUTZYHuPf+Rel0bnQCKTHYmfZZQ2aD
r8cMXeO9c5f3Yf+bUCqehlPPQChYBtmbvHmphJCNpACovmDw44XPAVztuk5ZmTdT
YbPkna/na3wWL4OCmxfiQqZArvQbdj4A6Z4sHBJwSfbHnImuhjAraLurTomU5WOl
1t+cyPRIxciq76rjtheUOUyKkfg2S5rMHYpdCyyxYkGCPMT6OFq4fEinXbOR0caj
ew3a87dHfY9p4GzQi5KseJe7ZvXhsoYWmGiSfd8dvGa9nKNCk0X/ltz0lHYwZIfh
Qbtet+FczyZ0oVhp1Kinki31yk/j/+loOGzuu3wTbYsi2EjtuItlzqYWl2wPw7qW
pRc/iMl5jeQD6Du1jvoPs3idx0XPb4pobSfOV3Yw1+RsvHnCCqvjag8LdqMEOmkz
PqCQld/HvuMP4oZDCx570h+1NLQHSSyuVqE4p1tYzzdMCKaIzZw8BBeZlOd2Duna
/eMQywWWVPXYm3wrv4dpKu+F0SuB1qhlkJoEcLbU/0k3BZq8UYEsoGd2TJp/HyCB
cNdbfnJB8BEyrExF9BW/Q7VlNSckMYV8lHwv6XuCz2LauyeVKRu/u11dPdzByl2X
dLDBfdOXHAZITEsj2MVt3Uwo2Q/Pv2Pezq2McJC7nCrgyP3b80sXmZRActX7zUgK
mT8gqn0jko27SbWy/VBMIHePFzf171b15bRyZPLUhMRTYcZR2NUNO6rH7FDmg/3b
hnHtPprIk6IGMhDdJJAyvXwE1wJkA3Nye4j6IHTISlDDSGVNhrd+7gMvk6MPlPyM
GxK/Df0Kjt9kSec5EpavJbSsn9wFXrxbIiHd6+Q0YqwJR6dXwPE09ZbSMHon1+a7
fnjhsGflZuTup94rqjLNOO/KgyTkwGeRcqzTWZE795rf+b+YRsOIQFrWWte9hL3U
/SBwoUQHcYPj5rhGLNtT2H9Rkjs4SGrK0iHpKXDI5PgHCPhgfY3OcnBCYS6AYiHN
HqjAsHmv8iYydZ+IJiNEZcPBrzH9Gk2mesQy0SBs09glluSlpY1TRzS4g5xF67dM
5wJySvcSsg+PzCfVB559eDIRckAzwoBzbdE2rihjG4Wmoooxw6D2m2xKVON3W0TR
mopaNRpbyCXHcskOt3jIyOnHTBGrA5aPmXP6fohCkDTIpAuzbFme33tNWle/xbdy
p80yzNLhzudjdh88ij5uxzDp/dcvEiQXOOsnSju+7QX7FiY5mDZrV+Rh74+rnTlP
/u5fOhJVisz6/4WloEoTBC4+f9t4zBUBtAi8wUOvn9O8KGmWnMBWH/kcEJM9rX9v
zZ6Nf50c6rWViYiIunaBoYEpw3RxO9rOHkbcraaK0a4pPuQ1K/dCFE0yXyh3qqxF
FYPHYCQRTbMf4fYv+sqML8M+Idn4oImahg/wQMi4PoJfhSbfhdBrq77/H7ro1G8d
rfEffwZN4zlSMBRwGb+BWWncyMH5BGZ6b7BRYQIGrLAhvh806mXhpYau5+cMg96y
1YrIaO30O4op1H03nE56Cp+f6aPoT1T8FvOH+Whqc0j6ZwLXZqD7bDUGvr5CIiX5
0ZgiYg+aGHivXW+k9Ida5CAUw0FrAcfpdN+AuayB+DI73idL8dAsBVE61Z11lUny
CJXiZS490BSH/LxhIcrkV70t2vAR7S+fHIB9U1IPlvP+CPgGVH4/5SoAT+e7PeDZ
U61kkIv/oqjzdGi0WzhCRSO5zWqBEghY3LpdsUMyMbBbeM2kH2uOK2M+eYYw1UzB
EqzMivYlEPAs5AX+fTEEt1nJUDXj+ttdv9KrwF5RjiBCeDA6kRBKK5yank+RERxd
afdc/HSGW543kH818VmeyzLfyum5fB27wmz9+rJfH1EBiidflV3rfs0nj4zCZ4dL
BEFXc63/wc1jgtJCdMjKhPRBYRNvdHITyqgpWbr6ArgUDZSHVIONmXR96gRDN/uI
HBsOAruvO1xeV0pXfKeh3sXNbVrhhV5mNENEEvYILfBk85mBIoR7tTnhaxa2CS6l
EIa1kGR6r8Qrm7W+xoAl7BqQ40swM13Bg2bSOioIoCoTwWrqLvTSNqXOe1TG9m/P
siZ8XDBeasnhobZPNEiPAHmkeU5LCu5QdMVaRZLgUE+WupQKdvMbrx2pnUIAPMmQ
w8TFz8EBZhy5h1fY6SjbqnTPg/e9Z9MI6txNihNIQKQkn/IbNaRqDP1I+WwnrLRB
RMkot75GgyVhuIK8/xijSzB1VyDQjdruk2gdsh/PPJkm+D98mqwF3h+AZFFFhhBH
UzSe7145IxDtHAjx/0EjHw2hXsCEuDe+T81vsTpptGowRxTR2GUuLT459ijcz9L9
XWA5ZbfWWv7+LlwwjLaEQo9Ep0+1H6ZthPE1EFo7b6fNRqosRtM2sfOsTzkVHb+H
kWcMFdc0YFM2dDwTCeZzCoqVtxX6kCveCmaKuPHn28plOVhQ3cF6Uz2pExWKUYR+
ZYlHAP/qZTSo0inxkH3OYFIrNATgLxSwCYBX51YJNo6yO2qBPF9WC57x2lQIvwJ4
xd0sjYw0zMWX0shq3uMGOqUHDw2F/+5oRK5bFWXZvvSeYa+upKclGHqmxkM9aF+s
p0n6UmaaoXI2KUjUJvZulDqRu6bnEW3tPTTDo/SQ54tCrTZuZHm7Zh2FuiRTUAzU
xZH9f0m5iZwpEEe4CtrKWxw3V5jh8dvTRrTQJ7C6Coq3yMSrGaCs84zycgZfUuni
99BABgQ9qimJuHSxs+nOitWXZzHDEJIjGRIBkriWCQ70hwHWeY+5xdtYdykfRsuK
OlkZuSZo0SsWcQJd1gumVMWPY2mOEI3yH9Wa/4YEi52Lnvvs/kEK8dAGGaUWto0x
ilbrxy9tRc40Ky/sBXalfontTcHpJRKVvGIC6gVg2UToGcOAqSc5Zttlvh8P/UjK
sRjwTvBFteW56MsvOBkKdt3udH0k7rtVrB8+Mo2TAi7EWIEske51TZU4u9dhaLcB
xWWaD+3ZDyXPjjdnlNiuX5kyp1xcPxjEKkMGeQnaVIZo4px+/yfBaTGa1zZ0LtHt
zA7B9p01CTxEOfxhyFP3qzrhcmm/OOWvI0kPl8ZqGdRTWjU1dP/AGv7j4CcQpkdD
svqSW8ZVPTRlbgpVZs/6W7m1rpJYF8tUxNh1oDv+vliXzhSNg2BEaGYeNQCPVHtg
d5dpUKXp6f/RkBoy+rHxiqB1w6kBeKUXcv0cx1hZCS0kqQu/uIAyeBUdUh07TKEX
RCS/+xJcNEtkIvlNKaM+olF54urLoZymE6FJFdZCDUX/OCVqNaXvagTRZDq5BqHH
A9UCRVdFU8oBpsztNhspTC2gmsieTe0Jx/uz4e4+nc0LBVlbDcdKU9NM7FNKQbeH
VJa7dWq2gdrbQTKzA+sucBMagj4Ts/xgJd/Uksb6sJ//yB7rcOJVKwAbsTKN1zxe
2x/GUcltNyb6pGbkftrczjdJfNjktJRjWrfIS1/JmuqEKqWJagnvn3Z8kTd4FwA3
sDhHoLccpzYIawLYbUfLjry8eXBowbP+ma8MPBT8sMqBL53ZKsXa5LekSERxI6Zt
2Z9wdFQPbPmpr9B9fZfuwJ+Eq3VgDhv2ttwL4NfBRedza5GbM8Vvhxs6mSrjqlbT
D6QRJTGBdWzxuTKwGFZX5MXQdoITEMl+pA3FwdYLlWZASPHc/EnL0k6tiwwsiT5U
khlqE207r3pyVRur8Gu2etCU0gvRRwA/MvRI253SbwW/E55b+afZPEXWKt+MN+ZW
1UvAWMAKjTw/RfwK220gmCBifY6u3uuySvmt0dTUcBkivZHLdmp6gJGuNN5Mf+xK
IIB+Oje2BaJky1TIR50MpWW23onX0m/3gJ0xdQcaQGWJJov4a5q+OsfUNc+7GmKF
3Xu8QDMXvOuvpkcxDvNztP0zIGMpKNd4aBjVVyCxH6enXRo/2W2P+D4z/tL6QXzH
KK4cBsuiq7EviXsmPGUIDgJtxF58sSpq53dJX/6Vx/iL7zgFT141VZj/xn15H84d
MHlNapsP2D+AHNHUr99qPOGerehrN8MD5ys9H2GSqTzfC7QsRONiqB61zgTs5g82
NNlBD4V1f1dmy+2hRAxExW3WMUMqDSNXzXDMUx3OU4Z3cPBnfb6ksC/mDkMdtyjo
+bqTKdtcn0mVSoqOxjOGaLR/HUQblMBhul2namODr81zmhgdwC687M3p7mXRIqAT
IuuBUNjwwR8lYQItf5iVvwyh5kxoge5lNXd6rXwpats52p2dUow0D5AJa1vlVGk0
wilEeaSR7cWe2oP6I8Fal8uDEFBBqV6h1uAI5hz6IRlFA0R5MN+EEH0b/oTw5qC6
Pi4zmo1ule+z7sVShkZaXaUf88bdO/mlCRVXc4VYoDnwnR2xUXZ+k1J/O/NPk/Ba
MVRCrA3TLwDVIzXCG5tInCGoGr/mmncrQmTyUPLUodZo8BzRFcIbwKzRaJ1Hxodc
sS4WiPYy/wBT57hFmtL+j4AeD7M1fT0TbcLnuCLrvsXQc7DklhcD1TIHGmF6kd7y
S5i4UsfC+FXLGOwV8i5LNdjtAQEK/jtFFZI5XJW1g2NaMyNe9xLU8jyxrfyDHyGm
QEMNlvuLWfoKyJmtDnXTbD9FloqHt9ODkahxj77oESNMOufb0xK1n5g4zIW/Zqht
Q1M9WvUkCDpk+Cle3Or98uIQIYY4Tl/XwHAG8lh0fS3y3+Wl27sl8fVPc+oPNLvG
bvkPoCvoL/BXEPj06/+jRGAZmEe0H3ItdxFmZAB57MGDtVjnYR9GBjKp2zQOiAkm
Sbct18QTpv0gYcgHQ0HexP/rtWUU+tdwhmyfTqgQlLEk3eC0cUmYGBQn/KE7zzVq
S43xoaO034BH7SltJR+YKL0xSzUmj7MOXwHnA4RubX+civcFe0OLpEtFgP4lLBzd
WbeCLHZnsurqvrQtfRZB2eNX3dM3goiXmqj4MUSYm39j+W82pbXIrOfpTw9uDdJC
XKwoHsw75DiLEYWY/kfBeqDFThxceKTrpXN5IszumfEG4hUqhCsMyRLHRDkpFP45
poMrGSyQc5MpIdoNK6tJZWkwxGNV6wGArG23ZHxMzqesLrtH4wYp6loMi9s97Cvy
+6hbrx14mn39qD2+zfnNbGPML0l/i4lJQda0JIF3EVoh2zv+NwNdRr4xHxZ9/eZN
mp8W1AAb64SM3t6vDk6Xj4Np7D4+Cd3sho7Fp5Nos1iivAVKT4Z1jqF33b8lTbXA
R2gX9Q6K2A0s0ewjevP35bYR8w0A4Tsng2rDWI6FFC4tU+s97w9RI9OfiOZGpGhi
ZGUJcz6gp6J08dpyVjG8vWDWE3XBJ2sepxplYMPTcBu5TrlTxFBr4Ztl+w7uO8Ig
T6hP2XbVczbB16X8cL5WyUQqhVqclkKJ57ubJhTqPn6H0BdeaeyTEmMz0XoCnppK
81/ZIMfzWKZz3jztOtmzLuz8Yi1/7NCVBUsUrm7GDhM801sjC1IzVz7sIJlz43ot
Ow3Y3OZQ2rkE2IrL7Dz25Q0S6xucKWhM7fYOsBz29xWlY9XxzZuY/bq7K92RpT+j
weaSMNN4IYpXWKkl4eiPvYjaMoy7fVfAquHTzH9SWdeed95ivBYYNUNj8+h3+09N
eroFhVToXFgdjeLsSiYDNMWVdy1ovzKxhXhkq7sy7OOAbsAmPD5xyCiLzfoKRdw8
f10wWXW9zHRv9nfV7BWlPGXMYXpTPDGrr3Awm8ET0Vx0JLpopZr+gOwzS4Cjzms7
uDqNBRHcRSpijWgUbYW+q9zDkPunVJYSXjFnOrTE/XiB/Wl8VPcroKHa1o9+pWIT
DCBFsDP4w8GoGusb3HVKxW8Ks98uJEAUHPBuaKpYEUPpIeYe4OEhhce3+HreyZaG
N9QWbxbU03LfyF2wcGNmV87WqiftWVrjeXyeYSzdifpbQx/fyuJiKci4hs6i9Csw
1N1tpKnRSBFJW8tYK2Rh/pF1uwg+EA9Sa4uz0rrzGJiLEDOymMieAe/TfUcDs2FB
Xc6MCe/QZ/zz1Ngp6Y4QO3QPIjaU4i6RAonmQ+Dc7+i+sQbddwcwhphBok9RW7Mp
IhCj26bQi2syFthUzBMsufcwqa9h50o/a28U97aYISbUECN7wfmjlgj883RmFldz
gpbhXlJrqAgAjp6RUIq9BXyyqC9yzuktWDgzIlt5IoyYUiW8FEwMbqcyCy6oQlzA
mqyfUo3hnIoityprlAC5tJBUxL+gbiZuG3MP2ex/4XuVfKYVKywI2Ue2h2xbp6nx
swJZAradg2RmHMxCx6utGGkhJAWdFHRHILRuoDel3GlRC2KzB0dChHtDQDmc0vXK
HT4XK8X7PsKAIoCW0QZIzK5+DLvICBLsRrjHR828LUPgT+ic9AXM93y2dmPdvUO8
qZNKefzTTvVmsK5bjzMvH827h0GRKwrPPEiFCpAbu8W6BPRs3DiGIK6F3FSw+jRH
WHW2yFrS2qA9Jmub8WPd5vYqVEmN33unJMWwfuhgLN5c/R+L/lJMxEJn9ui7RBjH
lv9MY1PBkDcKjQHs6HFhXZEt9esd9F0gwPwO5hFIbYmmEiUALDzFpfHwOqvpz9ep
nA5LQZlfXCPshI5wtStRUI6gqMG/w/z1GcZ98pYcNTsFIHM6h19hgVkfHf4VNfPf
6RSDZXVn4+RtsBiQz4Fal1TZuIKUopcbp/6V9aqBMSzaVS6aO5oIoSgQBSsuYcdz
+2ViZjFOxXHSY4pzdkwcS2ZBYswf+mZtDBDAJX0oMhJqqtp7SOC+np4pvy1iJ7Yf
hl+zE3fUuAlJ1KlGJAIPMesEXlFVtaYm1s2olVoKDoBmkKNtn9L2O/lOfvd5P4SQ
buywdOqzUCXHwsYHIC4qD/OkDaklHSJfbTa/byvGyhsP737zDc3HpW/iqSId2erS
fhps8AW1Y2RIZ7tJoTCzNbzXWOS8urI45yOk57jFlCQQCzD6pQfXGWogcUyh6d0N
n7fFW/jg5p/m6OxG+t6VVRu6te9kdDHnw4GMPVuoyC61vsp7SfRX9gHFMV5W7wMV
k5GXiYekRSG4CW5DZJqpH/VSRw0DM9NCjedSQM8JTfGukpnLhEQiL/VfRmu6p9Ga
u/zz+2vVN4yB4jRVQJSuY2F4OQVp1eEvigf7KBYjIBJ3wBKzCjfl9aLv2xfSH5gZ
b/creYoy6fymP+Hk5c9LKbkiKSqarxLAWR3wDMJJakeE0i96Qtnt8hCXUyEiLdPm
+eHrsy/wU5EkRNXWMYyA1Gw36MUGK5VI+2rQZ27X+jdOkcpOayG8rLStu8TmJMM4
lt3ZXeSW5Mpoq4D6uK16rrevq1Udrfm+PdOshzBdjX/K2rDefAhhivXxLeUDgLVt
9CugF2vJoCFdduBlqSsKqisuvrm797sQStcsdhlrfLNo+CgFivsCBaaxZ4SbGz7w
kqph6+0UV/LcJNJfUvvJacHZ6tbSDRbydJ98DrejAoZzkQJZHPW+oVxT7obF8BkS
DuW2SBJDrUIGg/K32wj5T2P+4Isa/SaWsErBmJYaRRr7p3WGGgF0UYt+ZKODKSd/
UiSFaOXpBK+BfQ4N1z4Qw3o4Twc4WcXcVaNF4YZZlpE4fYaAetQU3TnFc2LPl3uy
4OC2vLRPJipm3M3Yz72XWn9th9Qc3/+jVD2G2fm1ShimqXeJFkOYBQV923uWwIE5
fUPSDoLqI+8RhDCIQsC2SKgpRyHVYxsKjqq3qW3WcEQrTEFMW2Dm8ppcE7l4zdoL
pmzMA2hl9cHXzaFORlnrCYPSQ8ABz7Yw1auoQO/PlseoXgHRl02qArsVhpi0fsSq
ICjXPrj5Imi7Xnp4j8/YvVfiEFDOgeyxNrvMxD29bm6M0Eqf3mKT0TD1zjSFv252
yojxe+PT03Tc6A8hgeeDmWnVHDj07GmlyWJgssj92lH96MOx2021Ho/jjC/CS2mA
7R7EVKXKegFafiSZbdEHajpiZbjfuOjsQ1G11QBznz3TEAkrFUcKLnMz1cpMrj8q
e8cSXUdj8RaxNYPVqC+DnEPjsW3WHjLQerneF7yJufwgbjeTIIoIBaM9xyWgkhVn
s1NOdifjNvaIIcE/BBPa902Xcu6G3Wc0QwIahLgDWvXDDWRKWb3We2w3rCTn35on
ulD8HSNAEaJ43xHrpsbNmU0kWZspgqtf3GQQiXOyQ0mIOYSTTE7ABHGCs/4r0gaL
MX7Qp8Y4XmEVzd4Kbf72nURsANeUD6vJerIJuYly/2kNFjx6ZNAchVglz6adt8p+
CNDqerAWYYYlIxLKcBG18sLVnccAK+CARZ+W79kqesXJgI8MyZhup1l/wJofuTG7
5de57G6MIflMfuaGhJq6Z1PuUjSTH6aNTU3zLY/bmBxaS/RFObQZvvm6FgsVlEIF
ruujkvPV68LF6Z0veNeboYuAjh9ItDcZeMFFA7vowkrQppYgjpiBEf9YrOp8lGFW
zHBQ/t7m2F91+xIRzRyW0zHD5ki3IWmlCmh3drK+2aHbYt3YT/k0Bba1Hv7zzciR
qx7AvvFc6S2+1MNoTaZ+01zIB3uDjxAGrhA/Dj0k4wE4cH7Rr2v9wjvkW1OaMmCo
g9ZFtHtJyNFeyMkrhqi121NLcj+E/hVs+f2vykI7aIBQSdV2T+BHK3amXX2Nwg5U
cbOTk8wGTEYNKXuySbSjiZxaodoN6wdLPP2aqQxFhxBie7O0fbAB7qnq6RrW031U
MR29LJXjx+zZqx7L8HnH1kWjTlrv0Ji6rZ1ZmPJX+paUht6XeDwzSFigg4NubQPb
Mz7PxPiGRQ5UPhZ7rpGiTDLXjOmlKNgAqYZxpdzeCVj7cYgSKLG+7Y3clqDKwRRY
4McQE3ZZS4MxGOBtliFUHE5vPaZ+fmoykrQdSrjObAQzTI4hixMn2q4K0c+Grley
3uvdxnm9WA3M6LU/SP8nIDFCpL8qE6zemzEApeAdNs9YbtLZgVyvCdrNW5H8YjN8
IMWGmKXSjLzK8ZWRdX99/vC/Y6GMCB7xciLhhhnvBclWkoczcorH7BgBVkyApf+H
48EewqN8v7Q3jnQtWOXtgc2vpcEeXAC4DO7h7evGy5bNYvrGi+kZmIzIMpDZ5Z28
J+/uVOXqW3lSrNURJgquUu6PdRWeIrQcbYbrsmShXASx1FbcJQ5o4uI7BHYQYbbs
xFeCwr/Hnyo3VWAVhMqUBjeY5mfu/rUU5BSsvqEXVR0XfIATCA3/Vbq2vVPky+mr
P7US1M17lXFG1NmdXrQ27GNQEzLtRT5IuEDDieyAfcxn8K19TBKej/TdD6CnXGdd
oR4zxTVG480WDhZmiXA+ZcFLne3WaiAxnvB55dHn6SGCKkF8qd7tGHBkv7N5bbfx
Yu17AGwcqmnC9l7n+2p1CB17gBwnb99jH2iqfkcR1B7U4yPls6MXqrBFubqmtUjd
B/AyLlGe7SuGmNUyx5pax/YXgfuNH8P0hmqXVsE/FHK7gtO01uq2OC8p49HLzv3y
LmX2sH9WYF/Vq3sNGtKBvfIvKH6Ann2D8YYXqdsW1aj9dXG0TSVn6uO3EFrm0FlJ
WtxQrT/2brkv731FxNcPAXp/5wT8ST/kowLFuIt7jQdHLMBmQqhZitddgB7/RDnb
Z8oYCD5MFm2hta1pe6du4CNXgLia2eMnLI9i42c9O7idnWES2rQVPmP5LElLHo3m
SjLEAZ5vppno6VR2MS5zQWufMID3Dr/KsuNaYbBo8Mp/FeXkSI2Nfy5PWmGqArTP
Hh4S5XBZzXFCbYKFT1+oRkFpE4G8SaAU75BVb/+LIxXRMZpC+buFXM34Ft3e18kq
XKDwC7kP/MdM4Y+vsQgWi7a5rw+pOPG4mHiLcwBRKsxz1S2WmIL2BOfdXqqPDdOg
KxpN7g8KhwAfzRoNtVG4lllOyP2NVCfJWv9wx1Y6GbgOjp1+F2IxShgToJKOVV1W
Jj0hed+UQBae4+k04WEw1wvvHe8bdobbbtKsVoxJtWIAcQoUys7+0s/r3joC+K9y
bHL+6AjI5BLfIb2jbt9E2rwFoUqFvRuachqWtXiCvkZNWkJok1DmzST+1cX5RO0K
88/mHK/WvjIfFxWORrQEhpsAvDz/lyANo5gCzUPnutwQxb/vDj+iMrawpzZT08aH
5TvIPAcgePUZivYhLrjRdw7ye1MM5POA5Wdrv/uC3miGlg+nmAnR8KjaFpADA753
w7gU+PVgX+6CGx9npZcgeAup4XS/nxEGCphHtUt+cbSGFFNHrZempsujIcqULV6c
wYzRJG7SkPjL1RFNrJjHFmAEKj6rVLfzUElS8kFSUkcUN9SwdS/UYAOUq18AN1qi
Iw6dSB0LzuOBbsVN2zptZpSrYQiIoYLtZ4yZqnV9PMc8cnuOq6dXu+/uryUFrqZY
AzoQjrKa9Hi4Z5oy9yOgQ5QnFHN9uRTuMlXtpRJ558JTBJKYkI7ezDhk9iN9eIqh
A4tALpiwS4nTtfxQn5x0eoJmc54jieKz0v8eyfBo7audbfO8m2+PT9O5S5fumg6H
UdGqOg3CuqfLOwjDgJBxKUxniZzaiZdVdUh2VzaOT80xnjpYrY8vKdEgZ1Z53AFd
BKQUw8p9wxXsoOiCr1RcCXIMeiWeeJRXkI7VKGhZzT0W+zu7I7Sn07Ti2nYRYKPY
+BZ0HC1vWGsUAjVXKg3nFnmUJO9zwtYxbozBc5K1Y8Ho1dle69L3ayEE4C65BPBT
JeFMHwnJg13908L9JXPvDCagXj+64Y1geSUOvW2r3IkefY3pY2c+YU+hvhC9hI0s
3tOGAdZQ7PmTxc5x9/LCm5i2CqHkxk5YFXKM8ix/2rC+Z0WxbxfYfu3GYRUGsoTg
rWNGM1/PFZizwob3wgdsN4n8oNbOp59Ilgjm35QZF02hOeAJtX7Baem2jwzgYgkR
bNhxzYMi1BPiyLtgPe5sRpHpihlUx6J35MYE9iR1/h2ss8pps7fa1nrc/cC/jb0b
VrX3NrtM7a/VTUWMLAIESWIkhsKj0hVrkjQmhpeIGU/lP/W1Q/ZnIc2RwpiPNf2H
z6P552be2sOYUZCMiJUGty2ag3tO9GtdlaFJalKsHPFApgI64a2X0oNFZ/OfhjKN
gXMs6gHBpOJBiMEfr/A8kQw03GJTp3T3UlIPrpWAcOruovC+hNDlzyl7CE9+8+4k
7A/torH69UnBoc8b5NhTVFx2zgOnclBJwT7+tCETROodGAF9nAzg9ZVMKvEgh8fF
VeGjnVaZvplq3lsoyYkMNT/Th4IkhmyLELc/+Xt7+MaVccgs3AL2g2xuUnuqoXlg
3MZEITsLCozl/GttqsAX4wHPCV+Elda3tB+RBOw0Ww1bE92BSJgzhw7Qp1+0gvVY
31H1/sLOLDnTk/KT6T9sXte3RMUPQkZxxbX9xaxjuoQMhtclbE6BL5T9jNBugEID
irzLDAZMuj35+vUX0+dPbMaI70CbD+TuVbraClCafdsGHIKD7muB694Nyl9cKZkU
aJQxuG8Ov7iZscjsfznZvH41v9lg5BbzkF17SC/DSyohO4WahKPOBFYGpWSSXSba
+Y0xvmnas39qiAfAV0MIGkGxQwwPhritY2Esuh2gRVmx8pPx03RxtV0bMpehOH6i
8DSXq9YRFrz9I0b8tcGl4c5/Qi76KvDy/cvGrDd9UdjZiXrmUa6FnpITj8qlnULq
0yOQD+4YuqZYTAi1WxEl4hgxBE+Q+7QcrpH5gD2MKlaG/JzIB/5CdERBeCygZxjg
fo4KkqTVm0mD8iVzkGof0NcjJQ2/zFKGRpgPQDEr4Y7EcCycBmxBnTRywF8gsvTg
2d4sLlzXA59MtXJg/Mby29nh3boR30PG8hjNIvNokZdDSwfw3BZSyWdXwF/yzEF/
74zx5oAeVHWZ98sJX7yJvOoC1PjnvPTaZv7oNzNvq1y8w1pKlSA2Y3J998YKoZIm
xMUlkoDWiCaoTczN/upF+UOFUiOIAZcIKZrJKKh/hYR7FyjUeBNhN27YtvZinwnf
JC2spG7ws8at9u31gyjTpqcVvqTcN1vHMzWufaT0ZVwQarvRXHhKbiqoEaYjvAgA
AjkOJDUXv4a65X9cuD3t9ptzAtSO2YEKUg0i7jNCTnQRjo/PwbbltOo8NlA85Tgm
I0KVO70w3wu5UAkTGG3N5v+/5hKV524R8IyxXBkIMklYiG2aa7BqSd8gPHmvPoka
OKo6Avi83jHucYUz0R2WWukrBFdS/ycJA+BlJd8msb997qv1oxm/A6RTlba4WiiS
BMJT9qnjP68ADQ1iyi+/ghQlr18KXUF7I9n56f6cseNl4VaHOENqaA7D4sQoFR04
WEbHrt06xFgwMNaAYLyPnc+9ua4WQEvntVGr9xvg/O82o3Ye+Dv6xbmxsSiKqvGL
n8W4szAJQBG7+ZdxQHdNveqc/F47jPA9t1zqvNAiHBO0JVn84Hn11Spw8HwO0fIA
0CP8Mvp/cwlkEc/8cbckOuIwM1ddaga1y6G2na6ngeNKt1CYdNE96rCvU3F3DY1L
wDqEc6jZo6X3ZAmc0uVtkvGintvGcOO2ILnH3ndb4oi/CPEDtaxwrQEyEGRVoXSf
wTNOxZs9vSXJVA8XIczxDOz7HGTaHjstDewiA5Z2aR2Bk8KXOqeI8ozDudkkgcs/
7Uiqh3v0PmrbXngxUICHuxBMJ1Gn8jEAILiIpGnSjdAsvZ6O02IufUrI+8lmCLQw
LJaXIiaGFsUNIs5RCz9M1ATrkyJvJgVGSKb+cwU/MQmsBbDtFikw9/znrFtH4lUT
2ENOvAwZztwIgr1JvJSerIrohiYCKB5XxjspEr98b48u4ougDkPlR5mAmt8G+ru+
0N6l/T3+KO6ljUOuKq/tY1zp0z09EtD50NH8gCZl23dZUU82SDupUKjnTMXXwB6y
IgpI1Jg4szGCvLVyfyhd6kvjCrtLosD1sbrzDaIKmZKN47OYnoeF5l/FAInahlf+
fViVb1UrTCu8l5LgA1oaru54a7Gl8LPZfxsUGqH+TBgR46eXbKydAC4Oir9LbGuN
8QT/HFFayCxOys4Xui6HA3G0HMKAwvcd04JgBn3yVshUTlRuTbMdFmU8iuFv8ELX
g6zXDLRl7Dz3hS30d2XvorfQttdxoAg2RXYnoG4db8VPNKFMiWuZh8k3NtIIn92M
MfofB7mPsa99r6dxAFDi+8Y+NniGqOS4+N29N5z2av58XuIx0StH/kX6KOkba6eX
REmso+W7a0TcFRKWDoCW9k3th25iyfqK5WUh2gG4MKqvFFWqrF2HNxO0FMFsgJPz
M2TPiQluYUlf2Yx4lqWrQyzmO3j3hmP9mDEV5eTr8dFiopCktxYvNoGb6VY7UYo7
FUsM4C9EqYCbuEH5fqmfRQHXwk3fZC8FlWT3b+77R6vCMyWYmjMIO4vRNbLufoNK
m9Z3mokAOfvOYIBziOD5RzTUThKRXh7vvKb0zLAnISsQSX9e55CiT2Ufpcl1g+m5
xLNEr81qaCN3EksWVO6kfDVfKrUMT4lPm4ZalIt7+MzQKzy7vog/840cvu/cGybR
W2nTXryRrV/srfD9gXLI4wsJu7Od9v3CQkIsxJv0Eda8bisCHCqkWNlr+n1Ej3+K
DzV6PVQfTsDqt1/zI29ODtzrXDCXtFizoKMBJtG3ZwnsbucBz+GXoQBF6Aq7Juak
1EziQBYeiJ/9kn8wgWnI6KOwbGfXmTMGwF/snHL0EByd00a9AAIuFwVnD99+jfiz
V5BmidldGUJHRS9eBVzz8cO8w9ctEScDJWtV7mgOfo8Hcr4OZ7C5WTKQYKkqUsl9
bly2PPS3i6LTZtpk0ZehSPUra37AiZB1m8erdxUnDSrHn+VThmzsXbCC1lZQJ1CI
woq4wuoOmINVdczZHw/gq5ehlPZYZk3rk5PHsEl+5fLCKTNwZ1ui6MUDFmJS0U5A
DIkAYHAa0s+w5wgLF+BZZ0KsfY2h51u8P4g1MlbXUMHVRqUpVhdEqFsDzn1w6fGw
Kw1B6emrq7O/CJ2axWyuOwlL0qSAjNJra7DfMT9z94mvcG7Cx76oZSFGt+7cMWnV
4DmfPPJvqrBCRedxMZ3Nt18r5bs8sxoTXnrnRlXy0qgOTP9Ltw/Jx4veL3IoEzx0
D/f8cJ71w67skTLbPbZ2ekK8FULJ53NJiBxGrvXD7QHG9jCF8Fwkn8/2cr9KLZX4
dtXkHgn72b4zFm2Q+0SzTyJM8vXoZmQZ8GKnuqqS4PtX3GyhRvf7FT/bntvoNn3a
hYn1Up1Ftz1CP6OutoYZQrY+30Lf1QiYAT+JbkkhHEwDUSzAEAJZ9NYS12Xw+x9n
pTmcGKnAo8L9PFB7KroaZ1DihG/kwaQmAlzfdGbvVu+BRnJ5wPY5DCofcN4KnfcP
ExRUrZfq6Otiwo2WSdGYzK19qLS+IbituPl0H2Tbj37Ol0LvccbHsgdNg5nf/bwu
v+rTC7dx/MtXAlVbN/n6N1gBSETVy35K//Mjy3dyorLdj/XBJh/VW7e2kjCbr1gt
XgS6w4pU1Q3fAYWTh0uX0Jwm8k5nq639slg2H1WC8/8OZSpQvBEcO90qZgmM3QXu
Gh03oiGvJDFcX2woxfNRzLSMfzG7o2PTpF/b2cJPQc5gTjPCEinwEPC2nXq5Ilc1
J+brYMGgI7kUr8M9HyDEQe0fBXWE0TgVEMzQdoPKEGad82S84kOD3M3UMUt7SfEp
Ztr+6Wv4R9SHiqFEgCA/xaUv6SiTn9jFJSWLy/TpGkGNQnAjJr0kMrcnwKYy96ST
R2639kMABuaBxq7HJLi2EcTUNn2em0U0BQnmF1KEpkgCV9QcquN/xtU4XMUQBj++
CuXerQsTdgoLECLdFDS6RT8H366Q6ub0CdybO/3HFtpQfUjDe8lp7trBRF9+V8Ol
axy62gP2b2QPqetBm4mwvWLAd54Y5l6ANqdImarGuA3/SHf+8fYqbslQGUUIrrEP
HULsW+rdEXIKTgS+G0lj7BjThAUW8Lv4XYyjmyvtJ7L8ShkwVBJM7uzwP4sBZyJU
8efue5jnINtsmDKkPanqRwDMf/HFo/xwYMzXF/m445CjmkB/rK1aiPEB1iW6iFNe
RJzFlMu7OX5L/4t6TGUFTjtNrtNqLofwADQCdx+paMUw9pLsa/rGeYIkmCQim9Nr
oBV8bbE8/EeDWL3zzJQm+XVkYU0O/E5DnB1Jyb79UYUaHiySMZta9WKASL9nBTPO
j0U3fwGmXPF0kINSj/T0hztVtkR5z8eLcP//msPdVnubVOP++ObfYkODsiZEAreO
xsoYAZ4caKVEE5y5AyA2ROREnzatRn6AG+IAt4/ALIari9+MShmPO62PM5wkY9ES
TZ8vOCQslEWmS6sPkyEwCArWgM5yjFju+nO0jFwoASdEc2jjBxkZgcyELOWVe/Wm
sfPsnauRhsQNMNjElLAVgTfLWMZBzxSVaJ16t/vGsnKBaPJh56R1LoLTD/hrrJDc
0Z7DAlUAMMQ+f3V+mDtQjtyS/Myo7pJO96Hw5hZBdvTU5GOuC5I2XzFBzD3v6eKj
VWtWn8J0gvzDtAqa4MiqOA8dURNITFFflHAK5Uni0hQ8dWVEFAnbPr8c0H+8hIaY
0oVTpck/Jav5+jhiY0adhr84zBb4+iz3upSswjlLFB91V2HqFP5VJeeci1AS69Gz
eMThexpuu3s1F9k6yWlxIZWK2N4KfKpvPY37Tbwqrt3QjrJOD9WUxLXjkNaQJGg5
p30m19AZg7LLt/2P5xZhl7joJ1G4EI7nDKnzOYfzCthA3n9FmdFZPBgLpI+S9mS4
4fgPAZCSlpPilt/V6/CX5nzZFdDoGU8bAM2SobpWEWUVEAqwzCJrNOdLN6U92lyE
VGKXDf++g89SQJeJ4KTHgsx/Y9jjepcIbe2Yr1pOF5yD5x8igj/bkHUJ2HlKdOXB
/1gl5w1wzOshCr8qL/2aVo7lk816ok1EDPJtyI0uK8PPJ0N07LEr9YajRB0E5jcw
FX9hE4fJgQzn+PCQy1YcF72SQTuI1hYnWey8csgI7RYdT4QHi1OF+BKoUvAL+oZP
V/trcR9tYaqguz0s7wge8mPlzE6RFFf9TRUDUwlPn45+U7Ug5RubHMtiE1A9PYWD
6cbx/f/GgH9d9rNY1RSl+LnaYYXf6DLHM/AcSeEvWPoO4syzdWBK3jUb+E55O8c0
ERwqMrlCAba5JxjBMwOZ7CI6ca7PAz+dF7RCzbLlc9oK7FvtBSuuuHrzdg9iaPtz
s8AXjUIWdMSJd/pKLCNphFLXKLtVExElhZgdLUSyeyMg1qUbuHrvFk7IpAYZuu3q
UUdolP5KpqoWeHqYlztzi1elDluZ3O6CHSSOUoF0JozUbqr8yKPwx/qObcNLhxcG
t1aJYSavYqG5VR+VkB2MBXyfZTM28WFfOw2AY/sLSrwpJyGCDBVLDeEp6YEd8ezj
tfx+ti73Uab7nKxaJRii2ttfHWfPj7ifnmMQmqCe1/df5e0HqrG55HRHxUEtIBhw
TaKTz5xP/MjltvPt0EjOwNb8b3em8pfCfPjya5+0+SajpfgBCCWRdf61H1CzT3/S
546Ihbu3nlhPOrnGFZ5YmvIc1gNEYMWjDVi9WLR508fYBi0CI7FzdtIUez7EDxDK
AYN/WuUkMMqDrp1gruTqLZDm/uVr1dXSbJ175z5L3yzbtHnkRKcWJgle5gkOCEUr
g2vatb4WPGpc2VBJZFuxU3Ecoj2OjBRyRy3JKoGqiWlRtg5diU70MNP6mGp3/H/t
DM9MfxEDU56XjcW0EHbq1BLqDy7supePSYVaMoUsHQHUHvOjQgcXNOQgxGkUbDQ0
CuNqWWu3kEYlSyRC2Lb9z8ufrDMi+Z0TaKeBBwy7XA5YTTJkSLxAiw0qSQqSu/rj
ZEQ8jlsA52a8VRGiIT2SvJXmAavGbPPUvLRncN+nBF2KbLLOCywF+aYF9wL0jpPp
iBW0TUB59l7M5ldT0pAoaCIhKiiT88MEkfQrA9/CixjU9o4sXzsrRV9mp58vaj+F
xhllwxHDYDK1PaAA8gk1Se8QKD3mR0AQtxvTqwMEKjgRjlXyjpbwvMzhh0lnuysx
yJhBfFqqWosVgX0hdavhzrki1T6h+g7ngl52dYwrmAeRTV1FlBbZjO69jEG+RrjL
wxmcG8/RVF2DDHUsy443dwZfuJU2Yq8T77eMLn1jZ5DNA0XQmpfdfhdgqwRq2DiX
dlNvdUESRT9aU0nqEMJWWRFSDmhb4jg/41MtyFKC3oCVTe9Xlulj16zS2eS6gI/L
+sk4AN05GQWMMkpqN9cLaOl9RYF3kmT1RznJqhZnCjxgYdRpooywtcXfBXW/szvH
ZielOpT7gK9NfNqGbljac1I02fyVjDHJW8GjlivgVa8mO0LCH+cso6XY/ALrQyyU
fHhNy2ScD0JwQxWLWEj7WLDOmmarbCrjB6PJZyEohApUo1aIhgExBtZyjdOUNpqK
XBfzcYDHQPBgD2keMOv0BTM5WXjaDRsTqgcG4mDIiaAfTnCx2+NqxyBiLCwzAte/
gCejo8bGlbcQvpW2K47OFiECk8ec+PS6AZTD8V1JEUTXF+6GnHDONwVf4RYKglQA
2sqk9UPacNl/k7rn8ry1v13d1MMxrseTQlQqqbsmzOtbWvgzkiXMr/hpfwGAkpjf
Erls33SAdn2611viiWL3oaK694FNO87kymTdUgNascrgPtGfcouTr0wWOEYbqy4D
tS7oTm2eAA7BIOYQqhv/isn3t66ziv216E1igSSIrN8fyuXaVrSwd1vqhXMhQHep
UO+tLINELDen0DMpPwzrRdf3vIzD4pp3Zmw9dqB6J1CIgnuJtDIrgEUjWTq2W8W6
Cf+229HWvLX2ikQCGxq/XNf64XcmJsajYwDKj5Q/vz/UXZvRfjgtY8OKchfDMzvk
JsJRjsRY+nldqAK+1dvdyy5P+gj/xEI4kcFSxNJIRtoLPOZ46d8fVJww9DE5KKUd
QSmqFUbxpKEINkrAkTcpGANlH0HrFvhoCrUVjDa10lX4nHKIdzCdns/0HqE6zgk8
8Kd+V1aPJwf+mJB/GkSW6teahXO+JAzizWnq8MKMmx1nw5oEL8qzM+yuymHKniCJ
TcjlqmUKBAtQzk+GTilZYYC10lxAG8gQ0tBFhuHpKzwWij4wYRYysfEHmsUbbASD
UH3sM7+v6zfeEk3BfyTmtASVwVOtvvYXXg76UtVTfepCyYu5/c9QzpIjtm42PjOZ
Dwz4+pr4n5Wcr/bwx7ycWhO/RF5wSQYxW5iAOHszfnVIBvfKqNbbBqXdcDR4A5El
T5QZcbIbWEbPAEM7kMc7J/bSKrqn7+nMO+G4FLMYWb6iQx8A2RYWUcvm/Pg4+9R7
S+1olwjb1zb2JacZE6WAL2n3C4YwfCsgVsnof5CSyTa9kzabmcgiQGmAlmZS4Hl4
Bibh4c1TzE+owLjIe14FSEEjcfzLmEugWC5Mc0fAo5SCgwT/C26iA8KztXBDgGTO
8td7jIs/QgK0jECSovroZa32DkMZQ0FChqmJht/ODnwICFaBjlAIG2k0bVbap7KG
DTfEdhcUrCrCu2OSQxDH1DZKKqP6uzvQ5G83Tu/xqoyZaPb+cApH6dHnIT/hkMtN
+tHzydfTAX4Up/x7TsQ9Ivs/UU+/0pcwbJK4Dx87KVf+lN+81obxiSXAZs890Sxb
ng7zbA3/7HK991XD8sI7/79wJ07p4i6V9H2fWGqXT5KI8p/K4GjlO59dJvM1yTEf
TxTv2vlRxD7LyyqSYfddp1N5oCckyC8RGXsCtmuaJDtp0wGkS/OEstVP3MpaowWi
4gAIukKbbM2Em5TilndWV8Vaa+x/ltoLkcBGtd4sMNVpojV4IlpMbwEETPei67Rl
iDa6A95gDIQ3hCcHgSez1ltBZQUd0EEZyeC+mTv4zNLKkvKFMmxeXNyaQwQGqzTo
nqAQt6ny7qoeEEczazHVC10CINIw2EH+yUJr7qVdc+Knusxl6WaSEgXuPSAHljZi
62kcCVn3jAr+5qjYqrwd3XGIXSr0rU1cNQITlgsrhtc5wBcP1BFXOFZ0XVfPGziJ
j5qcfqv0MyBPNhv2bPpXVDCPWgRGmquFbOqXULkiRgb0qZ62czeY2KlvMtyG65pE
aF6maSb2hknMtgdU4MlJ4zbv7M5FAvxbTumrj99sJyjiAWo0Kc/4isEuPmzlGrL8
6CGdeivv1qQ6n5Y++ixXfU2GfO/pn8LscFznT9AG3TIXTa+990HtA+lLpt1zvb0E
Ffl1SQAS5Ym4chcJgIW2HSLJ1D9y0SRhCuFEQ1FJQ35DQ/jXO9Gnj1FY9U+KBwn4
/1AQ0v1FU2YqeC5q6t2uhEisyE6Hb5FDffvrCnuiBXgtjUeBKC5xLSn2PRx67Mnq
qrYEum53QpOpsVh/rCTj/y2tLk0Tt+pRAUDK0cDa3T3KkieBbChGoj2NCFyLPxJz
UI5DMUZ7aUFPHdh8vKNLzVRD3lF5Pgx6nvGeBD8vHrUD8WDlYH8kWxAvJrIYhiIz
4CzJw0mx6DZTr+fPEvMIA3VL1hltsb5v/iQYC+DM617Bdjk55mfIZFHOIdu/fk2P
FK5fITg0cIXbQbMFH4uNZJYIV5YGAZ/43qjVOPP8YwUsiaBd1YqLcyQZcm6zuBLL
s3WKuZXtrzUxDldhMo5wR4gthX9BuTl9X3LvkvebrVp3xznwTTYK/G61uRlyzJ0c
f7uYZdKIqWDsfAbdHVgUhxXi0evCP8bUv9P4i4gfg/LVLoN2bMyegd0PkE1lXOhz
/5jPLh8kXBN7vL2pNFWeIHjWsNf0gAASyN6DhdJBvBPWTgO72danoCXdfccqJm1r
nVbw1db2KZIwuHjT7FqaocAoM2h8iAKhy6RVmOz3vUTZsDkZzSl04f49HLZYEvzk
ixAd+jjOBByyxsvv41wxyaML+kcvqPb2eHotGnkoDzHKu4WGN1X5JzReea8LIi/O
n6mqnh3nzoDiK8Pw1TO4i5wJ2p96AgDVKAWfYQtVctsk5nHhsdlbNR3RHjLY3Li0
OYBUlLaYZGtqrx0S5FAXPvysNJ+vt6EwnFvv6HjZbgVGUQvEA/u3HNHshWz5wYIc
rWs4/amlITujRjTTwiFj3omIoqFc1xLZiBzSa3zxgMx8QbM3srTJevs14Lc+VaZR
LbXwrOHRUKcfVXN8fNczsySJxZ9jtM7fQgGwN8N5IR1QDbXBcgWHUaTF+VP4YKAl
nSe73xJMSsHIk8Fq4N0qEezDTqlqFRx+TWe8ka9thZA8BG/kx0VOY2RR7/QGosB7
RVnVw+O0ID9+6f2mduJzEU6Sh176RXlVzLeWYEkJkSP4+ggczUeP40B1fzXuBXCZ
1gNtgXIYi0kFS51fAsQMti3AIdj/gLU4tHAK+DaqoI2H964RsGiKIl8bMknOANUc
mybxIm4NkLViEU+QFRPYXjiEIKPC6gP8fERYEjg9Jr+CPD7qnIza7qhJBoldar2/
53L7zqzSvOOYPcYEQTGnoaLyrZ8wuazCZ2uM+wD3WfRJPVcG90BlJall5k22l83I
QEuy+zU2h712U9uoacdb+8G9s4LVaikbXvuISdVGQicuZh+q2OSmmdIdOMCaq7FC
mowpS8wZ62agorbmEsYlEg41QJAAyVMCgjuwexNEia5UgKtx5py8m/6ojxlW8W7h
0pVD1BHxKbb1rrHbbzpj2buChEVMfYTiMwDgNWVg+6HclVB6/EjdLAjJqE2qcMcG
FMCIDLdSV9L5mutRxLLw/OpH3jMMTN9ZeaGg93TZ6W/2OrAJJzahjUaLiWV2/WM5
PVZ3iQTqDIpG/gSoWmaQMHXBuArbJVDD3IMDO0XroY4nO8pktOGsqzTRzgBjvMR/
USrg1bhnyHg7BvhLtOwQllfOKAOTXod8MPpb//VVUoGxwP5hcqAImwenRktPN03m
UumWEXmATT4a0eV6zasCkUAbck3+Klm5mEQLzAoeZ3u3co2cpnE0Z2YToQUga0IN
pybgIZAmQFu8BMT6/SV84O0t5yzu4hBGds83Swt8D7QzBJufSYizNMnEAWCrw2BX
1wIFxLgoyjLerDWvDP+4lxNLYC4Quun2GH4ZiXC/2pejyN9ZyxftT3qHP/rrgFmf
6kmaJZEHINKkQ+hVEmWm8Conem3TxP90dRWzKqvFAHcCIlAiW3wSMJERlEUiBCzI
umhnUeFGOzxQ0/fuLT4Yj3vpYBaNLG+5NlBPdyEJjsmehyP89vgxdFsQ/7/2YObB
ZmHRM+hd0fnARsWO3msPpFK3ABEzhQweVoMNU1zpQdiXGpMuKY//nG3f8642Ce7Z
TFpr1d249uOpBjoXrcndgeTeGedwVvA8XHmmKEwVWoSmBU5lI4W6DOxYaTm9w6f7
ck/2DM2P3NMjh5hDIJlLVKjlNz+Yu0GG6Ze02iIvohRpQIzEMuGPCJtCmD2na0If
eiQsw/zznvBgTq6Ak6KqxWkbpUPApsVsECZeB0IeN//g8dqfx4XaFSGsNPJzxfg1
lPvZ7u5A3Nq8BgdpBFR+LPnHqhJLyUmvv4W45hjlCGdI3UpJvmTZN9cEY+dmss37
HKqVtRnFuKPXAGIX4daZUFVz8MhWPMFUDQhC3Pv+qi0wSQHychlOjeK1kMQw8jCf
mmvuBmYKb3qLl12p24+XhKOSq2yZ8Q5mVTlqBNEwsPenOuoeS+T7Sb1cSOCMacym
NQHFbq/hO2CcE+c7CaUfRGqhbNHAD2YcLJmy6lO2mapqCsdCuubsrQOA1zvngKSx
EIbZvZZsY34EMR19rPEyBNmK5OCtWDemS+qaGjsKbSRFyMuoxQZjaAGVvgJRlmsP
buyBSnflb89kUZZDxvmb9G0aTbMz21ohze+5KZTA4+WzLuwTJlpGu/1EwXPKeakP
Ys0RlgnJm0ZXf2LrEOb5MbdhRXEQR/2J4YZ0oyF+3eTTJmWDJPzYVhCAVopRCAZQ
lFyXU9TaILbRzhcRE+DOoyo6b/zVpe7eiKfMShhsWC4MhHzqAaRGmJdNVqI7iNHu
cNcagVZZvz0i1DgrHn3N1+2I9G5ZILHu21ALrPDrJwgfEMj/4CjYUhjuHPBiApjJ
wX7qJsKpccnMbuYaym6BcyyunryoUDTLzw4NxBFeZlwajaorjwZGhHIoD6mk46bt
cKJaXc2FfdyGHzTc8/wZP4Q3UQ/LZmta5sqCm/nxvSMxO3at33aSqNxTQQ+kbzwj
WFnBIGArc90pLRM13RIvrDdn2AQFhIh63Eq40GZ5YT8JoVGPMAXy28rhI8bYASYj
2Ilr45r63LhGgOS1MVFIFd/QIrsXUMsHWxygq9I7ygpdaobV5ryM6JnnvX1FCJci
Z6FGIZT/jeOspG9XUuet2ZFxAIlTJvj+yYPdv4aThvn0SI+M6VVsWWkcBs+BbVKh
Wpywyc6R8EDZbpndcxiRcC7WMA9ZVT5sXZy9NyrQ9m8LFbpenRgpuiwTVfNUbiH1
7K/7NaFwBM4TeB0U8TSn3NNx3Q1Z3sBX0+qJwbLPbhalS2MkpoHnvk6+0AENMT33
juUP40LjCJQrbbVvNP2XbgImSQmm7mU9ydfUTfm1xfjDjdgfSzUfVaZXseIeOEaW
UUW4iwfjE9s88+5tTm+eOUOf8T+OppjvB72OjnVPuMEyIs98yLhG8P/QUISFHuGL
FD8p8pPRQNXO3R3xC89UdU2rFSXa9+Iz4vKyTeupAJ6AIkeoSbTq9VjBzqU9Z8Km
pcCzTG26e8HaUxTJGwBnmLDIQTVERZ6b7KzArA9LjQs9RDAMDkkOxd82rqmBUY4U
KbQHlgkaP8xryitYPmoiM8B2VMKHd2v2E+3eLBrc0i6n2O9z+vGp2uNB3OKQhJFK
WlY7V5AskdImTMUjTRHiiOkPAE5sBccNo8kQcN0+m/NPMWkKckK9oGOX+Epxoi6v
kbVRTBB/dYl0mYf89Eusw3pNWawQJUQYHcn+Bc/Y8TkLEUdzqwxVMI8Ro1gO6VJu
9Bp30qqarO5pkba6KiRkCAxjuSfFjYcMCe94cFQC+sw3yx5P+0aHB6jJxbtHOw/2
AfHo7wqfVSZ3kQU7VfhVbCgWzC1jMbXoi7MrKleLkZoDoAx9lwzmBTuCXdimGsna
HxDu715PrLFb+ZhgEKFBBLUn8bc9K+yX1r7ptGUSi70x88NJo3t4VdvyQMa7/7fC
JPzYDXR3uPCCBbsKxRKf76Q0p4DFo2PaGIBxJ4xQFimW1OHMSEgx12QepkaPGJNc
UPEUiOZnIUdcgi+1deyCeJnk4cu13BCD5BQYq22ug2RrLBeZ86kAoTLHQYgFBs/3
QADCNtXqRQXJuhOVzYOPOKhPbM7P0N3geotw4pSNcd7rEJnUnz3At8pd+CPEbVVv
U24YimRIjbP3y3SpzczA6hidSLlO+2C+HRHsma8yE5pD6Om8i/ZqUGNvr4PjiG9Y
VoHJ5/R0Vto3djLEK/CcE8CdfqXxfTbOopKQTGKsKWtb6izl91KVc+weUpFbigQT
N6RA6GRNuv8boSpjWszQThSzZidK8YuRsSRQ/7haOpqLifqWUV0M3HzrTSmFlBMe
jBC2ctzej7YgrO3MlSzzfeTYZK0xbY15yBh9256ELy3BJaaxN5dK+3vKvExLxVax
XO+6UxJ6ZEfkPFywrbOqIuCHHJFR1m6doRpBQFys3kQspLy9n0L5KbnfQGR5/HCp
Ihf53cZSr9RSW9i/OHY65EwMnBwbnkiSdYkU06tLI8boJLbE7tGepKfohjYANsjp
9WqFP5bXiPsFpimUlvdOWpB8ei9v8Pm0pSV/TguE5ZLxaULhZDTUvqXMONlB8gOg
fpXWF6Qo+WkHp7hOvOV1XgmH1VVPA7z0lEHzG6/NP75bziTfHP1aSUrx3gn2XPcx
YY8dWYSwaBM85TKwdlCxxQOiTACCnI59OuKCu9WUxfd/S81+lMVMubMQyDazV5Xy
+3VKRDOYpe8vZtzi5JNqhvluV7ovwUVWTATP/jL702tjk6KFqP/kPaEsftkg3SYK
KvkyZqYD4bwhoeYjmj6MKw7OPNiHVerQmb2zRrBJq3HrySlirTLQMQeAMOPqVUjc
Qlw1OnzwjtT0TZlGdflRUVkh49VcXbz60r8oTDsXNM9WC3FVi1OJOf7Wi9sn5o82
SntsfeZpqwUb00jk/IvS2WVQBmltsC1/ZQluAabhRfOJoGPLZ6+5djTC0QJ0D8wI
wQNEmahOe/4Ah8giqkzXJcXZLQ7bEBRY6dj7Nkl318lxZQTEAinhiJIWAyOGwqVN
lBlrQIEN4h0TWwxh6e/A2WEiOK5Jb3aEuSkxRh6C6rEaglboDeF4FNmW5eACdbHh
in/g3Aixi4/h2kYcnMuBfqK3YL+smBE4R/AjpwKZN8cEEK+5/QkMzxVIlg131lAx
X9jHuPsJ1oQntE7RFb0Q4nJwAuTUm5kGSRcHtOIUdpWMjKtxCk3pc3iw+7EReIxj
QE8K65lqBm9dkc9lzzrWW0UFqmXFdIznKxiy6pjctBIchcB6AmDanBsCFuLQRQJL
m2YoGF1/pz2wbUZQHz/8MngUQ6yk/WOmtOAw4xePNVHUBxKwumw8poklDVVonI9s
FOgXmAENYg/3jRvzN/6J5KKXf6mQwotPimDhNmpTsDS8iL9PR6PmXH3ul6rdYW8J
8xuAKf/nHmhM6WdUR0jzpOe9kvS4ga7MkBQ+M34czBiuaNO2xkP2vmi6O7OX5yLa
R5c9Xgpqqc1zof6K9SRjQsVge3GJvf7pjEjivzHr5KPrbVPCekisWdPG2VvjSsNY
aF64d2q5jF8vuKI2J+6mVIQXULAZFO/+hqoSWxpKfDk0suJLj/rrdv9HeE/92oGX
Sw5nzPemNJwHMsbIMFRMNwBOCFK0sTAXvEaRNaOj2vQdXMzYv5V8nrmlUNR2S5Zj
cAvWhdPnaqiCyDCxHcDvH0pdOblwflq8BkxEtC7h4H/HxUtHNCO6MW7Z61mglQh9
k/zXccpH3H9vp1AKWLj26fE9gA7CODzaMaIpyJyco6yFF0njzXzL9mVrvWc0AYwE
sX9g8pEjFTZ0xM64rQu/uhep72L93T7PPR90xrx10Xf7pdqEaII8woX54YhBsiVD
0HxrrliNTVKjTgRutdnaNE/JwBH9oXOq+CDrDILjg+j/KfJBkVUwqePu0GpZODtq
fK50jZ0JbLvkhnP5LcVHRa0kGQaX2qum1dWhl3HLTlAvHSLQ+KQ4nzN9RuiqixR2
KL+W76wgWBRIAGTPurkZ2RuUxyZtgh2JqD53DH3FHHn6lUYcnzMpgRHMND0T6emm
G2p2WZjeCUPuWfbAEY/oX4u4f4sHFGN+Ip0CD6iNmvpjRC/B+OrKfWZYsvAutVm9
MGkD4uPoux7QHcAs7Y3CAW2zMvHFepn0GxdqDm24HESt9HuvLDgjcyvQ6p/iDl7R
MGMhrIkAYWKq2zjypUh6BGhCf+zRUkC8BinrDGObouujbKS4bnGqyOnojcBIZN05
K/6rX+DsizGXUHeyw0iQC9/nt/tL4cDsbBBOFnVRwpKhG/HNfOUw/Dovd8CoctS1
WOX8m+MWCLYqfc7zw2ai3hb5Z2Q/AzT9HcEZC+JZY6vxWfcrjRgTMNO2A16gpUfR
3VoqNUsesfIGVkJsGuxw3ttDF0SrD0twm4IFa5Pig8fWyIz81vRY4AzvByP+uPvp
WLYqSEJ0v1RHsN23mtdyKmwSdowUjWfNlarAlw4oBq31zfuZxw9cvrLiXiY+CpLx
OG9yB5tZ0DRQXbBin5mIZfFMMpUylOaZlR79G+w3O7yesqZuQs6+5lRtU5/PhwCi
woaFjmZAxUeDkif1TCvpNJlNnsLBkAzLz3iZFwdQ3SL9U4H9ZQCBOGnlWFUF9KC6
jawTJvQIJ3yfUFMSp7hGvMK5dD5lDrY72a7dYS7bJtjZLjmlIZlbj1kA/DplZK6T
UcCJS9i4ehM/TubQW7fBYHvq+MmncVMxDX9IVlNIWAOnLClvg9r+oLJwrjaHc6Ja
fcZ5NLudHFjABg101JUV7yEziuNgeYf14oJoIywGKLlNEevJSPF7g4FWYKE12i6O
mZ8YaPA2yR/uUuKx6DZkRbMwwFTjMouhmkDF7Pih0GQ6+GfqpLBdub1Jx3dGhRVK
K5VYQJqHROcMeRwtUygp7huBNntQONFs1t755VrAyWnz/BfsT22FbZ3PvsbwLdFe
kgXJsbnKsZyBL82eZNm9ENAXe++iFZ5krzQEDBSOzlllAoMl+509Yr7/LPZlQLW8
GUENLVGaqZYF7EZUeh+rOBLWQZjoe3N6IBJXqMFeWJvEZEr5hZ0Hcybb6+BT8Vsp
CooeFQ+CxRCv5XLJx/FWHowYR9oeWBrUGYGu3vbQC8cPXwoCcBeGjA0cecB4QnKa
YMuH3LL4JaRa9geyoW4/y1Id6h9ITpzAtGIZIwMXWRfF51iLMhp7jD6tm53LfAue
z3UnUtX/gxBjwSGHau+8XJmgYT/AIXqH0sIyOQpljTO9hcnfXIN3Vr8mi3P4fGOo
SvK5UZKfQng9Yo2EL9le8NF7n7xz6iWcOsZTAnwGH21d2QFDDkCJl0JysLrpA/BA
j4YPJu+ce4FnBDB3CQ11GlJ+Jk1+Gzap/jafblAw98Zn3XlqJMP61QvfEzHRBKBq
UgwW1dzREjmUQyzXQmvmjWrpzqG8qznTKAAuLHUh8habRT4f+MJrtTtWxmt2rWBW
AT8NhgxjUNDikBOuqK9zTzdzFqCkR2lpnq+BmuZWX6YJDYOhpNUP/6v0URUquDvy
NofhrwlXeqqfSaYjQ2v/EpkmPxAyED9JGs2PWM/rmjeUIJVayDvoYKU5SZqmo+P/
wDCZ5LwqF6ZtpWHBSRkpqkx7CLyvFsIPbScgCYcolIOTEBNIST05nxZ+00km0Y0a
4d/RDnL/C06MXZ2d3VQyezDRQUOhQYlwJ/fwKS1+Kazasqi/7r1tLsmTxEaFC5Nb
4efQtb8iKhM42kFc3s7Ilit6cESPmodeYUd5W89gj4wQxUjLO14KDe3e/Q9cWJQ0
7/7mQ24hUnkewCB9U6RuaymL2FlKG/DrI39duHkri3YJUcKQeyvWilW36hBUJV0u
VBhXwXliJ+ltoVH3f8sIje4/SXsG5TLqv78L00ibtaAV45krW13vixHJqIUW67tn
ASv9sqBEU/sVjzTDvzri/TjsHAXTkq5gQ5cxvAi8L0WFOdQDwdpQk4Xgrsr7svct
K4XjuxUrYc3f0eQMoulCOxt6mR4aGKIyBk9smvQqUopycccc0GUqnljMgztQR4lm
aHZYbQapMvR3WNjAzknd5MlKSLO8JJRa/k+uyAvUTt8Ty0FDWaSOzj1lYmXjAjGm
IjGAZKXabOOlWAjn8JHqJP9uu/LfrRgwARF4ukhOphXOByMbpquOKHMaTaM6PgU3
tFxDo6ASslUtTGsglL7wKblDTWOTOBmRL0oVDOKedvK8wXvDRpd+I+qhvsrhPR/W
F0bpoB5agwPxyVb3sXxc0TqkZXHZlo+NWsxd8Bzj2grmEEgrz8zt2Ou+y0PtFM6z
HCehAYlMla0ZT0lk7FOUnv0csJotX9X5167Ek9F7g83daA/dzn7DGENjJQb5ixRj
m/Fe8jWytSzR4mfHxKAavKJFOP98lXDqdNxgyqpzEGWD4ZG9j52r6x8czVrvwXxC
uB1R73GzjLBqFSlfDsdTw9X424o6+FzAZV9CWZ7O9CJhmneNlW1Hxuq6cKeXxnNv
rwJ32NZYqv8xlymm4WQ437wu01Q3FQhL0qINPO1xHUd/vXgdolGx89kbEZBc0OUw
gwY+h9mLITySkiUu7EAJV15ZwC0puFap/MkDmy4m0AUnQtetH5iO8mYYA6F70Jyf
3ZVSkxawnJZctzDeh9Otrbl7Jrlq4vY4Pzut0wfg7SHm79z8LPvlEBP18TY4oSLd
JacAnEYxThfhy8NOd7wORMwr2CR9sV88Q+9lEOF5etgYg+aR9Y1E6v1N+/6+627W
wUH7ICDZGjkOzNMsz61hk0x15u939AjS/XCxtQ8K6m/0Ga65GjZsazcJuNJvy9Az
bmmX+rM7pv6wIJ/t1tFlwQabILNd51g0dwYvRzqmgOnAKXMkvUu7oCgKPRlJemXz
bF7sxJh7NqIKMz9FRe3tEXBwC0Uo5QPZbvtRkmwh5yXfb7s/fk1C1aRkxD9qvM0Z
OtDMis7mzlyd4yWEm1psWXDkqdDCofSCSwyAxGxjLsQIqfaywGvbR83gSBt62pk5
xuuoPoucDLta+M0voxhvA3yYFhxHPUq1eMpuaBFM3GUqPgbgkONS4E+h3fxnTn3p
eImRhsQv/8L1sGAPtjx4V14e/HFlDeY7tAT1Kiezt/fCN87FcJ3f29zFDhzw/8Qo
H8113vVeOmtXIyi52YCbYDj1OKmCKAUvW9Wu3zQh+xVmw9a3saewOcer91GHgvvW
0+uQzQnBJlLGdt+vNgeAN73VyVny6kkbJRYuOZnGKafZbgIhKTZyNJNsZWm6Pqha
gbY3S8apb+x7YZe+RlYLn6oE78upKKnRvHcr1wMwHOvgKgIDMvBfrE523K3OoCVT
hfkY+GQgKLy+ELhfy3DfeQBOnKdXVa1mO6gd+TlWl8uDpWzyq6isXzI45l5l7O+k
D0ors4nOuvcpD2QRy59bgZtxaFs8eSkTIo5A2YLEC22lPUmSLGNHGNDw/sCeWii6
Bl7i4Lrs4uyxqPivG2pfNz5ItXRHqE0JkIhFDk7HGvqw37BX5Gt//xAyM2d6iO3+
kHj82WxGLxI03Xc/5e3UQpaGy7BtaHm2XRgZ8qZ/1xggp1y5pvJwSCsHv2lgdjjS
ORHqeYxUeJ6Xoeb0+K7Jo8hlfdPDSp/5cSbq7rT6euBfIG23YJgzfYCS/X0iEz0V
S92NJYZ9Sr/RvbPEHDE0D2czCqWvFSwsWY3eGsdteZRhG8yIFLRoN1r3pyhzVN9V
7eVqV4Wgux6/WV7Nxw51um9HnzM3n0R5ClCwpqizFSfUsck+W81tz7kro9Bd/duU
YHYUBHO0uDxg0Xmc8XtyUBZbjvIEcLSkMU4OnMhfIMIgngC1WpEhiOu5JfROCJmw
Q9lACvJspr8bwe19TufuNo2o/JiGOAUWZA5CdLGV4perIA9SyMlNb1gXzI5J+NN7
dYbZktEC2916u5bVjWP2+OGfSL4iQaG2tEfZY5D22Qh8xsmPO72fZuD5z0/3Yyx9
wb1Cx0Qvr1GZ2sQ0F5TywsuIT3vuPw7677HbcXIJV6NDA2GOJYdugNPMNyulGEmo
wf8gPEgDC0jT6vIKSUxmHGjIektj40CmNmn8FOOK+tiHuDEp6NzML0T82MrJ03o8
Swre2h4BB00WdYT+PauqbdJQ4td8yJ2h26Rxmk56dp/1gBGM5P2muqEP0DWIp75k
Da3uFrDG5R+1fX0ZQrdiVTz8sBF/6tzJoJnjePzaegNAGV7lI3XAzeB3guUlNknt
HlkbmrPdwfzXDXDFKSzVq09HHiayQi8II7SHnK09yB3MjaMKV25+GNiAi6vqpGrb
2jPsn9pZ0FwT2Jjag31IGpFUes5ci+F49BY7+q4l1Qw7xIc3Z/mC+29VK+v9Tsan
Oc35sjVBnzaSfLVd+SHcmErPlbimJr4G+gupsO3OAs653aKWAchTIV9fFwJ7LSpo
guxONkHNBeCsuubiW5Jls7xxTCfi+SLfd6DX+SPVgJphq0XL6i35ccrX0A9IQDD4
BtTA00Sn0pWlAbQK9rIQNKO6KkmIbfRSpFn6cHUjJ+YCu5pZBTFTWQ/Ar3jTjgKB
Zvv/ccD8yegMLqpJ4ogTAafmIFhjnYvRq1QDsBf0r6ucUtWzZLXYfOYNU+7sOoON
zkCajgQNn9yALdZlGCCwfzVe9OWtqZ7A2JZD5DX11VYaWY7DSzkSy4FpDV4fJJG+
y3wJr0Y6Km9bFBipzx8nRM55syoYRk2pt/4D24z7SkkUBuiAYiRc23tO7G/R3Plg
+fNF91ZsK8WtXIC9ejjncaR7JOSfsRM4ZxM7SG/Vz2rej6gStuaMlnrL77rq4Lz8
zWDRCKtccUIP6r+A6OXaMqmTRGd7x4lz50Bdjkl+uXYSqEmzLJ1QWISg7FwIbB8g
BYHR1kf7LPr7y9k6njpGZArd27p3q5gWKN+DRO1UYJRShs2D2+zHUIw71sBbVyyy
4CngDltUXDTTegVjDX37ZYmS1yGa/F7tpoitZn+2mChwLILzPguCPRn2P8GaeeoW
ql8wvEWOGgsqnHWqlFlDI8/OhGayWT1efMiiAcAcWni/WOuU0izQMHgolsYnEaLn
mpiEjr5bCKGnFwSuddHcN5Z6ftyXRr9lw6LoXlU3cMXFDhb33QfT5VPnzgKDRQtR
by6qSC1Nhq6882NeFvPh8Ui/EelGR3THTkkuyGMTzukgxKOhOaOsiMJ5Ez5y7B0Y
IOG7gdnDmUR1LGqMb+OPpOLAVf70DOUs8VQDf4+jznfuP6E6sJNY0GTwnIzP0QVk
i22T2WHERebFzaWklxFXb8LHjknjL0II+WR2N57yXva5lVWlpwZRJVmajdFonPNS
IvUu60Ec6atDAQm+WgJBPjNjXZdD9CTgcTKxWX/YV/lwy6MDZHEgsrKEnNoTGIgC
QboZJR6YQrg5oKutkvJdBqcuQbV2v3onZIZGDUBE337Zi1prWlZHKhgZT6Nx4Twu
4BHR7JnUtoffFuppFr9RehqKZpJR93udNf2A9BAsX63+eJU6q6co2qSmKd4v4LCu
25Wp76ACrbNhA2zUBrhvPb1P/tqa+/kOTzuI+6JP0kKHe4BqTHyjbnTWIf2T3iEk
AfS5jKab5Nth159K/U3LLeX95k23vWyUfvwOkG1/A4O0B6LiS8qRurCW2xcOLPxE
coUAsNzjN09MR2lW8KgGBn+D5k0l0qB0ErNzcYDKvKQClD7nLXNc/wK8ZW2wP+dI
cOEFHI/mtBZkJGKu9rRDaIrgWIN1a+m5+AhA37edFZdy0q/JrEHqDHQ3LyCnK9/G
UEyqBXrBKDfgHB+NzoYhDtqkGg3NBJE/5YgxhSFKmzUeg84NAvsQ7oC5x9o+RduX
FPb3lHNyotExz0I0HCXfYszllw+UHvbH1565LRDiiGstBKSGzPzIzAjzMSHL7/fh
rAIl3sMTWj1UaiOE7EsDZl+7HB3x1U0aOQary2ZkIxfT9FkTeMtxKBvAiqsgFO+Y
VVxH9IX7ItbSOOi0fIG5Mp79C8UWm65U0Z9Gi8kcal2Momm4Xr2pp/KuJhn3/Ry5
RKbihb0W6m+sJgHJOweLhaWDxaHK7SvlRcUAmWynwpEk7nBrEhPx7z6YU9gOCX2c
ddPETfcvN6M22nN3uov0E4C2Skh9C9UtjCIrHrdfqM0K6jRjjr+Wto+1D6N6Jwev
pmv4iQaF88gAaktrPbRAQIRH6OzEnTBls7WleeKB3NM1uGXO3FjA0DSvVeF0C3se
BaHSXbWfPlWY0zmyP8fxF/NVvv9V2Ad1NKkZmTSxCo3JQKvwnZvgxQxGrvqivw0r
mw7NeAQ4Argg2y/AEkX/CmhG81xeJgYG0rB1OYQGm9gX4iwCx5PKCKipG4ULDuSN
owoQt2/wJ6em5CEMUpjwnEYTEMHp/YgHi3hB2wdToYFxBGeCKXrLwtFMae65ARmH
EKcwCoISsCSzTupaqGgQ4Vr73MS3fc4g2iO33KlLeSmi7jqwsTIE81gZ/QuQGP3R
b6u6y3Pa4xn2225FV1OK4MKwndoNkmRofyjud7ZJj2d3mBtUTFfDTfy/tbBqRP0F
6fAWozLHzEU9P6XLKzyNzQu8PPCBzlO2H16cHgDSRe6+/XYQtR92vm2O/KLS59ZT
Yj84VEDMlUbJcY3P/9j05OQFQYyvY7eRn31Dl23zZVA52hZCWt8PQkNSMs+C5vRm
Zr36i3Yx1qF6QQNarTEqu/mu7ZPdGGaG9Fug0JetB1ETHRHfVV9/5T/d1rxwyPo+
bPJpSOegmsu7JR/Lw3zUmkmwGxfzofwGv/YAg7/Ht3WUsbxx7bAgVqzsSM+t1Mw3
i2+ieORNypUmpo2rrHkAidhKoejwT38+OiMeTJkQssYxFQOY8GTeQvxASW7hOpps
/C2KXaLlJh8GEHSjRXlTZsP7sZlY/lG0tqWvjwi+D2Qh2VuhixYfI7LrqHkHWLpg
HkBNnvPOzUxFgZ08QFHi7lFuOoYCFwtPf+N9MhWsEOcc+S2D4XVVAB9Q74TGi61L
2YCKzVxxeePBlLTBFZgXvkk9ro81eVlLXcQlRf66Lg5/FHaVEoFciC3e1gbzF2Qz
s/BaD6sgC+igaLuYx1gxGg6Ynftx+5qyvhDunIsIHwTtVllMwjk3tWlOwbfzfQpB
OmWfTKdP1pRRk55kbGOzwIpeP5RlYyhybGuJ/ptn9rAMVkCruSzRMBIgMr5FvcHh
egV4maKaB61AQkhSSEbr7XRKy2ErYC0gwS0PThmLGVuP9Dragfyl07r6MNQH3XtV
DVvNFfEGyFAHEoe6p6QjRFPwvtjGBBQrQWUrHlft8ywipPPR7MQ7JUPR2wB9JHY2
zHLS0J20E+9MladKK/JlP9RWA9IysB7HAw13ieDjtk1nkrcL3D13bh5X7wSmxSC3
bEn58zKZQLMzoAH6ewUeAjb6LXDOlt717eB2wy6YDd3PvF6EOv04UdyXzkDzulPr
pXM8EADFPOhbdmUJnxudzUd7+OuoFUUdajcFx4ZDJV3IX0aBOuNVS2dhsrnn5cfz
3RfTNIQChu27to97JAZ3Zs2d4kbyiHw0d/8L6HkllA9y6BinRqdll57DF2fyFxmA
arRzGuR3PX6AIq7/CjZU8LxpbFz8uJ5zhVphWz5Jsip9amD4h+4bHgvOQhjDZlAs
/R0maS3KPKT8G3VPh2bjtXplM3V22YQk9XYKGhURu0kgwLu46FVKJomltwMWhIIB
80hHHkgZM+2YouvGMRPYuisJ310WFO47O/o9k9NRpZhCI+qcFq5QUPA6P2KKsFEs
FxyzbDa4MrxKWwV2w6ffW63FvseY5fOswyLvaojj9Rwip1sNoS+6xBi/0Pspaflk
ee0CzF7XYNhhTK4tg/qP2smqbJj4+8TfDINnx7M+RHzUmKDc08CrQ5dQqcwlh5RC
aaOyd6kg98ebqgsxIGBO8O1Jp79Qq2EdO3iik6RQanL8XTQooP6n4q03iEUvrnEz
hP0ZVL5pewaRAn6Cxj6atCk61TKDhnivEdfAfEFSrjQfmvusiuDYa2H+461xow/g
Rs7vAbAjkESgVcbI9iHFv7RThp8jMNSNM8GQ03/nsR6A4rBUPQNT/up9VHBxtrxv
dpWHcIP3Ab833eCquf8ok3039EoF8JtQ3YXr7RgHWIwszswqfKWHsROSIGaFVZEj
4HtGmUcOn59Pc1KoNz442itJxdTH96aiiUGA7aJAN6RkugnDIkpH+eOpegSmaPjr
QnjLhGIQ+v4OilYts3WH9lYN94nn14B1gqWmbs/Yqy6ZESq4YAXF7ax9yS8/r1j/
koNVKwxyHk4HT0qbaLQp6M8GgZjct8iem6XNR+e6lXQ5b+m/JcnupneLCUAue6PF
/16B0itjn58keHARYCk4hCGIz4T/a7cv/x5sz0/9o/t/ERDXo28K7Hwmf1R26ALF
v+LSr3qRl2UAOpnabrrZEtcdaCzPoCTQn+tKGPLu8KpGvHy/HW4HRtX+BnAsiVTF
k1TGBqSy+a8CP4ZZZCBqN2GmE+oWvX4XUmsX8EydHhqKsWTUx+NxpwoooDcoEZhO
+83OrvHa9e0AyGhltiOZZm1gDHFdZp71/92K4iHxtlNGOUr5BTjCWuDkKqISNF9Y
V0VhRAhnsIU3MfJ+bXk0NnWYbtLlIvMSP2CtJ3EXRmrONRKpU/x4Pa5IRnliJhn9
YmiPAyze+0r5wL1S8gmALlypQi3xsPUnwMh//RUlOl1808vuux/NuIIOHZkX77YE
O6fAaCnNJun+0anyb2mm5fUi3MFRLd2PM8Vp+fylDRsyvEtQ/ovQ5Ts/kd8V7/pG
Y/9BOBoXrwlSDtiLWPSFLK8WYQfhayOsR/Lhu8rRwiUsekV/K+VxPCglwLqBrYDy
XJTNmmumAiDLdMumGaVIjkjAuQeNKn10ggeIkSptlhWCQQQpDXlKSwgn4MchrzcL
Sn7BtojR2adAleNByzIVCYZcKOzeo2sZEOxURnKYcbj9yyrU3b+mlkxTR23JTvHg
uc//MiKEqGEaiW1p+g12y5lc3B2+/fQ+JdnRCRyb8FYK4f/JsEGka7XnF9E4k338
R0z3tsTWEMjXOkIHWavt9c3X6X/+pZc9yMqUQQJOktIaQ6GZoIZNnWU2o+qu3BfW
hg4yV8Y9Hs+8obSbJrkrlJ780djyOkxRrQuOP3QfrPj7CGu5Gu8Dm8D+kZB4SUK3
i+NmgYzRWLTLfFflKPLRkFzxpvNgrM8Y3oHyPi7kQBH6IlaIdcSU7iDCkBpkxELn
qe1xCM5d+eCxLsToUHJvEfSTAAEiurWgnpi3MrUOJc6I3r9fPq+QjVDJlLfcZzXo
WXRHmp0haDX7fP8Btx41RZz1i/hgo9UcZY/WjBEutxmqMXqTA3tiG3g9lDxwyhc3
18cncO+JWqRXJkkzT9CVWicxP3vboAtQt3/T9DlNYPjKcs59NQ8jF5sfXm3ozH93
8LHJ7NPkC5PmZMt2HmXepbmlFA27b2YFSFcRjJLOUKuP2UaizPgFowpCJyD3OdIg
ss/w6sjtNVFN4muUJhPuZcoFYWvaeIiYHvVfBpRQ5ilRfH5K4TvAehx+TA37ZsD2
uktOcHaPvjQPFCg5EQeIzt5DkSXXCE69NKGW1NdJxcA7sWm6biALJEbxc21Zillg
ptCAhksRQI8tlLXOFyE67dLA8yHzKtCS0IUC+grxQ0r7jl5uCG6hOvcsXPC+3kJP
rblPd1/26dMc22QuDGMDWT7XZKzi0E2JRb57iGPXYNOTbf5RfdEeBM7bbb3RbVOU
T7JeVua0k+eLPt7iAu4J49ismtuc1KG0bwO0osCmjrHe4Wxk9m3hqZn+7lQeuo2k
Kuy7/qI25N9oqSf9xn7WazCfO+KaRr0vw4idQOXuRBzKwZUcII5i9sfDL1siDZwe
zLg4gzIG50tbOHnBLbY6iF1ppA1iMPARl2xUwEonLVFU5PQcbj+G1HO1fvRHzQnf
vD+sxndtw1MbQRY3yTHoK2RxsBVP49Z7HJGa9TNcQqR0Ra1YF9Z3fFDKFb0bbgSx
28HAg80YwV6Tg1cjD06bh/vxW2Z7eHJfTwBBU7GT+IpuOXGDJcVitpR/8G0EIhmv
I9A+p2QAqkv4s8w6KIfXvYibyH2dmw3hTkzPpa4jrGTKwIzdpy366cm6WeyHnyN8
tdFOZr7wuyeOXWFw9nRF7rbw1oy3gTcpsrNwnxShmfxd7hrLvhPsiXLpnVGqydYt
XDFdFAz9mwqd5xVP/8tpkDRvSTls2Q5+01Bd4JJeo3V1jvnOQIz5VsmUoMdOQQDx
PKoIhgk7Fr5WyuXDSxZUDx1G1Ejmi192U/HrxqfB9Sgd7lg7XY6FAZzqNEpjQ+2r
rJwujOLPoKSH0mVIG5PAaL29XxCHbCQRC6OcOnFPcA8g/NXViZ0Sm7aI5CbxADtC
9/7T8UjHmClYWjaXiAao9qDBetUSTlhPQKgtQ3+29i/oECNzYnoOLVMQs2CK3D3h
PMGtJvv7i9VpIAnXCeqmCBZ1P5BlaaWZnphbbsSsnmIanFXl+AtGVlmBtxzYBGGO
7JjI/0YZ8N2hD2cP2cfMGXQAOobhQhrKkLkq7k4lT/fKVgxv8DuB8JNRM/EfT2p1
k+USxD8MnmhN1jsuqutLOMVC0YO9SEpWGls4OlGRaaMxjwEE9s8iRH1z8Wy8Gsry
jmZzCH5uf13Yo/O9jLm4tS3uTASSi/i24niWuAgUk8tVsvyrgB7P6Uo3jrroE6m1
h1f4vT4ZxDIxj7YBsAnMlb1ceEJdoClJ9uhsINwuIFfhiGZV0l7SFilDfH2uZLuc
346E841odhHVGRt0XmiVV2dZzIP+srqVPpa1bEU1UHXWslxpntZmGqiEfL1jcX/u
Etao5V9jEkueRmXN13JDzMVKW9amp+iY0Y8ymNkqdnvkjFSBecWNhzs3JlHdhCF6
0gt21tAoNvHLl9JUlku2drxuQem5AXoMChZTbFfB453G31/PqVYDO3M3jhC8I7uf
LbsmtbqSmPyVF0vdy3TggCbPPIz0gi0G5zY8D7RjfuF5wgo9Kpa2oCeHqyh80sxM
8YxsVveASS+Psbn3utEPxciRvvf0e6NQJN9EKjppZ1r1Ab1Zb97qPOE6a0hdsxci
aAVjs+FWcSe0psTjLFFtBAjt0qVCcZ+hFEDKrQAp2Pe0CNZAWOeHlNJudjv8m9yw
OuhQaJEVNh6Unfjh8vP4VgOOYMGxKs+q+wVXEBBG4Fy+GNOzSoA3DnP82vYvOS2P
EB2ut8bwl70zyfTA5FTqcMe7KhZ39aZoaKywS651HBuLmkIf3sqOIwbQKhPEGjcd
sa7KSgFAbPbYAZ4nOVlgF8rY/kYffVf1yNWmlkp7xko3w5G8B/1IpZx9DXn6P80W
VwFW+TSKzI4TfAVWC1Ib241h90Ex5WlIN73TrkceZt/X6Oy6rK2duxDvwDQtisxO
jXXEVHugE6KXmVI4Zn08kw9kQ5sWIGQOT6uczpJYSmh7jRFOWct8wCNf1BMxWKXc
C6Q600P9xjyGa+LERq7e50as1oX9FGtsR3QJ4iiuAUlIT79H8vussb9DSPYj8DOI
jFK9boP4kz94Y5qzEXEsKZSDICjBsIhoF6o2X5nZvUOFXNW4LZx2axI9vyA1ou64
3dzZ+wKPgOD4sTLUhFGpr8HAkBIMwUJeFFJeVymTsyuMqDFqRuBXb7Ig5+SNFtxO
br3lFGL6zcXdv5kOh5ZuNweDUoEN//1gzOniDw5xBsWne253+HCmeJLcbPkgTw9V
q/qKto9jD8A8AESwdQJL4um8z3X4KAqsG/Ejm/SFKwgJCh+SkR+m0nw/pHT8B7mm
Grm+j4BzDBtKYxJnTVyzh2GbqLB1bCzXhVWz38tVIubJtKtJ3a+BQgv7hwgT3oBH
HXc9VLY1Z1ygEgalPMlESipO3eTwx3ejpz/1VJNZR5WDbKceZDgH2UhzeplLws2r
3M9/iaywRcHWxyBY/M1/cHjUiipK8+pZ3qWxT7Ibz4nMXuRXCfqpqRaMe9FAbDZM
xsrSXEV3h1u8AuCt3a1Z0ezuBpFbG5Kt7UqyAwwL1r5S5r4Z0KYRLQI6FoShhDgE
aJVpzoyAdqSelCbRNgJf0NQpnLSNWM5729oV7dPMZOCzqRfJ8CGL4s20Q/wyEvIU
Mam36RLub+VUotJXNCS5/dX7tvvxVZtP2UULZBfvxZxShfuKdlyaTygqkQF5mvXY
bByxAw0BNhVojFiwjv7YAxvUhUbhCIQHapyrg3lr2GsYi3SEzuUecilo+usVHrlu
4JZXfkQtpp0HWM2Mbr/5L8JaP7r+Y7Faei18909UiKtwRw0W4sAxz1krPji/OXW9
ud2VCmjhjChH3xZko7t65YbEWVsH4238jfyjANCrEzmI8CQce9NVd86HMLCbU+tG
WIMykTtJklpXT5hs//XR83SW8Fqi8K3lwgbvpIbvCJxBtuBnfO4Bou1NEKUIaz8B
1QCtsq2Xwi//2vfHaXWVxVx/b5KwocBmxMZbNnn3JN01+kfUuFDih5OBZtSGkkCR
y+cwHTr0p/4q8qWGdMHOnTovxdZAU0wrf5t+wEysG+FobqnBGikidNezsGZdubPT
jf18pC67KQmR7J8F/QvK/8XiT8HTKm40VAZe7bbuPI3QhtETmVBBo6Z9/CjiB7IO
4+V3b3RXTWFKWogsymCAFwGnI+zuOFvTBYhMNCLROGCTaR9mXM5ansA/aS5Jm63l
G4UJ/t78tLc7OPllyXosBAcYrD/cKxwHTye4GF8hCOQv63KFD4goAlGEhnUIJe5O
ir+1d8UA2fy4Ax/tdjOjHWLIoHzfue8jM4ko7Lyf5/gseqPkfJV4qJ2VeOiFJ4YO
DLj2eob5y6MU/aNTEsj0uG658ZLTHXd5vKegAt+K0ve/cGPy9/519sC8vXgbsvRx
A+a+HbJQwEM/El+XLX+J26g3yuNZsb+0FXZl2IJ5wctTceJmUrL1IeTnVM3r5nRs
qL9wIHrhvTrBtXDOJXYHdBCdtAo3PTluduDVE7Bh6ihTBk9MWSGJP+c86QuU+LcH
GRQNsJz5jeuzbtP9w3QuxYES7nk3DLj2Oa5pWPB+goClLTYiMUYcBSebn58yvYu2
yBzJzvnAl0c/jmouQgGidgaAN9vf8ciox07vUEWwIm6A62BK9OjmofZNQBrvHrmT
kWFpBBTQEk07Bg+Ihz2c7SQLGswFP3A2VlnGcAW0Ek0i0hv8YFFfW8kVd8WdQksL
8yBi1cxwxAJ8QPOayVwGIrVMR7RxX5Tln9j+1xRZkupS/grl1ovOMevXHDFQMtmB
1fsZ8PTQomLCmhmCsCU4papjaU60+qyQRPWo16Df9WjW2DSotl5RQ1YQLjUhWSTh
GrKtRPHYdHzyb5KPursU2zKzpPKEiHYdrgJDx2ZvntQijIIryREDkKi0uZ66E9tx
ULpy4ED2MIS4EPTRP1OkeVus4XCZAA9B8LEJNQ0lgrMvkVBiv1/WZkDXNdQor2jT
zar7+5JaBTs9UvrA7HI2PVksJhJDTey9e7r0jREAKh/frE6zIFFtbhX9XPzypJ66
9lj4vtkBUxrf70svjRtBjTCB/rsOhsTB6/mQ4TROf+9wZ2NtGMnqT5h4X3NR/F9N
qdZGo9AjEcZB8/9tMNtApd6PNnjM84Wj5tPIbxmRiMmdgDMXhKUABB/KQqnpCPwD
9gCXZ3Ramaidjr72F4JfX/Uhfr2B/UhCp0Z2RkkvrmhiUJRYp5W7Cth/S4mOi1eF
geMc8G1Ypeoq+UsJ243pnuWaA/SJFX1ft1tcW43nlNvFb7C4MNkaDcedPQllulKq
aM+JfqJdrxnRlQJLLl6cx0lJL6SkZbHGBUIOy1V6fn8XzraROGK3ETilZnNZ372m
NGGQDYP7u8YJP9Jrl5nmXkmjcgxi7JNNMizdw8DAIlM/9u0XgbPd3LMNyy41XrH8
q3N2sEVM2S/I2W29FJGqCP/Ul3KBois7VELvKhKGuYhLkjTDAGHIgqipvtWmsXPV
T4YF9vINKOKInKmHHHeq+E0YhuuTL4n1YBT98siZd5f2vqZHv3HYvtQ/5I4zN8Dv
L1ceyGrn+Zb+qfDqNTurOgTpZV862CErY2M+gGMZFOGJAlyzcHBF6ikcPWUtztG7
f8NLYOqgALXp7Eb7bDDzelC4hfXUc+YMltvnu7hbgWCPNZyhen5Z8pfMPNDQ29Sm
om84xu0NzileuuzyXrK44iN2w1m+cF9Cnuozh7RgTz22GmgvpfBNhgNeBWOPoCzf
flp4gWTYxEhI6G3Imwc6+va5JhYAN3OQHlQvwKKriMv90vOi5lWIoeB8VmB109H/
EB9Ikm2uZAjQ8nt5Veq+ncaW/fKQr59a+/jjErAiM77Z811CHBsUCE4KCAl9FVPX
uV0103CrjHaFBcHe9+DZz2vFDrOdZ4AQ6MUZ6ALE4aJiaf9qCTn8LGG4qES48muT
hOh9+vWuTjPmSNP8Dlbh3KTgi48W5dHQhcNiGgtMToSM0hbncTOS7ybfcoXNzimo
OKzqdaNvs6mY6/DbeeIi6XWAhqPxmxLj75vxEaHT9JqjR6X+PYIUdtMl2Pi1G+Hq
4/pRbuxwZ4iwOKw/0GgyjBoEyUiUq4Qo2Bjiw3ul7/Bjo1nXf2VvuPOrBd5dOewv
nEH0Wtbu1VaPBzGK5eF0MRUB+ZOF8juBHIZ9vIAu/Zv0kzNCbgYh7B0vaHcDFb6x
vo7QLNmfsdHTtFKYM1gEsYnfyyFAIgOMsGXhxVswMPVTZf04Whwd1NPBXOloQwPu
5yd7JUJ8bHi8hYf17SrzmGDer2zbLpmXv0k/Sjx5AalekBSJ9gNepmwpu/YgIAZ0
aAhC6vbZCqsWleSxDqtyKhxTA7vEthbqL+lKH6/RnnpbpXP6T4tRibSTwM6CArTS
HXzhuYTr3QMqugdnFla1QRCQsiPE08MMKlo/V5S1GiX+hJJoWTUUmEu2nLL/VJHe
RS9aEgzsyao/1+RNUEpZdjyqk9aBNeAus6/NdVPK7hUKVDW2azUY9UeFnQqw47t5
wL1vF7BfVy1ia9ELfkINXlM4+X5nnyzwk7k470oOE/t0p/yXJIk37ufEyTgmmTdO
mbSk3qSeBY0/VTWIanxD796jCnwUBYQhqxspGepzeMK729qzRv+YRNeU7tgquaMc
1d+axjSBThUvsJ3A9J/g8hcmVvkrMw60NOGM5h3JCbY8oe5LTaGB4BSh9dNeuJI1
R69QK+eputQarNQA02TQSTWdQb4fwGqYqslQL73s3iqCKqJlbloO9XcXW6PtBQVY
54NjURyq6ddwuDAX5lSozJuENhCoD4KtZYDeQkalfKq/ms+k2k0JWezWal1Imryd
qlHiN5zC7hurZJbfGGz3aqR2rpUDdAVQNVyH/coBOiKbkXBrC0LUiNG9l96fANb/
1gsoC70euxzfjqZ0FV8EzPvba0ejF70z4ub2Et1J4ULqTuqGAlJ1+YVy0+vCq6/l
MMMTmcjESlGiH9qNqrfHoiG2bmgR6tVnW9XIfOCdlUGS0ByXpsos3x6Wv3omTQYl
2rvLtuEPPLAbBSH53M3yww4CsBNhy7ZExpE3B8c+7/7isf1USkKWJRhArP3SsiNG
aRpG2ZDL8U3rtwY5luu4J1ZcIh9Y8Hz+3DtUfpcEQDe/KdjOTmh4WWNXtCGl5idB
yd8EDHLHRpye1dEMlS8DXUu7JE8+u6QvwbR3YLL86z/fpy9ZXibNNPrYaRlyP5Fk
QqcoAu0uVck7YeJ6qbGE5vIRDoKA149Arp2DdNzRa4oiYzvcK99sZYxS6Xhsn5vi
yPVgusmfJIL2vpSRnVHRbTQbJsTSRglcrj8X0z2sZw2C/sG1Qju2oAUhToz4z99n
n8lO/srEcPaYaUXsvXP2CbswGRsg+RfltA+/TVqZeDzRzdDGFBBeHmO6nqEqWXvM
Be98+uSVFqEvkufP9QvO+HiIzMc9KgWd3+oTHm/Xcg4F3dSZ3UX1C8j45AE3m/iJ
SVBH5K5wXFidG0iUdB+hKtdPyKVXuxlv1SD4Ev1HSTOiocy4ph3t89b6tUjo8Fec
uUTUONG3s6W4Ydp4diE1KlKuuh57hs/VhC8rOurweTkiEZd5I3Ikfz/6QqDhJpOl
A9e5q9YX4PjaR4sxnnw8rhmuWz5KTNgPqAa8YIjkHBqqot2Wnb5lN8Du4Qdda2fE
p6NtiE7Vq/SR/OfLy3U9pRcZacnJlfZ1bdXYkphF+SMnKjur4czX4c7bbPKRmGWo
BWkfEMZ9CzJfGgKBXErlXXKA9ebTOwa6ZoqYXSuAiRhg9rTiffU4h/5EtzMObQRH
upzrUZ6sQvY/ByJXIVIMB3KFG78MyTFRG5WeyJ/+5HRsDyTu2bmDsUHyiL+IYeaF
FMmxbrLFmXDj3cZ0tMX5Gt58fUc59rFObQm2fQsztJPBqwAhFHuStzGnGLQbSGGw
1ykreE6pNNxBFd4DAKrnhadvgb2yUuS2hyf99R1E1r8MQn3cu9c//a9E+o1mNf8m
kFQXvL/ZsdQX+apWd/P6rgV9Vf7O3USvTbbdZhyqYHM35ohw2r06rOVr8FrkBIZj
PHt6PdLNVu7jiQXs5eKgiXZJrMHeYeNbQBxQr6U8ya8LJ8suOVAJVR7nCOovWeV5
w2Aket6c+UGCvdUa8o/vMXfTWxZekzlq/8Dq76V06Xm8diRoya6LUjWtVxXcILG5
FTNAVryz5lm0gpxG1pJa19s17n6pneC2h3On2dK0/lcJRtMpdvWG4G/SCuvt1ax8
1xPdhfvkKuhzuqpATgRbKeDhnNOFndy2Hamf4+61Sgt/RLyIl4Ki/vFIkr5y6bEw
zwvf8pdzvxaQ/UgpGHCtBtnIOQAJLDClClMVVlNTL2wxtQtjsBNwPQhsjHM4aswO
u2LT1g2/OHmj1G5LO9fT3OHRMCx2jcYStZNJVYZU9PMnPQEJVkWjv9Ly3ANRkCRt
Jk5g8aGisWJOUVLrQyqvI+NdxbhbJfecDocuswHzFe4ghuQgHQ4/qzfGrBa+tBu8
1DUME5jWKF/DBfKM6ZMW+Fc5DFXa3g3SM4ljtBptsi/QseaxXiwSZIyAKBrkTdKh
XQhDGjO8+qiXP89GX8zN6kt/4bPvIKHo7yUD94DtFG43NVlTyH5z6stoB8WOqq+F
4wC/TjPXJo7cmI7ZT6NvK8m90C3VPZ+Qdf07Di5E3o99W9D2UgkfPddzx8DqA8fL
B5qlVQyzk224dDo2Q5gLC5sUJVHdbHGXF393pIG4QcLQp//TOVNO/5jG4Vreyo0Q
SziUOvlk3pe+azwY5VYP544EVy6MDAI8JtaJ6bjZk7TfMW5ZFWxm4oDW6IgzmGXv
u9Rqyl3wWulkCdwY8mitMCQNEBHFvPIUSUNTZAPh2vExonWXHrgQlmAP9rc/ZDbW
GCJGxrnC6AIwjSKe6QT4V/ZpPnPmZ8yqlewPolIjIfGC9pGOAMyzOhNDXWuyP3LT
WkYKzKHrx93dXRGmhEExx0WAG4fh7olTeihj2ARhJp6aISq5YNIQPdgwlImXHPS6
zUoAe20nu6G6leQQnohlayidfRfAaenfBDfAusAuJrFt6tu4S8Xr3fkPA8wJVuFs
+mjxjh6ubos3xqVaha7VcGM9FzZzyKgR0hxkaEWxFJ8S0UWyPd0w7wHhQIxdAaBT
cnW6VCyzhGqhfZ7V5rDHCCcWsHktmHX8zx9oXUFjGVSOTjMKOTTDAciYR115MMTW
VlwV0U8Ag7HfRSmpsoG179D/Z0srFoghOfmpunG9t1MNFLjGtyqvx0A8BKXb/7uT
Tp9/IKbBUei2hlZLIo7ynlBKEOFpmFLTL+RpjdYczPDmHu3mBHjfACpUFl8o7QGX
MuWpsavDn+So0Zc6GRZY6eck0p13a4BM5ONRtyDmE8yx+hQSdiMV0MQauQOUX1F5
WvHsHcfp7XzMN1XjdZ9t3MD5rZ5ThOWiZpaohR6XkyNA9dKXKb72Bk/yPsgpS99Y
P3L8M5PKucyj1A09DgYT42Uydti794tKwaYd8Ac9++fq9BY9Dt6LPfBYAwC0gWYE
q8Ld7t0MuDi3I0mF7i9KFtdnwd7nc6p7hUclYyYeD78vgRNBUgI5jcb1wjd84bK8
izJI05SxXXvDYUOWGsUroCMV5YuE73GSNFuhP/1GbATUCA8hOjHe05kx9qdt568Y
tJAL2XtPgpDsmzVfXwjon5r0ePc9f7zbmnBR+6rIsM2QTyuOa0k2YGopBDNO4kY5
Y9aNvlSJ57rKH5hzmpyAYrYJxKYeSCBdx6e4Pm29Cvrkv228SxaU2a8CjeZ4DHez
3Pyd4QxW17gka7bTnyewtRBanGvkWeBIh1/bYsDMmup65YsT4Qq+1yjdanH01MSZ
eLosPNL6ZhFsH+ar5DuSto3mjzXnkoZKYcHxN7xpHsp94pTOFAooq12+7E+p+B+t
MHSQY8AIuwYdQBMv0ql+QNkOr+PkGpikNrKkaiUnSMUHYZlMYmbfghWDnCLOXjEh
fIi+wssS252igt7lgEAu3Z06FM/O1q8/6/Yaxw83ZARn2xHeC3iDOY08E1apuuJq
YCCQcMRSyTkNW3eQ4HQaxb+CeSLoVGT8fCslGUlptGthCTA48u3Qxp4Hl5kYnOJi
ZVegJiuQtulnB2jw5/u+14RzmzIC5mgntQO9PZyy3a0+1OChG9L3FyHQlzSEY519
TCzWWkoOpxX1hPAcAaDRegtT53eBBYAyZudfgE57XYDTmKIsqn92NxYEaBoU8CYN
5EemsPNjJBeMU0sjAPcUpUsllJzfJDKUbp+9NJ+9Fk5r1S07SxsASCP9qiJqWRUe
eAejvZ0URA2JpdDthvrqUmsbsaq3Vl6z06IbEcle93tdVSmupjlmM/od7inLrER8
NHO/Deb8D91tM7UfI/Tdmas01vGU6xIL3ML5KmVw4sf7IyvJlFm1Tpuocasui7Sy
5DyMfQZEgxdi8VRWxehthm/wtMxY/ARBzVJFLDw6rUDA1OoaU0euzvI8jTSQnmT9
e2ANQSUfp0HX9SlM8z4I7TCZGh8v2U+Gozgrvbd2f6J1SvePjKYJ/wXFmQYYnzIA
a7ey+988uqMo3GkxNnKqlLK/VCZNWvyZ45KB1Z8FrLW41PJAeQkyg2oeDw149Bmd
4I5fioLAFaHXo/R/SGaBaJXszo25FwcfVyIBg2icCoJe368jCZSRYF2VOWjwYimr
t79bvD77H70gIe6x5wswn4np402i1e/WU7VN0bXHPCOPOzV9Q+FKm8a9DwDBpe9V
lfPA11f7NrNIqOFXTKxS3BdTF4Sv6xkmvhX69bKxmcC5M5DAzy+29Cscm7w9+Lkm
/zUdm/12uMGhoFPoEEGtqO68ONOEqvcIpggZ0YR/YWIbLaeVLISniIGUXsuC9DBr
ZqRgJ1RFWfWpmxB5pxb3a0c0iRmdvDHytTqTlCC5mJt0wD7Jt/zZrhGLOso/4HdK
HSCYOxkcbJ+45b1gKeMyD8L2azcox11/f7pSohHxNTCLtzNxmUX2pe3f53R2qqxy
wfROd+TUVp5f3Jz1CyIMazG4PUEZMWh1pMMQcVfFgstBMTQlSjcclVT2gTIvrjYB
dmXKircP/FjFRSYfMWvz8r19OVw3PiQwBqpr8MHrdJ3kVE3bCvNJdsanTSkL0XXw
Q5v2UvoWKuoglLhdlCDHA4QeL0KYShHyWO3nnmwvnSdX/XFg3y1BgmWDmYoTDIZC
lVxaGIbrD49cvjxbhzFGiCJezgPSRTASqkv1rFBLEBObT7dRXSaslUbh3xO1z5+h
yKeseEdji6dVZ1dD/EExO+phbBtvFI5f87v1NekRp3YLK//fPHNJW0zld+VhrSgc
zFdgxK1ohTPaLCbwq6Me9WT092ZudqstGikpHhsZiEHcHESZVnMGuSte15rDdIrC
9CJ2r1/dtlBa6VXx82ZK6eQuWudwJKndGmQ1mxV09GJKh6I0GQgQLCWypFHWbhok
OLSc5w69lEvu8OU2NLhPVllMR0ub3FNNjFqt35FHG7huDYmkbdlWeeGLPZp1Dk8U
1+WLfwDv5iaDqn+AHih7Le+jRlFAEXXodz4wQ6TJo5acPGvN/0xO3V0BIC24HRNy
tuEK9UM14trwTR1zUdyyJliwHvtG49K0R/zIxP0hSsp5CG4V4aLv15/ZwguNKYMS
JEE15UcxSQLbzVEall4PQV1mbYmi3D3t7N9P3n78NijeiJk2LFqQOh7R3/KODmDM
2lqNXw+bbeSysuR/Dx9Lw7x/wGWRvZBHrJUsljzY+PA3Z3BAAo+5hm5g4EZSStyg
bSTaRIq9FI6D1Nu2kCTZjvTf+LV1wTmgnAytkf1suR1tUDqx2JZi3egQZWvxdFbo
r9Xka6kfEdqmN6xOoO59M9KfrxhNnGRO7OiWwqrbAWcZsb7Gy4+m/nyP3a8tRw6j
HY3tYjxTxTORFHJ6d027FgtJ1U4K+kU99yczutrTbXfBSuY50f+MofLw2G2+t7Qt
oNHGxpKRBATXw4PmOWNlEPD1FRYTVQJQ+gyvvE3lqs2VgJIwmG/rLWvvOTGTYID3
hacZkbEOovqSBPfuvcWayZhfsvDp8N2z12gW2WDTaNohCoAsUwgTSFoLu/iZkkoD
hH4j6UP/dEP3HhbgKBnvsVIykKNWsHB3sMyaMql3LbzdjVxPq2rJ33HIlC7sscoe
AnHQ0ppxdbzDJVIEl4VHq7fToDLOUXMgmUfAhlwCwTcQQ2Jc0nb7QrRxOrwp0Z90
P5vzepfMFhHBGLHFD5mCS5Q5YKzdcGtx2B1rFpfQnhk05cUoHtoiNRnbyzSFciCa
YMd0t764Yy3lvJ7qbmG5sPqwEquN2DHhcV3M7seL1I/AtZzRP5tbkcXMSMMR4CeY
LLHeYhktnEfFXereWybY+Ar1G/e8HOVwKT/ofsU6B7FHtY9Hca1MHPU+pMCIKueN
IczOV/NwCNXDwdo4HpKUpOAu2vi5GWzePl22BGsaJo1aDDTCJJUuvZRZ/Tds+HcZ
8iJv6293Ki3z+mySUz0JRsUgiapjy19LvR7f2r8NlbA8JyBav0XV6bxLh8tOt+eq
XzePW90wKrdY+yGMMJ0gZAbRPHMdvWJA3eiM1Iajz81b2nDLOmTuPLj/WmQVoclN
guh7ZUNebvTsqxLEMd/uji6GVqtZ2RHA6qvAjx2mKNnyOWNn+q/J2TtX3Hsqlqjl
Mfr/qh6DIFwI84jlxL2Z2tjVJF1rzX1O6dxQv/nicV3mQUJzqknmURXEXoWA4EP5
W4U5/FDH57lA8HNxSfVfga67NgnYcpGHkoLo46fLpdIx0w6H6t7BW0O0FoXBVKkb
PwTonWHvn+pes12swZzJiwd+e2td0cKon9acAHeZ1kynJHXz70sP5BWuiS3mj6Uw
hj13GQoJGUIeyskCCqzgFDwCNcEomS2DG+slyf6PO82jI0fz4NP1deGho0lTjCnJ
XxiT7sj8xxRISZnhxot7ZNYb1bPMxWYfvSIu7/9qOqS8Hs9Q036T7RVmB+Y/4ITf
YRWjnzgxjrdRtWKK73wGu3OuRhYyQbzUKCHZk1NM1ytouzHC/1fVdmK2KXxIlxW/
si8o0lGiOQOj1E1XS4CwgvKU7RpJQq4EZ/o9a0yHbKtH5APfYsoA7b4GQnFamNXg
R3g9hNeHBBxhKEpce/T2THQFBu2i+BfsslM7+Ha9YABQB7kAi0HdZ7hbs3DPlmz5
A/MODf8okJr1JxYU3OfMOZ/fUmDZ0MJpW1hvgUKYuc5WdMKVCT65Z03irSlpuSig
fUmwO/M5Ut1Tlgoee7og8s1+Y09pjJMMuWN9L8q71emuWsFjB7YGfEU6XU4xtQvZ
OjhyYUdf31UFi9ygyRqeXkEOtZM1Pb1WJP2vYjU1j8X52jywBmXeXwpAWbLP1/3i
Fu5nQnc4X2uJadHKNQDnq0K0qTIUReIhQdc88R5xWhReYnarS2gdSMD2QiSGJgXS
meFoZROBm9BJW+lQVdvKFdkc3SgEiwhn+cjbVYeDEtHoJW4l1q8qTzhui/5RNies
Zrp70OErqLZr4dd1UStDeRRQ1PHSNTYk6Ygxj5oKRLhnDJGeerT4awx7jg0RnOqZ
ofahbReiX0f4DusifsrKO0VqhkaKRHXoryg11e+x8gRvn7/C3nV9D50pg4hPs7WS
0q3wCfED+rM74ODU1xRi2AHAUq2r8KiwYpSQlOD7gp4auCiuk6nENz24wzhpv6Zw
ghWVOTxTchYhCxPjBsE8JBy95fDnNSAY4RrtVwVQ0l5IHeAQER4SRlIYIi6gAZll
7hK5ljSZzhBVmHjEUwdCC3nn48fBDsGtwKo5vxiq4bsIm/8I+WwER+nutUbI0Nkx
SJncdnHTNLWD5ySlE81E7N1F5XrolQKRu5O2BY+KmISbqV+SnWDq24pRCV/Sca4K
4KZq0w7tpEAFqpuI1fhhVX94QXkNoOT2BKJMm8IYbS1ouX064FiL/9MmB/a3nm9F
cI7kaG2XXGXNXMqZ+g7KQIcLtoAYi/A7QLPzGUqToExUHxdED2NipsF4GfAn81k2
HlzrlLLvR6ecnYitN2RBiuARJogXLZ/Hzj9M4UgWPhEgJfvvXs4oqmB55kh1WMTM
47owwy/5rBdyFUzBRiKaEqcvCdjA0IuXi8T5y6gyJNwqbjDRkReVA7+5XNVGLdbj
DoV6H1R/XM9NjwP4eSuCcPtVr6prRuBW8iS/mk0lAf9mlBsRXSAk5I122RlcNM1U
FSy36YeoHMeor0e+r7TplSYZ7ovtnkEagZMET4AdS5xccNfJeAXDF3Kvkzv34mRz
iF4AOFhpEkQSJki+0J4KwTbjSkG3uMMJWK7vDWf4rg5zaM2WjTMYpEJ+CgQLt7IW
YuMdMOyOxgrYs8EA2oLzgQdisZNiNN8Y8OGZICcgSvsF98cPAWgj+XVxHN2kPeqO
APCmTtin6rQq/9XlzipnHcYGHqwM3HIhlz158hhSZTeG9mUFpL7hZuGdGBSv7ABx
PxSfOcGitQTQho6cOuZs0j9lqQz6qYMLtAWdvAUNPIereKETSvoRHkq77DmPtXR0
EL5FXLgvGcgjkT146KBN/s/Q8V32yRwM0+QoTjmWKbVO0+KwPZRKP1ymZBxy/cic
HQY3H2bep69rO9dBr2bXYiNRpO5A+YcotGDBHAuD0rbvgKbXAgtBcD2B5QMoJoq/
fKm8hojMahyyO9ch3lh1+S4kQg+Za9anPjGrkDdcdL/u6/YQEc55aPJgYiCBPQAK
pCqXiEFNLYMuNLzbYOTa5lqGfwe8ym7bqsL9Rh1d14CBQSPoTHPy9gsU/lmEytvO
BW9Vkaa51DExx5lMgAzy8uSG5dObVEeDxX3d8MN1BJpQSA8tbrf92ygPG75N9XsG
UhRF8vpB0TpFAu4hcKCF3eK1IADZ0UAo1pQeBJdAiViTlu0OFXH/iQFYh0covNuA
x+E6ihNXbS+Knnvq3MVbzf38EE4IuhG70LBlDSaewiL9w6HZxGOuulAP05+aShwH
WPvQsMDXyMgcFs0DiUUJQO2b35l9lxY1fpzw6PdJr6DzO3YhV0V5TD2Nj9RwgYBj
HoGzLEoiBqq1LisXclCyHEM24APzoQgRIjxyW7Ru8vWPIIVpd71y/3xo1+EJAITG
WS1aQRBqGC4qgZ16F9FgW92Yr41MxgrPcejjIsIA+dNJdLOkN4QgsqiCPPbo6h7v
oRirAkBmGJZb8+jimx35BdV9vIe23t1qYIUA3CITobZ+SHgVDjeJBtK77qvCCs7v
bTiAmnJceVhlHrZytHakh9h/zRYqWp76uwknW7Iyx5w1L7FLbztuBOEnUtRoGoS/
XDUd2BEMC0J76G9f5vOZPgitHpOUd1dSBiBKsnm8z/nLprjpkpXJRQqjckuaMBT0
HAw2HSmD2yULuzObJ1pgUziXuZB5xCizeJqOsbeEOTVWA90wkJ7lvCROssOKVXca
ThW2CdoFqr453wpgW36WvHFkllC0azxOuDOkO3vnzcPYWdYEs/aadmfMpP0pDsSa
RA+M6OeWqE4VVFybf27owzYPdriehbcgO1Ed6+o2XWjI3mTmZVgWJ8PYK7UoSGga
XrCnv1DMES65J3tDWx8dJLkp4KfkdPkPTiwl5YwVlI+c/XaTk+54hxvxhayulBXw
YHBOPRZtY0y8iw/24PxcPlG/ZFjSfq2FB4wc/ugfNclO9jpy5dLSZLxWeVGTfQpT
jFFGaANtiTHNeWDu83FReKGHQ4iMNC+7qlpXQnCIA/1ejG5eAxH8I75u0NwetveE
EUqeZ6Oo/h7/njEaCaGUfwha9YpEo/v1tPpG6fD9elEqWVHley/O5dq0h6MrqhHu
Lr4+PVKgWRoA6pz0Pz/K4izwlVA0uezNArDsSAufvSU8eidT0m5NcU4QA1EsEVIm
DVt8/7sykalDK6+w/An6mUjRGY2XuT9dPcU/2ZbT4aa5bYAQwPXizTxCtG8vcId+
UpvSduL/kRChK+zaQ1VqLcgKPnxWz8bCJBNWcatbMQT3az6pdSwZXiKEDkj+d0r3
EYZVOOl0cL8ABKtNugE3WaO0cnHEnCjOBTXWjI9eAjHcQBd/yTj6w4tOeeX3tgYP
ijKLeGM8YmAQ1BHz/a5x/mml+WTNHSoz1yX1o8LzTSW3bfvM8LBPfVyafN1xEePs
F+ggbLnXMNmrUSlT7skiKWCt0qkJM4QJLdmWKa9i1/ss9AOJcBUVduLmUpBykHox
VfnaRn2WyoSILwneqTH/7aiySpUgI7lBdgmiRSWq4OQeVkj37t3jqqGFhk3/9Q/W
oZdk0lufjTcBshuBK6imieyWYoNc8aJ0CkWPFivZ9hbqeB2YDdxdiLMJRDl7y9R3
KCA2bwMLhYGizZZbksL9zNWuwgdUykTc1DCeLGgCwxTZwCNF5qpXAYlmfe28CETX
b3r7jSJ49sEUo1fZdw4902WYsIC/er/CEtd8UwAuz94RDSPdpF3/jsba3C265Yyd
2G0eOdw2HA9dtY7wmSVwBseZ0wHZWS4q+z9HeIhJOlpzlkWM5i8XINEdr7jVyEMP
KayKkyR/e4HLpm7P53egsolS32O2R49d9WCOTdo4rT1mNJQNRtZrmNIGes288lXH
Aw/nHjKqZAym7uaFt3uLhfTfBLrsjRvHTubh+0kvdYsphUwlawrNB0J001C8eHTY
M8WbR/fgPU0XUrRF1n2bPsk5oqlqtJOcndOQrJvqiuz+42gTiObRtP33CkCHJVnN
o1g5Q5+9Ft1XrOkOCbikQbRNO/0EglaRq+EBT8Lg7lTV0pBLVEzvKcf5WVLvbR/u
VN7XbH+i3dR2yMaarMo9gM84HxiiLRRg4kO6jf3TCqk5SOATV05gQq2s9G+YKq5D
UbDHVOf3tKZISpr4NMC+FG/wXsORjB+6YzQxDasP+EZWXLKv+wuUDqO224R5xEIN
rJhIwf1gbOlduTYPWjH9rsl6gHVZEXTSvxC20jykdJ7QpmBZTDKNZkXZjbaBGRuL
IQ4Q5fB50EKfjHCaAuTuoZ3wbggvGJ3MD7XNEV9xQsEIbX4uTvAG9UQw47/ibTdh
ZVs0t1kf2d0FsKgGIA1Dh1mxYTK/qTWWb0ZjenoXnLsy4Zfvc2rO/8aexhe/6k/J
WSbrP5XnM8yzIQOVzDRei2qSQN5VCrYPdlyQyJRzC7GUyorjSdK401hhOAISy/jg
1UQhNsiHuUtR4sGOFhv7Q0LkIFq7NR5kRqa6eyFg4rsT3NlsH3gbTlEvTPMRvlXb
+E0Z7KLZGQ0mXdm7VzEXWjSMRf2pov8uu6VAb+c4NGFLNM0LfYwlD0uDCKq+Fca8
H5y/Jq0ThRn92o1GZLQjLP0w0TimJzqGqTeFRSSXGP/dUVfWjCC+V8x+a2YeseBj
f1dg1fn9OVTFOz+9RnyWkVcGPdDDM9HrUWkQXrhmPHq0PvtQ0/DBcAH6h2CnvARE
nyypSjfoLDXA7wLlXsQ/G/2qh2Ovcm8B+jU62BTe1g5m3G+xOpY78v00zYFNind5
H/NaKPcHsDKJKycPanTCIUYQb+vy2xf0kdH1uFC5h/g7d3c2+FuDKQS9cjiomKp0
yEp0m6g83H7bfji1TnYj5kzVC++iD342LEJOT+ZpuonFP3tUh6BkbyqrXinJmRFs
CJR0rPxyonFigbvjwxAqz2kicIXFvsBBK4lwXCGkFvz3+OAaXElCoqF4tPcYupOA
z/jGsGVunNyFsuSh/YSEgsw07EsXsE93/NriaMOnrpGyVhIi6I0dDUtBHdhh9vvU
SoxtLGf1397IL52RGZ4XbaQAwcx7WoO42LKZ9NDHL7XzbRJaPL0CVejr8kwS0qvy
8faN/orLojO+8uf1bSxIm1MJYZMnmbmPIGQTKXw1wFCusSDRynTrUM62dcIXlLTx
DSa3xWOlMUeLD0Yk6ZNu0a/N28yP4cWTehg3CIMKRVJxRQmbAt/odWvDHMTiEzpQ
Mexr8165UogSGfd3Be6WGxTSmEvfIIqHI9S+/pVW70Q8GxR7xaJ81PCfPQEN+HzU
YrnPwqQJdY+b93CvIOjHTX153i+veNw2z9FD/KLBtE6msMrrNBA6L0QKkSMs43ea
Ppa0RGlXO/rhUi6i+LKf+pOjUW5k4ZTvYN9sVBMKatW1h8EcKsqYAzVTW57zs496
reLZBFwsq/IxWhJgkKE+FTopst8DcoJUwX3cRouj/R+W0il74qxZH4N07nZEnARY
WzQ88V9Wzf2sH9vaTQTmGhO+qyzYj470nW0YR3/codoe2e0HqzL6Bl9GK02Izopy
9s3fs6CoVJbZFMlTa2etdBb2IxHxNi85v0uRPVWzVeSnr1G9ILYlPbaf83njM7cW
SV3sxFNsUo3Z4D40QrGLKgeBQijacCZ6yzQGqCKr6d6qdfHYhmH1ZxPzJpVkh7fb
bBGy53kb+EeY/voOgIEmU59SzzHjMLVdkoHvaaN1qb/Itdr0ZNJYcwSc4v3UA6pa
da+BTqqkBPB/cPkEaFgYfVIKKx0+E+VEqFfzRGAi/5L18h+wb/4Q5Yw9BtkDd7Pj
cSXpwRHSelUCdHTjIp8iL0Y5v6Xhep87qva1niPlCwRjuPGdy93rGs6QOTZMkLYv
2MHgzTbp8sPhqe7Fy8aGvQh1xhdk+dO0qZV+8Kv4EAeyplSnmGrfzpDnsZXlWZrf
quGYkDByvMKO3aaoGLlG46CUYmEFqvUeecu3fViiYyj2z0zx5lRCx+dM0efUKyU1
IarWBVr3+haJTOxUVu2g04LbOFoY7QsAIl81DFutaeKwdVr94hjGqDA64i2Jue+M
chigEhB7WvDQ4uKG46LtknLJfpr2gRzTuVPGllGaFc32doYMKabxdw6q4KRUwNJp
oRDkry6zpDpDrnMTIdRcaaywnUm7a4tNgy6IPwIrLhDUeICDOEhKVyA1P2m3rItz
6h7MP6jwx14QQZxjajpAdc7hZ5Y62jYAh0OXfHiwWOfAdT4GzMH8C5JDzydGR+8Z
jBqx7YH7kX8kHDgniX8uyenKAcg9GEq9jbGA47s8IT6uoNJGyA6Ue3I80gR/B1gF
/qei4wbTEi5yNVIOWrBlykD69L3XqwuFZwUWsUFPLEObqdOXvkFQO3lqz4CHSWyg
8COWWFWqdHBnLZGTlSPrzVx+gdoyRk5VaI18hSpLdRWXdAoKSqwU3zPAZWuMTpOG
75jMJqoNapEvJh+tq4Ch6+TpDXv9g2MGpX0dlbEHvQkXITlF6/SeMnvt+IAI63H8
voNdbYeSHi3fBG8YdEeYe5trSz35AlIVBg6aPzawXn+lrl59wosldPxeDBablWrf
WdwX1/fGNWewmdRYDHrwwxkG3g6PsUVLenHgbOUcb3t/0YNdiVz3361MYDOEQkER
iBgEgpdUGECWlZJ5cLUau7ThloIybbFIyyL4OKNk3JbWJZ2ufx/ACclEVWypaZMx
k0U28vuFyBRhMvcE6C4zh5mmAwXFgTsV5cU4o9z4kgHzjIpTovmpv+8SlJ3MwH2f
16odYaZ91xFbh1hDG2IbW81Qs+jwFp5BFw+kzfiShHi/+M4XTdlwENrU8RsypIZ2
2NQ3/wXzgk5R/6iP9o4GdWdW8QZBnmb6JqV1UrKFm2Tzme0o4DN+08zev0xXKBNU
hxKkdgevPFOtTEdDoLdGtkT4ONTc+KI9y2URiyXNKkPu8KIliTrcMAjorp+zjYz4
IA3sOxSVta/+mmWrHbzUh+j8OSB33kWZv26RX+KfmuLcl8quJt5L1gGVRgOWpFM0
et4M/I6+d/2tEsw6XzdDdtuT++wny+0KvEtOsqx1FLiF+1W28t3wz78PZQ/znZ0j
dEePJQmnC9mC19uS8g4PkkjwqHadZoNOYU65t+h44MmJ0jGZsWb3UrsnKwIOr2gR
5A0gRoum0M1zmv1RVE1gZrY88sBKc7kKQ+SKwTTfaIoDEH3cZVFpw0A32LEmbmap
i6ZeDr3TTcnm0LnJ+U/rpjlDy2mJFM+DwW4AIQgPuo/MF6VZDpcw6UojSCEAT9JZ
dzkaqq74oMn0GyG/cg5B3UX2N1UjOXLlLDCxagzPtcwBD4YLW1IY3R9pA2hV+Adp
CykIAUxEIPaUK9i7yhTJIQIGu0Vnx8PO797v1UxnEv2/Qt0BR6BsMn+rzFurfuat
y0NoTxMAyO9tad4nV/B78yFUb+/77RUe3fEeh1+8HFdoL2vWw8aX77s+WYUuQtaf
GH1nJz1va8SBhsvbF9F4rA+gbb123yD0hjycK04+7iQcNIFLaFVP10H22vB1FkGx
vutKrs+xwp1rcD8pdr7R0jG0Nh2hleGAUgXIePIyd65SVFx0UKkg9/Z02EsPkaSe
obWSF7TCiPmVndiSa6JvTBm+zYgEbWbfUFNyhUu9VWHCkRae1GquCbYc0OaJEjBT
mt/CRXxSl8op4uoH0/YVnbs0+tvn87heEyZ+yIr8pusJqzxqOfUM0hRjyV02EMuu
5oyXlisyDDglReICC9UhwFWgQueEN2r74dE79z6TcxwnMxl0CrBtJUcHIDQnqDKr
yzNUUarRUhGzKw7m4Ph/hx3mIfn+A156dWVpha6awiUV/saQTaEoCUS08w6W55oY
s9gVnLnbObjsRueyLdJjcGJERBd+sGwQDNDbPcpAUz3ShBOrutAE+E6JC7TkzsV+
2/0QSc1MpqPQFqW07f/QUymtxpwPQKvq4HHpiT/7WfV4NxDOiQ6KQilNvaBbqIIo
yI/mVTjxmVDAQJrxfwJ77J2kbhd0JSUbWxAf4NP02tRQPq/P+Z4XcKm/WgcbgSH3
7fUwF23/50DHZrXjnv0nLzulzOuculhxPPGu4fYLSWAgcjVQt1O+ceEatgyRP/Pa
dNK4VdTmshMnU8jWmLJbaGZDX8XAjULp6OKGmOxDWNTjlJlng79RpaxiT3p1vS/l
pthkgc1UmMO5KNGM6pg9jAO++pOihprYCKbCPYB04VOtvxfusTeUhkQNPxciDK6l
IraNZ6KTOYmSP0Jjyl7Oy+WNE5t/xrzAdPd33SHjIVK7lCkQsJHBBA7D8mxeVoGO
R42AVnDI5+gwlHmit7GoPesNWIgzfwJR2vj5Bht9sSuJHXxHWtWioBGan3DG8iXH
WQ+wUFU6kHbr7pUKL13nNkJSr9ZlfqrnVmDJ/Uzl+oJEBhQEB9BFwKJMpfb0xG6j
41Fuff7gzKx8IbarlHQS6omU0RGyv0PgSCdR/2x3Jm3+6RCUNUJI5m/jSqLRCOWW
+x1Ug4WARDFSKgEHoFBx3S59nX9eChRB9ky0tSsvxoWQRNjeHDEDM2pr8tnYRpeu
Q6ge73sJEeS6eIof+gwpAcfYKkSVPhB75IGEljgFp54My/vhMvZJs1IQgF4XD3qj
tKdEjrJI1KWxrD2tbRF/zXN06a4JWbKBxvrswHphXma2WNix15cPyUxBb6SFYxjB
OjvUTQQxsCq53gOE62KqiTgrDSPQmE9lKVBtSy9HGSM/TPtZzK2fkCSg/wAqJRQj
NLk1WG/tKx2Q3EHtcv2uhs+B6i5dbmLNmyWjZp40nyTganMK+V3n3TagjLdn8F3F
AbA4IWb+YEws7eNbSOOxaC5cWFAeE5vtqTm1C3+GcCTH8v0cEWIeELViSyIGZ3Gs
DETxlBtIsX6D1g6NTnmceBNy3lueipV1r8uFlQDuiYzvPzT8y3S/vZmCQfQ3B2Zt
levGW0Yo+rvYPyFvaWa1RNjmmmrXlz+GO9QOFUJLiSQ30c8bX7ntKykYRUDTj15d
sfajAJofM6CMUSYJSuJ/IPWB/JrMURDtYs/UtFEv483PeC/nXExdMBHcsy/rWViL
MW0GMJz3FulfyYAIStpmIUtiTAVXe4J5GoE22XiJKzXd4KVO5rDkMBwBiWX0N6j3
rM+0nSHNMV/91376CJLpy6GYU2x6/addX/exCBVdtGWEcmBWoX4yWUNuDX3hZYYL
bGISkcdJ3PkEVHnELDKpCa/zMFhuWlJrrpAKnNW0vTFRcPX4yfy4NHccqjONa9Nk
Dyn0IPY3GKwb4dkOxDd1WJ4eKOTOz/7p2VuJs5cmt9uJuth9y7EVVklDd+i4oB1s
HkG5Bu1TFxBgek+Wr2CJEE96H2EfSgwke3PfIIPr3sqgFSF3th8LDjAGVDlN9bkw
4/sJ3rQVdNylJ1v2AFkiULltoKGmPWCJFJN35F0YWwWb4rm6sEKSTjcs3NuPUAZR
JZwCe8kowVRtJK8QEsE4l2UiLBXErBChVcZju8Y+0g0NcXNW8Hbt+OgsyONh9GZl
ymxWp+HHAZfCH7wdlBfGR6L9431HF3MUUzy7DUp29L0nj6R4wSnsAKYQYLvQcHbJ
fOz0uqOLeqwtX6y7mEqZDwBQ09z9TRFLRwHB3W0cf5IO995F4AwHg+vqsty0O9+P
HC2KW8EeopNQJ5xJ1ZHB9ftiFLQfJHaJQ4lvp3HzEzlsE8PBS92B3F8mBXlFA8To
klLmqZdLRnYZHxeBBoh+BPyNfwuIONBcJIrUYaV/jP5GeM0qekC6E3+gOrmhXkaK
gPKF4nApgiNR6R2Zxna4zT9ISU3b+ewA8DSqADj9bOBAAgQK6tjvJ/vPhJmCzm4q
6uknAaYdQO/bm9RSyRVA+i6b12aF9t9VfPNx9ueuGsDyvS31xDoaqdFmEWTLWti8
2t7fV6SupaF4eWCwEjrRUc+YIshunWKotaKPlIa0tAS7OcmSKjOYgP5816Dz7mkA
zfVOZfsPu6Ri8M3mHOTpENVniZYWwxrjhK0kCvTGiroF8BWM1KILTr5WJrY89sSg
nA/iHryYbYVyVUi+1+L918oMb5dVPYUemDXy7FfmYCdIYOPBmqQa7B6Pl4r2S4ES
ad4JwTozIc+z/pJ+Vslog1cK6q8Lmyhsi7GKXA4J/pJ+PccrMFKSAjrJMmefyJG7
/BHDGaWUjYT/lLUNcsnaO/eYEe+LLLqJJW5uC+whlOypXXwS7hz4RF1v15hGHfKX
m9+h4bWnRwQcs5Z0XqUMAsZ0E5n4FhI/286DSCDzN05WhwVVsmy0UAb8bROnYnjM
s7B7ZcHnhYE4KVVR/wNnbOMUp2u2+Fa+VN6qLOa/Yerkb6o3CfJoKxQaoUlyZhhw
oMyfNc/1OZgAsS9RBrzgeww47sR7WCR2OZuIparUvZnPn7X4wL/ssZ9pJDEFHxS2
xvPxg+Qq1aRVCf6lzu5fEuOFm67cOc9YImiRrGEwJepO/zMkhW40Q0neaxjs3JCF
YFrkexyK00TMKxf6z+xLMg1KhzNULztP+LepT2ZU7TW7APJSvN1xxxX/2dgElOfc
vsBdCxXZ4QBNmU+oX0GN8vsu2lueFmFLV48sgGuiXmhekTnvG8AVxJD9yb+XO6uF
xPBrCTwxS21vYy03op7Qw2Ytw/6o1h2b84jcgj3/tMpBfRAuCARnlU15gibKzVjG
ulkdbYcj7Hd8TZv3OMCZP2ja0B2+0SmxyTHcqC9qlU3uSTZv3nSGOBXrWxUFwgLC
I6CWp4xrrKSmDR/VvQGeY4RFSUVkAbic23dsRdfWcmjBqYr0iR/XWgrPrmHheH8X
+2OUaxmv6hiC9vdcR9K/w4KOEFEeieayaxFxITUb+eTquMO+o2n3NwKD++TKxoga
benmRJJk74PiCsqopwQIghu8eBsswySHtxALrqOA6HrYMhEe6BMyjY1NvjlJDoEK
q6MiT+Qxw7KfsbqROC+3ZbdN8FRxsQK45k+AzrSU6q6/PwcPt9cFuuHBCCxcI6fW
t2pAJYrIniieXAvWm5knMzWR795ZdFqG8Z45vCRJtBsJCuuex5EqkEYdfbWIG2uX
vIB3XiLmy9Y9IHG38lpOdDzmlke0RQiMyTAy6YHrN35T/rFtt+9xkGPcjkP8ogbY
BP3BKO88KBcJSGd0fdwgTAYlcG+ag9L0B+UwIISZYBBy9C3PwqMGJBoI5V5gnuBM
OFqh7cBpf3ayhjyyKgxNDeByEncbiuNjeU6a5ByCDGOzBOnS21xyXxpu8RNwaouB
UowslCw/9+Uts41ba00DVNzXE2BzONXSsjJ6zNhCfz/mTaWqDmNc/vIfIws/7sQk
tbqaQ8VnlAt1LpzVDUc2HkQuvSXSiI0jZqMUXV9t468gvP7GPj/da9JevpytjqUf
8KiWoGFEVa59N8dMkqFDBmEI6EO4uL9dtvM8CTmweOyDupyhoWQXtTigOQj4mkAJ
AkIgS/k111d8KOgUUWg7HapptUGhxMWjz1p5fp2QbR+2PG7R1cOz8jo8EkglU/No
O+3MKcOzepcmINcpspoSuvthBPJSOmCfl/nbqSPr6BgCZOq3byGEVia6x3fdOXl7
fWQlaqRkm7JZIu3Fqrm4p28yH9upArTbBD/fV4nLyJFDu58K4snIo0AOvtlS9SOz
ULPjycC8e7j3Dvge50ZvWK+D9LWwqi76vtAq8h3dlIXmQnlWGUqaQgbLsYHNIO7m
ImkessPteWQTAPdrsBx/N9hsTHGEVVamVlQAqum1aUMB8D672Q/wJFKDIA5x0gt+
0R3PMJ1GRy1oVoFTuIf3ayUSQEKgzZWWpOEke7pm0n7mQLXTk/CZd7jb09I0MXXY
RcoOMLCeSJ6f8+ea8LlN+dXvt+qeSfqCMnDw8B65Jv17/FL2PfzB8HrP+LNb/laT
t1yPR0szcfW87zB+PvjZaQABVOYU1md3+UX//PEgE77Lj894Osud5yva3nRN6CCp
3oNrBu4GtLnotErUUwxTDlXGAl2w25oWuh+4dE/SgstXYjteFD1wLcnweMMDSqEo
URij/gjWw16Lc1FHbz0zCx2DKhUOjkxlZRkIyk7mV2bF5aEu8TCflgD6Xn+yxCJN
T7ZPVM9ccxraH0KH3nNbdlg2esvcKceRQHuws+McsXJIgUrvAKx5FlP4VlB4qVuw
wJc+5Ea4NI2KWwafqkS8wtVN2PezXBLFeLhE6c/1F45AepaFzI/5h822IWX8S5Hh
aqZ0QyaQvdOdPgqy+P5jA5MBJdsoaCdq8Q69ch/Y/O85mTuLVufISAj5fd2wMxj2
/x8KiBxSNfLzYATqR/rvFeTHvWvlGWa2KoAzqgBOfw5ix1dnMmx7sdGu8hs0/Ano
UWkUlCVtBTzgnjTVMyrFbDZTrWJE3+4nyIMel4GaRS6HbqKZE3vYZ+rQYgfdao5m
saxPX5VqSVm0CC19rZLLUCWV5alEGcMXhpH3lnn70193ewfW2ytqiytEdwD617wP
uZzUfafjpdMPMY8AEb7oHelfAjfQ3uCsq4GA7L+ki4omI58/Apg3K2DKpRO0wpXw
YoCUgJEEBZ/N5LiMg2issYMoS0r2++A7P3LeJwQJ3yCBq7xKOw8FcRTL8Twh/aoQ
Yga86KsELW9t2Bi4S04C1vdAR/8DVgEYVRJRDqTBD/PVBv4pHWSlhX4gLADB9O0y
mUWEvJpWC5gf7HJecdPKv2ThpQJH1K/I8DKe/OkYUuuunU7xfVPKZdZPQMGLj9/c
gxNOFu3WJlhgToe4INSnLMnU+gTdb3f7fEZGR2WCIcC4bZVkUscz8bnNCQ8z5Hdf
7Hh70CY8egfIl+Gx/csBOtFc/HmueLN041gVWEYTTcj7EkiZKCMm/8lVDZhLCFzf
d5zTCGNjhD8OAc/AUOqboDfh3IuqE6C0txomlAwJ6gvoL66lkTTuZbVfFgPz8x6Y
fSWpMpkxXZ65EncZUwgte4Qt+ZlEpP0CpV5RXNV7VHQq1/5WzoodH3k4tud+/QVz
ohkGXuDMilIGYJeda4KTWi5P3OCH2yNz+YsH8aAQkit+vDR0HxQg6m614rvxw8Va
AFJP7qBNdjfKhpaAg/R1rwRxlXZNR2NEM2E8cItUt2Hlz+4ypf0/wQ4oJaRrOpiG
x+SMi69cJKPN73o8IqyBBKn12xhUh6iZoVyK7WWzPlWgC0+En+zXfS+oRx/0f6Of
kl9dYxPgzVXJ6tj4hmEMQJ0Sr+35rL0+oyhNpPOxc8Una84y7CsC5ThYf3YRoTkv
ekONCVDTZbG1G2piMag0pwdFRmCUF3xiugemrT64Q0IwWvbaQFcZ5Rr2iISlmqMW
uyKByazolcix5r6MO1ymMMDc49J6fwHNoEgi8TUKervYd5xMBLvSwph1cGzS5R8o
uHF3hGW6SPYgjjodnl3BH4liCmnd15o3fNOFolaIZoJn8YkQdwJLB9lKYXu4f1RZ
fVcnjZaVKX46agTbva1Ve0vBmwTDOtML+4C+2xrW/KgbGV0JD8togE4MOPApr6Ep
VFw0s0FeCtsJcFM7j8LiKpuXXa67DhtGohcZ8tkLxT2jvZI6g691HNIs/tT7w2qw
bXCBCzgpbjyNzzsL1Lr39nx1HptwM3GpRZgtNubBn6VcGBNx6g85QoNCIC6tjttC
SsajsGIX42qqCWh13cO+P1gu9NeKM05CLhTR+uNNVlUzMZjygGnXv2iaJ4ZA4ekF
liR2P4L26Ija6OnqG9fPKGIEVF6Aqpplda/ncbp4w9wvGcIg5pKG2V2Th1OI35Pl
fZdQ6HsfVAgX/B42brV2AEzjf3bWW4frUbz/YkfzRO3xZl7wBVTqsVyihHTmW7ov
zIym+BRH/Gq4sv+gQDkHH1iPa3sLmmIACcm3ira13wFTHgUE26isMx6aig5S4rYY
InoijDSJ8vmRd4PMG1BAsQwuAgZln9gX3YvJMhzudPzNI3arFqBQs7Ib1hFf5u8B
wvfcgEUA645GRnCeqUUyZEVePLXv6Cfn8d1KKhJprGbQA0sEeZHT07mrNqO3skWi
M2JLWzqxyIzXpOccF5CmuUhnsLIFoykDtibPPOk2mmvu459Ob5ceH6Z6b+/U/tFz
mukZ5eeZyQj6asnxSrM1y6bi32WZQrtRSmFy8IXbo9Kpm4afeJz7PFEQtcnl4vkt
PjIvuSsM5Js2NqvxJfkZkt1M6tZ3Xl7oQYuUsSAJKpq43Vq1SQygTPmJrlyaqMXa
ELvETk0sr494oDsnDI1S0XFVYuYhsrW3Ii4DfZXjmLbBZ4t42kOjIehVPFF6aiam
XpGATgUtC/wU5qp4pMNS/odrYrfmE5kAdCJQLi5T/0JxYMndYl+qVTG6uaq33SS9
zufFWec1tiM2p3wldMMMvRlkwBLArJHNCiLSa9dRHyCIz6TsYKmvLLLpS1JCmTgs
EW7idrMRK5W3HjLJN3uUsLpJjArTGLBzptqKKLfUSLBb4ytYj0e8tRFDCFfwYa8X
ybadx6l6XJj1ZXiZfA5tbFzO0CpTq3Cq/pAoTze4RcN0iZMrVOWJFF2v+UB8hkA/
8Zk+K46ex6/Z4ASdU1mRLk39YS6BjLpAYktm5bkJuVLiGknn/N1dVb/aYxNtIfrz
IwrnHZJi7fTc1EXQWOyuxat/V+hWnUZwtK7B55OOO2dUHE3768R/iFa13F57XQNU
Y7GmVH0NSeGVJQJFP97eCUBqZRQ/CET6uHTXd9++DiQ0uLdf+1AvV4PIg5QL6iS+
Sdu5bsAo5TsxGRjLC78BuVYB3zgFoNb8RI4YcRV2FUVmPfBYRUO86Ch7sWggXENP
KhLFEIwShlHYqPzpS/VPl9S2sv2hCJOH7+HygBqkAH0/CmEtSVk3E0GHz2qjNQi9
qullZ972Ikm1IDkONacZUHr0AE/+OHiXqfieUSlSIuwB2YSBHFn1VL7XQdeWSRMu
zr7M3sGBaeggy87IiudVpDBHpHDnGTcfTQkpAmhCAazM4aUYxT5fcbinQQFWrC8c
+chd9QYMwrFZnGmuZIQd6fv+TdW/1sLfl1JAlp/43gPF26wl7Zx2V9XCISwsBHs5
oTS9GBfusRraJH6Wqnzf0PBPz4igvJH6bqk9Is/qOzz8PEm9rfeZI3GR5Mk7s/AJ
bD9f1sbosBJ/NEn1EursrXsxhb9QQ2cXgPGWI3jlVec4aBgLoS4V6V+LetoVJjGF
R9zW+4wpH2dUJCa065eO0e4KnLyVouS1W73Iv/PzCm/ayROndmHaB0gA9NgH0a7i
yzjIRgUEn4bRU3f7Sh8PloGBJEZN+HHMLy8qK77vkBcz/DWNYdhK7H0z1QA0W/Z/
OzQfC/9hLzXrA7mJP/9jhLwlUVv2T/yjdnS3lVDEDV0AZ4VZU+Zwn9nElUQbiydX
AwxzHRqfetTjppsNOraOtoebhUbagrvI/Jy/q05uRc6TivQDbmvaNWpBB/WYvZtM
I40TxxEMd052Su2Ra6BlLZzFLo4u75hwfu0liJjDIh/hj/iLp3Ep7LYtutN02pWF
sMQ+d7FmdctYdqC7WGTD1mxYsoqQ/AhIzG9+ZfVK8SBLSfQFB9G31wXaoFiLoGFm
W13VIMnlzWmHgfeNjG3YbMT/wMMbUbH4HoYtTrTqxfzby2cIE3PuMck0IjvOr6oC
BX57h/tyXpMUbwGNYcGUE9GvbHUY/9tIJ2bzLoYNc1sKPw+4QVNU3VRvgTY2vJNu
7gGCNsetRPWMC1qizLo9YKyagiSCEYp29DKaYY8QbMtDAFzvUNrRbx2kSIeicQy9
AFqWbOQmXs7wS++GXB8Q6qYVTB4rUz2kmXrET2Vbvo2hqfYnWD88CGZdBa98nQbX
RXTyeJGSGNbseYEU3LUnav0C0n59k9aZRgJbCT89K2InoV0GHZYq2otRvneunLVS
uM4aa4evTA2uwTdEr2LNBLxjvWPOaKfhRMvUBZZMNmJmvzPq0NFxxLkoObF0dx6H
Ot9/54bfI/k02CbaO0IbUKIHM2KadpeJbnNBXVKoVHYlMoowJt1K/a34EU4yGuf2
5tqMvLtbyeY2CeQNEc1GiVGkuRCxXvbd8wBZ6p0kMRl/5yTYVASa13vrrNc+uOgo
83fc5sfFZsLyS+goCbRDozCBIkq+vNajNMFjNgQzDUyuXnYgI80wo8fNN3FoR8YF
eQ6k2f05k/CqrmmXOlA8CVLVhTzhB94aEXX7rPvIpR3kBqN1K1OSahk16qrXw9OV
figXTJdL04Tk/dxu8YlkSeNHqQqNEBnr5MOKp1dWkqsN1jteM5RAQ10RxqjLcXOd
JJQPo/0DKXfYyNLKUm/h5C1M6oqipuLmUZOBKiAZhOru/w/d+4tMog6eZ4zri9sP
pq2LJk53PVW3KB82PEhK7wLD+RrRwxuTuGpJlksjolfHXp34FyFHSDgmVTk6LwDA
ex9Q9TSGexHFl0DYDpdZLYH6/dLbzrU5bsFXnMXKO54jQbA4EIaegzUW1bSgPwbG
KXqjSNgGuIp5s2VeP7W8y6A1G0eUNQ7HPFcTVeS7QeMhjhVQDfkPQ2pVQLcj1QzD
+nWvQXM/xs58vk0TxE0fKMdVicDvX8SZs4BumT63joaN9+LVAqYawuLWmodIqK+6
pbzbqLN7L4Uc7LVemFQvpAJKiqLYgrMnpI3Qc82EgcT58mfviGf3coryQ5fTVu/y
Ut9ehCTPWq4lu9mkvgACuhuDR23L9DbxqKrrvcnu8xrT5unELBT8V+eA/d4pRWbL
u1ASz+xYXh04jzURWOLUsWbhJZDbly5NsY1FJHaciBYW7oLgOVVc8wethMmehrJQ
tWi3EPXa3s0KSknvoSDmkIJ2WuiYb9c5jDF4HGyCxzLo7X/LAfvmG7389QvUmB3H
XpjvSgpksLVNucQLU0dxzEtk7OdaqKIYAEGp+r5cVAn1Yr2kFEKet0dFamYiAAa+
2KW3Zxo7x3C6HLo3b1Mkrzyc1RMqERVM8/Nuxs154n7g6vUeNMHFheuRJlSitlR1
W5xgqyhLWo9XPriYKLRj8Y2h30EK2gsp2ngrJmIVmGfEVPF6mbNeblc5pM546nwJ
N568vzPqgoFQ17/CQKBoa+Bp3zL/p3NUlOYoyKvOj1cFSSAVWHCG/RLtz+u1gLNj
EuJvRN30/cKGBQMfsBkM6jUfA/FoZ29IBW0ji5GoWFsdRUKQ5PcedBnVYEcRVbtl
IP/hwk1DUG1Ttq3VAxDCQxzU69mSbL9tg+ltgZL7ZWKLLXzDmvVzA1sNgM5gBKO3
uqowYXNsXX30wnE7ZZcGxZ6ajiYJy5vcgumX5n+qeVHaA5+096+FRVuorVLSIzcR
NS1e68wUXmtS8jbCvG94RoqDunCdmR0bd0lPFBCnlgKS5omt+rdxOAYKQUzCtcBB
CwDw9lPDxHVFfAlDt57kHj6OnzuBWWHisRp0jiHn2j84k2Jh61liHD9hj7qfeML8
ge8kYsRLbWdoc4BMPR1tb0wCt7shcYZXRADz0R/Hd4vbkCNEa91lfKwvrBNN0TbF
UDgFUQox885U5tvonzBxEg1UdsP0j7y+4A2CTwIAr9NCqCVyyWHaChrVWXr24oq1
zThjpuFhd6PbQ4vYj/oWuPh/ZI8egRC+kQRcVirBvnbH7obeE+JAUmlgLl7/AgHn
UBonG3ohwx9H483fdEJYhGljcSpPZKZfctsWM7hjVy+mTMvGyIBwtANZrLtaUmbd
LgIoxNv4G4IacPvqoiKsi+egjJxwjNGZHcFOeN2mZ5fPaMwWVJG+8q62jMFQcoM4
QEqu4C89GpsCTVlgb8/pWwx3cNXcn585f5DqqFGB9/1ntaplOgpfBb4PeTPZ7zrj
vib5x3mQtAx6mrIcz64DqHrt2enKN2Tc76wu8Kcc1MpYtXZuga0MGtNmjXBL2ecz
gtyTxpY42aEu30mEdboIkAkyeK7MdBQ64w7zUfHh9E+piBR1O8zOU1AOYMoslxoa
4GUk+O9RzAV5xUOkqRhhqQL8emSy3+NvJ4johWdsmQt0IJfV421LxbTyjBef9OUn
qvrRGkmWWVmuDXswM9v3BT1x1l4qSEYP6GYU67a/xHHlCXpZcKKLd3GblQo6wv2U
8AfZzH5RLGhTPN79z22BTDPnafA8CDgUEhjQ/R7p9WcjOIB5xqy5Fw7sOYUpCc3q
44mJcNAvfpMXcfFFX5b1U+Cs3z60rwEMyvYFYDmt8dZk+wk0G3FENQH6im8F4VHz
zyGHGeeB/0Dayj6E3vn6U0I7FR7OwJtt2I3164KUiphLnRonN9T7bZz6EslGFrHn
NMeHNqNTXGyHiwJWdnXFssnxXDgqoOujGZ8WYIL1wfpbOrUlSF1y3GMrCGHduHAe
RsbQYbg0BQaYWo9hdjZFg3mik0RpfLyv6oZmqU7uGiN3qBma5irOOzYT5yCeCFWU
RnjrYc2Z/IzCVWjoCVuMXJLmjarvfG+n3WEvTewdQ+oW8gbdb5kI/vNigFHyEr8W
4unJm7riRlsy7pM7mayCbMfCSwIIU9XAKazI8upbib0l3zBwT5UFMQMP6Ibex5t8
MU+n5dHrDz3beFm9dSSY2DlkJ/lEGaaQzvfv8D74MsilerVF64OzQUxrzZpOh2oH
izYAZSSX5kQ0ikywNwF7G+39QYBQdgjOPHRi+McDuboSP81Ujhywh8mwsnCbhNd2
IOHJ8LjGlts0IoLUA7w2RS40yeGvTwTxVvEcAQnK789Mr0q3zZd3hBtn7dInU34r
fQmmI8/JIBp8vVWuyUm82eXe8k2FqEBQxYyQQT3+OO0mMceRaiIEufG25mbTdKgT
4O/7f5umTt+dw6eCQomDOU/g+TMwcFDPslwC+E281vWuTA5E4WzqgfLyjy3DlfpL
WIo6FmsuQ3zsZ22NKJwJA128FtONRiuwFCIYeGWQGE5zCM27ISC8niPkJuPoKAJH
oICuHqaqMjmkbaqaTqgsLji6zdjUear8MxsaSdHKnG5VuN96/q1mDaO+x8o6WlEd
kT9nMcqyb3KGiFr+PQBkr5yv8rzrLgGjR/7O2Szs/ZhbOK2z3f4vlPL5px9ufy3e
AC0GyagOz4BYOJP8qtXz5YM52/2ZjWVj7AqXzTTKb5syqeUamzYfxnZpPPio3wMz
e2brCUQgzisogUQqWRGh6T28ipL9miAVdZGq7CYgMBUX72u5eHsQ0kkYNUSuMTwD
dQWz3SFDOMGH15vjAzdTL/l5PPofNXxonPm4EhENRd0eG5eXgM+Wm9ZVJpdyeoBd
3CuLd4VVGwtUjoWw8VKP3Zssc5FM9vPSfZzOdlpPaF1VhThAqiLp3uCbwhtGuoR1
+LWExv0D6PC3sGNWgHNUQ2FB1wtlwKP+SsGKTEUieOIYTB6wmDOFZCVy+Jlv7lme
7thERG4kNPFZhlHSASC5vPHXzdhYDky2ScBYjmCRQkod8z9ru+yZQ2PK8oWAYZ9P
DzFc1xI/lioEXdWmUIQbo7waBszfECsyhxXUR9Houv/APnQHJwODbIjIKC0/Dyqp
MbkQXIHb+1Ll7ZjUa1CLrmRCdp0jaD9OzoDClP+l4aopWX3vuSBKjz4gdhta0taS
t36+WeSf3iLgrrxFTxv+LMkYopjnH+zCSgdHyM9JrqB1pacJxajaZDshtzQGoTjf
hyfODazILqKSSkPm0hnj/Ec44AdL0J5yAvWBGCTzCxfZBDsOIsJM3Z8iS45sMs2z
7EaqwlOZnAflVwXdy9yNQHh/LdMH9XIgR2Vo3+YwHmQY4Ai+GOqGcPlCsQWEY28o
r+rZMHFrkKYDAuWm3qsSvOaNK7yIGTGzDgOSu/PJiyEUIedn3FP5G/k60+qNIJTT
1AMx7/jyL/n0+PeAZ3H2zGt81eaOc0BuC2YKCk19NHpngIESH6MZ4eTb5jjWpU2K
tbNm++VfNGfX6ycljiIt5DoHPa3yYDslM48JujTvApxxuVmKIof9HbxPtj+9xXNL
GtLtH4ddT5ii0rKJatGfk79p/8V2K3YnSP5Ju1OzyRAogzSmleq0bfhRz43Zy4MN
EXMFVDd52ptUzZOSj4P08HWZXSjBty2Fqdot9KRTOPmxxRAcAIbQGPl86aPKK/e5
2gYQyVmPJqnogEWytw+IFHRr5xgq29G8+jOPuYeTTxbblP3mmt3VEOuXiQtMKd/Q
YkctukvEprUE/pccCR5hYPsi+UE6Nago70NiipE4olTd19kQq1hswSwnCBEqMgRr
2/lYq3OLB740RjN0ojRKjokmSJAxDatyxbiGbIZ5rrQVxYdlxhxN/nXj2Cxxfc0x
E81OwspJzwfFElhjvCaxZ+tfI1lmKT+x+6tpq8W+AaxKdSpbu5qTZwPSrkN19iY0
Y63Gv4ojIjYFgHmZ7IUWEaaT5rFk0eP9PpRUCnEUFOI0SBoKonqsxJIRJY3Myn+Z
dInrpcB70QCZH/3vr7NDXT+Qgio5AVEHJlC/ifWeMw3g/eFmUxn0u/rGtbRsh6uZ
Rp2grCTQcBOe1Kq8cJnzwv5nfmnH1s7WLlSN4wmi1p7q/WI3X4FFSaRTg9PSVcnK
8AsVi0dWu1Dzyh06DXwAaVpC8JYvag9wHEi++hwAbGwhH50qEiZlzkYwAyN5qNRA
0B4lukeOq/J2v8V66zr9RgMFjLhqLOd2CzFPru6uWobxw9f5C7WnGBEt7dg4bjea
QInP5U6MNAh+r3NAIrMe/MvrYN658/zbPYUeIM++8yGde3ojwGS8caarslc1GWo2
wivDQSLDQs9TO7ya/VYbNGbxwbG9DTbiDYdjRfYqWExJYEkv2tfJuuaUZr9uvbHk
y31BRs5+GTNedP5+2DPdkgG6GxefUCL81XYgqMq0On1a/9Jdqvylu5bAXXioXMzL
Kc7VAEMxNt4TClHYw41rz10FsCY5dADpZ8Bhy6EMTTTs5YS6K9w5WZfBXJ5nTHwi
22lgK0brSDXnUbct+DchVRkMuEwcCnS4ThnTFFyXbMFSqODhS4IAJ76xh64bDalj
0z0BMFYWYo6VXEnSGDbeIcmmAorEGEiHrCADwLYstUieDGgz6PWKF71vZU+4EGdV
B9t3rr6hFBsQZ7Q7FtBfrJGb3GY+Apy4xOI9HHiU740NdIPYK5AR2rgAo6CJOSso
Fgaec/5vQymUuvIzx7DCBrkfacZPMamtbik2YlFzf4JyjdIHYJU4etWBBqifJJaM
L7y7kT0q3t1KzTDDKDygGeSJPH68rIHdxA+/4i3rw+TtBO01xv0yau3wsp0MefOK
XB6byq29/YK/f1d2vG7SVgt44Qq52QCVyc3umtpzg0DiqtJdHnXtQuhxFBak5kSn
7IYrCRwYk7UoZajTo5edeOk8REEaLf3ieFwgGA8Ew1uA3gXoYtb4aScalF50PPlC
ozij6DU0JMumhCUnyZFt+ZV0ZmfoQASoB/L6cBuV0tniX74S+quTGHeZaWMU27sm
raIj3UkM4CXnyFWMchOH/zkKKj61/nN/470/KTfOKwPW1PxlBcQFnf3z7QY9uF72
No1pD9IDW2zGgTfeY8/PEqtXy9Vnvf8oQr0s99TM4Z7SvMxzdgQjxWdaiL0KmcDv
M89hwKeH/U2teb6wzBJlOs/vNlJb8bny43X2LFunRcDDhXtESZnVKDA3yYMhKlrv
99m2rY35xUi+e+0HLoaKzvQ5/GhwgEI1yiKKKlaWgGtEm/vmk6qTOUE1qy5RQRQL
/6sGn3MwhRaC0m/7K2uf6QxyAtTCX2ZkcxC0wGIFga5rkCmmSKOn7y8LQ7SSq9BR
YpgIwypr6C0PEIlFo8RlaLvH7EC1XU5w5U10vB7ybMTxgpC5yWNQuWmNpWO3+CLT
Nx+SweIhrbw67Iy4AUIOHh32Rj6BVaOHwt4NWhMIlb97PaGaE+7zaJUoEE9RA+lG
MbaDgNRF9NPGhmGDSASqd75eawoxSDkagL8tGEY/Z31keKUvcE3nENME75aa0fMw
CmYLiyQBCbZz14E0aZdHmikRwExr/XG9wv54malBj76WvXYhyIHpUXoqrssJfUIG
vgiKi5Vj9uVHfqmquA3KpYQTsDq3C+XRv/klBnX/ZQesGfeUHS/Adqp18ak1jwWj
q7BQRyzGhkd8VNRnWKgTBCG3Ury0u7hjnplbcQ6n5MsUvJMZBmiFjsFNh5nCq92E
38HF+e6PuHcxH95j3B4FiJjA9hQbCZWTFMiK0wWnEu1ihHnyH48FX2Xs6GwrFHJU
ldJnd9xpxYO9i0Yec68ma9580M/32wqEdHQHl1om6xs3qpMoaPFSUQT2Kst/F9P4
LB2avbAyqAJ25d+oOuH+b1N5s0Hr7Mk3z5E6ALgX8H2GdO2jgAtdYM1T2gbeAp4W
DDuMtg0y/+YMnHKHIEiI3eeOx5a7g8denoFim7iaoX/GuHlDJDQu260raHk1eqNz
fIhGO8w3M6RtrF+Xf39M3woYm6YmKfQ9Pd9xLyhlUlrHdbZxAAyHxgLXRoIhDu2n
nOlN8BNP22YGwJuCjyqQNyERiyHAb6+xeZJn1iofIRL/V4eJoCarlpEAyuhnajI2
VmdHDgqeZe6cOGntiu58F8R5eM48m1P6ItuFllICriksL+8ov+Q9JI56o4qqEBvp
zkEDC5sRznPud1pBrJVKP62OZhvLYTlsUj9DmCD7ghOqfiCWBNvIcUgtGTQcz7E7
g7CNx/tWApk98ZaoOsE7aM1aF1ps33O5uqo+CL1OV9IthcstM8kstl1scS2clwxR
v4AlbsJF4l2SLP+pg0gedflqkLe8ay4s+uiqm3jZyiSfwAC3wR+RsTrh7gO4l6F7
SU7ogKekPW7yhZMHq7e/KU1sT7si4RQVkZKgDHLCrp7+RxwYk7e6gRru/OFInW6c
XtuzwtcmWJHxpeZP1mL/vFYTzWjDjT4sWl1cmLvYf+CawLwePTDVAsjKrdPWaHz/
9P+GJwe87BYyD0RPPtBd3AgWk9iOECJzkSo6tX9tsetXCApAJWd9W2YS0PDFgkdX
N/t8fnDFwF096FHoKV085vCcexHjhUhOJi/6oarPiIWKVrcPku0FenCEjvCQLW55
vdWotBNF3BxORz6cwPW4btKBD66PlWrhQGHH1OYWSN/pVkFfYGtgpjx4OvCwU4q/
iOf7dRZ4f9H77wt8LCF8pK9q/+XU887ePwoZP19gf0H/c4xAmn6DK9Ff98BE038n
AkoDO73M1L+VTVHIXs2nGWlllSimoQmPYfiIZVnrD7CXdpOfXE2gHjtgA6Atf+Vi
Qxyzzq3jh3OW36Pb7v+746WnM+n/aFPJkeMVU65B/m7UUyC0MHKF5vU9og9GhiTQ
QdxflLIiUOgP6lZy30wiKo3rwpkLt1EuGlUqrG0fni7BA+xwnOHKs1BrRcPPfkXU
p7TmGjiL5fhAGFC7OrtmniXS9iONWXvuY6ZryoqH0a5wQpuIwIpKEBputNA9B8Oj
ADuyeWDyaPJ/GUIgZ+4JImVihhHMPLvA9OClOzWMrHqC/9fnnlb61n9hlHyTq/on
W8JLaYVy5qrwkFS/13ntLgUuRBidRHoEX3WcDJ8DczOIoRXKOe5shkXQi44g1zut
cY8Blndqh+C8KXSR8FKbvch7POOEetrgO+oI6lwVVP97zlts5Qg3iKnoKWsUsoNO
DJhrnCGdzq21kBFfA/ngu6C4M2ZQF+ILkBCvRIKidLBwpH7dAGSoiE89KHgNt1/5
miGFui93hS9QlM8WX5UFnDlN14s3Au+Q5emeLFBCxa3OLs0mel/apXBd87ZOUgmz
JibKAvNi6GPeEav50M3ovTAh6e47Qf2I7bQBP1xpjjYsi1rqxnOfdF7sbd0O6v6a
8970O9q8DLOEkxwvULv49GQcKrHiaVEEbdpflM6wPQxOm3kDqHbJ5jYnblvYnNWW
y3wXa71E/VoCwqxTZwPZzbn/9LXEV/oWV/KZVV2JHcQCw60V+DQUMzBojmoHYJkD
ZS5f6yvXcnR0FDROdxBo+k8xK1aEDnasdw9WgSafrJMl0ZnBDTHJq+2Y1YulH77i
Ii8+8K+JE8T/VjZ7ccNJZBKuyK2uZHhwWxk/E073ah7Othl2vW3VQL1RspJamcZI
XzchP/P0TlLt7d/KeYGabAppAkbtnDr2u/usqPI5VUx6df51MRporTSk6tw6CFEu
tzygwIsq9qmJMJxU5nW/QZfEZ6glxllNyXuk0H13dlweCqwXFMcD0k8EkYlvXclI
kmPBvvglYZ42Jmi8sSMpGy8QM7qmS9E6wjkIGx4ihpHIu/XoIPVlW8KWXDLWl/Xk
+IlZHP6oJjYLlod5PLFb3HMe3psv9EAXsl519tgNt77e1TfezwrzJ91hB2xXDG7l
p2n/iQaKOnYUaBPpOBC03gR/QvrPoDP7vOscueJhR29BV4CXvb184FQL5U9hhk36
EVoj9SnNYOAc9VJdlG8hBp3bzVUuZplqLUDobeXcd0YQsM4o/3NABHVWvq58PMc3
VWJfBK9m4qbIXHb55RXLyfKXIrK+MBfs2HhD0GE+VpSlt75BXJObcx2v1NS0pxyF
jn5xRL2qd5TXYRJxh1F3MDEFRvvYAtsa5TNTs8roPs8/zZbmVYzvw6yaBu0DYOeR
XKSzlwqj8fpYusQgWta9I0SMDlo71ZHpMEe0m/hCHGxOsoySdodRsq9djFx5p5KN
i1s4PI04I8Ilr0k8psAClbQifvXa3o460lfUTdRArAjm/yueSD0EVZbh8vSc1qhA
V+ld5jCI0ng5gkJrnkYfTRM0cbrc7VDpXDtgJTXXn//VPMb9pykIWI+8hDcs3Ous
0Hx0/6cF5dN2fi77p4yvbLlGPiSQXmD7rDav2jkJ17Qb8akJZMGe6w0J/27esJIo
sp09C449upiNppzxsF3sG3PpQ7jbOjj3gShOjtmMikaR3HzRs+Ws6s86diwon997
zC2oyxfDxXGRpxG5XuBp//+w/XrdmgBilQk4GHe/yzZvOvNfqD3+b/rmYCLeiluq
6SsI3cUyKyGC2JhMzR/PI2cPGXsL38WNgpI6aX7pJj1H+ZC0BfHV06UfOksFxvzV
CgZNxsxFwJSHwU4D9RrW9oocscikQpvsav7vaC+AQczyzD7Ilzj8KBkPrwO47Qi4
5rJLF7nQp7d9jAdkd6yusM3BS69k2KepneUjzAPOH6CbTR5KbrcE5T4TCwsiUmSb
fiMA7fLti8W5E3H9AOUiq5vYmFLO6gxa9PrG/pPMZfazoVyDstTgPNq17mJcUPjH
BE6dBLXh8FXLLlaCgdYjQyjd1pSNoJNO+bft9gBDgDl8LZck/uMFuUJezUJkWngF
U/GxfNFZ0UV1NtkjPaXyJchVhdgUPNtnN+LQECDeTyLFPRxK85KqaDXVVNd1uiDd
xXnMTKajJ5UcCKTeQBJhfrc/ZoyNG178p107bomVMocbb0j/7pVuKLB6sqIwDQiE
KI/j5JNzHAR2Cr+GcsYqAY6DKDLoGh+7+Z8Q+dT+iOzOJgj0YUHy1dHG+rzHrj8v
gh2pnGzcZQz40m6u9HktU72KAQUWbIRoiUyHXt1Nm7WJRyJft6EnYGJlaO8SGHYf
WtTI/NX7vdCh2129vrFzwAatLI1dlCmVCtwNaqZpE02iZfaIyb+FsKWgCFPwoGGc
4jY/5LGMtGNy6h1aQQTKFbeSOTaz4tSGeN567EmMi5nPWjcEIZCgn3IDnrM2N9xw
yv+CDACpMC7U6PmU618AclHzqh8UTWoMsD1i2ZHCkfD2+IU8exRheJthRQymcbSZ
MEYACM2rQZAmUZcRUup1XZH7WPJn/IcVaJ/If3Mr4I+lw5VKq5F0gEfq8keits8K
FP08gsfaotoPYkgUzksSH1lmMRBlOwLJMyFVvKj/eysXDJ0EuCgC7tWyf2gnkR/D
3E3DUihOPlFokZ02HUElO52pDGlB0PhJXLhf16PJKX1uoHGvGlOAabHkocNa/UiW
ZV0KfsShTsLC/z1zCbtnEJCg9rzxKSm+80502ijo5GXdSiJ/a0/7leg+SDkXp7Ff
RTAg/TBzlbc1+C4yOmX7qQcDReIjCnhThEV1Dr9FOU8vWf97hkKxHTZe1mAFrq5h
ppapIjr9yxq1ajd/buMLU1W7evU1YmEYc+w3NqRPQzxC/r2dp6cvGn6jLTP+ZYF0
1/KUzWZNWRNm5hRAdcnV2GvRJafT5ellYLi9+VhoyZSkqMN+XhElc/HKKUz/8oGy
jWjOnZiHfqKyrKEO67zV8ZTADB9a7XICBt+zo3J3Jhc3zHdzXh45pPcy4wHosW8/
GmcVz+vBOIp1tzWJppdqATVQPNz2CTtcelNmMNbq24n4dISmKryuMfxnllU36dEp
UpkY/Y5TOu92sMMKK5mvsWCnI1nsicrYrjXFUG2eBiX+QcuPu7+iEdw2dOQZsKko
iBKdHkXzosMs9Z6nAkJkwg9alOxNZX+RgEQwDwkPc7Egk46k6ZZxI+K1wSMW95rd
MarYLf8p7KXNk7OoCyJKiIS4CGDJmRnuKo/pyOpy3eIgXPyIQjyiw/YMW43S3TyU
MfavVlolGBroWIR8lbWVrhQ3qgkzqV5tQzp68Au/Na6M6unGOjBQ/QdkH4i7VAM2
dkxA9M6VNqdqRnfyPVPU+RQLsqLNaVxKb/TmB/JZlG3MhLD5zd9NohKL35wjf/fr
4vDWWoGAFA3PY1KI0JwA7mENIS08PEIJgzYnro+3ZATVzB5BXOVtys0EOEjqZ/vh
WmHX2iEKHzHvWTlkzRLYkC5hWVUn0zHaOx9yEQYQdAWRijBiD/ndp0AQ95/Vo6La
+ukwyEr7Eg5vxAFR/2SBLfe20M89dwcMKroMhByCB1Ok7ccJUvvSiDQ7hyUy9B+o
QqrW5YKrt8drTUueHak+mtE80PhOE8VjWLe+0jeHOEEH/SPiOVg4W9VKUu6B8unI
wE1S8eErRl64b72tKAyliNTrnVAxeNRuAiMkuMxgNEGGKHCnrLbWD/D8/um4ArWQ
I+UrCjo7b+8iKVEgO0JqrV01grT8XucXYJFoMfp1tEKvdjO0L+7Y4to9wxdoXBvo
BmUYka5w6/1EXLg6d4brYaULZkvrZ7jSPcArPaA7DvkgODwhpIUD0Zzc58gz3KKj
yfW+Bi4b/l6GbbiFkuctWlGY/Yr02w1zaQ2n+kw54bBLb0YjLYqikCs/0Yqigkom
4ctdhlaQSQgovt6zvB6uEhCS1bcACD2ifJnvzktW+EfHXyRnC93Yb8aQsD2rP3E7
hSiI6Zg7MprkfT1ItNCPvPquZ1yo4pYPvm8tKvzGcpXa1kd6r7oZA+zMRD3ovbqd
OsERByH20wrUtNiSWf1j40Y5TlgP9WFd9tbz45XLB313tFqYe0RmoE4hWLFOvxiv
878Gnv7vvRlNNCDKCXGxElLPb43fQyiNL/SzfbmoP5tfLVXzL0o7huCcsVxDKi2w
D0NX03ElkxbekqznflO9NybGmPGs3Hm7uxE3q5+IyfYARQPWomksrkvL46xC9fO+
+vzgnqaDbdZnX6g4jZ1dhAdFrlalp7ihSsl74iKx88iavEL0bD3TKOj378wDmYqE
qUFT9D1q/9WnLVr1CCOHiwgzIu+bwxaR2bm/opcWJm3PK8eFt/KJmZtp3I1A9P5J
aefq0CF0hF6aZRhNxFSYHCaKO6ZG4Q/ekxQe/W4KytC8Fy6k6x3Ig0qYHlGo5qKA
MiPqdmIfUtBfc6hncByclhciSewLTF18pPcQe+ibbC1s0OgaRNCLdDmi5C+eOo0A
lgw0XTfxFcK0MIKgpYpT0d1hguURC68cbYsaFl+PiuO0ufaPqbDw0iFh76fvGOn/
zbYQfU6FqS8IdS+hu0hHIC9yodSBPmp2VHlolZZPSucQkF2d9yq9AIK4BWsQDeF/
eP/RgA+xwksu3oWl5pozh1XGmFVO4zK8nCKchrA2/rtYOohAXlFEVJF27KWXnWAo
J9ZgjopQef8mDMlJqmxESFrzT4qITClWcSAoL4fKRsSMAwiPbltiyFFrh/nt7IPZ
hTX83jmpbMyc1yssMYbwWeDzZD5muo+maszdtjEUclYDE5L1bPpHTjyULqiT9F0i
AHb90m7k1vzW+VHg8BDWkIbjAuW1tBPo7ec9cxQH4o9JFVTeAPnLEBxi37VAc8TD
yc/8FCn2h9ly1WMtxOAkgFKWBhhIm1QfIIFSJx6gq8TPIqps566U0OnqyW7GE37T
OocQBGnsVeRUqHufSYgaBg+TPCVqchp/XTqxQ6VNhM6r8qUR/oNjLaLbuYVfeRUi
Xmjb0EEDC3sJC5lJI1cXrAylyE86AjaIcuFC92SjOG52trHEUyHrXPzRVt/CVi93
eZ1+GemxE+OthYYWNuvrGbuWl1kik9nEqhW1Tn8Nr1R9kCQQYGGIKEj0V1JA2MHx
2h7WR8AeuwBTvIoua+Z4OlCzr66Rx6O2hufVb+pXzX3e/8Ux3EsJYhTAdG8OLeM9
ipcnXKPmsHdyFt+27QoYpkiOoDquFoVV1MUyyYgVypszfWBWO4fmtkH1G8ACLjJW
xck2KUKcj29ztA2X3Wh52aUVW7iJujgttvNO9aH4i2WWpHj/HkyL0oHtSfOtYLoA
wbARMGJJAM7g4C2xzYoK1uhvu1k0P2fCXm+3kUOSYp7F+O5m3I5i86t5K++wfAps
kRKEKhzgpuVT29GbJ0nlSr6SCS0mCq5KVcyLJNFNrREGNXEzDyg9QIpMBTqt3rEb
f6mJkFNU8ojnxWjSrF62GcZbGEXumo45IJLd0SFnn227XR87hPBU2H1qPUQ0m5i8
uI25vWLOGWiOWuUoejuZcURt3LBUBLPADVmkIYqsdFjPOrGXH6h6MgwdBSA3b4p8
t9DThrGU3vQigwebc03kVF8CS8vNUnLUooSGzVj4/jTZku/LZnf92HwBfeNh3Os9
PHI13BN7BLgdd5JC/8MInMFlJhCej2M/GRxLoLgGXY/A4MJAC8wfiRoFOcvnpXzq
ZpgnseRFR5Lpop7mmSMoUJ6nAV0+H3dBD1AXtOWV6+nA1mi13xduzTDNkywz5l/3
kkKv4hAoQbvfPagHWHnQKiXadZybik8jLLVkvLJW+oY7J/GZ0fOnG1XM73SH3JAd
pD6EeLD/DqG/Cs4hWlzuM3t4cmVyQygNK1j6yJpS43btBhm5TyZ5w2g25ggaVcO5
3gTPE01/clZZRE5h8nqZtPuP6yCNbrPIgZmAOsWAyTPuwZYYFvph2af144uYlvXr
YK1EC33gXHayxhtwKflCI4KC9QYEFLXmIsKc96Zi/MJ49dl2gC5WJBjIWFPEE0/D
AQIVxMzRtfjd1Pl14WesrBqZFTA7dlc/UUByf50Pfc+WXQQ0aTzFIRT1WEK88UVr
5U1mTo1OUNvAMOIMHsscFB25YtzHN15HF2uDwi/6TOUwHFRYQ0ZglYp+rQAGr0WG
vIvavnuy0oJzReui+VtLZPaDvIEQj3pGL5i3r+kPQlQi0Hr/SBJtdrb56il/br0v
NdVHSm3/hwuwtY4ScmYSxk5z9m8tqi+dVqmRxNK5P6eTDxqv3xR6laM+Dkf9k8hq
+JCUoj7EeZj0n2E6BiyUAV8WwMNOZT0D4IAy8LUE3qJIdrkoWd/tBjGhZliN/Iq5
92ZuuvwKK+OLZwiB2fqH270I8qUatqXo0Vt7Tw+hee/kHCeqPrmB3H49b032Moe+
rf08K4rE1aljIV6yDh3fXuGpgL292BOMdI9ukrbnfZ8UWfU0nPbSpOG1SQ0QLrab
GklZicZgBioLHZfiGOke1BGV5IiV+/maoKpWSlzEuNPDHMnI9iaL1FKqu3EV8ojN
fs10+VILBalAMdiYji1me4c8Wm0cTveit7KK5BBdO6wiiwjh7Xq8qhBLEbFQgx+q
BLtQGt8R4MmhrGIxqgSKvCKzTyUzC73u+Hglqoux1X8wIkWvr2NuYHeCEmBm+BoK
gAe4QWP4iO+tgAa2osjSZxq5LeL+KIls7eQD7OCDS6tUmnCJfpq/NubJlBVlXpdo
up28UhaZuj8cCWL9b505Pzh8DnWW1Ic8anGHVou0UUOohNvzVvN3nu1F8vazWTRI
1oe9ncNCK6eXHqfYxY6TGvQJg+rh83HP8VphDt/StMvgbRmW0ktPRZ8bIee7vjHN
R+11AA4VN0sqdPcTqfZWfnFxSV45EHMwvORVmN3XqtcnFWQbLQ41kibxWi/2CcDz
SyV9KdGQjUFUcxQAFsL9v9FFen//tOgtAY/2ThEJAJ2CwxN9dyKli1kAajKfkTIT
37nXPjdploUR432eosfhn+ZWFOHy1O11GlYp0RgPxs77j9SWsUFtwzWHfALad/Xk
eunD5teXwTSrh34pHj3BBzLTTc18jESj2TdEKZTA7vxMUpUvpm0V/P6KoF8zkThf
Nm4k4AxtoRbbdu7frbyRtD19+NTa9y+CVGMUeoHcVYyu9SSo7+rk+9tFpcoWzH3E
9o+xMaSQX1KYxZPWe6XDm8gm9HvfILKym2BhWC2ky6CrfGhqNci4xVCoRoiI7hdX
0kIXKSwEXOERB89dEjJe+UZmZZnbKz2h5AHdLBsErHu6ds++wYzt+8pDTdc0Fop/
RtIO5spCMCYnXenvXK3HWfU3wUupKp+QaurhO0Ln4SZUti7KsVhV0dwl4BGVzuwL
TKNtZCZpYxeJTs5p8yjfdcC6XqeA60/1IfkPiDQDZ5Cys8Ezyppqvewk+CiCEkPs
P/HwzSlLYK6/XOEPGZUyhSsSRYOz2P8oepGN/YhUpGkjkzkt5EDQQV5qxFkgOnd+
HIj0dDASHW9ATUGdELL3Be0DKG6oFYyRb0azvLxbzsjLQM2MWYzHMdZjnG0Rine4
Jgs0Eb/qfpYDds8xIi5MfgNy0t0fBQCTMyEzkNxiwDH+7e5m+DMFrrmzPC6dYhaP
QRGNswWpngbrSK3Ou7LwkyrDe4ERUhFg133+ROcUbqKluvQoCRpsi50ZvD5VZ3ZN
1r8zhGliu6dyoNlq6GE9Ua8/i0cStXDwF9DB9pNtvC5qhGVsR5ORijH0Lw144urH
FrmnBMAPaqlYnwyr8OBb+XATGX1zwXRttfr4rlTW+R0S8wagW82L6YAMKTUv7SDt
TZ0YTX/HffL4MjO0LFZYvQoLaGSpQg948G75t1ilC91LfEVkGLEvdwixV/WyrEa5
zgqME7XjM1n2HeMEWmw9COASGEsliReK3/m31koz6xTjKGpcw8NKG9M22HMQXid9
2qW4Ty1I9vSQZ92Pr6hr0yUF9CXZy9wVIB6oTzS4RKQEft61A0KEoCv6CsMMlNJP
Vkt5HglnGN+iWlFrvz9C8AsGBnxWRCEGY2JK83+zsa31/ngd4otMiooYKL6D6tzS
e4gr+MoyI5rmzQQVhYgLgmlVqGE5MPJTDvCchuaJAYlNzZzkqhwU+YMhnIywtl61
WdEQm+LvKr5sceLEdterqXoDpADgwOgyfpdeZAczs/tOSYwYw4N/z/IFb9UNTNzs
LOOBqPwksHr2uhqI7mCTdzzzjY/VA2fTWW6+6F0om+/YQ4r5NxLG4n1QCC8j7f2y
limsh9ew9R1CFfAcoTUPzM4HMO4GvNUGaQ+K6U1X15yK2sky5eGK+BI4IsC5RJpa
l61sLpgN6+hc5V13+7rYupWpGh1oB5TZgbkVkb/3hUcGPlapU/vhU/+/atmqOOwM
WMXISSee1kI/GyQCdinMWPlNwO0JPiK5qVftW86bruOrwSTDO87A0th3iaktrRK7
heScEn1KGjOGB3giuj7Ce78h4t/q3dlfSGovORa/z/Ce4HbZE67irc32j3nJfMU+
WTwG7a0x9WYiyKzX5w++OrvTPhJXmGf0/eRGWEfAMG3jRXsmlMUWV9oATCxuFsi3
HoeIvD2G1Sm/bUdMjnhy+Ifkj1qookQg7Z+dpBDZZE1bbtCv2gHFwuTZhtqN7X+3
x6EiYiHfgXnu9+0pNCu+IKrPiPJVfQPm9xrm1Vqp0tT+YKV5eVKpzrzNdgWRjcHN
/OEn3P3X01qEbQFbiC6A3YpU/3ZoWzq7H7iTmDPreHx8SwE2hDLYyeL6PL0H/X9e
NP+AwoB4kRcE5OebfxbNVMK46kfiW4A/4lABy9Lgkw4EoKZUGeqgQkyndrvPYG15
sJu5KBz5wjsVLOfOVPzqzrPBU0/axlYy6YH0uhkaSPSG3/XTzE7QttyghOnARRdO
NZG8YjBxE7dvNJ4bs7dwSdWjtozAvfsEu3MdVVQkmHkxIVTFr14bnrs4ShXm0n35
8LwlHa5RVKFDDGPEJr8MtK1Yrd3x6qSQLXVM6HZ+f940kAmJMkSezswHwjdwPQoK
Es/wLeK8MGHPdp7YoZu6VVZLThOIYuHud68haBR4vyAm6sCCmRtMv6DeUh2qo/yo
4FKcT0OHWXVFBTGUXDWmqyg8vZjwC5fi0E9Jd10PH48DO1IQlp4dC648I6SiC+ng
E6WPOhL58pztc3Ov6SDodgfgfCoi+fPZ6KbFfcTjOnHtPhTLOKdMSZzvJ2R+MwpR
PLMUTnMPLkTn6qAYeAav5MB0HD+GXjjdgDmmM860gijh4Bg+FDutC3wrzGvbh+Ym
CdkwQIhV4HiBzl+ux0usKmiwdPOT2Yqj1j60rjrH0xD3Og3HHXVgwLLF01Oyhk2V
2iJvhS8Vo8NQSrzGEV6w4ZCJYYw7yaEu/c1KQrrwZZdG7JylaB96ULriPVQnjlnv
Y4xqfSkaLLodJFpRP6K3nj+SwBEvFzseMlt3RqQXkuVBBMQxjbK7pHPvwDtPMLnq
2NYSr+7boNr8+L97cUROpor/1LlcKLD5tyYNbrlJVVUwdLtHxCg3bThaT9FcKVqO
h7ClFMT8n6ckS4VEVOJOayBBhcjjocDiU57LPqXFzjp1ywuD9QRywdA5vv7MTmXa
auXWemtruj6TS3Elw9TDcAPtKfSAaT1tjxTE2iqbuj6j+n8/TFoBiKnIeBHXfM/y
Olto7bAZFSUahjj9zxDXvin/8X0x6xqBJkyy78b4Fd5RFToJUpBMcg/VKNWgSyY8
m2c2OR3LEABjOrNQ2yqSIYQ6edqtFsWsthj5Up23o8pMEHS5Q4L1YhSJxZOyuUv1
z6vyJ6A/OsrF3HTxVu+e+19vjA3FLeF3tHwOwY5KTih7UVcYDAqIdBmkWLZtslOf
ylz307f7lebDdATqx8UD3eiJfbroPlzd2+5ZDj2zFExIqCCbzi6kJAT3iOsk006J
dUiGNEdm6XV53x2Xx/XwYw+Zia1zptaBgxqYSFFq7kpnARi7zApTlNaajuXao1mc
GpdHK5pZ+5Wzz0roMBwTEZZVrO3gpXBTO0na37kUMjKq1CPaES3EmUBuO+8rtu4L
HmNnMwt1HlZ8xA4kis+A0PqkXYUUPUNSQTMlmUQ8hCLK3qSAOlDUqPnv/9rTqhel
f+VgccWlPhlqzhz9/oe8pWw/PU9+qKAIra1iG4P/mlYSS96exhs8XDfUea17CdZ7
3aeTwpJhbsbZSM3fFRISRRK+tZJWtXApsT+Vjvt+WWfagM4sqn+VoCoVUozuAj7S
f4Ux/7EgLDCTjg/+728m6D02SNuHMPDTfcrcDRjvEEsx9M2LmhEnxacO8EYLKYou
78mtSjol7H7r7SVntEjj2PpoO1Fc+P39SbNjl+038oEclw7/jhKxddiYHfYXZhAP
h9OwjRX0sQZp4UPuTvqctwoFv4mmSEJDe0I8mnxWJKV1Ef6F/gX6U69nVZ1rkrqZ
NjTJ6UZQuW+I+GiPJjq09HEHiQ0B8RqtOIAenQuAFQ7rV2rDmlhHJMzaYMvFKS5w
J68afHBRr4f2QBQng7MiNVHVXEufbQ8kEs75XMaGwRjCLKk1D9qIk76/N+5uMm3e
4NfuP8ftiGxPU9OuyDnoMPHjGTRxAxvwRgt/6bgxSZOoP3xvrrmtzZDbp2uF69zI
SSdbxUdiUnaDWyt9bX8bUT+u9TH+WWl1x2o4/fsHvNmkVSaqFQK/zdPQwgRkWblP
LgguXZWClFWFA93TMCZXOiCVrZM5NqqFJBKPu9DJeWSj8fRtWGsVf9QPCQZEoG6Q
PqxfK9Bu3MKkhdBaDlfwH+UhDPzOtsnzXhN9TUtukhpMx5ag8d5yTQqq0m6kSSbG
qIKFu/Wl640RaoXk3jNsOLZKO5o61SmvQkSM3wiIbbTFQmM923Y/AeUlyugaRmPY
3b6yTjNb33lVTyDC6AIMbK1OSgSOXxy/5eGtWgi0z3llXowAl40ptkBPHLlzkL6Q
MKzXTfoe8czvTH5oRdMemaUNIJhCXoDuYTtk5+56vV0rmty3AF5yG9t0bqJdZY2N
TUZSC9wkz/VCGBV5YkWnCWQv59qR25vlR+QO9oMoKvV9AvhjFz8tl8kHdaHMSoC4
GcCJSyS26Cy9IRcq1ZUlBprWYBHg/cRm/W7H98aq32+/Avx4Mter3laGf5oL6Xde
nFj6fM4NBMPRLRcNX3pvf4Kr/KAlv8g7LMIN2WIPGKdltM1zOAufMPUapyeggJ4c
jPfQoAEI28OKAozAM8A7c9Oknki6cBTnLLbLi8AXyjjBvyXS+vApqtHxZRv4sgZr
idwFuCBDaSwKMLhMe2kWibvryewWiCG+jScOwJ51It1/+mTZnzv1Rs/z/T4lyUmw
sOUeXjUMxyGVRP7Ckh3SvIS/C/xxKAK8z6IUlWaW8NzHhW8tii9CdXLXo2W1lpuR
R54SpEyBzwGptCOtop447M77XfLdZRnyI0DpGnprA7mba1VDgu2E3vz4PCHCJvCE
FMOUrqUB7IOfWzeMaaFfghZrTHBmtRfGcdjD4f87qGAG0VQMu8XoXETc7AA4lCvl
QpA/ZxDaK4xSd6X6f0eyHPi3jF7/FvsBUAIfHbQoTI1ofnewaTDz0Mfp5ZBcRg3u
7+C4pNnYMQeK2kVRpc5U9iLO2zmHSQ4XyI/Z1vmFN4b+6Vfc42zdnhbf14POuv54
L/VmxUvOC7eR10H6iGBI3XUbyryTXz2ydeH5uMK/hchmWjFMVcsiEveojB2Bzitw
p894bXPTLzq3+GrLM0X8iu9rHdHj51HxqMyQqAOQTe6ZuukzX0Eg5TGQX2xsEiC2
ktD5+UsXRW95bS4Qn8HEF8cI3/2TzzsoTpM2mY2lCT9SpljWTdLTko98hXss1CqN
BhRbZajWWJLt1bLwNlYuhE+ABX3bqNbzwFZJ09eVinoXv2VmzZrABRbipCmm5StY
TPPCZ8HfFskDYpgh0Q0+uqfNf5tOX7ZdzCrDgjAZ+4oL/KLi7/4vY5DfvZRj5dje
CqK6FEr0gG2cJdaH475nzzzJkvhON+uyXZx5BajJ3oxib+l8qyqVkelcP/Bba8TY
N7JDlTGkz613un/7VU1ZdicLavFrBNPDHTlNjqB+6VsNU8o091DMw28GwDsSqP0w
8xi9m+2Ymo/lxjqAMHtIH1nbS+8yv+MZ1W0CajrcVUiSKUCORdkWXaVNz+XtMbIV
oamFOt+pLEZq4wRYzfLPFqgaD71yZ/4SCZgSBSmJbju9NurDLCrEMDslFh8WFe7b
5+N1V7fxot8O6QO5WxHEeTKP/XD9Rl9Jil8pxSwqY4vtl3W+Ixgzvv+vEOX0OdPM
rNC9NwbymgXmz5a/DcOzcBx6p5cSU3ajdhlNRxZzksiwgXWVWTAvexrokzjdJcwv
ULVAT8bmQ7jwTBso0Ei1O5HldHtZghuwOwT8T2eZ4OJFw+7jVOnFdVvzydEI0pgd
O/ZfskBTL1yqDNRDvhdoE+dsoFfaEktJib1UosqlxCVbsexXXXpUrLdoh+mNPjzc
FsclsSvodSmDCZdtObkGd/upKYPxSkhZ0pXpLL9RA77PRUO4OM8W5FS95UPB/s1t
kmzORy9fpK69dpsc7svNgITN6gX+D0Kz/qOLJojOddg4xGHwbNlaSyTp3jz5b4QQ
qNQx1TgyZB3UsrglJfc4gH39i45O167JDc116tZSCtFSiQx0tE/iBWRoGby/0GVc
1ha0wp5hrylSrfz9CisVe/RiFhR7U3Fuc6xcQ07WGfseCTHUu/l7fbTbi0rxgzc3
KKoosoRB20CMzqH7m8nFrI4+7SYyDdz2iqU/gvAWkdKk1bnMCRsYGtDllvTPr0x8
X/tHB3La5qiIerZMQau7K9MWHnaiDohCeTlDKUBEDn8kCWAc+VaIuugm85rxX78i
dA59puY9kc4aETqdiASuPDlaXyQTHxhr4IZfu1HCutFlCr+QQiFDkaEmrxxiHoPv
8PZMSodFV91DDo2hDZffhmmB9WLP5UVroL+rEdnEdWWynpIqfChRWwQAintOQed1
DEXKHpYdhaxnwYJjSQw1qZ9Iyf7l0B8hclyOecmhKBNjDGfYElZzug5cmGRGW06v
HM1K09sLG/xPGi0BggYVAAH1EM7AlDoBEaXbdQQta1aFtR5M09jCkMHkWY4X/4Ef
x59MbdUQ5o/pS/Y6ueGdCQkS/nOkATVqbCCKi5g17X+AqTWRMDea7YmLZo5RSThK
6aYJOcQZ1+Okv9zB0VrZ79pLIrbQwF/F30mPKolj6Y6eS+lm32zIz04it9s23GId
FixkAGxAJWFQl4ys9dlqFjNCssxsuTDEmnKt5vOOlB7iP9X6UxYXJbNKQWFmSSqd
Qi0L9p8eR2spSYxoM85DJExxatErkfR62m+xYqOoto33xrVREJjw/TDUsT/gsVwO
L+dBZGMVU+xPv5BOKjgzoFuN4GwJky4N6VZVjK4pem0NC5j5i5xma5YRWPZirG60
X9qUOy2ugLd5QfS4J4wMeJ7BAm/MmUl7Ckg94lZ7rFl14LKdzlPscQ/hZ+/gQn+L
t84uBI4Aw4kywWr4yAt5f+vDodM2vF/UCje3d+ldW6D+vdjGPaujb5rqeoYxZUoh
5HGLMAPWkc190LyStI0FydLHXvtRcuuitlRci7GXlqpyrXzf5D8d4WvmEqTk7lsY
Iw/fuynsW3UE4dJcaRLz/SITWPpTjHNAzbOlPmDS1HRpPVM5vAfdlf6WsPZjBQSo
+XB/pS8zifkHDNXhchQO/A5NiESuqG8hwt1JC1oyiBvx1JDZWVRgUKdDDQTRyb9W
dxSNfxziSvgsTdGeznzLeVPJe8d9oSfjBV00EYF0Plmro9fBFkm/121v3hOnxm1y
cU5gjSp8nX9uJZXjmJYiJeabCtdD0vjo5z4Lr/Lpvi5b9POJlrJk0wKpms9zi0tu
ahDRz4YCIEpBgXjz7GmZLHmjhBxA/VDHdnfiP81bGesvMODMJ/RtuuoUa+rg7sVz
4Wf3YrU+l0Hl5BmMsBrQ3WeHObjCyjqixYzw1gaZJydbalKgzC7OTEK/pV6lgm3t
2pQtIsCxmEH9A45gxA8vyv362HbqnC7rkSvnmcw/FFF3B1NDLldJU4jP2FsrhWK/
9pMmMs9wZrCqMR2cfcmad7WgPcZYCkvmKoyW/LkGu1fiaI7DGuQYm9julqg4OvD2
RHAVkvSEetDnxTRKqGYN2ohoTa+w6iQIWX9SoPnWHc0rYEOd4ePYZxJ1auZC8zb9
iLSWnHR0nBILr49cAEIExhHncigZkmu8lWD/qwo+Apf3XXSCd+nlIURMrv/cY0JZ
JkWApzzlDt4kp4KYzMynBBKHuGcEQZsoy7J/6GosI1opiM7gLR0OVta52WBBdzUY
wZ5wKpM1gMwsyHjzAQnVSLGzC9X1DQugM6bhIx2BOXryt6r/SoZw3QWokDvD6DqA
y/mmcPyQ/1smVLHpwb1ZAssDlMS41uW2EffFNiGtLiD+DADvK23d1CJmnvzefCR2
NdVKl6pDN40uYhrZyOhlkt5o6jhUvzvMeiLe36Q3zF5T8Pp4ZgCe0YwPfupxh56x
RknJtBMmSeE0+PBI/5hgl2W34c7OQt2kX22cEONcmr/4g6xKK8v8b4HpsoiXNrUx
T5eSV1xsCgnlHfMmnDcjv4jWLBfyM7m5b4w1u6J6qLCdc/FMURxEp8E81C5t78bM
0VH/WwMxggzfefL5SMVS6n0f3mag3l/GB+j853cEgdtXnR7HQDv8ZNEKq7WbYYtL
XjYau8KgrD4jp0SdxucCa4P80lVwWnmrluoO3qTYLStVVNJlrQg1vd/HXbAe3rxA
WJxhvrOT3+UfFhc34PEK5eq7Qy5zbYgq4XA0uAvGMPsrfhdL/uSqhddQ64zHIGgo
/jr5E/ODB0qSvMPJZdBkdhihyumCj5kYlutxEcwFsZBKpfBfM0T4+l1ikxViOHkg
WpoFPTkh2ZnIRrAUl9QdNTXrM2LYR+d6aclDu8tRyp64T1EmLDxn1LbPw/sEtSt1
NathxSpeQk+bie+dUCYE0DDpE1GtKGKvTI/U4rG0Y9ASkxZvQWWQdbAqvRKDqJbf
nNm28V4RxZUDA2NMPFGTyTXe2M8tMnghjTMh5tKybI6subNWhBicW2abQmueevIr
aLe7VqXr3TRzyG8Pxs2EUUwoyoC6znQ0ICmclFv61QXucW3yEwYoL+JJt0r3zdNC
RzPPDuJk/w6Z5UU0Tzsz7G7TagBjR4CwZCxWs3WMGA/Aqgvw2kl7/49k2jxjlO5P
ujfILPVw1fXi15XG7hoROPNXsayt8uMCzuvBxz1QdcBFQNIrXSNNlhSJAelSqhi0
GZu3KpEl3/BFe8l8cskYJJpnvJRiWM2nmR8UQ02B11L5OYD9A2kxs6uQ2isMZDeb
K6PdhCXJ2lx83Kl4y01vlIItJ86lNnNjOZlsobqyhkNtu2wIgWsI3kUrEEJQ6YHo
LIsbMlGvtUXf8yWIWr3AKvDgB2ugZFV6vtN9oYgG/ufj0AaqINCFTpLVsfHpFJfU
d2eY1nmH1U2vFYIxnWD6Dua3ooOAJttQlPoA+oS9jaWluW8/2ed0FA1F7SBBCrBH
wENE51PTtX+QLAXC3j9OrC39LomyBFH41B7PBWqo0KmU5pPs/6wKprAhfP2tIsPk
pdUwGf59IX0sAFDkdH4u6uh7b8MkFsUCTrbmgjvuq9aP/WSNGQ9lUqezBcBvmtUM
BOQC2IPVE8hMJiq54N+CsW0voGK7SvBHrLe6rItA68daey/9sKK4Q7uIYS42//hy
RInxxHL3tGRsXgLzqQ6pa9A9UgqnPWNmhSoM+J/Z9de1EvBYhOiVXg5N57uhps8l
gE4oxHd48MM+GRXRQ+23nbldRW6z5FpKvlDvWeaB4QR2pL/DLAiW/9oaCZ2dyf8m
zorP3eJfXkvoGDGB3DDBiRPPtdmyaRKlDp19zBCSgBJ0USHEtYMVATchFbWl04hg
jf4FjqFHcHPvk3GhS1slib4y6xhuuHIOhA7iWjdfjYR02xiFQt5hajDNOKfJO+5+
TdR26i9y53wg2FGL5hgUlwCKyNW2a2hauM9HBWJFI5Zi4QM1AhkC4Qp4OUDHjpFk
3fBLN2QvZICuJKnw4VjPA/Kh4zOE5N3OJsjDGd4bWUrBYvnEuei1mUO9tHm/1E4I
6b4dnVRwbtaOBT31fIGamg7oVs42mjSo7GFQIBn6iICcTbirbo4DGHi7Bu+2paBR
hpnBbTP6piTLwm2wHgZTwdvr0KIQUGWZR2KHt4ZLU+/sUpI2C/Wiqx3g0D1hMEnX
ECBMt2aZ2LiydFK72HZUehOgjxgobFrUXgkYV74aKWqaqL/OA4W7SNzbPdiRXqmF
10vwETRUacjHquIgOuxGrBRTqUVaxdqnpH+/nF3dEjAZuyE5VOYb6jZuyeFDVvgA
0lD5pFGFv473BCxptLTQ6zsC9p8R9Sc8uYKAxXGV4lzPLp595dvb1JrjuSFnqKk5
XIHBrWSSxlX3qI1H+TeHc72NmaF/avuz681GB1smoaEoXl3ZorwGw0y3FKLUyRQ2
u52xUG60LsO7dkTYk7+3V/VVVB5bVIl+TcyoV5617+qXQXo5OTO65QEwm708svmi
YbW6yVzw6uNE1GqDknrC48DlQFvrffMrD+vGjv7SGQBIC3/wfV4/flQtkhfPwwVU
1PbkBP8POPx1e0gHbWFhXisYt2aC43wY+1BeFnzRd0ZE2+gvFh2JotiesmyomJCV
gpbn03KrNyETIveKRwdKeXJbj0t4NcntqFKvpu5WgOWvKv4Bi9wDYGRlOGKQW4LY
WjI+tq9j2UbgQiE4H3lBlRiY4vbAgtXlXpTp50NapAWItLL75iuqMnklUaWNVTZl
cYbahGjhqtTGuiHpGVqnKGn1itEPPENS3WeSFBya7uuZBX9aRQ9lWMia8v1wjtkw
us3dJNYIFe+HBkwmjyq4OgqRbfuJnrBYqie0/oBY8qV9NlKWBwB5EgBc5etJ/fye
O9suyDwYFR7FVGj4uMFk4g/fUAIqGT1jq3qdfbmPKOR46wvWNPCGgvArxy9Ydj3q
yuqbifxpX+3vu2XDe7n+3ZrMnPZT4xWMyNZwupXNAvdzW0lPJg/vxvXkWAO+9FLA
JHgGt+AIiwHpBPnaCnQN0Yf4sEUCcVyBIKqpjb/EJP1KrqsCYH5xS93hX+R5xjUk
xS/V4D1Yhlpv+F/I5YlsUnJ3sDGuQIZySDmf2msjLo8TlskqvQGGSXmUSRXSMOEy
At8EHQC3rAAsd9oGd0C1Ji+mQDqDTgXXgp1rKNLDu47JnTi8jpeNUut3fytOo9MJ
khtSn0YL2yPFBkKI7AcqpBE4sxfQh3DXSXniFKNTvmhWT10rl2WmuwIx1QJKaR6C
gNh9Kvk5Qpj0zhYyfZEFjJWYUdRdt1KOUOhlkwn0+WD6rqeKQlRTiTtBumrL7gwj
sGVc6bDM7ozM2zY6P1pkUKhCXqDMVdeym6Fk1KeHcQZSJSXmk1DZjLGZdpfYDoY2
ihJ2u+sKPROnU9l3r2KV5AT3VuGuP2W4xU4DHjcCTEzM7NuX7c5g8ubDHpqfNCey
SSGLRzICcuzi18yZ1uHowRKzWLaPyPg4mAH0Wh+v0aO90H8gN3yeFTrWSaxfcq1r
/WXsgcUPnS7MUu4JWw5z1ROJU/9k+gKQgtKp7RAB/C4M1yuXTpFcJcr3Uj2NVSJw
PFO+7rvTHm8KGpJLByu+fG/vY0yKSQO3t+6j4judwp3lNsp8JpMTx5QjK74ARj4E
YZknmaORGSfN+5bjaG2KFfkn+nAl6pU43MrYo3pMwCRWTdwYv41lwZQ8VEi5u3fS
4qlWDDMpLb7/Df6BP+pvuzvmbYFcxq3NCyY9NHMJxvZcWChP5h/Cyj63p9Tu0K2z
apSeXYDssHeFt62UtfceOubdBs23APrcH77ie4ycbqXBno83J+iu4M4kueoRwe5r
OlOnjYh+cK2lfoImR8F9kJSGdMS261Lh3FZm8KhlrXoXQXAy95DpkPiRs4toPOWh
pm2Mt3NX6hS7IrSWDxkiFJfQFqyLHWP7BoYz730x1KTLDlAgtYEUSX65x0YWaC8x
iNLILPPwQV6RcqR0JUJw5GH9H2AgZiTQ5IZ2vehka0nuD2afPbproeQn2t6PohTS
ExuhESkTHvR9qMd7TBj4ZUWCzScZ1elU+9itJILw0C5FySvsemFjacEjO9lsV8KS
cSpTx0RG2B68dPZFVEu5mTPnKo8fZGN0r/mI1/Sv9jHUFR4BlR4a3gP7/n4yo4CV
wWY4XfwoGkxDsq1VjKNzjqLKeqylsONzS1Dm7TXS5kAG8wmvA76rMvHIyC7FCPhD
sE3HG7zA89UJXd7/2zeBRNecQiAcxn9FzmjCe3fNoWwpwDdaw5yGK5Ig9egLBXIM
8By5+zusXSiYEjojuGYfGqYVpXudXiB4dojL0dHNRolfB3EjZkFoS8jQ/cY1MYtp
CLCsbt1Fqlyr2Dy39KhIvD1mom5l/BiptQDsP0RGPG9CMN2uwgSHW3XUDjmk/21i
8mDwpmUdEMGMlS277sio9lyWesP7eGPZbNoCZqB+irLqZ4bUe0ECbsxX0RYxbQXb
NtUtG65U7lcR0uw7clL1RJcZbMoVUxBO5/RJTqfaw93EmAd2PHr6D9d+s89o/04f
+kUND+ttBQzdOkGFSswTVRH3zb+ePVexyO0JmMwxaMMHsaGd3gWZt67dDbrrv/UN
7+TxOVPi8AyZZ+PvMtH8R3iGxysTOnLpDPUELUK8H4U1E/i1FlCyD/uQo/E4Asjk
UNRHqOm5sRRjAO82EJoYOBfUJ7WNXOp2b0g7zENTWU12yZwhUk079RLvXscpiSFy
XgzBojakZj1jkYZHImgAT/wTL4r7KfcHHcmUJ5eeQa9xHlMbu5mwLeJtpU72roE6
eWalvXbbQVqa99T+jxxf4bmbC6yezcJtGHjpBdce2mo/l0Rq8Q4HHF0bP4YT4mai
0mqXywrcO5963rkcV8CwLrVeAhsab0g1aBmTnh3bWKVspyoIsYY+qGio6c9av4If
kPqEMy6Caz0lFczfto6D3f0N23aE7wJ9V/TX4S9G/h52WsZ/7K8+hIq5BtFKUduu
SkWTTYMmxKulsxB/Cc3D46xhJg0GXw5TefK/9+khxfW1bhZNlJC6TjkeQ7QQnETU
eNlbza1BvTjgVeYyo3BGx2eLfskwfXyUYcrprBGmSMqabvN1TrrxlKVmehOT3Hox
/oKuNxbEXx0F80xGKj/luxo4jyesLB7RjNlNogKKA9+b7O4jycEVrlPwswiKTKde
lmaDeVd2h3LoTDtwh9/LRajNr+Hn9jSrbOv667yRNzL60cMgH7o2wnRjB6Cpi6cX
fe9HPW8IgVXPvD465i9VxS1ZEa+isvDDBRe4sm0KjhKtKGDMx7rNP5dxSCvzG/b7
VJN94VIlwYFYRmKxCqHNSsVhJRpNGUBsz9+5NqAO6qfYPDGVrzxuxHuA83/LMadR
u0S82HwRAyYRKOQuPxfLrhC9QI7TYcqy+/ZVYzdfRu/RCA87ngzOuDjUi5guYaG3
0M7xJgCI9+Ybh5SFUbuaGgt1fs3qZjBztPnoFrTMWQwF2jCdV5eA649dxTOG6NJ5
qen6pd25QoHIYjCtRFYi3K5mCsKntLcI5D+L/++u+pSkpzabUKQ0v5uJL+whnSmo
qJu1m16md/vKMFL2VpcQNH8rOOd0G2BBzHIe2IU1hqXtW4U5ndrSqKvSDN4w5/bm
/yTeOg+Rc1oUonUx+aBYI/eVO2dnX9i4VSy4GWK5hjLGL3ghNe1jGF1Zbf7bPQ4P
rd/Ba+/3+YXnOVNwh+R3teI1+/uF5LmhPayoPAX00WGfNPICjrzCwuHx96vkF5/7
hOnb2ckGrUr9qTpca+5lcrVWDC/eBuLqKAzroiw1zvIfwTHIsuKq6sx3fLtc58tP
KSBq6oZt+b7FGvDaVvN9HYKzaJcmmxQgVyOIbWBmkrrWdIt69gTcUHddPDRuJI7v
YLOyiHzwAH/ighIjZJzufXEDoQsnUz/yM2y4U43xf28dC8S5Fp3Rm26JY+VKrT8N
YANkFdCETDVspNdckLkcPWW47KxwlAdAihgV11m/dpIfhFR+F3QHc47Qww2V+1M7
I0+MYUxDvr7J1al6PVGZZB2tIq4f+5Idqnk2q9Pet0KRxS/l5tH5Ooa+qufAln3Q
5qjnQYIJ4UFPCPEsZDFOVM9Y7kSp7MS5MBWt0Jt49vXq624GrAhkeJLq9be+QyoE
1MSX1OAFHasQ0fhrz90uVPGOHwtiF5Cce4VhJjPCBtDMFWIUg70n/cYAJFRWIVt3
m1pHQp/ojWTzaEWG3udSJZ8r+n+EKTHuiaC2WLeSSFmnEVUACCssgWPRcdBjhqmS
Wd6yXV16IeJokWNSpgnYI4AUHn2B1/n0fmlO4wV3vwVVZ3ReEPEdGGY5/plXIfyK
9FUlsI99yTR+u6ST7nsSZQoE11lv066/vXUEl1MFd8KhuIsFAetcdkbFaPGd3Ap0
2NTlG9lyVHmLC/MntPZOMaukI1TEPo5517FM0uu4FLewRc6xogfenl9/gbZ9P+xw
OJcGg314cl+H79osCq9syzpwEAAAZeA66SDYAcduhIdSzSfEezf+hb3hTtcmMZk3
rotm0jWLO2+ScllC65dakpZjCzdZkiMjoXP9UfPD3LjGgHnMj21y/eXemzAe/PH9
osBFyusvhLC6lUDeDLG4ZKrn1u5V+WAdNbBOSsH0y8PtazBVWtrYpq8otWKuwY8o
tfaxHY0h/H0jY9YeC89XsRNO7V+n/jTP2BFMaONCwgFaHCMxE0Rt8Frc/56vKvRO
EL1BV+3FrK+58dG5iYMNlkiCLyOnAKDOB7spqxv++BSo6d/f13oeUJsEalF60gx4
9ISspvG2FhE9VA++XFbZlcfUTtnNk6PqkxFVmLxPHyTxGO893bG+6jYCvGnx6A+y
jqknIdKogKy2oXX5WHERPaTjErKD4r6bD2LFb8mYezIlktFYQDAyIs/EwbMKq68a
KrFz/J6KoJyLY58GW0fQJzZoq5wmNQtfXQxKtad/BZQaRvvMT/2TGFaGnbM0d6mP
zHyz/7+/6Buj6g9aTTP4QTwH3Qaqm5cwOZn5osPINd5oXzU9YSByLSAGYdk5MWxP
WI2laXKsGfjYyv8zT5S+ggeGGZDIMKC66jCVitMI/6CbtN+IL5OeV9v4s0SjJ0No
HBb6Od1gU+1DYNVgw2sz5vDhMC3xXXrCC6/oltghT7dBmof170d8M+R+MVt5tsuE
sG9V6kY3uksZGPYxWFfEMMjrpo4IiJPj2vvhDOVKmj6VPmPN1d2IUP4dO94JQSU0
kQD8c89fX0POYPBMWye7CqA/vt78ks9VCIct9ycIOpvWaMKHIM/zRT5/HkSDIO8a
xSBfTsh4xdA1hEaBtDVck9yOAHPO1Ffvx1RceflZhbLIec5Y8J5lvskV4bVla6Xv
pYbiOOqR2NYKPBwvoNBT0ddrjeB+QE55piGQyCAbbv98HhuU+7jQZVSCPcTR/jfa
ZOnSNGfUgFEwV027ayjbAgh63Dv4UjdNQy+V/hw9C8lhNCOXjhTVzHZAZocg4Ks8
BYKcSQ55Yev7nzwsQyR6MmsEA8IFBQzQHsAtCGTX3228dYM+vqr0KLt9VFwxRoA4
mkw+BOJKs+8N/NQVp52Op3MzbAF+oeb8zwq/ft61N3xqJ7BxfVrbVdedlhmDyY3s
vv9IU2mCp4YtOc4wjVpM07NdbkRF7i1qxHNxyv1rUxlMW2n6NMHsNF4omqBGRHUL
iicqj0XQgSZSbn1wnU/I36khFofeMP3UdsCPSSlkepxnCaL89ZDrs8uRGA/kn11r
ae99xTEDgb2Vi/4GCvRCy1o+1Ew084qC9yv8Fyh2zZDhRHyJsit4XheSQf7yiUxR
KbycxsLPQBPBrTdkRdCuON7PEbeEdAFb6HQ9nQE61JX2OnOwAiAboja8lkVy71mv
npGNh6Pyfj59scZkpubWW6o0DKztqHrY4yxh7/M0kYsQic9Ro40SDG2vwjPVo4U8
cMZuTnbphEXkhWezY/TyrdErXG6dGV/p9WPSHseY9ageFrvSHP/mPhDrwMXPMaXr
c1XaNgur+C1pgdFaRfqbJc9IYp69UOumtZkqB4Suy7i9byXbbVC0/WLUxCxITn3g
DbqdskcLBTXRPLZHAgaUl35ffz6BCEGiDvBo5v73fMAxdXPUIMqV2eHRgj2QgViW
RjI2Tx5ivZK73Rh2HxzGPekZlM/q84NXt4QOskTLA+KC5Ii+IGBLVxYslFF1qx7P
+jY0pBqZfQhZrehwk0rGZPkgPmPhyCFU8wEQbl4hc0cxWJqurX5tqFDx1PO52MU2
xUg8cberPKkQLbYCUg5OWipCA6lMghThwgekDcUFyX7/brP0U4k+7tZiwAQQvECJ
6yV8fMoZlv4YPtXWhwAFargZJBcp7NTCzO+FzgBhi0CFJeIdJu8btjJAFPh7/FAh
t64jTEr8CAmPe9fx6JYUzo+Z7N4G6Vg6F6fMvX/GTSD+NoMYImdLRhsZaq4Mv/B+
x8hZ+hFPEiEjxGkfe6RNwuoxSZpFZ9K4nV6p/Lf6XWmzuU+QLQYnu6CU1NlUI9TK
kZCOcEAUDx9ewGM10kvFZyp94JaMo12BvmhSLfoz0gDP/SpTHZa+OS30PW68RSNT
RbdqRqOpAlM/emoiX51nZdN9GwFQ5SlhTsp+rT+4yiD+3rtoVP4InmP3dW3Npezd
3vE6aZ2/dybW4kEzGsDr1Fhy7VrdSMF+7jKWc1xv3a+JLZDMeu+oEvJn6+vXRpyX
7oKmuU1P+lJhWoNI+MoyfFnkRigTR4SBasCJftfj0ioPVLdBB4pFRO4xyGJHVaLX
Du86YCyVxeWEjlO4jqzzyhEmlLzHl7A1bvlTru8+TyDdrl2nW8lDiMmI6KzeXluy
fdQl89h3SSK+PUyGca/99jQ1i8VxYB8G9zmJcnONHql00H3sdU7nEAVJiORmZLEH
o2Z4HYbDqrMR57nZ3W9e6JShvwIhQ8bSPvk/aHWd2HopNbafu/UkG2lZkyBhOb+X
nTcVpwezwNV/UMttyj+uGshcq2cMScFyhx6Nps3U7oZRmW5/JBwoe5XKPSypz/zK
PXn2qhJd9Un2htQdyhY0Tyab9EduokUqAzt+/gjYCiDXWorSoWS66eE5Dsta7Ki6
4yI/k2xOSWi2eg/wY7ayf2SyGrz/KdESvogsqupdDggs0v3lw79lxt2dQDDzgFdN
5bD7KgAAOH7parlQMnrww38ofl4ObwSt5bgq3Gy2wPK/SIPKCQOwmdGBp44yg73j
ybky4WwpN4rX91UAHaCqZEW8IjrMdJ06R1u2R4RGfuPFj3aNBv5XFX4tjLMz7UvB
24Vj6fQ7C6bziPY/htFngMprqIQW2QjDk0Iteb3uizv0KLHN1Zp7FHAOHq1KRJRR
0B6a6Luvrh9tfC+mDkidQqoczNpq5tDm2tetNzvNkD0WKPDnWl8JmnFQhPpJ+CwC
2jemyp9trysaUut0D5ICrAE+yo4rZw2XE5hg3RYMTkVPkYBIvOLRqO5FtxDv418Q
0SJqNtAHX6fqm1rp5uKkej3PlR8fanNzzNdVq7GOu24tZq5jZ4R9CjmCrCqQcd3G
C3B2Gz0VbfiKFVWUmFslrXXIRKy30JwCglb/lWxt9vyUb3JyeKIZwyxkq2IuOyJg
/UCmPQS2qvWSm2cvYlIJ4gWFxTQlhQRW2e1abNTfTnSs7F2BGcscktrVmKdE5fYL
ApXTPglgGsQ+AvA35i08kflifpxsZT9GYtPDj7hwlzOkzLL7nNfuhnbXPrpQ74VZ
rZZhHxNjxhncI+LCr/pKts83iT2LTLPP+FurVWjJ1oEgrjZ8O4IQVy6wirJpxp2l
cdBqfHM35KXb9SZWf+zSjgOAIBAMS1qJghE6DOYFyfl0RssQm+LvB7L3jzh/hERd
AQMNR7+sISXIgzqaSJkeKFpgaCm5oGOrLSQADKdVrD9fp+DH6JnVwSiUrDZGHjgJ
C4+m3ZotMCbD4hwX1snGic9+/t/iv/Tf6LAfng9haQG+zktJRoNHxvecQlh1k7eR
PiXxg61PoaUfENdYizSyfrfoPRUj5lwl+FoovKHcL4pbroFQLI8uSRg84dfAZy15
zFAQ1MesLeUJ87dNT62ZC955ydLB24FM5xHiok/M8d25Pl4xIFEcaiIGDBfZmBMv
mBZGPAGg6vcQPFsGVK82h7dKOyrhYlCIEVAGW+wf8QZga8AfqyPNXhgrC5KvNVgD
KfXt040PP3Hh5yJq7fjw+vGS5SNw+XjhrPF3GLv0GjHH0ARruxfJezUxsM7mkibt
/zh1gCPkJZ4ehi+Z6h5OybekjFRMr4TVvs2rRU8uEzPCV1l8q1HAC5G2Wj87JlB4
lb8pDyxoqfFgBx5fed8q3p6W9ih2wUx8IQS6NS8RdklDgqBTgWSw1unIcncUlto0
2rlbb5PRFjZtbJ8ewrHRHKjkyIBCFk2Je901G3zgoT9i5hsM599VbwedEfrSrg7W
jvL/qpGmus9eAToYc6n6haqGvPzp+3BsAgc4C5nWWfemsZ7FIph65ckiVNaCSFS+
NU+AyAUBEcs8euLFU2es6INGqJFlxpRc0TmGPTgByIAs6+qsQnMDSQ2QER26/Bnp
q6AJ83FqefJglAZVQPkLxbRKPtnq7hcYHmW1wE5WrejC/jVRhSBBJXqRQhRUGnkj
5QXmAdSule6H4IQbHvvLXFKVk16UN0R/rKGS0Hqy1lTCxDxrrRR7AHlviEVRjFuh
3ePSEJC8hr9yMKmNxt4BgxKeBwUGvW1VmNbQMxN/Yr3Ru4AEZJYUrwrHIalskThd
GpZbLBgMUOYODBfjVBV+tWxeNd4LU4LieDwfgg/WF6GE+XYmY9Ec6caaomgkL2fT
VER53eoZ6+jlImzAgH+8be5OgZBYxhYNOBJhC6KsrgZhJnAKKOLcDQGVn5ROtsfh
jy6hOwKtF8eaO/OawgKKNeUqtTuMYrQnJWmTfdPv6+MtLTLw88AKdqextLlkerJN
GKB+Nfiidw3t8zT0Ncqqp/ehhoT2QdOY4uQdFTgn2G1Kx4nD7CvRxkiN0yKYgfYM
oX9DG0prjNNGK45Y59Bhq70SKIMveag4w21s65Gp77uoVF7n3CSMQ9Afr+Qj6iyD
oSiEi9lDLGD+Tja4+v0QbTlNgRsrGFK8/fKD/48r6pyQv9t0V+gbBiT9YVM6eCCI
caB7xQ4Sx4vBm0HsSB6RX1HkALeZVT+RHWO2w5AycPbb01pWWIepj8HdiWe5G95O
56l/Bnqs3/hKGa+aIINEe5hmvp4rWMaFfzXXnVP0qS59OJO6uZ1PDMIBSY2bcaQZ
uy4r4Xdra1Nqh8QwgqxuuwGK+OScvHZ1iTZohSU34NvC5YCourN3VpSWOVoq8KZ9
utptltbXLXhUkIvLHKhpSwvAcSjuT9sacn9ihku74KiWBl97pXF9gguhQ+xBuemo
ky2i+WSmLOqzmi69kmhzX6EAmnX5XufEP+kWBmTAK1MXdbSAfN1zgFzZe+ncVqpi
unIBRvmkegyxyOCYWNVLI6DoiIc/wlJB/dsgLnu8pJl+Ff9Serl6cBw+ppBisLgS
L8YJA5YYp260hqiQaRLzqbfSFSmmWvGE8lplkSbj2OVy39uif2sTQUWXo/cBpF3n
qliTrh/qMEk6mma9DggRPRDM84IZRdQ1/QsPhWPLc4nt8bOq2X9F/yfwV0fAFTc9
+/7uPIvMnlciWCMF3huTVcAkuuFhHtWIZmj/TjBuQ1VCuHzcUA+xybDSYnrt3fbT
7Vw/AJnjFXxl6oZ6PqjSASNpzAVVQzZ1pJ/9NT+rtglTGvFFP12wO4sqffy6bKmO
MffUf4+RXDqDrhom8exc6tx+mNxXVgJE7LAqDNUrz2FNuDitxJs6nhHoDVtbnC3y
Vuj43bgVq+BmwixbMT+04KZcor/PNRifGMnvMbdkXRlz176pcNsXR+R1W+U9udID
giH4UGdcUbmC90cJ+MQGDrW/kaLd29gPwx5F7zHNFutFBezu1YL9cg7KoIV4JwSP
rV7+zPBmUsh3CLk39BHTMug7qumGL54S/IczbGHp/Ds3CcvbELzjHszv4KaO7qNS
8VLhUtCq9tad5MD6GHpMiRHEMwmPiBqLtscozlQSMzeKQJPKHcAk1o0LzJLoAn/T
gS8YmAKOosjGZi6yj47GIRZbjOrtsnOWr+pR7d0bE1bE6P39EsdptKpRg29C4bEA
F5d362NuFXXvFJ6NURdL5RVXpKvA7vfiZvnxDn5lPcDFA7yB0PqB9dfDpWONrSpl
irNeJ2tdstyGgrh6QM7+KGs0C6TXk4T02TO3jM5gTvRJKPVp7Y+4Nz6Tk4bYjBYc
TsUitq5n5gQbKjSP/vmqoI5kz0DlLzG1Yi0zlH9WpCe5l4BuYXG+Ke6W0XfDtbIr
kXc8dqArnoP0FGhtW77MW3iYu9mCqbTXXWZrGbFNA60TrkygK67BRUCtg4+8NT1X
nD3OCiN0FeygBONGcgCupWzR/GjZ5qP7UzffqjQPCWnFMeIYrPmU6R/bNfzYBqCW
QRUgpCduRHFZzhZlLpSt5cOnD8QrsvsSSInd+SUJn3iiu0zBG+kcEGWTFjO97mVE
QBchEaYDm7vxGiNs+aFZMzSJw+vLObXvEuIS1Dj96uYuWTY7HfVWS3NVIetaPfR6
Wi5VgMxWH+CM2NOLXu576UZOJEgEGdDDOMrOfIYlV+ysj1MiyCEr80qHriEg3i/e
cVCqxTocJ1euBEfTn4LrE4mRN9Mqw8VfdEIvaAjnOoE51MyX0fGPwCIqnQNluheh
sM385e4aWQ0bCiQG5nyAXSOy/CxNgMjPyJhXz+jKwa5sce7eVK2PBgQtsSPz3jqO
NxY8SzsRjHFytEAkY8J9w3sLnMU3XMk/FxItyDY1mE/mEyI9eTVbna9bD5Sp6Q1o
Amrec2hy5c61F3q2yN8uKUUZh3+swc9tuxr88VD8rW2s5ui/RNih+DiWKQ9Lk9hG
LwnClcUPygbHnqjm+4/NpSxaSInRg5tR/F0vTjBfFzMbBYzkmuoNmcGfPSe+Yx5A
kh7UNCEJeWgM6CzDNfmIVo2laPrh68BC6vCZ1xSWzI7gpwQNIgHwfCb1yaY7tmgE
zgdZk5Vl/WRP4O6gztx4PQ6fah1daVuabIkGBXh6zXQibMj8kV3CTnE0g0FIyrzW
N+bL2FLzDD8j55B4xX5Yt7NbD4JZdjvRFD2QScR6akoiy1k+KwUq4EqSPXY7X/ba
YLYoC6fdmfymFwkbJEmXYfeBRDVARtjOOTmOKIb8u3tNFNPdlSKVgRN0K8Ztw59b
itJ5wze4wBFkl/+MHd2kTdqKVd3oy1qXfrB01QLn5TczZOdf7yuzyF2tnrADeKHC
nOBRyEBPeMK7pN9oxrzQjoqvq/epsWM3uMD/DzrpAvogr6KZ+Aoy18+dxP3S1ABL
tJhhSvOjOOGfS24OuPBQCobnracYelKosdzeLaztwtjYzosaWPPh+gYsz2M/yfDx
ASbnO+8VkfAKN7TAcywIDtmZsZ/5HEveXjyWFPGeAh2B12E5vXKur7gyiYPSckxk
sJHUn/ELHhQ8WJPTkGvsawThWfZozyNkvuGodG6G0Wb3EWfs+EYPvLWUlQz3q93B
3QebQz7IXIVHmmb+SyN2igTIheTWLLgN1hPyryG7tU+NNBqf7OhT2/TuUvvKoiIT
RsG3mvqDuVPFu6iVBwCw3gwORfyHUXsimhA0717mPS0dPuAo/71S2iCpE/y99VW6
J1hOqdnNKLxpu8AwyGBB4d7U0TqkHRO9m6K7PVCaUPlFVGIYGFiARVH7XYdrQDV+
MG4ESLuY5ilomP4N2qA52cOg+InvuVnwXD24yB0m3XEU8r7paxtlxJJ46Kwx59Rq
SKjSZIIdhixjWnVE59Skuhz/wTPvmZCQweQT8kRUipewMkosvGRIu7ym5dtDCikO
fQ3cXB+59XRGkHsbI9sNn8+ndUFca6HWTsKMrQSwPt8a2NqkNJkxO9Bb4GEJWN+M
ZgCIMFDt1YEeN3THyJz2KnD+uPfjlC+nBf5K+vN54j9ShSTAnUYDl25OaGgG0QNk
9mrPfWTiurWHRAFKDZZL//M00iiqIaqI/w8y2RMXEEozY0q9U/xllB1AcBDT7QW+
iRuxqHmbLNyhyL8IvnRThSQqj9PnUk7MDHW+Nbqvvo/nCqeY6ZItPFrJFIiiEwIy
wd9h0WcWwK8BfQ+vNEWKLg/BJxJXejHbGT+jgpx9/VQhOJKvMFaiwVZDaGEDtf0U
xds6D1NIwNZK+3JP0gfWecc15BkwtccsYFWOFVgtTUoTxSMQ1hcmapgds5ZuqMe7
DvmlRTsuD3CPW/y4vtVFM6KdRm9BGrMJdhNLlSiau4p08MwTDl/Jugpk/lDEwXvJ
oOzMuC1gftF/p9VPiBXGQUVdCdNWe7qFH6rZvQA75uWAeaQI8/Olf9uf82svR61X
BCwT3o3JthSYHlucWsN40y7D/3IbLhnR+5Ovr8Fsk74c0mENGxdNpG0eBgtFg/XR
GkBkKyupMd655toIfjbNFp16YX81iZ5cwlwhDB+OhfC8MPDxUCO+hKtzVeizN9bk
NJB07PhUeUIUotftxJ8umXJPyDWB38KSUtxXEZDnec6S/ronK3XADKkVcqjGPMUW
le6xGRGsibjWkym3ygF6mFAygtP0ZiZpKEP76iMezUo8iB4wiVu1xLMzSWMw855O
UtmxC2f0au2/qflKOCwpWJVu/8E0sCQ4XGAhUv+Nmt+9JA9qcde4R0u0zdQFNyAW
Vk3GDihEyu2HdKu4tFOIDWa5oLmqvtrU8/hTm2fxqCKf5jfYkecQVK7ReGlxsDxD
KGFF1SPIucEVznW4lk/9asj72StExioeyYkwO3WOc9VMVEmgsdZqt/BTzkXdQXKH
3lSoEjvyw7GJF2wJgqSuPnYgIMam3oBLEcoL1CmMLZct5EW/1yvsJBqw5+EjJb1X
oDvit/BEr+AbAzCyceDkM3xBWQUMtadBWS/Y0CUV1ha1mMlevX1BQmQgBAX2Wers
avt3OF1qsK2Tg0as9XBpLgmcsuB/YbchePgWaYhNQjEJSlKTVXV73jkdg16E4Vxn
BkNXplrBbmUI5nPxhnmm8NB86v7eLgUYQks8mZRsfO8SBaBKdlBEknZngC83INkd
0rBrDqXurJ7u7yvLksK5PjgM7fiarB1Y82B29exH+xnzNTE6bH//IS1vwYJARJsL
X9xDK7X+f8+I/ZyiKZtfVPUyPQsL/Rwk4yVVC2L1Ppcz0Iww1Crymx8LxbEwcf0I
i7D/vRDw3qbg3hSPFby3NQrfj8IBiSLf0pFMg2xMb6nV/OHFxCmiRDBKMkjjk5Ob
g08Y1uVwWogBQkD/5gWJvUGFek+N6lzVvajZmPCu5Ry3YE2izi9a9IO3firy5GVE
nC9r+WSEfk8W43TPSePhSjhrtD1ZdkYCtTnMV12GuqJOLYE4b3nHi5dyP5X5vGzj
oeE31iWFCVRRsHunO5crGKyizRoZN4rQuhLTcMqPUVwqMt33LIQPWBsQf3rYK9pz
LqFsjRS99WP+KyXX2QnU4pgVmIdQ0B9iDw6cxq5FLnM/UZRzAIzB44Pnv56IL5i7
+DtF0nHOGAE6eqcEhO3c0ajCLtFivrA5Jon9yNgMpFeqRvIwOzwq7URfSJ9C85l8
LK0I58VA89oaVM/MtCR4r0VHtO8KJeTyy3xnlBb1nw24zkwctazUD8KuUYINPbIq
HjCGMVamcH03/nL7bOYG53cRdilSrpmncwi7QJHjKt0rL7TEY7/iSEpp+6z63Yin
OickyVb8jxubo3CAUWYY57yUtha/LI32aJ9IbFcG4/ylU+z0JDXSPWWErZFt2rsL
BjamX+XEZsWIPE1YCHdaSU42Uiiwswcv3t4WfzhPIITmVyZtBxbgn4DLsTI9G39Y
PWAkXFE2No3rccOVnKjmV7N0xEE+ojeZ/zqzhYEJq1741UGhJKVVaeHUr5VVRYmg
tatKTa2sDqQa9UomlHJN+d+xz1XjO7q6Ec2sceEoXbXKRvUaD/aLFFYlWq8nZcaE
q8ptE3H8xSysqZi4XyIUCtUFga4cAMo5E31TEYWQKw2Ocq39lAGVRRcyxwHx9MJG
Rz8pJyQv7Ty/u5RdNooZhcYwHgxiwo6HFQqwSZhAnLOdGttjX3mBrv6C72Kid6PA
HMDUP3Kl3mYSgzyw2tV3k7oOM2wpsO/6UpR8TuFHHqTybvbiIa0AAytEJgNEPNly
2oSMzMESSnSTWrjMOTGdwiUaHwA2bHYlBKwtBU5CKudmDznyus2A4hCoGeYXcUPp
kJLSCo7PztajareRX0Dc7/1a4y6R55eGy3F0/+cp+PDst4SeH8B5tYjz61QD9wOm
yn7ujNQAVoQiy03uWk8DwQKfutK6e3H5WnXuwy7/lmJw4axa7CHsHE2f6HjGyVz3
ALxLrmx/8WXEnHavbRm8ajXdQXcQUQWkdiWt5LJpFHwKQqBSD6HMkcJ5qONBFp6Q
3WWDOTHt2XOy2wxOGAsfLZvMk3zlcsG6bVIDbH0Bxw8nRFP7/uqnUbVr+PF2gZxZ
eajDLZKbEcGy+BElhRi6DLz2GFXdjevtGY995jlxnzRfYTMSuI1UFJPxYdmjvEfR
SMxq7F3SPzoTMwI/337VoNTcskhuMEeyPtEEaILcbUI7L81rd+ePbZl8AJ2HKRU4
1errEyw8MW1qeFxn4DP7h3BV8DarZHVYyhfafb+NamlTfJLdcDFLTTIKyUAPSnKw
MiEVdOz73xa8mjH3O7LO6ZybckdDynp/n3ubmWnZ1cWVRfesXC1ZbEFa4I7aHVoH
HtogkbiRGKZDprlUcv8CmOaBY4fGgGcv1MGsrT583oES0IL3FtOQp2e2GqnHCPa0
QtPDf+LM4b1iAmQc5iEt4HnqpxG9pp8mgSrv/TTMvuQCJR0rk0/K3JuQbVqFaWUa
carVNecKRi7apAWXTPUcIA2Y3CBnUppnnzMEYWHGVVkJ/A5TMeLxmTNCOrvol7zI
AOIXSxK66BM6LR2G53MSmFgWxYZ0DlF3fMSmmMdQalwChxUmbBly5PQQqSczm9PJ
sV2A4eBNiTXitMUA9xurA6gRYbA4HPUekMpU1z1IOZe0ApjUzvTd5GqPbWLNBnVU
sdGJPVrd2pWMfSXI0+urX3HzA9UZTRR1FDBRvKc2cCVoZVDwBvFHlIa9GH91W+eW
wBQO75XMxon0MT1wBYDyTykr1/4eYJb2eUeUJnyZwd4NcdypdwsTzg24Jhxb1fH4
h8uLGJEE7yfJK/EmCVotX2PIWufbQIPSuY9CdnI6eHs3RBr48ZAgRtLWaf/cBajG
8H+5pcivmjpxQuRrglD+dik9P4QiDB4iMR13vM56XdwwwLF46LOvHejnrq/Nf60l
v9fl7TlAh/TcuYkxRKLq3Vyo1MGHfCCZwYeliEJ7gKiDNvSUALiRRr+h9c3w/G09
40VVE76PebFVClKbsJHKBJGOc1lxf6gy1yAChpJoL2mXlWoMrx+wc0k1ovcj9Aqn
hXVDYSojYoMYDFM9juZQvsDj76GhC8eSI69TRKz5I89Jjo3Mto1NJQWfR5fP232g
NpOigjNGzk+v/NhqKz8C2XCD9vJisdKSg8c90hxx8lEQJCrMX/YAF/qwK5ojyvJg
f4tdvfL5DoNtgQ7hexixZposD75+IY+oeMiCjG6KG9Szt5VKBRj9jyYllY81hSsH
8G8KruLJ4WxW6zUQWplfu7Tubi+efo+ixVyde6CfjfFvFc51MKGMRQzKHidQsT5A
4nHqC5x+3YEj0CXApM7vihn+8ZaLtRIEqxCFofPF/kYzXYXQ7Hs7Azyzgri3Rs1H
DTaTy/5Ef8ML/GHgWeMpLHVn2hbCuzMDqu6mZus3SvmozMP/JfjZnOaITyo0ihKv
pTmRfVOLtiuYqufgdIu9VwkKC2safIJ7tRUT5SQhueTB5z/mDTjFWYY7UvsV2IdI
QPzJPzMOtJvdcCyVbGsN5NEExKUP7Rt6v3cE/q06oIfNfy/pr8Zq/Afve+se/CxE
xT1NpiWoSYgStWsltEMN1+qpVCGE43SFMa2At+GJY2Xth9IBV40bi+WYqEdT3xM8
yzGoV+bM1uFO75hhm7TwY0MjhCrBoDKxtl9UdLe9+ES9VCSYIU/p/4vyLwKTnE/r
wXxVPUcFtr8T/gt7XqyUCCF4Py9hioszdnLCvCv7RyV0kYR3sRFtbz+IVvX3vqOh
aXL5qIiNomoZv9Rf1PM3OfNoO1M+ivRG0qixhzOS/v84r5sK4096RnqD3Ivc5Eb/
3mLEt2UN+RwRt+aJfNVY7vdvyBGG9VzNjebi2ZFsAoOXWT+rLRG0Q5Te03pD0hlG
4ADYFdJUfWpHLAjrCdMqh1kOS3fe8YGOxQjEWbc/WYkYeVWWnQkfCCiKyFuC+bsh
C37m8lhmSBrtPyyv3rsTOZurwl8Fe1gAt+SIwQnA5jfC7A3bpGK7nuV92wJOd3w2
/xGFsXivPxHJhAHHLUHNz57o/nyud92EflP7bDePZRjfrVR9gey1cptFA5W62BXU
W17WO7pGxCvIjeRu+0D11F8Gv9KXXrPdn0UPOUqDHvYjgvlmPf8AFTzpBttKrUoi
aV2srOsBgF/sEV9nmfaMkk6p1si3FmSabr2sAS2sL2Ldzx0kv/5UmPn7bSzZL82D
KfstwDE7EtO1rwCHLKgicWKJtquumyQTDuf30fMKvK+9HVc1GXhcaDqF9c+0a9Ao
pb4iv91j5Ivn9JVf+145Om7X9uVQpk2SwHY4wsfUReZa+7f06fYFFD8ycN0Kh+1u
vgXCfEdB2Kf81F8EWqWDwOGxpI5jztpLuDlYp1qAWO5YyExV8PhROMlBCvW2mYUF
+f1NyFks4gy4qpMzU2Ud2AafYj8/J3Bhg7+fJbIOVzXyZSyWktkWkSQxNr0bB6T8
EA7TNZuEWawW1vECDdP0tenRfhGG2cB0NMwFsJc+ndJ3L4augjqPtEVil+z/ZBy7
OMiIfgNBrkqFGoTITG2L5LvazI39UTSyOlGpXtlzlg/0cDaIqBFsiuP8vDNx1AbK
KNiVQHMZaJ8MEibnFq4+IgDUbHip8yOSxikheBHKSi2GAsAYVQjN2j2wb6uqMXTt
EV5/eZjhduBZ/QT41j0oSGSuomb3HHXoB7BYHpSc2YGqhMgkEusttFvTz3ybPzXX
rVe73RqfE/cdVwYevQdFDtpqFTT3j3hiHks8bB+1eu+OtB0WRU4ssafSGx5ylN2W
BixH1juDkpRrDEKxqVp9iPaobEkk9wSSOwsL0dYsjH46RoVwsfd1bGfiBf3Vh4Ds
nINljNYkieDltXGXh+a46Wbc7mtfEjyDxgHMl9HDaaGbv9vctE7mQceBoluVZhLH
GTBL/KtPyurGoL0AOnm7tZBtOpiQ3H/5LPutLwT/spNPHLdz5LYnGCm24bST3ITX
N3lNNY9pzsh9QyWIZKObXqPemkdyWpJEAR01ue75vTMRfDfRNzBrXPBIj6/E95il
lmicRDVjx55SIliP1zhg2HuurZ3Y0JMebWyUETvbiPpaMgzGgzKi7pT0N1EgLxXP
9cg4do84BLxwhTt5X09jkVhQuC9+ydlrwLrXZTId+7fqtI7mYDrsE5MqnaCrEXVA
UiW7QdJsnGRYbTQg0ElRB+XuVPENm1xFCEuL/DfkwL3qgGYKEn4ONaKcH07FZauw
DEQ0CsrkDasOccyV804x60HriIeC5N6EDUPnGQRErAn1WZk8WxLnFFRgI8eeI5A0
XVyx3ALcNEzlgQDw4n7qXwO76EI0jsaiBnFBbN9KKKTb2BXHEqMs2BuOSQwAEssp
dZjmQBxd7/zNN6R6FS35Jqwrfuc+WCptvcme1Ch1htpV37sWP++PY7MJGU436F4N
k9n/fUt9/jyqj3qJ3cDrQ4XQEZZe/wYVwaCj8cSnW+rLE6J+gbjtnoGiQVdgtZh7
A97J/iiGABosXMHPe4kcxBzvVIulb3bKmaoEM4tEw2hAQZuHv25yD1AAL9lLbnW9
x1xP0B/Pm8ZjlYIUQg6ILbIMJ/5u24a2eciXCoMUoKNfCDcpMSt078zpHXFfj1T8
vUfJs00BUYxgVDnVwA3Bs6z7WUd3AhXo+Ftp87JJKcwZ+qI5VBXFOMeaRrEtJqys
mTrMBRpnQ9rmKLOChQznEx/gta60dxjEia6kJSlEV/OBvu2t/MyH85JeBqDaMxkH
CG4358OBjs8jkWc9m6PCnyFGdZ7DngSHuJF17vNGlno0ewzbv+CJqZCFwTgwHDXI
QBSoPAJdeT0HDdVUbQjOflG0f2ScncM7TiufP9X5T66b7CQRamz44y7mtz4L9Gj6
YWYXqWUzn16PfDsA93hBPhTp6tkVzErsGCF1EMO6G7JuEIasrKTaRB8UWEQ8xNYA
qvYVKefuK6INCFARc26uG4PPkccfA7IVXf78lQloeibXT/RiViD2LkmduDcs5M7Z
nl4ppKHuaVTE7hvcFqe0ffS6q/XGOtX10pwYe4bKGLbDgGrGy8VVKKD/pj2ZkO7X
NBlNOtDn2wLIMw2GnQt/OdeMRQiudKI19dnzQWNfOjq1/47gS6BUWVuH7T2bvskQ
SCp22oKLMiv1Vo9HS4AyQwqG7BwxcGyUMbhxGQWRYe+vWgLpIjx5EeXg+OWdyR/N
PQQMD1MGD0ug3vOqlw8Uhw6W1uBfYEyJfFgCtBQoX2xFZWr/kNci3jxSCUKJmmvV
qsSycsKUK2SH5pF5IKJYFxzLW4cw4Wru3g/dmvqF+rSoxLGq6+uaGqGJehHGBpci
pnO94xYNFs2SBodG4C6X9TvNXBZ1juNp/eLMCkrV9WQrAJi+A6djsouWRcTbxkPe
AvHlyrOihndS6yquy9jbJuHutjpsyPPruFS+uEL2l5Auktm/Bf4w+qxtKfqzVE8S
jK/eiiIr9Eddqo3uqJ3fw0GYqOgqeFrGHAf1VT3CVyYqUbyetECozN4vq6Uw1zc5
D5Lp4IFGvMcvLshgzjGcFnjOm2tPMiRW2wfj/T3zBfTUtFUKIw6qR+WTJ6ARchQO
fzrDuKL4kvZe4VV0AjN6/uQFvmPJ8vCiLMGYBmucwtpEKQKICE6R5+kIFxelZDFj
n27nEYTvQxa3jtYNw7yvqVp4qcK+e/Pj3Ak8+rAMnwvWm5WVk/XPCJ0ZPQFIDwDk
nOoq/yCeR5DpbiRMwgQkkuZ3hiUmOSMZ1d41gZAfhvx5+lkR/lwxZuOSHPSGKOhE
FP4nSKB5LLUWXBihd964XxjrvCJ3k/aM03HFhvbF5+LZqUHczpC67qCfq7p4n3lH
W6dV40wq5wGzQhs5fIprjZHWtt2YL3OGJXVf+v/YqwJJAVzQox4I0czZB47XRiUU
2WE+NPsiUddy9ATyFcMQKx687YPdX/t4kYK7AeWbsEyYOqFE8L0TA0wypglKoZ5+
UM+kcvav7/xeDcXVpAEoNLyUNwrmwiLcyZWqNtXD9dW2fwDyupnLDGVSR2cjbRaZ
/a/kut2v0HYxY1YVOMKAiPRkDzucwQ6qAow8gNL/yd5knBlJWkPE+mA5QHJ4GjZL
V+TN/NXVqzMbn5Ihm30t3mtXbIRuTLlU3gGUilB8eW8t6rZRBzBMxMWOXwcbjs6y
RgL8G9oiGjWzX2rLduaDv1i79tmuvEwwiuyQVCOry4d1QOloxUSlH3s+kaLqquKn
y1BuFYoLUIrfjGFzwtaXULWFLIV4H2KYVxVcVr63AsbEP1SnlPpro+RRt02owyNx
vrSeEhPymH7muv+7IlC3/xnXYzNZQHUdzqkivSgr+k7mAS/KX5qk1TKb3++9qVgA
gHvrJNJyxDz9Epomeq9nhDZzxVDLQ0zFgbUibZH1IJCZXNcxaulnu42zVH9knC5l
RO64RdWbE2TBy4qGtr1x0zttrLCtY8GcXT8JTM4MV6Z+La666iJ+1dNKxLVRTzL2
B37gX5C9rm+8LlU/LY39sZpVFL/ut50aLqe7oeqUwoqebGg3Ds/fjqD5h9lQtj/o
HLZ2UiGnTNVwkpx/jfFLITKkL9FNCVnKOnDHQUfTvXiSWRKbTX6uM85dhKWgoMWo
jLAxdPgCJWMR7yFftgCDL8vxYXk3+PiG6FiMRvtlMS0ExtYqty0cAKRdyC7kJGjW
VOmANeQFVAQIarAsRe5RwvrLGEW2YGqdvPA6DwJ/VgDW/cc2cOOQI63hO0txTr+i
+ReDIEjxdymDkGE48O93J0b40Ng11MEbRj++vr/eNVccKhV95pX3xln3qPS01Uzq
PLA0BO9EROcFwM7ajoJic4dhAtCyfjNh0feCG+OqYjbkc48GkWCCgQmV0UDeqsuy
m4+rT3S4aPVgpQr7Za1AlzN07pFBwwrAtM/5UQHyrzRKiltzb5l0qVeKelsj7ooE
T8XnQS/xJN0WbJNhu2uEWk1duvhtWiylaGLV2upxflCc2Lgm6vIAlJXVXsUaBnTC
k0wT9E0H0XHWac6MP2Xp7e5QIHe2l8Fe8CiBoHFdIuOV4r+0Qa5nqgVxpBVr1H7w
brSjrSE3RZgtOhGqp4dY4aqekMp6fQ85vsdx2/MYS2J46z65NcEcf0xURYWQPN2Y
2OW94X4nLS+XYUpf3WMIii2ckr6KeXUodAPjycZyEOrG8EoYNfGU51c82/e2K0/Z
KiHD+1a5XIRB2JKMTpssxJUGOcvNxzFu/dBrv6IuxjPJoyuEpE6NaB4Oh/zk1UOB
T7B8YaLZuBSJ8PUiEvYP3/Z9BCfRSXIMmuNOlHcj5iY0raLbl1BOX7tkLQtSToAR
EYxWos2YHKmszTCu9UPqXTzHETeBKbEioiPDZIegc5B/lNWI1rJUQMoQrcshmxGf
U6Uf/9lR6eyLDYu6lWoJOihodJvFm1VpSCYGEs8OMhAFBlRpaqFRVtyAVR7zH5yk
i+i9mEq4XefhCnE1dBuWD/lbPCPGbQV3SugWpqYskwEjXXfYVoPWi44GIqU9agdi
zpu6BoL1lMZf3GVKJVY6yw+vbwmp9NbsKyqce72iM5DWVs0W3Uqj6GcZ2mSZ3uZw
npPS7hE2wmXQWzrXyQS319LVlk5L6jafXrQU91AEWX0ytfQg2NsyTJQvfhHWHsI8
hiDzdqtXcJVVrZuRzXxImv27cyuBuNhV4epWu+7bb3utVVQIK6Lyn0eonqHpndKf
V9uTQ34RxXJnmt9yJ9dSVp0FUjayhCHZQCg92O5fSg3yi+SfwAjhGIFMJpLaOtCa
S7RCKBbKgxDd91tyegUhFp0UHefzeULz+ayJptpBzvex76HqWhaB8gBtTXjClGvn
UAVX0nyl6pln/VpoXZIq1+gWPAGaPl3jyv/mjvMpF9u3uWYFFMP9T1erm/D+uIF1
0Yi5MnoeIEWww/jA6XOf+OsA2yZ+NM6ywq57dKl4g0epkRz2ah/WV2nzce8x2vEm
xVuC4mo7EeS5y0v2JZ/sDiuPNGiXPzLF0u/LsypBNAHCfYO7CiuXl+X24RxKpGca
2FssDf+a56RDCPGGF7DbbuJWctiMLRZ5UqXyKFuuz/fb0KvYbyMXz3npautrqVKs
QA6gNme0LFkvsj7U8cw5xgM6fcnkwVjRxpUicVrxVAgk22v85ArEbaBI6VUUcBkF
xVBrQ5VYrFVGmxl2qb/xZwP2cXwn42DI1lSIgjCAbMj0qXnzeTAAjSqluQfoJuax
5ToZhogzGUKsFtnHI9GKJqrPcRjcY8puVmpgbRQNRnS5qUqUvYhobi63gShs5cZZ
yRbJAkH0Oaka2OH29+4IpvdKgCRtogTEUEujuojpHkhHwe88vW9/ghwMTGAKJamI
L8SDsNrJPTgP0YV4UUdkmHXpK7u6Bbxxrij99YVJFsWmXWCE5PSWokqJf4iaZNgY
IaCRSreVjT0Zd1Cykt1qrQrkwxbzNnPRBMM8KVT4AboONme6HwNWQDm7c6HIgfOV
U1BGTkpTzr/RHNpdhAjEBiM2U1rb2JpI+VBONkx8bLzVbTtsx/y9UU9Shq+o+EMV
DNCbmd9YtEShsIF4j2daXGZg1//l7ArBD3UnFQHrH19AULCXyFTdcAVgBSxmLm5Y
b/Qj7JaE51MSLxxjatiQBxiPAGL8VtcMOX6Ou0cnUvD7SXeJ+TbKNVb5aqjEuTcB
Ub0IpXGgzyzAp5Qp3pLBbAvHkW/eUfhTUebc22Xklzs1PRHJJ0IScFcsqBnsViZw
AZrczPX4y6WtRoPcjIkQbnz1/sWkFPBVqjtz8aq9bw4Ync62OPnbmuajBjl+YQs5
ztD9+dHbJEQsSsMppROixcM0aejSh2qejXux45n/ozylWTkd8ym7W2Bai9Kcg5Xs
uNd8AClsGJskXVT8CTQLdoUXWmdoD3S3OuWnvBFWRpycG61qhpemg6x87w5jsjVa
qn1H97LcaztEJ3cxmi8ez6wxMpxMO4CinnsUF3ZyNk52HEzKnuFD7ovtomlTGe/D
BzrpxPE5+7AvWF0giDnVWjU52WOAEZqG5hYZtNE9L6u9R41mXIrVkSwKVLSov0y6
LxZF6wLFaOra3NR1IT1MvO7RQGz5NSc1DmJ/O+I6keR/SECqvt5mlgMcFRd2n7pX
Qy00uaQlE+4Bi1Z9VXBT0wTAvSPN55er2hyWjIv17jBlfq8duoPMSLPQufpZ5XUZ
d3l2oksDWRoKLnEMxzLhiMmRZcB1OHvBfVmu0h0cJbN5dULi08h1CeXBLSx+X+uD
KsKwLRqDNa0ybAnAVM5dNEY77PMb3wQCqzsxTNcqZTp36G0paa7teM3vI0XgZefY
9ZT9YPKMKyF2T+PzrpDYkrusa2d9DIUleJzQdoelzOSLDpvJA5NqXj1WR09jMtLD
cuQeUAw+SiX6YGd9Pa1oaOc4XDfn1SVx8xVn8H5/J68XiPOc0YWz7nDjBlkgXwvp
r/yLGL1+KiNvwnvTyCf4yLplaN01v6PYE4gsFxhutIieT572TSPYFr3OJj6eFXCW
kNlBluvLd2kEuuDGiFu94G/EyKi56HxaGTRVfYUP9MgXVOxJAkt0xlMPrkb+L5iU
sEFV8TbZChPFOTm+NENG5MTvz2tP6kek8M3Vy/E12S11IdKV2rSqfXv1wQweubrN
1VXDA7kyGrj0HPyX6F8IlGPo5X8glvu1XrIXuQUlNcYwcHkhNnUVOErHcACF+RWK
jaaR3JXOrWOs70ZjUf8phszc6s6v/4nRQlCWnorlo94V1D5loiHqLaDqRr7yxR5U
JZV9fHPKoL/07AfDAmZ8ZsG3qSbQ0BRGHz2im1LahiJdoOIxWNAeH2UoZBjLgdn6
iNHk6a2+JHER6C7tNz9vFyuOpI6wUHxneZbXHyjCOYO9opH3lHIhH7f2ZuxJHd+R
Lt0l4zZc8fELemxmErbnoBb/jS5+VfnQOq6t5oCvEt8TfPjx3FcufDRMgTFrl9/m
ewuE1dBToTToEHzB6f88k3S9sBjuYYmCrLHkHabH9CduP9nP3KQ9IbbUqpCE9XYq
sh0Q2g+dqCi/Vyf53D4bU0leuAtX9bGZKP/BdvkulPleVPjoGgq3+u0OyzqZG4Vz
SFX4eumrU7UMcDQPXsyWxEoiqTiVrgwEQvvMArG8CxbLPHSjJcgCqrVgZ9mC0FWm
QO3+zYs6CrgAVw72yn8gjxy5RNmtsn44UBp7VKhV05dsTsDyAYaKFkMj4VtEzmzm
56GtKVUPC0fkPXYwqAQ+6CvWOvY83jS1uanPqBJcoxkJnC5S9svGYv21zE7qrk0r
QGj1OtE3LTj+4PCKL2YA4MlkQExuigNXNRLnP1IIEsCcKZu+ALFgCh/BkL+bA2rQ
2vkAHPl+DdnmyawrPngcYC/xkCvqonhK1eryq0KNzVYR3B6z6nUO3qMoq7TShQUE
t45cNeKDD6Wl0JwoPckyLafBvyq3okxqwdK+5ibaqVJUc4cASlyaOAOvz82FjSp0
QgOsnBeaXgAqossh4Pef0NNH4qj1PK+4uzrrCPWcS66/0oc0k+oWob+TRTiDUw44
o1rmxgu0zCyFOukzZ4SSW0F5TKGYbAXyx7l/kTs0BjtUx/LtbQpNFWAxs6geinmT
sp87aBD9ykJMbzpHmeBnZ8OiN14Y7iOgNlf7dg6hL8e3ez792cdMS15O1m6WcGRB
sgUuGFAdBwsl33T8xCr/dLPmvVRS5mAXXHmD+GbG141parMuP/Fj1hVj534YfPJe
Zev6ahadK//5dwGq2pURzlgqvZtIERM/yV3RJCuBeplbENhM6unfDCooygYC7L8q
1wdCuLG2snLCjXV1Sv/IWrNJ8j1Bm4M4m6IMRFjbQZSUkWhVWW1TPP394kBL+XTi
4+28w9rsK2rLoaY2eaxAb3PtBOL71HX/8HMCkGF8tJls2nQEbn1AGnGcQLINUoWJ
Zlohm1zK2SmUAQUMnYjYgvodJA7v9X/DIhhr8OLgSLVXXgiGMYfiKeI7R2Za6hLC
NyQ2G9vCXy3OY8ZJ8fgv+ZMALNZgLu8p+g0xAksHZ+Amx3vmwl8A6z/Hadoj6O/0
ewjoUJ22oWIfJH6TDBsn763kgJQwjp45k0wd+XU0eHphSJkaXb+Ae3lRAta4jVEd
1ZwbH1BhOxjP5k6ojiJydRT9fT3/3ZHjry+44FpIcdiLLign8ABWs8FHO2bqARds
d5hOCMHMGll3LwRvtlfIjHVmqzcAYn8IyDGWWfXbOgIrs4E2VCz24Oxyh0B/HG5R
RsUmWula5MWCf6JR7tviId7JaJAw5/jV+4mxxtYoCo/XPly+YqmTDfaaeOSVcZjj
4wjZ4HP6IfxvHmXHts/5jsb1Jx5h0UxW7TRcxLNn1ry7sSAN0RvI4JIKz7+Q/gta
KwlmemI6uwn6MmyWr/t9pFWZAJCfcPkZ8AZMHH4NCF3FGRkKD4XWJYfP19AzJhR5
Fjh7dCZVFlhch80i0CkJSxYKY7fkgOdlBUYsoUbW6LlVazJ+P46uL3L688BwzjgJ
iSzuw7annOjzDTj/zFxRy2eeiqxdqafQE6BBr2V9PtUiRIzlpaZ2bqkkv6dPOnet
jbeZqtMRtHqJoI5W1OFRbPCAyCXF7TrHhLNVIDxy+muAVX8Em+uPDI0NZM3amOs+
SLLjR9QEIzXJDlrV6RnTDXd+18crCU/vNJm02rnFXStrwYWwWnZylOpN2mm49aRD
bLesk8PrZKOq0PjhHnVsT0FsOcHLg5V8ialhGJwflDIWWLWGIB3CWYSKWDgedVwx
oNo7Jmit3UhIwtRwI9+McO+j8Zp4cyL0/x0cn11VR6kkrXZvUb3KlvtNN6r14B33
PPK/OWtB9OHIRiHqlaKAc1+YCfMFdsAk3qDw/9u5listng9hro5O/6I22XC+Zn2v
SElnTyEXa82uaq4ZAtD/GV5LAYj98TQe55KH8qwdblTkoKLxxCSN9UaZZ/IUWtY9
36uxFe8v8un0cY1Btqc4LNtqKyxvSmVCOXxivmNGJA5P4j6Ue+K91ar7lak3vTfR
0GPJrxBgG6F5wxPnf6o59qymKLSIAUufB/8UWX+scqPFuHqy4QrTFtuu4UbwtGaq
QS9F09G6dZq51Py06IZUlzJZ5sR/M56frOfP6ni03Xf8lWFhMFPMdBfm3/DvbuWI
cmUakWENN1NsviWZqGEUexsxCB0LUmUZ+d73qUgsf3PMtCwb7tL5uuv825z9UP7Y
AYbF7jh7iRJzgk4FLr4j4BlUivAyChCdNqhA1DaMNFj2PHoaXICjURCZzEgaSNsk
0YURXBwuB2kzmXV1glMsK3LgBDTW5zcaMPhzu7vbQKqYT36zYFIro55CBaU17WVJ
hY5t1atHMs5PyYrnesCE9N1sy4yCasLSwyFppaw7P+2856A66amA5gVPz6LRg17k
ws/9PNZeKFAQmUznqODC1/1BsB0KkWRrIHasGKzmRJ2kghAbaKsZoHqZ7RKLP7l3
WZ5s8pFQWAYSqxKbnZKXNOFSKioQjTEEObCnM7f7D1ms8fr6lgmrNmXLgHS6dohT
VDzvuIvJPKRDtuhwItISOgSECCHFFRdlFWbrPojqEp4351SdV0JmxV9Wu/gRmeE3
qczcx/styxHoVtbrOoaoAtCoDKCsIoAgwPpNdkqniskg7fv3GPbIAdA2czqRxJuW
PqBMWYZujFnPYi3y31wp8KIRg7/hkITcrkq5V2fApT8YMJlJ4NU8Z78MHMmeUGqF
KN4WCP0XejKLJE7200pG18Vj3BZ3sJ3yBigYcvFe5SgvKNReP0iTmrwoRiVhV5wa
ISF/6bK7TLM8EZ/ztwOL3mMMeJ//XzL2wW1IDYA3cjv0fAYW+CmvGFuFyrF+rYRR
/27h+Q/RuyQz8X+LnjHH2MWtAY1p9g77QxDCD3EZQXCKQolJTXKqO++UsS7nDA+a
iTE90Ta6qU20x1qu4o17+Au68GFxmvIHL+5wd43msrn/WYn2qM/6op3fKjPcE85D
Vv41STz7Atj0BpXsRPyK3mRgi2HywTTtVgwbsPxzkukKrOAFUb/YMbnpUxiB1Uuc
LUmHUwfrcEYKLbXz55qEEh7guGVt2daZ4C0cfE8iUkvPN7sPGpgw62RSk6h162cH
AucQ0KW/rN7xMHR4coJiO6w+rOlNo4X0lIpvfjNHKdqCtZjltv/Ym5TmzF7jqE7q
tN290kaG7kAAODD+QZtan/6tiKqPmne+CEk5W1tA4TzcSFMmh7L2K2EFiRgxKwG3
QiJu1pgCsFyJ1fGFkaFtRFekbuTqDWl9O0ohuuwI81K3CiQuJqbnwbkfheGXm3L7
UOyob1L85mmmBa89y1rxnp+WHi1AE7ppByvaODROGceBS5IuLxEeiduknQjbrFdn
thrliZNTSQTo9u6WolcJSfNQmK+nOzqwuNW6J0eg9aFa9WKiH/qe8aMd9oBSBOGO
RFJKKNUphBs6gx+EkYvlvSVAMNe+bjVPylC6SCNVeBF9JNwfyeUWmKmPc73A6bwq
81DtH1huT6NJA7lSO93lcWgWb7zJTJZp4/OJJ3BtrNYbX00nvrzOjSYrKEOER1UW
LiWw2tWPxZft0CyBxQl7//8SkQHLRdmJ52wdBvPY+Yp6dPO52+l6wv6l4hEuV1sv
D41jgdSuNn8w7AIs1YPnIj/74vaJHBmV+ELGCwR9vxD5trWTyUQMlXIMII811C5o
1svE5yn3qNlegTrwK/yLoRPiFWfEQQGVQi1NmnyPVGrwGuZ5ZklqatNm8r4pYr8q
3AegOMRRYaEZkp9ifeBwbjWVAnAxFP7C3h0BukFErHj6A/xP0n1KsAUtGTVsM5BB
RIQlngOabtK01wC70DYJ9pWfkSxUaICN/W/LUP1sLt5x2pdRPfmV1xzZTNDRXnSI
rdRDE2Pi9sQw0YcOxJPZFI/Q/+l5SkJccRdGcX9/0to69jey70nr6eJaqY+WJLhs
UGO0KYFR0zidOCvPmMOJSpn3CE+YRKt+w5Tudzq3Gfh6EEDlnYx+hU7x0aQZaqBg
aGcZ9wlE1ycvpZvPf3WJuP86Rk/LymRXKWQahuNUl10edxzVe/oG8JKB/V/+wOuj
8YdFxtqgKKfjq8E+ITB5zfAHn3V2vOmwYSnFj73C6eJ94w9WZhQ+/VDc43TxMsp5
w1N6lK7AtppjbtMIHIEuqcqvDMpcO2DTUA1vDCCEUimAIJrJdl1rXdaebsS/qjFZ
9YaEePR8Jc4FeZRTFTmPEE8zQX7NQsVH++uB6hRLhynHGKAx27KB9ixOhCmcuwQb
sNcBKNxgNOr3qZm7vGQDrVF1+SqTajb9Y3x6kR8Sh7RYhT7RxIyQ5j/G73XZNk/y
TK6zIHXGfxfSY728yAjc+LFTcHJZAXHdHHEZ3xE6iluRyEtrCfUkqyj87KSZOEsV
XGYQCRVS4J0RtaUzqokNuZcYCyp96aC26Tv20VBp27VzKqrScYgVWb6eTkpUfblD
9ZUQaTltX30M4nGnAvPnHvKnYUgKLMsiUZdMxY+7S8oyh1judAxA8wNPbL4k3QnQ
wRc3bApCSCHwH3xiYU4R6M7tYHP08mVZbaw3DDKJWhVTjtGouo9n32r1cERJ86At
H3VGfywYZb7ZMC7XYWio5Uk7vs4fnwFJVIlo4MW+A+/REbCEOQC9RpI/EPLyOJfJ
4K1Syb06T3kPMmmqIKxoKRsyLNLgkdg2Uu06yEh1objIljtT9lu0R5MrX6nPOl6B
NuG0NQRbs6bT9RNEBrvO2jZucEOVHYjqGGrLvqVajyTPDrhhYv8li5P9kNQlbQ5/
IAZfTjfK/ll53pWQxLy1u3VHzsacBSXBpBr5yEaA1omdckFla0XUYeaKUDJE/2YO
G8PIlpYp0vATIqy3g8HEQciewV4AlPWK6RlEEM90jF2ll0jg29/B8I8/O5h0xurH
tNd7EPnqkJiS1cHnHvQJudPDYOnYfGb5Sf+UpKX5tXMIbI6W7KpqqkTKfBxdHc0/
9nrTm1sHbHJob4o+P2c82a+rq317W/ggxvfTzdtijcbtq9PcDdCUUSgyyWqfHrJm
y4uuwUjKuCzI1+jcrGaOIfZbehrF/uDh5fGxyy6xNvZhvAx0W2Jb4ZUhKGfhFPvF
u+/JExNwotW2QG1Uaezp4+Kx7QO0CS0Khdp5vBuXP4ywWygEyeQot25p/bPI1H7k
51r/modvI87t21lfHXJwcB0gpVBuDPG1GtSLAeHsvSFP+kbk+2lcxRWq3zZkLWSs
m+Unjp25YxwZqHwHP80l6Q9jwCnGt6XWpAjvR4CxSg4i591HEwg3ecpbZ77rb7bw
RzBy200gQIKsfiD8P/ldDwVGvzVgfR2f4hIcHWJkoUVPfyjeyAHBNxC5q/4D+Y5w
CV0xhR0L2eeyT0GQP8gUlMPGcX3Oz9k3OVx7PUPeUiapDltGWJx+9Onfv13fuzuI
X4qGJRMMYcw4FBNb/Vm9eYtRWY5HdI9TvqxBygh/QdpEFGgIsb6EMsGcXpkVoJMX
1WjaJDq/Bptc8a7JGhM+r7rn0qqcXSCWGpAVW5zOJZyodfxjqwF3/TbDUj32amOi
6197MLPw03izYl12jruyMfZ/niFTF147hpth2+SgXHaRdp9T2gmId432qiY92+Q7
wfBzuSPIrZssNpb1QjXD015B8EfXAKiAHXeAKzC6FBelSmRcFScMY29VK/lB+TYd
ZzR0KIijfTgqpomKuR9BLJQ6DVs53F2tfEJIVUTVDZhPQPvxSG6ux1HUXV0ZdZg2
MV+A/tC1IXOlOFFgFAmrRIG2Omy+6MOQedtD2nvABDPDWjs6sbjHCM/o0Ctg7DkB
g2Zh/tz5jTk3BRnqx9sEML9GqvfPOM8VCNTt6rjri7hrUh/7ID8CaP5jrumaYKKF
XfrsnRBUe+5GVkfrIK/Z/iL/DNR21qpkJfTcgWsCWPfj1/Y9dz3Shh4NOF2BJJBI
kaIDwU9uD+lFCYL86WVwBcIk2J9HdIW4mA2pkhXzqX1jC9lU+ooozXVOIO+XZ5s8
qJxH5N6zqqo4me/xSxGyyyRY16Y9Xh90Q2JqUEi5kmUhg0u8wREB3ogeX5XKGVm1
qlNgBM+gsEcigVLm+KlBcKyXfGweD1d9xPdR25wacGNak34TfDkQ44lcl/ykz80z
gMJFvfrYYqv8t4WWrulBcYhnInBSCrmAsLbdOYGreociZLObOevMzMs9gBiY8qKP
Ao0JQ1pwwJE+ZZ31b6SwIfoV1+xmPZ//V6qP0Be/oTCyTnPhEAD8XRF6D3w5RvkI
HJJ6NS51j62hMyW+MkKxrIg+Fcu7/o+bf0eW+FIWwECPHa+sHxMB93Zt9sdP68Zk
3+6AJcMBJ1fk94S6ZyjBrLNLAl5ITdubBm2Cy6sTnIjDlTaSCNO4FRZKgBq3RQUq
+mUq2WlL69y44GtWBL6Uzv5FWZ2oWcCcuYCN76OD+3fSsMSWUJ8sB6+nFk1BAJy1
luT8Ncv4bbxKtKlMitDBlVSWuMeNPXvhx0Cb49SpmJ/IYlbTo01X7qjKokcEJSwn
hBh/4hldLuyMa7o1QHroQukSHQCCgJfzcOYJ7N51/wUNfP1eMox9e2Uuckv7VyyK
KzjpiLlp10m+dX1oNJityz+4GVDYgi0FhrroubBCf3M4mGRqUAyKh3zlEIt9DeUK
mH7pCgFQ+HzCecqHqgEjw8yAFgAFaou/5StfdbIkWHX5esdmMT7GhFaH/M1bsGa7
Cs6QWY6FZJ8szNd91tGkev50UWxgS6dft8FiXLT4bYK3BnwEh1zFtxn6jKU9LrKj
fPWV5bRtkq07LNfEn5ruPutlvA3J0f1pD5R9ChD4RdqdwGKBwgW6VUJ/Alio8NGb
ZEMoOawa+Tul7qByZ6sbTfj3vL2ipRu3SeKE4ZxyCJvHAnTAQcyRh9N9cdhMn19c
29SkOgd4J52s9HomV/1y7iH9Je2PT0Nr0XjoDpKD43ImtNY7Uui33LN18AvyJwQF
SM8worUmgittrZqDUyHO/BCE66GKN0xqMnf0EFWooWSJxQpMvKk2X1jofjJ9+aSg
2eSP0B3XyBebHDg0gTtg6/enwcr2AC6cPX164Ho63P6IC4aIW0UsaW6mh8Wv9sV4
E+XV9l/WtOD3XoQmwovV/RldNfViKECijAturYgbP+8e2mckF03Ue6AiFxUWqGhm
lAHmL8gBbucNE4kmxjdaewjcyqCiEaIE0DUsovvIdVUCoPiY4d7FsfpQc4KypVOF
Fz0+0Ztby0XHe97NdLnraiEIzbaWFbCSlQ2T0/0aiaKupqFlKNmWUMAmkSM1BaPc
OGfe9KwvYya77syN59+vEkJvHEDyRzWBxlLI5piXLfyutjxLpEE++DyqHIkP9ulc
DFSFmW6SUN6Zr2JgOs3fTLbQDlP7P876/vfMAurix3zSBeIrmytQmJ0PEmVHQ9JF
nurFsTKXhhPyydJyBJZUCdN6Ks/uOMCxw+qm6cuvTL0RmxR07/NO8xmR6Gq4okpi
mZYpkFdiyB5bHN0rDBHJUcEN0J5bTh+q1/31KiJvvnpJh0SgESbLRWJJ4Cvca/JE
GbyqS6xIeR9PeCtTwRMhRcWX/MZ2YFqykkhC61Bp0/pcYNLreOCnB+knH0b7Mg6l
0HGduyNmag4DqNdHhuP2Mqwe3R86u8UPwxQCB0c1mXsO1H7/LnQoaNXWOjKxNZPK
jPwhaxPB63gQ2FBuWO86wxJ6suQegNKy9HCiFAFtfIZvEmWfcX4elS/g2vLIlP1d
nmvgt8gK4+2qehGDR4PD50RZsUxck8dkdqDmUdoS8RmhcdJUgtj0n7SQlr/7F5uN
nUVO6tNQhb3yXwbQnU6pjslt8VnpNbCphRLT4ZEYji05hsCrwzuP0CJFkpx/nkmu
mtuIBdzUb+KpRCIjF4mSqfzRRvw7t5RIKyD4/mGg8Y6KptoeE2UhUmzLh3PbtvU1
eecsnyuFX1J7hYHAD3xaQ/ALcoXA9/lrRwiQ1DHXqmRN/Z5HTGir2Mui1KS25Zjj
GJRR+WxytjaQ9nfz9ZW3XZvIxKtRlJgLpMXXUuzUN7rHXISEhwoA35jJeeGzISVu
PxmfZT5rC85I0UT+C4Sg21RzGhSww+pB0YYuyw4tYXzmsqh1mMJmAdf79C1QYhFB
Uj8Phynq41Q2CHCjdMlPpdLisp7Rp22Sn7THtsxDQIHu4zdK27IAoN1VyaiqqMQR
jpoPPkNKsev1sVQCcusIU01ovj/OmxKKn48d56XN2+Z4d85oJq45Bsp0dIVYyjUY
IySogqEZqfZTF7GsqQ/bHUG0wdXiaWyj7JsY20RPvXI54YOITH019tlXrI4OCgPB
BwnSN3ZJGwdqa5rF6wkPQojfpywUzP7iCGR/KmeJRmUhODzbAGv8ZRCgokR0TRue
2ThASdF6y2hR7jLycrOzaiW//Z/Ib0+K475b6gy+7xUR7JyE5uOrEHBtmL6xIboA
mTKJk8flN8S8+/WJmLYVDKBCnpJPdhv6qd8TEFxdGCTFvM0wyICbytNzCTJZ81M3
X61CwXjEZOG3jISyR1r+9i/Hgq5F3fQFiYhp2E3DXKKUg2AKCriQ89J6Zp6516LA
FiImfgFTOHL1HNsErkPHX5RIN+X4kY7EOFh0GIqDcj5q4fxorwwdIpqnxJ5D/dst
r5C+oHoKVs7gB5zCwhdbtOAjfAr8hbTxPEy+y3j1jPBZC/+4QjX2gI2J8VsHersc
3hS/EB+/CA47zCvUNl3ARb1WzrgtNO+Ndu31NHLsNzVUCVqL1WVz8kiVKBHklYBv
duThp7FG+hF24DmpfyUL8CxOt7OL88TtvQFn7oWsrf3VJLqLsPVbZa38KiyW/40P
OnQZj/cxp1/uT+iQXc2eNjjVDFAGyk0kWeml2t0DF6G/3IfOZ7ypZBDsvaWu5+yL
LRwi9YykV7uHBa7EOugaOHoBuyrrge5/dxWvTEDYUfg4ZO43vZcIvavfNArupqZ4
WvzmBZfqBO/obGPHwJ5kpidMI7NLYBL1ad6zTytYltyUcVyrcLOvd0Ex1un040Ll
XDKnLdqfqCayRooEPcupNAAmZjWiJglefCyiCJFdvLmeTLnpwejyfpP7ovJyVoHK
OknNbp8WxV6iX5xzxJgh3Ddlq/kfnuSVbLi0V8JOkgpD8858dzyKqHNWWjQWylPV
Vwn0VlgFYFNbjCc7E42Ijk8lrzReyNxvQWCwK8G4A9WvCPAReyM9GS7HUviZtyF5
ytzEWVlupe/OIlYf0f1X1Z8KNt8KqDkbW3pmk4J13KA7Xd+B3xq7yDYaZfEC2cT1
ZkzxSRBU+r8yrnBrUqAFsEHtUSprLgM0dVwwJOnDLs+uydj9pb5+dpsHbTwCZyZR
R/dMe9qrpWdTqIKvJQtMb/BI6T9rLZv+u3pWil/KwY5S6RB3sOPgTg/hrcITgqfm
ioEkNzBAp9CP8GzeQ1kC3hDWMa+q4uqCEz467/4YdFup2LTIW+F2kzn2hppqrfGl
Zyb4NG1aTKIXYoeAL7/HNJ1LQxqRlxe5XAxEU6hZ5bNbFaFuetHs5KOmPZe2s/D3
LuAv2kaCCxhlnnsdXJ2L9hLf2Sgy+7/gvC+sKJSUkNkwnwE9fNCaAT1Sv7i06E8x
B50/ObY6xgBMHgEJHA7vepCBdpK7zRHyAINKtxYlA4THQQzNGALVeJ79fKQmmt5q
Uj73uLrxQNTJx9HJg7TQLp7+IcwPePEWYnv8B7Em9QqK5DjzPrgvupR4xnSdxK/R
rS6oGb4MaxryYirzQJcQqlFKtB/yB76zzV/RJpQf4DXAHLkGCOLDPUs3xcGjWLcg
VffMkcnXacfCzGQHE4S63oscy8aOsZYup9W7hYdXiW4C9+/egh5NHztbC7WSVmLF
lfakG6W/oadByXN9ts1urdvv0lP/fpe0yxZqabAav1u3L4weF0NxMW7ofZKk89YE
geWl1WZXwIGjKcsO8guTx8bMXVY9LfwwqktPPob5ixeLsKwlZNrtZPdo+t9NWfXC
m74MEwyWMvvj7HX+Qi8mg6dgz1Tgmu50+mr2s6X+woOxrzycTrdsMdapTk5QJkrv
laIYJCiGWlv2Z0VKiE90d3Gs5TMmtb/+ZsL0zvhQE3QZDJm13ThKdDZIJUabCTsJ
gUybnuMAeSCuN02EBxhLadu/Fxeld+McqrdRp+WnrnCAK08opSaIIQssrXXhLMhL
Irk7wWjARHhYDxmBSL6Kf0L1WhHXIR1oSny1E3wNqfaO+zV+pyAZnlZGtVL+lPwh
EW0zADUj46vM0S39XGIOrIzjSjoKFOdYqCUZRy59cPfQWBC/RZAwIhIGEcQAgo3x
eKJRD1EQD4zX1TdGNMRE1+AmtmauaDgpRxdmwPFn2hYQ3mBN7ZUd44A+m5Mt9hmE
+f/GH2/LbXtAusFyiYdZ04H5Fs5wk2nU6wU7YwgSfrpIAo+h++LSarwlmMJqaAkk
dKXnR/kVoSf1SNLZUewDvvNpKQTvis/rVjuBLPAaCS3XwiruIyepnacZ1tj2tCfA
3/zzASYAwFb2ATVE3CfjDU/+fUtpnI+GJxqtAPIe29tHLJFyejNcc9/XrEVwst4o
3ZNJA9h4iETn1Z2Js21KFqQAyi06PKZSao91yznrXyLIhu0KppITKAPfOSpwmC4B
r1r1cLi3CjZKhTXunqMfBq2g17IMFZPu2wcwHHijuZP0EshUvw4ppzhdlcbOcrQM
ywEVUCWXbb+L1/Optufyctmnf/YGnbyI9uRJDBGESJmqCMbNvhP0O/mtH58IJXvz
oWcwJasZo2cFVA5n/+ias/PvZ2kqyTicgvUXxyan1GB4Ma22BSdDCpbvqjgI4xDu
JX691Ak/HsUhYQaVQGdeTvdlPTqJWCMV4r8f7aVt1QSUK+hBgtIkopkZwOe7ixVC
bAf6CR6cfxshKkESH+4g1tcqDUaVWPoZOCNIts3J4tXFLOFdugJm0uo6OuNoAsDI
0+RqnO5rKTZ05/wcovRxLclucmyrNkR5pQImh+gaw0e2N3DlkiTcWVXozKAIJ70K
LU4Cxse1AgZCOwjoXxPhpw/Ocefh3Dxryx9MixuJLeVCCSBC5UfQ5mD5MOA7dXC6
re7oo35kWEjC+2ZOaaakjH+T3cmRNbPl7kWnlw99dCdaCl6Eev7sEY9W1J9L30kL
ugXtRTzKxuoYWEKzsof9xFdG9Jt9AbNAOA463YbeNZmPfj6ys1CZ+WHODDR7KZ96
oMpT6CP3qSJi3fL8uKzPPipMqfL3PbpxvN4mGvP20exr3oXCAO1Iz3bgoevBT0iT
+4lFns7n6YgQSRoELaGl8nkJtYLz9MGgzI6q5aNigZbOGx0NF4Ez4qZ73F3/rOBs
c8DE9kzYVlPBZ+eevgfK9+hCpLAvTwRqUup0uQndnvUfU7pHw9LIo1it8Hak/Eg4
d3XAioM593j1XCvrgnWbPrc4KVaOFnU+vdPoxLtogSZCVR6dKaACVQV4ks+KZdsX
SyKWbyFI3Ewo+oVd7+5BVnTIxibFOEzCmyuK4fbykJHzOhfddZr84tiXQhsQCK04
mm0NrMqprJpyLOQV4BlMR8CF8vrHWpThZYQfeD5lrpopwvlD/K2ktAVTzvTHVTkT
MHODNWlMZEDTbhk5LQirYHkSUWOAfnd/eOG9RunmQLXiCmvfMlowDfqqa6eSdTUX
3FtKOsW1JI7M0l2FPvw3eceWqFqW2XyBkSVEenS85VTOCLqx4avK2CyuEzkpl3dV
517kEs7RxrLMC9qSqbdUUIWHzSXXed46eK5ZuT+yevp95EgldaujqX8h6nKXuTMn
0aVpzBmJq4TSexb+vRoQ/tgq57cZLQdCFkPAC7sAM7H1PNh4LA8tpXBafSZyNQNg
1zthf4TvSwbK2HxVYacHn6WbvQc6xObDy39xt9QnYaesOzKPDdSOot0HuYlXG6Eb
Z5csEpxJ9zZFlOvrXfF6L+icujj7g44pIztPauU/VWw2sQbO+miXQT1z5p3ng/+8
IkxvkYGc1WXacr/vXwWk7F9hnLsUK4rBNVe+eLTuV2uMmRTYewPvdDXxZjXaA6F6
bT5MH6X20GAgVWnpCAl3OXeyXyfEpTDVF1auBQAqHuEg+bBax7Dj4+yuycYqS0L5
PgAInJB0adyWsBDJITfXRzcSGJi0//dyO75WrFuzeRkHu46cRbQMXKfmRV6hxwZC
zXcB1atfqkJqMUB3w7qIDTyFxVmXungzQPTeWaoBavha6ZmdX/QqEw4yMTx++B+N
fZz4c7b3xMAlQmGDc/ki6lDXnLPhD+J6UnbEaU2q8WBLmWqqKsLkEkL7canKX2zG
ays/zLEG8HtafDc8nKeFWWVAtKtWyYWxttr11S59g6DtTf2CC2SB0QR+0in7DNGC
1ryFCrQHukC/J/BbQpgLKrbKv9duDYnbRJEi8Xsna8lIDH/UVhnzlFIRMupqhEC9
2Siz6y0ZuN0Poahii9yx0r07shPArsqdKYBuFSrfcw8911IT9OC08QNDWGaRE5F4
J8PMhXZEKTCCQ6ebVpjzAt7pvHaPgtMXPCHE1Z7/ul09zigy4zDQLri/oSpfWLyU
HQIFoIN/s7ztS2nhNPjFPob0kjyNXkPR6OFvZp7xuil++XiRuaKAoj58mFbEujWd
IrtyIA28HPr/JTPST1ibqCSi0odHLv0Y5bAAAOEdKaQTxvh564u9i3/b+cTrvFHc
sfMrSahKTX+6trM/VQFilnkpFUBKrMpcEdhaIExHZS0uzep1+NLddJAuKsuhjBKT
rAzbvLaN9lZAOB5sxlyqCcubKVdICZ88pRZGJJ100zvclbuYYvX9980dlhLUCO/S
sS/O1o/T+4Gmj+EI5YyeLxkY7zO5nPnXF0IQ+/diNzQR7FDzV2Roh2U23kS+1G9W
bMXeCSbbQBjtzYXUeLz76s5CbaDRgVIbey/kuZ7aVY4bM4PpWghvCj1DxHBOZ/8S
S8HQEmsNyCHRbDHpttnYkMBngKt3vpmbt4fpkiO+STk3qaYSOGJtSnRi//usUOCW
k4IeBMBpCBcodmSC9TctkQlQI80USQw7Zn8y85mzycwf+lNMwyb+IdtXiv0islfy
yWWRCIVV2ub+CByS4SIQ6ueRxkZuRZnYW3/63nn0XL5mi2vDarZzixE1WWYKrESa
zoencaTuQxKp+FVEaPxIDmmZbd+ZQM3eyh6qyjQVGrFNS+6xW8U4WlD9hHcyN4J9
YVerfK4TD+R5vD0bdwsuqplnOzNLZ+JZAUHvzWgfb3Yq1PYORdsoNQTwqHYxmLZW
E/AOnNJIUlur558RjgJsAMHAyO6Yy1Ly94kTEYPZYQ/T7aRFnW6dyXsq2VPHx8sO
Q/Wh8/mrisIm+3LT0vYcmL/1J4z83QGEs+J48XEZXn5AS8Nbsrrc4I2suEfqdWRy
5APorV0aMl3qUOZ7wBC29eTfeq05avQQo2CCSVLQBQEy2n3vRoUedS4awcLcmvJy
wxUtDosfXwEk/KsJOts9/FMzssoNQ6fLfVVR8QYMLym+KDN209+NA0HeM8M+pb1+
va8ww9EmRTYEklVr1o3uAavPyX6x3YXdfa2WVJ+bn7phoazS+kEi1314P7aGWWwp
Pcif/hlPB3bB80PVc94FSnDTWwVor69RSonJfEttCpCq3PHDAk1sRRp/FRd4KJI1
xL1Gin1s6iOcPQELx+vd1mQ+hFAzrpPUOBwd7qPcwhevPF7Wi6vegxCz83/so2IQ
IEXPh3Lk0C63vOlxn7OB1f+ajiYDsJefxGPkTNyIniwDDljYvBh9yFlgOVjB7kxW
sH6VZADKHFUZMsbYZVAQOc9rlew3/YhX2J5aUCHGSZsGrJY7ZT/0Y837cOfKH5yQ
8SA9qW1jPL4lCuA8NuLBh66hjOc5clVOIG34Ysol2Jw9lPOT4zsYUcyhm5UOz8EH
txB/CcB4A4DXMzikJLD7tMfSFnfRrDPO4PftlT7EZ3EOEzC7BTgce7J+nf18Srgr
qyFXBKd2AhKaXiJdJpKFNn6aNDnTiYpYV6MfNYQOqDdCroIDBMnwn8Y5FW95QS+q
pdDU+vWEwNEQiHryLKciVgek1XpcJdolImywcHusBhteomqvIFDPyQB8Bu8OB/xO
2IFbvNWQxCpkBL2OsYbObQXF57OmFa75umR5eQmnO/WqpHGMCPdWMKLAPSI9nyni
EQn8P4MIpu3ZxYExywozROuSmHr5Xf4d3APuQEipFPD3d1Lbt4pJCkSnfHv0nd1n
zcahrPAATyO5fWOX1Aq/Te8U4849tgqH7gJDEA0ZU4kU+hssw1rbDVih0S1k3Mjw
lFqnbxJTspQLcKhfosz5Rw3N3vXh6GN4PzyJnGPAH0prOHpmPY8+xIjAnpAyTWXZ
YXw1qTIuAnke9EAh6ykdUwI/55Xu97MlZR4lbxXgJ9YsJDwKJgAB7xr735Uo545O
VrVu4NY04TxG1XmOXxCQTV6vUbxIae21S6A+baSsCljcS9SNjjBuZJSyaArrZWlq
pUlYegk/WGHHcVHPg6uoDoLdarOGKsUfV8F/H8GRvXqnlNQj4biBFPPWofNA4xhm
rCULnMBLX9rZ+nihvjd25SNqGeMNX0c+WH+Yv2mPOcX5l61nF5SnLxxdY1Posvuh
YOzxelDGMOVgo5sShrS5V3ZhIIAyaRNQhL/LgoTTY3tWpQY0KFtrydQZ8A/twsfc
SZtKye5HRlJY9caJXHQW5Fgbn5MTsGwkb4xfjjHLNSfXFvcKMM7/0Aw4SVDD3Nbw
/e13kJOqEE0JE7PgLJGsmqgj2+nUT6U9Qi09jgPEBpOysJ7k/9CwJ8gDJ4fvJooa
sfUomxNW47rGXqBfslfJmRgsoroweaaVfxrbApwyDgdbuK22iyITKt6TsCyfp+S6
1O3SViUP/L1KPQGLkrSPVUImi+Px9khx3GCXWD4zNsWr3tmbwJkvCtVzJZHQrv5W
XQaVQSNNZ+lRArV+VoSOwgiXxjl6qed6xYIPcgnlsuZ0fuHQGQFzaFYWOa7DJ/Rc
3zGy9lGycmij4sQIFAMKoUmw80IyO82r+GUMhfcYH/jSIHMSiNfpvdz6W5pdjifx
+6RXu/NWH7CumoJZ4ABKuNWtgW/ZQFbiXSvs8hLHpE2+M3fBKZSmYuE3A/hoBLO7
G8nDSFBUxweWVyDbzyFY5UH0xmMvV+funPtE4dI4liYPedqK0kT8fb1C41W0CD6N
hMNlVpRohlOo2RN89XBDuanVgV3kho2SVAPnppvHvVEKwh16qSJRU+1DctGL1175
VVwWya/we69yLH5j/bq4rVmne74nQTngi3DtmmWaTHAHO+neBm0J/MDuiV7wORSz
4hJyv6rN6RBuU0ZD4QZ8v2vY4rs6IXPNFjRfq5mO6AEHYZ5ObJAHO1C+NboZIXlc
P+eZ9tTDh2z/p68Dr/TkKzk/odUnBrx+n5stWkUDfs/Z+d3rXS75Fya9UWT/VqV2
9vrVxko3On5Cz8e1qaAOADLvsBCJ12Ab4sBxshO32CX9+BSj1Nw7Y9LfcVzcxxlg
dmnbnBbyazvUUS0DnJ9gcdrBpWN/V2/66MWe00PeTBkCLcvaf0AM+Z2XfEVbV3fP
dBCrH6cyUqxkCjmtb4db28VIYrFYsN4y1Ayey8UYxc9ugC9FlmNho7N3wJEq0Rvz
wUCwW1ucZbWoQUDp03/NZP0ps6qkQBcXJMh+kzyshXq3KoMpgmjbKpBMaS/XB5Ct
bz2VjJZ8OTPHqDB3SYXpdrf8cfK9DcXg0IpMruVTYSO/mai0cmn+5cU/LP3D8u4g
aSsrjAvLKv5BPqSGdU0NC5lsvYCBxK4ndMJOBVFZSxLDRlrbHUCwUFiCK4YVOsN2
iyK0qeTkAlRmPm0tCDG712B/HD6zZWDxwBSdydNUAzY7rO8LCFvfe+sPHbqEgHO4
T4MQV5v9FBBKChOIMHiV5168oxq4u7EBc0uYqAgYMLUNGzG74qb1nsmaRdU6pSvf
vrxswkVEZfqOKq11+Zk1DrAj5t7MFGJt2VFyM7kyet31vVMFQL3Zmb4rYavQk9/V
99d8Zl0DguXq2On4BzATqasU4e/qlFXFD0FOQX6CVD7L8cPFooUCDExmoFHy/YmJ
+ReoDsnvOdLJR0DdK0OxjFRWqiLEQj1S5NsCekuQC1i2eprLeEuIovmchZJTQxft
GkNw+7C56Jn9Acw8JiAnGYqQDcsxANtkrzk8U+yOTjktWTHoWxkEH8Smg67KSEX6
e3mXBlpEj4iZTa63UFFndm0JXTCIMGFaclhqKRqZO5vc8wMeRghD+0junmF2nlCB
FBsTZO1RA+mm/3zhKUXvf4luOH1kEtlaLPJ6L6S3XSE5eBZ8zxUgfLmqkzYhvSNm
awxZUXiBMKTWfULDVjxjnXWSkWNhMOhOLeEAxdsvkguQKlahq8KK7SepaS5tbiUg
v9lrLoY1OAMa4ujFUdod6wFklSbOO5X8eE72sTegPJDYYJGPDBEZ/XgmulAHuQ+Z
FuFF0mT15MdAx0+XfN5YrGaaSE72iV4nsUzqjNe9q/HbzR3iyXxOc2/WQ+DLMphe
a4VRPn1TsFQQIYmmvD6Z2wP8kuA4MQm6wOxVGwb6ZygRuyAy8owwsuuuvJLfPKzc
qdiKaLjLFepoOmvd4hfiiVGWmkxm+paiU2FJ4ukYloSiptN5UjcjYxuCd5crI0l/
pqYyOMuZ+MjBHWQYHFFwgugVW9UfWCbqd7qw1m0qbFAoLRNnow8TAja0Cw26wqPE
YfCraLYiOUdULKESvhqfRssMmHpoSDc+mfqWA1ydbVc8hzQJdlW4nJyUf2wfgBYz
EJLrQHO78b+/s3Ykx7g3BHSb+PH6AiqbvNU+Yxhpsbg8ThlyqQMCIARK7xs++OHD
FDwbv75sgcXkRKOIOqLSfgvKGeS1j6tqmOJriFBkMLxpAYEd/tOmpAUvTgfk1DVK
1uDRUxutKylh0i3mVa0ZQhg3urcJBQAmAw+5ezypkcwj6mfwL6C3KTPBKNWvYj8g
u12fe9bnNo5XNVnYJ1S1teSlKl13EvKHW9QLBxRh7i9iyBTvlrhsqEyHMLgsCHLM
5esQleeKR0Ds7C+8lsoHgqVZc/h6IUn9hSVloJaPx63CHBDRVUJQrNo/uQ+8ldko
V2pqBlF1OaJ5E9h6RqeIyBQGX8QhRSEo2PVm4inyxzWQWBqRYjSeaG8eHjxw01Ea
kvsdB43mDMsJNkWbmqeYFM3Nw7B1bR0Ah1EuWsFwruVk3LOskjMFqZKp+P+yQBsI
xZ3wVZLw93ZvTVAGXMXFm9XCce74pm5xkAZWZpsPHKHT2lVKnhxQzvcLdLsT65Sz
BhL7+StSTPXGknF4vI47RtdLMfwc7LLApgCWmMHJvctI5N1MPI3H7wjCmEdlSbZA
sCQ+ssP4Qi183ooi5T1tAdkcLzwDuKLh2V/bs3c9okATtN40ZkRxe/anosbNhjsk
LGUzd2vkygID6gwFeS0briPuXdfKGM5k5jfhQxugHIkaaV1sBDcnSArCjTcedFuz
auzToCPtME5ukrjFSf7+J9wRmATAptN9jiwEaQLNaOjYM9y6S2Iw/LDVPnuidA56
ykKt1fkhw9AjHXYqaXEoMZmzGROKjJit9JLEDHlNn+wxRGLX1sU9gfcl6HHYNQ5H
2fIrKVd3q2MW1y9BcN+Ts+cx1WlYc1jxhutfr75F8QqvLOgBRWAr75b1GSP+pEZk
eEyp3YO9TRRrtaBGXNYXsrFEDKAakSPvhOSGfl1uHUISb78O3ntvbBXRoJDOI/2P
3/VCvPuwZJ+zXQOCx352K/4oUaaZL/MhGdj0i3Mnz/V6erFet0JdpWJ7Ig/YXPYM
Vw7IkHxLFSuDzY83jRJ2wr9mChCrSsId5AQyNvfgqRLn0oRQGalbhckJVuwRIvqR
QNOGFF+WDw+cPhb8j9Ak91jgAtyHQXuYouEtpF7lBKF3YJMWBQYgwyrmyrN3IBsm
ujlH5sNC0GpJtpMh0CjWAxiw4bVMVxyP2cQrpe3QgO52xlg0CMYf3mgmLv4N2gu0
VFtbzlsp3kE+RQuPyrokPSwhqwaQnpLAe6KpsPBp3ZGu8h/gF8QEQHrBALfPvgjU
ABCIj0nj89oH36zDO++blFcU6IzNfyRFbdDOGMXm6/GPvUbbPWpZuiNqEOs+rUh2
VN/JenNmuOME88BVZqpoA5byOLUFwpL6DTweCYZ68/g0/O1PK/5N3PkNDL8dSFrV
boTqVCMD/5jXP4wrFSp75Rnr4knvYnKSjO5xQv5+9NGpEGwPfj9nvYP1K1xY2NHx
as01G6/sWpfDCkFC26cjARxw7CWcleBvLeNfb1xsQXRzR1t34hIJK0Gb3dII3jh5
GCQ4TfI6myaa7a8FxAua/qeI/ekHrZwUUDB1Wz2ZHt3NRr/Wh1nso2bT/NqXsRDy
2qiynzoSADB2mi5KH8oku6bggSVQabTrNb9EbniL6vlySUD10PAQHr1ThLrioMjO
K2GzvkBIutBsgKfZjM/j3Gl9R+z6mraoOV6P24/kJ28UvkPPWMHtNG5IabO4EtRs
q5xjZLUS9hREuxJiyYr+SGnpIA3QxDu74Q3uDf+Ds8/67yIeYnz+RyKYQGAcXW5R
YjfjyLnHGrecAp+0hVC9FD07z0eTOPCr9Q4/DVDEAc1GmaW2C8ZoxjjAzX4qQy1d
gh8KIIly4EdPCTzYNfAUxBwrPCVfm6bDBgp0dcZeVJ2g+qD4nsIBn6BKWwSeuHjt
8TXHncfY4HioZ6+OkWEJ557bAabDlQxo5yl9447+sjqZQdKXhO0Zrn0hei8k0SR5
G6bgrH+wohgWHJtB9Agi3YS1qO2k40sGs01uMQjGPbZy/do5y4wjka8y8MewGeau
x4se4jqlpy4JXpNboZmcTDv1QDDwKdZ5+qZN8me2ahq2+EYFQ59ylgPxq1yMTK9w
RWEFRryyvVRqSud60VlwKgeWfM3tMiipV+F9m7CMddk/hN5hdjzqllGXquLadcqi
vBloeIdYleU8hECwHR01HyJKC0h8SeNqdoUYgxy2hWVyrn7jsBDG62XiYXbcWcBj
6ytztT1VL9QWvjR7LPt5iPFzie6z4BWuMptoaFTzoI8J8jDBzAxeD+TSycaY/8ng
6kwKjjVm7xaS3WeR9U9rcUPpDosnWA3sU2G2LBHbFjJYp7jx8ZNugD6eTkOiau7g
Xq9nVVpmPycWnCXO+XZLH/l5OrYQ5sroSuzNack6EgTzqL2ByqdITYqU2jFuTAxR
8pIXk3uwRyD+/XzY1YO0C6/lglAtr/AV8YkhrswNNabTAeL2ivF9liKJqBhud7ZC
edgWC03k2B3W4cOE0fYE2WqyfU+H746eGdTJlUh+BGQN1/DOryQnSFKrFvpC7O+D
pl6jCHkRirt5VeogZk8Pfc5ncFEU/Mt+QqUql53QFafOzNVLzK1ebI6cM3/38me9
FLlEuzy4f41y8gF0p0NdH0RRPgBMsTYcWDlFErpPTSVChGF9S3tSx0vEN82oI+iU
+FV+ceMNthK2wXjwkbv9IJsVIdHswB+V1LRDnmeAUEpDMu31OpYQe4StgD16nSNU
xaI+4+Bc4WQDfqh1FhztTTq0PvCZN9fDzcyu+U8+3upciKzVWkAtClyFkjBpA4Cu
jsa5RQZFUi/pbQKWaBA+9lLe8hsncasnn12oBDq11x/noHROk/KOXaZheEO2dTSf
XhcMQlOxKirjMOp0enkfQyddVG2C9qCIzTtaeaC/GrZXgN3f6imKIgl66vc6FDil
yXUPEJ3EgCyQvWocvnNAGqbb6IYjrZa9GdqKZFzoicQzcw7kUUqmDGeAekvv/5kB
xMpaX4ys8szq/mOnvhHUPql/Qrx4hO8equggDUUMN4/JWnUU10hBk8ozrtyPnmav
gNz0WvEoRynCW3KZKCbfkOGzJPijP2iFfr2I6yIDFy20inKPSqG5CNCdxt4OhpVn
C14Kog1DISxRzMvnmLN1CevfUT23apxf5WV450SkfV0lDRcLpHKJElwpi977kgGq
8cVWOiYe31dDEyKCSxM2H/k1x1TMkL1vNPs6Mim7+W1rzUR4tKHNQAm7rdMxKW1B
xEm6KW02HGVaEsrV64ZzVG81Hy4ezNrZMtxq261DHghcusyL/4SwNkziWBuUbgrZ
X+sSyQ/mJDrGsjYVf7J4NM7LrNKdTpMvQVZLu5ekvE0hgg5Z+tyvNwuqob/tGAgx
5i8Bbc+FGPSJoDBZuX/V1CnBP8iLc8Log1yI84fIDUX7Uk6qRAb5sc8DhYz0dibZ
QbyWzyQjqQ8a77OZ2qUIlx8yi3ZiNsO8WFZEzBOKGaDCZe5Mq/dXvY3neq+MVe2f
4iZq6cPDFiTTh+pj9DL4NVmqjISSl+j/gaXDvkOsFuknpVUMrI9vh2jast/eRBVw
6rILfzUXtm5DAuaiZzIKnIc8RuVYicXEMdsgHv2FGrU2St9L9tcP9z7nx2CkT9l0
kWMBfSx5BpAUv4LL/1n3CzZVZY+5P6lql6usdV6EOtOVeIVhKVbD8CScWk+xi7cN
8UyuCnwB480+XXAT6E5qZ5TadSM1eXtjVNA9iCOEiqjROmBU72opu+LzqwL+6ddk
OOZ8SFuyvrBd4GY1AMwjjPpj/vpLy93vu4HzgQ8/55tLhqQnaEjojkl+fmlPP6w+
AFj8eSYqwAGNCm47oMs8STp/2Nl+/VqlBLhbpAZqeS19FuWkI1GDtfTAmha3om1x
WwNQb2nv6/WmnkzlxkFlT0jOlXzoHgZyNy89v4HlvjRbXTB6vsiYaS101ttJfi9m
/tO2lIV/3F8pJVPc62E7Dxd77vvxxl2RcAkpYa8stbMgIlZ6FDLje+mNC3tP3wIG
oe3c5jfhTXXjeKkKdFl1VOhuRE7GOFMWnY/ZvKgjXdC26YZM7ZEJxsUXn3h3dJAi
zEaZSD17iokyJ7Zf7YM/PDv57kJu/PNgo0MDmSUAWB44KgCuVPADObwRdH2YpdPC
Gq9OjixCcUz4zayZHrZtw+oe0TO4ljj7TQh2cWV+ah/1SENCv48P7aRe94oISdlH
XuMMMILjxhW1j9OTIYwZEEErtMTj0idHnjCClAta0oNHC9rSzVbxLQIen/It9iCA
ZZmrz5l9xmSsN+UH1ufT08mGNJxdhsFDNM3muddJOWSdyB4Oa/cUCcyDnS6zX+ox
hTVy1XK4udz8zwcybSj6G3944UhLBbwJebx+V5Zz7AJftYOjxG+TRIKyGHYGp8hc
1gnLzfA1NrRVx3h5Q+FYggjI4YMvomWeduqXSbNzC0wn8hyWahoBXC5dSq739unk
p4WvHUyMe6swA4O1q46ZqthHBLDuENgfLlEeEaBtKlQBHRWW1OU/59eqhA5vYBSI
L93oDnGi96FbJ71rkjymm1m6RuzpNpn3n7mZhvPSJh90dTcr48WWqS4p7ADKsJfR
ZvCbaduj2xcYvdjB+FtxqQnKRG8z9oHkV1HVSb09iL8ITtEz6FWV6LmUravw/fNb
jhxwrLMOEbgROiCSGJ43P/iFl/DNT7RciW3PihPPwHjoMSVdjSLT+sXAbxyFyZQw
b6m5Dk/aahqYRx2diJ+Dtpws0z0R25BS5AJ3Ldqq1LlxxxogvASu44LWe9PVbnHY
vWvsUcnoGq/hviBdCEOef1NUornLxmRk9apc0mlnvLROPcyU3orzxtXxJuGC6mIZ
0FZbI+/HXDNeqMQGP6k+UUv4yNtMEI5OkVO30IZ1DUK6juYlmcbDKYtQXIZL7MHO
cA6a/Qr59Hu8YkQ0cOXTp//08UCcHeuICltj6lfbsAU9hCsr1bQOJLzS7qkCqJX4
dh46Z+VF5Tmq5+AVNq5v3UL/F1VElwy/CHdhx/vnqVsKxj8z22ZTOQiGf7jmcnDB
01skWIch9YuOK+YzEuAnpRLh8j1WnzFHa0AmM6NT1lpc7EqWmIHZGNQA758DT3ER
M3QAM3WeJj5pDRLCXPKVEeeQ3OOt+i4DV2bPCcTOeS3xN44NTlwnhAXfs9ryijaA
tRrJMVqQAxfBdKDjuxx5lcmKKRSIW2jsRkNMV+Un6QAPQcjBUjFg/xJALIEQuLaP
5D8tWpfSiabBIZjGNExqZ+FEFlMAZ8G5TnEVPUSrMWtJ66XpUwqaxd7c9vYQfiMO
9EPhjU6CJn1x+s0WMbtHwa0scoRD6zcYZAKlVhfLwwhmEApo0Dcz8xMoK2D4h+6d
xcu/na9mlqR/s63OFDmyS38mI6NP7zxMohbRhY7iWJOxtayddAfVkA5uFEin6Utd
ZJr3dAg08SwzclS3Zxd52byoLxDvnd2q+L8fktznzOxgA5QXmBHBThKvbAYgozVV
KCaOULN3iXbdUo9kSSrV9alHp4/ArBnYO46RPX2rym+Q+fePQUzNc0Z/0KQEd9j0
9l3ynZZEOBegAU5KD4CuIOVvW9EQ8L9EwD5c2zvhMPuF4m7ls8RwSQi/6GS9bXwx
GE9SdoTQYymBOwUDs89rE70/uYROgKAWepXVpSm2G2IntgB/OJwr+xP6mPuJKDyW
fu+jONQcYob66OV0duoF15bbriy1dF6tot7f/kJCs/T7mhrk50SXzd4pKS6Uo8VS
pe8766VGge8ZJMTp9eWBm+eSP+ial8cWW7z/LMIx2izr5tDzJetTS+C/TCU8tOa8
LXccdR/wNvX1MwhaqnKJoUQEVCrLPZBjq51tn7+QTRlf+Mw0nULuh+ayV6QfqjZT
PwviMu49PNI4CcBOl+g1msHR00zjIHz/DJNvKdVchePg0wliwMZlBI8bp3vTGXoS
zD3LaaaN+1Pa6zeOFTViTHs+xtjXNIR0Dj1RbNDzuIplOK5xbLeB1VM2sxeCtHp0
tUVcbg2VbnFCdPXFP7ilI5WWNTJDLvva77TKLMhk9BbHn5P9hJCSDAMqnfQJR1iq
QWJwV3Lzk6NJrNl4DgrNKzdecUTusXvPfDUO2+AJJI8eUZuz34QBQqd6vn+whCTw
B01gqnC8Uo4OG1IQ2gv6df/J1/1/aqOSeLHuf0ZVcyaGdPmca7iUPRHEldw5RbXO
9Qgc5jnTcAyKyI7Dd4kXNiYOjnFq5Kw6o4Q5u2rk4AlFF+XLNW28AySsA2PqFoc0
vhxm5U022g156ToJgISgv2+fCOb0Vgdp25nzRFcCD7ksLdUHwY9H1bnK1e9t/J1d
qjBLpxin53Pu0/TkrFGXsA/25Gw6PAvTX14YFG0sBSchUhX2xLij2fBFZmWm0rRj
7Iw4uczyV5D5ZZY5sgDs+/myVL+QHWGmnKGZVWgTWW/0yrXAQTdf3G1d0qWZI/he
n8wi3VbB/MCXEekkyBKigaEwG8YDkudZNwyiEwSzEeuRs+eL3TYfnsDqrB/S2QSN
JoRSjcGovdjd6C3AxEkTI8V/XgQhCQ1idhh8b8wgrL9wMnt9tty5OubHJ8PEyomy
l5xUpRT38MZNuXx4E4OH75sbYDL1UOjdEdJ4BHigmh2Otgn8q3Ex0YOj0Yj5oyqM
sFryUi1bhq+adpPeIS5fz0bSHghmDxpAbb1zLO3h5tNvfkC153hEqEHgUcQf/MXa
83b5U298iv7sRjyxGcnDLseND+u+Zg2MHX69HJYlv99y25lSH9FwyeHtuXsidj8x
Jz9/AlTW0ZTNIK7e3bsC5hJaEm/FF/fIqOmuV0lw+Rcu7sBN7lhUmrR5RmWppfb+
0Bfsb/yHW8T8jBGQks/rxa+NBnczcBR+EdHnqPTYRBvU4DnsaOnk/A947lwOFxPi
LUj6Vf5kHE6PML2MI1fKt+f/5CanYN0JLSZOYbsnF/l8mjHmCTUThuItcxiAg061
sTl/5+b0Y5YgLoCQB4XWy9bngvU0bvI2uy3DBj5A8n/5bo5C6aCSxM7WAc7BAYAx
h9g/pGP1IOoFs0l6hlDhEXo0zswjUXcP8BQzayQciBYfvXVjq3xxK3u3IJV+lmSV
4hc2WY9fxogQdCy/wvGd/lm0EDoaS+pXk3biLl8bmI2WtiYB8ebqtHzetpUM3SFG
vdkBwPiY343hztFvk/CrjFU1fRQyAnzLW5O4Cwt4iGT3XKtj/UdWA7rXsl2mqR1x
tZQaBAtpaSdUtY8j5H13JaX1vTLX/fH19imMyfvBQZ3Le7d3cI14X4mnuBdpDyY5
vZT16w5rYHpVnQFowPyyt+YhhK+0HZYPh82dDnW5tz5NcZAefeUV312AVtHVYcMD
zdxFvWbGPjEdafOqLX3sDO1DDIfD8hFpcNsrNorJyyxEmZL18Y/8sjlLqynNHhXD
gJu7i8RkD/55mGXhImUp8IuACMJihBDex1w6Q1X85bgN0pZO+7P3BT3sQ/geDWPZ
E16gKx30P7wWg73vq2Yft/gFBep2XFiooMzQo5yEpKE1NIjsLVRzt/ARn0d4LM9M
Hx6pF2qtHM2wpNr5Sw/xzNXVdeY0uDAHNdkyAlvgt3yX+ZsC0jk6p1m5Oup7ARHC
iw3ggkdHYwc5YU8m8J5CxnA08bLmsknkysW+M5QmY4bv8URUeZPErAImzhAKyOZ2
ZjEf7OMW28onw9t9lBTjEq2TD2HGt/yX4lpXRc6ITcb594XARwwSkiv6YUcfnGzN
ML7z9NNxK3EeD9lofEYNhyHI2suWkwv1N8/Df7SFT7iXLFcdxlO/Gx7wZ8JWDvte
9s5lZaWgT/DbyprBWJG1SFs+I+B3Joc0oApjwH0rOOkpk7VBqHWwX8NohSEcpfAz
9YasxaAWBvD1OxHiH14nlpCAtHV7Ln+gMXoGT2gDwYoCJ33u13Mn7T0JRP9I7Aqi
pd6K60zOWuNL7PubzPBvrbEctgG+rxsxkr7UMVdJM52pUquM43DzRuCrvoSwqFqL
2j6b+6X6Gz46EUz3oZxMlaKKDYE9V0Jj/iGtcIEhPSEyQwGSu84qrceSh+88FikS
SfkpTtnJUwPHcP2WL4xgKJsW+gFCZQcvLwVY0SEZxFqnXyxDHhgHKo46DZk7yFlX
oAjcv/kWTrN5iP1NabUh5bNSG6+u4N1Rj9mOyJ4HroDtNI6CyAckF9x6eDYQwfBY
U9MuLRDSpehJwtPbzJmpFrcJdrEajG7GjPWkAaPg6Jykf9HOtdzkJOn9SbMzOVo8
B9r8RcS9JSdvNxMVgNGGyxir6SRXqh1SGatlsXipjlyVnE7t1ufRv+tx4pYFDa+r
mySNU5FCJ+Pkid6vAni/T6sTLUuWyFgmBAexlsMBYlhRIdyygNv0bC8yCEuqkuk5
cEgC+y9fagRfMKS4T7LNYz9giknC0XkhL+iR6CazJlp6opLalUS7RGVZsKIDx+Ht
W2ZjjyvSsh68gMm/3rFyj19IuoHJ3od1a2go+03kVGAb8CecubLWCuDgCFdanavA
+YzLbAPoPRJoR8UAeK8hGSlNoSXHodcqJ/KfFE9JnWwfD27QtWQD6GQQK7SF4/hv
soJ5YF5S8ExA2q2QZ1QJfgucY/3dYGR/0LIwhBh4SZ/Nf/nVhE5iNog14unW0rn2
YT4eC3YjzGrgfuDNSw1LJ0hkBRtuRbbED2MXtzqUimO0hu32xuQgGXid9LxYn6FO
s7XC2RPLtHPDruKXPWJv83yFG6JATt0nlbVYh/StpYdKF8Rt3WFCSQsSiDVulbbV
GJ6G/7RNMO8lkcfRTLjoo7TNL8IQoBFW0o9W7Kr7NMLPn/b/zh6SwuFkWPtsNNMt
M/oSY2GGe5P/vEaHvu5PlgJ7bTyYbWqwvWqNZ0NC4TRf6dimTuRf0ynF6KIg/XKV
SFzReugSamMy+YaLJez6d7QIcAQtZTqYrR8R3mXNtzAve4y6YFF1RiF6h6fdid1K
uI/0yiZeKwHsvoZR1alGj0a4mG6soCyAQL6e5V8nBeo9G6iYDJDQSmpr/ghNO4pC
NuShkkMFsOf69G6Nxc0+4msAxAbnthEmHxNpWXGv3B7+mAOLwYdICjYh2iU04rbE
pSho1ovE3dCE9Z6wGK9K8Z3BkuJ0SEBJ3GXIjN1c73hAe9ptZncZi7u8eWvgnYUC
KFHA845g6sj23zdOtVX43TGN/N/sTc55IZleDNwWzd1O++icQy3sSO0IJdbsyy3a
Wf+68ihPpE9dKNeXQ3SkDqMcIjByCRZViL+xs5swSOc/eKQU1QgzPNfr6zCDbNe9
YhqfnDQQ/v0CjOuQFrhKRztaIIHz+fGMFsczQXVkKHXF+RaNyh/ZxUEHwF/IrCBb
uGJzMAIRQ/FIY1DDyD2pNVN00x74+g4c4STnrRsO3R1EzuB9POp1Ni8FZydQH1Nz
VMlFCbLT2dck5u0Rh8WJvwVkFv4fHNyuc2a1uY/njmYs+dyKR8OoAaUgcgXNzFi+
O4zds4H1p0fcPbjsaM0M/LEgi3j+siFA5zQX1AyipHvoqKd3VVnizJFqH3gh+LkS
JltuOxnidOfaygHBopYXHqR0Q2qQkDC51RlMA2UGZcTJsO6ki6HJyyxHUYvJYcuk
ovBV28znkQ1HdmVsgMnuvDOLa0FmSacaa5/A7niL7+JCo549Iud6Lw/orqUB3HGs
mj+jffQs82yzaLxzuHDVPt2z+bmVb/3+vYkVREdhex8SamtGb+klCswuZDq6LbOL
wX1kx/q/mTqskD2XQ+axWpAMXdxuO7t8J43G/F3uxp14oaNNHdsWFwgHgyUrtXeP
gxHN99BaFUymGLxXGqFAr91sA3qcA8ZsQ13sJ+pkBseP1aJKIjwmja3tOA+8W9jP
+lwwst3G3AiKwEjLJrwzbqn6OalKC3PfDq8GiUmWfR9Ko/WUOngjnXTEw+RkJWY7
FWmglu39higv5Wz7Z3T9x0d6CQS4Fg7aXjhSkfDKGVEgB6bNSWKBTYpCpPRDXd/W
/YRpDGvS98aWk/GHQotpo1TthjkueNOKwMp4lOYiKc4Z9JYzaVGSBgV5pT7Kf87F
yZ/RNGz6Pu/JbreT6eN1Q2itSaFattWO5RwX9nMw327+fCl8xiDHPpOEezq1DmOh
QqZO/EXb6+M9LRddgfeucqFDXUBZcXPjhJiAt00EDqOHgh60VAGah+lNUUAHSjJz
kA8jPYY3Adq1EG81vlk4DErXQ/CaJY8e+zsqOfBZ1fT0QjoW24+jdfQJKSGuucpP
EYXo62GQDpuzw105n8rDtv1MSRA4To3B8r9kEG5qt5qkSWuWoIgs0fDC42BqrhnI
244fS6Ks9KP0xndEZ1xCTqYToiaoJRfE9GMAXC1K6WreDJgA27ictEb21VqTjbKg
6vf1/UWm5ygqttYFqB/T5Ea1Wlb9LNW+QDoXyvESIOoHs8xSj8OAixD+fSkfANXa
UaWiCjIu0LzxKi3tNu7b9d+hqdyqTUxCFa9fp8020Vgj+Lx2Nnt3xU5WXduVsfE6
8pas9MnmjhQsvlu5F30QOdx4S3vSqndckpOGHJqKuQdCbZvsAiXMnznCYxI5ILc6
l+S+93a2bma4STwclccUKpAZEJ4836CDLBViE+0AltkVNGmqQ+KV9Z1o61FRaV3U
7hRtlVQKzKnW/fddnhpmrIypsO3r200tKnrqUXCh4joZGAD4ZtsQVOn6cg9Sb3VY
4Iin11U9hr9uwplADcadaNyr16tMoUGUuMg3I62w+6PhhAMWj2Zq3KQsbOzug/kM
E3tZc4FuWCZTptZjvVhzfQMb0MYA8Q4VciZi5mbxh3ejOnuNA25JvD/F913GsUPR
i8fCDpuYLKU8SNwjZ8A4Awtdrj32u6nThnbNVPKR7IWW1B0SJv8RmBDQB2f4wlAr
ey43pvPaegBEgPyJwryUTldhN8qIYx10RJ/PckdT2heNlDvlbgYq3zvAHhBqEMrT
xiDN1PSY6P2JLAqrU/8Fcej23YjldIJaSzpqIHmaEhuUh46LYNBPqeE6qf5f+FLx
espcbOmetrj9guXJ+lg1+0uch1663TBvhGwy9HjmruMIXYdnIa88fRjv8AoHhQzz
VkO/YRCLxsTzj3noIBaL9icmXifCoFVCf2VlIbw6apM4IZ5+RYYgQLaquATylQHK
A6++4nGWyhjWNzsXx6JJEaVvnG8Y/YYKcEihZ/Byd+RMU7E1uppc+qmqgxeiaO/g
Yu1716zZHQb522WBhnrgSGR2SVN7z4eYviuNnAJXXsG5EFIIKR41cdUeYbRAik5O
PLv3x1TSwj+zgKvJvclPDjckuDZGio9s/1itKDFNIuk68s2ILs+Ezff7nCUrI5W2
JV8uCbceMdRlyGXtr++xpnpLsylC6s1Znvt2JKvBdyCo3PterCcxwSITiHO/28cf
lhBaTfuu0H0el60gA+QxbJMnFacwCmLyuvCJQjhpfBxRpfh+kMf9qn2knU7aZC2z
D7db91Ae/388XImkO6vrosm14x6PZhbmHAm60Y9P0yB4RH2HxXDkDwkRkmzaoJoZ
he0fbW0+/zbZM8Szi3PzCRVWA3bJWqzxvADYWAig8CSK2BmSI8T15CTBTbF2sFf5
Nm9kSj9XbkZvb2nlTIXmdcSM3jYe1ugvY5N4E3ea0050AKpO+WNf2r4rQO3ri9nM
dhPpTlWuE/C4WiSasQTtvjqO2O0AuR5dRv4qR4xGzrw1tnp6C8iYfCgewRPn+7Y1
LaY75cNw6m+Qc2f9QWEpybCmS13iZWkkhuYGjvWSHD2Pn1qXCGZ0eu8GBTRnzhD8
2T5FmFAoYll3Wq6QFArnhZKx+j5SK3HPC2BcBhUziFxyZliXUwKVtxyFNNQijCBX
G/dGQAboQBHa8upsOk1I6ybjChhqZ0Diu5M4GO7DuFERQki84s4dOU4H5oe0R5lT
nVnxdFBpeoshCh8jRB0co8jdXI87gb3cOI0An3oHdciI8a984RCRWrJKIZAlQu5w
90U1dK4cTTNCw/Bpbmv2luCsEMA+FcCODK7nwwtHIbc6E1s2CTJ5y4nQ/hLi5Y82
Uf4M3aRyZ2QIiSLWU/rvXQPk2wRQ/vEffE7c0cX4lEY0GtbOmOYslrr5riqzLsiv
ByvHg73nOARNIjeEc/GULgKhrN91zCDPrIQfGgXdvRyZv3NWqBaYUU90HwVwaBUb
uGwqYRXm/VLB0ydthShfSc/aR8wwc8FR9i7G3okZ12z3g1KAi7+XQlT6DZhgkhQQ
auNjbym45AEFpcQhuWqzxutTWf1Cx6056f4kAhejKdaosZCuG4rdrFORPjuc4bqz
67uFpwFTb0MCtG3dn0p286poeuY0mK6d7toMoU8NUoe8uz4IcgYCDYh6I/u0ASID
de5xo996SPxliNaDN/L5mhqfZhNBEcxaMbD1D6rxa9H/tNVj0FtlxQqs/pgKNnuT
fhomzvQuYG3AfPGeIr8+wUZ0cA8aA+c3rKXHQQ8a/3O5U1Kz/KLWLLB13kAS4pGX
BCgArGbhvHZ2ABhKF0Rmpcj5uvtJge4+TEiXUsUMf5NjydKHujZzUdPDiHBBktxM
fY3WU5L0my7QV5SkYCdsTavmVl62Y6eNVVmsV5jkQjjXIHf0ry4F5Tf38XgyE22q
C3mUZ+i0IXt8U+FVY5TnfDSRWDsgMrZfn47gxvTR1uykppKzK7Te4+to4D4HJ/eS
h1ieC6oDRCp7zbnUApsl3Jelyee3jeZqfFWZi6uYdyByWGoIpW8n6BvCWD1AVuhh
YPolYY97uCEyLzq4bQTtmTuLZr5jVPxNQbtZvCjOkcQHzTu6WnMANeFww8hW5yik
oUE5Q1uaqLt7A5vx5IxW/P5mN+werJpkiTTe725r1s5mbxU07nHqjYF8WXKDyMFR
nKoobomBg1zsbBrr3VRRokZqwvuoavdrO83LVQhccT2SRImNOqFRpIZcE23IjmT4
ktZxJBWKxFegglENmbDWdlFmWisWCC/O8gfTvw84Sn9Y2SE73ElsCQqUOsRlaCcv
4RxJ8hOTh7JYei0diJ6CB1cYxOWXJuAzY1rCqUJ6A6RRzd5LJA3/pxJa6g3HgTZp
1g+nnsavtvmSGaunBt45HahSV/98pMVlelI/axllE8sQLZrGH9RrWKbnqq5mWdee
JUWrFSTjqJuO7BglCjzMMQzbEjNNfM6Cm6ivxx+ysjxuOidSb8hg7iWohhptueb2
FS8G5V676+fItdjyPGl28hmSKPKmuJBtCYTXXBYZfSVkHhKPds4ysxUvEwT7LtBl
HhAe2XdnHvfFCkmSlaEvLxyHOLsMtT+Wg1+Xxrto11JOkwxGB4SdXTDrtQXa+vB0
N5FY41yLsQEGV67Wtlz/8udIxVDLdGnKI+1iGylwfFs8q7SJ/l1VpdOo4D1zfJOI
ymgd95a6E6iZrcLVX6n0USp0r1ss1iFOo+0MDLHYRtm/RSETND/2wxmfHrxUuxpL
gdMsuzCx3X1UNMu0s1wuE3OLM6mSuAVbhSwwQyXXxTQhQTAi894ZL7fjyj5CtUkj
1wxpEnxQ+2Llp1yCaYA7AGuvYAw7YQoNThkp42ZkyaokfpmZNU6fPlP2NduFU/Vl
dbLLQ6VWng6AXs21rtIWz1TnDipoKNFDaJMXJzgiV9LHUxXfWHM5KvKCYl33zGKk
5p0rZBSi2BJMc3als01QUJttP/nIo1USMxAQNiCBWjRdKX6Mjpt6CwT0zXuvSJ6F
swpGrvHRcNbbFEXiNACXbTJeu/HAStBTeRgAu529wPNTNqeoL2zxEcB0CYh+XC/J
+OxUGgv24Emg35nW9UYfGQ+nMW3OM2Bs1Mfaq6O2EqlKmc9o2WUunLBTyDXgRpHg
4bt/0OtTYpmI7WJ+dV7qWSq3QxdQ7JLg5iYJ2eMIdDhBtWbHs6c/uM9KJujoKKTz
r6ULQVFdu4/kmGeg0J4PEbrEDjuJY/zL09bXy1xlEOpceMFjs4GiBXJJXxMVjyCA
h0HqG4yRctaeX3ti3m+Jw3YEgXXikQ4H70lpB8N40Ng98H5+qzPZSzHYqDiOg5tp
YsO8v0lc2d3A3i84tUaxegr8CARWSvAiV6kMHHk2TSwsZqnButeEC0sFaEj30W4X
N20lf/rvWXlsbcP9OfRw4a2PkGZYVOIJZOF7A8bIjy61bTyFYDL7ORslXLggZbEP
JXPTuY1LeWsjvt9yyDJjvQ1AcnLnrKwg16S6wSVefHm3Fj7mEg58Ho7aJR6OGqSI
iW+7iVbUbB+ry58g9NqOoOxgrRd0khrxH7zmBrHSRsiA+JfSUL/+p3slIptDjS0t
eg7nkhLDJ+p3cgKdO1u6pk5+5Pd+ICVWRlX5a8hYRPQg+sKzo74AnF91QWpQ37In
y2VCPM6SnhLxHN0g3G/4c1Hn3g/Gh1po/bsijCvWeqmDwY9QOLS2oCGa27vZZnHc
x8L4F33bNh2RUrlf2tC1vwNS/OhccxdmIUBWzH8akCbCP+iPDrYxpPIm1zfK129X
liolVMf99n5Kl03yIpNhuAoBSooB3dOsjzh8ik695URSMQZBU3QPDnxn7PnWORAG
r9T1H3yOJmMmDHUEW/2gGUtLGWfHfS+VAazaexCi1QQw+jLvJrraanBEmo/6+39F
HChj/GY+M7oVOTrQiIxeI6M6HaEkDWIk3s2NqTQeAppTHVrOo+9Y/lPBg3LyuGSL
icSNW0x38tY7bj4eZGOmVIWJqPiPUFMf3qcBbwje5l4h9oSXuax+No8CjDTSxpQP
K+l6jLrkHy4nhtHScu1jWy8zH0dKuQ9uKcl1LFp4k3DO70m2734jDvb1IJoBV5cD
VNwubHD0gDIJ0jKM7Ja/mVvxwY2HNmP6Xu1LlfBpLCndpfbkL4X55aIxRvTWqJIe
oSyNzhxDCq+ada4JjTMs/h//d8NcACcCfJsMI244Mwog61gLODpIjQKhSaJxqJlG
QdW/cnMP+KZd44GjQtU8Na4bb1O7VOvno5xj/z6HhajWFhob9BGh5Bbw/lz9r19j
jyB/Xqqs0ZPsDfEfTbOsmkgO/6v0CltqhZKemnwDuuAmLNJkJTgk8ip4y5VZlsWQ
IMKZHdTIEteZH1ho+ocyaiWW2t+iVnxy86jy673N9Tb3YqfxxSekdal0/2X8drHL
EUpxcjBsfY+RA9czT+fdJnutmVxWkwMtXOEBd2elGKegJNNQLjP+4AvVKu31WgY5
0TY6LWL/v2XR6k9MO22+qtvOpUcd2GOqsGZmk8E8pSUkA64v/1EVT30jP8FVh9t6
BdymR4d2NRvngp2dQLZ/QrHpIwWsNkT5jwfSj7d1bGQh2mSYdfqb+xjyYBz3sjKs
Ar6PeH7FcpVHe351VD6zeFNsenZrdAm7DCU4Wwk4MCKJpgp0NgVcA6FnM2GRi69M
LX6mvY+dU/ZGsDWJtNlYt0Bq6Kj+YazrYy0LI6co0xb+9cN9yO/o6iOD/ek0DYvA
OByPQ6gE77T996J8VI1Oh9hcqvLjHUEUfXa9rskcQK+2l3a6zP6REFlrzxZkTBPQ
C/NyReqGZyNkozlJMtd918SBMkedNb/1SZDmIVtbeMMFYVhG/z4s3qRAgw9LT1YX
HMWbN/F+I9wZjgtEPu8S8xFdE8zPvvgJnqN+bBf1PfDRpjU7phj1ic83JECbHC9z
zsVW9XIAxIahBsme/CCaJRxyUYxPBIIo1ZezqO6jnhCBMgcv4LRVvHP/oxqMSBj3
Du3LDc6Lt22nTuYEoc4Q2onp13UlqOhH33U7YvBbF4Vzr05dsfJoH9AvsMaugwjA
ANW63bdNpwDXC+tNoSyVAm5Gu3klDPXwgCic16sQqO/aj2P5XRbLYfXDDVN1If4L
qcdRHGdz9Xa1RTvNI+iCEOBvDQYeuieQwCszK6QRXdxAdtUhfIiMhh70fhdYwFUu
mUtSebVVSwwnOw4Nl1uOAq3ODoECLpAAyihHgMZLHTi8isINQgrQ/vmxrMVekiJG
s5fj8p1pQoJ2BtivZq/KVLKqgxxVG6KRV1SCdAOy8tdWAgRijY2+hp0PXT/71Mrh
a0WhsdJ0qhIRxVrwQgnwuu1kIdYYLY8cY55QQy5G44MV7plfseO8o13Opl5tcU1M
8Jfq5+faK3FfiJb5Po+PbYqQojziic2nbaUJyUw0Xk8azGijUyWPoLRgWgx98V/T
NCo9622dnEJ0v9cOCp25fI2COd7jclRJLJYGmM1niEtvyjDEZJqyCZ45unL/DE2O
cW1Mtnbgn0TJZkyvpvkX1HoxlgGLQakEFZTpt0D1FS9VFno77/NrmIQ5Fa45JZ8h
Pn9OLcC8PWn9EGpEvFbnhDuzoYWPSdBi6uropOl+QPh7WI8d+2LKalpRoXD/kuij
REr809tQrkHHMW2QymOK7kRBdHzLWf8DCXpvkzMhAiihFc2yaoMc1M+1h9yrzXV5
7EAanocCsVS07vPXYh/V/xYk1oNJmegcn6oTKgGoQzjDQ+auVuwKdxp+cNF6XzCK
UHDyTKMl/AtpyX27sV2ZBhSjA0fpobWiLF3Ca4Mc/3EoIevpmrkb83m5njwBgPoW
IdDJCwfXMOjzZ0tvGKYD5jploX+QAqOLDrPZyNcQCw237Go4+uWDHMcEcG9e1Paa
HpKLHtxA+osL1tvnOUUtEP6aAWAjhfAGOb8vsJObg5rzURAsiX2xhSfj/Xnm78/r
+IXBrg3Xst9Xvmp78sLmsh7W/fuF2hJKnzjjc+iWmByB/El/PD1wkJbqK1gsXAaA
4hLFoKXOZGyTQoDY/wnLNrHcM0VhO9kYKaHYKm1ghIU61ltHUoE19ON5mMYOUO1D
jASf0uqbdHBSpIMhHaTaAPiTvDIFTKqAXq8K/4EZ0KZzmNOZHd8Evm2rX21G1V1Y
EJRI8a4AKxqN8vsucWInYe5qkONt5LiGp6ceeJvUKW8wjA6rdWdz690YqBhKDKPO
nSxunycvxYj9JJofpW7a5t4F3NCePvUecPtokEaIFh+x+nJGCftI5to5zEFO2Wxi
oVGFrtu5bO3EB+jNlc/V7WeLzX4ipFjc8Ow1+024lv3s8TMTU3tQ9rmu/M23qz2t
7UDk6Ed9b7Ohm9ZLqUyTBlfIH8w9Y0M0ThsPQqFDiDyvSwwCBmbN/5MlX+kWVlnC
0xpegEKNJ6AR2KTpaQ4+Qg/A0MuA97A6jr+xQuki9+/vXAGL4bPjEFO3KEBFm9QT
yAP6efm0amZPiHYixVG0p160O0qeJtbMXq6VGo+U15yq2ITQlCUpimmQn16NYc7z
DJ+SvLwtUndWTCz8X+g33uV9xziloNz7E1GwNoV1BD+5WsCjlKvgsrYdEarX8Mf9
+WDJnyqDvU1ZhRWFKUmGxJRZObbgPLQ9V7TBjf/LCg/pVhxybmHhEnXsCUSt6Faa
EIuI0ilfC1DmggYucixSKiFvvaJ+11WlgP4dcykR7JZG+BqcXEuDhsdmXERrpA/k
FASQHMu3aoe26GzAIQnrYGYdIrpaLoUth3aQHe60f0wfYuFbNDYBqMIVBwXqx21V
skYMUvD3kwtexGDPAXgjtr+IIEDxbTOmnMdjGkwFMT2P5ogHhSOaNj4Ebd2C2KEX
m+i8ysHRc6Tj3jFB9sKFB8LBX/3qeGMnEDDqGTDAouRKbxPsjD/+0p5E1Qy6NDxg
0qg3x+L1d+aMXU1py/JEAsHEbpKUmugsOCFK0cnRsqJF4KNHi6claz/X+2PW3Lub
LwQQr9nsfnbTjq45mgRB4+9uCyEt4l9U4taNsCUBDMwt/7YG+e2uIyGLbNKJ3iPb
d6CA2qmNWbrcV+Wu/JTV8T66M8YfD7EsuGiXYlJPT8iZ33049BwTZS1+DGUEfxTH
Hlhfjh2iWApR2+IzMy7mYeWyWB4fAQZdLir5zcg92vGPm0xqu4Slt6qeI1izNOw9
PqnLr+ffQ7TY5OxS8B5wyouUEIVyYN7HEyLwF3Qe5LRUEFb4DTdgjAuKPg/OeyLm
6x+7LFZuJrFiXSGlK++BRzc4PN/KMczUrrJ455a3A+7j9sXN7rT0zfzeJoXBl+sm
gs7K/Boz6s6lBEVkgYgxUcXvKkDrqykuCDmYKVV/OghnLF01O3F5u0X0cWiV+SYK
TX39UQ+vbHSoBjPlH9hITYdsTviwRceGMrOvim1SCTCnvhvpbOjin7cEswDDvR/8
czclsHnhabhvoUtcXHA1qnNfnAyIco1Wmcckyg8TWQLZtw0pN6+SSpH5UsecpWin
ECHtqXRORiFBAvaYnk/3PcN3mjUhy+W3B0nlouA3gkGus4o2p1AnQmHXuqZ8giTR
ZSUAcoE8QpuAMvvehL7EUaXxxMoy/VRjiI5Cv/D6wB68zbSCSSYSpeMpQxiFuVDv
f6P7iY9rDIoMRqupZTVRgd2Ysl/0K9gLhCSVEqfY6jG2PO4yb8806Ue2VDV7Mpbb
jSNxTtmvyKR8x+1uAqFvdLmDJVhaKPQmd/BsnUhh9T8aAcqRvLZ7v+rIF2p9bD0c
IOHJ8D3u/f+/PCPqOLvNxBBfRck5xUPiPP6xkoBXpDggjVOfCjBet+Ox60mHQAhm
IrV7otNUABjFjqyGm4uXboDmp8AHMeXOQz6/5/WNYZzKiiUWaOBAEWu1l2BnWg5I
BtdTTraGk8LLPxT3ZDZrHGplHTRXbRi4o8c1Bmq/cHKWHN+zDmtoeWP33mRLqML8
ma48U6X4H9yXpDSLaWGUFutIf4sY7lFdNNeAEqTo8kpYWndJdZ5QJh30EXtmxoeZ
vpjXqE8Na9rANNDkvxVIS6ciQFZVtY/q+iRg1UptXIk72WaFzWkqmOLiWmGjiXyQ
lf2TOzadLfv2wlYT+RaNkYQkgbZgXTu1tJ5tZpnKZZUyb0iholgwrqQPNqCXYo+T
Br1YzTdR/90Mxa/lYTSw/SIHPeBu8eRa9INo6+PGnhgY/+ffvLloFXvxbp3b4vF0
4LiFFTvzjvIOOVCOa7GPEU6cSxlrm0iGq6CmpRSwiqRobX6jqwvqmG76T4BPTDkW
qdf0EERoFtDbV1iwp33w6rOABAfw+7rxGPJGDue+/PCE+qUY+lNg/Ep+TcVv6BBn
sQO0n53vqdr2pVwUUC+QjTRmEauG6hzrGBVKUZ4ftEZglN5w680ro3FF1BVVPSmI
T23FDFFaPMyr9F2NUbFDgSEt55GgwbVLhxY41eAFtMv6cuBkewAdhLNCtQ3RJSjv
cUYhlqV0Q1cHpDp7jBgzW5WVtN2eqGHhmuYjqeJuoYkPxF04ca9+6mQQDf0fNswq
OVmUqkreBeZlBzXBe5rhmDoQZA5eazX/rRK78bnfjY2hbKGPS4G09Na5lgS4glye
gVh8v4h35raZ3tnfHa6YiECtEgIV4WPm8cOddZbrfhkzJRi96LlAC7O3PpHDKoOj
xjJPupF9KHLyDE5zTCVW+GSDVtTHTk28+isM9InYKmumzt7Dtz2wwEMIffW/T1Lj
BQKGduEACuFmBLacG/pVX0QPEZdl3k9aDgffpyci4RFn+hIjOHdT8hY0nLN9rPlP
s/W/OFB17mLUYiTWZW8Wm0iCajZzwh5xL71Kl7QFjbYOPH4xbJeanEawHZZdFdSh
9gnUrLG3z2w74bJJM2YYbE2ap9bVbBEJBJ7Id6I67UDuAhmyZVj26yy+5cLK30Es
qoWcBp9QkPhArKqjvjOHP2yscbbLZMf0VDYW91qjkJsD5UUxb6cwKvUDdfg1un1w
g2iawqEPUT+y2lC1+EnuAQfEl+rOK9oCFYBSp2yQeIA8tEZFN/aOTICTUgjXW+Kb
WjKOARQH/WR+64UOqtX8M08LgPoHreO/nCJLLNPn4LuglETic3FWnJAdhVUPJ/Dk
dEREVmFrCMPzJH6AQcSVPCdFBpq3o0Txr1Vb/lc9y65TSP5FqQyxwZJW8/pHK778
9YKQdpRkdAhx/0GeU6rcYGLp6lzpi0oZ2U1pXG5QuKK5RTtIxL4Vj1Wd+cvX9kFl
yQ02qBz5boPZsXTGB4nGMP2Yy1hZ2X+kFjOkSmoDRhKcRl8JN1RkGQNjD1eo1RTf
/3G5m73A1uS/aPsti0DAbg16l7lxmRnEXPjdtwyHc2PgBLxuviprJujlxLT9MTh0
bwWHJd4rEnR6d0eO5Z/w5j2d851x2yymF1PZUghCI9Pv0N6/ENux5ol60zFpd2Bx
yJVatJnweKahoBid/o6LZYb7rkTfK+2YfgSmGxkwTBc3ilKQF54yRjnOPzY7JZQ/
56E+XSuJX8e96XErbiNVg18mD026dR/G5iqWGLCh/9JHI00OX3aw3X9CMBiMagJw
y77AU8RbcDMF7DktBQzvlYxwa8Tre62DsX98cNrqib6hjqJp9J5VQbCVUZuXzw9e
/Pgy2X2cKU6AozWjnmhj+IyEYn9D88YrPkk8GKFAYFGrTJHPfnwjsOKhgGx/pum/
0fF8ATJWhW1kkgbIORRe5AA2LSjE4n9gEcp4X5yEkExgAdDK+IxlRygce2811ppp
uicsQOQqG1xuzuyYpnVdk5C06SiFRfJLgN2T11sOZXRVGB2pAbPpT5Fu/uL6Pql1
AV6lwtrmuQLh2LaB7qJiUPIxlQtK622sd4ahFn77o4eO65kkjkZipkpI1yEekGMf
dd+ESG9a2KHPKI/Zz0UJ1Nv5/l3K7V6WMu5XFD8355MONapaiBbJUIGlQ3KlBi5e
swfaHX4mkKXsOG3YBHt+/+8f6gdDTdwm4Jx7QcuOzvlwdL4OnhLWIjwtk8ufWJ72
kMLo/2h3FecCZGuasypO8rJVVqEBY8XMau6juGAewbMHSbjZ42eI194hHhxR8Kg6
RoksZmU7PHDeo4HplruhaL9k8AJLDW8XqKOa2rbOOkYyGaLomEQrEjgQSSfz4hx4
s/fqcxqRxCgv7AQFZhbKlfmFSGtT5m6Gk7lNEXMDQLMQHY9uT90+CVXNSfLoW6EL
+m0K9O5uz8SJrx05GXKZO3/pwzPV6exmmAB7Ql57HunNMXUwbc1pJFwX2qwAueqq
MFtaEjkyoropAgJdF2UZo1v4oVQbYzwIdoan+VADUl/uukGrLdiqkJJbTVWtccBO
YB2rMHJu9DLc/uwOr//avEQ2j6aC1XpbRcHnSNkEom4HkEPBi/IL0gaobqSCV6qM
VXJVcyIEN62/wAU+i6vreCbk6M9pnJLzTDWFWz5pyfzFb0ACFAjtJRqvAFg8F3vs
PhWjcmN6yqfUkW79ORbFz7CNrY5TgDOpI4c6z29JwQMyaC1J7p498XYpGLFoqol+
kuRZsrlUzwAtOkdFo5XZt1IcsvC9qiick9HDGPjtl7kxEZH1tOPFjF/0xeHlZN+g
NxBdCqb425HNCLzstxQOeaPWdd2pNEIhKd/Zt9VzgPhCxhEk0dP7PN3FImDLWWxs
X4oQuJowKmjMqEqNuh9ttDdwOOMhkf8mJKa029rDv4KH0xXYet7UMhSd4PcPqmMZ
BqidJGKYnTalbkoFPZy/kc4bkT5DXJyOV2rEyQGHlxvFqAvkSK3HdhFo55TfVAZI
SFMDwlmlv28ZKtixsBDuwqj1JrPNZ1/IlkviJpZgIzbmDpS9M+PMLPHZdbuT/8nS
knFBjxS4OgkwA3d6Euotrygm3O1b5DBM/fo1T+OirTrfi76+pXsdFOfqMaFT5fo7
zzMMmIe4h460c3RJkCQmmh1Eyzlk4GDyDIYTWnG7a3s9jJVJn6WUTGaFCyPDzwuF
g79ROnEpl29ZbOa6D30JU8sYsI00m7yG2y8KZUqBAo7DQtF7gGUdbVOZiueZJ5OR
4FM1mYz6iJsO8sueuGufyoefjve37xvqytD4x+vgWotYXjSvxeHfwkSvK6kHyR6k
Rs4u63cbAggwHDfMMg7/+PsiHATGKuTDeJCoSAykc/hMJHRttysVVbxeMFqxu6Op
OHPOy38frUesZxVGYvKYTWkB9e2UErQGq2iELzoeYWQRA3zFnggmiW6AEb9SNskI
UIfpgnOfzfic3oF4V153DoPp9ZvhVlJCQMvo02kmXl8bpsm76J632IkgdShxduKH
YzRby4vxnkLQU9VUlinI+fSK6P5/jF8F2ped/bzD6VBAFxAJWxr6ws5IE2vbyGAr
icSXjHi2gAKqCRtIg1Jj6Yzsmujf2+ETDDv1owQtp431K7QM22csOiFkM6r59oDh
CR8XeN43MjBKp/Nd41BK1yQiKjZlAs5B3FUeA55XHLTCJppSz43QDVSImUi/Ovje
nYYNBF1qwDweDNnRc6byL3ELaT6kA8usAu4mPcf3ybGr0wPDiJ4Jla9bGeiSDSXk
eYZMCsvlMzWre1sU6E7Mr6xcIUKAPcYDPrRnd9PQ5eCnx/GSYaWMNtdx/3CJbdIh
90kglPgmH2yfpEyMh9EOwaRzieVTpXkA649PzZq7Fiutn7/oXQK/XOeHoRG0ipAt
3Y/aFuj0AcXWLPgbMZbD7UIR5+rzPByu9sbBCZiTYLXJlNCpqxWdjZQ0FKCj9nPp
PO40W/lE2m09SuLzfVuKrrGwVHDG9oixe1LO/nmmvgTwhPGMWQlkOHd+XdY5cfFK
dKKhfCwp87A3wlvVowOwQh9/PxJmplIzx4zNZnMyGgaI7NWQY4JBKGe8jvQKzUTB
Yi9fVMoiOAxBSvy1bXeYzlJBueK6ArODtwGiD5TnVN3KBsk/zn6lJA6RuQ45k5k0
snH6u7WXCSoXnYh1HyJDPqb7JRjI+pQjSRmThLUuz/Ch/DYBBGwD+MczFAbFqm0G
pRgOBTi4pg3/4icJ4BAPtEos8SGOY4rA6XaDlYhYNDZIPt4uBX3gwH1buuEQJO5J
MT3mjVAjfYhCQD7JoKI4S80segXXMjx/n7/rt3l6QadgtoedQT8/lXI9p9Eqo7+V
SmP/QB0zU3UTrmtWFNOrfyTuGKRaJT3PDaBH/vL/gx0m1tyPlJmgk+hmZwoXg49W
d6fDXsgtKp2n2gV33QqWdkMS6vqHxc5W95+fr4qC3gYzCY8hUqObENfNSfNZfkLE
bIYeuQVLNlhA3vlSq6aVpVJDaIoyNFCijakOcowO0kMIRPu43h4RH1w2orANsBuK
Q5FtNd1uOG0Fke5N4VKQf+gTBU3Vr7Nd/piQTsr1WUCzqqOVrhnMf3dOf/T+/TEE
FItqxiFDd4Wn4hsOv1pIDFNyNB9dN1272nnXN6S8VqjnXmvJVOdqwM/A3Zb9s3aZ
juqzqb7zHDSlhZSNakhWIk9mxL10u4ldEiVbI6G+LJGjaYxujU3lmKZvLC2MP97g
TFkr2zHm0Xul5pxCm3DZRotAAGgs9v3kz45vUBmtEhmv05ZKlcVNtBFMWutCgFe0
iG/0GY527NLHCmprtbG11Zlhn+doyyERMXes8OmDpBqmhs/Tom6u7Y1LbRO4qCg7
jsTfzQjWvuGA3wLFcIRN0cL85BLJH/uVvEaol3cWQ7vMOM1whQj801L75kfmYDrJ
xspdMgfjDga2k4p4KriTUusKruOjDv+teSZTJ0MIwYd5ibPgH6kenDxiYAEohL75
YHuRmLM/FkHlj5jPR845HbVOk9mJEgxZPKBldPkmvP08mOgG8U8U6RtzAa5yYTJZ
Eto8ixGQTiRydvjjD099o0kYV3cS2+EK4HAX9ZWLDQfXaljMa0zwQ4xkrvUxmbQ9
Z0cNjJ1dpZlM8DZDU6w8rP+T/sDF+qQLLYzk8Ux2xiuhJXouPUOoac78gkE9ERBH
Bg1kk3G47zmr5Vkuigd20eyKZ43Oxlu/Q6P860uFA7f6duzpI8vTv9HYmNSoJV1F
K1xmF409lPmB2hIJPETlryvd7p1mEYygXcBUCendjQvA6UIcV5x5bh5/fMxc8ZuM
wlP4A8TFwuejLAN2vQBl0y28sjUJ+AWjWb/hUM9Ld3yweAZ9UxGXwHGQKalgpPNM
cgokbL33nm03WYtXp+J+o1Jucc9i+1N1ae9UV18PqBZDy5a4pmhmPNJ21mOjna3b
HUhNRnBAJ+fNTbNbzrg8cLldv0dyh5AO0CHsk2RIXu4+GAhtEW9Gwe4xYFqUqakn
2aq8QEmbxFpqRV+Lcpaigx/EAtN6jBdSFERKkAMIYwbTkBdVengC7v8/VSU/RHmj
7PcjvYv/iq5ZbPMiH9Wv+ZvpAC7Tzk3SpTCdZVyuRLOQKI13/JCBulWioON4eXKK
vsIpSYhr+x+Bd3MPfs4R4EV7JOpmCZmf169j1R/OzgH4N4fdkAh8yTtqLNiqJayh
3gLwLEM8+JjK0bQYHGRVUMq73Iv2kgqCvdMPpyXW7WOUbpiklVPFeJ3iL1VIEQst
yyO6MJOXvL4RFu7ZS8XrvXmsngC5I41FaHrDSUbdcnLzSl0/h6v5dLRTpSFUvAaK
OVO8vc3upwn6qj4X4pf198GlcM1mK/5+sQ0nZ0THjAZR3I9NaM7OsfMFdHoIdVt4
SFa9dhFJlW9w4uuOyJCbFXYJyLHkoPvM2KlqIodr1xI16S0IWgH1eox4JrWc9+zi
hGOzj0yRChigoFM5oapOVnOOrFG2mL1q/zsq4vtUDeCahGZJ069DyUlbyyZ7JoOF
xdZNMnDLZDvBvN4YFyO+0S17dUzdsLIVSQ5jdusotW/7ZjWmHIRebZne0Oe28vOp
fjXdH7vWY6Nni31sw7b/xbZ1lzH0RpsvhZ5vOCTFSb3OkF3oVhHVo6KlxYRWWWj4
h/viwhoM1TJimfPBdC/4fCeTeP9WjF7FPOZXd1iXLz1mOTTHmOczTNnp3+ra71AM
SHkNUM66arkKEJ+IjjJdeadolCA3VBS7LZKrAT1MSJN0FnH6fpAMx2zoxFLE/1QZ
hW4PfEIVx0okwGkUXvDyuWs4TnzMlepaLJRobdq0b373aZyEb8m8nnTdm1yzqYwC
OLkRddrAUmqu6rt7ipJb2Hrzitmkd7xB/yzb4JjW+00U+Clf2D284R6HaB01qjLT
SN6LZUa6D7GuD3wq7a1cyewt2AmLMo0M4pT2nDQEt1c4wG2tVkZTj5hQzWpP3tVn
HquMXnoN6tnp0RbnI7dDpGQ2kAw4yWXw9BUeENZeR1RNMKkYgknT2n4lchfIY7t1
27o6YJgWWrdZZtqwECw0VkJPfkcv8ksH0U/sXTIdTZmuyGSk32PtNAFmrfozck7z
dEUVXi3e8a+vcmkLx6YiNSFrX+lM4US3L1HSO9AjUGPG8lreQ/16BrZx873qxRID
n4300P6KlbK/Jr0WQg7R2Xy8R6vPIpt/rIZqr/B9u3uVA1TyLuDiKTYDguL2cnwY
ewUyhfT5PuCPDCslRkgLBLZvVYaAE1EniHl1oxz77DjHmWUMFOuF4Y5ohIYwiyQu
5v/g5m0wPNK2KYaI61JsEWw6E/GEBR4GnxsABKfLPiKZglNosRCtALO2ynEkO1K2
xta2TRVw5sO7ncyi/hW9gXp3MPDLTzJj9P0z5v3bHstdRm+NLF8J8EW560eX/lSg
IvrhFmC3fd0BTNrrjw0cYnBInDb4ycdwpxnFWoey3D8BLn2Dycelt9HcQzH4E0Ua
2mh8rTk4NrmSyVW10/6YzQeb/NxvLe9PcleTSFnxz+Ba0LONyW86rv1PUhCCKY7C
Rlr7VqKemYeVDtDt4eWC8p5ExP3cetramclNNUHeVVHkU4+Pa8LVo7jMGsg5o5XQ
xjZdetTc0XYnhiSVGjDdDXO0dCWNg6UlK+cDYNekHlxGTfGRa8Vm1kphSH3PvhTv
QY6YjxuA1BnAKDQo0Idcjy1ONqffDwIyIOaGQbF/U0GPYcBxbixuQU5mWOGXzv7y
i8KiWsHOGu4fxDl8KyQSQoF0TGAQ/1CrS2XLyPYvsbJzPejyMhPQ4WZzI9N/TMy4
45canY1C8izR5HE47aBKB9AaYca9vpJukxbC3O19EO4Mc96OIeavWf+NPW3CbIG0
NRCcZZUID0WFevzCp3qhduuprn8r6JZunVTd2/7VkUxvF3FQOfdQhWaf+QsbVzsM
63SbW0UoORdeD9R+yjqGvGd9uUQYW6eVQ3qYDJCUMmBZ+Z/aQPY7IWf5DIzJRvd0
6EBH954cVBzTtTq4a6rEV3FFoMnavHB24RcVMhvkZwQqm5OBrihtoWA1sJ+97v1P
DXWbCShpK43JH7uXASUf+G0uTQMkpa5UucOx3waaR1wYWJXnQE+H/medQpaall2z
ZGYZPdHD8Gj7+GCQRmH3BPSd6zkkatIxpOKVOKUFNyo6P78IbTmTAYKkHyDVwq/u
gjoosh17XNlGhvqof3vA7mgEiV3o++HGPZvpOQ897xrZezHrRVkV5+ieu0NXx28D
JrVbNVSaRuXA68PeiY5de3Od8JbiYOk9J4vC9WsYQbmb8y9s+9deNxK8iEgOwm48
+QVK6OGQCIvvcnCTyemMv7Jq456fsEyI5Q7vSI1ebDz81n36y+F96GGXqKjP/7Ve
Tnd32xbpMR2IbCdsVrxYJKlcLmVGNCTCNlNzfW/KeA5fsAAYMlk+4IYdI6UumO0o
LbxgsB4kAvLS3jYMfVvx7oZPgc4t9LPP4nJnBH6Ydy1WZaQSl3psO+t8o2nI2nTG
24GzkFQOlyXJBWf69tlEuvBlEVqn3UdqAbS/+btb9tzrAXaMmBykn7wsAmK4cJNs
d2wO43QdCWSc7fCDjQNkAJw43vFtnthAzw360xy6e5JEFwrqLYPOo596wvcpwF9t
hQkaVlLw3Z+V6LDCGqLr43ZL0wcGkxg37sNO2HElXl8//pKdHsWRJ8msHMiTqZBO
sMkyBKNnjCj5edl3HNmL44AngRRDmlE4cpOcOjDkibYdPOVKXyfe+BuvU0+jX6rs
iwKir2/cvgvvBNolOh+ZOjWcTBRjtPgmQpLO51gRCx8aGF+zy5/T1Yb9MqaY/ia0
ZJPB+oOJikPbbQGS+z4AWSgUidcvxhWQrULX5MSYJP/ouQwPOrfFPdu9Ug5mVC4O
kFb3H69ScVnphZHAMukiDJvf7UNdZG5pZ4c9LSMRSJqszV+e9oquMh4AvyHjtmaS
Gscm1CybJlkpMWIhWqWOtBBCjkKMKYofQSYjJ0W5tnBAXusRuT7KJVei594scXVl
BTfzaLdwT0Mf8+kuvzosQXES/mtTvPxD6yz/SmWeRqLi2UBgkLC0JAy5dp0cnTQ+
ost/lUeuOiCUAB7Kms475QKRlVdF4tCNOIQ28dFoFJ2CToyuGHo7r1VQcFqEa12T
lc3Ol6S35m6F3d2bk1Clos6GR716HF8sGhKWYgQBiioD9IflBNIVa4DlSyMvOc2T
2ttSOLNZ7MJ41vKb5fcXMQfSVNq32l8K/sTBT2+GBS7XfY//7jHr2gxPAC9JYEYx
YH4pY2FyT8QfFGaldGHjPbbqx+ShOslw0QfAidxGPJAggKFqCL8rNXsSfHP/eDDa
PFHQQ84V4QvsSAEV7yCYMiIkh7wCyEW/9JTy47Mv9yhuvE2ieIK4gcOBhj7lU3CG
3zviiLlrE4NeZ++NEfSXnxHSCEFKAuna1NRY4fu41AnsB+Azw172Hix3vM8V0wsJ
gnQwQfk/XqaW89YdTKevTNCmc7tX8eWJ6rgr2kqGE0xEKXTeYmQhtnyMIeU4wrrh
0+Z7ZJX6BDAzTjKyhCELdBhgCP55jC5wSw0y9Y0UGP/mBE+prDumVTd5i9axcgNH
13+X6jY9o/eVXciUkyKLDJcR+44anu328PgacRlALcf470QwDrHQEd3C55ca1OFW
D6fK0nyaY+vpS7KcUjiRmxmoGbUo/vJ92xdfTI2gxnblJXY3obNVWxyRu/vu+Nak
z19ZedgDPoU4gPHYcov1AZVeDC5FRcD8GXngxL7NHebOwcP+Z2syT8gpSBsC+nzX
vbXbWsTbkKMJNrALskPDoKiY+ei+5ML10Slk7rDQG5ZC+UJegLzpnkbBhsnNaakZ
vbG0lJ07zu2h+7FDt6TfR3yTxVklO65KfAOUA+DQV2NfYK+0TbWiGZ1bkTTB1irN
krI7ClnLpdX7h8E4XBJ09a5p8j87jE2aJffMMj1ScelXM+uoeTNoDqbnOg077mBx
FaADdxTYFqBR6Sbg+l2j3vbuydxzhV0PWI4uReTT8SNB+9MJN4BwLwL2Hyq1WB7b
ocI0xuocxZqpe5h0d3FOIDHTsf83ERjHRpgSQVsrdQQecdn7enYyWug5u8dnulhQ
3pJotektrYiMElb5IpOUvO5dd2geGvHccBlPY5iLKKuXUU1sobixC/lcilpGSyRk
PPsTnd160vtee1STAYHwPP0O9+s6xLgMkAp6mTI0V3ip0oWhID+Ejri3BqXB6ZcH
MVtHLw5CaC6f5/p5+3beEivV3ix3bZzQ5bpZnfSlBL1JUZg3GiQ9dTGfG7sVrXSy
8FpR/NV+n6NvF6FxYdZrCa36EaO+G/DjTFh5Ej5dP+OVyCqhlBdPgtZT5dHQkwQv
ySdOuMilH0Q5ixQJJszl6wP97eJRM+R5WkIGUFv6oJ0IuY7cITE3esHf4QB0Q3/a
I0xByGXXtKgTgf029dNxJgCExVunEaMk21K1TrKtylhW4O6LG4TciDExo3hYWvlb
Uix9cBAuFNRPaH+dE3vkQE3/ZqCa+F8577GcSs7pRSoDaCVPJcBgtioeTWwS7WQ6
Lzh7kr3KAM+PR1X0mVgm5mcOTrVzSUn4NgfPT3PTrtd34gvE0SpfdDo6wt7GotCq
jE6yDpUaC9HLltxPAV+9FchSdg+/URQYp7mSh3eRsPeD/tZ4B7bgT1gLU0iigotK
VoyvutHCzA970hO5RKzNmlMi2WO0VbFdOdal6/GgYvDSrNkgXi3vaoHPGuzM/GP5
4v1JBqOexUv6tZm/wLS6kLfx3MK1oidFyMWG3QkekbfAOEIAKhzZGElMGF2/pLHs
8Z9SOdze6+T4hMw1iuWjRc9/gJmwH0DAZoGb7eisqD8zSYhjLkytI9jHKlAfLkMq
DmkkOHtJJsK9ouzD6uwXWQwOyicKm+sDluXO/UvCXaGnTDgz5hPqT38EWvA9VINE
IlV83nV/m+RO0qhs9+CrS/JAPlf7plTU4JvZCngh171NKc5eSlneZeufhzZLCL3K
zLLLj1H6OS/fQ34eitVVTDkeFF8/F+MERcrK9Xpx1enntvA0DyJQ2teBFqOKJs3P
+lasJvP3QlE0BywlSvQmM6ZkXg/SGzfYW08A6LOcLCMW0mPRVHD+IQJbnOYD92Oc
5EF2OKwnLHrPNFp2fghE1OlE3IhXdpGh4uHterQLVgbktA8DpoRzqcrNLgfIu5oj
tyNZ5ekLVhGSMH5QpsAH0nkhGrzSQZXTSyWscRWk59ie09O4pL3sOV4dD8KUbI+J
MaW5VSlPImOcaqsF7WSOp60gbg3aDqTrMTrK+m1PGqx06pQ8u/u4+ALBoRLipzmT
K65BQLR3yhSV5k6MxgFQtP2YSfc+D9eVKhA7UvE2UmCb6pmxURZu+EXb8Iz3LrEA
03Uv+LeDU5V6qwOQZavLsfu5cQtmxPWTNBKrHo/ZvQR2NAc2ziUNVNF8uZ5sd89f
AA6nw8w/BBzQ9wf+WRlUfdbEupxaU6qMGEUqPRGRA/D2i/UCjOZB5E12bOanTTxs
nrXMnTBDNEjuQa/5Y5gf0+tLA7e3yWio8f1i1POvYe//7ijJYkmn8XmApw18apl2
1H2cyortOLAtn+Vak99CHJnQK/E7HHueOat3BFXA6eopBcZKmx0o+x1z85L9sT9E
xiAIa/p2MwqbIUgZjcy48zXtT9IZk1yhBC5U/WsTuKqBgYAapjfN9/gsB1JmzVmu
bD4K9cJXSgVNonF4H/0m6k2Fvys492B0FUc4wA76B0cTecrdj+b757Nr/ATBUFld
SaQK4bftwIAr1D3rJmnp2ivSg/ShGP8jYesGgyBl4T9bN+Z35q1xz14f2k0Z8H5n
+kmmhhV27TXi4DWt+k3pqsJtWtyxdVS1+mWCCspnnlwRVhQQ/e7wKcABxV+kMreM
R3iqjEZ2riSe2c4MXzOwBNwQ00M8mXm8957bWunfKTyZEzC5Y7y7wWMSyhv9lPts
X56iA1CTxbCvt+HdWHpRhkl4Sf/fq3RbdhgCWO2gxgj4Xc2jUj+4/aANrKSO3IRS
eIK8aYapmq4gdJwhlCSm4gXSmxIXzOjlg/BTNF5Sz6UHuEzP6/cCpTB+tnGVIPmx
JEUtWG0qPRR1Aau5242uWV/GkofdZXZ9rDDRhulZK/JMmUdyjuEcxIgAa4CxUK57
9y8+Tz4ANpsvjzVvRZTUl5n8bCzFFjWClr/jKswA1BMjGSZEbi8A/YVU0dzLYyob
8KuUUuGUGKoTV50BRJJFtn2Va01MJ2Kb8NZ8u1uxRzx0F/s8XrOo62kgqsiKGrwI
j8psAyG6IxKAaBsHsjU7h6GlwRhOy6xotyrQ6JVm9SXvN4Dqx8j5KJkCdmGBE4vO
g5pqJHeIfEisC2eizxEowr44vcmoeL7RvDrJ9nKMwC2KiPtyImMiHQqaOMzgzVcQ
mXi20mJJOSJT3SbxIZRjGX9hzq2MCO1VUAWfMsHQQ9oYm3kdWC/YdnPYaeLPY/gh
uWcFQW8OSLuRYZ1CPHz5rIzi63bj/H56NvMM9UCtAts25UbLUbgdzwCBH6VSv6Tr
fB8dlBQvhNoMKCLwqPvCm864nyxvEGsXdF+F/PTPxcQjbectEU8x5y2+VgShrzrv
XsFZ2RSo8qtfbTVFzcr9bkf5Hd/l7APl1UCSAsRy3wDk6lhMuAF0tuJ+DXGLFOm0
hN65ycycSXj6QJXEhA1Y13UCtMyOkSYYMjEKf6RNrRETSsr5+VYpR5rfoVD+wm2v
adC1PxxNugTa0Q72z6L119M8M8x4efhUlov0toK4aXJKu8mdQ3QD8QIKJVpFi9J/
sPuIdoMcx+JhrujwwIrBPn1jgiOzeAWHBvlb9j9gho0XIeFFF3nUB3Rg89+nPHql
THjmzndhf4rl+zaiaJdRXoRRXgtCbt9V9gso6ltDe0CHq2jqSNvQ6PC0AizRZBhl
MG89tRrUbjqwgJt8R04DQSG/CCTcVMOfrg3s5p1bRewxFIjuM0RptlaIOLs6nnnr
6wpFPr9okIaBUjvZRpdmknxI6W5JrjZdUsc588LpjQ8/bMqMPz/gBCxrcle2WUIV
SGrjqpYDJqPxlfxUngsrvKQx8PIfmbXY6gUZgOPmQFZvklxpuuDNavzgKzLJ+S+U
0ip6uig3iuYpe2/EWUQWKIWGQZj7aIrNNl8ZGOZWrofPb9d1YStbHCs/bk3Yi2o8
LAjXwinb3qhSbkWejnAUvFYFc/+C97iDMp9oD+WlQYPmQXAmVyEozzvZU30WmqMO
5i84jT78oqUxefqubOmQq68aS7EPyWL/z3RT+0LtIND1Md6wW2ZqegRMJ6PYM6RK
lOsg9YoMQy0nNsrcW6iOP8kQrzH6r63VWwNSHz43aU2ed+I8ykomp07FIlb3GL7E
m/Mu1XnrP+khhuDQiYJR0asUFEln1La3Rkqq0nMi1b+glp0v/eEChFBvTHJC1Vwr
ilCV0R1p/eidikxxx4JBGAVvxvtkATrbgVQCC5YfD99EJzdM6xFnplEIvGQ+CO2J
/6nwz0nvlFsQOrJYCKjtkedEMTaYR825mg27QzDreHxRe68eaa1SZ9Vl2WfSh1ij
+/zwHC2OvXm2G4sr7KmuqiNDcn+cuk6I4AkbvMpnIaVIW+ED7dQ5boydLYC9Vl93
UK87oBx6bYDHeKbwPXUTNAnKVzbtgzL6JVPy0ANeSMRj/9NBZPbZ+FefRA8C54BG
72vv6rahZvjijArlAKtWZ18Ulm7NQGv0IDI51rSTcBCz/ILailzm4UsvlH5ViyFz
IYkB/B/zb5hRu/eJFQOQ/1gFFb77diey+/oYMABHB6Cieit/BPqDMctjzSHV62Q/
KTv0jJ3FbHmdv/F8SaUukK+0q2iMjzZp3LiEk4H0ILrIFwwR0rxGzKU/g5x2PwzZ
3554pJ+uZNuRKW7++287ssJT/JpE2j4qLzJD9ufpFHXa350BrL2ZJY8j164PAMtI
7bJLWXNTu0YQdWNUZAmYctvgVmsNNhQV71UKMX5diodpvw5dBIPaKdZbYC0ES4JD
J7iPcJ+C1iQpV87QAtEfpX+C9TICouAm5/I3g9AtSZGl292zo3yEqdEah036Eg+2
FCCohOk+f23lRbB2sPZt3oSfQT16PlJbv5NDuFZawVBwUGtfQ+G/KxmhtEK0dokY
Lu1IsTmDnWlYUZ69JNNrC4ImHi5zEIaC04D994yH6FtMjfnvntXcd+PvvzgS0s6k
IY9LUjbCGaB8r0wKXCM0105+nrY/my09Go6u+EZtZBq0oKse5w9U2ZE5y2E9UA9V
+2Ij5iDL4eQJmE6pq8o6e9eyLurCdrKb/EdebWxNO4+Md30ywIgWK1m23dcrxYC4
vcInUOVd2F238EtG5UBdDpXfsfWfDKhHHGFeFUl3jmV8Yxgts1RELWwRaiDNYOgD
R6Xryf9QVU9TDEoY6nZRdokT6j9GiAZtBwlsCZAf2xLbqYDZKSlQkoESkrO3sRIv
ONM4udfR9/SoPmM50xZlgm2SyYEHzOlrLk9YSVEuKaB4kEFQ5x8j2LljlhSTX8OY
uNf+PlKW82GnLrxaryS1/kR/kjhc6R6DUSo6n2gWATxHBQATl/PvwwuTNkGrO9+i
MtTo78S8m82gnIuSEl3LkVQKE+XW4aYNWGYndR0cw2XKjsKui18p2K4ouL9j7yxf
+3WZjEXhkHkYGXA+ss3Y+WTXHUNUAdthT5Z0UrxjuNzY3BTq/EYu8VuxchZwh0Mb
yzNnCk1BvahnfwOp/8jTW5lbr36n0I8UtOuXJDQpaMzJQ/hJqGtH91JXa5XuW2oG
VSHqaBSJwayzoQsVm4ZM4Ue3JLamr5eMZ9LtRKiEea5SjD/bS7CXtbTxtRvk1+ld
FXG1DK3rAPe+166FSZt54dNh3GX/km/mcMXEL13d2xqjqBS9vgrxoirQ1x5Vx0er
QoiH1uYa5W+EKiietYNXvGk2rpJrop0TAdVWGSNe7915yxbLv0HK6CZKcnphBJu/
ZC47rQ9/gXkyoV5q0eTfLGkf+vSo7IAJpW7f3gkd1Ogo/8UpC3JpExztBf6AxqYs
1P7M8JbOUe7gg/RaaTOsYdfuv3qr9r3rak+4iOvLXNB16dz05blYVJs5YoAEDhFT
njArwZDSMctKQrlwPOGq3/ONE1bJ72y4S4wicWLm7LwRYVqhvaTrCpcZPqpPZQX8
We41fuwwjeGEEzaG/PH/LuvawyJ9hm377LAWmIv87M5pMMBIKv/DEpBu/HZqE6Qo
8utpV+jxn7zrnshRsUys6q81M6Y1XEJzZ4s2UJmGNcJAkA3zzvh2948q9NsA3qoC
ZvawQGE/bYH6VBwMvjfDmsEACr2idO8u9FBJpGbRUdlXvv0X/MtxdnIfYkMwBnuC
yqlGdQapIza0kQiCqrEQWmzq4vQCxCicYwWmy1JZw/LR3KIaZhKl/EzpjlqFswb/
f74vymai/1LozYYrFlkCTr5ZJG1j3qa8+H5AnhsFbws6+GtiuFwZy/CA+rw+j+Sz
Mevd8p/NRZb7nR4Cki7sXIZWrSjT9qSUATjr5fU/7hMTaMTanIj+GlYHLfdzM6GF
caT/x1xwg9lyQaA0OBOaW9p5oqiDAlz/ntDBUlPpH5DJd5/2gtRbUcmoMDiG2EsY
6crs1083Gy71ucm7UwtHSJYNVYeLELk/rD4JAtiHpPYNZXgtmwtiDAIs1aAmV5cG
RwTOo+RqJ+S0jjT16CNk9NnMlR4y2dEp4XeKf5CnLGdMnGH/ffLmumwI4fmaIvQ0
uHuN1lBULkqWJERRkETB2DFLVnSUd0tm/dn+wV9x71zQzRi6aVKw22yyV4r7XMuM
EML0AItIPBJdEcnZlABnWC9A8tkTORtNRULQlJ4pIJ/6LT5BpuxkdTLel1BToouk
sLVxd4PClHJn5qYb8H0q1kS/GVftXlVymb1Khw8ouBkGB9IrBKlWsbfW2ITz2EJ9
fmcSE/FOKEXQ7xs6lfEax+mLFacE6i1geA+TMn7lgIwofF3jYFcygw6zqkff9OiA
ry8ZesfZKoWNsh3k7aH1EmjiKf6kTJCnEx3kxjEFM5tyR7fdtPRmiBJ09RD2ulfT
BIlgwdECPnBM/UHEu0Zpuyl87DPWy4cey20je7j1+Zf+PlxcPY/d8gWXbaCTkCyJ
UJd7H8dL4SeSPOjSihXujm4ykUe4cjUdAPIbspCdMJeCRbtJV5HS8p0Enqrpra9m
LkfC24XweuHPEkLrXKO7xT2tqcfDjc7qiRHhiG/chEIyWYM2zkx78ReBVZNDeq6Z
SMRsapEpW9qLFBeh4fKOanpgVCn6Nm9MAb9rRL1Zc4SjE/a69IbRwj4uMxTIx8il
sBV1dyHJkoVsKmtFEYUzwcZnw/6un7NGmG8ylroVrDTygQaKWpXh7mfZrJZfxWf2
sR/Pn55IDcXKlnnM248z+gNC79V1oFhgPB2BgkT2yKszpss8fDerLOd31h3vW6TP
1eDXolOVkQ+psncACUiFL6AZPm3bnCyu7W+ClFq4Cu1X22RAk6Ux6gxxJ0PzYYqG
FJxQ9ucIqUk87LLoGF271sR0mFXo959KMqPcs4eq8o9h2NXHK6fmGGBwWJTM9N2A
NvkdDHIbh8v5t4jvHn0NqZuXL5Or+85R8RrKPbAwnCz26C8PaBWSAXIlg/aPaWOa
9ta/p2vxaGfnx6IZoGHVoJQp3gAIw2cn/MK6V6v5ga0reL6qVpUt55AgTXjFl9zQ
ernIIwTMnSZzTjcksrwfMr2vHldY6oTaGlyFzMQjRLk/h9vC89uEZM574J7bO76A
wNFem7hvIE2dIwvBrIBphbuoSxUNzce005GMaDT8q9XjneTWQozZ5TR3kFLdWNsQ
TKmSEOK5oSRDydcpwNf/Mc0+8A+ipojFj0axc3/Hqj0XsqAZhf/2zGi5JTtjb8Wl
OZBMGR/95h1N0YmepCHK5bKCoJCJgMDryHhjTYPC/2poaMlz1YbZ/ECFX4mCpj4A
4g9YCNQJPiMuANiVPTGHcw3LFKfAvIroW5EyugVJMnkiMAk+++I3rJqLvwfuNpSQ
vQK6LrGFhBcd0txJs6xoUO4GfeLtvV3CpKdv8mLRhrxiGkWT1NefnNJKZXzvZWrv
KfHydLhB6MMSvLVpbusYI0ftrJMwynggL/3D485oeYZ7SCZ4cyylJj3chPDdZCDQ
6ddcn391PUTTK5jCI6k7krP3D96epGItx9KGOrw3hyK6ufpKDtPl7iRl1Cot9HlF
1ZetsSQWq2Cr/4WdpQ/0V/hJEqLJoJ9anm1Dvg9EA6dKDlpdGFWgj+KXMVGin2lS
lp77rdt0TLzmDQutiKwcBhmj6LmrVLyRBCdhLFXYcRCOO2bRw57saxLVkE0/rcxt
dwf0Q1hQwhAUUKwfU7TxZrvkQ5TdlluzyIdZUlLuw3etZv+/KtDbwTrR74H7dTtg
HdFYtL11ctIJWRDw76K+OQCKCDUaF1N6s8fyzxhQ48feOVZgp96fHIzdHTp35rG8
JWZa2oMi9MVMRZxRTWNCArWL+GCjglui3nI50OMfW0FRLNAWvvE01JntKNHDgky8
Af2ObXECA67rDsIvyOTq2ivJXQS38LCq/Yi74DMPun5yqDQ6jEN3pvdaA4wCE5QY
4aXQFhWMsQ4j9Gfac29CyWCKZdxwOXALueil+gc79n2dshKak5Sx8mRd9E2kMq1b
B27PXISntBnrgMmJIjRTJMRjNlDo9pfYpUo4jGs2ZoK4tjA46QaRYWKADy8IEk5F
jBdPphWcyywMfaq2lisLbsW38rTfb7PQ9l9Y/NRl6bPHHhlYeF4uAq+FoeN6GZTZ
5fj5SBinnK8NJbCGR88WSwPH68fgnxBC+y6RFTJCm4HQKjtKDKzMBGMNcnsAOPOj
Y7zPWGcBct+t053/1J7gNaAoHz3mgER96VVfkTFWMmUiNgM1JwpSEI3ve11q7+t9
+tdpq2gqdX4WkSPT7fD5+n9iiq3JYyBBByKQ76rVcdU6BRe/RO6Ih4nxkbSROjhn
Qqsc1mzpzERM0hS74VZlaxIEq597qKuV+euEVkHGGg1RcvszP/Jvc4TLCFuZyN5a
i/dV/yA7zDmuVHZODplszB4HyA4ba9lS7z1vUyj5k6G5rG58N9J3qx+CPAOpK/7R
AnyFfZ4daFgOq+BbkZZIU9LfaKu5xiwEErBRZSZ3cTy7w6YGKtoYA2X+PoT57rsZ
MfYdXpRNCdpyV3Ozwx6HsAh8pwJJG3y4Ksjci8uncfytUV57vA3BhiE5dGpqjT0f
4VkjYsedxlFMVmZCyD/1wz06PLzf5fr+g0eCMmhBba5rw1zbY1MrfZ9Fcp8nBMYi
tJEv7YNUoADM+GhXs/kDypFZfNFSRhGT1/VCyx7BRI7I+op3b0LUPqF2bkRdEMNe
B/jDbbI8rTOdrxBLelIwZHTs9T6urXlAGTjWh+nSIwcnuD28pY9ejOB3KrylqXZ0
rSTARlKmWRL9hQ4rffqpD9jGLlqwaJjgzKpn3MAollGCLohL8woymNEOEl7rw6r9
f45jXneM8fWXtCrCBayyI966FN1iQNW3dzLTaFcLURsnawMhQO0pMCaaxSsoGkdv
khwlAAWAw3Pmj4ILOJd23Bt/IMWx0sjJrrRkkk9081LRfPIDt6Bk9tloQxXtJcId
4GgUl8xvkLDhX2GgPUz9uqYlWpO6qdQYLgG27Tz6TY6jXGNl3Z77FOj61EnCpdVR
FAPo/mmRQ7NNXRYiBj9gdTGfZLtU7FnG2yCQ9vzlHLK5bg6RMn/WxS83zLntV7dw
IFQ2LVr4Oaaj3KkFcjVTN4iUPJv1bGcNQmYVFIfYvHtdZ0Kv9dMANz8XNSMhywq9
bpq2gc3/v7B1olfPreXN9JRKWVuZ1P+NmoQwjBTsmic6xOgicH8y0zLhMYRe0quh
M00dO3plFWljpUWJTW9KGzAtHA5ZS/g7phlfv9JOyhpwaBe3CkFH6T4QyUOZTBVr
CItIC/uP/qpPcZAKtarZE/BIn4S9zxUV2q59nKH+0GIcVtSFw2xhCyP2yuzks6Q4
VUN2j2EvzocYU4oa4lU1vhscIAA5u7Dys0EHNLhDl3vyLgJuFOCm8Ck/Qg/mELMf
TTD/kKEbETht+UGIAdIBis0IgLOFoNoJr+tpfgXPn5IQ9UujbRj9jsXs6/UABhk0
DDhSxrStuWD0zhP95Shm3BnjxYzPV2kggHI/J0GibtotVDWuMsPJUP8ELj4QX7zY
kms53Hnq3ukOrzRwZQj1f8Ghs8k06kZRBFuOqWYZEcTYUYhAFdnVbWK8jlP8UTR5
sOBHkf5lcJSHFQ+hqdXU9T5KAf4nf8W5wdUX4bFIF1/UG1c/Sfk8YaKpRhpvkPlA
hsDocAwJS3IctLXwY0+29pZMzxNZZgnXOpVpp1MWQ3uiFPWRWkSzeHt4fxE+dPee
27CB9UU9NUw/9OyMF0Oj8U6aw1G09k+JiJPYBStRvjemM66daktenbGvZDauTQ5V
y1YIMC7bsi1czMLQxwYxzeASplIgYIbCaXXSmrEmwBkLdJLLH09mEJtgTACyg0AF
bz5CXtHf1TpsfhyOkg666Xaw6Zy8sVO5h5Tg+GNtGoUkg4y68fb6QMc3trTUfE3I
x5E4zmZQOgQ9415Edu7xYJ1AanmBTbk0d8mQ6upjESfU5IT3BIIhx9wr+8euC7aX
hgrV7P1sVPznqoXZjhA55vj4sajZk+Pc5Abb2+/yQTPBgx9x8qcnpv+kj1edwTAt
HfNSJOnXwLAdNxJi0H5Vr2odZAV3+tBFmgwYFVGUh+G9m2AUFDPkUaF8ZFnlRn9V
odrSoTjlyzGv+5BxXA1KkJy+CPIoBrWEkne1Sl6DsuPSLbsenMEZrj5CQgNQKGjy
5KxIYXc1eTtC1mpJx6ih/67P/3xrqc98nUkcCcXIlD9ZhSlB1psxvdF7sI1KWqhr
SOMR3AvgRBy26SCToR3iMWGgtvuYh2AZQan573+F1cgg+BkQyONMh3fr8bSRTGGv
ONWtqOvF0COBPDA6lMls8CcDnr01waomzpyXlpdq+SUbN4pCgO8WA/h8rer/K/p8
OAIqjQQeDr2P4rS317oYAUKa+QW7My5zlRzKN0k+FPPsCqvqZAc8JinEXdvRDBFN
3mRgwU7qzL+Y556JtK6jFal/2R6MvMDAys5v4dbhakoha0kHh/AdLAVBTcJ09YZh
dhqPDZ7pUHZ0D7IdI+KF/nANtuVdnq9r44R2UZQyWrBSmHnMcayn4xlZyvjqEje4
hOVY6yDEPqm5y6QQsr2YLKLTWy3pJJa/SXZubpzwoy9d6koteChCymO6lZDYUUQm
etCyJNElaNj7IP4rZHQayapdTwbsr6lvDJ7LZgBv3xQv/I6mTK8ZNY/EUTOuPYNY
G8HntzFwqpwZH1MM8TC0dUcvxORj0PlFxFEXJQzXk69xLvuBXDlhDcJdUncqwT6k
apxtkh/9sQetIgItnhf/8+ODVyH18Q9Hu3l/hoWmPoXdF/A97NJmseMeeZtYeCgh
EetLPoSY3m0PfWPePnsVmDq/AgT5oitt+SQI/zImmbxIV+c6mu/xV4Bv+xxEnS+0
aMKw+bh+c+A1xjIC02Slp8PgWH1E2F7rgauNHu8ynwpLBZxcqO4ms7UFQL7bfjRz
D8GQalNOZ+67U6ScPEDAD8g3DCc8JkDjtsMIRgX9+6dRfTHNypH5jcirao/p6jhB
IBpUK2CqiTP8hDtV8gqxC4iN/tYh1XxWdEK69sj6yw4yAR76Z3OM5hLdlzJ4/35j
/pMVPclML/z4LkJBoN0MomQhZGqHpElmDjawVss4VONFGQCsC96s4Eb3QYIW7XrO
zxQKGuaNCAzMDjdwTCujrT2xfHi0BeIXpci1SEemyhGpYoIvYL/i2TxFeENC9h7s
tixF51s19ysUveMh/Y142yolje6VFB42ZSsV7q2rgBWUDg2CJfDFRLPJ98dKYktT
Eh4Boen77Nxft5M4h07XxqJNRNmwQVO0cI8ReVwFIdPadhZPoKLcBwRxEWvzpvBx
bWdMyQaHPaWEc+uokeS1vfJVX5uAIvXuNngJ33Thx4lDNsA0Ne6uUEkmAl0JM4Gp
T8DFJQopTI3FCCIIKeohF5opxMGKleb+SLNlvz+Dgv9IE6xKdjLi8wHOYe0SvbS2
IcqTQxGmPak3qIxGkL7iMp/12sbPatNc5CPjemUTzrBIuQGqzqGeAg1iahbFI1MQ
mmYoA+bdPiPOcCkDd8BgrwQLJCCApAiMBwVF8BXTYQWmBzklcv5/NGxxLu4GhqDT
Bg5+wkn49vwUcsewHhYl+o/e8CWEXSISQPLvqxtuML+i9++bZPWOQX838Yl3gzOV
K58uIEh+O+j4DLquiFSRPM+TDak6jm0qNLIiqOwkRz2lbLtKC/ynf5xSaLn174tn
GjxLa8qyncWa3PneZBqotqUd0to2krYSRiAqNgtQlJANzZa3ROXJIt92JUV/ODgK
jj4+3yvQCeiUUKVd9gsv9ZX4+4f+5xtjXY4eqt0tr7gS/97zbddSuPN/1iiMlmBa
/LEUYJRzhFd2Xe4ipNdqRRssRF6Mlzo5IJBNPKDikbfR7cazxaK9JfGcOmbObASr
SKDnrgXk2sunbqfk8lNeiMJsgcBvpoW2J1r6T7nD9tNfvD8CJtlQi7M3iw0aTZm5
s7upvGb5hOZMytv+sz7Un2Yfnuj6mGzLhFNrTIStFnoaO9z6kzIQMotSnGQeEHkE
a9OBuLosi60rZeZOoHWy9UAU15Htm4DxxTeWxoI9HTr1YCsxq7KaIwsxYZY1Zvaf
/SotvKpGVLw7aUoG9h5xC0ADQW8GQ++TaDqV7bryBkw9ncb3J6TtYE/Tr8wKfCoC
8TlUvmAqoCnQyiBppp198Sqn+d6sGX4HYkTFkBM8nXSWjfJ1UnJohBHbVkyVrJEE
pyX4Jpfzcy5Jz4GxEZPUnIndyXWR12NRUutsyEZrGOsW19zCQiZ6lBsXWjWMT4vc
k+yqQCGqCL1nKc8TYfnfo0EE0u7EYz5+qt6H84i1goZ35KEsKmUJJgIh8PX4cpyD
pBMiA30SRT3/SY/OrSrHqMhXCBkCdnMfBg5HfwDyyCHb+2bUwWhhCZ8IKkQAezpw
Sru0quN+0I0WUvnZ/9AtfKD4aDDhmuuKvmI0zKTs4HC072aTmfwdkVPcCOzUT/lG
5sEnRT9dg95Ij3vGtjKUZExyVTy+9IVV1mUH/bvee3FZ+yfFoREsVVVI71CKnJfo
x8F52OJagAkVyIbSJvevYAgKw17KaQ/nE1AhOw8Vo71aVVaKYDZcbB9thLg931p+
Sl2N+hZZtZgAnNzZK4VFDYgxg02lZ0QMYLS20xcnFQAW51038CGNh6CYCSQJgGkQ
qp1fqera+kt0KgfX67ZrifD0hWhoSzsImfhqip9jgT3GuCeJehySeVXuuoMpt7DE
97xtt55CmOYV79Fmbj+ThkjcXI5pfzLUBh69s98B3UvMXoR215J8tEDsOehibaHe
v/9vKd/VeueJTPD5j2eP1b+cLW6R/ySWtWdDIk10rO+CmVzZuFQnN7JGLJfswkOs
ZGisaVCRChco9lAV7GK0PUl1ftXIB8ymFh9IaBMklg5Yn1ArrO4WhDtx6Vu7INMX
PBuU5XYmCHrTsvegqPy8606FFoTmYqFhWd1mquYdrKDOmPrWqNmtriTmsMPV1a2Q
R4yqKFnLY47cuY3sbr8K1x2lNVDsWIIH6mBQdJLLQ/UlxTUgmboM5D8wo3ZCGYoD
J3rXirbH6EYWqzVF0yOThVJEmeLxETonmcF/FQTSSJrEZE+8bYvZpRDmc5fbu2hF
Nq1sQziJlLrm5xm0hqN8qG+60K2bhx8Nc+XDjUPuwzp2YiUup56WSlV60tfRxmn1
I417I5Xb+7J3k2uT8eDphY3AkaY8utL41GP9GYr9xR5WwWKbwnfAtT93rIJv1kAg
zUXKlA+Al03bstMoFOpc3m+DjQAN0dLtuc6q9KyrwQ+MA8SwHK6wwlyBmk9TIyTo
9IPr6IPP5eJbqjqPjs7jSn0HRX4WIqPyzyIVA5I/cAF9ImprmXUQlHiNYJlfrVuf
EJuo59OOi/UcltI4UoP0T+n/3ElZvl/XuUu6r/l0qVCRHjzPyhgp1GjQLPmV3nHw
FUu4p8Rybqj5EMOVVmQIHhTH0tYMbW91mgIcbS3BarXkg5wlfjznX7Y0mjqN+I+V
Yo9TrLxeVQxGXfAcwP6gw/G7CwfhcvwTbzYZItZ9ej6kerlODmzYWF9PuOG+5k6S
4ovHJSonkpiZNLej4AhYkyQVQO8ur5alDD5SeeRwdHzJ7ewpqYUGZKpqk6St3njt
SBUaLCL0E33+quim4bxOM0ncauAmpNXxSGmzwk1bZDAAvFUmK6KWxevDdpv9TpmB
APCor1o0IZry6ukZnjkoCx6Jrbg00inw4UT71qGBaTEduuSnaV/7s7PUSoHO28DN
vHRLHoqpS0JiTktIjMBC+eATMQGMBut1Gz7CV39aqSnELIPRQDmjJWe+pM289y7W
u5QDlzgq8dpbVcjXnuDWGOxRy8fm0l50d2/OIQ/YCOX2EWl/oN7DKjOHWcR36Qas
qIjtqW7aYXfl9ZjsC7MIPiB+702o+HK1+3ONM7L3Mo64a0PCLCFBz+9ZSBaKcuPk
P8fUtEXRHTQBTSNz6Q6Ls1B+p7qmndOyQ56U7bwXWsIugyCccl6CFAZR1TENaQNB
OCaVkBd62kr/vrDuf6L6s/KvXnAT92cGl2VDKjFZoACmm5nBDfgOnJOQmcLoXneR
+5Sck8Xx8C7okKXbPg8SImmlEkUoSHebbt6eJkMb1BU4UTr/koKxsG53LoniiCgX
r8CTa836yA26APIXpOpNH/fu/3wSUXPEV5T+o1aic8AkbgaIXjXDYKYIEoYDJ8aM
QRx23Sx5VloKpF2kUFhug8DM/EoLmRTzKyFFWQ5wvy86qXo+62o1iYR+SOpQPune
YHQJkOWWxUe9BJyjtgzQoHSNrKrSs1iXqVIr+BW41gfMD4ObWOAE4Bzl9Sd9bvuW
wd6c2hBcj4276FEXNx6V9HVrsqOy3P1V9oYgl8kjV4txGQg9GI93irX70B8DeGEb
8ku2zgb3+CaFOSpmkPBRSWX3MlAGb9pP/ZIJ0xFpieRyFwO27FJthMaZfj0y2rWZ
7kS0rJ47K41BlmCeRNEDJL8E0BSka3PhW7v7xzxvPj1bBUwLeJaqe69+ExC7uwfv
mpMKKz0XqNBcl5woKahbOPd++BxZc52IwupETw+8Q+U73ttMex6RlUNeRATcgXZ2
+KBj28ln/b0G8y7MtyGfg3ByGIJoqv5W6RkTOABBmFsM+nWjhFAGq3bWtKj3CUmS
RNXi2aPzHMKKDu748AwveN7mrysSHA7R28mFGX9i31wNgLi8zgrbOttCSwU514vn
tTREnTzSJz+AuYMz1y3i8FU0o2NK55HZV7CIJ8+SAbjWpfOmnE5H0CB+DJbuaKgS
wr2vPeYzfsX+Ce4acDHNbnzewxQ3gACG/jEEMAOHwKh+cJ0XXmHhxj86l+o5v9sG
8a38UFRzuAvq9JGnShqinUZuE0jrD1qnYbbhQ+22LH+rsBwgGvlPTWKLiCZM0Qwu
uqk7Ogy/VxhONlYo1KTBARKb9RT+cpdOa+DBnST9zzSduqq8GytH0bZrh3obowPl
r8hcV/zUg4zTL1ysawPcLGHSTZhS09bgyx1NXznQTqjUFgbA79MGBwuB6a7foAGf
nNz+EEI9suPwaOnj9ISJ9/lnnuKnUYJsPwb1k5sA3qpDGkDmUwPTnvuBagXEXahr
R5aFEuqvtNZL1RbDzl5U28fhdSoFuQcBC31qdvdncVYaJGUv5g6C3DuUNReWm/jf
qLZWXs0w39mt93d4uAG/2kyd6T3FWXX8O1j5+RrcCxDOm5BbbF0flCOi3SoC8Us3
7ip5aDjUxLv08wQMjVGXlk8dVRylFh/1B1gvOraFm443mDuQDowgJIldaSyoLmEv
fHjXOv1qqUCUOHQt/WwQQ0pT1VvbtOh+D4E3fWjYOIldKie5aOFZLUjUdA97TUTr
8briDlxTgUGg8g3p7VNTA7Qvg/uWAnJm807g1Xe9/zuLzZiOOD0KaFRtXY9uQhIH
dJdOfRm7JrPW4Q41ZVRkuaSHdzKaS6WKO/zdkuS5iBS3/Re2tVV0lXPOk6S3VG1t
vNpOZ8WiG6ptaST/lYesULn22vGNmjL67Quh7XS61HzZQv0EeDpjVUISneal0ppA
IHtznTTH4FTGsKIAlo8j3TQQO+vSzyL3i9YB7hacEBesOJGUHBmvi7oBrAzzQlgs
jbkAcGYbEfPIDkia3huIrPcMuek7b2NxZmacqntR3Ym25nXqxRZaRMaZsTSCoDeA
mAs1VqAPCXqqiADIJUGB/0LuQ8qoAkvsbIaO3hb6GU/DucT2aplUyLYhgqCNQRoe
paMGJDiE6NsgLBevm675S8kJyRMxmU8eSaPJ20uBVayysre4UqB+s1M/loT6OxAT
ClYJvkuLuiJVsF7IufDl4kFR1UFBN5TRARHoj4jpYc28klAh56TksnMczUFTYTwr
cFbCCmK/lFnEOjghmEK6nqUP1DXrka76bWDz6YT+V+lWpItndQFwVOx/cFI++58m
7E5FXKh4ip6w/ITHgBeL9ECOhrZhZ9wbMSckpvTLwDoLE1yduIoVTLWSwKHFUqar
4iHB5AdYbnVp0WCMkvj32C+6zib8pgduoTxb2ePH3N9V2ZppuNr3QBgZ+fR17dD2
TS235YYwilYTRzddwqYd6+rIabTwIrO+HBp5s2dkxh3SD4k2SW+zmsLONv9AgBa5
uyjuSfKHsP/9XdHinaPlcu5ticUuvcxi0QhO7xzE9AKJOnUOMxRu7IaGtDHpXaWZ
2XIzMpf0XBbgARtjOFxNxCGAGk7kqRrKpNZ6NPREv7KsvERUJzFjlJyhIz1IGSkR
meEo/oqmD6H3tRdxc8MB147+ltZgN4bY3ThBbNYOn6WEPSeXj+kKOD39ewZGqykv
iQL/S5uCDtbbYcYMFFcb5fAzBz09JSNl0en52tzlfVmkKhVPo6lWVJ5CIAPmeSXE
+YgtjWILhWxM05bAbqcDuq/lkCkmb35RH8ELORJ0dCpFBRVeBYDqOhdsf6J394We
cvrMiRbifcQe43ebSDeF5Z8nwzCkytIoyECuMNoZT0zXz7rDjP3YM8p4FBbApaIe
dM0Lo0FFHo3djOb9p4wd+9RmLTtiIPAjYBmQD544v96HMBNgkTI1IVKcSpUdQAtD
6wSz1WzayzrSEr+1IRJXh4mYiDAgl1JSY8AHDyZsx4SWik9fTgwtbNVjJ6Y6wV7i
xaoIBlLs+9yWjP557c60esJVhkCbEwVIr4sel93fHMHf1T88/w/WXZcLqM/1PKqp
VeHYexUHPxYeeQIfyUvN/RhVfxOLhURCBIcQyJsBrK7RiPDOArJY0vFdXavbT5I2
tvWa+25WFuld1mYEOGYIvUFkt3/UTHI21imA2piLNqXyOVE1FN6/ifkoO8Jhiwkp
Fnx7zTo6sY2ayWagR0L4gv72Rs1ZNcMDe6Nu4P2xsTpyAW+ovPU1/8ORnjo+Tfoj
LPyZINCTPJ4SoPg4wHCTfHA6VflHJgk5CBgPq/LcjsIsbmr58JiiveNJKdVqvDvv
yEeXaI6/bW0bOPXsxdSY0pxzK0rL/7jatg9GWP2oBeQp2n9E1ZtT7K+seGeZ0TIz
usgaIng55PWDDuxnFA9zwPrw0Lz1GApF4PLa/hIVLf8MMJ1yVkpCRW3JcbJGBT+M
GbP9yKN3aow96x3pkhtGKq/8/xsLbiQxJ6U9jhVkbIicDBMOoIMdvSAKaZUj62qz
IdSsktCmZtIr/jA2Vh1Y0/Th26suIy7+vIE742EJBHxwTymoilMTRjNMZsLOSYt/
1+Zv79cSu3q5Nf0uxloBhNENLlFA15xO5Gipimg2pufAMOzlP5FwAAa/n0tPKKo+
B1ArIUI0633aDkXMRg9frgipHrbKiEd9AeGR/EQb/aspHEKgnzQLeIze3VKNmGLH
U9+yFwfbbJcIO4fEKpQLkErq+ZnyJRMHZZil3jZx6FG597rW/Rr+mQVbTbOlBa82
u6TadcGbQ+zR/GwPThJOOyqsmTRXOjRrsAYM/QsHUupWht98bADV5MDiQHelf7ay
jIyCPKA8ANtpt8qPWecV1ndZQCG3T3tIt3qOWnjH0Ki5QCLB1oETp4ufZ/W4cO9X
hcToFSd5ORkIcov3TOcmze7xL9zSlJbs8XyDz7xiOOdnqbzq4LOkmsRBNtiGPCPU
O5k5WLgaoRxoUu0QDKqGl/KOv4SBriW5KwMm+whmwN1HSdh7Bq030RRpPv8cpHCG
nsBQL2nwo+ylWoHcSEAfvAzU4APU4sf378vJgyDz+4CVFCwd7IYuSVTkhkwAn8mp
DutfzBCVVdCAfllAusDmSZWgTWPPvQIKu7He4P96Jv57lJoz1tnFT7NpmLyUDXRA
dD9KBt1Tr9bnoSubWurkm0nAF4vhJyxfctj4czL3cJIXlGmqEvqRq5qbyDmfb/ik
9LlttgBIZGjPaQ2t/VaGabjKCdGb24DYWygYqxtJknrtu9woeeXERuKyI0Vy/wvC
OZKSFiM9R8GozslHzdyzfHXBVoQ78bG6bgpH+egbdkJwMOAOTjfVR2gYC2r2Td64
QaB5FjgY7LZu7LH96uomslhE5lYVd9TXJNElnJGMpwzlFcy/UYOpUzR4qV9Bax8P
+NJ6eNij1X6MRUe/RfzpUk1JuNlcH4IKNzS5zR+E29TRY7UCxU4uQAQttXwpzcaQ
x9Z2gMaBXX0AlZSatNXkm9ePPStrTGkEk5FTRzInOfIjqZkVXBHnGi/OXmZE6rCF
DWjW0xGMNzxnZ7BbvWa0ruRnSQyJF42LsxUF6g1ury+AJ7V/ZHB49MRBK1oVVW/m
Bh2BPlQTLTBE5EwCVR/0A7AyE+NBGdhGwG8YXFe+ZZ65tx0UkEEZ9zzmp4M4DqxP
GRctFjSJi2ylQQHuBaWcHNlX2bgi4F1CBIBNpJ34jqpVYDEZT9pyGhrtoHyAY0B1
D7imNzpP7V67Hoi8QdxfizYn+8p9qrKhm46ELc4aI5AO4DDyE27BnAeRaxXx7px2
3aTLuQ5ifYmhDkSXofbFq2IRNI+rD+DRxd/mrTtQRirksjEf2ibE0qeLRlzisR1Y
cSacNGmh81+15IOrXLoyckPhIDNeyC8mgmBvBO2rCVa7QkXldVNE5dir1FZmVrwu
/WLoZzkybyzFEOZug4aGNem2JdFlEbGsX3Plm876pCDjSOymrzyXMs08sDptlE31
QmtPja373A5JptuPnAU6Wd8sUX6XmlcVzVtvP/I2QNaYgggkLY2fy6+Qvyrig+45
fZBx/+CbCTiUVvgHYSvJTyWuZvGJ+toJ0YvxDoA9zWp1KzZMjii8EiffkQLJOrZk
csQ4LO7Dwb8pniykD6/rf+244P68u0REbE7qotLSZ6/Na2XU7rG4ohQKxoCP1koV
IN2dLFIDmTVrnnZBT8cblUaGHpFqpVjjIoPqWZVpYuZwKk5cNVzaJVGM7GStQdHX
z7fp7cg9tBweH9+5dRfwGJLh6sL9oJeHJ3j2xF0MODsgPNXNL0iDOIHr0hsMf8JF
r/ulShUJmlmX0dC8Xe+8q9Oji0B93DGnODpGOxqslCevu1UV8gE76eWFOyopJ+iq
+fUYBUpGVgxf7XCKa7YkoskaOirn/p2PtV2e/LSFA6NDrpIwz1WMlkWwJ9MjV/3H
IMaDNS4y+SNe5d0KhnxYm+KjFXglHshtOXFEkXErB3tWQJrkL8lrNFEdzcc9ovvV
BK1q+ZXRqmDsVelm50B/oXgFcBviW7TtuxMLU+DGwqkrBv+d3P67G/eUSo1CV/Je
G+BbInrC9kHIQbYWPq5G3DA1UzXGPc5DUlVhtwqn94h9Liv63l0tl9sWMqlG9SG6
s/fpT4CnzRClbQtKjGYX9Oi/Ajo8BNWEPRYxukAv5WrIy7/kO5Sf5N/Vy48XLF4X
5PdE1Un3b65KkH4cB+NcoUvL7mfp70NKrqB/tTiJXCqRv4lHuwole4sL/rsNZ2Sr
JzfG/OF1eYfpHHXZxRxGMOZRY8dJq0THqPu2IovmdF2I1t0gT5CRbYp12BscCjHS
WGJi0mbB9FZ3VjfajqASZjalMJQOSYb+ctqNqLBs3GH6OVoaT5lK40KiYA07p4i1
utHykyhEXUxI+NjhAmk4EP7xHFTG/yRW8uOCw7E7jK5GwfYfn+3G1ArObllXHSaC
SZJi9YDIeymEDTIEP6hxZ2jikM6Si0UeUZSzln0Via4IB7dTcn0yKoErhi+jNrBh
fIM0DpO36gB39iFTd9Ba71+CGFxTRi8xye46Iqr2ps4NUycT7Wcz28zsXwAe78nJ
14HfUp2Ohk4JMVGtu22Q2V0TbdHq/xMUaEy+cAlkkiakix+J5lhOYmqfHwRleb17
HEyt2vnCg9cE7qyLvWC+aaXVZWuSSQ4XBL5FBWkCSRJVjrut3sgOiieBxNS4q7hv
cy8TuwSLSV1JmA5g0PYYaxPebegZz2k1Tf4wXltS3MTyJjn88FbSx9ywu37OmpnI
7iugkMmQMd5mB2pV856fzQscMIzd+PHMxQRtLNxbUTfKPNeJzv1+uCRbyh02HuXh
hJqgTSW0IyxNm8WgxD8+A4d3vEdjyp6PGxQGQHS3x2oKdKrOFV1vpz+jJYgUbq5A
IrPATbIs/ehgxwsDek+tfg+XnD/JSrDI1VLPxWoY9MKcYZ0w5svi8WOTmkZSXSYi
ezlhRe7g91i6blzpn9h1YfCpZtQizevdNXAugd7KGZfNuHmfWEKzQaP3Ph/ZPJ4j
h3L6yhfF4zZBxBIxlSAWuutJnpA9Hprw0A/IUt4b518e36N3sdrkzQIdJe93XoYY
lmwH7+Xkap5uEmuiLn1BRR4GI4nLq+AUdLNmvkuNdpAnEWQo0HxlEdEQ7Dl+OVgz
NfRSCg/X3IS+POr/LVuAPPyfXUrNJX7HeeH2exD16TMx9rTPLVWCnv7mH4wmlYSR
FsSUzfpQWyWaiUoDULInt9WMGOI6xmXYihpsb86xzcvYBZWnkp7Gvy89l6Fa5uJ6
7FbBRWzjhoCMcWrFC4xhvjDmpWLmoQnzPizXYTqiBKoK+++9RXwmxcb0ssai+niC
4ecejIPppqNOhqNErnH8c5d2ejGHAm3plMElB/+l2/YPaylhCMKdZNQEe1swDaQW
j1NYbWM+yeaHuqAtvX5LcLQii2YRCEBLBb7Wuwz5v+NNgLdBWyaHxv6pp/UHEv1W
gOCvpF6hG9MlSb58faSf+8OF1auHZ8+t+jIhdHZHNZ4HmifqJY+/cFDyLHiZzxrI
USrr4QrK0KqJPsazJwu4mxaH16fgoqKTnF6h0BrfSbTFYqgHTqgwJCDeyNToGggw
al+1sqrBUGA3KgQjoLL94VASP3IDCiSn3ImUuCW571DCeCs7xxkoYF0MC802ZusQ
g0o/p9+BvFy1fqU0wJPIFUjLk6knnJ4rpYeUGbfy02bDP1GkBPSxqsF+VG0F/nVo
Pao9eQ/5yU31xG+T9h/5a5W5veKGtpRjg6WW74WRk18Wd63e3GAOugkHsq9d0ztk
W8Y+9lWuAIEzq6f2B9n+zA6ydQWBeKB1zl3myr4P/muswmoI0FrXrM8X0ZlyN1K0
7XRohd3GMYh4EFMfpP5FF9fDDfjkfnpnFKHNnrTqrRU9wqXXe/SWa7VuMn5o8nM8
KCfKlae7g4OBSrXzdGUVd66y1EBvmejPbiXPFDlQTlzuqb3mwMld2f0aVjYrMPM9
PwQdlcXSoGgpBHPpoNsdeMRE06vSLHMPd7WQZVH/l4lU20OmeqBGNwabVtsGVuxL
cLw+UEkQZxnXKuLYEmnFWmgUp2vAFws6MceRBb/GW8+6iUmljoJtdk9e9S/UPIPg
hBjK8OBBjeKCCuklwowi9GBvmOpzrL8RkgX7iMxwk1Cqk45c8GMMdz/1rSkpJQj2
KEsSLvHDjHb6gFIxoyxhLBlt3GdxNynBRmvnswVqPC8vDLBDL/EhW8jtOdSZBuf+
OdKg2u04X01DC3jq/oFUMOoQ858zRUBY2WohzZiM64if8NAw3z1xlivD3u5BNuim
Ch5QwPbSGTTH3QkYpcfcbdArpQF+fg4tLh6aEDtwu69ecDid7S891erO5hXVqdhR
jPgFvQaCt587RB6hT4UdLGLSmNS8tVVTfX7ont461WeveOwLEXQPNFB5t4KaAukY
Hy0S03+ucf1hYh0YSZcBHfXPE2llq/Q7lFGWCrqhqrdfToPH6HoVcFcLVXnEV1fk
QVFjsVCfR8tleDaDgm/ILH0Uf8nK1pptFOuCXKAZctKjNpplF/wHqR5rtgmPxkwl
XGg9KQFXeylStsVGHh1oxOMhyJTwonRzAHzxVh1b/IqXybO4A51HUTuvhucn3/s1
KOznh9HCDj7pjQZ1NBdm0r/LX9GAzDenQV7GZ2Eah/fq2jeFH1n+0bZXYEdDKIDP
C42/uFzZWzNI23ExszpG2QynWYoNn+6L9Go6WjCO5Eaf4/1XWLa0Q4hezV/09P0P
mXJE8n3IxQYtO/T1w61cRDT6MREMPzHzkzREmLDulcNqVzcSwFVoQxvudc45WeQG
6UAFq+GtnDFbPktkp7XSnCSL9LiFHebTPKPq8o0CF8eSzltJ1K41O2gIbk13TC5w
3pdA6kkjR11GvR5owjNIAywLkkf9F4PCF03B75BpQPoJ2oiKSL6pMuZGCmP18o+w
z8F4qLQFD+GQUmmXJ8/ZNF+VsCvOPMAJEGaV/2quQP3WW85n0P85nK8EAqYFld1N
OSbojx3UhKUm2p4fNmfwc9mc0NBfRqLrKSAK9AVCAcr5RPF93QQLIhB2Xn4A/WdC
PLRhQ3BUAPVOXo8dowL49jg+EK6qkcKJ7ASGpzY4XS6qh74w9+CfYss1QOi+h8OS
NCFCDXEEvxjxeMnZaqFCdxw0e37yUnTpOvwNdPlbG19evC1Abs9fPiEQQIB9vYJA
9epFVNz8JSMZrJVcd2z2/CVZ4pVz81yUSd+4gV+yQmTuISpIAAzCRZr1OngeeHND
dwdoIWXgV0e1cUXowmrEWghwke9TPEZaTB4v7/5dP6d/pdWNOlEBOmy3xGNP2YW/
1C+Jcv/V8ztOcqvJ6J0DKgQAi1K2dxSWrQcAfxfPbZyz13fH0YMeTQGmqJhlm9yT
CI9ZlgztRd9rFehfAfkQOTHh2TitznfS/JLcr1vbBk3uB0Tgp6Txs6wFYnRFizJa
hPZbDrfcFqbdhP2g4ZOIDRFnMgV/S8nyZawnlB9jTBFMW/vIu4e5zS0jnxFXla9/
Jt0hZ//zbMPeLQdQj1GOIhPi9gqE4LUeHoouJxVIvBgsjc3OLQIdPzvBfH0Z1hs3
cv3gIZv+TY2oAsbVVUjOW3mybqRGQby71eVgoggiD4MlL3j0CiiyfgubCjWfzkiH
Ca2K8GXuyDuf8Ze/+rEU01Q8c8N5+ZpwCCuAlF6Sl3RDLSxs2N8XnzHYqM9dt6d1
f+iD9Do73l7qGz+UsXPMGwLn4POLvwuPyyiC1dJvHmSDCypPJDZA+yO1UJ00vIUr
QHJEATz5L7UUDgM8ZC2T86gzAVUymjWEo/1NvOzDJNkKC5N5ZJOPekSPWPqzYKvS
89S6nLjfjYV4u0SMsDxn+b5SrEgUNQ49NZDkRDsMzNzlkeiV1qQbHdQixmBK7szp
Ftxd9CmB9rUb4hFqaojVlsFY9ajs6Y1QoKt4yaanqfmdgpUREq85T2ZSbmbetumA
dj8fVGTZ8AhZUZo28Utb3U01cGb3jWP0Ddv/GAsCRjUxARzHy/QBuSikpj0t9SNM
4MgZc+/7kNZgx3U8cl9QPlchELhSOT8zGez1j0Y20b1n9Q2ioLWxgctIw3nojghr
shL5neRsoNZLHWZ8m8IDZe1f1sqZSvEKqW2QaiRlO8YF0D+JMdv5I/Rn8lX7hRkx
XWMvs4DilFyedhloAABmz+l5y/w2k0i5WMJQ38ot3KwJgcnMUOAVOtsayU4mevA9
l/+MGslBT+QwVVbhQ5xL9JVRlf44W5iWGBzMyB3XHMNrNQ3HMLofO6KiZG6auQA0
AQItceliYJrSJ7IKiXMPJ89a5jOsi03UdgzQY1536uRPFDfzPdTkygCMTbtCTLcu
rT+7rPEgbZjst07H0cPTVzAEkTtCfXrgpx4YbF/pqO25rfcGCVy+SuFbZDANXI+y
1GtiRQiKtD/ErDmj9wqAD6N7sfqnqLsLvMMS70CCCQRY5rskyhNoIRzM3OloUftg
nVyOJfh0LfVqiNX7VZPaWNs3bPWAU1tBxJTHTR4j9IWH4EVIMmANEDh20nKrsc3U
0pasgCDL1gncbK6+E7ZcB9miHjgi20difXbNImoq1KSe5WWefREaClIt/V5eAVEy
f71anO1zlhXP6LZSaqh6fgqjiNc5E82s+OQhqSFA1zt0/StUcBosWkQA7Bntc0wi
pAydb5XgiHyXqbYyeL634nilejMB9SFzklF/IHcrXTxkoJBi3cgBKd50gXKR/D3d
gADzOdt661YBCs1mQmO+ROt6BZTQnqrqC99xJOhIbgExQ19yEwJSno+Q8E6556Px
ujt54EpT7NDx/oUbmOvw4l7HWMxaEw9nfSKmoZ7Ieteon0p6ZlC8KcfbTWnCqDAI
ISglKd+7iZlkwINzRr2g0zCNxSoSXNLOVxC7u7/aTMMDQspZD3Vu12kX5HSP8BKU
LqAde547oIg9NLeZNWPUktqlbVnNfn2Uk8c00kou1JL4Wf+17M+iEXDU8gIh+TJZ
mzxXYuq79UaOU1rmmH9YIxKpu2k6lR92QpZ7F+uBTCD1tscdQ0Ge/8bP74SoPxBG
ho92gxMThbRmMKvWI1GmeIR8WS4oMhDBfwta2FWsOfEI4Y6Faz8nhel5oxZ6EVA4
C0q4n+FZMAGxHVBRJybsXfFJuIGUsjADkqc91FFpZgj9ttXl+BBcOc+J638b5hte
s6ryTDbHR3f0AgXAYnkvcb6MWYrRNf32F/h4kVfwv4gAdQPviVvlA54wbQ/cFyG7
jgIZ3ma0NN8362Ac4jmYfVqN3NODu3QotUdypi1h+N9iVThcgQegxIazPV2/Hp83
2N642040g/0er/sBA6b5Ek/mtiJnYwdgZrX8x0nLmmQh8BkyroLw2DBfdqjBhWsl
9vNElsoCbg31j12ytMrmXW8gVgalXMdUTWnHySzmscOF4OXxoo9PX4WbOQl2qglh
89Z46CgkVKd+MjjS7kWQCFw7HCPjvfJ0kdMid/0mDnWWwc99Uti52vb14960zgxa
O5CSf3drsA6K3JHGfVMJ8jSS807TL50FXntcT1BMrs1W9TzJ/VDfkxwGP+X1z50x
4kTxKrNCvh0p7djpl07konWQkSSNosBKpSgUsW5I1Vr1FG4AZXyA/NzKMMHtR/db
glZYDLECgn62TKf8t3vO12T7SfE9Flg7PcbKAoCW4fUExDwLSvUsedn43Jkjaih1
UYPcrRSq8zYQC3rz2T1/SYTw0pSSiSfVUDeFmcZgWa3BgFjGfW7aLyLBGKmN7aiT
li9AAB4/nSuFOcJDgB1C8GE2H+bVT+Lx4mXE4MtiB38JXcK0B85zE0vJfzI5i985
KkRmpYve0b/ofG21/AOrf7rwYp8xHNOLyT2LUoulapC98SuImFgYweb6yWwWtN1E
hc+FUxvjcokV1qoZlE5ctGUdADyDBqj//SKk5PRU2Ij16rIr1x58Q6Frs+qZ8EZm
IYJL82OhgwFxuiRN7vhEyz0AiMnHdRFyye7FemRDj9arAfvfOGzaLT3MbwtAO3Bo
KBe57TWvNH+BvFkjivcA94U2CUCcVT2+rYyodASS90wmmY3EPp8wWSwv5xSJw1Jn
agfYjYA4BnK4IbCewvctGOZETIpwzKvKxpSMGGltAolFab2Dqvxytsg7QIJR0gj6
fkrjvaoeoDkg/9ZqQ0edlLE9q/jfc2f5H/AfDHGbqT2t0yf4NSeb136lA9TBJ3xx
qgLvKx9TVDAant1wRkZbQqLpquw8RGsdLH2CgQ3S88dSMNMUoL1Yb1xoea8Z7FAr
UAq+gZwR3MHW0GwYQRjYKHyG2qp7+qRrN6hWQA3A/TtVVfhO17byilzFyk7xw43B
Dpc/LpC5bKY4HE2tvU1M+SRaMHiJ4x4dpYrh11wGMo8id0gL0ibKy1ts0NXn19gh
ryauehH7diq1wmyrRB17bBFLugW3bp9/rCUXmcHCHIbFFKRG3YNZ44FEccI+CRVl
fa3ABDl/o72vHFWHqQefVqtoK0J6ZUqAO9Z0KpvufE6zCPuPzBoTY862oXMCfliX
wnI6HIeBmuSQ2ugd2s+G7EicWKhEm1PWfR/qbQyi469aajQznRGCNN9WYyaVACFq
5Vy6mvkC5fXBDRKECBBbktlc/m6F7T9CtN8X7VIRcppcC8qf2E3cJvuYx62s7B0p
gbZfqCiuf6YMx+Lng+beH3tY74YWiCH3qNxvliVnO8cwJpLnpiVx+KAYvyUhZkPO
On/KAogPfSQ9Hs9AR8yO7x1Kdha+lPZC/iZAg5ZltmUY4Vc/vqI4wWtBI/daNCPY
QbH15c1Jd5BTHVnQkAbOCIbtFAuxGWN4kcKWgGgAHZ1xQyl2DntlTgNdM+BoVNRr
0yVzF9fTVZG711N/j6uxgzItVEQ9ZKbVDstJzU4FDB9I55mNKFXf8AUt7eSvZNTo
HLdU8xWI2A/xZqqBkfAiIc3hGv7ctTbnWgdXb+3L7sEJoiYUnTURkkwRCW9rGBJG
pPBPkxv8HibzAVAeFNXUSB7Br75atm8YPstQB/Kgo3YTUgyJQfzOKrRG32jOgOku
Ro6Yy3m4yXwADAGxQeoKFXyzvrD+ftiliQeD7s4RoP73oK5Y/NRUBSSM05g5CUZ7
7mUqBdFKyKYm0eeDvjg+HBtL2XCyPnB2kh3f8XaWz/z3Nq7z4GVrfbxwBc6fHtfp
reuZywdwg1eUqZoQLvnrYTILiHx6BTU1avCZ0fiqLfm7/OsyoPu/8za2CHUJHkU6
beXY2vEU8dL4dTpAzZwI5hAzq1AnRlveoXOyZJpKXlV+P6BXR90Dyjg+jmzldvDc
3/LqXY+3rzOL6UG1m+d+7oh7oI0A5R/6t9/FNqJM1/qEHjHFyR12a7HxkceCRypU
vvroo3LW/GFiqKSV3ereS54xh9QDsql5E0hns4o+8iQadXV5GrCLT+BmkD7uAB5y
hJtYjKFnmchSbdMndnt0Okuzz+kuebzZKw1tYRBtpPaI2n3gkIXR0ZBhLjDmW12R
7vOB8TLDW/5IKliGaEhkzJXrxFcAWtBmUijmN3kwmxzAnm4XXviEq2Sj0kwVhQ1T
kvBtBKkpNGDaraZuaXL6VPKEv4zPVKZIZCnLMTveW2zSVT5VXasn5RE+ZtJ9eD51
geyPiEnEOUyE6v5JTPIoDX9DriAv+MRpGpictVRdUg08ffc9mlZvZKwnwOWyOgz9
A0G+RMflxKYSwvZmsXJ467p8BHhULLu1c9GnDJ3ArMyml74dn8SgwIzKI3LexIaT
5L8BUkKj7OTTrdeneY9LKR/5J4qb1zDXG4m7WEYs3HoW6fdaHO08R3ACc81q4dd7
8ZiGidet4wJaYhtY8ueApNDk86OvPQLWcGQa4KWmIcW9LrXGjt/E41qD3nfRfgmq
sutZ/vbAt3M/BR4tjlRaK0umLtGO7TaPLwC8FztF8HgiOu/ahl2kUEACQCBVlLUH
cWsFYHAi0dmJ9waj5hz9mRYldEV+CAeVCZ403aQlARWXd+laTy28xM833Q/HLHYb
1yDk07fiE5GVi8khNWBVZuQrI8k5stWH+qn1f19WHEHvyue5TUnYeDyLjAQo6kZs
uIR9ZNVREJIJZy4z8apb1BUANtXQRbbjvU5RyOO3cyecElHybUKuSy+mIN02G7OM
0U2a3qY6s4IlVajiGc/5hFfYi8IFBlAnS5T54Pw8Q+7cznSw7EPNpZ+q0ksAm+WZ
vP3138NKnLpNgJuDLslDsqEVB2cESExxY2xKqKwjsHubT03Hh0JnL7VhO14umpMT
yUEPzNAq8Py76tJCtd9OK/c8u533mheN1pmA1cnTVlACZD1CHfNsy9dNZat3RiQf
LC1V066WYYMQp7QfFlO3WoWvnNl1KpLOl/Uf0UVq6AowYyAFBEz8QOQsMEKh6eib
wVpLNup9eJPpt6uRs1zdAiHa3plyWsOCFD9cVn9FLuYkXeebB95cP0bvY/6MApWB
uDTcljoz+Jwwk/o52R6Y4RBj/EW/Z9E64cSHjUYrCAdumYfpKQCYT77OKniFnAsU
XiMkyFfQvdBacL5e1TVXQkCHBtBgH1nxykrmm9Uk1DtiDCjBaOaFik4TP8hXwIQw
+XW2ha3BcVJ7eIBGVXR8qsFqrKxkqLS/AYEGZQxMX9QWSg6wVv6KLJhpya43ZDOY
LZLboaU8BPjlSDa4pKt1q53eiyh4PA70K6GH5RY1QYEDu9TvC3nt1QOrUfL3ctaL
sEld8Kf+m0Itc3hgCIhBk082/gWDTATv1q3KnUAg/Rs5Kj3DRo97uy1VCjZY0lLi
QgAfewK8qu/HztY7GpXwd7OmE0uDbRBIxONwOVDpeGWO/O+LXUgEfUxG48AHntst
IC+PF2CdwnCs050XysjlZ/lIBMIx7s18TJV+hPQAQ47kGC2QY7Qa0k0EiGLyT1So
TYkUSrmuq7flfLDQohF1WWWeGr8j/IMW6JsGIczM7wIDwBKn9Fnmb9h/0I31XQHA
97n1dyvUeCA+XYT3O5eHwysdFRfkPWLg5YnfZm+iJsl/Tcq8fyvnJQYW7ndpqAmE
jCQxMGbCm/4vPogS+XNWZNDMcYWNadAPgx3GFgTmGCNu4BMg8IM9zbdn2sle3pWg
aTWBOrei4kvbDy0vj/uiJWmHqG7bw+yjeDOZa+PoCjF5aVMi6iRBN3zVDBXCOizL
xs3r4d2oiHIfhKz88dbpTVskIcxkjyCWNjqUZ4pF1NMH43eA1mwS/fg2roLEYESZ
gq+wno0n+zyOMTAoqSMxhFk+kbIhTbQ2bpyyj4pGTWKbqFnqfQ6T031X2H+dkR0E
zXGQsX0EAxuLktCPU2LzzCFe2j7WYNjGMQCJqONtPALO+NfxdeSKXNJtBsp3kQ4V
MPDMc4oP7QZTU+8LrKSeaFYhZBeVGHc/+S463wQmCAx/y4DdJGxlCAkiVpMuH6WZ
Xf2GwrsxBZt8rEfj+UpOI0kmke6cYe7oFNhoZcA8EeOvdqwt8v0GMAtwkhnFJH+J
3vXWs3BgVbHDFtXBoRNEcljg5fpCVKZBlbgec81lyv2PotbkA7NJ7nQ5HnECOvYT
sYPfTzSEsvmFQaZumukIgLg+RbDTwCZMSaieAt4Ta9Ksd50Reuj20WtiRHO0OE5k
vA6jgmrZo613SW9w9YgLitaEAYkzwKxdoSZRM0uH+HfWQ2CaqPfDfLWK5CNu38Ed
a378uhIhWwsAQlTb4FOImkyylSBC1OJQPpaH4Fw++CAKF1+XGdtw+l8sM6TM+JYL
9ZxcXaNLHXQTzs/mzEJHlxsYwxjTbwgQ/ObmD2nP50V/ekQWfm7tPHNB61Oz9wPz
KJvfbjxxXwtEgFZ0K0UHztoEB8FXiLDer+4MYA6MaSos0NAou4TjUYeRs2AEmI1k
OqPTbkInwJQ4/x+PJKrygJPnE7KmREtj3YeYbiF6DblUIp6nlwkW95QapvrWSuKb
db/UXWA8rf58f2NRxO5WCC06GjHMyfl0xue5JpIbHVOJv6/8qCWGm9DISuBStZHy
7fz4Hs9Wdi9tbOJ5f3QyF+++q5ZR9IOMMP+rJIVTPw0BbM98TyVwJNMJwNxEeg25
DhangNwjcY52oIEgFgjRIJ319/vVwr1hsv7L+2vHFCeMvtaBzdZbuE5nmSGaUigt
MLaiHyBEW0t12foqcJL1cDFkfRxJf+SElFT8rUaGa6uPHVSfM/ogQiPkFHE56bah
A1eR9vZe7Y/XOP8p3wXQNT8HEoPLdCT+XYParVJxY9FpFyf+YGEfc6DuV9/yu06L
KQU9YGpYaGsfC/qPWTwssKozJqGNz7yT+f+c7j6PsVc87Iyh568sU+uZGFX6N3Ii
BXyu1LmS5iQYUAkxDPsPfAcFtGn76QiRNsgKEx9NeONbUdb4FWF4Z97B8fmD3oFW
Bk07bhnYGK7Sdu1wcaTfVD1LFzYlKtyYkHBOaiGjPuu/uSj5uzbXiSqy+CsNav3z
IgMuL0ZBFqVw8a0VqZt9a83x91nr9wQbqoBxM2vyjbwzvaV0Dcyzi9PsF7SqxBMZ
I7aN6c2hPlIKWq9EdjC8G4VIc2UrMVAZbTQa9cc338qgD8oTZ3IWNRX+lnckkbAV
nJ7uzyNPJ8n38Z2N2PSWvobrCACabYH5voRUiu0BV5CRjqnc49c/vWHIY+OGjZrl
YxyIEPVMgnQLo8twBxQC5yrkK7/jl/lW1qVP6Adnn23+tEjXxWn2Zlu0u4zy9Kp6
KOlqX8qmgVtF2oJPA4HyfVG/lZ0whMYrSWgrQCFELfVWnfnvJTjKOOtyLXfmXvuC
mxIxlVn68hlNxA0I04pxpXXHU/Brinqx/yjDRRPcs3009mcNgBgHX5vz0Z+UkiGt
Nof8D4H9lwjZaude5qHP1227V2VJXWfEM8dl7SoTX702lOZjjzLSrW2AiS2YqdYw
lK9tw366HiysXmZmFjdfhxQUF6Rj3502mioKcgJ9TkJT5gVg0gV4QGEdmuV2EGRe
kHngPnKmTiy5XAHeaaaTTEqvuz0JXomkACDnaqdSfr5rYxqwIrdqk5/OEkrMQ33G
jL4WUpZHUGBkdy0vsIEmk5ykc4QJl1T+h5UJUoIqkfic5oCK2EVb9kYP49obhD5Z
ERdNNR3BNMcD1MFwhgXTpHEJO8MmrksQ8GyNJp3GGZ4htNq8dbO0pXnVBFOJXTZQ
WFvysXRb6EQbByJABM4nfWpxy1yntbwzDoZOyLaUZjkcP+u2Zqdk2KBIt3Z5t/2w
bK5kgBE/aAFJQz/4bL/ZmYUrX4OuKI6PH8U4GBdQFGureYKSGB5HEXv8a10KwyUp
gyD1/oymnms2BmyyB48LgvdP12FMoW+6p2fu5omnHLShhNS94S9/QCM4NVvFMOtL
oG/2Z8A0IHNpKfWXTQZ37FLBzDtt/VvwLLoZB+2kIBbFdzs6ZKDh1hJpzr8w5QPa
BPyuJxzMAh3WUDSA4A3TjNaENqjRz6w40Sv3RiBGbyyJN0NrC+yyzaCGcrjnsNXU
3DES9EwoyxVvPmuwER6wC4EAo8uEULoPi9VGbAoFyM5Xn2d7tsjjsGa3SxJjvSmz
tB2ECYEFU4YqMGZFvANnClkAb+xqCBdLUEDcVmp6txXJJxMK09bPtTAO12rG0v+U
Sz+/XI1JXwodTLA3bM229MCinNXtX8cwCTUz/rR0qG+yMyxrIxgTHfGUM+psX8g1
WSeoxXwp8Ey23MWUFzU9r9OkCcDmsTQVx+VHxvqdOIALClVCAONSMbcquR+dSU3F
c94rUC0oT7DkwNNz40Tc6Cq8Z3mMdeEGY7J1jE7MHqO6SXsfAkr4s4s+MrlP9IBp
lt3bRH0vJTBWVzV/Algm98GfYaASIXy6HCYUo/21eKUqQB+ysNE+UVzE1YRF7PBD
PJ61/060yJHlW7VeNBTjNmoUtrrdOTvKGSXJ2I34FEv2cJpgloBBBXhUjkgJ1Ecu
xBzlqcpB5rgZzrUAUO1u6hLlpgka5O+L7B0wJBcTF/5I24L+3+mGw0Bf2Fvn1iBF
KMuffQNrCnLQsXwpidVT8UVyUo0Wbyq45krxlTuGHXC3X/HxvbnYsgg3vGKCin1B
UIhin7Nbb4Pob3Z3e2lVqGjCiVCvwF4O+z5EHhd/4YtjDrpEjsiyQ0CQeknBbiUy
Pqog2AS0twyxQJVinwsqS/n00agDDz3k/xCgrTuXmxJTRLJ6wvyWMQYmdZGu2WCt
hP/2WOQyUEURJG7dT2ijH1Xc0fyk0l9NhxrHjJuh89RQ3Sj0RGerxhHwzw0yhNr+
b9bMZAw+jiBD3vCuszg9jNRRub+Lpg3EdUBTXkRjB2iiom2ztAnBeq8wBGEMvpCr
DEGA8JS1/S+bwPV3eYSrpitQtcvfuGxHbv+1e+S2FTltrykmfL90PBZVzEvcKKyf
YaVzmqiHzIoNmUpefIqlXELruqOC98b1v7mOlyYu53xTsexqx2g2FUP6YOO6IOWG
9fsx22Oj5Fk0LTQRz2NICZUGex+qvZVnS/9+MkRgQ1NaSTgHBtdTh7THsmWf9ZMw
vevjD2wusndGrJ4XVwxMUgFApjkkEDePx6WTDkjYVC3GucdyJQN/HEVMvNbz/qM0
umqlizxx5DhM8oegmy1QU2NpxyH56fycs9cxWWIN6sZysmg3HRRVFGW0RlPQ6dfc
dO41wSrYoxiQYAJLtdtVa+d3tPh+z0mPGWm0it/wcJ14/09QDoaUTiDWX6HND7vX
f+U3MX/A2t7++6rk/zEIsVsmAFTCdhWr4u59EkhQhjcqvnh4c5CktKkWFSNAZSCX
TlYVOIDXs5qYTJfwKvifHnFshv9FODObAq4zMyXuk2LdTkCFOjIC16tFsfiVvze7
mrPJLrRdxBToK2GJU9Yx7ksXsgL5OcYndnFF5wFh+timPH2LD2J6S6h1q9u3OEIg
ty/MiS559NzLWpzQ0pN7tuoDwXCr8kI5LgnQSCYxTtVKKEZAerSCUPjQtv7HT/y2
LbVbs0dOTRxpV8XeEGWhEFF9+9i8zK71SNH7xPcIvWpPkG7UTUxwgGZB5WACVDsO
ombE57yFvCwy3rExYyy00MLSI5f8dkhjxpCvITKRygI3eQy2XgdkGF6Qg4KBD4JS
14NNkDfpaUVMjVFd5dd7i99pQUA8q74kQba/7GTLRnc8MOnfh8cjPXFo5t9sRgAS
sIzkFLqVbzdMmDuwLbauqccXzBkqkJwWuCQe0JDCBxJJfyipMrdjUA1l5p65psB/
CHVxJygK744NLE0ff+OoYfSxWQLjVCxtdfNjZ9Fv96WXKmBGmynqtBwFcWWlxfs8
LqganPdpNftPPB5Tkt5aEVdWpGhC8KjHylC8yd/F9P3JcX2tTNn8F1kRvfnwvIHQ
+NuDlNJlIRPrD1eyaq4FyRIBMirBfqNFOveP1iSa6/CSSQeQ/NMqchjU6WF5WPDV
sdyAFN3k607tt7NhCJSqGaioSuR23BHAz+tHS4rWgTs9bVqr2BJ1B5bv6dt7hm9K
Q3oGBy5DbiL4Eozifl6KSOclij3ishAYQhi8QSxPKdFHQ7k/sRfVSVuiMFFDlyqa
Md2VmZyvR56emQYrmzDTfKFGkQAQuzdFY+EabWMvsuQzAynn1io8oDrmB5quhDg8
jURkYkRJHre1z2/y6zk1hxHcOw0SRF7Zd4jPz09WA4ARAumm5DmlJ0O303mf9nPM
KA4LiIvji5t0kXeFiuNu1YYWjb60mj+eIFJ7OM4MwAVYg1vyVrXOHjI6pNj30GCU
CipUbsN5Vp8C24azlaVwLeRiPvpZJTWPFPZ6Pyjf7ZV9H1/mmhAx2ytQNgN54Rdl
LumnhdoDqxB7mkHJ8x2C3c05/JZ9SvA2V37W3McJKg3ev18hC/xW/DxuWKgfRgyO
crM1+2GgXljCueubNgSEtfSnwRLIdQtmFwwCeUKImeb6ofsKGr1TjO69ci9gE2cz
hnWhyCoCsuXv4hDeXQmI/+SxF6d/zPRHj6Ie/Z3IpuU1fvv9u/IKxcgif4VsKc5+
LsARx2Tr3FpABjykD+Fw1VnW94zo43yWzVENpwliKCSzYEglec+bTOzJnyQ+LjgE
yNMjRGFPa4YJf0ALjr1nJr9IEIcMPyJbY5MHsZCKIFg+X+Vl9HZsFdAQH0L9tByx
dJ4UPyRCpkDzFiwvVtIm+wGeQglMtygMJn8vup2h4CbJ8CiXgIzp4+Fn1V/k1sqO
oM1AzkosmLE5MdXwIHpQWXCBvYp2tpLB4LiqISzqFP1x0fHKZbAg0H+pG3/8b06E
g3dTDWrqsy5avi2qlPspC/UqObFEsVbamfsxBSQvE4YRKHm9NuSEMcJGu84CKFyK
tbWhNcmqqDd6bxb23Tyf76Mb7hLZY/MOncHfZZ+yawOZ20cLnQwmoCOkNWfsH047
9wGwqRHyrWgPCPCeiXnhmVMOKF7vihZ1XtjmMU0jyetqS9D74fj2W4YbaPwBm/kO
6ixideatyRhgYApJQp67QbWZ5S8ajPv13PN1OAN4SiPAhS7TxSUMWFJpL3AU7pld
LiX18vWsghxqh2eYp1EZGKcQc7nmTP1g8WvNKUDDm+tJGkLm7LW5fVe+FrOBdogl
4Dt3QIrsTvEjHey9lKcRbGcLSz8euWT1xcOuV76JCpsR15sAU57EWVcgGKWNc0xK
kjuZJsWDSBG2rnDVrXP2gF7zt94tEdqFwCjNOczVBzJZ5HbmdUvc2yafc3UxHJ3K
zrUOc4lJLhl/OlObEiSHz+dT3eEgKvTdvayUw42fnrC0quw2A4j/PtjRRKyG2Guj
FNzRSWxekZ+JQrwAPee6NnBtek8q4o6yHh2RCZeOqTYISXpxU6UqJrGOUIRsaBUW
JdOYqbiis0+pdo1ly2F7vn/wM65TcKnMUUao20zXWXwJ9ncda9TpwUXEDKuYfggj
IhU2c92ZOVVIJN+uOdBKkZx+P7t+HuAGEAb/r5Gbpb4mgoRrdADtvdZLUk+5XecK
72lv8vHlhNijvBEFKuKuhkfSF2duO2m9w3rmBfLQQgHM9bdhK4lZx2gCQYDTzvYu
4ckQfnqN4jmY1oKO3rT4RYs36XqougQv8MS7mLI3wtn2fq571My42YV90rk9AGn1
zXY1hOjrIrHq+/KwgxB15lHqdv0ZdG1AVmHjS49MBH35yUPqy6k2TZ+c0v1pd2wl
sMcIZLIqnTL9vNb2j/yXiDN4+OYOHagDx9kXGI4Zioojp4fWMlOcfdq8ovev26fr
YS/tyl4WsyRbycjPHs6PRnXO5Be0/dHAjaLOc1LNLIxBPwSOgkuCLxfTKgq4LHXE
myGjoZ0NcXloLG36jbbjPdXU/v68hopi9dEKQZCh0Tbmg5mEebVd5wikTi6IVoGG
v4yHtY5WGen+VerMX5I/QsD1mD2b2z25iyHOlrv5LjGFv1GS2GdzKh9QMKd/3a3U
9I+uZ9C4LulcXzJ6J6c1pOwUX3Id9k2kzEzjAzWpo0fto/231QaTGRAPst2oDpAK
Idi2ikShGKEW3ogJY8Bq2KHtTQ58WiqF9odz+b7bYBbvZk44LtAOk/ZUrUshsvic
y4OfKaWvJGfPnTwmvWnnCShL4jZ4OhFbA5Yev+7rh96fghEj1E/ED9EdKJESb2jM
WOMgesS9lveExkySFTaxLF19PDT44HJ+tyuyx/PtjhbBLc5ETYYBbeXj/Cph/8Lp
IRJeCFWV4d+x/riwOBKRi3Wh09hU1fnqjly/TbzGeLKYagQjKL+ZgeUfigZbFxX5
Ukl90zEOLz0SvSm81zQvMdSWVRPdjJsCMNQX69gVvB6jHbVOJlAMKHSnlu/ejw4o
wEs95Ydctee2t0EU/FI6mlj7WUSoH8rP2MjcyJSv/Zc677OFAPQF2/6deauPOTwU
EtQ+7C8M5JLInSXKsbU0WLZPhurfCb60Ht89uiBDhiW4oRuD14OQIAFC6BATsFFS
C0qiq+r4/92F1pKeOoIikB39KO/53m1yUGzogUt14qXYwwz7sZIbQyb6E7hhEJvd
3yq505b9bzGW3l3TgsHd3OZEXmKg4i+fbcChqFe22Ktf+2WEylhuOUNG7e8ph9O3
3RhfSON5oEzDrIuhdIoAQ8rrQFJnEA9XCp6D8VKfCPfNu6JJul9iCgIKFzj7n9FB
PP3PtskbUisr6XvjtBlioKehBJMcvb09tGQJjeSuWSu5T2Emwd0PeOnTCf9Babqp
JsKCANr0d2QHe/ChDayPksSWWxMmvG3SwTGeB+AQyexIDnv3jeosPX0FWKYCjt7E
jIGUW/hsN/42EKhk9rxzsU9kqRGi/vHUYcyAT1MXz9m6o97W5wco8cUfyMVfTl9C
hfvbd0CDzti4Qpxa/wgvyqRvVOOWwmQjSNrWPXgFAWKOJVDIhEg/Kjajnqdg+0jA
1OC7B00N6jlLIbDgGGHVXujYh2Pf9WYvIEbQvZLrNCDnZT84uR5EuGSMgtWSODUO
Rlde+Kxmu2E4nmhIMnD6SZumIKBojF9JXk9kp73AB/8B/GLak54ItMoHepKMalvE
wpFgecZ0KqZFfrOg3Dv5WLSWNxmcdzeetx/l3hmWlL55rbHtxhHBFNTq/1mDgKD8
pO4ukQ1RAdFE1Rut2RMfVng4R4dHrsIAyyRkdREphhyF2AZhxSlrKkFI6VBS2AGJ
1iNaIYR7wMbB0HL5r9AsFFABtxQzxvDbuH+DvAXpPhZL9Bo4oETGL2xZbkbNpk5n
1MeKUWTqZ2r6Ygklag5PaGbj3KeAg9sYcPSB3YmVzzVX2KQH9cJWrCD9Cv/RBcCm
yEDrPjkGGJlj04IGZTFjJblpisot8CeMAK4NYeZGnLbv7e4p91kk0YuF4XNX6wPT
G+uwLZDq8T+4KBTHz0JB5EF6qIKV/yrKvhsGU4pYSh206HICMNCdrFS4Y0IraCrp
cDcYeau6rdjnF5X89FeL+gagzwTYw/xYM7+z8idDpgXq6GwEZ2nkPVJsPSduUCDA
EJf/0oYrMVSTE80cPulSD6DanJXGfiyWdITAURQdVN8CrzgjK8S5VI0IyqHkZEW2
U7gQaX8/4EcGUSWAgpVpPZ+I5gqoodCYd3YEyyLdE0RbGwzFTCb7dJZ5F4seYm6+
DBtea/7iRX1dbv4s4KlIiUH3rtSeGZfbdPpwT+9zfeelhXyYyphEr7hf3dg6JBdc
ODzeriVqwug4lDokZ/uZVDKv7EOtCqV602xNTkPGzOBFceedWVeonhYRvfhL9LAG
mCoqXhdRtbFakLxNVM+z45ELy0gW2SGmqB42/I7NvHcA3wpCPU8Zrhb4NtRzoTFA
UxsiJO9rdoz4ESBVHnZ2oysFgtTzocCpoJyc4mgy2l7OJ5UPoIEB7vNXnQ2zT62v
snhOJdP4zx1AzpkhjJn2QUEEBQ7Cn2aL8QQ5t8qI3I+cKnEp1pbQKYwxcDpBSR6/
oEP7ssdH5njbXKLPxNMb7Opq50Hu8IH9Lnr5TSAb/sOSjI4ZDufj0cgY8AoNOKgt
pTarO3o9Hd2yQDrNAB9UVMDyB9RoMhOxQfu4Kb87IGySPArO1FNecdjccA+76cy4
D04IifelA1yMoNdyY25nJFQFgRH/yU0eF1XgGj9ufmM2HICKu0zo0W8xjLjUHKdu
/WPOIGCdMXKAl1OCHZhEIDaqMyCbm/FElk2sLgqW8IyG2zEi+274WUa+FFx8gy6q
RtpO6MMjvQJWI5R5KUJ2eK7gXaMUCRuJmILXpo6/Re0mT6rMmTiceuoG+UCsePR1
UY6gbuG6GYrLP7UxTiBAJWcweE7jwSftbFqMhBVc3ROAQ5OOP1aaD4OtUn5qfGAG
zQoHHRrbzFK5DDfE1FGO6U5nP469f1xShUV2LQCjYo+h7vmPQVSniIqTqOxwpkPh
LY1xM30KlJKI1exVEak/sYM1Y+PYKe98n2dJ3mANHErbmkXmSzDs0dgR8cGZgYXX
PBFqvbsA7Vi4dMnaRDZL3aMpoxUkYV50NkJLdbit2kRGww2EgNWWd/MCNCp7c8/5
yU9aQHFqXtA3IpQ2tzNiatspaXP1KtMRsSHioQDSHq8QWo6Drg143zXyNBN9BWWs
ciT3bCWDT7WM7+xaEZBagfconN8jWwE3B+fx7SmMwKURyj/kQRV4oz68WraasoDG
XXT8B31tOflQkkbPsS6EsoxXFV9b1CroXRif4XIikbgxqRpTV3X/+o6ibz1N27ps
AeJfHSjJEzH9Y1FxmFN2mvRuqoYyQkbNLmy9C7XmlE4NXKip6uaGQHN+LqvpCPwR
b35lKsqY3WodfKStNq/JXO/sQHeydTCQMZfL1TBDtE4ElccEUic5pIkdQjWpAGoA
IU2QixdSQHVU4wNRoFdTEXr+5HPc8GVmJMxmJtXfVNd4Bpv7AbbU5ZQOxXwHZeM4
NrE+phrPpZ+lHjCjqBODlPqYrlHCqGJf/y40FMQG4OdrnbF8R2BqkjL2uQg3MMKR
ep/SuY2LUTdjrZJ4Ebx0tRQee1s9F9ZdGDb8lTZ+taLy+UCWnrbmTLjnm1IVMWKu
Z6kCvskV65deW09K/7jWcjspZrPi3Kit/DIX7UnXlSbbhWmFLShUhQevb8TFBZhE
16d5kGn0IyyKBqqeX+qi6HxrPBCeapl1vxZQLhnF48TcGdjgeJbV8iXwrocHCKd+
5p7TjnqEhvKVkvERwInkegbeu66hkm5nBX3Q+fdMXWjkSfzRvJfhZ2OEoyXRQYe1
ZVwr6xh7qmxfhlOjXfPfcvC/XcLuVYyOpiW+NfLbveOjamEEwgDqRdp4pKinRexP
fsmeXxpEvJiSOBjMEQ06+i4rQfBy1Zku/zcGQhei9Gna32Q5oXl/wRV5ccsLe/Vw
5qsYnKoPwzZmrfqROCmBHmLFmRH9aeeUAOnLAckhUWMiIis3c1ojhJi/SjBTuwxi
yYBsCHjIL/uvaU6BDRYgtjwblb5OgOaCUpy164H0UdFTO11n7inFIg1uwG9h3AKS
1WvmaUoDL3ZeZB+I46sSlgdYipVJ5AKd9hw3MVewudKuARSDxLAzJxnfMmwKQLu8
4MvfxtgBsHTdg/iDowlylhRyWZxVUmF/KkWzrC+4lQsT1N8k3hdIGYFrY1rwumZD
B3Y3bT4mdEhkWVZ54IxY5F4wPfJRN7im6Z24LCygRapKOPlRovXH8LJMkAgDV8ei
eM9rlZdavg74RkzCertc5rCF+B8TtdTXRnG0mkxXdrg4tCvHzkWeW0NLHknx2RGL
WIj5Z8XNLPE38X3QkXrfcQ7awnmh5UPTlS579iHxqgZETmEJCswM7h1pAj5dRYZ2
dXB686+0T5v5I1+KmBoU5kq0jTqDyxaalyQKSSXy5TYKGh9ZUC3mdt1BOfNELffH
nVqCgu/fBftNarUiZnPE+SrTy4+3mLcMk3LsFTPgANcG4XXJHMwvkMV7IpxtXMT+
RXWAog54tlo8P7ItiEr3qkU/476zdH/0O1QxVqmF7+wTCTMRPklCIv8YYD22u1B4
sA+S6d3idoN6y6hmiC83BWIRAgTZE4Op1LbjE3v45qK5oXCkN39r4cQWv+JwvUFH
+1rjY+KPp8REHnnN8ZOWZlreYtsh9mWfZEeLXcfr1zHxVx6n8ot05d7IjjxRPiaH
zBh8vef3R2vq1NeK79ywfc8/ZUAoeA4vz1vasFBvw6gb4NafvOU2efuUnQ7Rb/ga
HGJM2Rejmb8GX7IxqggqvkmX7YSWfGm9lDkYdLvp/Z03GcPR2iiKPmbRGsNCGOud
KoFG7AcSs5EiQ/G641oUm3NrM1QrasPUGOXCYge3kS9t+UuKLVX8y5ap8aJMGIdD
m1pLUiGSnHd4ipZfwj5qH+/ghKcSKZjSoBrCvWpnF3d1a6VxaQYprHYfV31M/B3P
CqD+i6U3TEwTMtFMcxAhrdgXXziHZ6oDwNtOWCjzHiV+/ZXh+z7EUBMJCDQWrqzg
S/0M9pKBzjVGZ62TdyMqDICt4afa9z22ZJzBmjIGgv/NiO2WPlkk04lmXpJGDqn9
x46AVSGIE5w+cOjX7QmAQy+WrskKdzt7xBWNFqLaToJVUi3MFijt/GK6W30KFLqt
JciiVxgIAf1ChpzzFHxzwjy0ACDi0k0V/H4pVNzQJ0/VXOYOOZer0hryKBAX1Gjy
pgci00nvq4e38oCSv3w5Zfv2AepR74RDNUwia2OD5V/zS8GhsGMY8oA2HLPJMdon
+/HHJzv9JVjw8RMzBeQ6Hp7tjJBKFrPz486G71kGXGzhxIb1jkbw62+BnkrmWs6N
cMZuRv0YgVyCOVoIdc5ZK48sZiSoQY9s+uA0drWU+FDJ+re8RvqsSLXlTpR7qu4X
iuAxojBKhiVm6INjsXxtmsAhLCpQcLVc2/BKzLUz03eSHE8CVradpoN/SKx4Wm2z
JDeBWuTTIny9KcvuIw6YKufK+QSwLfeM6cx9ZK2oZfK/UZ+fJQxCnGLDyOrtLVGe
a0cgIv2LrL8NTHiaQ26hm6z1b8ogSjLSn+Y8CC6GOYOiZyv2/w36mX9QCzbyoeD+
q5+C5EmmJu+CSCn/pQvL1QN7s3CvHPh8Pf99m6r7TtXXwdzZWWUALbKsrWn5U3Kf
t21sgmMBfa5Wm/EGt3vNvYWd9nop2pJZJkzA9HyxdFka2vY0sZBpVIJF4dyWEw7s
Dge/t9Q0qedrQYLRzf/lQf6iglWVgaY0gXYXQRy1Pf9wDg1pG+5qR8o3RdajdiRC
D8injEzDTFRbqTmsk3j8HzL6Rt6uwZmCig+sFjogm68Sw66Df4sEe7TJpT7IlDKu
+kiRePIv42iyiXX+R4PSkS9dI9pTlYq1+TmSQbXFHlZzjOe34VgltffDdpBBW0g9
fqswq93o1k/72lLNQ6S6HtpT0y/33wcPFlqW7wG6S9oJTpIDXuMTndo7NqOxou6n
mTHtRdzwBxFvQsf3wAtN5NWU35Mca4FQRYpwYvxAA2510jF+TuKmTLIVGXyEsy9T
wZml+SmhmBsgyzPy8yG9N5ssZORDZ2KB/Inq2ZH0wdAwL4vBOZdMG2iHm7YoV6JI
5yisoC1vwNnK/hwk6Pw2kGVaEO5SAbYmGouOVeWr/u5j3XfMEMa9xqERMesVxj5L
M/YXClb0bopyL6nyx+FZ5JYOAXxqiY6oftknr7Gpu/syvi6K3ThOT8ul8VHbxikP
VgRa5a37nMoRKgIH279UUgxQiWJST/LeN9xqOuvrd/+etXmu6j+TANg/BQ4Dn76X
WuJzbnnCx2kTjRG4pqEweKY/fkEyzmS+2r50HlqgaBS0EWVu74cwjEi9B67GYE7T
BBQAQMbEDQLNwZ2n3nt9w3/bQxhX3mL9+O3s+WyrfxeCFFxNzYiB4NTWvSxZcqn5
u8Ve1hutI2UeusYNfCXUQGzMZJRMVCC2Cu6NbN8Z0rTqvid3f59Q5pbJEOc1iFPi
kCcKqfVVYYqWNzwaVOmxC3YnEq3QcjE1uLBu0wWG5TimtVt5w+Z06GHJXQgr4prP
GuAwmzmBX6l8muL4+woN9RmIrTTgZGl5ErcDqNm8C0q1OxMDsAe+Pdcc0gGHnSSS
ej6+C3cF+jtP/q2kfvGkBYyIZV2Ch/kjBBntCgc/6wTmjARg1bMUR0Pco/DQ2ogv
cr6rl1ZjeKGt4CrUAQvtII+il0El2T4a1OgMel9MtT6cdphG16zDjbjzy1UV+6iy
ZtgrileK2iq3lkHqtS2hPBrdv59uxNIwgjPE0WCQ/BR6lqKEFWdttSIwKRrLv2ZW
5vLD5RgMcKI9AQh6iCuxQcppB5ABjPzLd70YmP9EECf9qcQ8gQQds+Jauw7DE6oV
eEOb2uL2HUpG1aucVehru5ngI0cx86+z7mwE/a4N3zgm87bHroNuhuQ0ICKpoBmo
oHNuDibD92X4wfS6kCmNYcSjEbXI/OvCEREg07BUxEYddUqvoO6xJMo0yFEMnMUq
r6gR3m5+ehTLSIP+yP1dChOUe9gdsNPHKnsYcCJCGmJ87BIdSJvQ/Gh6FAaQ8sj2
m0oSOOrpcFgGsS929zezZ9lNl1H2qtA34eF+NC9H53XZnwt7ZcMKD1duPrtG6AUh
rRu6SiwOC7wCEUNIFv13fccYLq76My3Ms1dHyGtdIGttUNsTtLX6y6ukIFG9PlT/
dO7XwGSPukls1Ya00Dm+iAwVi5ip/tLtDQPEyIlYHQsJ+yjKKBWA//1Ab0T5qnVb
gBWWNadEybqri6i6nMO6MgJTYczDqYXbyEFq1+jLGCyOOQO95NKnfSSPZ2MjsSOv
isviVymzrt9DqgjNs6Zrf7oRTB1kavTeY01Y6xJ38tEY0wPvflIitavfu5qWEyfx
ToO/GEixTSC1AwVOF3WtmiRiSBm/9Ymv2W3CpxHBbnSfIRaaHSBAmqFEdWDTlIli
7Admxjseo2qaoJh7JSyEAFZp3qoRVmxzEh4DAEqB5BuMl92xGQOF2bsmdeFqimZ+
yMRvmxRras9mLV7PFP+lFCTQj0o7Lc1knl7ACS8NqJkGu0n0lmOcHrl0sZcC9D0T
I5+KXAt4yTzoUJ4Iyr657K3RJ4+n7pwjLsx8UZa5kRv14u+KqyfGc+r+XcwPm5N7
S1xWLqdgc2pyMq35+jzZwaWrcvPWQ6DToMsqKS/E3SLPSKZgsZFoSwpsNgQpgxjC
lGO4ksqtBw7aa63Kw7bB6u9+CgWmBmuVIDhkYeRv/d9QaBpZbfsNltjbIQxkhlOg
fxtgo1cAxy0cgImXhfGg3vwFY9D45w0aPO/slLGNLqB3/0EmZPeDX1uNFo9ciwES
d5APyG+4rRsUyiN01QleWhpmkMjjPirCv5AL8iGIyV7BquI5JkxxIgXmTp32HLhe
nzS5LFI0Xbj2RHhWI7d2Wia0Vhgw1sehvBV+nEQLBm1Rn6/HSw12fheSC516PdGp
eIm7mPqkYEUeaHk55/ys0zkm7eNjvvFkdoUBpXYp6ZLOQhZID3o1150qHSJ+k42j
aHjvs7r0v73v5tUJ7zpjCwBkVmUxaUmjQUUzWp13oMkhivXbRS6aCYCXkr3tv9OY
nOoZW2Pk+bTxQcWyQMV0YdwK5eDwqmOLBNeqYxjkiARg7WCZH6bRoorDq/JfHGW1
owi81z4TMCf1dhFCnV2dFaQalLXV8QJFXDVomjMX7oMjtRIISZHTHWJBzfjDovc8
mqU0R7IHNuUm6bLbsq/ubHi67En2qBX1KhVHdE4AASEntYCiSpIg81oxG8978VeO
mbcG6CODvFOhWjB0wZJHgnnhCGXo2/tSCVZ+7Na08z3ICDn6nVg5uaXoqAyNjtCk
1VC1l2oHC614cLcV9bskBBlpZxUJHUftuUZBxhPROK1j0ovdo2hijKOE3KQP83oK
N5uuO4PjOj+vlaq235PP0V/nc61XsN7HuWTMV6Gk4DLSPzxDLsMZVHHz3IhJfLpD
G1CTq8oBm6Y1CfBSdID7Y+RRPclJf+sFxl3uCvKh+4dGzfJ1uUjHb9I9vbKDy7CE
2KdsVk3OhBLB8lizpkLXJd5+GVF3LRe34T9isnJf1LF/Y8Yqh5ZnEks95V8wAFWQ
m4gwXHWmBMzWc40Fu9UdZWX/iqIezfwYdr6L+gmWaO2Glf2DW9OxBAOpfAM/VHkd
HtLw8StxR5jT1ZyU+d8eopi/8IU/8Cj37uFe4zJ+JU1B/fa6DVFtfHfjNVV9uqa2
F1eMzU71NugFuPlSHlfRNvTFjIL1Hc+/tXO9Izyn+eB7+8zsX/ub4NMa/Z/gW4Yh
I/FcFleFHYNo8uv8fK/y1tqAv8xsm1XejYfufA7nSuRkmKYIyVVI+CK2UVy+dbnT
JlgjU8pDcsuFpAHGMLelD37LHjVKx2alBjxc7v6dIAs9kIGHJqlT9ep/TRM0WRkc
g8Juwrf0d+/pHUh7X206pIUxO1m8QHCGR8Djk89oHU3fbDR0/gA1xpzD7c862T4S
AAz1R9ezZZ+PhPG3niFCsonEnFSdQU5GgklqHZgAJWbedUq0JzP6i5wyVy+Ccrlp
AR9XrHA6Izts6Fk4Eqy/jR1hfv71vrMUMAdgivKviG5TfkBPZ7tPhOw1sBEbRU0H
CQZhgjz64HkSiZhbr+baj6EUjyIuZZMEAni/LsAf6GUnSHoTBxR17h37Xe3ajOUx
QZNinCtQ+CMKC/Z7sOIviQ9p3K61RkjeowLbtkkfKhSCJh3AyPi2hLlfq7qd2+hG
THE4+FiEPYS7B19EINnofM0Wv2HuyT94urDkCPEiOJ/iFGfp2YhcgzvZAtHEjiru
k/NhRaO/dtoF7kfTsxBi6KdBQuPJruiGk2QjlS0NKIBO5oF7PCiu/87qk/AWIxxE
Vgv6140I5nIQJBpS+Oq9fALKJzmJPjmfz4KGP2Fevx9LdoqZTzg2HsxF0klWe0pb
LJz8V6C5O60RgkAIrdU4gBiURMW6uj26KwgqfYgEvWDR7urEKs2etkwyPUSYfQ0n
pGhoFgMv7wOh2G0MnRCZ0YHqrju7RTdYv88PbEiiLV57wfKAC2B6uuumnWBJ/8IB
sEwIvffAV8Dzl/sc3w8TDk+zrfXaaW4dYW8w6IwgTzRTVssJ4S99u3zmHmQNFfz5
QIt3WYys/qQc7eDDVYGY8b14wfbChrBb0ht6Actxi3VOeALZp3Qk+f7aZ9gsjkfJ
c7SQwy3pmsX3keEauPs7kMKPKEf4tBkih4fXRzVQHNAMya+Zj+wYEhBjDlrSypjk
rF3qkMCI7njoDokSQlwQqoE3FJeAiQx3wRTyYqmy3Au1BC1du4meDWzRw8fBahvi
NRDn8hyl9axHuy/Gx2lb430h2Q8dKHIAEI33m9DUah+wqSaYW+GTFihFHNQLQVtV
UMZiYkdrdjBVUJrGzAg9j8NiuZf+H2nGb4wmlWg2zaPOzzHNZ+IfW6IpUUBmzxqx
VXuTDyaZr3OkF20gnAxyeJO7fjwohTIXgKT+44fKgIPXggFykwNPz5aI4H7x0V1n
j1BWpu6b7d1Bj2f2P0StTT+ipqmPUZm447qZzaYRyZdmsYfoe3NBhHBzVWldYp07
Pvzg+rGat8ulEEm44zBe1SppyJu5Z/0dc6EJ5w1JLokQ+1eeH6/y6/z29lY2E1sz
KCOMaMsMT63PqPDt7Z0StMOtss/7a5hPuZwdLkwNXvHjg+9s9zGHfxAczGi8UFHx
zYFCxZ+LCvT+DslUUuzjW3B/h2NmDQPbIcoVUcb0zbZDq7APZRznblmK/ERWME29
jK2LTT2W67OH/2yKNcV84iGPt9ImTfiIT/DxCcDDB+ksSciObn0oo3iFznbecMmL
n2WTWsh//wu3xT8nDimpYrAz1at+4Ayzzp4g/haHPKuzyNDI78NeEXqcAfzNdyJD
QRozA5KQ+wEgVZR3Kt5oWdHFJMPHGHXA6T2NKuOy/HcGgpWesl9+4NIBXIkdu+9D
fyWsfPCgV7YwVivZCfLQMe+IYOOGs2cYPbxetlracSp97jdk8RLGpzGiKx335Q38
FwyI3cpTKNj1BkWjiK3iaqyIhn8gZxP4ddQIT3uaYt7q82zATcOXWb/YeHkr3Xn2
2783MBdAkZ9+/UfqHeu1sAG4Vsw/CGtBBMrj0xNuzGKVHPwefuP8V2YH5uV6ziWf
dcmbH0Vi9a4RgLt5wAM6VuKOro/jcAOEp2OycAgptq5rpSsGYQwF8pT0JT4E9V7f
2CtcN+oBvSujrSInAW3DUu677K5SLIyYt9UM7cQtdFVJUhbvuNWuc1ZPEYTTjEMS
vXISKu6nfKnHSu4kFLUGcRuupb1kbnNrmkLGbQZtNQlEHhecGs3q64wuHYWnc0Aj
epI+Gbjlg+/6bfui5ymFuKKdm7DKkMrhRCQiuXBcZPG6RUbC3+PFedh1Ond4slGC
DqEyJqK2v06JdiySZVX1HG0rG9hzQhF8o0fOE/LcaSXd/q2YG+VA7FVda4KZjmxb
tU7Lo9gnOz+wZvZgLJffyq3rNxQJg9BqF0Y0/6CV6UHnif/mQ5ocByN/ywd387LQ
xYEJE9Ix8xIEiTvRakc09cc1GQLKkBrPTrQdy54MqoCL86kh867AV1qqbHkS7jro
u3b2QNdEp7UwYf26eRFQIC0EXcNMxYi3EyLSrYlzzD02uky0UGsDWvohYosaVvaE
oYNNtj+BvBRdDeJItrIHToyD/YU61icpxy8TWYeknWBEwJ/BqVFn5UJDmT672c4F
Ulh8gAVLJL68FHL7+SE49XN+XgBM5Wv/WVg0ryCha4aJqmqjrmhTGM8fie0bhMh4
Tlrf22xUrMDgG8U8HSOyCogxbf5izo5OQs//q6BqS+1othr6itE8Ukh5DxxCmyGb
8ovXvxz7PFJNZ10eNhMXB5MOdsDnmay4AMGi3JMfWV9ICk7OnC8EUoME7rVLEDwH
QBJ1cHdP1QEhjoLm2s8Qo/C6UmyUR71bCs+hLcijqWktbRRkz1xOvy4ZiySc35gl
bq9RqqzVBcQkbZ2LHsv7LYYLu9od/FBBf1gjudhYZ8P1iGThBW32swXCntILOsuM
xQUnheZkL4k3wqTGxBL+I84yQYqd32EadtYqT16swRDHhnePWN3KLYtRGFB1Fwq+
//QhdVll/Ng066E4onTInpYSmnnMJuQ1TFMfcXpwoezrp+qJEELvBLVGv1DLk9Ve
dO74/qenhrVwbIJgHRT6nFsoWkcOgWcWpjR5wwSnr9mKDuZz/X8G9erY0VB1xuUp
Ii8qNQ08QDzPQb/5/89FVDrSu1PBNvjnlswIEgM+VMufxQ8Vt7tAId/W345deTOy
QPKkVxaDDkMVZNXim2R0q6fbBCrhqwlRsggQG/DpKQdYR6YWxWHmWqLs9J6OWIzD
vzoR8lAuVqwStfcOz1D+64iAVut1qmXMIkLE7j1iYIU5ll8n3z2B9mPv/X5Lipr0
gDLJA/hhBSEUhgMq8DEkxh3ywpbRauVKOzS65BLVulBt2TFu4ztPzwkmim6pemwl
Wogm/BrKJb0gPbhEKBHcH0t/bfPRiJh29VnEuE6sUXC4nzng7zU1tFQZ+80av6W0
nrHR0u1R21wnfTzJpFOgps3lrFa7/IVcfA/uIUTAeJxn+5D/GMwjbDGVjMNyxxpx
+M5YiqXZwYzSqiYtk8x4XryJHgAlvDgyAKtew43+HZ31xphzy3XYatKFOFbl8XXI
JorRsihKiJOM4fHPRyQEVgYXRK08vawvUF69cXLasmIjKIABGhditDUAfMmLzEnr
vlMjOkhlZNcNYLjQNeXIqtTtDxSfggk0HIpVIaMGijr0fTcDXeQefKtJxMnCXafH
es68aqIwBYXNmrhT7OTCAjdec8HyIT552qvznIoetomgBtK7uoWwIwqub+Bk9hIW
f1Mqrx7xisYIdUamYYNd8Hmq7oU6WJI5vp9y1ePfa9dRyZ3d83vKuLaSZCschGB5
3KQ4c9GeRZgREkD4pNhpNtM+lDE/BBm5k25Bgt1pNzQmabA9MmmsQyiS3PnfnGGA
JU1oKSqP5YCiqjtx9HyuVywpu5Wk37lOmn4+s21yuNCB6xLxq3jXuqWDtDsa+Vdm
ulSJ3tNjKN6LifpUmTvylBW1BqCIRPN0ma+twJowZ9HkuNqzKVf1qnbo+YapL82V
a0L+iz4frNYQa38uPMsafWvy0IE7dDFv439sHyXfBlNf78aNzF1T4N2x5m6Krndd
NivRlRDSykbGK+LZeJ8nTlof+iag5IbtsDagnNOQU5RwIPbm/BwSrxMVuEhb6OUg
cnoemPgfGbCR8c/nR48JrkejddV3iW8dyoHkohG1GQ/swtgDevvkwtMD6Qg/g/3X
fsPIy+BAYDsJxHZu3DJejnSyL0RcIztJYFL7t0QNyiZ1YWZbbv+TghJlpSESFKiO
YVNtxCwBgcUxILcpR4w30SCVWsyFYbj67runIoQbFFqPPIqUK4XVATHHMNGWHUJI
irLHqqTVL91lcKb/tgX8noLBR+suMmrT+WGKlKlhkr2s2TUzHrV110Ftf2wCVWZr
QFaZjs7kEM5z8eu2sPU8+1qOPnjzXLBi8Tg8WKOxT3EJ92j8Sz35p/qIr+G4fCY1
20o0z9Kq0YwOnQ3H7YdqjG344GOg5/XxoPjDfMd9F0wA6ojK4Q2mvYwQH6HUROfw
9Q2WouIURoeDNfC9SDybYj6/Eyilg1EV0apMgphQysdm11YvuAULXw0D2DW59XPc
+jYrcpYQ80g4SlP8GA9IK5Mr6fj/W1NZ6TaxElvXl8NMoq3yThSzMlVgRk8QqNZu
KBj/Wlg/HCnZz6ZsX9yniQCGCztXyB384/5JFk92JxvvWlw52wOtPnapeksp1p51
EkiMGLJNRsFQamn6gIefd0ZXbKRG9/yShiYsiXi3YNMzQ78R+HQx0MKyj9gUdinb
l8d0X3vUHaTnZmMIcsrzmXfZjdOl5oog2WrTwMrLEh9+N1ZdJQjGaS2xaqiF3Mcc
Uyjr3LWdpjKb3nhg+QAFUHzpzlkLvTQY2gfwXS9nSCBthzQ+eZoCFTUQHNr4Hyd+
tlkEUNOF2Cv9SM/zVwBrwm334bFICINnBbscNSzOaaCyrg+C5jeqeyrCFC/jDLWj
lGzDSLcH1Pw8uTZUORq5AdTiPP0lNtgv7bbPZ2SMF4BoXHs7SaBdiTkbzAPINI+P
CLP9JvqE1C/1TbTeuSeKyzUvSSSCo+bddXR3KBTiS1u5e7f/krHng7D52c/Cpe66
z9s5DpYosbK4+hy5cHmUbYrz/r+ks/NRY07sVULEaswjGNEyFVe3XXKWEta/tYIU
tQai30F5rhW6EsrM2yguyuH1k+5hRXkc1kG6bq7239oWmaQMGNX1wI1PKjBnL4yQ
33QBaKSjoXlmiBnkiS7tLpvfojmJOOeT3PWja///225uk0T6q1+l11l1IaIph1Kw
TSzrDVPdjusxzEGUekASrVPbjxEP7eTklJ/l6cTYn/eeZrqjbBzB/sRrYS9RvPFG
EAQn85mYAqOtX2CBBxigJTcwqnMcxPtNPK5bm0Qd+OI93aSTxz5oy1gAVkVlNvC/
S53YKU0ZD1d6LG2yIoKA1EHxqOnjOGrhGvgd1bLHzz6nVx6VhTATKoz32IGPJ/w4
nISWYfom+tdRMMT3sJY1CPPCEH5jcxso0WnSzkrZLnxT6AyDxYfPUWwhmAB6P9Sx
yVR13Ujs8lxwsoEB3EdMJlsqjLrx32FLiKEpea+nzN0zKhtr7oNUn2+a562eu7Cz
ZI/dRdtZZ47ugDwBPoF4q1RXBEJ85oBYlmJd6cd8rbTBnn2Omg4uammXbeiLtvMS
nUvgRS8gN8qv6NfMm6Joh7U0aws2vxawE9u1e/QIfFYCgVjb/Dh5tq+Sb99riZrH
3ZJuzij1zHGPCtqrKp76MT155uFc68nwWe7soawrE+jLjgulFAF7QFmGHX/1CW99
3F0MzQONiuAMptI2DBBxy0dLL+A96FWCLzQZDrqG7Endfdu0v30ApB+FDQGxi6OA
sfH3kJ3yROt2ZSSeziwkswem+aZpPUSYnn3QPiFhmCO82482Fb2kOPLI6+/kXI+j
P6fc7gI+EP3WK2q3HIxQrLfFDm/Qp8dASLiaqbZlM5ArvMpGzoAoSnmUSRYAAeFS
LLXJsXNqZRa/tsARuuft8rNl3X9/PEFJd3G8jQFyAxsxHnLOtQGeAj+kWUfu7deY
8SomkzcUquYHlfcXbvHxiNuhnbAZgg0OR7VLSIJKYHNCx92MbPxcg9nigDzEkJD7
El8r6VsAVgEuRlJjCYl1KDBvpzIiNp1CrQGDtytZL/vGNyjcOMYkBT7eTy4vxBJN
/eMyvNTpgAcvhTxs7vYIQYHSPDVougZZzKUsC6Y86yP3MfpWGlGIaVwMgNm3VCgH
MYkHtOmCeSuB1AipcoXt4VS2YEp5QVLB3dknquooj2HsT4WWsqSOuBgK3XKt7VUK
cUQPTbz5U5wlGWifyTS6Ygvh+zI8O+FtS0PPedeC+pfwzgkuUhkGQgiTp7DqiCeC
r0MvZPvm851Dk9Pl5dTd4Pd9yAVgDy5nEM4nkyn+JSBf9Io1evoJdxi4q4XiUi61
i9lvt7fYjkwBkP9xyobNOkyreJUn5cjgWfgpiaHF6uqlch25D6c1TyWYT12lTOQ+
aOabuk71HY3di31tCcqwbnA170+goJn9LSW67PCji83BRGs2lz58pPZSxsg5Z6wJ
o+cAWJlc0zoW4sjzY+f4Mq2PP5eGiBG/5Ey09Q6VquwbI3Y4HY6E+HFOMuvId9Zu
ExZuKIt1T5nnAuI7SAiyrcF1IakPwPeSF6M3dpT3emKMlMRUQZhxFp9hYAdVsJOO
8FlFzBhUvffjQlLb5O5VHjXpTQFQOxkT8c3V2t+x7dGRoz+KpAd4cOPmkovej8+V
isQOwWZIOflQPvolVbvRdGwT2k8m5jj+ljFhe48WIpjvXY9eDQlJzHYKMDUeYJTV
UqN0w3rt38GPw49LpktMvN2Gjf9FBdpGeid12M12epgwr0lLhYaNkcDkwYsig0RV
H0Ywctxy1r7cJrUiJVLTyGCvRyp+Jz2YtO/1OK2spf05B8/ClMItMHSHLuJNpVoK
znIJx/TmdG2ccbaJekIkT/4xEQfj5EwTGRxlYWPt3xdVX/EWCpdFRLFk59TSzR5R
dKNxaMAbXVgv4UfmnVjTmIFZ9D8lWMg5E+LZC9qbw4gNgh6n0FKNBBl6DiBQQaeJ
evvjGqkh4OdKDRi6OSyQAcQQocH/ihlaWjf0k0y6UCMw257juQx3uYKmu4ecM4dN
bDy9lWFO885iPTBRAt+bGg7kR1KNdozIoZUI8jBgcPCB/MGkwnPBjVPNL63xBcWl
8uYtqY8myROB7Zr2fOghLAfcKnD7mWVAQqM/wCOqaufrvJhO5tleqBZpny4pSmYB
npYHv60KfQ/rTSQSiJCXbQfvUYkgGzyIJ1BdXbk/e0q57TDw0P9f8GMB4IKxMcCL
OJZsA9qPIq6gYy93CbRzi7dBtc0orB2+h86vSRtEA7Veyb5gEVIgz8EW7etQNL4C
JY0GsYjpWQ877cfYgm3OViYZpT/gjTrpsSzyNgUtfgqDWBmmxHEq9GEjamPuXA85
GFI98KOeUyLqkAYsgt1riZxmZsYY0RQ4r9Ey8pwHHgACCQXoLTK0k7Ooo6GQlE0Q
+H7EVvWPptGPDHxzEmbDrAN4brdNugwEOhlWcqsx/9w+UDYASUK1kspgU8dQMESF
cJm+9whvYBc6B0zUIykSs9QeD8QVAB/+3rK27EsbUAA8dU6KI5WR5mTmUXgBVMnX
4F8pinC/u3QWqNxt2FQOt+lhjlAUnXkJMGDLmuN/2FAvGsaH9R7AdaHlYd1VdEO6
6AMcwF26hSqIDqe4f927+GTdfKlyxpxuff8Nj5gyT78EVO3olQ1QefYx8VouYv1Z
cSyPwJLEXKSX0RLVU5CbkNzPQHsKD417qRcQN75ZZ1A2KrErDkM8siFxnMvU1jAm
dM2LzPQ4BtR/KAbbTbt1mXXyqHuk37EPbVE/qG69mPtHYRKOhaaxhwXoDLafL+mp
rip70lL26QESmmAXy8yd2JWz9w658r0gynUd8oEVF2M6zSgLr9SQyokUXuNslz1j
/QAAl7h34f/1X8pcSnGHOfvs3wZjSyVPmk0wj5LYiVSJvLK2qCu3w39OIfmOVqFM
juSUzd3oEc6CWmuEcF29YLrKFLcVk9jx88vVVKpsZThe6RT5C0EOxeAArWnWBQpV
ZJvoP3C0pWBDmJhxd400dyhi1/ymsBhnXz3vtj4/6amN8A+sQ6AOPkfYmeu2EVRA
a1rnMnGehdNCRcVVWdSpXHO+GCdZD+BzpRo2pHroZguf8z5EBzswj/PyJLOx8JCw
Aym+MEBmfDn5GRjBdnes2M6mr5ypUL/NDw/YMM6O0/njk8Tguk/JjggeAxtIeUGA
aty13HR7b/KdLZuqiZjF/I7Yeo6C+bH+fd+difUVZMg8XFHX3ROu0RIq8nakcxYx
gBQzDbmod10aXuBaA3okF73rf606Nw/LK9MtJmIkTRq+IRbxX0pI21vl6tCn4kaa
8ZgxaaIfcTvlXWZtojOr0yQX6BpaOmTtpfuS3sQ8m/b5wYbFggmeI9KJNDlRSpIS
TkE+FNhmF2kia9Getq3JVKXSR0ldGDZmj1AOJvVUUivuRzr2U0zlTgDlKH9zkcss
JyPvVaZ1YvkTnecqRFQoeBJhfEygrQBBAgMVc1epjQvANP55DpD6GhwRHmMrAu/b
QjjkkvUkeAr3Kr+MRpBW+BGl8WXR8yVb81Nb8jq7X2WapUaUfNIrNETAU2HXAS0C
HJlJW8nnehPu0Jd3f80ize3PudSzN59xsbmfW1KIdGiBCPdRTBaYu1JkdvTUfcWY
ejBx7QPdScTfvPnNXQPq9EcuBA0NsKzas9tQ2YdhZopKl/8HtXoNFl18aSCnaZ9g
gBVmUHq9q+U+Zk39R8qZnr40pX865+5mqOvmTvU+eSj/XI541nO4BKTTqYK0DcSR
dOHEIQHEmnQ873qI/rPbH8sC5eqBPPXNtG36rdOmN3VO9+05ZQ6BADjEoywf9ysD
upfUUDHD4I43jQPuzE7HXwZDrmrZSkzaGH3zRRFQPpKkXNsmH3o/sDV7pcgAsZan
1SZf7CYG4bBc19i23yjLu4rfLxYa+RUeUvHd6/FYtp6EIQh1rdentmjMT8rtCnnl
69QgWIOyMBK+qjheSuJ2aDo74PRFoDBmazMPBWzdadhFfBhhjfU4zSLWFgEFvtrd
FbtL3JAe7yK87zPKZI+u2Rbcz5LCsZmPI8pNA+o/N/QNjmH/eK+CuWATxjD51Qmt
2iGAvq1LH69l1Qav7/QlXwG0DlYfDX4xCuUwoy6AsZmAl/6K86flF4fl2zdhv0rp
wj1x9uSh++NfakdY9Cqpv1pTyPMlfi7YgT/WG7LBOnnEHIWBG4r+wsGpCmaWKNva
XYPpt21xOZ3NxjlykaVCXt2TM2i1rpkzCrFQAc/uyDQAWq6/nttTJEY05i/zTfkY
e7BIUubAUmgA47ueyXjFWy4gSWMjN0wg//SmP8Eiv23ss1PkuEAc4LYqV8jxx8ya
jkyH2B1g5Wkdq+gKqr5ujAPRGnPAT1oMBcmazmmK1Zo3m6TLoP7T+gVIivmBeisA
/UiGhXEGcVgparNcld/KhviBghGtlhRqhagF79LUGHwVTfUjaZGQqljd2jKDuvWK
j1i7UfkSCaPgnsA93MArjd99RYkIRCme1+hiXgey0Sh5sC3XMHfJf1MtgKfzOy6D
414gYEaxYtfh6bK+e9F0+dUt3hSH6kJSBpyWMHi5Zl5lrNdtg6rLWci5/8qi4DhD
TfAG5FVTp357D8YFA0KWhS2W63227ldEIkoNgTKeBJIpoSbSCA/j1MZL+yZ4K2nU
53w5Sk+aWDtLqm3YKtsvew6CeaGUzS5WbQ2nOASXGeN0xaLoIweZRyBURtdAB8PI
VWlVA4eFoUUWjFMgAOmqgdk/UruwjxeEv0zYFSt6skJALfhSIRHvY5q4PTDxOSUw
lj1VN0wJyt9K9XfDtP6se0IfSlbfuRNUlnjOU/qTKLWhWm5/s5XaD9sdvJReS+6y
ZQ0TySRptsFL75ru3NCRyi7qdfArDwVGCgFawx8C3d5Iu6JKNxplQTBFDCnjaSvm
/kVXb/3UaEIFclcwfYll6gJFzXVrcZAESsAHXMMu1pwWnhwwfZn1ippEBYsqbB3/
V0YROrk9UPE17R/pjHMai3QbK07SHtp3FDzsh4hM+M8XESR1S0qnQo0ZSIDJnv2w
DRfaSlYCl4pjN+CfFE9j2Cd6mIcxntAT7tmaYEViAIv9GrnQV4XGYjw43vT+TX69
d72e+y5xeLqS07gIKvkTd5j5Z7UGIj4pmueIel2JsgbD0m5sDZ+8mD/uhuJAqhAx
hgm1lEXOu6NKxu5KTDYCi7ppoCcM2DMFxnp+wQ7eEH5PKMLXTMxlkroB4+4MPaKX
3/BV0qPA2TM+7Taslot36K1gOpghTxdkcMuDP33zpKeKtYRXL12kK1K1gPBf3o2L
qiH0YVaH8emKPpRmf242U7RgMDsmkG9YKqEl3rucdbOotuZ3KnBydP/l8ommWLQm
9MFRQDzk0RJpMWcuOCONkewLZg5orYQXz6X+XM76uPdfIKuHcsbaITWKqPQmkQUO
4C6PMJCupqmnmQ8YQHdocCZh1pAGRZKbbypObFqJeXfyKyrE1QdNpB3PgTh38UH8
r7wbiKSmamjbUVxjXyGAQMHXLcR2kFKjTk02MqZjp+Vi0YVYm0J2w+8W9pL2RO4p
cPw8dkStuSLCaFFU+dN8cj3BX3YXLkpeEHqu5CGLGfnUSEK3T/wSZ8HfPnohdG9A
hgntabVtgFKHt/qSpM7ZQuO96oIRcwPcJesCjulK0ky3GvPj4IVtddm+v7k007F5
g2B/DU2407aAkPYmaIVTqMjZspDU69ZNXViqh409RujFdi0Aig0PXYnOyXvtDC+p
0Akk1Jx+DxuWKq7r6bUJrirVFh8Pfjykl2b94jo2Y/npEhj6eWXp2RJvAELv8sTr
P+Mc/WCZhe0bENAtu9Yz4MBVOjSw0cTfEaje3BSLbByzKn+AM5MRrqiMHkP3ud3d
q8sSHyDn55xnpEeyRqFyPFcb6ALMs+cSqU2O+b4cpHorDr1JjZf6YdUXQwbRP49B
qhRG3/Fk9hVBGmfwOg2Q5wHomZ0LfBqqK6sZenq+SlEg+3JOJbGoC5VOqUhmhQ5K
V+aw/x7J30kNN9vDBHGI/0Yi8Er7subQ/cySQTme2P7xoVz3GKBvfA41hXFETiPC
nl3wrU9+Ku2C9sxHl2p89+B5+RQggzQXAOOOI6D0xfZpPePaSy29hbH3B68q+I32
ZGEFa4cR1KLFri8EcYcRxkbWXRVi+sf9CfBr4E1nf1CdtTCvKuIDlQolLT1segBQ
zxv+RZgur2Ywj7WHJbegyQl3twCJ5g2NhbN+VqoFKmThpD6Dd4NsvMl4jFztKxGv
KNbMw+U3NknaTcXKHfWL+iB28jd6DPY5wAVwERlldmHa0Ij605iS+6Oa1FVU6uZ2
gVotoxc2yTMFQfPDksoa+sHnL6MtLKNLlX/ZY0oDd8TxZMUQIKQeLLzoLdn3YQl6
xVYmedQQXIMY0ox4YldiRKMIFwIarjDklgyFK9ZirFHItfjFJnPowqgClge7TYYk
mkyxg4bPVBpDjmXwwBGFoJvDZ/JPUJXAmEVKgNXpHMZ7iEmPetW8xbfa9wAFpief
ABVkZl4dHJHBDJlWwx+lw03bzPYLj2wV2TJrNnUSTo3ksnwJoNlLolBeTskxSwfF
oyZa1suO8u5MQpyqdu3IFkFfkUZSdh3+VvHkz614WQOE/m7POLUKN14rHUt+zAdg
myvu3qq7uJEHGVem4156BqMxseYAZ8wmsooy6VPnEU0Zs9GfR6zv+Xr7hmeb1GZa
IBHH9aiB4zXx5WNHlfxWn2tbvioRuDrhGe65GIRtZwM5EGbWiEKHz2KF0myb+Tlq
PCSItCOMuYO9u/000m1E7ofV4XP52bTaHMx7K4UFeU18GKtNgPCPp/vICPyqg75Q
iR9sSlCSG9+fFiPylBJb84ZdgSuC8MlWY6/uznEUy9QyVaWFVAWynGip39sspqM/
FU+tPqEDfwe1+Xzztl7pimx70HuMhLn+bwc6FOlcKFl/LHyDHHBSvaOS/G07sYEE
uHgeFaVnyKr01nRCHO4rLESGV5gONz1XrIL25MczrpuFWrt2XgKEJCANQ58JnASr
MEuEWilDgIKHXuStLt4yr+iv6T7yGihJGHPB5P6+sDr6O+d4cCTSMx1nGeYZyZ7M
t8GvXpdf1+ZdNCqokI9plylHQ7nK8/W8vxsoLJCv2f2BycyXAm81CbX4RWJkrmRx
SDpZVo3OjzuTgOqhHafyC9Q5aZyu/FRS/n/SZyg82uJNqWugOV6zadZEetwwMc9H
IuevTqj9AlnOEtzfGezMEO6XWDaAC1oASNvqlE/zilS355ps46BnTHnvn4WGJv4D
XeDxCgcSvbqTX2TRWikwJdfR4njQh4gG2nD3FLeJejDrdaaJyEXX6ex/z47um9W1
i/rgzVRpJ0/xUeY0VklpzmB2j2ZAW+f7+yL/VWqipZY1e87XbznZjvfT2aacileL
Xuy65tW9k3luJURZpKa/HpibELQXYDa1EGjDOG1zLCX9XIkgC+cVKlDkQMKrHKcs
2gxEo5R9Chrp8cir5gm04kc0RXutaY7oIbEr38dp1rCfdrxZPCO0MlJM+FO+GsPs
ZBG/pALhOs6sxzv/Mb/IYkGMgchz9wipmNV5uwuoEdhkQ3IdkT+LbTqmhbE2+7mF
7HFdJhCI9k7cUliY4JCPi7kiIr3XqHIzGaFVi1ziQ2QNJvfK3BTfN+mO6mIvU9z3
Os3ghMf4R6q39e2Mldumw59PcSf8UVMng7keOGxqCrZubqL7SARuJxEQS13tKeBo
uXj88LG0KCzxEfwzF5HqbxH6PwFEpiO0SpX97/WUXBG5mwbtVwuvvOUEoSgt8dDT
KS3MdhE4wnsTTZG8K5fyIwAUzi0l2HDa/SqZ5wNGF+gD4Z9SbfdXPrtIAX8Kphh0
+DyXcRTZXXTQjdkryDPLX4lO/eZVx4X+a8Dj12471l6ZRvK2VvAF2rSHB2OWL8RO
e2j6K4bAdKNDTQD8OGTydrNFmK7jIXs47f5yvaYnYkgQVQ1TKr3TG6+LtDhxJ+qe
xAPQWCIpU8u8JEe4vRgXBNL9/HnYg5+0W7oEr3F910jHC8+SyuqM+zkX9j0Dj9J2
42WdVfJor756iS9FNdQvDbpw/uQGizIxzSrE5Zjdp//6+1oHyaf1HVrKanZJjbC+
oqsqnY9QZHXydB8SkQgWU4EsQI+46Na/Cyl4HdT1GAWI4NtcBN8OOWXlGnuBGrlH
qiL5x6/4b+rE/rbwtLEuzO3aBGyWdSpHGoPmk+PE31x1eCqww9YJLagodtAHED6n
fekM9qCxk2FpTQBfh5iHarCV9B5PRbJV7OzZ1eC2KU6r+9zhGrKJiqy1z6Q0Jfj0
6bll0MklwrPOGJ30BB8tceiZdBXT12DjNIfsKRdbDq2f+iG6M/Wj4VMhqm4X6EyT
fBNn+LAAbv0DEO/Fu9NF4A1IYUWIu2730BeBtZyK9RTsF0VTwr7I6tfa2nt4KadU
wEy8rNFK9GhapT24KnYGAKTF60uTt9gP4CSTHmgUUJfb3QbmFZBIi1d8f3qMwL9s
srBK6U6mMlRvu/BC1hmng15bPHC841pyA6RgF4H17xplGubEQIf3SOuEajCEY/ha
8iImPVafesgz2pP65TTM6MYZNM1h36AM/gkDZxITcxgKQwSpNVxAmgbjlG1+n/Sj
4IUww+6+0MWkFqH/OgUopSl+qmQsMwzfW5roqAaGobPxZWVmeaGj2AJHtjIZK9fE
m10i7Y0WMTP9Iv+4VWb7cJo0vCT3QOChgsBV36BzsGxthEZe7fY2BuB0V3a0OpZL
jKRN+M5H9H6bNw3b2x23x8LgJ7w8/UZ5T4LUOJsphqDCRJBzjhVjo/9KjG25ZcZ4
Bgt+EhmJfEdnfK3Dhb1Os4BXwMvRVJ4J3STf89Fa0tlyQcfAllL4nOp6ItnXBmSl
ZJHXFhHWgmRI8jcWAek2garYWks1dfaxfmewt+HdHAvOXeJ5rQgKGe+gNI/8vEG7
arRlWyL0wZMeXkHaFGbVE42lnrh3Lk5SpULgb/zKY1sChTE6CwhzdDsSgJpyVIEF
6EtxhkhS0hyXudugyWQzAIHGycDdnvTuQ+KvaP1fsXPyu6py4G5UAjoKh1rPjuNH
sb0SxGi8ycAaoFZk5cQjstjegQp194oRs3W2vt5ndegYuyuxt8lP/2/ALwmntTMw
Y3H8efN0CSvSY2ckXxVQzZNPwA7qrLKAAHrkA2wBUl0oadAUDH9KzfrlHycUYQQb
gqbuFthq4KsKpMGK4SPHBCuY0fRDzXIo62Tk64jDPcE3FXQbzJY/w0x5nZXBV9SL
QMyN22WJ6QPPGEzxnySEnfIebQ9jQrZz57JRoHDUak1YmMAAJcpbc022a13D6wF8
jhok92kTD+xqQW9D8vPzQXMG5I4SnKaAiS9NTJ8ugRKhDmwCLrUJ+ENbm1un1Amh
+ycSg+aajOKSfiDuurG82vPBAK2jEV3jUazG5LGEohqxw0R87p1GO5d9CsLKarl3
lFO6KQSiE45c2L1+CxW4I7aA/j7tUyJL8BSxA/eYUqTwiOpK557rA27G1dWg6Kis
OF/cupzxijbxdA32r40v7tS6UihFl8caRQWFz57/UfYxttS5GgO5MXvMQsLJD6MW
584S6BZQ3pmII/sqtd7mgrdjkwT3OG+gSMPnGoSpHAdlIk6HG7CO61kfIfm6TInK
fJxh5QtJ6AzNmoE6N1UDF8kUZPUBCTqUGPnd4fZcig1QsBgtASod8cbpxmWKuXB5
NL1beLK4ce39vuus3c430v8rGAjJxVzX0wzv+iuGdQbfGeZBvUMbyaxyb4dt4T0z
b6nW7z0UHnFJ0xGmOazNlgajz4JUiwuoFk3IAZUdwrNNP8MVYhEc1wvcZtLyKyrD
4kxRrNfEYJVkseP6yamJwsD2uqiUswjsYXQGDGAzw7fJf8+YWRHdM5nZgg/sgBMe
74/3exm0hiDGIA2Yt/bx75B6iY4tbIe+KSKWv1SZhGqZi1Z5q1lJOGU4CkOnITm6
/jgpFOdaMydEps+htHu/hi86Cx/Q4p4gIisRaJTbKWcegRoSSPGo0zdr50BBY49p
lieUnKP/G/MQNSWPVjRGnOWVwRLLP5fWtLg1E2/kwO9G92MZUXxUQQF4RSo8iZXk
7K5H6BrfQ82ywSjAfMhrmHwoSEniFkUqLITynNNUyW+R11eKK/lFODir1yhWBAeM
pKBmrbnTUMMpBBtrUX3psk9/Rn6Z3t6wO4v4uNhIFtqbjjE54zdsQI1cHaKAq+6Q
LkpjQXtjfnHS8cuqwpb6qxgMzFb6kBX6MVSUBshb4m+sEBMJ6w8k8ECuD8+PeSuH
4BYXieSOtsMcW0rHjR+MX1TxDr7mIXSsI9picQkCNmP9OHnmmRvB4ncwNXbz6zLX
kfR0OQFj3bm4fBUQJmRBIxXJwSjYi+RfXN03s0i+mtzhtOEkvDYGgZ6eJdq5aJzA
JWrcdUA7gBqaZ2ajT1Ny5ROYDslXaz1RL5TQS6ceGBNV0VNhVkaTbA1srYYt51By
MtSZ5/O8yCpTspKIc0si1HCSqlN7P2ix+hiQ9pkU2ow3tsSBuqAWmAwGnW7HInN3
j0MrCFKItb8pvgXK/elXneAA6mZ7zUVXzTZduuBMZSpCyVwsGA4ssLL/GZ5QdGjm
oevQ4fA7gOM6266+i4G65SWhnc2bnoMViJq703WwwG1YNd3BnK6VM6DPBzhCc9w/
SFbeTHcq+TL2dFhnK5EYB9AnB7XGvmG+qc5Z6XrcafEvRbkYE9/4AGgu7+hBHcMn
b+r0Z6O62+u3wXSFIvEAx5dlkxyBTbr9Mo47E2FEJxHnZn/lVQX94SQjtzRtSzy0
0uazuQx90U39WdGwauHlVLJ6B9seP2kKwyv4BXUtaJsCTx5enosYqp2nmkYlFhYJ
IRCWmlriyBnvaucf8NWTE/Siv6N514CZqj+BWNp4NoHqLuTJBF7JijQLUZdxMweV
yel4AMAwU+x49wsq51M9DwecInLf7Ou2XOn+zsjy6x+zSjXAGu/g9Pycndc5aGzo
bJBmnKIrtkPDHDQXzge2oLqkqiu+ytHSl2cOXOLphT5kopL6zA0XhNjatwZydJ9l
yJdS6mw2kMDr8ibf5wqrKLA8YsG6BkNdd8I0cajr5ub1/CZ2kbFd2bdDqC5fAAwY
tmvrG6d6vrq247C4cKF1AXOwrYR88sqK0YIya/r34y9qjrsvBEO0tVydjSEppcwk
hcJiWnoovKJYSQh284+YYoOvxJ3h1X89FrxzdGdTp1cBaUFPX4IoC0OB9qN4h0j6
3DODCwoP6nYG+qkccVrsjGWuqstbr4zr3vFQVbaWKoxXBGkvee3BpTTZ0SOsoOHV
Gt/NsDI3lsJdCVFfs52FowdxYdb42JwbFtiLe7RiXkp8uJBaZDgLy9BDdPHzkG4r
SgwYhzWc9XQ4tUpEOQVGDiFLuQ2M+ZZs6zzCE67jJKUCkr8nm7tPkQHi4AuFt12t
rshX8qiKZimuiqDXDSUP8FVpfjGPmJ5I3W2dCsm194+Vb53+n/cJ1IXjVLIJdHRD
etyl/b+PGO52Zd5szuJIOzUdWKRqflwviPpawxt4joiuclYcLHgDKZKLf8JqBf+8
RZcPWmQW4tb1cA04bGYRCEoSN+xkD8q3H0dbkoffB5fhkYXU+uTbhMnF0TwiRmXV
9U3/TNewFw3JtWYeV/ghAIQ6OjS3f7brqDqhE5BteS+ZOP9SH2IH3l07+/AfBf0L
2cfchdryrL8/oSukt2baAS5fPr97trcifRoV87b0xEJiIrLXky0TuLWvtynW5UCl
JIWfpAQ5nGyRyWwwAU6EgceEyE1kteidRAMk5ZLusYCqkIgcn+oD89+Pwiir8iUN
7JNkGP8swxrz0J6Dz4VQPwII0LrpJppvAQd0an8oPrFWKK8hw2IU1pvluBiuqCNo
0vsEsvDZ1fo3ZW/FFFax+mPTiCKYuvj16RweAo/TaTQIXfEuww5FnodH0Ta5N/ky
Xaw66eyO8H1TWXEsmLw6xfh/9l45vVLzSa44oSSXmN47ZabPbWVOfH8fp4erFU5+
adgx+A2JvaN2UNai0L1hGItSgc55YPJ8lHvRQtp7Bak3QNorimYqvY1Nrs7FSSbt
AtHnrtMr/kCGcmGx0smbb3LMO+10c1jAu8XeAzIRRRQFK3JRNj0O0X2cud31CM+g
bSQdRi3VvFawPrbm4WO/C+DmexfpyPC3aBbg4aljxyt8VgBMHSB23kBtyxVOOVB0
boJXZGvionAF+IoRDDLwW6G963vHD1BRngC+bms9vSRkMO7SjeshrAZgeWmSODOo
WT/P6EfXto/5v8jXE1w5FEtc98H6EHmDUmMhZeZ/V24LrznUcrE9s8/OhPmZ+k3k
77+BHdFwlYLnYc7r77CCBsOEwpTclJ7EKF8dDqc317QNqM9Ija+Dk0dL4ViKs7Z2
Yr3Milg2nYvofAaudOrH0APl4lJ30H+uRC449IKNQ3QSIwUEyhUHJkr8VmzpiUgA
/7NOtvNnsEXdS4B7I/WL2583UKkzgaqRjvaUpVf9GRwj27CGhBRNkL8ZxgISdWbo
vtiQC5D4Aq74KYLWEbfaCrEa6v/J8VvvTEz0LMuCqxH4MyWJ9XDglEEmgXqqkNQA
AES3+RVteuq40n2gSHRQmLBXtj0REczNJk4xDOt7rtyW7Dypn4OK5ItQMRfFS8+2
sQBa+KM6q8cuKMbcfpC9TeH634y6M9wWGUpvQ5s0Oerbve8Fg7StNEKuWsJL55/j
Lv7TYYnrZas2+JlR5iEa5+01XAvu9YYfWX8qI8+6FWSGKP7Xlpn/S2dTEeuUgbSu
+X7mXgpaNJ5qREvDP9Kimk0kENv4LG/DXnNRKRzsXpejj1l3mLi605HNgKKF4mDs
j+W6eZaKATqg/lVvGeNqxiPdw0JGkc651Y5FwCrl8gdJgsQ9YbeE0XePB3sixVqe
VmHavFg/tJrNxJozpODSGrcvyA0PZED0dHypP2S66Rs4Lh2pUl1nEbYzS47za13Y
5rBGxqcGcBl1PNmGaOZ+4/+GIbqx5jk0WmOBiT2KvbeKxy65sijN+d6KSWoCuLtq
cMvlpNlcoS2srZBMCllzBpvu1q30vnq+IlYJzUI2wfKhdk8iwhDLI65UwurlOERD
HHrYVbtoc3pD+42cR2PLASVYVu/NZOlfwPDaNGirYJVJ548TkBK5cvJfOIm/Taui
P+7i1nBeLuOB/RQplN2bLeIN5l3IeNCbVCixk8qm1nC6EPV/jwNs04vXkv/W7n3U
v4qey8RWhj5yFiX4DUP5q/fyA52TRuaEEYtQpwjJIFb5I5cptl+54EIWtKkvA8qE
kWbzuUd0wPnp1+QQvSfPJ127GQP7accnM4p+FoUhTaikrSPKPGUkcwRqeKyvKHTe
QBIZKs+Yp3dH9/USRx8IGykjD4HgH7VjgFBKURIRDRr4JlhVrm2uLWI80ehqhE6A
EOkqcL4ddfOFLdh4UEITEVOEQZ/EICJiLK/uRC2aaj01N9SQPC6kNaC9CtiOUaUf
YyKHSNWvejFUCfa9BQyVBoECWAzMPa15wa8A79Z0WLmfQKFdHEp3+3G9py6oRm0N
B8RvB/hiDEVnjUFM5Nwo4gQWPRL1Aovo2ZMoBqpHs56Qr4MBZiFzAzPFLWSpWX4D
2ZCZkhzMiQOPpQpVFNvRUsDpUzVndVFF6ZGzp8b2ZEQo8kS5kZ7n3i1ZBE6vjmTT
SkZlYY5WxpuuXXUp66Ep96pypZajhLFoYr0DAHR0Xa3MK1v3mtYDngBgqrEMCJ97
axRUT/A423DExL5mtsNP5SUnGS9wA100xh4f5UPyMJSh2a+m3GAtFVa3XzzWu7+Z
zpPVjj+xSjmIew+qwvykr/C3EJMXhxJPO4ZDxr5+aYYQHGYUhBIryfsvwXWdBMWG
HLpxMudCOcG6ZQdHKSqKEAhHpNMwH2ttR93C2vcwKTl/hZqaIm46VpABTxIBGuPo
OExvjW/w4qZm2XKGoEkKxuWtLKnYQ160QQWjYdgQdPyOYmaHEq3I7O9MWdQY3mfv
ZQ+dBpGvx8aflNelfHZYBvyNG0+PHDFDuB2Xk+cjVo++3Cu3HB0F7XHc64tQkYMZ
8WAOXXV7wiwqjTikr7sEp/Yx8fxshmf9EBEQ2NUAkPmNAFhUe8AhLkNjvvepgdk1
G4Wq93GGhrDpZLirXTwX28SbaFb2iptzwb8lqg+dlR4b9bZoPV4PkqIlDU724L9B
mZQ+jwl+7o6DNkVd9D7F76xaikAlGT4Q3R/wxW4vRCHPLvevgtjw/5aLrlPfBgn2
37VQqqAgyatDqKJKaZ5fZ55lT2Zc5KtRID22d+tmfuOOv/uAWvm+uKA/KAZRtuhA
OXNdm+nhn+b5d+0+ywpGuAkNrLjvcP9hAEhkGz5ZlzPZUnav5D7zd2T+Q8jR2BX8
mQhq7Di367wkYburKKUFEtwLB1szekHekZtRMDFKHIeE0ScNuTOYrQPwdriQw32k
B9fIkJby3cnK7L547rSVHNBnHkf9jcjLRqC1Hy9J3CaARKZG5Nd2f7iPT/nI+mBm
MbX0twvZFjxbISVcRLjvCO4HeuOTi3HnLByWuVtTsZ7ZN4eMbZOPVmdSzUoKT0pM
+r8yHt3LLDKt2v/Cqz236Z47djE4zVxxTmI1NULSx4Wktt35O2CBJFS8r61aN7PB
yQpL/oonz8gGOP0EMHS9kKB+y2R0Cpln52Bwpbh1pgxgtSHRABGRyiCPEW9uJbd7
+JRspoMyald7SRgBSNigBc0Vjfzwuf2jCeOmZqxtz01JmNkNWLMn9Gww2qSkyJEW
F+MlsB/JDUiXo7rQhjqbE1FEmKDCCULU9vVBXBld1ZVb0rxQo3nkURZrJP7pGQ9E
rml6OktzwDEmV8gGKNVHPFEfk0EGkbj2Dv83gZl6Ax93K2mUIoeCDsJ0Z6X1zovC
4vryJV58X2cRoR7n9jDcCO8C3mZuiYtROfySAlxaK4rYYYDqMxEpiCzfd7LvD//8
0ldl42Jwt4/J2y0fj6Z+/vVphWgZNOtlu4uAZhCTL50EzJ4+GnasVQkclRk4sulk
W/bBffstqMLkurDAkHB0lLVzOaqvdoTky8PhjUq2fv8MouobxrZgS6+1t2N5u7oK
eAwwgnSa/O6DWRd+DWxg78wD7N0evtNzX4M/HTwfVU3LCENh1bEoLEAhASqDKgCy
ge6sSQ9SYqVj4NbhHA2KpIApwbOkg586Qww/2Qq/wOtDLxLSXBMAjRUVBEMxmYy1
Jem58yz9RNwil/ssOvR1q8O8XhxtyBepwYF3lYyZ7ZL7WuIsM86XdcYHUSqDwUpn
epgsH9nEQL91Gnfp5ufTSiOZjKrUWBStgqMTgEA8nOConHBIwrA98PnOD23JCUvD
6isBAwdItuB8HLbBVVdXz9gEJThaRYbcoYurIcUKpdj6fF4P74nCZO82YoEqUasv
r+Vj2iB8DYFKHHBhFgkYGS+JQP+tbxsnz8W2gxk8TrwOlKKEBMnLPK6xzKsKcuyv
5/1mbd5XDBNpRGVKNnV9xQorPp5tB/bMIaC5XWC8rALZMKSSI16IYMcKBRx6pdTt
RqUlBsoj3FsFJ++NFJiHxJyfpunFrOpPHW7VB1At5mkxc1TveJ6+NVGf/gwgFPb1
Z+hLBKfD5xt6XJaTd6KODluzwNgCEclFT3waHKTfb8MlEkG63u80ElgDN1TX2JGu
WgbjQKhRKszU60shORoDYjnL1+F/O/uIerMYRMED++NbUlmKmvqTmP2I4eoy00WI
hMRcxgXB8NebTrjYJfhlL2kf737xafXLHUoGMQ0POFZ8eIAoOAU2iqLQAodvuP6h
uPV6B+o1gGk1OWus+QDD0gRhVnB6ui2rTilDYde1gPt/TH7NNvmfwgg7PVkWJJ7u
yfgBnvmBr9QVNYEU7eamPobdbim4dJuC4CFGByIa4uS+GoLAFZSVXPfEJsImWps1
9CS1p0kBmtrzldeGrS2Mzx+xivCb/nV9Cic2T1JH68IiU6z4jtKeShDlzXZ2z7WX
ILO/Y8Oe/DRX724WYB/zAm6ja4r17Rkiqzsoxwg5T6AKhMY7LzuKlZwgl/0VbfTG
WFLz44EkTNk6nusoP8DLJis7yDRrh2ZMtBdcTKCZHPV2N1uaXVhDFwKbmx5OBwoJ
TWAfYEJ4BLRpR+cT5/vZ8M4dVCyRmHlLb3k0/cBrI6sLKgg7zgMPaa2HUiKlqL0x
la5HcL6hZ+VTet9yAXwI0oOGlw9jlQhtgODrBizJOcFlDNdMmQlnVR82oZStMKW2
LDXMRBjVnYljzWF8BfmERShFVAkdi5A+ykMhZGT6sG25O9H7e0+FXbCifdlgEp7h
EE4HIljdAy4qwYV6JxUwSasJG6G8UMiIS6ziK5LFj8xG6wepr0EjdhYGRFjGu6OH
Q692nU/yqFR+4mGeuq/AK32cYwP0nc6r7vXkAeJiItE2xn0g+ifombiDnyvZwb0j
ykVtzPAF5llKL/iDuNm5GJGYPCiOyQnJthZYO0E2qWuALw6ZfcY+tjKh+zPOphRx
vTJd/G7yQFEW423habBnoaF0M8hWkRkQvILEv+wY+4hICcvIPlRKmPEEScKERoSO
J66Swn/bJz37akyfI7F8TMjBZ1oZNSiywyDP8TunmKXGISuKx8azDGx+nC3zi+eK
lGU5AdwgtrDnp6gv5a6BWwuwCgmofTyQr9xYawzO6ag4s9ydQVDHsTJNt3E/8VTX
VSZEGznv4i+Lxz+ajUwvIpVR82iGz761q8cNz1nL5qPFTBHH6axi6AwjWs7OU7IJ
YpvrRW6xnS/Hp2eKIFPgTqNDblbro+V1f8CWw+R7kHHuBq9Y6qGUPtkGu7AlAm6f
XjrWFAmRd9NFb5L/XpLIsYDYe5uDLR7baa15+ObK0+CozhgLePUiRQKSiyG1DmRd
/UCsQMfc9BdeXHbW2NH5aYEzeeH4tzdei2GnQu7d1oyy5djTmk8o25THBRlAbLfZ
VZn+dns9kC42PQ4MqnfuH5wgDnLL8+VFVvUDsAhdyFBDqIgMDvtPxT/PwfdH/hnV
BXBLEHe5XtW5SdFSOSqvRpedV0Q3U3ih1R7YgS/k3GVfju+6vE8m1IXDO7AgddAk
26P8qIqynOpdl+nVTtijs9YFcjvWqBUBOPjfMJKZDPDYpPoldY36GM1v1wwqKUeG
ToxNGOGsIRXeJg89u09SFYyvWazW+hb+VZ4ybCJcooifqsec6+FbTu7yqARoN2du
I4YkJMQZvJaUPox4mhilmZhq7bACOanTPKR28FhdkobrQ8Z73WE91CBoGe+PaCX/
qix99n8oHriffxnd5BM0HZMgkBwQz8knBKOThsx7zqw/z2z1ldO9qq7sBVszqRIf
N+IwQT86+hSx6YEHJZawH8jC3zEvxmAL3g4B+6aZ05gZvMdhIgwnNgaEQBxUQsiJ
D8q/xUT3tSRvXHfIWYn+5vb6+qVB5ifzzelw4LCGip2QU4aZXRhQ8vD1q3f8vD4Q
u5gaS+4mUzu9hD0bG1vop/lAtV31r5o4QA3iQzrFTzIk0vuGRsomEAeI/oweeDje
/AqWgBt3X+sxEvOuR1f/BQ2mjBuIwpN7E8bTeSoTi1Lft2LN9f38r/QtOFfGsx3e
pbboT1eak/jUGu5PN4fiA9hmsjFbn6vUvYTzaAHu474tDyq/HOY5ScMJnShWTiOu
KeUbceS1thRiJTM/2gxzmZup5m23Ietq2UYxKkyt8FctkuRYQWdaX8O15r2uJ3Z+
rC4pFuGk3N/S9AU1NffJvgsH681p3EIe6aw0igV14FMQPe8FT/ibYA+mv8tXykup
sgVGCPzhFJGK7GdDoRThbOGllxEDNytpxPgFzvIT+9tmUxzcO91atv0l6/V+1g/1
It+Og2IOxn5clJB27IogPSTWoDjQOy9dLJIIHO5RpHTau6QwXvoutUglfa2c/bXC
djIlfNySYAz0u1u5qLWQuRhxh/Sb1Qk11pXXM+aqp8emvGae1KaaTyIoXweyfbER
60SH5qAHrATKSfw1Tgc8PsGxz56Cj+IPQ8BMnnLE/P6/WifnbCzzWmcmwWy5/VwE
NfA/4lyk/YhP56sssW2A4OnXnNHhq8PPVeUPZNdEHsnkRDvGPfpD32LxiinWPphS
mjh7lLxRkE6llqblQel5fQMSS/PtbHR0zfCQhLkfDRgcRrNVsJ9pNeyQf7JgiUet
8P0DQdM2DuBquaAJ/3wigItFWEDmh6I3oFdjfldhUc9UpOZrTTJ6kk2mYWJkcvqK
/4nEkOmVXdtKyIXFUA6NH6ea5H3TJkJ3Tb/Y38TmJ0oguuDU+TDnkxAinUwI5/Vb
5skiU2KidGbRwUhz1wm1eVm2r0uKLmM/p0Y5p5B4lnSvyodORzHb2SQVsjVUl8nu
b0RuZ/0OQPMJ2FQtTNdMOIMFeO8IIHu8jZhxLzwUrl/zNWS+TeWO+HOIBzy0qRXN
Zrf36vbYU3j1fz/ZQX2QdQLBEJd3VQvmCPWJODrYjDyo0aNkcKh6mLD2WZ3dxegH
xCX8B1E9dlB2U2fUbb3+5GVoaQqwG0FMtU7dcGcGfEsZlqPofeddfYPGwJWt+ov1
XwvKK7HTbw9fpSo7JYNIRCy969f6JyIHWX2jgy7hVnTDi1W+jqOTaH0/Hlhav7q1
hBdP1X+zmMpyUzf/vDJbVckFn83S3s1hOd/x98RNw9KrHszHkjN7ZPQ0BAOStY5C
kjWF4x5HgjANuuMpYt558sLHnRnYQ7SKwSvBwFA6LCMMY0Rxmgpcz5CZ5uymGTmU
xYSHo9Qrfl8igEG0LqlyLkH8x9UXtBz4btNN7DW4JM7bk95EBLSHiv2E0GUqemtx
WAEtXG1gVeimKEULI9y2ihVy7ReJz8DMAs/npDp2Vmv5xBgqiu1QwwOxNpb2FWSp
ba8pXwVVYQ0mK2iLjC4vdSgq0hjhYBh0uEdb3uas+toYn+pPkBaBszo5zh0zR3dk
d8qYzr2Aq8G0dhsOG308blwlA3Ius9x6q3evKG4G4w6ONS6SDn0cVvt/ZVhyt4um
yO+aMN1cNktI1HPYUd3ZtYUE80Y28AiSuM8K90Y8FPYqwJtQfimLkGLBRABa4wFJ
wlOuEHO43IpcB73jJMGZcTIdeDN3ddjEuB0Ez5HNaMrwCdCbAP7310UwEcwB2pWG
gHE7XHFQehojFdG+lkOHUNjOJNRLv1TAcXgIuDRuWnyhOo/UTJOEDdE5Z0dQvVk/
EjSpM4qaAFxAr0tTRyUC9mHu8uij0EbFYAZ9XqvJEDobyR7wSEuyppYkJ7TfmTZH
zjfY0oeEV5h/V4hF8EvYmKvkR+6E5HY31QbtZC2Io7ssI8ytHGlYllLrBjFmbNlg
1PjHBjAO68Jqu2w9EuQ3XxpKTpqEoewU59uHM/Xhai+gXfIFOHDxGW3tJ898fP4i
/6zE7lBZurK1aRUR5CAvNop8EX1nkUO8wLASk1OrXljduP2Os8+iMsY0/Iu0Wotj
X/FYwB1RGe7bfNafD0Cgv7YYrT6n7fL7H2iF2d3S6fdx8pKBAaGnOxPmRIELp0cm
hG2bK1b2JiVpJ3wxcP+/uZbd3dtH8l6gZSeSkCqTqLnEEXl02b+LjXX7IKZoBt7+
638t8UkvNZV2zuMT3BP0oudOJccHnDHDXDISU50U6fsxkzkrdfAfPTffXlklufzs
NH1xfj0Qh2q/z6RhtsrV2VG3giLZfnctPdpdR41RN4uRXNZOUkFEqmVDJDJ7D/YB
oj3blxLccRvI5VlUifuUcxso3t1WhJ7kGtq94QpgeWmZxx2MXa/UV9KlsUsi0tVU
om+F4hK14A8BkqOBc+q9y6bI8LvTPmNuOySOgX39VNrvUBSO/Ct3VAbrhFgPSpzk
B9WSKgJbPVauBfnBl6Ib3GYlG8nLxuCJBvHSK1a7aNfnlugbcN/btglnRsBz6EXN
lQ40zVRngl7jTJ/3mvqfKHHctya12KdFJWCY4cCx0hY7uHhxLd0fY9UvuF1C9aMM
ELl0w0fRsvUZp9aYNGY4Yfrw8XImCZb8QoUmEHJro43DRc3FbzdvlRN784PwFjS8
nU9UwTdNQHm6gCaGkIA2DwmjtdqVIBnNlNAryWjTQoiBoSu+kF2kcQwee3Um1Y86
PQsZ7m5iSVYsIRscQeVgnOmdBGR/gECaFN4ttus2nJCNtmGEWPkv8zUBtYN3cpjo
FoA9cnnwjzCdPkV49ar1cRjJsZIhJMrrubBEpyddtGCH7YwhhUdhvN4LUIWTIj9d
AsOGNJEHeveDfxmUsildhcKiCfSnrn2As92T3lMo0uA0B2JaNWadvTbmD0LGIuUp
6yBMfjaI7aXjTVBAMKWpGogAVwKXzTP6kf1hB3mhMMgyiweh/Qe70P9sO+cM75fQ
LtEuAy1nbz/J2p8vgbRL9gdqRkPGtLiQBJw6KXyWhpfzH7oOPKOsZ7uegcGCN0C6
ghtY8FUrT/CzubuhgEXcXgNOzwHPMSKX9VyVWxnMGOfASI7AOZJ69IdEOCuimPUD
ubSkmDpK98ptGJhiJXvixY4gg8RIQPggwWV8GoIDXHundlXpvxp7zebHs0UK8tIC
VtQ7icHIhY4QYIVdG8lStevvajfd7Gowg7Rqj2EZg4IVviAD+Qo/32fx4CwkRxYm
zGdOBTqI/NI5MueE63Kvd1/LZuiv/xpBlDQxIILhiLC0cp18eW0tdInGLEyvw14T
+laqlybAJ3WjIbvePmfXHz6MWIF6kMreYQgXgcJug/5IQgS34ThCyGxvzcnlMgec
nnDo8LlOTmjFc9SSBZxnglo8f0m8HWLK8ndhKyXa2not9bQ1JpBBI2YL4ZuXpCky
hTVI9jnAmkp6/Ph0ooi8tytACUYc3OdyMDxkHEvLAEY7G5GHcMsFLKnAOhYVAqL+
d8qNOkl6HSi2YsPu1As5IHXuhRIbMkbT9UOroyOF6RWlitRt3vspJB3xyTbMPPqe
VlaP9G+h+UoFReTiPjM0WWXvxLwxcTfnzHlC8DAM+Fnw3S778V43RddxJ+lf4bKs
my2lRrJDyJs0w71xBo9CqlRWZiPVM6VRarCh2IpRizUPynPKDKbgh28BSWVn1yGI
Y0vRUaO0SMm2af3tkzTJyJyaosE9td4+w8Qq+oC4TE61eEGKuSot8PIZg0u+d1l1
n575YBk3LUTWGxHia+uSMMk1XMwIwE4lxyyjhvirM8MUHLqGgTjSob/2k/OsZe54
qzZfTGtpZeTexXZrbW4VJ9xRS4FnA4ipQWjzFkDFyzn0svq7ZWiGQvrJOLS0ASjW
dDsKQq85/r11sGk6Xu1EgYwCpvampqadzkgXYK9W5DfPMgtKoYuolqK2gM6FxPXG
bODqb218P9fCe4ZQVAOVg/0LSOjEywsVp07Ey6MK8crnl3dqjEHMeYkxgUYdKYfk
PUcXmtVIAr1qlDhOtEjDb92OZz7Kgf4OJneZ8usSyDHKdytnzIfvt6hdUpQbIKuv
pkOKE+fsPHiHvC8gsiCAuKeDUSxc5UdQCDsCcpmreXo9oD7E9nPHwsToc9bJfBAQ
CHEZSlemK1rQ0jM+Giau6aGKdSt77Ng1Dv5v8mqodBOKExbBkMOkEKLfD6l92FdO
wPhbQdiPceJtPh77KJiLtlj5OXXKk4MLOEhkl6TSLT+ES8bRq0NG7/7cR7gPZ1WA
ShBKcql+KxwcO0CgjfJxIDkt3ygiEUMfpvNIpwWdcWiirkL7q2LhkTGYT5fL4olr
JiLJ8oq/0neEa3FPN8HMrZ/E07sZyGbsKdnEipklNzAv4BRkkX9Y48PZc/K0RjjP
0mzge452t5C7RIoNXPzkhwapseK8WZL5AKclFld0a3taOUSANQ7ESepja1ognTFw
qBwm68YB0ls0+GwaYAewxgjhJ6akd4UX8YNvO4JLFaXDRg2x9KTwH+nnfijx6Dwj
O+Wyjh+A8tFJsogtgUqO3JqNLnltwFyykmfqa7L6Z5mfh7RE2GIp5oZj+5A+Qh1P
LhijpjF478iJjnnUI6TGukiyJgtWmpRhYgfVdedWAC+FezPrO9qDTmqO3PxrVU8c
kHiPUbQhct2q2z0vy2s7pctDZf6LYRptuGWJX+kITp0WsCOJ2Qv+BQmYz0iELDkj
xtfUfaMns1nyJVjv4XRiudyT1JCHjtv6gs4zq7zKYjbX3Fblpbg8LXdoOXiyil6x
ivaFH5EHDUWIbZwxvtP1QV/qokz2i9Wa85VCwIFrWlVdnane17YCqxoZb8o0jIyJ
9Y6jIl6OYAEf8rCGO+AaLGpmD6LisxvcQWHUito8uRDQsa4HSYImTcLIYj3ywOJS
rSfmrloTAs7winDO+PMkVu8KI+FnaYmWhtM7LxA0f9vR9lv4xorNpMtHvzkSzeQg
j0g1zJvtYm5PFPi+F9+h1ljp66++GiiqMd1uoVUK/R88peeCRCR0STrSkdoUNawx
hXvqgK/18BEPztKB4XAakKOsXtsSotwn4iW1PiXmm9ljyBILf2Svb3hsr7xSYK0X
kbgb3cuiTnVyupI0yra+KDO3hKdQrrvod3+IbmKjRab6yXSnNxNkQBKOEPAIC/ND
ZqRbl9jm2LFJqjz8InDcDBf3iirH28iyDC573WfRINLS3jgWmtT3Lp6rMJk8G2nL
xK6b6MiqS2eUMR0vR22fqpEdehBPcGRfKqEOAnWXzibuhaUR+f7f+P8z353t+jag
c77uKMYHqWQWp43x6CVoqAWolfKjiUCi1J4Cob47+tS/nRli+JLNe1cBVRx/r824
JIgQmz4b/378XAYtsWqQCK4NYnks7i5QPYIOvZ70R4WFeGnR8mztNBF17MnefYUM
Pyw7xEAHirkv2HLquXkrGvEzdAtDQOQUTZdLWarGJi8WDcP1SSky8+le7TcIbgQ3
d9OwTLeg9UNT3fgPc6+vsySaSGGdSjOII4cjJrnAxM4pP2ifbu/NpgdNIJghLIgM
LmrG1SyGSITc1HQw87ygdrZFpJ217eCHbwPE2uwe0q6VPQSGCwN+uNKIqxuzpp+7
v3D7Ivjrwmmi4R1JQNrWY76IfkQEy5WpGLnHL94+sLfo7KDb4eeyFD3+uznbGF+6
4Es9kdpA04mAZ/5Wv9rVyy1O5uJc9Kj986Pp09wc2mRFj2lpSNogBJznyLYYe8p3
p/WDsLNnAOfwNQ8HieM/RL07oEKNqHEYZrzjI4Q15+6S4tNb4UBv5wqNaMm10rb5
O29h2drN6h/cRm2X3Rc1EKkNn4BJwsaaHG4bERs1Fenhi0Rkt1aU56g1HWYlOYi0
jbJ3pzWVIEBFseR1DYz3VNJXS26DAVdgZ8JRQg+syOYmSNIQf4PtFJfGDvRzyqWE
olXGEekL8+kN/9YKUV3/V9KrkbW8KdRkdZfu6+STTseAuy3vCnGaBa5wDWXYazCO
5K3qWz8SM7TT6pyy9BZo14O+fmc8dtiKgYqF9r1OanuBaWOTdSRD6QPmSabF9w5u
SlrZ9dOFwZy3ZYcjjrYVvsXN9rV+XmdWbKiFzukIyoWMJfB1IUuWngB2wJfUZPPC
9QRG2vdTRYTF7FXMSFO6lNTglnyPJRPAZ56nuX0qDgMke8uqP7J0r4i/AOWRT4zI
Q4iri6n1NbPeNfVsmJ8d1X5zphUw3445H6DNyxgYFc3Tt/IcrVjneZwj6CQ2/i8K
8pRxbiflP7pjApZKdj5RFf+c3fxCt8iTk55L3tK7qSHDc2fTuzaLjtRPY+UpH9VZ
ErL/ruxZyYfBlJBiZgGO4jBf5/J5ouWXqSvoa2gCA0pXCTXkF9qorXqJk8ijcKL7
LBHDts/H/X3uuD8dZz5jXy9kwYwfmeT85LgYcgcIz+esPba7pPMC4fs7OG00hD66
R1dwZrERu+PO7y+TFkPwDLcxkayi4P+o4XITf6fAjfZKELoGHPJlbcqB1QVHNzqQ
OL10EPZUZfjD/nBkueY1Kjh5LD/bhFxZT2VPSBzC+4S/nP6Wau066owr9UkJzmCh
zTJeAiOSGv05hJQXtHIjsUfodkbHMW23YpoCZp/REZu1046wQeUnP/dUSzBmyhxQ
Z4BE1Wa+iMiJV4hFh3qsvNWm2GK3DWDS44I1qLkhXIL2asLLJBSriqWyrRYVp+pI
mPgSHvlNp8WMswULgrWL9vT48LHr5G1Gse6UCJfpGd2qdIUeWqKpEmCGa9TQfFhz
Pir5K2LypBg6CeXClnj6g4ea901nwD0CXLBFUO8ICznSKO/DIR7oKmgBzGXtSqkf
5kCcAsmURwwWoLenXvhyDYUEjUk5GeTFSYEj1JsqSv+3GDHYEsWn/SV5qV/8KSUe
ncxmSOSaNEzkx0RDZ+YsXr0OmqGy0FHLP8D4twPM6bnqYmaOw4XSMRHq3etjjQH7
EhwC9t4CLtBg3Zi3C78g9RfRp4eJfEgLaferPaoiFkRCM+HDZ5tq0+rwIitdxwUR
46GGryQb7Wkq4dVGbPch2atIoRZGsR38WjrPuf+Z9IKDKnu19biXgNRD2I+sdf+o
0TV+gF34IsWFlIfVR8qrFyz7053wkV+fSMPLmHYmTzo+siAYynjtJdPVFHKDIGL5
a5g+L2wiUzNvotYHm2VOHbeLb4yApDoxhGxM/2q3kujpNIg+LG4EM/XMIIweK7KC
hFLJQEuGeZXVmRY7mgiEtGnjAQlaZIUvCLP2nzqRALoCVcP5JKQnohmZBsTL12kF
RAq60TuQUmsaR696tXWw2HBJLf94fOFqYE5YcJMl/Ernqn/zxpkKEr1fxI/YAeEi
2tQK9qTRZy9ZTdXMxFQXsR6hkObh2SxJsOigaZUOc/WMWZh9huedJEH0L16Q2c+e
H40ggNZWtTWQqLF0NPDcNTmkBgwQtfD8JsdTrss3PxBURb+0Q3DrKj0XOX9Gs7LA
q9V11ot3fkredb65qEnwu8rzDlNLbMmwTegA52Ayx/npjclynQEiXsdpt/BuwRYo
2H/WVCC/yugXctqVTgnzxReN8KjUWW7KZPEqZB9HJjxkthFBes4F0riD138zaVj6
loEm02AuUpDTiVSlZQQvCzXsR7WM+b/bD1AgzRFh5UQjhnTsgKFJA24vg5IrKPgE
4xgKxVcgYjngvluDS/F2NBYI/RiV8TAsqJMtUIzHQR3DU0L5Ch0otJlO+tj4Ev8Z
ZA0/kYBUvJRphBiJ9wFudP8CmDdTh2PEIs9/+mTDo8KOxje+DlhWeqXU90NzTAvh
rofbcQZn01rrS0VWmSg2UQDXba2BvfZ1fs6X8EzbRKCdOHBr6oT/hCk5/1AuCsGk
bCSwuYW6OiiMENnWpb3ATNkGoaHEEL1bCwNAiydYanQyG2aKzNzG/nkOn/KqoT3S
I0xVlitqfS99/y2DgSartQ2Men+58c0670sMGAZKI/dSfazI7I7/rkshTcaGgPgC
zEzsQ/dcOyC1XLvFK5scka5FulzDm/DIOneB1Fpgrejh0z4Y1Yx8+uObVAALbF0F
pdYk+Li5QvPcSzpgJxXq4F8ZoW4W/RfkZA1kisruYopt1MeT+jkWdT3yTcGNIHY8
AbMWwGMGMfxLSMof5L4sANAAFKlGXfJz+ElUmikzmKPymljL5zti6OvmerQnG+uE
mBB+eQ77C8Uf2+7PnQ+u5Pje5kk4GwloJgILSy3LkFvSLQK68xNANTKxtRBNZ8Bi
f3aekewO+1lNYpqL/Um3xsdYJDMyF+tkllyvRmGv5r0cArDvKGp5gS9zJityncGp
NrNwEY6KP2d9CUprtuFKt2+ymev70b8Vo3dIR7rKTQH0mS35J4kRTPSfbMzu92ZR
So4q6eDUESXOm1Z2ulZw4Uv0+E8E2Gl9DMTHSvWpmm+yLh9sApBxgBl/SyFZiyQb
jzYdhmvcvLT/4u+Lj4ByigpIjOSI9JKN6oocKBMaDN5+uG7WqSr3T+KHGIXDa9ye
nBfNnhC1ujYdRX5jqvZoz0mKi3EZll0sne+yalgYz3s4OCIj2zK39Jj8jZPPgDBk
OywiUfVRZ1GRJOOSu4SVwhEkb6PFb56yRtkRCcU/F6wko927US+TGRHX5nuKyT8H
yVm4KSTmJUaXsAUqritAFQPAB9WiWQW1pPwVj1OAI0DbNVbWMZkLPbfhcLAagRzZ
qMRgFbNPbUfs/ozSvmuuGKsepIKmRBcnRXsC/677KJejSRejHyqW3riMsWWr+NTL
azXMJyM1w/QRzR3T3cuSaAurQGqlanWGftfmOX20NlUdZ7p0PZiy+WJrXb7NnCDw
LzcSxwfacdZ332q6duUNH2/wxa0eCvu1vPx6nl/4dMdcg/nZQSkICCjbFzwmqWlL
fv2qDjzQOJ9tijBhutjR3hGzyM23HDy62eJ+BQ4e20rJ4LGCKRK6Wib2I7WMf/7a
CuLZwcZ1vaJQ7etMtKmn6WhggYRp03ddC/bAe4qMclTNONxBnvnOrtsqGss7SpOw
zcwiNO4rGhwhfn7F1dBRXTj6YhuVj1MrTk8nEKGyWeI9eiCSOIPE4EYZIM/1Jbm+
dy0aTjVXUpwxXyB/7szo3Qudvq2zRbrw89WNL6leb3aPlxx+U17xnfeKwS315Bkz
Ir3vn2vmOkDrQLvU5fyWA9f/jKx3664CXuXIf7PfOHSVMZ0MVpZ7V4VcLEu+T5Rq
uEmXp5o3IYRFET1KMCfP4p52ughfkqzv/MMdmWIIiO1xAA0qEvbO2S8YQCYtoSQB
ItsHuqv4h6rCGk+TXWkcbozNbaJ/wgKicUhYNWbNeI6sByuy6XJ+HdTdydkX2K5I
48/WcmdyhdLSw9/9PrxpUQfH0Y3Td6vHLalBc6UQ+eFC9vw+d5lcNzGtLZ/nVK5H
KOFbGrWZ8H3AgVphZWLQi+106V6EZ8DNKtI7HrqTPRi5J/esVVTPe1oTeFeDiedy
73ZMxr58eTAypJjl2Q+fFw/tgd2Yoaw7/alPsjOZOvHbwWUPIZ761RJilQDA4oFI
THOptpn9YKdij1dlltyioHt+nk2erAD2EXoOYcAfDctKVIu59tTg942Ws9CgyuDP
cFsT/VvfiujyGy8STmUsr4oILdxelXvYsTnME7ayigdi6Sjkmk4gkRpyVt3zYJ+l
yZo84tGEKg8+P7YJk4OcL4kzLIdeMiT//IVi1FlS7TmqsmpFiAlUbhh1cUaLd9kR
yn8PgTaU0wX62qWGwCCPt8mbJVkfPE7ZZBG29DeNtHTAgDmbshOPA2mNCHfGbEdP
qSobXlW7x5cc/+E6AxS3+2O8y6PYRu+xZlTfMlD8jLDp963UDIFsr533R13U9dKL
idRC4vNjBHvl/aLeCW2hMVdphFEJoX/UYjhRVEONw9vGgWjzHPbqWY/IwQnmvDkZ
q26X8NDBFcz9LiOa04mG8dIMntOphCIk3MjZ3BGtmF3JXX0vdSpsCXhkklCXB/HI
3NF0pSr5wrpKXt3IpiHmZi1k6TnJKZ6bDBzmY4lIRw7rBI2vi0zUMLjcVJ0U4ZSQ
w8DpQRftOQiLG/3TSabPlcA2tn331IMEdl1IKqsAcbA7/sd5cog74KV9K2XcUHuW
UrOVwUTsuTTkG5pgSqM3DVia2ZAoq3c1fxeYTzUDSEQTj424RgTqHN56jknLCEjX
7+AjcdhdoWAtjeMKrrjRrisVIE6FHMSzQsJf5NhjA/Lfq9LNB0iYnMGlmQnNjNCa
UL3P6oAabLwNkAUT5znc4wwBtt6opN5bzOUqMzrQ5aSNpnq4zF5gKLmIrKA1/Ddp
mr0Rt/gLYLTWm5GeJhuq/E5KWDpT0xZQJGE1YzWjLxOrnEROO7ObV8+GwcEMH1vz
z4rzHenHcocigTUAWTkOQ0iJeEVf0IGai4hwNOKMrkytaWo4HmmCl9tpUBMWDzqK
entWOe5NQwTUieZUbd3jYw9gXF3BuUNPfDChyFiJNzUbV/XMvBi+We9XoJBpmpSr
fxow32FqpX5Oap0VcXXxk1eFkoFiGAWJp9eriICQJ5JREYJZv3y+gYEX1QTk1ocr
89BXRReotLRov1AXJz408CPVeXz/GLMVQ2Oj9HdwuvxU+8qeH8U6DoLBrhliP4y6
PKF+gqZIe9y0/4WhXJ8fNDxiRVjZOi2WB+rRtOcOzDzO+tzzc4hnv1K4nLnHTS0i
XWABI+e3BmoMafqOLfVA2x3Txs2bA9bggDFgdED6/FVFSqsfhXizFIbjJJoUim1j
FUegu5p1ZkF//owWg5rZR6zdSBeKTdJow/yjdNsWicBX1SKbFk1FVuAgkEJxsxr1
gdOJpQr1TBfypDv4f9tRd8+q1I5BDMHkrRMcyWGMR7qnbQT0PzBF0gRnXKMszh4K
avGxkObHjw2JyXTaWQRGx0wn9gYzudEBKwH+Dvy92YLuquszUOE242n5qnG5zHDb
b4G7hQKRrDZ/pqKJrm64wcWtIvbfHFijtFZFT3ejn9TpR9FP9h8I4tkDsoH6DVIj
OBF8uxAQF0suWgq1ZublnEQvrpkS8Y2zjePKJqfKPnJDBo8Xt/P6LKHiNezalnmv
k/Jyb/eWblabiDMQFht2xf9UpntM94HwGzL1sG0Y1ld3Y7WkbytVwq6LL2iSrc9b
tgtSbSSxEG9jncY6W/QthlgZPgk6IyAeLU/t/YSQYVGFbB9Hi0DH06wNXExQtXF1
alejxOg34BR2WHgcJjbWN1LmL1uw8iJ/zKD8y38imeUVOp9fmv59kS0yhW27GGVv
f1xtfb79Q9/4H6KRrPFqnJizpUwkE0O6k61PyrLq1i2O1lkOPSkKepeDNVd1eU2K
J5YZn2W+h9A1jj4IhawwSgc+WneWLouMvRPUWemuEjnKyYBvUOEWFkupW8UTduLR
HuM8dN5NFpvE0Tb+fbl2PZqIUZ6upRRdwUOq5h2ky7mwiGDTs7Ur8TaC1z9Cy8pa
nIiEmp8I2l/bpd6vP60he1QtSFTtU1bdeRCspjzi89u6QPwmU2WBzsDw2qq82veb
qlf0pVimUNCxok9dvxoLPYLQDi8aniwhAVBZ02YwZcegtsS6VsrIbO2BXpnQWHzc
eRrZTi9y0EOcTjXgJPWgUPA2E1+lvVejUIFWOCLVdBW3AqzkqEDKWtxFDgDfhQak
xH2dO+Jt+I95wVG4V/9HeUkwvCDjuvce4xy2htoheLBedSWp22TQNGlofuXcz0aH
81LEj6EjfAwdXnbGTg8iJbD+YWnRq6YTaQhqeEE9ZYs99+7z4YF12l6ngklV7VLh
QDcrUcSuNpNnXI0VRSQudQqMGPT9grVdeC+9etpUB22pRueugkgpiMXkoaMxTXND
TPWXcuAlXvn85J3Xp8At8cJdDLCkX6yuTmPPE7wGLOkfR0WAZ/ObOac2kmA75YZi
AYng5dW9aUFiPQUyIAYbCHU9A2NdvXvfXoCzCmqpf+CA5lGnX3rHwLJcPyvs+1Qr
luJEpUsror11QEk57CeyHD4ZBNJOgWf2+lvod+hfR60Bhe3wWAOYOXNSsv0t60k0
CPMbXVN6OfY5RyIm1JTr7pnR1Eqnh3IuRahZvgKzw0YkI4WXft4+IfH6Br6eRn63
q6NYoAV02e8wMZejkJ2Uj8DQ7JYZy1PZWxB3fZD1FlivJWdGCpKacwS4e6/nm2Rh
bOOpnPdr0LlcqK/9J6lYA1JR0u7QjdquWdHJNPTXhtz63804b738vwU6K6djWHF5
43Y0dT7j10/ubH8EWTkBmpiXX3zIEjOluevTt29ZxpFOlemxMg+gRGOz2Vc07OJm
0xWvyj3KZ9VzFybYqxTLKEmttoLu+jyxrVX7lQ06qJlatorqC/n97fM6gYWvbDe9
znFn+S2WK0LEYC45u5VOa2Wt3/SGF7AY75ajRFfVa5AS1H3Fk2UxGW8oXXT9Emh4
L/UHy9fAhfVv+cTlMotfu4jYXSOdWOSNFcuxbwlZXPXfhwAO5yxmDoQDLr6im6U4
qYVlShcvEtKJY8EJD5Yv52UcBHXVFEBkHvEuLU6YLUaeGmu7PCI2ZmhhwV64gDLV
FCQ/AG2x5a6+JDozESc48RePdfj9pUtjsD+PrY+vTH+l5QtZVnsFdGVA8GJ3dR6G
XNy0EaNU1hQaB3niWncJFvjGR10DCXOE32PpTguI0331c6/rlLoaBjzf1ypjOV4X
SfXHV9kKsqnoYE1DN4tVkLnvlUIFQmHWeNMxbWRftr/aKKd0i6pjUtN65jyebWfw
DReiN0HgaJqx2sjaVPHcTOGzmyu+OFYpK2sWC1W0KwrQpKU5D3+Is4if5rJi0cHO
3P9Aqm8M32inaSTDHpdGjCasTF0qy5POGrKQvYPVOEtJz+T5EbmWy78/wxDMH8Gt
7cup7DnDAqMX76y3tzyD/hM9eRh/ZMbpjWkWSM4irVFbXEB/Odvw+0zVAyRpZobz
T77xSxMZRVRRvd/m+rdxN9LTSQq1zn/5T539WUXJU0WbJ/luXNVWVMavbJlWDkhP
6jZew5LDrQbAGXwOYagBkGr/hRqK9GgiIyG6vpneac3QLeBuwG95Rw66tGHI61Yo
8VjOigMy4gDFZGmQpXkoRo0BRC1HCs/m4iqBarqbdbqvpfSiNNRydF0mE+EeQiYg
4r5ByXMfcko20/MZauTDp3aucHrn7sJzoM3xleilcF8ayiednK9b0EqS3SRzIbTw
qoehOwgr2LI2oaD5fYdEsUpanj3Y2KhlfGIkNUae5EsXYe9jPT9fBH4cMfLO+3k1
uTRFfQBl2D2v7xdtE1UEUFlmvSvm2KAvt0ehQ/FtjQVVp3z5MYsigA1lh9V6EZ/0
eHXvpLPUGuDYgbfX0uatvPJcaZ0HWSP+RT4FXwqZvfmtQnxPjiuThsm5qha0Qb3r
iYAPKDU7sxZ8ZAkfJ8Dfw2IVAGk2/he+c69Aho2czcdtymwW+4VEjxtLUt9n72Jv
xGtd/uUdhbxlnRZlD8+7X74w9opHG9MO46/BgPzUNhI3gqPxJujXO6355LG+P3Js
Qs3Ay9tveHAVkivpulXSBAD9MQuGZvbDBA8gQ8U3AhcQivwlqRdIb32LM+EWG5gE
dy7ysh9DcpeJPj91kCgDLiJ4jaGFdbZ4FqYL5bP21mEjEXeA4Z3TwgkE3jSdpA+Z
JtgqMf6GqIU9ze7AEJaCKAfCbHldqpWFbnJFAQ1qzt8cxbHaBZgpApbUvXkelLU0
oOZkNDndKO6hYVQEAtyZOiwttSFak9Ku3ntf4GKixy8y3gqivrMOPD+lqT2M4H4h
r7wv5MWd7UTIE45P0AA3VqpXXkIT5UlPB3QTrlSW7REDI3KItKAyOVjTdP1xhalO
Ef42uljAcle3F9okio7JYdnWlQXKbjMz/O9MgoNs/mIi+wfBdn4dMXUmVxb1f4CD
9Bhh77f8iAoBD61b6Co6tixwHHWIHn7FV7CnFa+VvsoXV14T29REgtVwFvNLtSBX
aiqJnxbxLC7EitIvY8X6IiS0Cht5b4ag9ZN1Whw1uoXlYQtzkLslDkKP1p5yrsc7
e8tndEnwgv87GGvFCc4jPblml1A8/iHPh4xTK8W35Wq76oqslTtC7dwh8kXXeFTR
vdGJ+ZC7D0RyV2RWH2IUYIMJEsjDPgti0RZE/3ir/sF5RAtTRr87TGnKskL/1WWF
RXlZ7Xo7FXMlo4YsrKQ++OkyLUp8M9S0N5XIgCnvk2CgRHMBVr72MDUCjBI4jned
63z44aSdwaUIqvNxxMrAi6+fFuvgjijO94eiSuSyQ2T0Vo7L9u9bjI5lSwC2nZAc
A8fmxjh1K0B5bgxxDlqrjRBKgXHkNmsdjnw3Ithu6Q/0/ENZ8Ui99dvP/C6wbxG6
kgTW5ZgE/zT/RSx3CQqLNQCIPM9p7VS9aFgLaxvOyrc0J8NE898jr3BOGa+vs4L6
qXU/uSahC1/SLUZyp60WWCGGu/MKo2P9CG6/+YKXxj4Q/BtEk2rK/cVkgy/iVu8F
YVnoLvjGBEisBcGC2HP3i44BuhZuoz3XnArFZrp4kcA5So5QsVlEyHl9xp4zd3fJ
npu3zvPVmqX6A+3w8T1SvLANUmu9EPv7Mbqjj9C3KFpiK6x8kChaVYQ/u/F5O6Gk
UwX7yHlB/gPfIdZL0rbos+WtCDjzg/7v08geDAKWG+aZ4v8Rp5WL5EkEGte1fOCm
M/xIABa28N0Dr++8F4VEu5oGD//hALGotcpwIYzrg7OvhrshKtlzkn5JwlgRgF92
G08pU6GvzHLhrTnvBBrb00PdzBKxdok53FPv8o9vCK5U+SnpKYTKtEyPIjxCxenu
mZuTxqqjRNpPmV1arqry0RFNp1/yTwelWo5l3MvEdfD8fvVrobppGplhUMJPbpAl
du3v2neE6wWHl035SPyUCFm3R7HTowfJ814RFESiFlQMPG8rGO7zMGoTdwjRwSii
zja3GlGnvnpgjC9RyTnlLPwDQrS2d0fSkIe+4B9VPDa/0IG0nHcraRaaQEt2Nhyr
A7H1U3dcNeHI5lizYSZ2NMyt44BBnEZvf8xV21Z5bmYcJ2i3qBNn8EbfP67HDrNO
TOZCGePYGSHGjpYkmsfToZEpP2r3dfmiZboofzucHY7k9raUAQ76aj7S2qYc9ZEi
zM/DdcpYIv37Oaz16KFpuaz/TLt+YuSmEb8L8BZxFcKIfWMH2P7Ga4fJWZNRCAiq
VF5kG2C4b01RLhJzt0lSvDXF4CE6anBMwnNfPENj3no7LklJahsd1/aTKlLaha6x
KwtMYL5Z4QuuWhyHfxYp3MadlEHZCnvdNPxt4MXgYhg/OnQ1dy1yygb9x55kGypi
bIsfBrF5gAfwtM81Bcga0acIX2ldMWioEXmYmib9nMCTUMyjob4HdnE3QQFVlepZ
BNd4c4UmTNk+9sZVId9l6MddJcp+FViNtgL9IfvtyA15YUJ1vTBRtomuRIMvXFPR
mNFD+32RjW7qK3k9e3KNLuaEB0Mi1YB6Nhbtmizh1ax248RSWgtdxifsXTJSkuc7
nhMW4Y+3bdy8CzOYlrCSzeJZPQ8ccVSLcH1Ixxmo7swp9iAsPZhVhabUtpaAgT51
SpIEfY2pNKFf77uwcWNZk5GLjnL6jNcW8rs5uiTRpiJ8YI3gePZa5RG1VLcaHzag
IcW/jVcHeM7htUocnCW5oLBK3HNAj2q5+hvxxF1F1rvtY8bVAboTvKRZ9gT5SPfe
oKl18NHnqjp25X4/UYWlQn/xywmRptZM2ZRegWwAgxi5A+gKcHX6GO6EzPFERflY
fT/7FPH7KprRXhvPsstrZmSmo52pShdavxYo+yY4ZSybcU5lNp5FwzL9P7MvGDMS
8myFYHLPWmJyLAYWKERpBfTeBaC7fwXj4qfLthJuSGE4Aq701u1CdKRtn7d90HAp
CocuOFm62pQBKau+l/Hcq51Z2YT0xrsk/cGDPSIMWAE2sLtgO6Ovf3eRHTuIfHvv
9KGCS+kp9ZrR/DzDz+99MnkU8UVyce+3iXZAvs8m+fSlYxrOapeL4nP4TbVbZdwg
HkYpJB/Qnnrprpvugxhscbg8H1JG0e4Zv1WUNcESnF4YkT3jX58LbvvCP72IL46E
90XUKmIlgu3wu/hSSr8HkZVLZuMWTFRAgepsqHrGNU3/SF8mO4h9X9kVvdUZq+RK
poVfFH7pYqOcQabUgbpZMm3ecXXaWA/uk3vvvovt6vx81ixe8Bzg5wQhTleNnZ6c
j3mmdVtUbP0BdlxY0Ehdp3SMAwQKnr132bn2NK3RlM9sHy7jaEIb7WhSaU8ziRnT
ekxFCeKk+Ks3safv9EvjlK38i+OJgbIGuz+3LaliomZ+4PD6CqORL2rgjamZ6p/q
jfmyXWs7qAdSwdAqwbteu9lizNthT2y9/027aAyXLnZLDZJOUyPVhYe2ELkd9D4a
ywoPl3pc4c2pgGr5YgHA17wvyKbWklwe9opEol9RP160J43y2QfoV6ZQzWrL0B38
MGXl8+CGhgPqi9xbmKL5MgyCfVPpJyoc03yuBdgjV94QmbWxAOZvt/bVagm7bfUI
OIylH5zWUljyBYydytpZRC8rnqr78CT6YeMzbAdmqbYzYnjQ1jDB5+w87qbYzVap
xaH61owc8DdtjsgXlLj0JydoqUKMGTLcTn7L5yoxIk7HkviCnGBgSpyWybgmjqE8
QWh2w8KBjrzOYf/Dp/yRwxvnEODF1SEdQSxTLg2aFZcfCbOEJbbQ5dKXelitMR6U
qkP2gDqv55kYVTIosW27LllVByRstdVAijT4LUB/xWc+5a6mcNs0KcnZdCGNsGT3
Kkb7ZoMsN0yPmOVd04OcvuOOk8qCqIwPXqYTpx8MiLMlfd2ozXc2sBOL3I3O9ocQ
ChRJM04IUVfNDd08OCM6DHmou3vtKpfrM2idtUmyLMnILlv6dIGt97QAhz+i22PX
GgY/Ba84u4Dj+c1SS2hV7gFoNiRMwU4Cb3T7QHEsJs+D8qd9mXfr+wdOLq1V1TLn
x6/0WAjnnaCuy5UD/FttJTIulzRsoktYU2O45Kr3olk/YzY1qYfJWFhAUII+OwUp
vx4LYpoud3imTT70SI9rFwSKxM13+XVrAZl9+wTTyDOujC10KHatgkmvHmrX/K8S
CirRqi4fvFf0iSmG51tTSchdGDe2hQagkJsAOYzCt7+Ock2AO8tZI7vi+AoXu1vG
HWFM7fE3HgRnGAnbZ2vO14Bvr27oLLldQqN/L42Svbn6Q7VKMxWuA3PrOnHVyO6P
Q0KnuN0oJuSar//YiQ9PQMTy9aQSdBnpjQysMah0E3wR0420ZN2oPNaLZC6EFo8m
AqX6jjSV32tY1l1zvGhSZ0pJPNi92r+5i/Zl7qjjBmc4Jkq24orNVlOMafKLPFx2
b19aIeVwWPNNC2VrujRlVOso4d+NP2ej6bkN6FeyBs1lp7sWOBzd/aIetpUetaKN
3MDUOR1BuVxNBwc/OwN0bCyhQ045xzqw6x7Yd2liAWfSrNYrk7Gw+fiGHUpCb6Gv
C2zwjlAgQtZCABlUyJTEVO+bq7FXZYd5sWxOtwbdmL8XIGuT/fZHEtxv+EL5bWdi
vCo2WKJegze8Tuy38vnMyKgBhswefH435zz17hHejJOCKK3tS3brqSyBkdhZ+xtX
G+F/4MaAth8eo8+un1Hoq7ymgqnDcr0mdONVXfoeVQI22Pu50oRSNMnwW6coghnu
+BHi/oT/1VYW/iMH1XLxYfP6rxktMI4FUuru8Sn2DMJqzHzDrXwkrxnNIjCSSSG8
wZcroCUB5WTNzgDqe61rjECfe3g+gnXp5O4KkzoZ/IbLWEBeUKfU5VHv4kQTKOVY
jU4gd3G7cKOw4TgKQ+bZjzZc8oRQA/fWIgM+NtOFNpGly71pD0wAJ+z/hWELatYW
CJ4F+Ep8hrfMwbwwyvDfmuBwo3fBvEyDDzB7tNvljCeKnrwxjCLLIA67aOeMwCbC
TPIVMZja5SPkapvK1eNwAGqnDuc4SowyGiaJIvj6BAt3Go62Z5G+FiR8MVaxrUWe
ydlNb9AByjI5jXAAggga+DN877EA1SE/9S4Mtj5o/w8T2f3sGrYie0gmSsxDN+qp
3G+4XZBj3AS2gunCCKZnBMhB0gVcN/wvUiV2JDtuanMiwNuI3vvuZEuelRBwW3aq
uqioaB1DelU82xEFG6YduyWGQyZ7/rZGccj0kKeqfkkon1iP8N2NmFqihqK9TZX5
o8dNzcRALTUcffQIMJ+gEvwnVWpbR/FcS3XhwvhBZLJQGKuacWKSqTYhY/gAo6he
XpNZJv/LLs+foCYCsjI1kOGUHepqNI3QU5NAKJMDP3rb2VD/QDLtEHTHtl+Jd7fi
H66kSjfUZZceQRep1/cf16Vf6HbNK+MFmrjjqVB3Ee1jJiH8oRTXHlgMQXP/0kX1
vGfThrK+6bSLJN1XuWH7ir+rJka6wGqHAHDGIUYH2GsFutn3o6Todga0kCrQhvL6
QxCjZVXVW8/Z05xrXRQnKmm09X7HtSePYbNTX9N/O6DlTk5S2IFHtnRObMmHI8iS
oDpDzTeLKR5GFC/LAjQjxawYWYeiMoVLuZhI/cTSXx/SLErXCzd8xs+pBjBkn5wl
6ikWrZyP12aKtxoG6Gm1QsS4jQB+SbSh5XGWy6L8doM2voju0/gABswlgoYz9Yzl
bCc2LnsuaE1TSPyrQnT/xTzXLX2mmcjUeQ8Skdstn1favhTD2TKiCa1lBRZZSacn
CKOgCRpKQSSH6f80HK2MX8k6NtZiJJd5Sh182IstiZcjP13r34JU/q9a2AEi76zZ
XJ30HtXcWlYV/dGOdcub6JraY8d5t//Nbs68EAH490hoE6VB2ytizIyIUcEIudDt
L/NVSv6LqX5sJRLr1IYvHnBGTjnwhZjAsI0GpEGWeetxjir4YMHmu0VDEZSOgAD/
gWfPodwB0Q8zM8cw0Z/ntb8OP9vXsZhVwY14XR/GYdhCIb1fAC0nzhL+Jw3qQhTk
iO5X3sDjnxrWUcjtvxdNHcimp20xL3Plszqwo7KCdKfYEAkMbhrpoKHRHnUvKtFI
xIZ0CwXhU2Cprym4uWhsh9odIWhKxGOS8owtD43ATP4dSrkRxBp26cPcO/vJyb0N
1i6eWBDfmHtQEarfXmSSvokeeBsRgEeMIfxGzPoa9avjn7VduH26rcfYrzVXGwcn
A6sSQifA5c7V+8VzXfxKyYfTMtY4zgtAtvSIBy4QAMRl4pikovzhBTax5Fy4ARxy
0sxzr+M/hjFIJEMXTec+jKr89FvR4sELqooIOfyVhPUbD0ujWvDDH2C13c/yfA0x
qF5FbdHLZPzO14z54jIt08TROojQGu8VHZnb2WR7L/lEKbNlj6cXYYL2BXrpvoj4
py2ci0Dy37RJd93tCsZb8iRmhzGTFIzBTcD/Iou/UQ++YT39N4xdZNlI0kvgtdGZ
1vfofYoxbV7aXoCKAH6HmpnbybOUn87hapA0gSB3ZZVWta7r0xQMkg34ufw9KUfZ
cmXwqAoh+7BGj0krQJvrid5Bp1vy+6UykoHT2Wh8ZKi+Njasa175qY9z5/JB8i5g
1+Ir7uY4pb92WXLIUoVogIMyji/hM7aBHFwn0HfxrtQ0Xh2tju0wsdvZnShjRai6
NXoc4Tut0bSFPtwjz6ZU04ubhg6Y8LZN96zTKfad9lS7oBjiSs/9lgTRMWS/uX1M
I6Yq9ciLY4q4gaGRdGVcgPpgLl4mKuQnlyLCMqEDrRGWuNjWUW02DLpoZNscqxTC
+q+vycmRUqJhUdAUTuPo3fHMbi7zNbtzECqWdydTdVTkvlzaKJiaw2FBjWwsp4gL
o5SwxrAeyv6+9jGzagpi7cL2DyYtqZDwLrAnGexW1fF5XyCwq+GmSOTQX+v+OLxl
ZmNgmoDNd2SdYSitWj5OmJXE6ElJhmdKUtPGovSt8NOZdfWTque5Pg6MemrlFUzg
jU1xdXA+emfD/Q91vhzfD4IgIZaSRDV8ekqJ8jgtHn+9vgFK/3U6ojG6iHSmJ+GK
IvpYrozPSZsvCN3hWD9kSu5ucTA4yLEn9XsNu1sn2JfyEs41qDpR3Ykhy5rjpnYJ
r8QGSDfkFSy5u877bMkyCF2Gzrohqm+O8JQvXsyRxwo0PJ2SkUD0z8Xzo2rss6lG
5uhitREsqZFDyVhZeedTeAqJ+s7aUw+vp85xe9bCaOlZ4cprQamfomZjtN0eZnAJ
i/vf7UFW8JUgTOqd/+CyFI8lRtR1udyyZ/tpuJkql3B1oLS2zMe6nv7/DeNXNEH1
Ky8WVlCOfpNEJX1xStdjW1em8H9vFU1Wfj7muK1MJIYz5md83w4c3eWTUYzqVRwy
NvQKSStT1EI8mzllEtUV21YTA9yom+T/yketMVOWfTHnUAp8lC21XKWUF+m1H4Uz
f2RDK3ZHtVyqKJZ9XxLMMMM6ZHfSNrx4zhK4qRM0V2NXKzX2ii7Ef/CBe95U9cAY
CMIX/aIM/45ODxAABIELRENz84KtbrIPb8olUwhKaHRfwkyrRo0uxqAUVxaKDD32
uhAap4op0GU9WRp3inKGoFoF4jHIhTETrDvaG8fyvv46L3rxmvzvzo4Po5Ayr5uX
v+diXh80TVdc0yUAdpjsXD3iMnnipNxoF2KuHQYEE+uhDYuyLiS26/bOVWfcowp6
sJXKCg4MIFAeViWjKet+mImLCxJMy+7UrH5SXV0iN8rmjG9hxdChmZCuarZ1h3OK
F9SRf0Nzu60QOoQiV+KpSXi76V4XFdsN7tkvj88zIwzY/oCFO163WVj6kUBD238n
YcBSl54T9esYrVmOVMvQ70SBTDiCFDdsDHfWE4JB9AVOo+BidVz60m4vth+SQtjX
0S7nyPkFQWJx3w3iGinjso83rj10uEs94bKNITMI+asc5O1huH0RiiM9PZ2Llyxw
nXeLLe2JkT5RaaUkAk4pJdCszwQtxPtxPch90SFLccqNPKs2GDa8RIhVNRqvhIF6
yg+ptIo0jVADT9DxPmvB41JA3qkOojHQmXR7BfJFxk1pU9Hsbt/hBo3H05JRQmiI
VksQNJf/4rLisZgMCnE8JkqKnZ9lp1fxdCxa0GLXe6zSNUHe5NWQjFmpw8B4/mSP
hB2SVJNJ+K0ZoyPloe0yVnawBcTEy1oz1CkslYIDVe++nnxEcyeiWvo15k5pO+9T
EbVLEpLV8k2fxH5BQVAtqiA8TQBFLPCqLSayPMp/5DRmrPWlkJ323+TvbakYK+6T
ni2sdyylqXSnycQtnsI7TsaiBkSXAX/z3y/vW9ZyLgXnTphV9BYWISJm+Njp+EVv
tAi6fOWeQxBnVDX0Us4kHcA/wZfUmASfObQ+G+6qNUld0IqbmE22LCWIGT+uPy37
MAWguW4Ef7UKjKP5KrIvRu6TKG4oiyE1dBYLKxDonzCkohXV2lJRHNAxlskBZbMd
tMyWEKiZ3bCnaZcNhL5VkXvOOMKBsyBgZDTpc1npGRbMgBqkke2voU/En9OjP3Qq
1GvVdZoxzNPVuuKsZ3dxhzxiwgDcnQD0V1Rglt/LTfUb3edlgYFmR4NLxh84/KnU
TW1JfeDrKBHV61nmpBNEWDdu/Kb+ofYOVWKjqzluS+/xRGkNPPG9xGnoJP+MMLze
J3W25bQVH/z5jeaY0M7UBW0ADLp6U+LDb8TQttrGGAHA3LORd5np89eWVRexbhOH
95FO6kgXKjXZIWq71hExVzdtm437CBCQ4H1Suoz/LYyhmb6kDoM+ezyUuGL6K/bI
Qiy3B4jpm9evf1qPXw/7HxBqIUIRcww8MTMQ2N/k0SzveDqFxist9pCXfCuJiaVE
arvo9XxpJCKV/q72MzrnAiL5BBD/L4QQrtIlk5F/cVAPyithwk93ncsz/Z9Lt5+q
jKePkUGoo0x5wInNZvNT6q6srtXphdzLXVSzhmFVh/t8kzjMyT1jkw0PXjLu6NSD
higVkCWsFRUA4gizKmukD5lOt1g5El2aripV1kqrks6VVx19g3YygzHqSLxocaxb
loCHC5qdX9M3+iacngBuiymBpj6/+bx0Yb2xeluMTWvJw9W1Jl6ZomkePq5Tkx6w
ytzn/KnsJgAjT8agLyBGuIGIOOcmySuV5xxlhK6Do0jNpaU5zrOf8gpBJfHAzfew
Vu0PCBVC/qelrngybxD/syRlsFYi/dpVGziqJcEYv9LrHYQfUiNgd0SsSddRwpNQ
UKcxfyUbnpwhJddQycY+ThDP5EmVNMi1holuD9QRCQ4DRd92Fl5u3EjcPNITtyGt
jrrltJKt376tl89BK5ai/YGICZ0YjZljA+destY/gGMuTMjmodqCze7agT4xLd0l
HWpb60wzjpExx0nlZWp16vLE4Vtt5lPtUzhgZzlDQpqUUmTCloAuvtI/Gvu+hi7D
IyynkNfFHbLW9TjRZPFs5ErJb26Gv7U3wwPkzzqHuzsuI9fz+VsuxphMI/Hi5kB+
FcE/9JCp2AJ0wh3PH+Bdu18TNPfct5mmWCBvhIrBw8xHMta4vQqULrSHgHHZ4K4N
pWTe17CzruoW3F+RPcr6DBv30Fo5PKQbOJyOkvfq4Fto8Azo3Aq//NwgSs4TOQaZ
aA0eQx7CdYxIN4XEa+5irrE6xxjVzATEt/AvqqSSYZiDELstZEyp8MN0yoqilOjO
ezLSyXcDdYBZxNly34eT6uGGNzIqum4zQs7acW/Dx4GgjlOtOenC/4SjKUtjAqw6
vH2wN+2yjUC5mPi4Kzp84kTBodiRs1Mlo7GoEoYM9Ki/OI390piBYur8+f8YkHXO
VWZqFBrpyo/YRIcfJzgn1xjG6nn9Pz0SymHZhT9OAYHq2ID40a2KYdI67Zj35zoc
el2WPMvqVgaOiI75hYmvj3JQsgTEPrihHTOpm0Q8QlDMmVIOzLtplCGVKwQnXbSm
n676KH3gGMPOppU8BxNhnW2nqWttzQn1H57kOo3DIx8QE+7+ToCRFqD+LO97Q21W
MYlfWACucPaejuG5mNmErQilnwjuXQUP9O/nYN+NaSzxWEt92e8a6zRUuzywpCw6
CsCjprilG8SjLkpW/jKsX92AhcFH3XHFUCVphTh6KfiLT68It4Hd+8Zaw4N36Ixy
i2ruy3RyFBQCh8pAXrjE9mEx3Tm/i+ldp7A63TFLjd5Q+SZF4rxJdFYGsrziZcM3
+2c5eiiiN22LUnvO5f8vfGMZa/OLm73o7bdFrrkFymO7I/qLBlXejdegFCVU1slF
U9r1O1OX+V1A22UqrJnFFA49/akjWnpREKDb0Ndp1hWuN5H5EUlNTeBLZsmFEVyl
eMNAjhStjeItYzB4LzUrY61E4NaatYIy4YVYE4aI3cbFtnKq33V9dBoidHkVbH0v
XR9EpNK3Ub1XoF9b/JyLExhnRwF7LuWNJ+MQk+CsuTR4OEQ0UeNBIpY5+Rn4KkJ9
ynEX9aIlEEqvPkRbiujSda/kUIKRxpENIsRdTSHZ8kN+zg6gTE0rBV5wgtie9kbw
GlQtQELLjLuNDrfC8FKdwhccOOzmB7kjdtQuqe2Ov7vIQdvTEkcyZRM/rN7Ohntm
gYLi/IUM6xZBSsSbEP0WNZqZP3tkmYbSWEEpxn/ONTI4zAMa+Dbp8zDlC9iuHdP6
Aud3NJO7UazS2nItFM+FgexX9jrVt0wgPNCbOxHTz034DJl2PX+qFKskG6EQyq3e
kC0rbfnYtNlUN/cZ1P4IOBmXHcbSNjgWsBgG0hPDv9vdp5XJiu/atzWNBMoBoUBE
8PG49Toi3Gy2b1Wg/p8c/SDTWvwVRh9+I9v6XVyTDUw+yGU+xO2YZ41hWIvcw8x5
9AS6f7QDDmfPSHfs1LUoilClz75uuoKIn+EjALfNcUWbfdQJ9s5h6fWuSsJC/bkv
zYSaEp3tDVQjNURXot0iSQ9ZqfLopyrKOpwH224gpLzkv1EmOXXyZwVnQ8xqt0BO
LN/p7qIhpnD754zfkdZN180A0p0Yy/T1R1GrivBe6ebTx03f1876KoCcONfxnI0H
KKWGon8PaHvjMfeP2FLfE/Cnk8i4/jMmCmj55Sn/5GC/4PtBz3ceuMrt2Ls/zN1E
6THBkGn/GsQQcvxFRouO/4wcnx140E/JrTDUTYsv4Bx3YPbuPQYz8Ghwp9n9P0H6
YCa7Yp1PHZMV3WWhBSe5r08LCKSJ11neUSHkuOB+p9eyFWbOq2ZvnNqonqv3WFTT
2FcfKCNrc2aJdNk3HL/xHyl6itLqEQDDxogbabixJN8r9wnOcYebQquricUZFSLC
1tL0MawhDeAFnc7hzJ20Jf1wy787ePXYY8aRcX1m6bJgDeBtJs5Do1K58W1bSXLr
aOGDY8shaBtPMJuS9Ogs0ep0Koz2k7ItJ1dfSmbLobox9+N7YDjyPffd0J/jj3F/
as/CT23Mex3RwafUQxGcZnvIPViYrQ5bn9HGMEmSh1OV+SpA7WaDTIHh3eoMJt5J
6Q4gbY3OfpqU5PN9yjouKIl1TNACACJqkZey2Yahi4C67Vrg2bVdkoKvQ+oV3EVF
wr/+hl4c7QCXam4s1DHiOQwXus/iT6JkC/O8RwinYTyUX2G0Cmvz4fp8m5l1SpAJ
qGR2x8LvzfBFUtgkI+FC1EdqQ+IqeB+/hQVWWP4KnctmjUwv/OWqANbIsXAAxH5p
TgVYE0x7Wsf6//3KMDbil+IRFCv7qImv6nLPwVBdPWxaKJe+QmbdYAE6ay28r4ix
nMZdyKlcCmT9JQnJOBQf8qu2MkBWWxO9t/TmQ93S5hKr0wesE1af3Z8LBqjucCDL
PkgKrXDs3VW9M5ltqovf+2jV02U3U0O9SajqJUqZtDWtUeDKcGmwxdi/rPSzfpvL
7lJw/7OQau5Zb6dUeRjZ62fhB4p0OJB76EUxKadpuuSGvW5ZRCk9NRoBHOgQw5cz
f3yVLlAZiL64lr6Hsxq24MQ0bCC7hxzJOnV4cgc7fdi3srIGkKbZ4zrDWf2cj7Mg
RQ8r2ULMoEjZKfZVCdCtTj/cCgs5O0LjbEUzOTz1kY8XZ4RObATMuAIRZyzYruhe
yvMFskrOHXraIumnol7nOO+ms88HbywN6Nn9cBVnEHrQc1TYSifaf6f20RNvTuiI
/DAHhJNiszpj0hZSPHltIu7tmnjVcbQAfkB8EMCidgHRcllsAWXOD1alsq98jgOx
z9yi7UpX+Qs5GttS+FqeAuZ2CSodyxcRpBOiddhC2AN2KhNhw30H86iQyU9xjgOE
bempfAmeUKviZOuNhueZ8HJi+Mx0AfHFlKSZ0RATrrnd0hQMV6QBjuiXkE5GpyCY
XPeq13CpFnXzWu5rcnBC58gf5LB4aRIE6rlDKDp0W/GABDSoXY0ACDfnUnlfnl5f
GjFSmrbbsGRcE+AqvylEGS5PyRS5qFQ6B1sI3YD4C3B1ihrAadCpYOKvEvS9Bb0F
MpYlYW5T0xNHlXJGkQOHHmcTyeNRMaW2YcFskAT7fB47HmxNTDBu3lHXKVd7HLI4
6eVa72QiX6iZfHkrO+TUb7wEzTAV7da/ubZuQsKKqr96hcnvdOKpsNnMzDb0SOs1
lI2tXd32J9DT93d/nfybBAK1MhydJCIxTPxG6S5AutTILVhneFqLNIU+BBUwnJ82
NnLbN7Bq+o8ZXxNg7R4nNFkz0XzB4be2VBKjLHRGC3jfD7BHDjWolcIVXYNJdcz0
OBsJhj1Cx0KJ/2MwwJvIzDTnGA6xYnCDxZxKT23QQheVL+eEYQ4f60XgURGv/Hcg
XafCgbutA9S0oEohm1NQXk3ZNYiZViBV+c7iE4VnQ4TKjynNC35QggepgCaFnph2
euKGHBBe050TaleHaioZ+DjCMioxpYrvPFRcxfEVz8u7W1XwpsN7Vh6v0hoVJ7r9
HGovN3iUd0LuScw1hWKehefj5T2+2IRoZcTMRUGqQf/aVwQT6MvgH+6fiNFF441s
rn25lMSa6gjNwMn3nlFuRenRKXp66P+5hIxgTj949EISzyvpRj2pzMKmczbtU0kC
Rd6LOXncR7K4EFXaequ0F4hAViewUMQCNye7G7/pGlQJkUsIa04zX769xVmNDNFF
xN11/ZWGWTNlze2w5KgSeqYySkTxpkpOOVBrupw9w+CXWyer82igJbrAswfdRT/5
mpxCLcTvIkgT/uVVm/WjjXCmcF6D0WBha7R6G3fzrxeGbtpkeqf9DOceDuRlkMk2
nBh8eAewp/uxXBiFPwiZfDA4wIZkPqfG7vji62AwJklWOrIlTLOpiMJwQERDnuPH
WtsP+6DwZ87O1bDxJ1z6aoDU2wZHlph878hgcN+rt7YAN5AQDlZMULa0STSDAp84
4y3Vrce+4jjDVImfghR8fZg4kgyua2K4McSD3FSnduYS5BpYE91FxOXutgIgH/08
uJJbJ7j8jN0jexBTyZ93WqNZJIbA2lyanh5/fXjCOaFgTy0PhQayZfqvZKOLg++F
uBetW9u+VC1NjyfIqetGqgZDgxTlpV2j6DzxHpIEQOoGDwPbqg335hZxKPD2XNBA
lm7vWaoxaUsHa1bmvG1TA26qP48w8L3AivlvEOLkfnPDa8GYNMRDLA1d4gN4zB1+
XGYa23P1qUmMAAVYUn84jqEsdPBQlF7539ll54DvfkWyvfGFvTTlQS4hDgp481dd
qLTQhmYdoXFQ8hgJzmnmFbG/9Hd67d5SHK832rQ81GcsoztRinr9vTH/Dd7RnF1w
3dCtYwrn3AIjvrcm9VMV9VJCMPZOp8XIz51NJ6u+cWGLniO7kZ2fd/npVZplcZRk
lUBhr/ohKcHPnC40kizAOEI06Avx6muqG7LJvMivI9/tQ/92TGzuVQpaqT2yZ7Iw
oP1o1poBewYxnyndmlPh0bnLW0NWJIEaj+W8yIOgBC/pwe/uhdS9S5dL777ssCQZ
Lgl+CRFZ3Vxg1yQrhP/z3GuQ0KLowRErGQmvENTQQ58/6f0Bc4RTGGJm7F2xc/tc
HWV/AoDVCa0zSoWISVGlRaoV90xsbjEbQqLGv+GH2lgJkKQ7MPFF782N0QUAdgLB
Qu+Xi1R4SGA0aT4/KfhRh8ki9kSYK0EPrYK2ejwXFZV5e6Dc3AWuBckeowrgZnca
e3ENp+pQvvFp5MaqI0/r/oXjCj9xb4tmtFpilwCp8zHQmZVLBRsjps6puXepe6I2
e7K6lhW3K77KetKMJnecXApT2mRHn58bcX0c5Egr1MglJaWJAwcuLGsl/9OKGulL
rBuJeAdBJxy+F7mhYjH0q6lhWruu4vQWGP7DPi3EVX0Imn2kJd2RPHVVKbm2ipjl
N1hq+87HWpH0OvvNSY8ywfTK8YFQw73pVqt7782MG95HINcFNCUjJiy/BwvxsB2y
f1eUQ7pyXCC5No/QAjoTJGpVSW7jExfKhZk1nMETEvsSSFPiNLLi7T/rbeR0y8Zr
ERN8Mrj1lcOHMtgHuz6mgqJJqevzNd/J4CyWyZ7pCKCmUiLAuSQgWBS2vxCf2sFt
qtdKH0fl1F3PFlzNBzt6Qb/sg02MSULmAsOvJ4XQzb6rV66rrlHClAb9dKFQ3wFU
Vup8KCgzwAVGSggXEwKq+vaxRV1RQL2ZdsyyxrUrTlU791AeR+kI310R+BBiDt3l
EBJVDdcGXwL6JN8yELzuSBioYHIwprIAnjVLn25FjoxevJHnqaWYO0ZVv3R78P2Z
shs4plLv9SQMWHfJoTFCp0oDaCO4oiRQUkaG2etcoKIO9X6En2BD9ODWLMy1Nn6O
JlYHKsekpmfhs6Uq8NP3KdIlfVm+l03fYORolBF66iH8up+7shp28jJprXu9lD+G
e55h31qlfsSNX5spJN8cc/wfoR7UjvaHGX2RFE8A7xc1xzyYL2j1RKewfME+7atG
gG7NAsM1DHBGHpJf/51/EqnLbHb2vPSBg2SRcTlXs4muEfvUG92WJ8czPo1Lv2KG
aXMZIpRRPjeNFwerFzGUGA8PjXN+TmbHmDIysw0WbehsdLwBr1bSDagaHtB96tYO
fDX3GZ7gAKPb7J9Kl7P9OI51kyliWFMBECO5josBmH6ZkdRtlRAdC0+o4tybWsMR
OLHtsjL1sZIevzxhiyFUpNjymtLHRnPAOyH+OZMoYrz2r2mGjmq8T+AF/Ujkd05w
uU7Wf5fuy2IptE12lzdkqUMuIrJL63N6fCWrcVCw+fGgTKYLxnF5wU5/uzZW0rM5
trZqhtf3bdbZXIev9WMgMsqVH9o/kU2vE7rPz/B1yoPDkJqy7bS66IpSzRKNqHkb
BlQXaE+cYXk+lowrG8hCOXffvURzbQ3y2PBg78RS74EF9Oq9grPJZLY72/J3zKV1
+ASLCGV30LjeRBlzs0zS6ViqZCeH11X79Itg14J6NxuXmXrslzL+XEd01JVdGZHl
Ch5ZAGxAdDphtHtdvhSZMlrZ4RUmd6UyiGwOLFqs30ERG/U+7Ulx/rBt1j9Qzg5T
nsD0Npn5TZB9xJ3yUrPZkmbQKSep8KvjUVT9m51WNJLnku8WBM9Tsuuc0/MLT5Nl
uWq9vZ9L51oAcrUwwhXX1zPaBNqSWWmlLcq7rpEZRq2aqEqKivnR7DgC6GUdZp+U
/gXYkckr303d5QyttwmG7JPCxEzIzvkzYwZNbWretvEmYASFFbcFND5CIVGqnp1i
NutpRmqEL1g8znWVPr6oB+n0a0k0EXt45hoY2p5MiOZ/9UqbjgyTGjEpJPmxodM2
/4PgzTUK+k9BhOx0lvj+BpvXHWsCmdJYdrgf8PD2UGc3j/KpcbA8D5DETC3f/myv
Q0ufMqb+QWvbYnt1Bx9k0GoVFquolUEyiyCkHxkZyrncB7AotGEAUM2c4OhDYOYT
eFWI+J4NAHmrL0RCSZ0embBL/1FHMi38lB5k85+aDhHWngv/p81tTYYhPh1dwoxM
Z49W8/R+MXMETyqX5fNQDw8dRCKi4mdJrX00hFI5KBJeJzRdc13tGycqKCBxjRMc
4FPo98ZqNSB72+pW34zhXKxAPgWekTBZYDXZs6xcd2cZcczr6596dL2PUG3Y25ht
H92JwT1sjl7T7e32HtmolAogshiMnXokojyAeTWV/mnff50Rti4LgTDlVy5ANL6v
siA5ecqMcLZdevKvvs6CtyelYBClY6PdpTIeaFUF2RY1ToTckwaMyzJjDRylpngd
x5/p3GZLbKOuZEA1M48C8R6oDiFz6a5KdhVSy3R3tly0i2GDYL5W2qOouPh1F393
RIC6C0IjAPq5rHJv8uIC60Wk01HMaKbvry4SAxZk+nHHRSCtoz6CNFUtUuDRoEEo
gWi16xNSDdJ3052wuoeqJhN/sh2v8zvCLkXZAJ4VtSpzBluox+GWbBo6VocVve8/
za8XmcZdMwew1lkqBbG7xOy5PdpqHiFEY1+R95bh6cTMWWWL9FqmCQdInuTltInG
cywVHpJ7fpFc0qJlCawjljI+xW0QRyqSx9TOhyGdxGWKow6BW4TrmEeVzcce4uzW
ZgerRLjpfRtxNFR0xVbdCZyRzutug3Y6jus4dx7NSuBfBWzKIbvExzqSZx0bQoGt
2/5uWvsotI+7DSf8MkO1mAHHcXw23kYsTiIk3uRHiHUzzCN7LZsnIsVBLGLw/+o1
wavOu9xGWFQ5MfgDROmvk7uMCPNUzS/6GLLqR6K6ZFPh0U4jIcYa3ggIZkIDgDE4
99QmElGycRQMaRT06ZamZK45LdZDHqfOtz4VI/X4HE+yRctPc+nC3ajvUWduJ/5h
r57K6ydsyfQAB7t+sNCBMxySUsnFAq1sTBqDSHG5mMjxRW2AnLztslfD9uhZKsdO
PgZh3r3T8YMv/ObX74QiqZg5JM6DTLjmMua4zpdRLttwmZr0eeQo6gFQpX7ggg7w
vtLfML4XojI2hjC+I51KV0YDUTJqazkMdTDlk5S0oLAiDAOsgZOCyDwlxYhOs3BJ
gekHNkt2r8qS7d0J7PGrTLMTPeJ8dylOnFOkjeDXpcwUCZr0UmOiPTbL+1yXsAIV
eGCOMk+aIJm/wznbrsW1mnyUq78zIPCEER0iz2jouEeuv3ZLerEMd0NVqv1hQxYz
6IbJihTIhkZw5bT7KpGvmJVyhNrJlF2z0gusFdY+Uwx39UlTPThZmq+6aPQTFhlE
hhTL3A2T51+N6xcnsLrablG0hmfOAehp9D/qXWLtBRdN2JNmu+39nr8ogQhQ7rcb
52iVt9hTTr7ufYEBjFSHdpj4ZWv26o79tpX09rYxXVbXTdsANXV0q0Mz84Y0l5zF
Xm5sgn9JUWOX8oXcz/R32eA2zA2W4vH/+pt6SueZAqqI5/wOBOAH6bPxG+eT4hr5
pmPHRiXiphYv+t1dEskxu+7UFo6lOFuiQpU2M31JS+b+B0jHF51ahUy5PmA0YvFW
BLadg+zKFJIsSh1B6+PI4FQ01DsivZDfJB7TLROMyjEY/spUKKF5z1d17DvO/EM3
Lk9bLeiTK94R0v+XnDPtW/GJ0cugC8C9lGIXJWXBOvtHMUGcRwViMkD4gTc7ExoL
M3vxkON4xJd8n0J1HeOg27H+ApH7f8VBNplNyjl3NCB4cqUXGUBg8vCVxcyTdsGy
7fwZsA7LY56LXLFkdzPglIVWlRSrnpswj9hGWfK4qCTr3c17NHtFr6I6eNa5+jY0
ydNNYpZl0KAtFauzoNP5lMXo9gKk/rVoMnGUxFrT9tB4T1LP839sy5pnE2W52rvE
FqMIhGEcf19w7IhPVAFStyNr+TBFopaJ0WnuJ8isuD0o0lgWrw2ehVNgw2MC9Gsg
1E4B8ayfl1UAe7FqQf8tIw/r4V63/TMFF/7b65WQ3B6QUBHUxwaTXjLtsHi09Pla
i3hN04AHWqkBRojwQ0Qh/YuC5zbRt2zRz+mcgVl+3z4MhxsTbIrqbLCZl4c8p8SN
2rXQ1lM9rnq0x2Nezwg9c/eCSU2vUyEKvjB38ICl8fKyRowtxpN5/CWGziqoSFm4
451Rz6L9amKxOv98kQN+gkP7n9Kfp4eEZFfzEkDsRbHcioBcKe56cUcyJUGSTMnl
4AGlYfGHl3mATK4KKJYhR0XK7Z5Epymkoyckld1XrVWQtCyn+Au0vZysZF+/r+F2
tbcodRmFcTXDiJI+WBJ8KEJ2xizJZ2rJKdd7F1WKrvtMV+81nUGQcw6XgDtXjuSk
pq6nqT00ktEPK+lJ61tcHeByj9sbJg6x8V9AnJII7lI9hPsixjm4u5LdCGb3m2Zu
ZFQKTIhV6O1G+nBZ/Rp0AAFA1mRtdczulkykkYqno5qZoVtTwT8dikzj008MBWhJ
qnGthMNu5DzujObrfCtmMVaPkFcNrpzLlEAG8nZPI1w9lh+7hN+N5Atz777dWDEz
BhYy+cXqxTw1iHMwSouYEqdiCJEHD4LRe0v6dIrqgOtezMG7746su839ODr8wPh5
gXXqVFIxOGzzfhhw/jFPk564+BJpt+7P5KRsemHmBChxHDlJXT9VspzCthcQDvs8
e+S5WT2a/24KqIehXauVms7pYbjADJMCGLV7/J3kuCVDjF5zFtGmSjVd0CiAvxdN
9Y4dl9SfmrqJ5nu8Tqu+ETclN2uuA1lVsrS15rpmfU7jeghUIzd3QoHn62dOR9WD
oXoSn3e29ZSnmOWLDnmJeiCR9T9apgjqLsGXOox49BQwofKu9nSYmrIQXCTFlSpt
2GqFUEsGO5/+h4Uo8px5WU3zW5bmGiLIVHl0Jd/JBoTpaS/iCn+l2terZEPkvhsL
1BiAne8mIVCmqPM9qeIW8lfY4cKkD4gI1gwrXU4PcTm/6CYy6iIzEXFq5OE7Fpze
6vDXhyREv1KeHqiKaQ34LhqjmzgdDmfirNLpx83+7IVwU29RMuR5Vk75JYMEhXqN
pPqEpJmqzK+PsXn5xEHJEfOwINxZTrRP5KeCFsS6v7b52SFZN9CuKVqw+Oput44b
DL/K6pcGSQCaCoRt2OLZZxBlbSvEf3RX7wq4heDT6LdpFfXSRjFBG/VWv+h0w4Xd
67HDnYjA+yEeVdMobFbMTCkxeDgwK+XlTF/afMRa0y93iKCArAId0EzJ3Y17SxcW
I42Q3s9609xuZb45U71cjjvTDUFK/YRbzllpnUFELG5C//E4GWRXnEOlq3tKVfyt
ReD0PuMIAwOAeP8KIr3clYHlJogYFWuX0ukfZUqZR9tDZ94tnsJ3+khSTlnl6c9c
6fWVeMj7DVw1y6W7q76jI+XCQJJ2aNfqEiWvf7u6BfHhYBgdwlS2crDv3H5Opfdl
cJ7fYhVSm+ZwjGN5CdN8RZjxyHhauYBPz3QQEmbLmg5HbtI18hQVfWs7spIsyWpV
IecJOlA8/uF7qlJDFFwMBbEWsUHwFCvMXF23XZV2uk0j7Vn81lDDOCjAWwoLILFr
aVn5ShP1FLT4WK/W7R62AvUuqRPXxKrGwMCMEniV9+zqmI/svxOlCTYq8xNm7Jvr
kf77u5asG2araspTQmplDMtnmjnyx1Rtcdpz3o7fzGw99Pvu06B0EJRMA0rTh2Pg
LFyvctFZpsxzT+vnbbZG1HNglz+f0DMe0rPP8cnCjn50p12vuGRYbupCcYHHpDcS
LVtsXIaQ/h6LTUKvOUvFYuQXOBc7YhtF3PmU/7yjYbJIsM76vH9m+Rhwsm+FhIHo
A1n7Oe355eU7RXspCnzEmVPJY6dKvB7C4q6KlS0AqL0x+5NOApIulayp5wr+9Xfj
ZX5v3uCcnD5GWaFD6BYOIEvqMPn4vXVMcpPeYQ854tU51GdxrGdfOa+lATekjI9m
Q/69lP7K8Dv0ylm454PxAb3EFMyZUgRTxItQyvB1PRLHGz7rXe78QWT2zsDNr80X
iL0RouO6u2hosW+5+pB8L38ty+U//BV+GGZligkDAiKo0SymiJDisWI46lrdjBHf
T11QZUXgfmXQo5j7SXjuscPN+9jyY2K0eni1g/taS7+UAqgbWfWtTPeYR2lGSmsf
mxvgQYLfgNIsWjQrbeF6RUZyW/d6+f2Dh/PUKCAUtdahd9N4z/7JYgQuelAEW7Wg
f5hxUMc2DJRWg9q2Mz1VILrBIMfj35WbAaPIZdRCACBeA60iY9ofRYGJIeLD2dLG
u8LfB5G8WMUBxU3Yr7YXAOx3zQJg9ZNu8v9dyjKNHqOtauSap4jd35Xq7ABIfPff
tqaPbIYKV46mQCqV8hNzzVEmjknq1YNQIorg2oJYmrrKIzDw07eBiieVABJ5mXcn
S5N01egUPBdSXZFG8u6s36e0keD0kKfBbjZpnXdeqLfDfkVoD3vDFAH47HaIuW2I
6j5Giux+x2ZokIzjFKiSH+iD0fAMFMa5SseorcxTGjSkvDHnoDgjfs7RYw0bPzuJ
03ctHcX8jJTzr9sPVyYDpqz9qZ+UpLck+QM5QxRXxhpp4ze1sHHmG88MBQLGxcb1
6N1wR9wfP96lPndliiA0exhLqJe7MiInuFvm3McuVsPhBjYAWQUwkRx/yA8ffzfE
ndvnG5pJMoC5HxH8VI/qtVIgC5xHmqYO5LWAA7PRXVOjSLZjIrhEKrwNI/YOLTRJ
RaW76EzrgckvFUgyRh5Myq0+ucj3GHjhXsx7G9xVjdh8tRQ39BCNR40yDJDWbI8n
OvMzVoC3oVeS9cxn3xLTAckPV9y4nAgEiFMvnwYhNhbekdXbPpVyg8rfgOVwe3ja
6WrnyrkfO0H8Rs98kmdG8UqJ7K50nMnIY2dEN7m3mMyZtc8yisca3e5oTHBGn7RV
tzxyT1p0wXLaziHG13VPW/rJYtiTIK1SlzrFs/Y5hVr+OSClpfOiue2n1bGc6frU
jnFd/74azcofvk21KB1+D6hA6mKCsgRcMXlFEhTPOEoY5GPK+TotCDj/06/vQ/MD
vpwi8EfUXtQQr/tUGXCwQEecaG0feZxQGhozGhZFLh5y0eRCN5D2NYB8HBAklVrp
kTPQMzZZ2SETI+O79OByA+EQqFxwFPD/3NrgMHSaki7qZ2tsPa3gHX/96YdUpPPR
UJzb07f1ebUrkjN34Cg+mdUX6XXTKnZt2BddH97gE/kRHD2nghEsx9rW2FFUsoof
SRBDC4nsXAB8scMZsEEFBSuJxhzl10KT4pZ3l77rzCaVNloOLXEou/LFkqlQVW5P
YMGqlO3TuX3f3HdNuBsQEM0oTIO698p3l/HKc1fgFz9QkvmAWi6aITF9uZIKXmy5
LBLrlLS/dH6nqAzm7sNOhgneoMH6Qy3cAARw1b7NBBDak1eaIuE5j6oKitCH/cpA
2Zg0ULDmXV4B7R7NWJ4fnevyu1mJRk74/O9BDYz+CjkZMYMocam6cNobFvIZzsFQ
baLTjuDBojlFwBKbcqVVuP0qCaYImqYDRb+TeX0+OTL4s4ms5Cubh79nzL1o8031
6+8a3uAn/xS5mMy9ziItTus8evivSdP3bSuqxOfmzIdsND7D5111gmrWEDqJkEYE
dAkBUbs8BlHVKtSMm1Ps+jSJHPE4W3MiOP/r2oVOmVOHpZRL79ExeksBa6YDOOhM
K+wciM55Jkfn9CsarxgqYbw2a0lfyKFH+n71VvFQD3EimZtcom/tX0L1lG9nfJMt
N+47E7KbOxfFX4VJXwwXjxrJqvzihNaZBSluOy67hkZ46QJFniK1heOZJRVNyOwV
bT0q+9/NKUT2OOxCucOciK2t7Fm5SeMnGxW7UQEDhnbMFK4k5ohgSg54zpfjDEqU
x59XMkZfsG5sV4tdgXxi4YT8xT5vUBvpoKLqdCOoqzD9ntrGVZaqw8LTVXL/juhN
WoizS4E0zCoppQ7gJ6LFCMsxYfB0U6w93n0+uTSeS5STw4ENbmOGlvVZhZbW9o1r
SBJfCtVH7YIets7cywyqQSgjgmyKEEBdJzwquWdkVOXqK49gYGZu1Pn1OU7N+Epz
nXMEPmD/50rBV72o2yUKgSujPWHABT6ziagFTmZvQ52++LeFZ8xVdhi90s0EVrzY
/sOhFbqVMhwXNCsKXt8NOpPuW8yU+aDq3bR2p9NLX1Y6v5ku6sJgoWJrGXhTKerq
WciTqBC5rhGU9xiQ5AkiarZI77jb+YV1PZAGtcyUi6Ax+0sXMb449IxiAaKaDpyy
FLDuEnRsyERI5HuBGCOO8uFG2dXEH+BTpW4AZlA3cLMtzIam7MYTNvZ/Nl5eCY3t
EoKiOEdeutWoPTD9/D0YllKkQOhj1Rr38eLim/fIgagEdBQAuR1Ju9DMCFOJOgcf
U2rONXOR2uj/1Q9ZBFhpmMG5IMmi0i+h3iEgdXNmo0vUchkTzVCgS7Q71hT/ahpH
ljGY956yNtTEoifsj2/QMN/s/0HTkW1Jx9Lpsb7jKhGjVEIihlGbRiZmfvO6YETn
cfNYXfD+VGsxnnJV7LQ6fIGY345XNLFS8foj3NAEUcI5nsc5p52vDxrd/4jKG47y
asaZ0v5zoKqU2KzHn/1rW40FQiXao7tK1JCy4IycZ1tAyE6EohDTx6ryY7ieN54b
MhV01nLdisPLpuO04JEAxVekTWpCiDcICpqDvz52+2jYMeUWF1y2HVdQDDZ0SXQn
VsuJ7ORyZuvyhN6d1sl6MJoXDh0OCpVjQvCVPEn+hutVsn+Fql5b8z8RTue6chOx
/MNMnKbxkX2n7XtEGKKbv8qV4kdUID8LMk0qx3M8C4TX9j+i2L9rYrcTXHuPXZyq
Q2n41VWaeDQqgQBalY4BioFgcSvRY4XFkcXIqt/1ZJX8e2IHuDx+WviDaMVpbqdj
vma8z/CGy6FE5RhZu9EgEmkkUBauWk4nFeQhxiRFR1Ys26Q/I1NkCrOwlr7eb+UD
cGhjCm4gsz+7Zs4X9ju77WtZaKIkE6zyETPwE+pvQoh39869LcdCY7XpJJQWpjyH
mVdde8YGiHXgA9IBdHSkzGIdTBh9iRvFgKUn+ZTtGUX3e0lXqlb5uZe1+lC9lAXQ
fwyUbOmpc9AftV1qs8Wkf1tdMaDT3AN+5Hb9c6XDor9urTz4AX2+R8+aE5IMDRyJ
cX+jImvD/litlRYpg60iO6mBe3Ix99qDIF19BMLL7MEXVx0YIHGMY+30BG9uKvHa
rbRd17+A2TSRfNMnePioBdxQirPmsLs2xSkzaBcIm75WxVuF2p/FAX9TDB4ApirL
G9p/+LAYYzTs2o6pU2TxEYc3MxG370ubcI1TkeCPpHM98O5D1P8u5c5DD3PSQebw
LIY7A6gI64cw9TrTAHYGN3AR/eRtEVB1uc2x97mxGvFYrEQjSs0z7bZjXvLArEzl
iybYjkntTvGRiCPPrkWjeS+q2KDdes1NDZiLorB/VzMguWA6DOG738VWvchCA4Aa
7EM1xWCOqyLPQGjsS7zmCbcxnZFWa3ewxTPa/x0qWiE9fauVKQ7wVY/nJrZZ/YJG
3DdE2FQcs22/6TZ47oZIhmKhRcB5pIQcfmg/xFyyhZ4qGtaXjES+Y2t1u0782Dm2
LVNbxknSIIFWmwVmJV98MCc3ZiWYfcOw8aoT2wrcKzmXDwcmhYQee3bwuGerDWZS
ZVKuA1ULpODqTLtj3tqzbrK38F+aB7L/BEHnmASy5PCoggyD8Mqjs9zxfZ55O6uc
GX2eMGP93b4xR2/pjoYkM1zR3ArtEQj/JFaCB1G1rNbBfmmBznwGB/pQQkEC0Wu4
mDuoqLGgA7TopzwQ6oVkvbBYD+YNWfdVjJdCAPnb/ki6yDPD/QRxdnt1JYGCyrTb
zvzHXTBwhJQMKqDouaLK/S2vMqc+hULDzHCuzEBbGd9aMpTdDRAojVqF/bTZD/4U
prfJq/OUL3khdPAM7VTd3oSSYyNCZcERShcmB5sG61fd5B+3RVY8ww//4cyu4w/z
F0ehK/JyryYBQdolWfLqkC+CmhFtlBgGE2ZR05xoy5pxgM7/T+mG4G+tg1fyCiFE
a2dfftqR/3a6dBlydyM/T+Y1m+JYejCGmaxSEr2i9TNLYAdDWtf8aCmxymnawl9y
e/iwGtSRpQx2U6/U0YSCi+iDI+EcBQH7JjcNneKohSNtN03XSJU9fvyO1V98E/w7
mPgcsnYEz2HKRjVo+BZN9IVeb19DJr+o0QxlNx6jPl6odGGAYkO/q8CH8VNpacdI
R2p3kI8LGFphLnxi9EZEKgyC3ZjELkWyxp9eitmiXtVy9IF4Rmo8/0sHVVqPaMfp
rIiGeI+HT1eJxTxJZWbqfKwWjGZa28fBdQVRBasnt9u7jqCPI699YeZBO/G0uOCv
9ScbCzkt4uLGnm2GZ7KFxWrHKp6Rh7yJSOxYmptUHKo4k9fnylmw3s80QLtOdsQt
N99PSOjZKYnp0bDAnNpBH7TNvT/4iHSJaWsOoJEs05qkyFUh7JrVKij7Oq23I6rC
pGuPhJhcMY5R74PY4hM0t8zV6WntWGf+PIOcq+RV4m4/BiHovTobwp+56M/JpMeX
lj3AWEKmOt2+ylATPv4k3/YJWMH8Rd8rdySJK4Y9aoFjmT+SQNZ9XLdXpmi1MOeZ
m7QCv27NhG5PWr5xsLf9ZoA9ILj1YnjlIinCuRlxIf+l91fNlKrf5WwethfrSGi6
/je5tqJvfyuiFhbkViPm6aj5QAZrJY3x+Va6A9D5rL0LLveUI1Sf6kiZfsBj3QDa
kMhoND3N311PyzQCQueltufWZYLsKtUr3UNn1/2C6ldTm9clvb8sbs70BEmTSIgJ
s4lwOJT7EoDKmnzfb1ESHg16xY4GtVmiihFZN+QqeGAy6o9P7bl9jFXJQjyXzNk/
NV1XkowJlct+R8G//zqZP9BIp0Vzk36P+YNU3MyNRwMRwVxw+GNuVfYNR199GNzw
FkEpxG8abU351LGHF+6qhSm5iZt4B1UbWaT14pnfTLLrYywgiDQiLtEev1+JKvCw
QbFIrq7O1qMIMTF3qJ2aCMVNQx9uTlewOEvHrURoyYoYLIHoPzFnPk5Uees0CRP9
NucCW3dY2gIEmsfn1DSxanGyGUkRssrDtFIuO0po4vEWpyYJP2IXAhYLL0b7znhh
yPcdhJ9ngNCaJdcnPzbJCqgwoTn5tHlv0T/mds8rxrCEC0K13yHOG475LlIAns3W
d5gOTW6TJKmS0H4qVIR5aYRKQG8so7CjzAftAyQtzOlzGXBYRSMo+luepzddS9M+
xRPCcCpFZtpvKdXHIQngyAzGFgdzKiqm1oyfaYG73iKnFyxsx53iWRYBUw4oFk0t
1OC28gaJAYdSINVUKUGYbD/sdLL4UIbAU9VEwbxBucBTtFgRdGGgr4sN/FmZ53Nr
px4QAm6habSZwVOd1x1ptK6gXISEc9ekMvb3Fhtc5rwGLfUHXScfYaNSztFjPtLO
VoDvdrZnLxCut0VJ9q2/EpiZOY4RyC0x7azdyfhfDPyKXx9Zpq/61MOc4OS1sk4Z
iso+gpLDeH5BVkVsnHaMyj30n0DsJI4oFyIe7VGHN/3TRBNEncjcRuBBE0CaHLnt
ZFmnVaus1M25xeawLCtbuNSpicPWzOxlH1cWtcGdtZmlO89D5Lyx+xzpRf9lBQMT
e6YVhnnsCAbkEYgSP0+ijWGUbrjEFChNQFz9qDqHAARlx2ItbcKIDZoGtPllSAFV
dy5sBZsYyjEbKqTIWN5qWOiI88piG46Wsam8rHhQ2+n0FNPGfGQErZDXwwMLQEOQ
h2y4A/o/zukUinhgo5Q7sUl1HL+N2Y2kr5wqESHAQmKQTM+HMtdbCruQ2v9AkRhu
643Smt7sGaEsqYVBi3hrwNTLUeITJ6BEQPSz45ChOpIeT1GmiveNo+Bi6ky7vDRq
y50+PvEXyMrs+qJQxWg3H+KUZHamip0goFRcaybLonMaae8P7rM2Q7UeBelukHAM
ePJoQt5FfpUBm95b+tKbknrDZcvySYNvKK4Dh80srDg5at6i9JMb7lnvAvgIzDNd
5e1/HXNRkJadN1OptMRxuncgFacKVEVVH0yr1dAueJcWPDcSqgscOP4jofO1t3zL
1QJ1OK/g4y5bNZV+F/UVy7UIMc35Zv9PsRvi0lFMopLP02phHmWCDkuu2E+2Zk2J
aRd7IgPmtUY52UZGfAa81Y6Imd4bP1x+O3BHRAmA/WCRTzqgcG5cnSt+NgUWT9xk
f5lnRuD2mk7ZvuR/8wOANcJqwz7/nCwd3rz/xTyDIIOG1PFfl0al0kQ5jW7O79u5
v17pI9nLaxcwQAne1QYwJ6siWLAs7hBuZnDImlqIDaVzX83pGtV0xcdYoNNCkIaz
Qr9P2/js0qcTemobNOn4rgtv7AX6DTT7nXdZL8uSaF1bSsCUj+XlWfQXS8AdGxV2
4RyqfEBQ7V3mzWNE/VQiLxdFR1V5lxjH/SY638CHYO61HUgjqJHGVZ6IT5hIKbrm
NC0RlE8BpQHzOubItcKU1ZLNOiTcpyRPhOWezK9gMPziue51H7cXQ83G0leXYAVz
TgEJF6Q2h1RNIbHT9CSNRmW9PdH8dCzKZDRLdK/UuL5WoNK6BhVv8pMfswRpwjNz
optgd+2qDBPmtjcZL/7iTxwJ09ZaOQicyLsDsL1eeoPzkNk0MQKKeUL7Q1cCrgXW
XBvAE1Y/zMHGNqpm0FXY5wLRKGXSOM91dUmMydoSOMmznCtuI/yk290S6hc0A2oU
J5DAj35qZCxzfs9xSLJi/q1wJCPjmTz1bGmxySDeRYi74qDbnuo7ZD7KFTtQMlyq
EJfogzWmgyJ7XMVOJjDOzQoqUJwZA6NIHHjuViIb9n2TJkx6HGFuqq1+NEEUlTSP
GRyQdpLyGdxDGy9YkzHUXzfqTrMkSCbyulFuazrw/nWIMACOQaOb7kgoNkYivGVa
DkUrHU+lVGHcqI5RByQsNPUZ9EPGgGGXkc5OBgPVI1eh01SkuI8j0xKWg6OwKeQM
mXiFKmv6OQx3IObBzGtVj13gqsSLiEfOh3zN6U4TUcBneQaowJrQ+z6YFB+gv487
DS0DZWz15TI7pZmk7QbLITkmkCJ5JuXC4ci9cwwEd2r6byiiHsSmIA9JTJUPE/3f
qQQYqlS2hDVb9/kH45/VG8rtijQQ8CJfqvgcGqBZ+MUQ1wRH6mJs+fYPbcWi4Z4+
epEObiHSYeW639N5uHfLpin2+bMPdysRcwY+dkRBCBhGLNSac0zE0qHKJNaMLu5+
YZg0xebbrvDmSMN2n0ml45zygVnS8JbXu8w57SQn+WD2pz4XI+9fYtQq+XwZc0Is
Rsdo49D6kSZMM6yWgxUbLDnbpqsDvltPllKcub0RZTbrq+fk51dYgzQA6fZVYt/h
GzZsp2F6xcaQtC/aIgsJrKs/DggEEOAIzpcEmnroM3qr/1mWcTvEoPa8lsbN8H0v
7hFOAbVFLWWSQXIFU8COQNHYfUfsY2ZxnFO6zRxZDboE3OGNVQyEUUr5+4WG6Yjy
IfhNQ7Jc+Kqb6ZmMMAmOrJwL11RrTtU7hE73E/H+fXY9YxQ23+FoDPRpXbbakwOu
bjPoSZv8yfWqrac8RbCsvEBBxcszKus+BVkwOaYOldlvojA81WGDrZkPRJmFeZBn
M5dT9xeIFKfQ6k+q8CGFbhbVaiu8pOyWl+/1rvO1mKnf6YIoWd8ntQhsygFClMIX
PSoQcY4xCnKCN9o1Wx+48xuAIrbwN4EuScU9+AMf3rr5fl2D3uAcPcJZUFbxmk4S
TfuyTpgbg146c/sC3bZ3Zig0gtmlGrcRihZ7ysHU+16QbHejlO7BnqlyhwPzBkwK
qW9dQ/RTf/zFTkyplvmzmoYegJ2mzSlb9kZSuxmU4u3RJI/kqpTTdkO68Tzq57Vu
8QYL3H44S+F3JzLRiwtf4OfMR3VUqGal6ke1Q17O3f/IeXnRjkUzWqYAfeNA5qvm
m2UlRIXf+9BOrNaaPRYHIq3jKTgRQHEkz/rGZ6Kb0Bz0cLoS9Vq+3/5+mmZ/stkn
7Ili4c5rSG9iajcVtPkW3RjmycF5cGzKpes2NQmhch3RKGA61Wjk59A0AVlRn63v
l7Kek5ABpZDUgs5/h53qZGSTY7Pf0htEZll/ftTWPoVncqgFTZPiVf17yhwc+92N
B3jKREGzhjcnSwEczvIp6esWCNEdV7i6c7gNkV0xXJzRHoLB+61QdKhaLsXF6LoO
uHSzMFsIvDZfeaMJHLgYcwwn5kogkJEdNDlPaGZSw9oGjItvORD5DkEZ8lAcavxt
xICKq+LRpFXNmq8dprkyBgJZlx+660/c9Frl9EEAiiweO8csMu1Z+iSMb6+cz5Tw
KL0yAwc71C8YEGdto3QSOBKiOubuQkBIfbv5R/5XWjhIPUcMPN5+A1QIGc8x0hzU
EhYGq0fhVSPpG/CuQ2P+H66fh2y1vOwRma9WguhnbE1H+GMswEdjc1ud6/xwgrsC
n0xRgEh1tLswtZH9Ly+tJNS8gg/b7+ww7iKVG7uFPl5XdZtVVK+3kpaLcySgpq20
dLpsZoVaeI42M+ONtYT/hCMUI5pQEVBFCYFFDBM6vVOHhN6CkF2NL8Q5EJkv4Vju
7ci544Yjflppxl8yVzlgOHL67IPMZRfUz3YCArMQ/2AXoeLrY/ESu/wpbdZr9dHF
+sGskm5DMbAsfe7D6TOx7641u3zbj69ui/9ouK3kY6CM0h3/ZvyViL6e7dFfCC5Z
TeIzaYRj7lMnchkIsUT9LQ/7A3vBJLeC0s1wSki3eGWXCrTglpph5QuTSkAlX166
Izleq/12o2haDgp99gBtAPS4gPQeWuuKso+xVvdMoH5LvrSeNhtHTOi4R9Ffr+sb
VEaXDLgHcqyxzkrFjqNRDy5927+CPXlXFE9AZ8G4NujquWHclVXVhjiAG/E/eHzk
ALiQTMfunQtC/50RMd2uuhroeIgIQU/SKrNvN4P9FrZJAHvHo9fkS28rjqssRO7S
f9+cuJmm0dlQ/DKzkwbK/sCvzUWsW4gzoXC5kssxX3efsTwvxt5Z45tvF98WfU/k
utxQ4ILyX254LVnlRA1+n3r6Mnu173O51KknnzEEotf+/v7wG71FKxuZ9DhMT5HX
KuF5h32LucA8KebSSP/VVBOZQRQez0kb+6r0dUhXUSs59opZXwbKcSbH+CcCSd5N
G1qfdB8BHSW8M0b1Lwbl1ot8uj0Y253244GJhdwy7PmBZtjo5vMPC5zG6aLIBJqB
Q9HlubIQ0Rg19ulCSZPtvUAEBgZiwzROd6O5bqhInp05nU+F3o99zQ3G4E51wosl
4u6OObV/0PcUxg0UfB5lbialbqrDNwCkodKYbbeH6hkanaPG2D1pMDUn/5vKUhKD
wOCS0Zug/YTTg35opX2frxPLJpYdjv/KpwwQxwEniavmrGEzJvSWuZRBqzSXX3pp
4zeyKiHUJbrzPCKj+MJPvBiAAOPaUaV9oej3/wXHAXAaL0T8VnucgvtszYW4lvRd
SmnJ1lLupPaRf9DiDOA2sbngW7tNkypxifXgcfNeA3aivkEp6mPdG1/o2/9+DPp8
3Iaui5D0IlLglBf83QRFVhA7gYKnj4F1s814ghlG0QRNP1UuMpFzcerpwpBRYH4A
aguakS3u/dCwfiAx5tx4fE9l+Jd6gwy8OoUuZRwH99PRlTDyDsL82IPz3fvOpXwP
oLDNYzpPg8Ibi4nmEkk6/GMxhaMGFasQM5ydYYwL7B6zCDkex2ffz1/bPj3/V/Kz
SMEGTl2gi7Oxlp9rT3VPHgW2og2ao4OFQ3aheUurhYq5X5gDd/Z370RRq0tY6Anq
W47fceU0gGLmGb/aW2lQD/wZQtUgLB/oAhQ4tFGhCkm6kCbfk7MURejWF15bVoVg
NJaIF2WYF6gJjm9xkBhSfGv5ZzShzLxkSyhVitvyrSZiiWC/rGf3Dxfxl/b8Szli
KOfKItEf0mFIbQm+cvQvMOOXvR3AnEV/tyrhL07JpYzRfNVrpEVZDPmyPnOBCy/V
IZfar9NgT53MUq6mmfp6SZWA7xJndYf1MxuQDEgUFyp+5sLkdUlJzAfAaRjb76Sv
brNPZMWoleFy/1NR68P5vuxyxltCCSgXzqneMo+5l85AKY6pLWH7yXR1RpTBrFPG
oxlgG08BYniLAzxiFaNyylmjLZkqCcXAqax2nLPIGM4WYUZdp9cjEjciuSeoxQOw
qEvJv8BWM1+i3KVQiO1d67HxHQEAPTRkKlRSd/A96XX+AhNO/3muU5N7a0RQ5wC8
5qwi/D7wVpU+e55OJPW7NNpYnNxS09qdV87LCZJW5QC0xvwhjHfsGcVb+iUdirfS
8QM13REi4lgX9Fk+LVg8JgPufpTv9WGZhKNfeltW4vGaduKaRTjM7H3aQ7GqR86a
RpskbRikYf/8JkuNR94S4h0NP4jazSBJ/jQj9aW56y9+vyZAXIF2UOK206GYsXPX
FfrYuIpw8CZq/7oKvpCcUtOf9Q348CJ7iHOLsabN9VNE0ydDTQB2dnM/8yqsVlK1
GuP9DIrgW6aIz9KZmwHqVRhHfP00t5E0vscLBvXvuOMxC4K3poxorOoIRXOzhg3b
j2D7UTumZ/s2W9OL9LpyPe5phxiz4QZ2mdYQziEZ4yd0nFvnh1NyKoLufBBIiNqb
fxFQBvBzP1cjmCXArWjAaJsFka3y/sB34X4E7xF6odeBkD0IuIu0ljngnYsjrUvn
clzzvh8nx7fs36r9vhqWgPISqka9h/q1FnluVJP9W/QMPaMemassPxp9FCaVjW1r
RQ2fZiY+4Ydm94FPlHAK5nmEn9aKNp8hlFq2PPqRgkAH6BLUopiDie5FYS13civE
/d+KoxbBLeQ0J53jEh9/p571eBbMB9YFTIaeKF5bIvvXjK0roaebsG+1DdzjxEON
f2i1DyyrCq2geYmDScBDWfjFNzUXoJJHAdIXQnvj4IrtMY+LrcUpbiI3h93893cN
uzVfJKcSoWcFk9TxT1RH1l/h4BPiBMPESgZ/uBBmPWRdXI6cNgVCmZaqGL94z9N7
cf5mtnC+iEqWMNjz3Io6Iz9CM+Hj7pwYNwlD0v3uSWMb3afakYa1YNFO1103wqPf
Nqg+mlTjExh+8lHq0vhh0SPelK0eJovINtpDzDK5GnSgWhGOp9+9yaop//kwvFny
jzjv1pNljbJiiIEhbcwAkQx45drg4ugJSntXSWIxkNdouZI8eGcSqRa7sJMF0cEV
sCTJhc4LfKyUNj5xdFQ9oWSCAztjK+pYrEyN4NRCaqwhrWJgdoAYyOQmUdm/tHVc
yJ6a8yLJr7hwd6F7JlCcJdE3hHou9TFCfIgcbEd7Mkq8RTUpbTEXIfk7Bq6iSY7G
645dEASBeu2FohO140NRZ3Q6kJ1cLpNJ3aeAxfMDNZzj1aTNuAkM+3jSG7LnikWf
UObIOeKbzM6Ro2LjGie66ZapD08lqxs7rsr190Zh4s8truWaae6ZDB34VOu83k38
vzB3dWfx32ALMGENiA6ikPfFi+mfvi6omitxoz859z2NMIwTNb+3Rr312V4E3hP6
fwnd47shl7iLG6ED+faQWxEtHrVRLbbaemgn7RszLdNogH2kBQ5hmLxQV/1TpTJC
vrh5cKatmQpvyKkEi5Xtf+2CV8hF7k1PCVmWDH8WUcS7rqk1IYnBgVCsehQXejd7
/NvtZdRhTZXxyV8FCxEwdF3A2+KngDOo5fsQTWHahVNRu7UKgFmBEEyzwj5HOfTS
FpHF7oTRakrTGInM/CQANQxkMe1RN7fCcRHR1DDqiwH1XTHVXG7wD8vsHnxwle9E
XmOa006St5nDdkIsXGLn63SyDMpANDRTqQG/M/AHCx68QNo0BNgEA954BM7gPiTM
r/SNmWoZcerxbdI1eMoqDwMGvyDCCOsJ2EevIaSoWeRRb2MBBSl92laTvyG/mTd5
deu/iOlsJnde7kYGUuF6NJ9x+dmHtj5w8rfhkR75J5cHCuskfxqysVOL6U2vsFHW
vPYk3Ab65qeQuAiCqomKeUAgkQNcIMA3g6GOO+IZyKLaMDJ38CmQm1oNNFZdqHDA
xQkWYrWjBArLfpB9H6CFyshBG1smJa0f8VxL71G2pWue0ANceP+i7z03Hb4OUs7n
y+SKBU67I//DPbZmEZZF1Z51t2XFlCTdUYKWn1l3VILZZQh69EdhXDILeDOZ3P9D
DB7IP2atEI5ZxtEHjlgD3ZiDy3sKiPF7N6Yy9RwlL9k+DzdW3VeEhjszXccJ3dyw
xtCy6GXVBIjaPDHZps7bPS0qqHRzg8XF/ESIThNXGNsThN7Nq76FF+T7G09EwrTt
HyHeWOWdlvd0jJySuK1z82j6oNTw9eu240vhT/ANUgQk3tqf4ok3730Y0IIhXbDL
3V9filtCdP5XYXAvDuDSOuV7mZMPO++aGYcli2ugx8SHc4s8BG5KIzixbIf/fECZ
1+N7CT8nuo7OC2oyvnaE4Pvy1dIW3PrZXp8uFiyTmPmg3dnTLhtsAgy3bQtRygjB
taJwPTXt7KfXtWPeZkZziaRia1PLu8qA8DqvT2pjEORtwu1aZxi3XMz+fLHiOcuA
znSI+1YQWcwUhcD0MwyQ/jhMw2iv7CvvYJ/jRJ+901cP3tdsVtQnE4PleOIMNeFZ
+cX4cv+oRCwRbPpLH/qTq4oQC/RJB6+igm/jlJk5JAyXNguMs0u1Ulu4OnUv7pDc
dY1/GNAB/RJNI4QdRVKm7p45Izdbibe45YwB1Lr+Cvi7+XbVRx8xqWfe8/JKIozn
oCbdUM3BKiQT0DWkz7vvO+0WfW0LH7OQI+yOPNw4OiF1C3P4I45BDOQKp00rTEni
8vd9YPgvh2MR2D4oyOWzwvZ5d/MWiRqy0JXAx38BcmhzTGPz/7sNEXS5BjzutbvN
Cl6XZZVSe8q1bYlE7ku/Nh7O1IMM0UIUxNR5zniBZeMI7gYKhyqeJnIv/5CCGNY4
5CfDL1D1vbz2lJJxUsg3cKV1joQhS0QvlYa1YHc1EK8cd34VMXvQgYsvZ0M7qrRV
6fQUiFAivl0550rO3QO1bmTpgyjap/eOZ89zG0oa99K6+Q/NFufMq2EfPfeTsMwY
oXc+yUISIS3ctMWoMFjg02orOpsUf4ZIiMpJ5UtQG3cw9ov/HUIVNOfr9ZOWZyed
l+frBy8EmaV4XoueY8RgtWeCebwwZCvXZbUWZ4dM50C0gCz5zj22+czfAZLeSBql
06SKNaz7RtST72Pdh9uhZ4P5UFtoO+sPeyqBYS+INFzyDGWfTc9F78QrPoJq6nvl
VHZJ8Hh7y7PJBWH7IVY+ry+QVX5HY2w02CChiRHzVgVhgWrxND+hX8JCkU9kzGCF
zVd+d5fwEbDA9hppWA03PiYn95z6t/eU4ZT7Vnme1bVPDTKDFv/ka+YeraPHLGWy
SUU8UhvC6HvU/dDfAogQHTQLZBjqhGOXO4Bim4LZuOKF99327KHErEof1fLh51a5
AmjHASO4XH+2BTvYHAD3Mv+QUCAbsx+qK27SYkWOd6CNsLbxawdYjRjTwOu95cgT
bu4aeYEM+WjeS84LBlepStnlAcKm+x5xsOU8H85p3971muKXxSxDNgITbyFBGpWx
TGPO9dp/8x+MY2/+8Laeg5imgjg4orEG+hGD4gMafRl9INw5fm0F7kqMUFTgxx8I
pfzKyxvJRf0w77nyrFZyxcSPH+CrKdymO4P0NmUhxHQv08B7FzJN32Cg+c5YjFtL
7K68HJyj3R9QKPfIMEczi7+0JL+Fr0sc5y+nmekgMlRLrTOs1N2OYkGaLzk7q0VO
eBabicaRGeCMlL20ZIFHTwzwvF34TKZrI+UBlwntvFIIsnA6q2WiCMCBw/8jC0Jl
4yrqbktQbYqFVuyYmnPFJvSJX1EbK9BuENkZtZRRIjKp7cLuzznqxgiaREZmymIS
wf2P9pPbI857Ss2aSusG9986nCEeHmQkLn7bdcMPBfXbyZFQv7vo+MMHNDprXva6
NUeAkxgP1JYshWqCsKnkl/ZvSFcUkAGEhLeOKyx0jUeSMShi4JXbs62w4aWfJBnJ
/6PJ4dgvtLW/H5AtGSDJMljqFVzvD+oWtbY8n3KGjAAML37mfuOkyYib0TEqOiLg
EuK4NpY5mgEzvYOnyUGlGsQwc73Noo+X5+tPoLCb+VHN7ibMs69F5U0/vbh0nAhg
qjA3LGeGpSlWUbby7dtzGQBV07v1zkLhsN01PAopzmvdFGPNj6nKub6Zbp9BsUt3
20teNjnOjG1wy6QsFV4GomL2EbyKBmmw/5wQUFyrghD79GXUYjwcineHEjiRlVUw
kh8Zk4Y1/H9rqqouWYbr8jn0/24Ics8JO6edt4inlE4/aozMLzodgoXJPcp+8nk6
ua0fQTStqvUGE4UYrnVcA/nKXFv134kGzXT+2hVmkVx2Z6bLG9ZtTCqvTeS4zCTL
OieH3W7ZZF9lTxv3sK+AxB4NZmBkd2XmlDTy3mEYkfIQ/FIEr2eq2Dig5vKdzqUt
64wEqsUgA+bbMbR6ZMQmIckG8TNjfsqDziTSMDHYetMLlWL6bB4mhMUiqzpyZqqg
xGCbBzDcaJAApsHs7SdcmWr9BV9y90E+iwMsTqKpsXaoeDSM34K7EYrLVaplX4FJ
9yqy/dc1wI0SP+WRiYyv0c9oIo0ippRHGTaJVfHXaGCgmztFwRaOCZzg2IYxZGyp
iN4nRciCaEZX2i+JCDEYffiir8iZ8i8Js4kx0oDGXdniQcDPnYulNab0HFviSrd5
6d2YsRnZl4mxazJbvl2qgWW2owiWXJH21XE1U8hTZnxcAFRWBNBY/fw9QDrGPR0v
XEmEpZBn3csP3kR50tCqdm+l3IoJzxwwCNyp43aM3y3JzNqQoqQCkMyJUPLXTmk4
QW4sCVgMVwBov8SHrthigzUehIr5TWybfZqHRdGCd8r8+PF/qaSyLxkHi9USEf8e
7ijVjAmSMMN2+/AZXGzl4Gdtl3d5WTqI5S6Sqg4kzZ8GHu6sCt8MtkP7Xd9L8M/I
DTDlfUerDjpa4F2u56ijskC6tgqZRYfRXegXpHTEJ2nOZj4/1PlLvzR0lhXhaf0y
Kw8tvEiZxNEq8ij486ePqKMTDCInCwx9l3vBIzdmMTDJI+9ZmrhR9tWvkcGLPLVt
4cev9Dh0eiSwgmaqX9AryLnssMEFOUOVL64CkZH6gvHJGfDGrn65m/+oSNMs6V67
Pj9a92r+yu6MivmNvlxsnvlTcbl/k7VHWAG6oKjzSq906Yh/IH3pf3ZR2aj0NDr3
cYSsyjFu+7v1rEMHKDvXid1ILwBLWztWTjkhpSWPObW7ZXzRB2Td+1rUZx3Kszrj
JMLQ+4lldB57oABCmVWJixCvitz+xopQilAOewAclsdlAYzVR7EGlZrARUzyofHx
FolMUyr7O3I/gPiJ4EzxT5SZc/M8S0EZzpX81LHgoPcGqME06DFKmx1w2tTPgCuB
FfTlPNxF0v7+3JZm0OSfDBsrmT0hfcNuCFcvmqx2pLyk9hBNbQOCRcBvvhj43ZVb
7LwobBPt/mgH65jLZtwuZBJgTWvHinVmB3+yOXrdZvPTMSapbuD6msiYdAub6A66
9XUO3NPPWgLaXXeLRfp00e/7QWRHwIBwuu+c9eFQjgQ480xqb3WCofV3U8aj5N+O
W+jpyihnsYoZXf1SPWZqWbpfzKA5lg0T4BDlFoz7LN8Dg7Fe/hVzw5gyGmdS1KDl
olMUo7TDtOoZA+ubKClo9/y93JMCcpa5BBNINVVvHZNJZsRlDAPsPtjzF85EV2Pi
IoDwSBglEZKDKQvY/rjAXLuhmVQNYIMxi4tF4yOIT9D2C1gqiK8Zd1IEE9Yu5Rgo
px17m9fzqVNI4uS/ACZlioslCyvi9dxyt/s30tzSApLo//L0MX1UnMaHuPGG8am+
kO15Sg9W7c/I6rsaskjybmOuZq7126ZV01Mt8dL/6mRVEUqaFeVV7swerDMyIT2G
U1ewqtKaNdmz8xJ8/lfe74ptRfvweJJz5jQ80LqvrpA982t2q9GRBb8G2MVncyjK
Zi8Bqmqx/sBYxLHYArBzUvr1o7OwC4I/GOVmWgjq0P9XBNYycHkfFPCwhpq7X7K1
rbfsgZOjc8h7VivhMzZ08PLGOdoLTJTQC2DeYSfGqQVProTS12hY+jwtkzp4G03j
v4X6KngQDkT22wxEt74yJU5Dmwc14TUX9uVxLXC9Xpqz/7KXTMEbTPlEp2DvSeL9
LUcxxJUkR0gRc0/7YVCd5t3vAx0ZoIFsLGsTtvUGcdB2/wwg3vZaPpt8UfxLy/43
ESVRUjPkOmV4dRa4H2InNQfhd5L8h7XGMtX6JGDXipNnym9G/n7c6MvIVTie/sZL
PKUukZFo/iDwWPu+Bycb7A13G4YooK2xiOqrRPDON7HC2u63dtqDLhy59pI8CKao
5Mf4BVL3J/IsYPBAA9vbbnNnNZd43SniAzSfPFhSDD3ctrGZqIxUvcCUf2UuqMNS
DGtNJkjGK7hF43wD7Nb7carOINw+0IQhrEgRNad23UTEVbtx0ZDqb7eyzL6sCDog
hyeBHQUYsVpYVE1euQLIZopBXo3Rd9aXG7l8nFJFqPFfnZWLnjG+z1A48g8yYHkF
4Vo0XODbjxQttS1E6AgXTaJOg0eiBVRxf0qYiNui+yJ3UpUWMyyYfwkPx3i8qMRl
JxU5VqvFZUbV30/cZEOiBihgMHIcz4Idf1Ll+4Q6SinLVBbeAbvzWTNAECFAbs+a
W1tHuEHUPnFRN/CwCvaQKUQ6SmwzrMXsb/F0xpCbxazeu8VEvuhGHkahQv6FqqRT
vB1LQ80RAMq6gkzjOGo0y9DofR+Ay4S50rL/zrx+umos6GOVQb3/FyDp5huKwRP+
QjmvU7JTXcUgDLACMrPbhXgar3bFSk/ZyGBtj/xvyOjyiuTdJIqKTEYcHDZqpKn2
6uYCYmi2QClrnfzoksMRbd5I+VYd1sCcgL7veepq7DdZdzaPFpTkYblfFYrbHTSw
1EvR4MBb0VRSdNRkfPlMy2/67ItNujNuWscOQziHL1P7mT8/O2zF9SmulN2RV/Kt
TmT+6phgbnCVcUUWcaKztkcac3wwZ5MmiJjT0IlUZ8OpYuPb++4L7JkzmpEsF/T7
izn1z2lEqJseJAPaaQ1VXXlUhR3yqk0AiJM0EFXFe5VWJhppuH4jNNp4zyElD8SF
/pxbAbb5vBIgEkPEzONbRLkSkpCrnOT51XESbP8Z7jkoN3lXBxdsc9V1fCdcXUYO
R6pEVpihPA0XAAlk/y2Xcz3uxtLzgQWe5mWIJU626pVnAY7ZKXoUViSYd/iXgXby
Ni+lviaR1skIRo+r+zVOyaodAhSDmbzdD/DmYPffgFFncflfyduqhv+GDcUoZzxs
Cp64mz/H8BVLjPKWsUK55tbxdv7i3B2GIn2AVY7DPX4ygGkr8UDTY+6t95soWgaX
EMYiG5EVmmshoD8FYaxn+83JtDvXB1c3TWKJ8GVucVCmchRnsJFtJdQqLml143gA
Z0Lf3Kzmob+iLWebvDCcaGxSAL0OXnaLFniIYz/7hHUNBqr++8xprjEFncpjfqQA
iLP7/b45rPy/LsarmCqwsiAH2/ClxUIxOwxwNXuRYhkanVfNrDyy00L5rDgJynlS
ruS+tfmflJdFsQbDUWIl6mlPfCIbtlatzh9FsjF/2tjyBInyBvjRt1Yor+AAaW3L
53Woxu7Dv4vQxn4nic50AqOwLaYLQTxeuheurmyUnSJam4flPcD6IZQqU2Qn3YZ6
UjEeTPDZvl/Fa5ww6Vzu5SxsU6MkuAbAUBC4fz83mS86+WLw5vNc+A2bNGCapfDA
W41kLsioP9PxX5Or8yAplsicIR3tC+2mr2/eI2Enho2w4EO7lwhQzUJ+Aou+1ami
g6uDB2NGEERG/GY2HU2xDQCcWoaSmtZBnk9soq2WGaIabpEkVxzSqcNG5PeAOp3G
IZQ5WBNDyrLwycXoLHi+fv0EM1jI3wu8bkZc8wXc9dROdcgXoB3ekTtAnieDMAaM
N0N+A41hKi2M1TiW0rFkpK3KInjOAV1vpUW/ReFUYhCW2XoZ+b4mYZU5uLwXfmdK
XGewjclozWWK+pzn7GXyrs7hNIki/FwuCuOH8n4sk0oEDlLLXTD3p9UntTgx0o1L
LrzktS26m4tzvk8xtsnjJ2FbiNUBAr7C89/9Mi/j5nM1RV527QOXzy43kQiPD3jW
5ogoLGvz3+5Iqz16XtWfhBZ2890tmXvB8LGf5FEvRCxLnzvAspj7vlaJdjrYr15e
fwZf/oRxg40calZCZwuofNxuFT/FQ7IfnTB23OBIgMN4OdroDidUtyMzwJjLynzF
HhSh8u/qB8DUskdF+/iZh/vLDQHg/wCk/feZ0b/kNWLBSJf/nA0zlG5GGz4loBtS
H4PwJbP3wdIfJOYHxktU3WYwBYN/pFa0/WKu3pXdSX1wjEAjJD+xSjT0P6nXbqFT
+GHGuv2KVbBXUKFkN7lmqgRJRLH5xWXNQMqaejtxC2z9B1ONmRAu+UuiQs1SG49l
UC5UFdRaKSjAKe8XRNH4HTBY23c7OHYN7sQI9QENEg3W1u2uQRX6gXqfiYRi14db
Cv9uSi46NKXjLIn/wmxxKLC5OxQG67HLg6go/r12Yki8Yi0rbNsNGLFdVPtDOjDq
KH/51G+GZhtLBHpsobitYe/4MmjaVHTnfjnmL90DiPtZZa6cjLLMx+c7vEAO33dp
yO01OvaI16gKZqHdZGfehy56YY8MnGW7L9Od6ccmBelY+eOByD+SynufX7SpMn77
gpn9VDzs99DvhpEDRKGglgvi8W4rK3lBDQFzEzzIFxn2lAuQiB0Y7Cmeczc4z/wj
bPQIne3VleaOifsQ+6bMuzrhhRQ+II5NVHqrYKPTxF52O0IoklOzIbnEypysTYpm
1OyUQawED2IePrGAUKUcfYULQSnd58FpR9WRddNSVHR2/nplXwySKoKAKlQP7rNt
6mWvdOCRaQStvsmsOlqXVxQkkT+r48b9jY4UkHF4R3YjWQpIg/37UdjTM976SDXy
HN3OkuVrdnfzM9/4Vu6d8TtJt3l4XCojTO4FCOLp6aVZlRSiyDbBF+FnQJHYIyM2
iKxdz5yIyyrQGyIpJQvPxM2VCA4mBi+ZMqqk+D2J6sITMe/5v9guoHePIhhAjQxI
QR2EzP6IuWGUP1rWvZ6XvvZghzFMvKG9sbF2VxwonYWLh+5LCjpIwHk+Twfq3W0i
7Rh2yMblCnpeKNCAILqPPqGnicB4XxVubk/RHE1dMtdJlz4dsug/S0vh7dc0Ulhe
FmWUTmwukrkNUsWEKq+cSLlUycTpN9ZbS/+QTRh2aX6dgE2GwGDzEPNj5Rs//ffA
w/qdv+TGRk7FN7n72FewxLpYqH4G280KQVJ1zi5z2EymYnGKxEEv2tO4AB6Fl3Xb
2o/W0M/iA6zddb03zf5twizXVoOlRqKniwXO3dpi2JQIEsfHBUYWvHUuHYfRUw1j
L/RgBSEnsLXe2kXM6UwmIDUwxzOT+F4TKSBi5I1DS8RCjpg3prVpjy9Nmzy+dJGI
sl7fDvsoaRt5mhWj3RASqdIp07WUQ9xj4WbPlm/ZlIUMP+4f/Qv45McEkfOYYjCE
t+tE3OCNgovFVa/Wdhny2WN7TmKB+IXps7+wt4admY4pdOKpaMEtFnei3rVLookP
qQcZFseiIexcSWi3wofoDA4vWXE9ZNVxh1Xvejo0wzUFYLQMrDxVZg4Cp4VczMN8
PhK+3cVsQpH47thPbvgYCKyPIY/gim4umxs+3oJJ1UK7ykZdel1DX2buvObL+5xi
inn4benqQyatz8zXWMVQcUO2I2lvTpigvKziJxvYt8tFInIySTJ1w7C3EV3hXUIK
YqQMbJuismOXS3M3aVBSxb0tMtDwUG5wZWrDl/WO8iAQqKDJ4xc/qbf/MMggYTzM
JhVU6/iZsdVeacHGw8BbdyE6sqwRmauXCQSBCU3wjoOPrk2lhpABn8VG2PKehCio
sI/aaAlbeuT6DhOhqiq1JNbUyDvYclMefWqgZ4UL7+hgWLP22vYJpngI7A2WzP3w
mRMTkmQMgVeXGs1isZ2oppxkgQ3WGTrQpK38Kf3uFWNfDuHFCDu48aeQs5OjIqtm
Ns3Kvmul01L/I00JD4mDuroaDnGy6jSpPgVq+fCmJtP55PyGgjIoWOdvcJE1SswO
gXBLD7UxKHvrz4EaTfPFsGEXzeWzKC86bYN7U9ZyGQQ6i7iUOgPFQK5uVGGH5KPY
DnlsCV9q3UdQV5xBfwjTQnBMBFDKuVvcE9s5f7AsbuDrRwkS6o20zAQJOX31MLrp
8pyWMCtloakQhYlHlKlMPKGseJnAelxVJ/bPgGad8VCZC8ppu6vKHwvoQwChDKCN
/8eoQxBkTdf2eLYLxiBDGMKWy1QTtWpc8LGPNvCdBo47ZRCj1WYKYURk5Ual9pVT
wpQavmGTqV7NVlWLQjIQfU8gk40HRD+tEMyPwIPzliJfzkinkDkROIlwSUGDXzLd
ju25hmkMJmFkVcu/L5K8YsT1n7pDR5DV5dsvgqeDc4hiOB1xnRU9cAUkdr5uyW/0
jkcrDY9Z1xTvYNaZk5nOT+ZwUpH5Cf5k9cFQCfUTZ8TjGq4rzGV5+UIa+34Kq4Y5
gC8mO5DQlpTs882MtgD7sO6g8yEkUrjF0VjVPIpaNqX+L5Oa3+WzP3/TbeW9drrb
qPND10ICFznGa+nsZhlJseVNULZfCb2kP2fYD2VCJXIZL1TSyHM0kWfFyvfw/Ppl
O6RYXQoz3w23NM3omgi97qyo5o2pHcOm809JgVVC/LV8P6ERrrcygQma9CUYQCQS
iFBcNU9lZk9r8ztg8oVnWPZ9+TOkwrTPbrcnh0iShEOkcG4uXGFhFiCzG74k+Za9
TUqmtMaw2evI4bqpPZF3nbMM6vRJmtT88Zskt+X7hw+iY6sZrng11RypW8V/gTkC
9RMRnEA2PYVFEAZIqqI8qQcXQQNb1wlscOuNhTEREStaBekDrgvXY+AadRJ4qXDA
/FkKwCt0dTrziTxxaqJwBOJP44mE0bG1EiVwWSo4dbILUqlP9NjjDWruaghF1oLa
4Kmu33Sop+UPgV0YuKP7T6F2VpKkuEJYUdCUoyAv4r8KON/wtbB20osQuEvuM2aH
I9IzkRMtMNWFss1nexhGOG8messLAORQ1bKOq51Ddycge5oBwgaTaQCIi8i110iX
zn7T32JJv2OeFcNRaX+FDSiI1eHaEnZCL78220JvZXFkwvIPBTPnFkCpxRR2dLA5
Y21ORUap+WIua/CnkMKz7Na79OiS7F2Q1aYOg8RYD/V91QrPzFX+D2Z6zH1OiayN
LAE53WOhdCDLd+UdzV6ouM7qV6alplVT7fpDBGtL9XE0dOk2UhAlAcitpDBGTuUW
eAKNvcArCvAMbmxXG+csZYXRAK/DwIQmHP2BmZJILBcK8A5JZZG8e6umhko1j2/h
g4gjdAjW9QUJyTUvuq+AChKUeDkmO15G/o067f7h2M1J5igNfsS40RwEQSRgWOCf
9vx4AKJEtxdSKDSAgcxG05qxJgpEUecihAyFq6HSCw4rK/J8UwiwrTRQ3oU+HmYJ
HXCx0XtVtv80g/33jygXoAcUfljLeHctrO0M/YfXuoVdmngQKeYQkwI37zg0eZKj
Dj7ubhYoqurK2vdLFBZlwyD8SQjX5I55CV4iFHcM8SI0y0L5mtltHXOSbAY5+NrE
VerX9TaemncYOHkiWB4I8L8x36UYNBr+/BENdWYDLMAQrdm31peJED2kFU6w/JUZ
djUQAR3Vqbq0qydsrgo/3/ek0GZTLTNYPm2UW32V1CIbtC4ImkvDPKfqYZjkJSwx
tsgIVxq+druMsrJvTlqRQ/WoTj+qVG6M1hTSlmLMF7bDtonpxzVeRHxez6/j4vP4
JrKErcSFIFtrgd3epsvSVGfVhxibMxT2rJ8prBXK/4loTkAEsy0xUbCt7Q5arJVn
ks2cBWXjDG/HB6HWcw09hoL1ECk0s/+LfY6TpWZGHE7jziaQ3fYkT/sQl4Pdwiwq
A8avo6ih8nYntyGDH4UzQfhZy1VXR/2SJoW3xSvqHsFaIGP/itmh7tNGvE4evb9f
dg+eRyb1MSWQLGfWCBRzvMMLngFly09+NxysI7KHyoFC+HLhW8mRJonC2g9hXPj2
IIpCCj0EWBQN62nxZj24RU/KEH/GGIw8mwbLNbK53/9PgCZRMb48sOwqcOLLp9TX
jj8C44jSEhFP3Rlq0oF6LIEbaJUx90HWlrfK1kp6Kj9yeoyJhyLWtF1ZJtOB/xEq
mmyRAFoFDr1LaF1kE+0dkM2zC/UaySF5G2X09UOn/VuzN4/5+ve68YZijhzfZtaI
g87SAkv3YOdMhrJK3WST5KHwniiHq24naiUkRmR72VbXb/OISGyAA6CrDJCkO9G3
aZhaO3db55zscs/9sNBkTivo8hgov27zYBlPbmuRhfCk6au14AYiahIbO9/6+BpO
mDwvhTr7+u+JzAu0AOVxZFesXEBSm2puKGVIOfQdrKms3NbSqOYq717a+aKYiS06
zEwasulq8qTE7a3jBd0PADXsr2KHhH5c1fizn/3397syRjI4zWkibHCUhgvrtfss
U1OVrj4sT6oTnwFIn/wO1YQMGhEQ0HoTdyL0lym7newJkncPKxUEXrKFKQEXXIOL
qWr7X+hG7Rlf48HNHzj3aoozlg1BI0gIDOVEODsaddd8f872NnucXf8q6uGtwAxo
NlTaxQO3ptg45913PzaIeGsajjA1jOXfTXwhro49wq2GMflnhf/+BWKMnNdz5t7Z
cgs3d/xGnra1oXygfLSSoaVgKey/F3pJGocKzcEW3IJuj07Ujyzf231PkYlzsWsQ
bw134YQRUFwIQtgSMFb/a5wgbGWfgJxhsaOlliOFKkBCZwgRScI7DggWezm9AX4t
HpABjQ1QodY11s7nk29ysPP0fZO9AHRhbrJBhDnZJtttHmv+yRDLN6l4T/MQUIKt
m5MdEu47PUxbd8rpXTqTAJ0VugMEi+pxSRPODPXy9LoWhU9gEvXDxCri4eZE3e7L
SxgzkQiXi2RWP7eNjPKgzfRpeE7VbSBWEcV86GKLIznL1mIHPNT7F7G09fA/BzA+
H8Wky/oEnrlXbpF1lfGS37WMDjB3B/Ndv4iaLy+Re2ZmI+PAZBWPyjRhBOWMruTP
9M3qKRW26ERiCXDlbGvrcCg9WU7QMiaRpKVnsawWeFNeAq09aTy4P7eJZVDWYz5K
ad1u1QfsFEb960ENPnJydRgpSsvtVTJQOm5GExYa3wUy1c7umlIG/I7ipgGpi7Pj
Wz8s/wzlDh8xYN2nOaNI7Jy7bZmT3RZEuQWyTKl+MQZtREmpATgL/O2o5utEjpoK
7CTQj8pIgsfhC8WD3sNVO+yZFTkkxAit/2Ra+Zyu8y0WZL12IeNhDvFvAtwDBi4z
t6PcPIKDCz09/ycbvsVjij3/wQUoU/Up8YXZsD+ozjq5ltqrWHE43hgL0y4hv41g
EGrH15Z6MDzLbyYj5Kadt4iR7yAy581kZZoY3JsM2yxGD7+l7fbn8FwwkHqTbiJg
Zleyi9Sd5yPQHZO76s9UXcQ7kMiEUUq4yE+imTTShk3TFko3b+Ygw4uSfgtU34dQ
3As0nYp8jscMW9q8fuHfRbDRATRBXXRK3hWfZP4OIjipSHtX/mpoFzG8JgAuDM2H
KgAkBTwWNAAQlVgL3SW7E8UT1jQtXDhNyD5X6JEIM4h6Ot4QFi4T+RY6p07kkfPW
9AVbqfQU9oN8EldhFt2cu1ahJYM/Rz+U2qkf5JJcxw7tEggIPRtu9gMEp2UqD5EA
ryoK9F87VUqEPXQkCEU8mZqiOBCd8RJ+yKeDA86/uQOhADZ5vQ01V2lmyW/SvIvg
UF55BQGgU3Qday5I90plXg1q9MmMNTBsG6a1DbQ79DX8QZW9DpG16YctePLUvEzN
IrrYT8KMNwreAgkOLtFHCzCJdg+bdKjO0n1+IFuEEPagezz1i2Vw4KsDVygWlwO8
Vs8NIvqcc0fw9z6lfy+S5iNn+IIkU4aJULT6wP0DOHOwwxhdQgmv/XyzOp/8evxv
DLXjfAoSN5IkOlxOqa+ZY6+W8IAWR6QszbrkIhjlVBAIEItTWUoXV6DP/Wu6mdDx
GXlUoAnNenlZWTUo8QG+rsIzWhUrIc9dY1D20tNAgKLVNi6HUckwJfJ22TfSQ56P
V3X+oK/fWzJbBYfV9zG8jiFUbhRPefaBXYi1w0tTUeKK4LgXHez0qFdZcfzgiLJC
87bqUuvpPyX7tb1ZpHiXhxochV4LWmtWZhsVi0rjtvfsTR6dTTlm+On/psbHvjsp
qg94Zv8NX7fy8d8rdy0KiQdXxstSYWRiC94LUvEj/skwTOUpqWuapC3HbyoC2OIR
rDCUYySqHJfIiKu0wQsNSi3XSkEMucjTTIBJj7+RWsob8oFW18JTf7ty1wA8WIBs
XwdLs7dIY3wpg1wDHG4A7hyQkJMAblolPxPkPmVSkWDBTHQkTodmRlKquXimL4rC
Y+BhVNoy86Kt2akDcvPQ4+tIosJVOkQGIg+FI15miYqud0vQsagVyBca+yDBof0V
6qdGMtvstHsVm0XaY0L/hdpqi67a7Lst68jnN0eHKVSwshUpQrbaWzXHkfyMJ1Ne
P8tmYvUMiM5kK15ow6ppKGx0NG0Cqc44wYmmGXkXWGVBtcjs5uO0XL85hZnfjgHP
8gKS9DJNxEJflYoaMoqYvEW5KbOFexOZGSEsy+Kw7FoxMMPlJkTfpwqn+b7/18v9
5pw14Y+Wg8LnESfttIjpf4ML0D/01P1CUuHwnG7OLO4H1IsSu2zrEsCZgcnXraD6
4G00XuiGFs6Br5icllJHIx5eIkO1gIHBT8BaTisq/0qTuyFnzcVIG5exVEFdc0dh
NkcKt7mqtaB606ezQx/CybV5bvv76WWPOmSvZYLAbU/8lqNvNTLVGKClLfR4LBWK
LAsME2hby7AXp7s4UIOpylkSQ6Fx2saWbCGZ7EBw+O5NboKreCDFLDDlsJVBmJkZ
FvZfsdEXe+jykxwq3vA6PVQaTuM0eEdGnJc6qx+cxVIWFM8aQKmxq3xLtvkYqQBB
txmL46Pr6opZDnI9HYCDSoZwoWXPmwru1fbVIHXZjLhHVRnwrbKGRhDYo8N/uq/e
CD+43SbPJDd2DpomBFg5dROIiyicrAjlTeZtjpKLQejlMWEJE5NZU09Y2fZBaJuD
9xa6o75oLCcX7Wbkgxq5/jqAXUh5NWK5PuZEx1C25LUYU6RDmKT+pMI+mAv634Kt
TXESlu03VydoAfR/eB+/mJhZ4R0rY/k6Kg0m0YHYLaVOjWte2obetSRTQ7kmipHy
mjyXlipMKZsMT4qKacuYo1C7DQOlyne2NwyOas60ma/xGzbsi54DQDjLCX8UWF70
2zh2YU+T5kFJaWTNT0LR/kv3hqN7crHhVKJnJB+PFTDZnerbnYTA9rAzTnpEeeuj
WENIeM+6MphnONrxtvaId7/Y5DtJ/ITgmaiTpYdYwwh0T0IzGVsvhFQ0MrPZZnd8
aWhQ65oMrR0bUjwDRzwsN5g6LNQgeTkKi7NzS17DKBG2XuAIcWpD2hH/d6/Ikn4r
cixZI1AKExmacKQUsy0MlXpPgkkawnVvW7dm8efEHmhX8+VjzCj9NpaJ6rFzKFYR
yE7nJnJOUYZP/n9LMp4zM7pjmo0KF/+k+RahhZV6EY0IPM8ESns1vAZj1WHvAr8W
JjuTjcFY8XICK9qrAC8qcc+vW7BVeweR2CWkWncF9uRbF5SHgKRHbrmJmbRwY8BL
k9TbGFYqmlOGA3IUTPxQiVVMC9RgnQaNopkXRtyS2SiFWBWWT7QJrcFQ/AYKRcEx
BI5QiTJNkk2JCLxOzOtb2CmWAKo2SIu/zdk0bhGKSkqFY0Lb+E28cuwf2hDICiov
qoYVzz+mTwmV89PaXjNZ/ZQdra+O/nLoEZBh5j8LdaNFHAv+0ufnMCkKDYfhZJoJ
YqwZColi40nZ7l4btRwLjAwX/iMlj5G3vexWBeJnlq4gwv7qJz17E5Y/Lt83+KH8
8cCfSgQSFFR743C23Lb3pA68RuC0rslVhQneNkw7SLneC0oiMvdy3pq47fz9qYcj
0x5qmYM10Nkp+iROIE1bIDxUHjScb4l8HjXnDO7syAu/JrPglSF/DGt9817Oe4wL
RNeYwt9j3WcWLmu9nXdm5d1EmAmefrUYtBrbQa0dB0VE85Y8rCbBCJRLA3OivkHn
Jyz/KlkFlNEvdMB7TkKW968tMxMaLT2Mp1joyqDi1YjIDDixCUpaDEIEbqMYZMSx
a5axlwAdQIv17udMQOWon4zHZ946y3DlVQai3mheQjhs8cg9zS++jr51e0FKuC/I
zrAwv3+z9eeh7GRiEd0+v/aJ36XaO98MWiiAek0P1z7F4Nf5A3Mk8tIV7F4DpHVB
dW67FGomyHcy6T8LV/R6a34gAGz/BIKSba2Am1nurlwfH6cj1Yvs3+DTumSSffFE
mmodWfd0EZBjlt6SLhvnAQhDFc6S4ePDAuar8KSoWappD19rT5zEgMKKoqRat9aB
WNPzq2yqAZZNA25NL5rtPk5TTlFRSLE2pu+T224AjdedsiCSGcgzLLhRTXny6yqL
Rgrq37BUtBwjNRtLs7IMSfUHklGdpIemqjmXYOR85t6gQRLawaVH0AZnMuW90TTP
ekFMACclpk0+IiB5dLBlnUe6SOmAmj6KxJ9C1CbElK19wsTDCoo+X080s/duSvAG
RdGbMgKO71MnMjHvZtYhsQPYrl6witlAjeifm/J28cvr/uA3mSJyLAor677EFtxG
5J/jx+1DEuwmAhivqh4ZXMBeM4QfSLOAqdQyEkm+TZbANckxrsYI4Nwfdp+7hudd
79g8fkxhwqj4bqlldT9nZ7sYBAay2245Z4CbF1MI3Z3Gl9wVkKgPWbCTELXa9tTn
XDSPQB3DGG8K5ErocGGUoZGve2qw8lrCMxX2ZsZNpOK2UtYGeBJFtLRMLtTC9Ak1
gFkLLYfnJ6bJ7JUjcihEJX1O0ElQdyY7cEHuJssiw1pjbMS4RB52b+CSUIyoHrFw
BRc9jZL4CeVzR10uV8HyiRCtsVzcq2fPGD9h76pZ4fcY4drenbzGzJvF+pQz5fJZ
13N/qiUNQbn1B0l6jMfAxX/zzaHPBK5UowDWy7NeVf8rdXq3mg6h2DT5DScDx0A/
mfxRK3zpyM/q76vWoi3z3d3RkCikb2fE/N2COP3heWtDZBzEWOhu7qh3M3lJE+k/
/CI+ClXTCikwjdgfRTOCIDWZ8qeT01RayqNuteApQ0HDUsl+rzo49Hg3fcX9GxVw
vj+TkFmwsP7dzSjhPmN6/QK04nW81/ERktWGdFk0w1eOwJlRJndeSd4esWKh9wbB
XVdxfUcrxB2hNTYOHlnJXRzaFy6wChGasVdkh+b7WpYR1ktr4wD/zkrGBVrwYACW
UGgoge+fxfhJyndyDjk1oXXVg1Mu8msETvJrtTXCjX7DdNIwTBSa5qGwQfdf1KGd
Y50EXRQ2pQCqycyx+3XsacJXUga33k4k5v0clpucRgx8olBTDrX1EsU/Z6SEDfCk
bPKUM8HrGlInkh3sC6Ad8EG6DNke46zQlk5390Fnw53rROOL2dJ2tVrjtPNFNDip
MtnxNHkZOyzUex2BaDjr7LyBRWEEg7Wi8tEfoL5L1VNFcKZbuzj33G2TWpQyJ3VT
6JSCNWeNJz0zjr+VeJ4Y8wtsd2y90Jd4J8meWvpIdLNi75oMCo4+bpwGK8pNV8L2
u705DBNROqraNOos6WLnFwiRnK4QAOKyFiI1tiePRiiC+Rw2m+FgOOxTWxx3xXFv
VYuALhA5UNSyhaGWGkgTeE5UfJPAntzzET6oUPRUKxeL6oOwLsaMaukO/oCfHrRw
4yefPkn4Ciq+7Fu1/HpC5BHyAUCy8qKuqlpQ8LpFYbZ9Bm6y5msaV74Q5ALUiKG6
oQV6iksSXXhAyf0JIAJ2AswzSR71DcGK8884kuaXSOCwPZ0boVHeuj3TQ8a/daWZ
hNz1L7EtRN6H7R9faOu+pL8qhNHM7I0R8E2xDQdbr88AFys6WoF/8g0Yhni2PfPv
zFC25rD08mXFaP1xNewKoe6M98L5sgH7TwozO2P/JDfVg8Grxa0h9saKz097iQbb
wfXFcQTVpKqXNkenZpMncl2+VjkouJymsKIYIecBZ6GaIYl/wk5RbVQ1gbp0oisP
/3Wytb9T/IWKZnobggeiHJGOqtk9GPSJK5Gj6kUFog1mww2WO1EJBlkp5iYCDiLB
2lsgiyh+ENabvHAj+DTIAY/K3xPZXhcP8cYHkNtbfvp278Baxs48RJ20fe5wtTd0
tKh0EQAB717dw8PoeVE45UYJWntFQ7cu64irEEYj1efvXryBNhnf+8JB0jBC6vSi
u7hCXJoLgP6cGaOZ97aTgS9MKxT60izy0uTqfGxFG6ZeYhyCOz9TzTpvE4EWvuNm
04+9BAuweAB0lUWgrwf8q7tFM8O+jCsyVvGNtAhORbOSFvLn2zTHVM+SQ7Pb1C4G
Al9+j4GvmUFSTryWXsn290s7WthLAxE7JOJRbxwfkWax6phKJ7sBjhbVUcpGQE9B
sBLUXUAhRBggLNn8xL32Rcfw2Ffi+Xt8t5zHK1QjvUhSuRkm6mCdLidozuL2HkrM
aGHdU14Z19ka0G5HK9zYpxqpI/PyQy161b3JbtJjErk/WIbdClgShD9t7ESJLVQu
JPGu2qFL6ecuAOLir4C1FM4YmuFiqh7/SnJt1uo1+LQPugtXUyHqSmX+MtabQuvr
FIGuUMbSkPbg9Oc9pFRy/l/bidpXQu4yql5fwA8aAMZnvwOsFJpffbfNh+PbPexD
F/WTrqKqkztbxMnY+vvrsE/ZgJZ/vwrmPpO9tBdq6kLeU+OlfGh5PDmbeJ8hp2Ty
cUSubqBc4YB2DfE7SDC8ReTptQPtnwJlMYpoZntQ5OKZGu7DcjrfgXYQaHuqeBgA
3I+4zBLiWmTScHlRUCSVV4BLhCRo+YYARiLgVFKIBsCUHkml7zw+Zk95QCTwekjB
/lkOdYW179wJbICBRbvkF2aeiQIB0Cl3fG3vzWGlcbrDRPl8ImV/Wg0UFmJ4s6jM
Hhx31wjjL6DYQbo1cG7VoEuJ1yN2yDuArAZv/xXT+b7/uW5xa25nnNOGBjymjdmm
r6LTBZMCZkIHzsk6yeqYNQ8HJZhaYJM9cCo+8WOczEkTku80k/lsf5K3EnROTXYH
duBQWpX/S9xA9M61gKOEuV90qfp28WFeEHaLV9D2vEmnelab+pdlcQ2UmwOYiCWd
8jhnEeey8mUZvCULXtJTBTnj/02bU6S3lN9byR3e1cqTjQULbLol5ouwOFN71d5D
m9wjGbp/TZw6mNm3iakmpsCHhyITodqZ+ojTioUOfisXlO4jm4xxy4v8V9hoIRSj
FpbyBRsuapFyMHg+hU7m8grdLHfEzXfpk5rvbNp9tscWcyfqqgoy+rQ+uqB73vma
fyhuL1zOA4VUGIXA8guBOcu1u+WO+ng+zB1CPIt+qjYOI9yvwEK4S5KPMEPbjL+Y
rnbINEYld49WiIXe9XcGLaXnI/dOuQGG0f3kfSysp+Gnyq1Hpjj/QiNmvL4v8FHd
CcBLOThTdvj2gymuoL2uDPxSH8YDd1cuHZ9pWQgJVczy4ummGWrCmdjbndznl92S
YBlPaEP10E8CKz1BSBeP2goGwPWal8U7vD3jUQsSBqXjIB+xb6gV1rmVzipJ1AFh
v9ZUswamOhS/e/z6WKpT6nWVr9ltwI/4GlcjPqE0iJJ/ZOpu1+cW21bqOYCfgLtG
HeXcTMNFn2R2X1ExuDknwuJiQ9SI1I0JuRzjxopE+ZiRS/jItHVQP4jjyJKsdxp5
Qc32pooa5WaXWYR7UZglwQ2ibS+ZICs3eyAVEKtsbgoX455cW8k7PnpwIsE6h5w3
0qAGNqBlPcqrt+AllQpVO7s/Xc2tKDSBvfOxT3gAf/lwfUfZCULepl8c1/CY4s2o
8rhHzjh299GWLQ2UzB9/bz8+H2TMh7Bw0Q6JT1URb0JpHPniVdnB5O51gCHXmXYh
jxQm2+TFRkccGYemtuTvI8QUDXrL2YG1Zh1b7+8mQDCWuxYlC5/UmcrOXHTAvLLj
a+W+N4gu2IPeVfbf2virLYowKd3PUWMkLC4KwT8Nw2QkFsHT1cErTjQB5dgxT24m
/NWE7s5q84mZXAEi7cdT/oeiJTt9U+S268a0LXIZWnEQITdc2P3XnWmf0Nzh5LTg
1UNUhqKZ/utlSCNJyw4kbgcJxy6R6TwJ9M5Tmw4CEkfZgJYxVyOtit1PQaZr7yvd
Dx0+KSg2h/Amg506DrM8QNZU/qegfh7IFi/MFpFBz3uyY0NVbu+z0mdS+dnc9xJE
IkCbYKi5zMR35XY10LYhq3+ZECLx9FrmjIqnylleqwczd09uxZGgjSFfml24bT93
U4KuThEIjw2Q/G/inL60M38Y2LSmH6eLYShXF18WeQtTH8rVCpEJ4smxlZtcRPge
T/3LLvzid/c0efsJTW0e/lzc3VpQr7Q4uk2AFbcJGlWY/JCdzuhS6Pp9U5MbLJCN
ZTfFJHIMa+JxIKfPe3tgk/3E2bUbQEsTnMPbT69VKsdzU0ootV49cow6EzED1OJp
5KXgHp8AaunysQYGWE2nOg3pLFOMfLyXC3OALSgtVtvlf5xAQwnNqJ+jTs/RzqtC
Rzb2PB1eRtkL8MRA1LsEH3UykHlSdoEQyGsphd5MAXJVJxO+OYZpU36iz9kkgBsf
vrz0tJXysuC1Zyia1S+emNTe7tnsYDPtxo3jtel5mOQs02J5Xrog4fPSK94nmifl
n/L7ncGQ1+gUVFxKRoK9H+bcuCovdBWY2FsWtjWUcbamf8EQAX8JQdAErn588BIz
SOcw4LPlLUmCBQD9jzuyvGTgvmj1D2cNVlwg4RL/x8C0+/+gSku4mdsxRqEhN0kS
GyCUyoQdN7krwTDxHRPa6fmwR5pn/yiY+h9qOt0BtIFjtFmRw81ZSUPgw3g7R+Jy
jZGQBsxlIjOfIRAxwkjwz9f0bc8ETQj5U9hoJcbHvPRHOTXakfsfxcN1+I9fUqoV
v2A8TOUkrovl1zjg6+nNNmh/ZEhCbRNawlLCrqldafihyt+ypZ1KOkKzUdpvJIYF
OWLeYaU4ln1l2/Lhs5sLL6zUNXacIt19LKbeAQTfd+WoQq8bpjGgg3Y6HKcjZEIV
HR1G9nykdn7r/tsYpkypFdbTgmh6Cun/hFULaO+J7WQ/YRmp24pywbidCrB/gC+/
hky1J6jnVL4/YMamHfGwc7RmtvrTKlUUAebgZIGY2Pycq0HbdKs8EwWA29/iqpeI
jQJUYQGl5BNsCS/6EtmEkeEVletI6rYA/bDSc5aAacGVMOFD1Qoky3jVY0ieS5sP
K9xexfJsP3uks88ohSkXjrz0kdxSuLg/VGO16PpnKqbVDcDVhT3EEa/r3XtOHiQJ
Gg2wFKlSV23yQP5F2PVfg14FJOvjWmPrYqQh8cJ38mTENotkXYfxK1HqN7L3U/EC
egFXC227tNwe2E10qJ3QCXiYPSe6sMMZ4LLgS1IOcAORIt8O1QegPsRq9x4pDEIX
Wx1fOKajQBKQ0rgaTvzXvdt0WtQUtNb/mLdO/M2xtD90npdAWpOiELdDltrbdkZF
hgWMllpIr0F6kl0ubQoWN/Vx1koBM1Neu7dDkAyDJlTQVDszTUZx78gFZKpg1ZQe
bYoycAOUfDOV1nKPcSi1gcp9GrUE6uY5dpcwudbcIyQYomfDlPPj3zlUkLfYMRa6
LoPsPkNSTBWkZUZNYbTdhl8c3fZvSBA4SEzBBOeeAncBva2CW5k8XS9W6X4ST/ZQ
2ooDtHUKpmEzFKjKkMrvwiWuQH6CnDDjWCtt4vLNPneQzeshHGw1VEzdd8U9eUKV
kgFv4z/oEeIXp91+3J6LBkitPWUCQf4AgDOD1av6W3FnRjW/yV+gGTjVhg65KN25
Pv5z3d/88TBhBBR9AuvBIVv+HLlF9Wk7S3jlOiGlW2Kz5MesXAQZ8ihKFrtfuLvC
epfnXiqBK0Ji9IxGPrmkxqz/sYq+efEEgHr/rICEzEkw6h0ZvlTnOTOKJ+UZFLD4
i1NgQ1ixYSnxrq11LHfrgq3TbeL0zwnbX/x3qQNQvHVqIZhlTVqIXLcesZiZU3DE
BeL9aEGploUEnWPWUap9r8h5/FkRuZ2xSrbhY+l0p1GIjgAJoE/HqUQfu4yFyKI/
qS8Twb1oEW/i/EZbyUlHtZKDZDGseXt47zLW1yihxIE89QT3h+Cm3kEoUP39q6Vy
/c8rcI51YoqQHYgHUfK7eNESWxuu3aN38wf1E4PCZeJCgjoVuq6tAhdQO6M32BgP
QrxDr4IwenwxUfqnpfn43KSbCtmglDYIlQTGEtfvCSIX6seMu3t1OEK1G+bgF9HK
h5JjVHocGbKwgAyGz5lHIiAwZPCuPvAqL2X29zFdvnn619hb2Z/s8z3yjBGvRYmh
3plVC8o1MuqpIhgFVPy3nVtUEpR4qpfriqa4On2H4d2TWWBX8JnsYw67QKWmOpB0
HxedbwB6wf4JQmZxclbbPQFsjKEPjQCQLTB7FJUfWULe6TKOvoVZMonMVqPbfB48
ayNyupxHmKSjlhtrk5rzEyHgZ62AqwqFoRXgmowU8k8QaTpQKh/L6ajjbvmwNvWX
6LYuQyAQKiVLPDWB/pjmzKJ5TcDuKJaDSGtemP3XL6BfFY6VJRr52PDmviIU7fDM
yU3sOExyzVOVfpwUqI1Z9+oMHwMW8tSX8FUSbX9JuL8lQTYkdjBvZn3vOKc2IhJD
SUc/w9Jo2Ik5Y+M/G/BpXf9rTvtjfqsrUy0oetSmppI/cElv3YFFNy/ooWms8VlK
tzL2QdG+iTcv2YT431wGz4kPSU3Iy4h1UsnFLCnVFHHz28rtEoeuZC4wDCqrdw9r
JdavKGWiho9aak8VUT18BOQHWP5qRDmmpggb+ILSGuG/OExZYBLluRjW4RV8D2mI
VvCri78/2lF0ePVOcDhFkr9DV+5zJnr89kR7o+xLhhZXp04uXEb9IL2G+ZXxiyEV
9MtDQhexZ547O5EVKWsOFrlO71cNZfgYD7O05XYQwlVvXSBmoVgolCbbPrDfd8E0
zEsgwW2ppwRPDHFxACMJZR9Wxn+gApESMlGQAqeLTbEgfn6s13yNp+uBNUhANVa8
X9b1fKMBqP2c3VDLWuufseauzii5MzI8AEX8CZqLfo90iJRPrhfTP+Jd3epmGg/j
vG4wcLcO+02pV1xUdFuuzfG3eLF606OeFdn3SRkXJC1AmSYSh7M63VA2mQ6ldqZ8
82ulBJ4jETneyKarBvaMguyQWjrnmI1/QnM83rElAFMZOhY/ek/u5aEi/j2cTTs4
SjutU7YfHRr2AM4JeIbHIiLYkyYKzq7/EPLx0Lt1PBexQ9TtNv+9VtOSOCPJewB1
BarCgxn2czDG/5Xqq2Ld/uGARokhqnXx+rJlBQcqAomAPxLRcPSWMEMKQS50Qmd2
4pDkKmeqpWHYQVXkeSspTsagKLHXaJbHhoQhuxzvpA1WoW7qomM+dpQDTQ3Q1oo6
xGNjjxo/HiHp4awjHFMSJkA2HOy+CXI1BeOPAEzB4JWo/J4GkTKkkcMhdP1uC8hQ
GYAKdXQX1gp/CzGIEtWLaqNP92Mh4jUfsK8igWa3g4ESh6hufcJUnkmXwe5klePL
vYqnRPJu9KNOQu4QB4NK48BZ+mU3oWUQL8Uj/4gUWQJupP+xWExpvKPUTaQpuSQB
JW3y1MQE3o3ADcC9kJUtn4aY702iG5pSRkAI3USX/fDDxi2ml83WcoDy18eg/6XI
/JTCe841/UFCBPw45UOoKf6umk0ExSjUoBndZy002jSgQFDEbmF43I41fMFhYaOZ
4DVDkJH5pQhPtT3N3pJjA4JehGTP7cS9P+8ap96LUwBTCX6ufDvS6R5WnDVrs/1u
eFTAobBXMtsNGxYdoi+NqGBSr7kdsMtlcnMa5XwEMxRUwN8j0gB7YW58j4Rrd4Oh
4KTWRYMOJt7tCo0rvQRBy0wRTVcDxmO4o40nPzJZN/kp9/bnjSzZkWxXmPtBtEn9
Y42+G/yw4ekocbzl0GvZ0rXvIVpv8sy8/JIP3KpYeHd1r7l4c/MYQHYEvIzr7rN0
IEGwPNHoZ/hzJlqx3jZSG1H/eSZ1SwIh7C3z582+zx2ndlrDnuIlCZdsnZtvPFTK
ADbVs9D7AWL+zVzc//4aAc4i0+3DXtoI1fEFZZ3pkyn9jgyuMfLBNPSaQHUqjPXn
MeGzw0IRMB1Mh63piWedAp5fJcPwDssA6M57c/7GBYCEdAJGmMgysnv9y4NiESlR
YBr3iG6eRQTrKDC9elUFwsgDwJJNAxU4XjdUgwMaHCcIUfXpj6Dto8TktC23Y0XI
+nvQeg7zwWab3DI/SivS3RFskv9ZmISI8jzPZUGxFBVkFOasD/ucq2qgEdofh9Xf
PLppADPkFtqVPrkeBY4IACbGsoIma23phx9qfO5GXLIYYWSDJZFMm6epMUja1i/y
v31ISJWFG8pSY4ywc7H5bK4sdjsm5A9lOFVzXgzKIubbDw7TzQqgBNj0P85tUHhu
IXbJhEsj/Gvaj6bGtSgc/0x9vdW6mDeLxW4L3QdgjEyCROQTXkplrnllJqvaIteH
LsV7Is8DrdIXmoP7+uCvyAeRRIgjgdCt5ncFfBR0Hee/pHSAND3xfiQscwCjEVZ0
EZYqNPVQmTRz0SV6xq9zl1lvFgl/srWFsCKWZZj+OhxfjYWI0y/bqNPbu967d/zU
LPGgtq4EdaZQPsThylFDI4BbqPO6exE9xyz2sLRhm9Z0GDaLjkyGYYA6kG8eeMmp
9L3U7MrPiCIzj+6m+RgVaFcKoM9pA/9u9DadZa3h9DYaCpY0PEoB5YDUaV3GrTSP
qvaO/nCkDGAn9jqKZJ4mqXSchkZQDYxpLhi9qA1IwoFGC2I/s168S4gxM+H+jigp
mC0FpT3FT0O5tXPy+L3mhqnp+DxZJhhnCdVxnq8Y2rbSCbv19cxawqsO2k5QTbBM
GK1QuB5T0msM7RpgTGywD0Yo30sGglMVyo0TUr9vW7zcTrakOIJgVCVDlvE9rfb0
U+RIh0BFnhJ8Pr0orwY3PQXLBi8wMDdOSMCodvj19utTrPhiR4wnStgBN5R0O7U+
st32QGVovF2cOkpovtZmDkgqqfEqDu9SfZTK3WIaDudxm20RSDCJRs5YEF4JI9TR
2VZnp+wtYnOGM4tqe9ZRtDj2x6YhcFp59yw6uQw9JBadOxZ46acXc2BHZ9b/nDk9
G0qONhA2lgdk9KMK6wsfZ6fZgw6+oDlnmjdkVOPbYz0/BTEGYGxiqqHpB1gAn68s
JCsSi8b+WG82C4x4ps/IsO6bfNSbhVSoSOvszHvprQpXnR1FS2VVwkElZu5Db/6C
XNOy5e4X7cGEHGZ6s6jjIGZQpUXQjQgzJIXCnuQr9fcjz4FNadISyTep8KLt/4XK
OZOn0WW5sQhL+stugnYFhhCWk+mDPQvlMYZwF88YEWmIVMVlZk4j5c0SO85D8cNC
OMGSewyxN47kGP2oxMRRNQFB56ogNYJye2YX1m2ClznMjMBh/G6ZZu82k7I9mSZO
5hS/pNmBgVAN/iZeR21zqpVZ1m/lpVEuhZ4ahFGA8/SMuB+UJtE1ZGTmiafnYGtw
YtjsuhH3E7OButuJZ2hTQUsyOAXQHKY3FYOdyXdBzwRg9Tag0LcAcAyVR53oS3Bd
YpgN9q1VnqWItlTrSa7Qtq9bFyjxooXl49eytcUw2GYeA/sGmIEf5QiQbaKIwQxa
o5TPGTQ6ttV5THww9HJC8722kJrdjAm890wbLIMNG6kf5vNSifHLmNgbeDRTY17i
sKfGzwtKEeWvTEEIjyXTYRRTs0q6/OH2pRYOvMeG2V+6ubwy3nxVM8MJt81e4je0
PYFJaYmZ82S1BXA7qenk8XfcQjedOxJlZfxA6xZanF3usYxtm6kXmoEQRZfwIsnv
FP1MFu5zXKDZ/Rujn8nf+paOCHhpNWVoV6I9tVOW47rOc7vSXspLaOo51MPkObtA
yoOewn+XhkcfUwqp0jxn9cjqueAJZtpQH0uUA/ZXDoslA7La62EJfqJebSelWQC6
kvs6t/I61jkJMPkT/RYstYtvbD/Eh+sTLwVoBT8J/Pgt/GuwqwtX8kPqNraaJ68d
9s6+Wfi9tx3w5tPcn3U0dd6kzDsRfSpIgegtf6DavQCgukJRQGBGQ6JRMQbcD+ic
oMwUg3nCYsX3ikr+X8pe3JANyaiXZt01FPVB3kq6SfCzMt+eE9vhYOBzj34EVZPy
Vs1cplY8YLzIldCdOCoCWnpczrMLw9p/88pQvv6XDya8zQAn3Grq59bD0D41dHCD
L80LxzZGkHlHp50a8HCNsFPUyxN/xPpTFc1hnGr7EJjJ+x44N9tYeGVMkhgYgdir
Wyq4EH8XCTIBHaxBqOiyadlfm7WxO9aVcYBvgrT3qoXxsHtd/Xvt6okaNaEFhJvu
yvnSxBA6Xx8LzIQkKlKqLZSYyQSdDBR7S650hg8tMaWWSdM5MSd5p4sW4Nw+/vXd
xgWjdDUdwMs0dzTDpG1wFBeKudpr6hnHOP12A6bl03xEbi64hbfuiq+SkhQDGz9S
FWjaNdbKB731ShmXkTKViRVt2/uYyFjfC85TeCQM0tf+kbMW1Iuv1VShN4eHRx0Q
Fzv77h9/hZ9LEbyCTjjMxOmD0pZ9XsPca6NZQVUNsajklSA3C4mZdbP/dzjJbeRs
W5p0v3B3Mive4UVZObKa0fChm/2cv1ISUCwD28bEbcvjj+jA4PMJLkPw/FBuepml
Xrq0MtyWGeietgVgNNJubdMXjIsdKmK4xMlij3QAsn+M9h8jMo17sEWRn9cEfs91
7vh7CIhGZFyW+GJ3vIR5LPJnYzx7P32xKAEVAh7ZgEhqIfpM38+LGikwX/hb2RIB
kRMMs2C2E9EuS+dug/mXpomMDUKkpuottKUysY6KhhZEzHNI4Cakz2LvZcjFu7np
+gUncK95vVhDDVijPYX4Nq1KVzHMKgLGdBfIy68evhb8HeB9pM9EPX4yeMJUaIm7
RuG0lGZW3elVIruQNc3QfF70NU4cdJlaI/GZG9w242GFEG43o3x8tigXQk7KDwuS
+vUfndFdd/RGnor4rwikL1koA9GmikSsdet/Zox3s7963r2kG8S4+HlYD3ACVGUa
ftS3b/gj2Na1BTsuMMUjJIHqEiJ/TXZQCwyNHAU+teW/EXxBCpC5IG69d62Y6iAe
lQ2a0ESXQQB2TISqVGgKJFEAooem2Nv9/fFkblGPdpwDnCXYVueAgVHM/p+5rwfj
QOu3mul5709MvAYM5wIU/U7BZdBJXukcJi3Wbz6svJSI5FfmxkaIqkMMimcAG65A
A10v9GEEygg55rUqHVekqepcdiPsBJQxaNrfIjgK8D/XOftxASUdosneKDpqYZ08
v6b2O6XBo4G7mkl83qmgSoVT4QsS7nUEE8en2YDg7Pu7iC2m0Wt96gz3r19CrUb/
iUK1c8IpiS6ZVCXl0i7REHKaEmNqSSdDqF0uSEoKm4q1SWFKMy7RTrMmV02U2fGk
HlrqpTPhEY7TVY/aD7cLhS9XP8+HwZKGKj2wPCchjuckG+4nnp4RLak7AHaHFX09
GbFPQHLtbqIC42NKFte9igSV1LO1YRznK22EMEwaZjSumcglXuAuMjP/XVoVWvDR
LHrbl7eXdPoMjmnHkT8h0hNBK1Up1sNeMQ3bMr6AWmxckI6SqkUSLLklApis4Q83
PUY6Pcr81pFVABjtwNwEt6z8ecodiCwhRf4MOjlYqjiwpzjtsAG1GT/o/nXGi+30
rvAEZy+6igHeY2wFVzCDN1muC+Y050/qHjB/mYdX0CC+Z74OrfJwgsO0orV4mdJT
keDHt9oYinloAq2QUNrQdJnPgpHbnxqFIa51a0iDf71CSJlhe3afX6AAqaS5fRj6
7JX+stqmQhNIubnTHxu2M6RWhjYpxoLHyqZmgMPRlxQSUU9CokRBSVtX5toyIezS
dOvOVIqLupviHscyxxLWTkAoqMLj/S2TkiugkpSHE/1ozoAy0n+NPU8j8NjlI92X
s4U7JRbuLUXUgB/Dn9N0cDn+Cpqcu/4n/QPTJmYaNsfKZ1D+i+1rH1PmrUEciGs7
dsXsWSXwTIL52bl2cIdYFP+7HxWsjhNaGGmhIuRNkoIncz98tP5JVooO8boiBfcW
Sw69jUQgnXahiia0V/2ufOys7ATbamzOi74XWsMWt+CgoqusiGxVtIVAKaCmraig
MmI7awRe0/9zZV68NrReLwVcvxaS7k8XYic/t6icxhc3C00hUXfFCvZ06YMykjQA
rIkINw17ZRsYf2NTDMrVYtX+xFSFNpml7120HuSiv5AJJjD6cq4R6q5iED3vSjvg
avjUQM6y8wm8FgF60yYKmDCzoZpHe2w/JTFnxAmGt6swVn1++KhCYtOOS0gghjKQ
TlHGR7ttoZTSJabRo7e0BlENoJxHephAMqTXgM6gHYydhO7uXJlFKaSMzuAad1gD
6J4VfL0AulAkgbi06hhWfdbmNctcPBbtHnZyh8LyVq8r3cqu6p1tqfQ4x4EVPg/v
aVTSOpDfqF7kUzXA09c/3iNpzj+HmapFqg6K1k8tfzm40cF3tneRKtCFeeExFEny
RTbfEazFpDSMQ2K+TVNPDwHUKrMoFSOHiDTjskLLPY7JURduPpm2qQhSeOIuSLwR
CSPW/S3BZZ4k30vtK5y8Ok+omibxT6ypvoBtE4Z33CFyz25OIsc6RAHgOBWBLxz9
ITYU3I+hrQQuECN41NHC82BslKmUiHTkSFCZ2ZsJ38gvX+uijNE3bUdk9LOY5Fn4
OXCLAG/9mKreMFmWiTDxbmsmp1Jaktd9/6jz6OHliB6/ebpbElp1q5FrbCqyftwn
RBUupuxOtj3nsseEuAvG22B1tMlX/bjJ/bmP18qGAzMQDNPhLMA+4OFjVcU1L73R
VtSKVNx60wo5iyDpjFYRmJxaIJHGgXW9PHpKwMBDGwY7y9/FHMg8ujKMS9HDNzbp
PHPe+K9zvUFG5NH/BLT2kd6JMbrcl70BxzDSESw3hh0pbWCcj8LIVaC8y3KIO5lJ
YzLzOgOKA9USugUiEv5XiWEIEBAKKOmJH48950hyo6oPbmPcijNhR8GfN05x+8KO
qZGelQSh2qiaS+P4jawiPXJDf/L0bD+BXMkx8qZiEH/bcd6BKBfM61aD0akWm5S6
/BghwiarJjMOdK4weOyoxk24vJifmG+b+Nq70rCBOVeggfpxSlyVGM7TehT3jXR+
yjJ5o50/qsy0Tc2xHJU7fxvRnk+1NgdAhjBD3+V2lAeJBKLiF1IuBtphHsuKerSQ
pMDM9sbn0yiFKY4NmgBVczqFtKSyqEvzCvLqO0Qtsgo1NiD57TU5WzIz/ET+LSYv
rLrmuj+VNg1nXysacwNlgz8HA2R/f2gpskW2TsSs6ay9VEpCzGw8/3IMObU4IVzJ
+mu06XT4Io9Pzb2Y0CshO+4BSrlQH2TUuT2bZuSRlzVLcNolCSninSb0CjJ3vuJu
r8VdfZB4EpMPkWBseXcwsvq0aLY0K6tc9SexBYMcermLRmt3wVXV1iR72SHxJqjS
alhc2Ph7PZYAa3x66PqJIpUDlHmg8yRUWMqXJjACls9TksKuAyvxOkGZ8kuCVnJx
6T5ZGf92gpxnnIleud4SAJ6WnJM0xNgVwbD/V7BIQ+5wxM95Dxpm8XwUUaVPFmBg
3mtOnLyDqNAlA4BcvQ9KSj76tPWiuuq/jjqsBIBVVlnLHK79u5Vs8iZU8kezXrxK
r8mgdtu+YPWubo1X+kzb1o+KlFDAHzYm0YpbcCwm4+6ftYMw2wvFV9VFdx3URY2Z
EZZpFbDnMAeSLPbd/s+4ZtJVQK7kw1Oe4vRd6unCC9YX0hvLpZWXm0aINRrVwnw5
pcWZoXy9nKxtuLkkw12cymbaj4ocPdBCxMtfQdpRa5dP5rRMRyT4CPKfG3NpYjeH
j1JSYBpSGSJmI3WZ9sJ/gL86qilefM2jP56ZNwflfnnYL8WxQT08cMvOdrR9qf5X
T95R8+WIn+Gr48nH9+ITnWhUQUIp5zx5KhBCOgL01fbrH04FN2jn8GQm4EGMZpJY
B2nv9wWlwUGYyEn7+QlNCA6+g1vl8QVq8hruAdZW715X+cFzkTZaeibgWOMOocFc
YX5lvQWGyWWExUnPKCrNHYI/N8Zr+Q0xlQDzDKsJ0V4XZ14Fsuy6vGwhdlU0CqMN
w6dSo+it3qsaTq2ZWc+K8dOyxxcZI84mVP/P513jgcMTtriCNNnICk/VMiIq2Eu+
dEQ/g7P8Kj0yN4ZE3dWvp5NYvwMjZvFwluj7HKOYlJcDAAQ8LlFvm00Ec9jKaQrU
3iamtGBPKiKErSgyt6UdFb/EX4eqzwW2MoIYaCnrQR1F4x5JuDb5ieE2dE9AkL4/
WxF1iUd63A5yqel8im5vzxPEX0W7KedaEljgGGkdj9adkKUpROkezp1fkQlDcqEa
2Wt39s8Yxqf+Hke62+nBv2Q1NTDFbdicIHZyMiX9SW+efeDPsqO857IXTk2FRaGo
vipT2odvlKYQjVZRvrLp1LTqXu3krqWHsbyyN57o0NdfXKIUy9+9NsfyV7xAkJ5Z
Y9V/GeLeOmMZnaZuw0XX1O/NllSoC4GjNqfr+1BD7KTf8dzSn74XD6tXEjz+amYS
nR2xbuDI/IWVnMRjP0Y9dGDOhMgDVV5qPsI9GaQpPOrScWcq5++R1PBnPffOSiTm
VWB/XIIyBfqHew2RaZpfh7xLsM1mxCIV91WuFni+EnCEHvQ/BDn4384W7+bLk6w4
DvDw0zpmg84sUfgqoTZREgQeETk6wmBq6Z0LjjchrCrQpg8gXz7xypxGyrXi3dx3
gpwkyYVxyHFApp4kYChukO/rFgxGYCs02IeV0REluc24gghHaPn/Lgp58DwVs04I
Fg6Fsq5VAxKj5RyOzf08yC8cdjEdPURU+/kJtTFp2VbB2uyKExL4dXwSp+A/15YQ
pRsYT1RSeeqDVLGHbpTU8OkQoMkzN32ZhDhqUXze36PvELcn/3EkK0EKdoVB8JC9
HFds9tI20TUiGSG5kV9SLdccONlafobhIUH4K/4VVcW9UNBLUrw8QplIPXfa6pIK
Qs6RaMYoMEE2i264QVSnLXPiYOjCxplEcWdh4QwvUeHbXUk7znI+KZifDusgDAHF
F2GuT8QT5ZD4dg0741PTjqSHvgUxG+QmOD1VwT4Pf/qEYmdckpNXZHloQKTVac4y
kc9kih1A6Y2eWS0b/ZsNfkEKI0wQQNhrsvtOJRnTTn41Ry+4Dpe5ofKAOpEELfWW
1uLOIase1/OaZDA1baMxk3rPl+YGwj9BDrPEsk+CuIXGIyBef7g5unpnGoQ9QN5f
Grc7LD35PhHwAn7oBglzvhKTSLFrJGi+0BgsVO5ZlVwCKzipVKkRsYPajGzdiJTy
UCYenj84pvzdQtCegRXD6FdNBUfSX0BRabT7sgpLsRz48fKyatRBlrfBPRRSZNiS
lSbm3a/KxX3hq06WbwwIcss4ASgBIn4R91z1objvTb2K0wmZwg1615NpNkU8BH0G
LowtqCtshCy2PUiCvz0nzjYuRN/iOVfnNiYDpDmRJVg9nzZLh8YdEO5cnhDjkA8M
wdsI6Zz/qkofIFK80QPZ8jfiahfZN2xdj6jIKb1fBEkCs0yF83N/v0uS9PIkIB0d
wDabnMAH0jMQUdEI6+brdmJKrjLPfXufQTuD6Z5Eknp+giZ5THQKKrL4wCfujmD0
UC7y2crMriVZQ5Tm0qObPFLJTDANdo0a5ZmI5G7BCJcRxV4XG6mVpvN7BWis6J34
dBZ8BGoAOWv87b1TVOST5vX1LO8a5Mfnarv9I+rd8Oxqy4AO6TBYo0HdT4nWboqj
aUJSphpFG5qMvUnHqbQE72zkKYwfiQSApPw4gK+G+BkjqP23QBQINHB2I1iNTld7
ENX8KIzt8NJSZtZHof1NEoRMpnQ6GHvuExE5xdVytVHRJHw8xeOMR2MeDZY4nzdf
3GVrClCx4ePaiJhsEidvvPM3IiM2x/AKtqcDMS6hDjXo8Xad8vhdbRQDiXjoqFG7
C+rVNSsGGyLNw2IyGXMnUQ+ZCMYF2pVCbex6xIvphlnOcUW6WdC9e0NpSEiiZH1O
UxSCu8tdVxL+JQGHTlUpb8tknjVIUUbtmyNjPfSwyBOWNEV37cdG03JIEdbz2yi2
PWo1MycVtdPXZemPOW8AkLjiPkx6QjjV8Xhfuwz9RHZMsLP0XweoWneYAeCpOulJ
4p1sRB7PHu84EYagNVdO5hvd3tQZ2ZLxjCoDphRZB1EgRv3kVIlq89x7VKyHDKOa
RDO60eXlH6nwL6psQ+RKzWhT1bSfXGfFqTRv4v6/dyDHS1/qrUXa7+IAB/4JK8i8
44aaoC7s1nf3hPJnGxJkZlxmqcduUvNrJz2ddSOJ+jZ0AzGElKzmcnga/UicG4ft
InV3CwBq6jwdj9JqAdC9FRPk1ez6DPl6Ip6wSHSN3+HyZkMjF65XWB56kzba6fuo
IpBllpmaBFcY/35ReQANW6bLOTXgxYtY6/BVFj2Fx9/YyjbC6PnwTHCxDtTgHE/9
HgNPlnW3mTYAyzcbOgcTZTezlW1s5PA6YDWke4imB2dCJughrM8j8VNDQm2B5Cg9
Gp2slXCP0bUho1We++/Jqu4Mz7EtKQyoHhSYN60hVQh1Up5FdDEAQY/vpmGd6ds5
pknKKPmeDqkmfj+Lgl5Km/vLRIOMp+pxPJ7NfqIEZwX0NCi40fY84ukaRGvRxQyj
rio8k5e2Gdq8iMkyPLU/iKOHGodTuScWN8CUHXfDxJehvJKj2zBV+2GHjxUnzq1B
O7oMBidIYOUk9liQu0I4UbiNXLCE6xyJyEYU4TyWvgYgn1NHvrvTqovQ8udIkdAA
rF5HsN06rNIwImODmBq0wiHVHKiMWQ9JOAKE/4lXJ5yw/clGmy12odVXMJmzQxDW
AaRvuAyNYG9SYIS+vOMOtRC/RrK1R4vYlfwZluFNHbf5Nb+qqcVehDChWxESJnLt
F+JU5hkkwp5jwMIEKjbQtEQoVDsQDpmLKn34FkFXIjzkk6yHu+BEXUbGxlQVyOAL
Z8mNmwp42/TSMrRNUrtEKGNzeYU09jT5xhdKl6HnSI2yQs+HdVU3BJ52wmXcY4+d
abzD2/Sn+UzQHNVKrix+P9jVwRm0228x66hWcVffMMe09mGsG/0ZqGPSYGUcU3Ys
llHu67JuaslXAv9Defecl2v61VBc04oA8WopnALFzLLqfovj1uOFyX6/crboB9VV
hh6n8at+7tuwjUYxevdZll30C2Mj7Y+tfFmIcUUy35ZQ3KCme6ddxu0/WpPgb0ik
MaolVtJvr4Cq+Ik1BscJVs2140a2ORrVUdeL/IrGrZVjz65LOf4agQXkftsmHoGW
8U5b/Hw9tIPhytJ0HM9JHPDt7GebUuSGvI0oYXio/N58OJAXS9x3iwdD4BwtDqxO
j8KwX0INr79vqrAMmH55grkTcRVg3o4pyrSQody4lVJ/SiPioMUp2zeuzB4VAMWq
8z7scZ0KRD7vBU+PpmnIhfAfjS8XCP4r/YhgTWVbRdjQdc1B+kjVnJ4zOpe8/rA8
K5ndpb/Z4lWAmadO27fp8mgMralcEO0QeYRWw0VxV/y1UUu5RO/xLWDuyiIfsJXZ
/f+aUZNndCyp/mzZ/j/u5YTQhp21ZeRebImDrSUrQb1dSZUZL69BaP9Hla/OZNN4
vTO5AFqcEA8ZJTq2UZ+JR2pf2TK1yq37ukT5P5tYr0o2zW98D2HaBQm15ID5mBzZ
Ld3zLGR7NxZ/ShqHUUby3DKFFGIUZy0/Xzkio+n41QrlbPG5msPC05S/g3tkKBsT
WPPKZV3/ugm8v2aByx9Fna+DOgijiIbT64ToClIeVwB6iDa1bZTSAOeZtb2aZme7
JAcPY8ML5qyUBEDdeixVIb4X4RCAJX6WU026jPiaKCYM9rFNGtpaiHN2q3U4CDGx
g0+M53SfLQtsDUSMc83j3ilcVNbdjbi4YitvzLD9JEeADFXyXK1spMpJ00FKVl6V
aX9MJYrKZSbeLAmjx4VUiLdp5VhSDvZ0bWxgF0EHCKuIj1IJusAG4abRHrnVYOPp
TUuo6oCEWgp8fbu4NWdc9f5DPM9kEZQ/71qMmdyJ57y6veTfOrfcbt35k/AUoRap
Am6rnzGmXuCbzWPw4zYX6tI87HgT9K9EAZBqjMX37zMiiV6M+BgxvpANqSNx+gc5
84nLcRkbdElPAjON8+qXg0AfCPJ6xvhxPuyv5/ooSrA3XL2laRIUS66mTz0XrJ2x
EhlJTqhODKfJw+m3FSbwW7q+Npe7MwXoMpRJQir4osFXEcX7tTuLY6OJPivPB8Dx
0TeuIGUMNVyu2VsIHuvPrBCO3pokthadqDIGnDH7O6S51KKbtjjW55nqfxNgfr4J
u6KLHEsboWgyVAqeqfS65YKGZuvmg5wDxYcIioJO39y+6HPK2QJEsEMpoG12ieyR
IlsX1M7Dtp79DKc5TmJeaObebvlGjmGdJkuFaD9mbHwMJdTGGZpqDq4karcVSjJ/
zDiAnJyTDmpaTalNDyGro2aBkfEmIWfJGUGsxWk9hUcYOOqoaNriXEH1G6RdLgFW
80dO5/qvOh9N2oI4HGxSX34JPClnOjmGRab50FdpdavMNJ0Js5pWRnWBRCm12GEq
KKWy+u0DtjA5PvoRAyzMbAFljRS6JcOtSLgCKRIDlqW66T6B24iwC9YystrCCKG8
LgUXmJKrFqmE1ZBU3HepPPj3q7B+js5G9cQHg+KEPLyPNVVX+yvkt2HBwS9V4qNC
QVzTDdjblYZ892hKLOSnkd1PR0126Z9HXT7wmIUR9+aGv96KptNhrfp8hKH1TjI9
eoOt+SjoI3GYRXMJ9KARU9tjNhYyRJ9qxthG4xmvbJ/SWLcdRfMNi8sbvM0oBQVM
uvDXu8VI0Z/b2mTAMVL/bv+iqJ4DCgVmtHWD9gPOE9VlSD+jGvB9Fhf6Pj03EZhP
NzNIAjR/VVXDlFuG9dgAZ930Zo1CZciaDeEhlns7h931YmKsPizSCQEaxrh+s1Lh
2ppPGmJQmPEpWg+UHy0jBdTIj9heplCOdxbHvPWKlHduvQhfXupwuzgYnQd149Wl
hs/Bhj+/ZzKIVanp2lUn+rWdbMBrZbjZMXw5GeXI7whgYHqijPXPHA1nGi7ptKWt
kHnyKIwR8W3guzewFqbR/V8Q0fCegyDRtPoAXTxYEfpvWOiHLYF5TtPEmCcxJPX2
77Wy1kPihMYkXngiFz7OHklDdddZvvF7ttKJ5X40mqnYzSby04zUVFrOrotsieJ+
QfNTn2nATcs+hMePUssMbOVumPE/5bW3/f7YqevWcr6ykk/x5cY2K63QOzv8OVTh
tUbhwbNEFPPzgQnMX3DZP7I8WDneyUWHICeRgUhz3w8eAGgI7MiFvuCZ+OL5z4c3
ALAf1tXZ1IZn3Lyo65TzsCHCRAq5NRCmjqcx00SgMJf3JO0u1Wp5qQTnxCw3iJwQ
6HQaxOdYQ6nyEIPt2gdieHRq61dJK/LyBSm791qUhl6tofG89DJ4YsO9U4rT6QkW
74TQ2sHsGHPRcktfBf4QZNll6r/jdPHXG46Zh3hVoPZyYD61csbvuTkhAuQf2t5k
dI3fnOi96NR30Th7+a4q0ybLuxHqJvWYF3xuNj/wgNbOdCHhIey6vEstwD0U4G8b
grAsuGqx+lwlgR4aK+n/mtFjwacg638gH2PZwmP6C3c+4sXClGQI/2msMpECzZgv
FSkMkaFsutg6Er7AG8uMCokeZqukrq2RS07eqp5eGFnH1bngiiAN12PAGBjVdSJw
TP0e2IhQHKwiFX397IXlV4yEHaUlG0ZhrIiXzU9faY8bPY5Zvl58TtyPf9eBZvnZ
BsQmDTReuT76kLXc2SC/Xkfk3AFaqLrM2Z3W089pWYyf0gXO8WYwxQ6tBZaVpthU
sBZTBiPy1d/aktwLhR/457mL7u4TN+2n0c4E083xpBk1mN9aAfo50ncs9dN6+P08
T8F4uBbA+3O0Mnlluw1vVwpSrz8swJemOoSZSutZYy7/W8EKEBGJmmwasLKK92cY
R/Ux+D8KUyjawkJHt8sTYUZgXrYXZY3ony294EIMo8F5CZJvpnKQCwv9kIrtD8cu
ClfqYrihmf6NiuiUDpbV73o+MzDXaF3vEDY8DgdN5gLu39A002MxUG8r1aaJcgKO
x+CwajG7E0sdyTeRhp9LSr1vW/YX/BUzy0HhJUJIMxWGK41Z272s2vdoQOmPurpP
Tead+CERujB0ADygUemm2kwKcua20c7nJUthMZhYfDJzsOA+2tG9z7JF/1c731Xy
AsjZ0DA6B5wdC5DkUWhSMlE6UX+mqnaV3g0Tm0LYd4HH0pWFVhty+t3ezHYh9UQu
FgWLgg31RE9GG2vuYKUGy+aguSMRO6rh/KsyQPDu3QrXedwMJGrJWpvqX5XbHRkC
1nAWvaoOlHBpRU+XRFIZkbjwERi9wEYBgA3lVlqsVr4fwGOS73GbbFhm5yEWRUTa
zBb09nn8jNESKOzG0qeLM5lF0jQAhfdlk2P5ZwKRXCimBGJpEyy/dEjGIzfmk2zG
1ZfDbFGcQR20aMyvSjozFPSaUZ0oUlEF2BThr7lkpccsFKam+qWrja7DSQw/rtTO
ZxYURmCLz25yt2AlvTDNw0w3f0NYbnYM9ZggKf4AO6SMucRApSnhfV8DfRRMoq//
EVwo2lWb0UNwaa6q1TEPec8HX+hpBig6w1yZWdRvITIDm5BHXc000Bfc0F4DF48Q
m7ILlHzc67tfSqz2JzIiEtmbdnOycsmxAz4hMJoUa+vuCv8GcAs9aUbnbvlSoRHX
1DS5k/s/g7A/lT/YKpTLIoMZotkfMeDcVcw8YiX8nUEWF3lj2SWHiE0yB1j6Cn/P
FA5f2C1m+oHmcWjSyKvESUgm6RI9ltu2Y+5yv7nIzimaQJAcpHGQfjYb/8Na7jm7
xKB2/srYYU40nHoZz2ZtDEmRR5KY2lZj0/5HJ+TyMBFCMJ0u6OrBtI1zZ+akStWp
bz58TT3JCK29nr2OG2sKAj2/jUZ1lRZR9n783hVAKad0FFnayMLVSqunW6U53q9o
uqfmYclnaKMNkK/etfrpued2/KApuiF6Sm+f6nRfW/F7HwS/wvXGaxpo71B2BfpV
dSvUb/t/v6eELqL3vS0mHmPa1pCp3bT1tWyLNufRC+0NTmyRnJM2B4SCZTyne7q5
4xP4Py3rDxa2JjInxTEyA4W6JGaWGjekL8vFnEDZ97cBp0+vik3eZ3WeU54qQgMr
hww7AhKwKt4AkkaoMVDa5Wej3juu+iRTsRKeU8QlMPxxz5OUIopDzqxrwMfQ2NQD
dTvRTi3lxqg3mNmGipd2k2ZgxOn5Lspu2fIcoGrCCOVj2wi7IJEGJMDHL+lSh1J2
Zr5whyLy9c623u6IEmtzwSMA5eGGVWHdqRm+BherNPvQ4jWjRnPPDeRLIgczlxQe
9hPFrNMowiIvjB+8YX1NjU3qRdqs4r02ZWjpoKb+7QY3/Dv4Ce0DD5AY/dFpnMsc
qWaI2084wfLEb4fJj/rYeFWkq9fMWTgjP/e+XRxO311cPuLHYo5Yx5DUJ/cwC+qj
CeKBZ6Zl4KfEDunBgg4LNW1P2J8HMhnOCGJ/EUcAMMRHeiiIOgR//kbZtRU2SYnq
67QyBdoLplrRXMztLci/q+JBtTGwnBfL5ixWMeeroRA2g5k9jcPX3fLWE3jstwNV
D3lT3IhsGGN5MXnEs3jzi4vejjg8wflUpcwiqMinxNsOhfODWq34lbAwH+F5dSbL
EFGjUL0Ddcun4w/H5ljIhzwD9s1pIK6I2YC9biykudL/4RDyAdYSUkU+UxFn3g/9
34oVbmtIPu9QSO8BLRizmHQANgcwkHwU56iI6kkDSeRbETzDkiK2FpUQ4YpWOUtd
y/mavQrAxOH8j5OiSyPnEDg1HndGEBtGYSKxvxQc7WZ3MCTvkNGpQRzcwgWnJupp
ypToZqJ6nzt3nnHKHu74fifiIJcSFtNdeL/cFxD+eqeNTqcXsSuiDZvJPnyYrVUP
w86BCy5IsOp5S8fVbcZ/Ikk0BgPn1hmKOJfJKlJt//RELjLsnnMHb8ySG+r5D5rE
srVcMe8r3zm+D2on6wP82sTUxtwyK2kUggLpZsW72wDLCLYc/CHfOaYZUcIb9zLr
yx3Tqel7C3mUtsdoqiwFoMK1Spr4qv6OEVWkQZRq/tfhIILgHgg94OJIo2f/SHgO
oX5nLu3CH2zS2nean1hE0EPHYLDs86d76XoOFISCKedlVoVYEHOIihfWHIAe42mh
Hm+IzQJJWHmWJL9B3FCvU2BDQE45HkwRdVmeEzkzLc00bBl6ZSC7ubhw8+ULv/bP
filsw9QqLmw7DQLhD0LjIgPFWH6GKSchVj/f77NfXjrUYVGE8gmJf7oH6F9c1sju
PEclIUDgOYhWhXDYEaIcK9tyZvcfbsJKwRZi2Hp/RqnzX2iix5r/CTuf4LMR57+2
+40YnEVCE/wFy5VW5UxBUbAhub5KM20Pl7PJ3vIQovahIetS9g5TCBQ+rzLTRPt7
PTG2ntFtjBpzqkma43yssruTFbivoEnSyPI3x+keVn6SCL94PszBc27xj/KqafMU
UWyYebjaZKM6TGCQLTNq8r57qVjLDIHvUXfh2O2tjkrdLz6ubkCmRXV0c3kY6CJN
F95wxy8mDonqQsLrJPYwwMaRdkNcxrE126WcXtInyNjsUbeecpPENqRH8coZEOqk
ejQ6rDyw6C1AfpNfB8F/FJHSqY5hUz3xO/bgD2Yb5MgIN04d5ZSY5i/3ms7Wc3CP
TN/EFMdX5ECw50+kj733YJrxgCycQl6Kl9AXOq0HXppbYpS8LKy1SJ1oGkj1Fg4M
o6y+yrVFcpjaTMAek3VPPl7a2E7qBzIXKw91rRKNn62pDZmzrInAceMGiJnsvPjI
lXYuiwZzz5X+vrJn9nzZZkNYJ0fb05jLqxLwA+3QGA4ualMCaEqIGWxBJZD7azYa
q7OtJU25e6kNugcFwgA8tDJZQnE8hhhmle9JVAl5K9wEj23uRomtO6MV39uON8US
PW3ldR4GQxICiuthQym/pkojz0hctlgXL4bfcZ8hMAUutZTlpGyH83DBH/9bLjJq
ovLeZAsJsk6EgdX6SYuKkdC2j8B+GLob56zA3OOYMHD6oVuqN08sYl7VSL/7Wm3K
MYF/VsXSU4w95RU/1HJuqoPNySPy6pYqn/jkBalSxIo9ReHbVmiZywkrEWWaR5pm
SEXMjNYwL+769ViLxq8bGe7W3uTC57WhzqpORfM4Do9wSbucN6NmJEyxhyn/OY0a
liWGtAjsejyntpGDHiqiV9LyoaacD7Li8RNqalpe6jB6J4UjJ3UrOn39s+PBLAQv
Dx8Iu8x5P41BsMVa1Gek+M49IxzUw05okQjl+lTZJ64x9p0UOYfvKmlKRbLFT9Rq
/pjT4Kt+eqOeJq5wLkTVQEkPpdLXW4NY2otfLuRT0FxB6ctlSoU1UjAiZwlnD2gb
7IxO1E0+xJv5Q6NdOEzuPQpbut5SAdITzTfxzDdNRx0WjVi1Ht5G7vsaVsmM1mHN
sCRU6AvDdZNVza5L9R/yflkEz/ACD/n7NrGzC6yYcldj3E9VfoeRXD+hs4yo75Cr
Rb2HfNc+lcZX21pdYstlIVpifAENXQjDJYC4ZlKj3sKBEXMsM1ImqcnZqzwlxVry
M4Du9QAnJ2op7C4pn3G5edCdtpQyj4MpH5J4yF0cXrAEqlq34LpIIh9wiKsnjsrG
QMTb3sYBmAY52tmeK5Dib+M4KQ3nXMkhgJPzdGBTGKCpalYKbOUM83440jNRHFSH
0mQnFkrE5XQglQ3L2x4ZNba5lc3SnNTqrSG9/1lybGorY3DQoeQnJFd2Dm57p2tc
TtDR6N+T8AOM60+7D3Y3n1r+NB0bbYR4SC+MuIeWTr2y0G5VM8DcUqHxX7Y0ccUL
DgO1c5NwopyazWUwXi0QJxbDgBMfGgx4uBlQxNR1vrxIsoKl4VwdFrBuV3EETUtp
NobBoV8xtMf7jERRSPFUM6h5Bk7pz0ycOv85x8ZA71DIne1wd8ugZphNB06ewS01
obKo4zxFjC5NYZS2o391rx97jX1dp562AQxmVKF4LfVR5nzN4tm+e/dlc6qc/ozi
AN7erxnr/KqqDti1I+DA1ncjVRp/orWsoSqe6NneZZwlrw7g2uir5EJzk4YeT2ZS
PRSCDqHuCmWetGCje5myua9geumITzqX7ucCaG/WaCA70wDvWJRNmTD3mvUbrsPM
ewCTXeWWNT0qgMHZe2EQ8WjIyBQClLcV0I/vawZholXrO1qr2io/JDhtzOVVeRU7
YKmNggDEXz3Lv+FLPbOUoH/2JWIZd1CzDE02ZQQCXbKqWhYjqBCyYoo5X3OoeVke
+IningEEdSDxYEbiHfHiXPdPz92VqmvOmiIy756/3oeGIn2ayUzzIksHOoBy0tIz
vDwOLujsDFEADakCYSI4YM1B2bcBJ8vOjQTLL7gU4MCd77JuoFe/GsMveFVIGvbh
AKQA01p33nw1jnC1V2utQANEB29btYMVCORn8EG8h9AXYXFRo1teW4NKZpRrqTog
3IFM8V6xC1uXPr0TOHvKzRauoo1XrICXXdIocOJwYbvDkXXJpuTO9BOSo6+0Rzw5
KaaS+7dy+nGn9UMKXCeUYObaK7BvR3un2lwCxHpPQ1G845nv4TaBm0EWL4vT5tkX
PuXvWtY3WE5r/M5OF+TmK9EFntD6BqwfX7ZeyVymGtPEedPWSPX89/SHW9+ytr/f
+1W6A1J2txwSLbOxa3v9eZ3oVa1itE/2CLiEH8uOJx92DC4T42wm1BqW1CZiacXe
dY88gJAqwfalfXQm7+i1+EodQziAHbe0J3/Mpi44gyILeS38Ee3rvNBsGgBbPmiF
iiElH4lcOdcfsvJXrttdZTxTFP06OF3Q7YMOGxNWLUlqREiOWjqu8JDlUDjzEdY3
fBUchy2xExymGUE/soVn3z0iaLDfUDRGe7hVvX4UfI1PtZk/siKLRlZpNcPsrLVg
hGYPMZhROICTcF0JZB3RTWY4OTz5H+3Y/edJL6bqfbBwRMcVLl6dTA48MqgwttbE
p0i4UUJhVHx8i5zSLIgMu4t9kVqnL9sabWQcgfkv81nFY2j1NOi/zeXjS+9Ue49Q
Nogrf4BzZtTk+07obBvo2OYpXT8zMBPVb5DTG9A0YrsyLsHDDNXnzQjgFzdaJJfc
TUPMag+ozH35HJ751xH9kr3kvwMwHgQ3awZRnGvmujcMUgpv425i78MTVnnW0Xn0
750nASAmMxehO3UUMs98oJR2yEkaYAJn2Cpzop5HEXycRkgLYqSQVdKDNgsNLGDF
xr/q9wp0ib/yIBnanPN+GlfeOma165Y6yQaR/JQyX06fwJhsEMX7/jSD/xu+ebcU
VFzdJtSZSRyCYM/2m23quN+nsfvkfKjbH7V8eO3p0ojEl8XZVCjvA+XaN1JPyB9C
iN+a02N1Rm/Gv52LkgKiDeIEQv1zl90SFJL0dgDjH27F6WDEVbsUsN5bDoS8YtO0
OOA00xaIzJBMUK/84bflIu9EGZT8BgV/iLRqzEQzgddM2OgA9mIKniGJSjVxrVeF
ASuIfCAE+Md7a6ratZa7nIMYPBRFZ0iX+8u/S3DKYqU+jsUhuhTMeWlDJgWuYpLK
aNGevSJUZtU/5+LzbvnaeiNFRcDg85SyDZ5hR7yRJJR0fokn/xiHwJOL4gfE2V3n
FM5pfZPJpVHQseEYapxR+Es5RC7psbyAdFIr4f6ap6p9+2UtBxYlxXIoJPEMpcDE
lWe+u123+MrOdp1IwjjlvZGG5SiWtQLg9wQVQ+hU9ufjBkcS3CO5Y+W9meKExu3Y
hDCtli748sl5he+2skKj3F/MDl6sEFdKjjLqrLKxmSEras0X9irazEWGVwniaizq
mV72zZwEy8brbR/Soir2MDg6U6W1naPbquecTJgEJpOOcXNkikqooSGZJLP+iE1y
rrOAIhahTUHcDTtvH/nwHwccA8uDaGFNj9cO+jr+ddGrF4DyIg8jXqFYtO9VirN7
Ry/tELFfZPsfznF0O4WB+jrNUm4a9LKC2eDCdMXssGMgn9wBa4jSFxNTa+wxiNTs
iF1eIepxJj4NjuZielZSoN5+DLhIPjraY7hcKZQClWuwIONK32rWIuYNrXskFroJ
vK+cvp2mQezYstPKuwUjU5wOwKP0Ec3LFfQGXfo/jzpwDMtTNL64dcY4y1gBJlpZ
PlDT3MQuqKaliXQM1VHtvHWvYwTvYyreV4HaxHyuIMA0codfZS+KIzot+xg0jzdC
Txd8x4iZdre0Igj2iRxXhsqSR5Wr47//S/1/zquiRKsc/cznHvC7kwKffrP3aG+0
7TxbjLbl4Bz4MjwMclFWlhLBCO8HHWY9yKjtJcijh5Ne/ciWTqZzjCe5NP5Uff4F
tnI8H7QU0lzP811OIUvwznzFt0kJ+7gk7RcOsZH1JGLBFXoVYyHUG7dTtnQBh7mX
wkCgEeT9YkoiFvOHCNdBkiCZb94SRO4L8RkUhvnyDa1rya/0Hr1GBrIKYq3Frs2N
UcElP0hxisJQR0y3u1N0akIQvDIrk0gbPv6g8KVnfeuPBG+aUn0r1Btg3xwSl8iG
6wLadQE5jd1ZE887Qj9l1E3TImMNwHwAMbofYYJxqx/p/ZpnOUA73UyZw0gwiWhS
hRpU3m/NlezWK5wJw4bGAXMaP1ZAr/R3mbiBFJG2hJ5k6avUMy38kv0ruiMDP7Dm
EUQcZhKgHsubOeLclkTMxYXW/rxTbFMHon0wdZLOhAL+OkTVskekrjYiaprQzAjP
XrROL2avW1KvdNLBkB5ijTsS8Nrqew/cy+7Zm7zLKh6Sc8akVyaFDq2Yg/iaszir
cJ5ZBNvDe/W14x1D45a8YJkqn94vPQrb/PhZcSe/vYlbpMD8qSjPGf3a4XFrS3UP
TasLSU5IeHHu9ZneqRthHGKXeNDq2uRSJAQ0n85W9D6insn1LjdF1VIWLUSgzJ77
dX7p3kMIYHvexHOB8BncLOyK1z8wnEHSKVl4Re1GY7sK0NcMB75hbc+5A2Wy0qOK
PyK8B49W2L2EjsSPnl/odDiRtAtV4HQMsbPy4QotlIldE1voyys+5Xgaa6V6k9kg
STV0a/mXNl53qDj7TCTpAN8hwy72+zBR33QvRm6R4fecymTHyj5pwwXh3NFcgFvz
pgwj5XCofj56FfkbyXe+Mm3Bv/7UYKuMQ2OzsaOeLXJiL59wzwIK8jh0Uxag8gUY
EvQhbuPNb19EQ7rrAu4hdV+TxYUuNYsCVIGAhQdF7fkwodqUDSZgDVeRBOuDPY4I
u9p+EmVuXwBhY9lZWJhqpZI6yyZ3M788UnQHhwEyV9YUsz/PTV6HFE8n7lZKntY0
Qh63WqwW+c6Mv4wPMKM5Ev8lNjMSZYKcu/bEf0622K2mSX5Y9cbO2GqtT3DTZAA7
n4LT6V4ycYFk3Pai/hK/PlSjAaMUe6E9czMovbRAkiv0UX8U1Qxu+wuF44ImhgXM
SyVf/6CgDwVerdDEUcylhDXk6wsf+Es2Lu6BNmb0WJew3kArnMoAe6fZbe3OStgb
yxEzgRUJ3XdwnF39GHwm3zROczMQaZdFe68FMDCvsH84VWnUKfVvgtncK7idpkQe
ZGD9c1hb9YKLWvqVm/ANs+ytIWJHR8p6G8nzNLbvX+t6dO0TD4m57tSKAxZLCGHi
wurgMZqHyXFnyKXbhG/2dtCblYyGp6MSOqML+jAUuDEuCtFBbmdUvHhqvoOHDc0F
AronpS8ilTsNKjb9qO++aUi1raGKQVLOi0PG+WPEAur3f6v5sValI9rD8azCKers
pHn3jh5Tjw3A2WUWp4RZHEZPoE6LqxyyxJYC7hCGexWMOrlVXUI8YXUfxTtWp9dh
Jgez6J3PKM/QBRA+jBTCjN5XPvDp1mkn4sGQPdLvtqobSY5rXWwJCyXMvhYNqEd3
p5gfXcDkkyErg+DwQMuk1T5Mmca9DQzaFqdP8F07tewqYut4tIoL2Rfc4VfiPBoD
tqNU1OjZ3HSZKMgN2CjKkcMavTWFZt8wiKimARY1kAtZaaWiHkYa9Vxj8nvBxz0R
6gCBLKCZV7LI6WR8bbDIfxvaR1Pfx+Elo1FZgpd3hoVS7JpA7363zCOjfGdHoxc8
3qxaU0qAYf/TdrJZGY2aqoYV5v6AT0z5xGKisoJVujLak3n+OxornUnge8NLwtBT
dh4elki/ePXkzj3rq9wR/bgUKRYZLPL0uBG/NAmEywKEkEMKYl/Kxu6MQ1coojfc
7LerAjEF6Nvn0I+8I/6vd+U8/db+Mh/+TZdzts6SeJDENxyMwnUDxdUON3Yfr3nb
kGBIfNy/Ga00fx2AD9osDIA7uwWD1B7B1Hh1OcQdghEwfwQLYSG6LlqLcSyRySRz
0Je0RxFcGGnB0guNLDQpsvbZ/vF5tgTOlfVYrek4k/eFf9aXXTn9P8N3WxcRxTxF
pLx2pdOwgixcovF87lsAM6dFWYjbL5/vZcmkt9Zn+jnV5mJtK3Xe2ksT0MZoaj2P
rw3omuGQblQS08KphqBD2q/CnABPF3F/CPkUz8nR9QNh0Ar3ue8GDZyQAU5qxyVn
Bx1FOMcvv+ZIecUcitw5V/4hKGDlhkq/3EgY58DfguI+v2AnkygxhIRddSl5WfoV
AJR5JDSre3OcVFJ4WFXZZH3FUeK/jYcj0YsJ2glPFhW8QI0DlIf2Pf9S9l04POlX
kpCV19RrV2OgCc+CSHofAqECp8GYTB2R9U/0dyTFtrIvPmahTejCfE0lgW3wO146
xemC75XJZzD1XTId9IH5QK7PuGarRDUOTnj8tA+9ccmShBRHACccRC+3bmk/7ku9
Dq4bsI7phxoDPYlvNjPMgiAbLzUY6Lgr7VkSPgsDKCdTYYpA6hB3E5WiKUZBfhXp
l7e7f4lRnSZsP7AuRZS4C8HzS4MDbJVyZC2VGAF8jzhSWGfxJiZAqqNHOP27yFXs
dxPaVsnsaezqniUuquxlZ2dZPmSjGMFBe1oA3C8U9qrUjIpDhakxm2nD4LOzBCqc
iBExaYy+q4euxF1l6l2gi41iqiAQOfyUYvTTiHPWzaCkVit6sszwoDQLfoAwNwvX
KOiSCuoRlRyoRlwBwufwkf/WT7k4qILWFJYRxnjb8dxYeXqBP5fWec1cS9CsBwU2
62JlQA6USGd6GF2Dct1CkKYUZRcLVPjbZs5hqoKJrfZ+1jOQ/aH2jVYAMydPf89i
PXpPlMt+TZ5cj4mqT3VqvLRrvp57DbFu/K2S5TgNmXQnCEeO1c63wA4IKTMEabUW
vPaPHsDw72QluRTJqwloDAoqPwMBWBnFFSQ0OBo45TnRpX0jWbcCcOVMzBymO6Nf
b3yLg9z1nZI+XLLBYw4MwXfKnKZ1GC/4mMRj3xS3Nr+ZvC4Ck3nhnWh9E/bWb9Pt
U5fG1urDkzxOv8LU8Se0wFqWwx9eoJT8tuX1j0ZkDXPGD/jhBKm/Pn4hMxZnBoJ2
AeD8+jysuIWGgHM6fyeV+sAzNBJ5yI5s2x8Ex7ap2XUhVxWnQ/cV+lbiPqgljep1
xHsk8iTn0t5ryjJYv0qpncQx4PHFKyUAKkq3aGYrpahs8ocZu1TjTtiXclihPQWm
fvsC5XXgzewxwvyZJ4xIsfLGF8mfPUMRKxpobLTz4HAMhwyu/bNxQgQ0HxA+RAKU
EKpPEn8y6TsvoWEr1n8N52UPKC3ORag5AANkwC/xNSN7TPkOwp7NFJfpqoS94QZR
G/jMaAPib14pLRj369P0AHAWsVYHJdNYfXgY1+pyPtvGJ4MjjeFA3AyQDeZTxXCM
libikPikJfXUCiT0H4PntxF938qJKfjic1IqOLGvhb4J2duedPnqmITct8vG/7ez
AMyWUUtOAR/1MPjTmlPjKYa7OVo8eZk3RnxHbMP861jd0pjx9QoWfTF/SrLEPkMw
kLPYt6aA+4z3DfKouavnKYemKI7vZ4Xf3gb1uv0hfgNiPiWL1x/EyWStghWlL3E/
OdGNko5iaJ5Q4lGtDhyfJ2haKIfO1EKWVWR9ATU4xRB2442c1ikyVgGm/3gwo2Vx
98ZdL3p4MmHiIEpT5fktaXuVPKmJUNObRPHGXv4QGL1SKdn0nv8Gy3vtOFDeOQxh
CY9+iTBSfKtR+nGhlERkWdLvggPU8LwYb8cATqdpTNJgRmt+EnY2vCxJPIsLTU9n
NXSD/dt/kVzWBq+fXO/xWTsC0oX03DcOYLwKmNc5rPb2bADkk7XiV1BjvsbN2ymz
anQW5tH7pYaAgGpQSs/NccY/WjdQNNBFILm0rVHdF6s/LPDZ68jBD5B56o57ceIU
Zab/OVihVrCOHjen7OfW65eSLnXPCS6SUEJzeuLn3fY7/UP/GGrbiYtQufsL3cjo
QRIHel4C3fVn10taAM7FlG804f6aln/JIU97gaS6G5yvc+UqlklsD9ixUQzQs+Tq
z9RA4woztcffQIJbN5kJ0DpZP9gCwpc/30i+nmt5bc5r/J8P57iMr0v83WxAVQvl
x2wfjRJZFM87JxtmuCxfbtq7IqDJrhrBXCY7HrrZ8BzvoWdtNAT7Ootxsmq8vnKi
D4E684vmfN93zn010fUMB6no7m9N7/llgSgVGbGOJJvI151VF96gb30xaz8/4j7V
pwlpg3symrO5oPttIOoVypCkXGjjElo+cRqHq1bX5JtAPjtwPwUftOsvcA/+XL4W
JERGF8QO62p6SMSMfgYKXWZaf7UxLzlRxsttu8aerFdfhoEcshQdt8YYonc9a7II
TlKXCMjmyP38Bl3dWlbPVdOOm0rGyg1LCOJRY8evPyUK1Y1K0Xgc4qNq5M3h/jK6
2jOqmpfdm5Lp+59DGiGIyJPquBBu+X4b1ktTi9i1Qx+GNenXWKm8lfG61suBKiJ9
ghy00TrBXIBZAELnRjTFaEOutjQIXZHMixNVHFmCUL0vBwt9oYhBcbZ9KRBBjBPX
UwKzXfu7N2gdHHzXJfYRGSZElsj7UBDyaRdZT4gAh3oui6vHMDGwqSTgUodsJ+Fr
e/VygH4xo4x6+RuJEdSL8AxSPV9nYjW/midoecbt6t9SaZb/yaG525m9xYb8wUH/
5NzXtRefKPh0r7SgLa3cd6aO1HT61j4We50YePfReW+WS3MhrPel2Cv0StU+CWqo
as5gV5QZoGQJjeTpedPXP3A63riMeig+eq3OWQlR9S4yvU1/VZr8cbzuHw/Nbm7k
X62UIo7Xfa+sk+NVewmAMiBDTG6KDlPebpq5PhDOp0hc9WYc6J1gvQOArnplMuXZ
Ocuvkl82n/TjxYlVYexNDFy56b0IBLpTrHnDL4jo3FwTg/Q/peN0jd1gCTMBLpiv
uPmJgS77sv+WHIxEgVyoHO5gg/x1BXXW22g2+OC6uY/67W56ElRiWKGDQ8qA+ujA
vXSB7/xNO3LFtjz79nuSfG526FSgEdqJqwsR67NT6F7iRXIiPuYFqCBXXieTWb48
cBN8Agq4YPz4EoKuTFHdkx+9SccFUBPw9RPQs8qC2GIX411A0xBnN28TAwTI9Vbi
QcycgYRwcvEkPeOCLIzVWTKjHBZEGYYRPGxAnAuZ/G443S05yal3VsLbhxZ3zBID
Ahq/yGu//aFdpgdFVoMgMGgnGLI6xHLKS7vkvVMOPxAUzeSTZDtLOPNGTONbGHPy
9o+R9DwQtB7sMS+MLS04gsxaMDowikxagdkIbWFIVmFPSM6v9X84Oc6IcoNb1vfO
khFI18R+D6Iw73v70+UJadOo1GVcjjqk/GDQotL2rKNt5fl9jUAn2Pp6t/v4wE1L
6caDCqINuetzHAHkeWWZTtOuFDKCo9QDejBy6SmL1DgYA/fYaj1vwmHvhLGWTdxd
50KY24YSbqyMufV5Nk85Z3fYDsZZ5c6Dfv3+Qm/LrxYRFEaLJN4/jzk8/FRtJopP
SdrUtebe5f43IhHaWiIMIqh9WKWYyZ5oxfs+BRQvEr6srgXerbfI9QmYFBdGeZmI
/YtQjbVIwr7CfCN3pktETnElPiWzNZ+p/4Dfn32aZ4GuHxxDmXB82iePTom+tK/m
E1YQ3VUZSB3mvPN8cKaYsJfkwWqYBTAQlo104AjRjtYOr9D+A6GWpZbDIeh5/MPg
Awsz6pEZGOO4/IgiIn4cNRmSvJDZZH3JGU+vaVzAFPFES5Sfh+zV4UT94Ouk8dL8
tNHBRNxkwTelvc9QHP9lurJZQnYOngZbdl3rGsoBXSkG83junik/7/o5y9Dmc1jY
ZFwTyOZeF0oN145gB4RNzV5Fe5azjlxiFWTxgRDmVSgx6Pjhc9ahoe2Qw6hVXZBN
1zgzRVvIq0iSdjPXNAMDXiunMQBMt4eZ/VdTcHr/1OfTo64SOtyCk5EHhgG//fiT
ryXH2CEr1lKldrO+fVdQPHUDjCdetWiq7/jJtBdzDSpZk+UNDMqbjKHsdh9bPfcK
lRxp3hnKBxnl63vYJyX/jw+UbzNaQx+FuJVxO46A/rEY7i2tyT7iyhmDJ+znH7IR
x6tCxZdQu4cp9V6XFcp9CvjeIJHZ9WkG6EGpCHDYsswstschy4Z2QuAVYnZfvPUf
BqWAVod9wTE0bRQc1tY6bcXC0KwK35NN6jJ/IVCoCUBNeA7Ua+QIx0MlAFSfZrVx
EI/eswEYqX11i8ZlNcIH4wkZ67oTFeFk6qwSVHcbqodvcAT2+TwPWH/gllYKUMgx
EVKs/Bgi5LtLt2nnhZFjfQQ15vDjstTHCiHtZID2xK610Pe/BLR6dzXKBgHFUzOP
zbxGrpm+HwhGbfPWFJD6fh776VQlhDlCO4IrfWOOcWMdmJUBUfgYFB2KLhwKIwmU
RZ+geOeaDkxdc86qNx8msuV861ZqIJUrmQEX2hraKPROIaBi4l1a8R1GVyQFImg/
C7u5jKxB2o2AKEFsVd103q17GrgndiPUSyfOUFA5mIHyvvLtI9DiYZYIzxruM0ae
3oCYCy/XSaL61GutQ+TiGILkiF36UMjdFspZzbEgTgF4jO7j8RTXzfZm3kRwwV7j
2sBT94up9CNp9MKJK8ddoTHo4lc9eHL5kCWZb5Td2CF6gWY0b9PNrxPHTE9AYcWp
fH+tvPyxYX75m9FLt1dgz8Goz0V2wT6Brtve8PSpdPnUCi6fbSsBH89qvLpsPrIG
ABmVaXDsHSf7IN1DwhvhcKRisDjVjZDmdAD3csnFvUSplFcpZf8y6DITfRz+FR2E
3C8gzj3XHRk14r+yiySVFzP/mbE52BFfHr1qet4LciEzmiLHr6u9thC1Fv/wowoK
mOEbllHvbCEGLljcEiWbXPu37hfONK33gnAQjOlUm6NkT9A8hUixguMYESUuhggh
wQbRdSQE/hr0CRIeOMPGx9b5Sx74fN4HMAMmL33TKDtDnZik9+LffUnh9XhJabS3
pYM0SS1aLTenLKy1RpgCC+QyB56RF4sOr7VpiJhy2qZM/Ytjs3QiCCHFXBcI6VQa
m2fTE+hps1mVqz18k8XRUDO5N4EKazob+fw8iTBGb3DVNWTeKBb2DyGXnFKSKsNO
iOXKRp3A1ZsmLZ6oNZ3sZpirb/xLgPn4cnQormHGg80lasiJNNWgZGbUFIzCyJ1b
dmnCKQasPvqI6DdRbgB/VTOjQ3wYM5earuVAYM0b3E+yN23rOVbxRiyhZQA4ImyL
lNVXFVso4xIVc14UqsQBkkwB3RUVrtdmLqOPy8oxxiqSituj8kL3MIHx1DdzZo/q
xSDJbIonZ6nA2k86z5X8Cy5DJsiy0Ab1Eniw4GZ3x8LoZ4ht/diFUtMU7poEdnKx
eVVrGRR6KJRlCxOKPRjcKN2OAludita5INC3WHkkzfND+jvaMfgPFpLeXX+jW6GD
yfhXSd1PVfmd8SGNj8XVDXGsMUyD8ABd2778NBig8yUuBzeO7P9X4fSEy9gLR8xN
llqtRw4fbmFKTizpEy0sjZFsE3DcXEM72WwgdI/f2gKDU2+nATic4vu2HQW9P3jR
S1pvUHgbvgpTofLqrP0P+W2tQZoBajinV8ffipBvYrXG/wOg+S76qdA7/flgNh/1
vS5wYoCBA83xBBbpbuiYPAbgYjXkQPSuN3PadtnQTr3VF52+ieq8+RGYOGgwqEXL
qpMylK9RHbauKrzl4g/4R8c/U/UZ55vETHqIiNdkgrxSMEQM1Cz3g4CrwoMBjSnp
Rsrf5C5JNbVE4fnym3ASHcOZv5HkSZCAH8CpO+6giAlQ1eVsD0G3nj7FxDwGQJc0
tLoqJKAzYbntO4eF0Uo44m6tbcz6qi+Kkr6TraDAC9/YouqjWd1HXrH1YDhWdKFL
K4l71tQxj7MHbicWM6vaaDZepgF5N3fTRgGOIUeaEyKyueleXyT6/KwakvhOC3Mk
MHeyM49/Hyq8AxOvLb/83/N6FkUlTIbAB9OuS2ZXMFTvq+iicUxFX2EBMn7+9H6T
DQv4uR4eEhOpaW93gXH2uc6Lb4DKbLWl5bfjeRnsv5CkBGLSJJ11nKmfAAEtocFs
iAnP0gygTCeFWxAj1qLjVJyF6rqKuCmloM/6gt6YSIv603abQCPA8fw0AWaS9VBL
WpJjO3tKnqcToW4Tk5dD70hGVyj+XtyRMFbFflCacIDDS9sn4gb9pSC33BpqKNih
Z8l5z4iEdDuA1lk9o2KxoQfop0WPwWFwooT001GUpAbS62FySP7/mDxkKP71IYkv
NDU0SeJnj2BISxUH8GxcKCO3BqmGqjWFgxTzLp7J18uHdVFa4/5DzLZjeKXoVqlq
mdFe07EJOd5tt6pNs1XdJZ2LG2G4awuJ29ruz3FDpm0SmDuXgsQvdsfWtlqhslXt
P78gyfrH+WT43mPBec4zdYFnWvlceIyPFaLKN7uULszxYuFI/7eZ8nmBtNCuJuJm
e96yqQJJQmxgCethCr4bFXdOyVHIP6IcOyWNMw4M/OWk/iA5gPwlm4UUejI0bYj9
wggOZa1z8dVfYUdRlJVaXkYoAHaDuzFIPSwsIqvRIQyhmfuWGIUvGi/qaQQMw9BU
xlFkc7+Re8RzXSdAEF8h/q/OWmcZpyW8sQS7l5W/HauZ2tbfr5qL3h9a52jlWqiX
03FAttsbZgJyJpwUNlUXHtZxalF7G1jv3OkIG3r3UfjNwarGKHH/bcYyiAjm/NpI
X9jqRc8MP4eThPIyHejua9irM4cgzXZgvtPFn0CugFMBPlT2kiGQ11DfL6/faAoW
GpJRpEuWONYzeI1kH2O+oKET362mipzb07aONTDe18yK2+1Qjimp1FLXLdgdaPQG
uFBc9GbubKBpW5MBsvqIr5GTmdFHEDiiXZh0kl3Q10E1NpV/FPubwJ/9lCQ/2Q1W
aTVv6P0OgEbCZsi6dX45L5D+SmuqNQ5kTZR/1lIomerVNHezEEyfQHhzLMVTtCG2
uRwSVOxRwdOCOcLyVrK4Aeg0nuKQNPjdVECZ1bSDt4CTJfSZSAAmo3oQXzXjqoLL
m2yKcAe9xn653PLAr7s1HDd7Sfd8t1YtGDNySku+rIvXmT/NX9qpziwKDCMsGaZI
HDsp69XM0Bi+0VNq/r425UMveNKCi5u6m8gDlMTYnKB3dJT+087Vt7GaIFTP5qPk
BCNQLqV74w2fs4cRjFdW3jj4u/BR43OQsZoxgWEYeb2IBfFtkX87WUbfssIQ+fn2
eUyNWqboK6UBLRpvh6g18sOABQDDhndmnaV53mZ7yP2yUrmkQ3VSZGGtLQh6iIBX
Qn7jhPnCNurbPYm3JyAQeaN24QpndUtUpGXr/AVqY13TFRbxs38SSreYSIo8F0S4
9o2BPlvcVwSCsrKVF+IWyP/tEsALRVSQ0TTwWkxgpD/jkujjcNuvL89G4vagttRA
oxse7sRs/06lIlG5Gnpn6W6VQSgY22DIgDyDHJSAVansH03Glm9srynueVsk2y1m
RJBrYyHyULGP6MfIOSiJtNC5M5nNnX9s0RZDSXIUbnRKxw+JZHYN6G6b3hpx7ren
pbZtF+IigwVdAWGoRfYxlgj+vqMbHo/AJkWAA1ggV2gq6NMwwcuo5CqLBkiELbiA
h8XMHRxWzH73ieNVaELsbqmN1BM/eDZBcPI4BaBH4wszVs9lZpL2roKNQSnsvJaN
XcXoIG3VjAAOF/9SSmTe1YzB4KU1qaGoYz7MEdhOcwfxBXgklYS2sXKZQ0qbkrFi
h5c1uAHd9FrlVTZTN4SwSqHQdEOHvBOnAlu3+CdhSRY+O7Zt+6JquJftOBcS5Ffm
rPOoIXlI8iK7Q5JDOmjr5mIvfRhWRYjgfreadVl1OKM5YjdUAI28OHdEGZ12uzvY
tvtmhuANJsn6SlORmusFArYTPALhYKXddfYNk7t5r5Xnlwk0AsVESuNOlH9MaMHw
FQO5NzzWQ2MlprYCUeDE3s/ruUXCECflf37tgpT1lkZqaGQcUwRPlVMAoKD/RA2U
o5WTFz0PjjpLSToFNylRr50pLFggo/gUIDHSYeCWwj12N/F9n+MMs1sb49YH+qlv
GOErn8+v4oAmRHLBbGo1Pa0L1gxGmTmlQ9w8OeqY9sZxnyPLWPkRwEn7Kldk3liP
ToO3ORv+dLuNI1n1/i3pu9MaAckeTdLCZKS4rjwRghBN3mOr68B3Me9yE1WZypgY
mYpIscDWu9Rs9+tNnSACIuP6ajXQy/y27u+cEkshamNJ6Ec6zWFixnYnKYdMJQwS
fgGaIBVJO95XQMHo1pJYJhaWedcFQ1adW2cCvUjnjTItS8zPUMNS+ZkQdQMo2s8A
kZFSLyQ9GLiHF940fAAhYTyNc//Ng2an5Rh5XNORxVVZE8Uj/B/wpvSHiS8rLxhs
JFl6sm6y/IUbS4L3CRvLQfnvvZDeU8u2J5h86QtAslMPcmB2RIRBlFAL7ig2XXXm
bgzMXepkk1vcvbHWEZT3uCopMNb+bEM3EnrgfXNeSUIvuOWPKTxV+UIInaoUjeIf
OhgysUdTR3HknIZvYg7W7+dktHozci9KvRxvRs15W93D037QkPnJH3JbBBqlPdUL
d0x6hL+1M10YrQiM2fH+rV1f+uV4soH7rlEe4b6bd6+SOUD5bi0Uysal+Xnf2DrT
TEDG2bVe6fvjGXUjODH3L52QTffR32znspASHYEhTrM+1XECHnwy0ubNCnXxdtK7
+ta1QFT64798xnrotSycJyTMI7KIqkvwcWlCxGhflUmZ0LARKF75tOZIRlb5d6Ba
PI3gJvu56ShDwguoVnhTMAJzL72g7fY8syu0X3a61ud4gpuC3DotwokkJwY1+zcE
gaeppEIaNLg01VMFVQtnCvoLi8bLESXqTjTbfSn4Kt+ZRGbUaiJbSLTEoZ/z3N+w
d3tJxXZzMQpT+1AU919rNEKN+5YbgLu6WO/CalTx9JbAPIlC2ZxAsrUm3v584WVw
lBAQN78J7vRO1LuGDDoLlNxtbrcD/1Z54UMAx7urWdwiTldN0vOlN+WBNHUQBGD1
IVf/UYf3E01INCIHCZ9jhyLT93w52vFshIbLo+wguLIrE+U1Uy1FGnXhDBr3ZbqM
rrmTnvUnPdhevf3nc0EG45fyeUnwSafc7MtgsT15UWSYjn9Je3df6bygPoWm5/Th
72R+alpwUJZm9yIDUdk+znwlaXYxoKZYGCMKck8Le4Pdx+f1jEcZPW7dQvDKCML6
BcbiBM2TT5/yDbx3xYsEMGC6MjcNqQZp9KYpc6uLZ2hpsv/C9qVuZxaxmPmQdWL1
Miw86NduAO1pIGbLp8kps1+gfcGPkLZIl1Bu24fj3skJjFkIHJLzcL6hgWJy6afx
zxO4CYPqUozhe8eSBlQlXHVeP+hAgWXZ4YdxJT5sFSZUPRYRQEHi5qfYoPEUud00
nau8QO2Oa+5T5FFUK7KngHI35IKideqEmc0o/QL1Itbu5CgXK2huEXV36Ro7TGk6
K5SvMIH8kfO7RagZShcS24dFi+ifV+H84/lVV1iq2vQw3VihibEP3lnahUnMONx4
AOOze9YwhoA5x2ieiZ96lqomkKFSgFmfRmZcEi17rs7Zpy/+oeWXuTHbII7KJbs9
JDFduO/8NvNbfYF5emMKMD13x1fv2W4jOlCoCxqVyWNNB/n/KLZBI2sI8leUziSt
G1PjiloDN85kWGPzDJfkFVL472WTkOtARC+GWu5TPNqp7y4HAEgrP4kYcALCr4Da
Fdq+QQUW3ZgKlTLWlQIxPFahPdwycTLAutSulNPf2q+m1akBx8F7RbulU6eCmWt3
TeN0WhOYFdrtBUt77pCMciux1zSXwTzBqC3AIq+oWFOOZ2F4x4SwfsLLq79TWCpO
wtfa8ZNYEMwFRTTgPhWJWXsvgpurcAoGfc2dm2o0WLbgaBpG3yGxCs8k0GdBGjTD
0yToNzItIL76mHFSApvgagoeDiw3yTqgg/3ttJuTJu7FJSKrxQ1mPbT+xncUyvfP
uZhH/KOS3htSfz1pKBmaEZhMc4MZxTT70wQ1BgAGG9rqcGMX08gdLy4K1N5fEN1T
lXgKDkQISZB/EcLJktzDKhbUo2kkeuPznEc5EzrrWYj2wmwFxwgiUChyTMsx57lW
XjKh/MJ154WIdqRE2xEtnOksnFbs6UOTu/h9kj7tMGBsrzPwUZoUeD/AlKO4f0B2
s/Ui2XNjBwvDHScJnZxgwcoawYVtfk8q+f4rzun/srJVK8M/jIygqXX7Yoz6buUy
FkyRsN5p8I7TCts2fzLqMp0ObrAHw7sIMqQOZI//t8Q6kPzM3eMTQz1VTI9GzmdF
Ajt8iWkTra32zn4RUlOa7ApXb0qx7knJnffcARd+DQYanPz1lSVyrZOrmCtzR2Na
WD4iCWrsZT+IXR8JSpNZGTQwadKZzn/8fdEhh0JhjZboeNQTm1DKNoLW628902DO
IzJQgUBophDIirhjU9BuCoj3MJkowgVAUJd0gFlA7O4Te0d7H3Jj+E1+97GmTi4G
V37q/Clnv/7KbGZXjawx6rNhIGxizlky0mmj5SEKDq1BmRR3tXI/h4ffBVfk462A
zk8blmTLSkfkLafxmk1UYn3Fcyi3Cf/2gTZNNXA5AtazHyO9gQAtmC+Hahl7fYj6
fbP0ChX0hAV8WYjsvl1PrFdEDXZupwR0z+BtzwV8KfQNwf0qOm3F2+4iGU9Eoa8o
3aopBVBx4qL5Bo/r2WuvQzw/vp86a0c43fvH/s0A6WJu6CkEhn/K/ODgrzXUavpF
GalLTnNpg90x97A0zHUvwb5dkCmsuGgb3ArnAl77P0bphSXeNpkdGDL+5kk4j3p7
7hiO0h/Z7C9tB0s2dcGQyoKXeH4fecEnE+fS1TIdiIUKX8P0JUkbTwldkvR5UJZS
ikIAG97clkD5BbDuRjYNQyezi+dYntoSQAoRgxxFLRrZ82+JsEfrLXZJgOboSvSS
Wc+CFXi7gw173+ctDWEZK3pVOCo5loM3Nf6Bpa3y3B5GDbTY530ojOVFcohMI2B5
UUg69JPqqiT9ALd2jBeKOliU431KC4msvweKlLGucb9gvT4jwyiF3uDiQG5lIPZ+
Pe/xtW3msP2hV5q8hzkmusDeh/TRkpvBPvD/3lQB04HD870pXiE1H1bo04ue3npA
ITcCvLbQToNPzGEbBrIvyM6DI9MV4pUzKTfog7n7+pKx3HxoXwZT+FoZLfYNryed
/WwYYSeINMeeX5X8S4L6TDteBCsRXsZ0MZ8EIwND5XWviFPAx3lKLxlvTvucD1Jw
bakwPtWq5QF46Wnn+KfQoEQZ3me8U16lehRBMpt1rj7tAFl2oPhdHu5OqmF1U7tQ
3y7LAV25xl6uoLBR7/+XIm6alP8BJLW3xGGKZ8mpIP7LTuOTua+gy5vhBLmirDeZ
mw5iib9j9gyThwRxy4IUTOvl7Soauzg3DCSm8+dhMEF+skGLVvJauH82Hf/pKCXt
+nz1+OORmSk4x/5vzrDr+yth+naM6hb0NxPSv46pLPCQiLoJAjdBeFtPNeR6kUS+
ukMookqEgfCtfjpu8eRsbLfCPcxskAYyYMC3Bqb0hPY9dr9GISdBt72kCGJ/ileH
qRAxFb8Bj9ZXQ/eQXgiBOyioTPT8INPvmFcmBNdpvG+rnkvwoDm4jOfYHOi/70IF
YZpw+ekYpQI3BuSEmH/k8cHWEb+MneyeEj9HRJ8/DYdKmuxJ7p/0ZoriE0+4znuD
hsZh+IEUc24nUFRvQTyX1qxkMhsl6VJIPuQHGod3PG4N1l1CumiU8njnn+/LVtVF
+TKsDskqPSdGghI+S2ImtWUGP0zEbHp3GfrQu2pT6B8t/Ir0P5ueIEHe1OrB9bK7
oGcEOt/EzRERX+5UxvvZ7j/0+q1VTGXfSvkeoWev8dcZD24ZPEY3gRD4dG/Ad9xo
94x2tnQL33AxLxYEy6KI3rWuLLJuEOmy8yelgXTgHGF43TdSKQOka/wqmesAhNnm
fW6O0XcQ4W7vrttJ7Ic3NCSIDhAQ8uZegLWKjVdWG1tkK4JogZmRb/QRXKQYZZla
dnrsHUUFGfQvWSYlhJ7/HQqwaYZCiHhKs8k7Gc9svCWAPjYL2hSJpVrgvXbSP44h
Z+pww8/Kn3cM1NYZxOk7afbHl/wQLO7PZDQa4qB2SA0QqUQ70eceidFJOUXxjFdV
W5ba86Ofo94p8Ojj8x2UWPc64LT4naDQK2c1tUZd5/97OeUTwISRmYmA1ZkW06NN
rj4jyYYJ0FUuCx+g0ZVlZjmx77T1EGcLBuvode/csMhZ+VF03D8YI5MpHBARKp1B
mYv27xRnJ+lWwctYeNFamy7SaghgBoRiG3Xad/2OaHnRzFaXLu3C88pLbIqRajhx
J9WXMOGg+K3l8qvlLpZrnUNR3OMXBdWN5KnCIb7BwG39MjKeVQ4SwGyDSSABGgg+
rsyNiyVPfFPyN/IywD1qnAiY96vfeSWooE8t7a4Ceal3rgBMjaWUy1jroMWsDqLC
vWel892DpKXlIJVitPCn1BrVgVcn93yefqqUVgXURxt0PRWqpCm+THMdB+FpMYLr
WhtoK2hGz75kA+/CJ55KbeHUb4d+z7c8F1hyKg1sqDweUxR8G+zUeE4V3td2JPVS
eEpRdYsARwesh3Hh48O9gsd9Y29eCPI/v4mOKuD/u3a12+43Qy1NBVetO8kbQM7A
kA3cIcn09U2vajkeSZ0d7LDBKXS92f2R6tDe+O0uRnewACkN6L60mVW0t5ChN3gG
gFfrDFihAdvzGg8k0QAdCibd194SIe0vFcIF1/ZGfn68qEpxSCVtj4GzycCkImc0
864RAWJyi+FdYKfp1dhTNl2Is8DxQ+LxBrHo29oQ6mOAz9mj6weCYxxUIDSe0Tfb
Tjilo7xXa472M39A8ce0qGRO3zt1GUGRAM2U61cSMhJRie/zO1DpegFwIl+BQHPP
hEt93HaxfcJkxTZb8iZ8I0H3NSF+HTdKwrR2uuawTzrSHBtljojyZ0VoVlApAhZN
5M1eUwFe5GHxaq0DvFZnr29oEKz1+Xulvcyegw3X4XX6d+z7pOC7E8yUBRuPSeOR
fSp8Lv/vdW7jmDMOrhfqi/ULzoIncQD6bL0OcbAdcP3Y6HuF5pcuDNhncuB/Oz1M
u0IQr9Wx6hffG4JMF4+zkzbXnugA+0SmZwpm8awmk4qliyGEI0jlqx/S7Sa/ARae
aqaHT466xPJqOGKeJ8dzuFioYvJmOpWrCZaoOTQ/JDbz0wzoNqcGOgp+7rDSurun
GPbt5QE6O/jOub4w6T5PuhNtvnzusGB1mLJ44YsVPGDTQF7laOm7DEe9pdI4MBdZ
XxorsgDePgElJfkMveu48Fnyu+rR6EwCQcr+w6BaLd9YtwAAChKZr4A2tkkok0Er
AIR9yJ/917TqcOfed0iGcQDHC4LC+NDIF1lejv37JGw2uGxVfP3a4TxQ7kPPFTp8
mm32Ch/jCcqjlCWaCoq7vekzuLA5fDzyQgwxiHmYyz60dPMqfO217l/NAHMfi1Wu
c2m+zutqxp1qnyWNoms+rXbyAd0qwT5/O5gbyKGHOmiiYl3H2s5XPovC3tHxM/g2
bARUNJ5zhpm7ZMTXzF4AlskVhMXt33BXyHZd64ZkwA7h/0BYm1x+h3aKfNZvsCv/
xsL84XMS6eTRxTHmBR9nmq3ZTBwQbT1dPzXeT5rNW3/cNlo4lC9HTOYuTuQZxV17
0nfZUPD2wvUhCmopkimh7hqUzznSHK0pUljzLl/If5iWl095/V+XqjgFasXZw5iZ
DKAbftrIaXao5PuyHnZ2ht5GpBdCpHN8/fuL6Q/kFnXCbmv4fqEflTZwO5gWaKki
8NdVvwQIv+lxbO7OmwBnZbFsc2WNYoEANdyExeWSKawIobmu3feszWZtox9HEcA6
vmwhBmoRL8o1SrhD02GRWQPzbLRu+cBMUtOm5K4qUPH5nZ+cSuT0MniM0iDBsfy/
d+FAHIGjaI1f056d8Ws6obLBvuNQ9JSg/xlfYjKVKdqs/XYfoQWb7Tql1mVgBrjz
8U3keeKDwQK7bIQ7j3aVaGrax4bX97Pu9VoU56CkcTvjWGgEhYYRWACrzArrjAVp
RssRMexIWl6pB5U7xjkDTl2vUVIvfgxAXMcU+jO8aLOUOpUPQWxge29f/nyZg7/h
KO5LJvvlNUjjLE3urwxcDGnOyQU04RKewZsCzmHFNkggqnV90dOqJqbbF07w3zJj
JA7lueOBUUn6Alh+EhEK8VHKM0c617cbTaHs2azn9ZagWIdKIIpauG6duR6xL1yj
2Id3sCbS/gg/20ZJ81MhA+z5pVGj+ulqByzn3lkVDt8sNOdYWgA6TDT2s/4OYQ3r
nSQd7M4cBQC5+64ugpsMNClhDWYECnWXq0X/5U8ZQmzngThBlZ2snrfPzgfDZv1R
fIBs2mD+NOfJJyhOE90dEHNpvxpdPyNhF+T0Nzs+agIKeeDHHH81SZSWsABesXh5
xt9QIs2H5RteHU09wgRyP5kKMLnDiirMR0z9J//VgHheHiyXW2YX9tRRaL2B2Dqu
TBn1VnHNMJe26dA6kewbRWdRB0ustvlwLzv9sqa/JX4D3V6giD4fHXYQ+zY2bw21
Lg86NUtshULI5/fS/5BLV/XoB08NSxyIbjo4C5W+meO+m6kCjsY57dU8U1v+hNFv
aWenca4dp5her9n27oj5HsHwccgy04eSggSSSK3VZdlLjlpA/NOTPmQHzYovMkQL
eGRzWrTCzIKwRySfryfAcFYZnrJ5M/QNVnYFnPuy+L1j3t9s3lUTfuTs7dtPJubO
8cGarRdQ+3f95wBRyTTWRqFdAfW9xKn6ZfyXSfkvGPF1wIkHzu202j9tlAcnu1Tn
Gk9N+aM/RTe4HeVMH9KGJzxQiq1HlxvdHan2UhNuuL+BTagzOJXe4hYw2bwmGl9o
mKt4TpzQM/uK1d+8l+54ZQMe8eDI1/bKisAUSbqhWw39iRuPlKkPg/9xLqwiD8Ws
gYKeuzD9QJGztbhlQdRpR2Ckl0+1H1cwSCdQvoEPT9idnxOQB2kpMQkahNqsR7/d
1QKMm79uLqUa/wpDsZQn7kE8ho3L79+l65nbApRKwvhtYARq6iydat70mcYGDYNy
UkG4zPoAYYP2vLWhxCm7KBBSufm1xJHAP4jVvRzOW4rcd86+kSl+A8BF3gVQsWRR
Pnbd22dtHK2zFP+kNrngVgqUFRhgTiOZDBZjaAZXe00ss7njlzYF0l6Ip4kyKMQE
2GsEY/QaxAG69DsgtzOeqSRB8vJpPS8fBEVKa8oOBJTG/da7tLiVmoA5pnYmxR5Y
27fNGKmoEkr/GRXBnOlJNA+qd91baQgQMdHRCrSq4vqiYKSsD3ZOIwgTHS+a7Vn6
Fj0As8IMH3DfYmOlh4sgQkUKLUwG5g+MC3Xhoa3+zi17QvvGndW+9qlQn+K81wEu
hgHgHVld/PiO6E5+yMdCHHYw/aLpqIwWHeEHzHp3OiJ/30u5ooN4GrBRieN3vNMB
UJa2vnbzC0VJpSZVh6CC/SzsaOUV/faXxeF5oYlIP3crW/r73rrVqjjZGSKR+YZf
XnzO+odfN/QLgEnw6sJ8xp42Jl5j6N6MT1/m5iTywMiUxYWHEg4sGRq/DdJPJ/kS
xhs1WIAg/T1iQaulR6FQN528OXcyH76fLuZ0tF2FlISQUCwkjBwlvSyaKxRiZK0H
ZrWlq7S+yj/J9gtf2P9wjupubFF/CpVggTgskC2jNJBAej/J+ROykWNBPdZt74Up
TIyJY1bTUy1q6LBVxPdZm5PXE8zEl1b+ECk4oIDmXVz7YWi4Jj4T6KtZhi8O85vq
LbNYllin4svkVynUSuTv15Pw16MUQoGqpL710YWkzLspi3ifbQtgj5aPvVyEUKOT
Hl8cU48gt49kDl9iGYs2PdVfebOrp3T5Mp1j7+yeCDONVxvN88hUc3/vBtX8kly0
KP9Cuf9BlCDriTru6bS7quhCoGvViET3ab/5PawOGwGdQK/41m5vj88ObNL8FSvg
4wMOt3di/KO3zYY8qnDH4QQqkwn/cLjTo8tgiMUTckbMkJzoXE1KB4gwjSztUPS5
jihlmdO09YQ4vv61SeJC+iiEmyjTR3v1ArxNmAuWKZs+47DOEJhTc8kukBxTau2o
7tuKD+TIWeRZrUKMPUlWAA7wmGAheVm4xnLHipSTBD0yJp4OmiKr3B7asQa4Pyku
ct6wRovdn3dNnemHRwIgilxtx0nFRppLAtQDhfSFGt40S7YlTMja4F+kKB1QGgZ8
6gX+odub+Rls+E6J4+P1KOeW7hZ2iQ4A7G11ffIl3bR7+lfqswwwmHSmvGx3kZwJ
jiR1KLfydVSEzP4RJXoYrr/5hyM2L7W0zBDuCQ/BY9GcvM6IvIaQvuuFoyj1xK+U
GHh53UIO9fL0mgfC2CawXEYLpepwic0ce3vyI23J9R3mqQruC8S9vUdl6aEBXOqA
g0AxhAtx7c4M71bW8sseY99KwV9DOlx6f4RgfhrPNy+gL572h0wW9XqvMoLamRwl
nj1hPb5j+Y7ILnC79xpyY77Y9NWo0vQwG00a+n37bOAH217l9nQ+qnAtsnVaDLF9
HOpMtdTAesJe9rU1JenSurX8njsO1Hne2pz2bHg9UPJ4LrWaGxVloAqR7X11WzQl
X4MjMNwgeJVZxXJ8T+MkY5+mUWYyrudj+4GFVkWClHLODjmqzIAmbTLTy9dUOJ19
BRAbE/Q/WR2kEL3s41pHYVAYsnuEFaFj3H7RvFH9gRs6CTI3mWn+EsC7OXFsLaYK
A1oZ2QVu3gGy/YKU8ejyvni4PJqqp0lVmaVXxhfDNaNc089dwRahuhaQ4UwXMQkW
qnkZnlR0Tb1Wh9ZQKC+mt6Z4cDeq5feib6pQnyA0tveW7rGGeqdzVwPFHyalvwTt
EJLMdvTdnkaOKvCvuhHCgn765Ocr3HfCzuC4ei25/FLcUFJ/n++ulMr1myaBPRBs
sTMoGh0JsTDGuOYjjnTwdZarmm0bC2vfAHuDghFH4n+lp+C8XWr3xeDEEVx3vtu2
Vpa5Q5NkDCmocSH0nb5gKjb/rXfGzHvBVjDo1rKDLeUUJ3K5SBMctUlLDaZlmOOY
Y71Ubj+WeBGqRwtZEauxL3+F9aFlYeaQy4MPizIyIHT7ACFlPTn3QQV+bGto5W5L
nJRkxhLt6WQ+opslkDlUZIgWLLVI572//9jJuP2j9jE648OPs+4nhRiKm64/l34r
LkvVnQsxwj8aRY3UClPVfTeaVADoCn+m55rAG0vGXWKBJnQ76aejYldIvbqddxLY
XkNqcSgtYP0BGniBejtLdRt1dDz0H3fxvN4XWPtbU3M2SomB5G/7i3HJMoFk2O2O
196izMlUj/ygq0edoFYDQq1IPWUyJMN6yW/FIou/hUQXgN9ELP5A8x9u5IQGIuY8
HnovF79WUXMz2du2vZnEdHH36xa2txuGB+TilZGqmeLk60hiJvLk8q7LRzxQjC/I
NnWIHxClFNb0xJDpawiGYasd4YBjzQOg9Bx6owCTuaGFzAVM4LVH/+yRGtz0P9Ow
9blVuQHUR0qomPx+YQyKMfeh1IKD4hrfLGTUB5408oiId4gH2UJT2Lg73qVYSMEH
1JsFewBjbEhBeLrEcy6xdEzOJWtIzdfsWqUF/ZpLkcAvtZD8P2D1DynEi3WfkAlX
G/Q0b3pvI9HzFwHLM6dwHwNLNxhkA1QlY8/Qzuav/Y6q8YAZFLlSqql1MpwmHxxE
+dSt5qFWebZ8QPhxh3zzVOssE1TOIallhLTcJIDb/kmUpYuALQtDSkcb/cAmvA8e
EKwG6DuAweY91cLmLxXDW2f1zX7lRZruX/sLA2AlaN8/E8iB/TWFrLBXLsw+xx1x
s6d3Jr0l+S2NNFhv9rbPHzol37VmvhtHMkIejTwfTa5pC8usK0I0webfTWmH6Gn0
1kEM20jRydZxyxC+pCQJ6zYKK1/2yV/sPCT3J9o8flz+5xIbtojxeBrseSAYtKdU
JdRxpBN4xJXud5O1uWumAq2y/lpHcbOQWPvJhj0Bt+MQk4ytkJe8QMwNmqpwV5uk
6qMy4mx2fcQXhT4hFzgt7JhYUR3cP1mvO59MrT/tF3mYK0OmlOILQpwZwOaa+myz
PLv5UVQek1RupNMPaRCPBHgrk1lNnlnVcnVWR0rgf+X1rmny66rN4PapI+d1o2po
wfTzAjADGpbuBjXYt6r+9o/0eIYtslDvI8sujCHTmEKwdUcOvbiZhVsAfZC3h5Si
LybMWwVwMGSQh/IH/qeDpg3OoI4G27msBj9U3VGtK3UDHKX0pSTEFVi1Lbo+3Ceu
fTI0hs36Iu3Xs+20z5F1HnSLcPWtOB7jvc4UNBpqrdLABipNfkZaOj6HmGqxZITT
84y4daqhWeBDD8jMaiai9f0f7hT6tWxgJfoA7gmcKW7JtXXZqYQVcMPLngsKei6j
uAolHCn2B1i1Qr7S6pze3gktncJ61BJl1fvwVYrebCxXlgqgYJoe8NmBlI9Pswal
ACm+RS/lQJhZzsCqiWt1Vd10n90evxLh6fanQMeGwL1K0px758dF3Mdcf41gJ1Uk
Kx8ztjYMHSqOGkat26xb0KLbjmEfs+n8hV+YkMEKL7T5Ty7JUwDqhZhaGL1kH2s+
Otech96kdI0/3ddQ0G2OeEfnlRhZv7ICWWaQT6rHfCKEzPsumEEKD/kry+D//j5a
l5tHKrfSIcuKqjJALVmHoRRfeeaGLJcAlzOkPD+gfBG6kb/oES5LAgHusMj//zAW
1NPL5OL0Vt9hr7XrfOYi6q80/1OtSjgKBCGzw82SkUsBy39I7a/Q4y+z0EWVU+Nm
KMQ9tMgO/7apcP2GQIeS6ceBTySqJOdBLALaexQhymZwaKKN0tbUy1EQx2W/U50P
bOp//jgkH8nI52nwRJ94n9BVeZZwkLatiZz1WX4955F6z/zZrV6mbKJRSrnYXbeE
CMHhLo1M0E2/JLlUtLJPkghPlxsluoEB5GAA3RGIjXrPcCKKBMWyUBRE3YmQu0XD
yp/XmIGQFM2p1NClcuakyJAgNJG4zTFxp/gp3B/5vvLRAeTM9+OrGKqdwcMjOVfC
qJfs+cF5JnOIyLhrJDevQuqlrcsDYY0PycyI1p+0hiQ/IWISbYt6QvElekcqkmAb
0qfYTn17GE5vtSPK3/xo0ujR4AyV48VUn7VI4Cdr3GwspIueNWWkT019/Hi7nBA+
1q7wvVpjy2fUgBBkqWQWORrfevbwFRCdv5E34mNg4T9CrIwcUwyis7peEjfD7PAE
U2+qBzdIKTeeHKonVtZaXomDk9hv7db/O3xCSsaRllmjmd40O6hlqFFrmJ0ugSGe
ytPdbhKvEZwfvF3rmX0DR/rOKW7dccQXRCxgdNQ7jevJzCi2OVU988poj9OpA3tb
sXsHP+5Txo/bNfYw9p/P0R72nysSkgxKHeLG6+kT+Rpc7ccmP102/XI17MooKbOC
3kXKxiThKla1altxqGmuNMUrt2Trcu7AFwJq8S6i+f9IdwVpf+A4SVM01NPsx0Wr
eyRquoEpX21Tn57bRT76NJ7cSSAUof7MG++4Nnf3cHyiozrJlOxOxkJ58dN0ma7V
c9MYj4azYBUByER0Is2lXLa5UMtetqI5u1lh+FqYfHuTuivHF2oKgpVg68dc1uy/
05BoOkCVspeHwVfkva0mIiW3C2AvwkuV4ueHpfe7LDEftP0Y5/4uwzjb/myntqEu
GGNhLbN1wkpmJxomLv1rVZnT9zlbcjNB/8rHVGDDScYffTpJC0nfyp/GwgjA2F6W
7bbDJedtaKzC8/8+UbE8DfCmps0G+yw8lpT2UPFCT8U9i5ai8UxNG1Lstc8z5RRI
mGrzrN1luqed9fJ2/qla2nTT3aXKFASDVr5Z8y70mKaOvsguszO4WIAtAu2ztcbi
T8V40u9Y/dKs+1+IvjFoQSjgYEUu8/4g+KJV9jxIuKtPXL038pOrsA1Fkl9CdERN
rHDWw2gGtK3X2tU82MjUNJpOtZ5091J0zJzCGEqjS11QVkAJv3gs/RPnO02VhWO3
vmgMnDAhD4x/CXFkPTmHLINgrJvlPaCkXakjQQj02qmjilRT81K4T//M48dzlQIk
CREMDfsDmccCZwQqasvEwuTRUZcJYNEjPFDJ1YutE2HttFxqFBhHvYcrHN7ZjvJf
8DdHkybzgkcB13wBwI1RxeFSj1l2KzKGty184VKkRsJjnzkI+HdY6fu/8P6nZ1QV
N+p4EPdcRLbhS2/L/w3DO/qQ0TWdPXRx3Xi1gnkgEpX23jIZJG8shf2VFKplZhkN
MhotGMmpO5b/Mw+KDVMd/J5u7R6CtQtd33NMaoH2bph3/nxRPxxUE6XDcvHPFMQC
qC4WC2wqDMpopZwde5KajS7K0ollzSjPqYgsD2j716iS8ZJYdvmMil0k3TOlpEc6
3dc/4lsyuv9ki2K8pxg5NMSdzDbeLw3QZDmzd6tu0Q0/xMkN1fj78H9WGlYF0kKM
P09NVrTjhOHYQhKlB548ZJNUg7KzCEpOBkyUhW6iLlnBo87bfhZA0yeQ4/9Ucll8
pIToFIF3hgF92KDa+anYnPgUG21NGP4He+ioSB+R2udY1fKN4KCeVgTkHkOzwBVc
zF3Fd1XrmN5ODOhfbRSv0tZMyuRVlLAsagEH7fvhJNJJRDpof+ykORoRueCx7KBI
S6rap56O+IZWuOTaYdSJTtCd1hMARBnTxXHUeWFg8+js7FLlJlvryb+JwJdQ8C6K
67o1ySA7NViHEUO70+fC+WzY9oRVStbansNF0U12cAEn1H13xQ94xO0dYuOfuA49
lHkvR1j0RGhVjZbEFdwFe1L1tKzXCja0r3IIGr2z6NCSSGRT46ahSkdpciPNWqCP
vfxrDLV+d3NKLgi24xgH39maWIEm46+EMkKtqtGdeWF9+REDBwXJCV/uxyRaAC9h
QP5dyYUaqYBvhhtvLjTKVsrhqujYpYWv4GJtbwztJTYWD6u10hgqxsaSF1we4SWS
nKODKxGggJU6FErIoYh+Lxs+216TFt77b9aYgCv5ktm4ggRmF5XjYs/wAA+QUmN6
Dcz5j7VgWcR45ZBx96hYbU2FDokd0qdgwq82jKyJxraL80cvDoxel1SBhIXYf7Cl
G9QIPCJtXXPNexxUQJk/Q3RX1QoYUZ8Bb6pq8YF5FvlDBBXwRSMQJP6KT3nzNzYh
yIBIt1+m5j2ZR0eDIhh5qdhO/1NmId8SFN6ja1EDBq+3m/RUsNA9f4dSILQEaSnf
MM0cH0kcq/Tbpu7ZME3JBPQJyPClwo5oYRZkLj1iT3c04R98ZgVHUHFuTaxJBQfu
eevjOCPEtThzaP4yMJ4lznzcNtuLhjqAeSXCIpMdzfhBQNTxXVEiKIsoacjO4Oyw
OSE6bBnTJeZPYA98wMAc7mqGuxujFm09V9Iwy7iyLkuFprk1d1zkc3F9+sDW7Qlg
ZZoFDYFzULAuQTLIQ8sN87IQgXABtfPmoIzT/0B375nhKDIxZrch9VrLoSsJMSQp
1qKH1jOI4l09lO/5Xnk0QUNgniWO6GSupZOd9pq9v7DdPI1IKhJCuARQe1rt9Ozf
JNPwostLnEjOHpbvn3+O3CmHKi8mWwI977h59KdJq/b7rRMbDU5Hv+3fWIkBMdlC
mYpdKqSTK4kh/uVGJZBN1lj6qL4BYUBBBEYxBI2daS96/d+Lt0E1naHRIH5qOkxV
Y2vHtEpmr3D+D1Y5h28yhbKA7FihwiAFcMhhuYEmeTE2wFGQykPw+0bm74lI9z/F
VNZwGd48C1U0Wglk3yI624NH6OKEvohO05c4Hwbucvd1/wMW8tM5Ah86PCpjALBX
CokN80Q4+CmeyGUhI2AYPyWhval8mUV4uMSgbBRpdRuXhi0xS0mrx5b1rPTuh7r5
PlVPybWapOzxhFSvfS6DIdWkgMMlRVJSMWgMGm/OwyGgV3oG3MXxnp8YgIPsAcgQ
FcuG91HEbg6HyOSDlW58lwiaNqU8KGtKugt/if8ineMi/7jBhUqJR7envrmr9/5w
tnWk1diQEl7/1HT8j7dIyiymsTJrt06eb6u9UZ7JLIZKweASTGtnh0biC1HPPwWI
8TvveNd11bW4enPEgRWsBA2UrgDsi/oxqS8Ye7JGWaQvuOmRkzA0Yqsk1JihZspg
EJfQl7ltKqF5BCnhrVIe9CyksDyTKPLZfO4u0AJgL5xTaPZIZz2/A1Dlr5Quy7/W
QifhO4quxrGi22Df+zmAWPU4CAYkExjj5R8JbS4x5Q62Jqw+XOjniHElEWZiVOi4
faeEEqzYnj+3h3Mcxa0adfqurBGFLaYuvc2tXvzvdS5vrv4FFWZAUb1w2p+YFeFJ
PqzEWcOEqayNTjsNWpsoPzgRKoEEa2XXAAOBXzswYbo+uKLy/VA/IVVtSF5WupQM
+/SIjrk9PHuiSD3j41xAYwTOCNpAH8dqjdG8HXX+1+I6zoef6bVVD0izc421cIGi
2UYRRkARj13WbaXXQDCseVGd4p2Fzu+SJcuZgO0ICBCTvSEEZQS6L8DgBt80ITk7
UcReBb25XkL1Deq3r2nW/z6Ng2iRusNuEFSJcY4FJplnX0aIum9xvy/SKBhWc6oZ
Dgrtx9foNHAYWNFumpTiQBUA1uSe97Py4hkG3upRNCZOXq796ITYx6mS21vPPP79
41sBaNBRO7uTf0sM/vkl7tjVTghrwd/de339KWhx/nsSBJaEV34j+MAZh/X3S+dU
ml9ga+24DtdLtzKD0ucxeujPTdzUoO1sZgViLV17fHMLxmM+CtgzI9Q5uait1x4T
NWA1fJgRhIek4JFB4f6dH5ROTijsa5Lp4jIFsTntN0dK3p6egsPT5ZLSlZUYv0rq
hX6VfXrBX95l2OdleurDpgFXPVFfKRlTdD3c4P4Ooktt/Dlf5e381uOHYUcGge4S
aEYNiEK/vMVTdy0ugfFd8RUnGwsi2J8fmp4E9/REgWcOLB7h19ddOpmQXkINR3SI
GtLxPZE6LVlGannxkt1JnRd3XqOOTaTuuknBZr6hA0FbAUN+4FfNUTh5HIs6mC2k
Z7J/9zyRMWSysqV1UW0USphUvZ0xnHSwJF8FuekHD/25MBfq1ufdmZcZDx5jK2aa
FwJ8cbVZ3a+4DdJYqb4c5yC+b5WPlqIMlzzJnsbOu7l2u/InWg+dDynfIwubGYUy
ZUUcFX5m9O8liRvTyqbl/Ex6ppwdL209wDaBpNAAAB1v8r6B1R7zjExRBIRe0Q0B
g8Zj+WsBHr94Pj7EDeqEf9ZwjsmwQVzYZiuoYNEDVyZkjFk5LxPbmu6DSShhQuWF
G5WS2uKTodQ9myWd94NfNBfuv//2OQ0b8XpLGeDf0kC8hzq9/XMebXUJj0JVeXye
3tRfxFkM1yovbjaR9LfSWFj68suUzzsN9jfEBCvumkTZjz5mbZ5sQR8nO1eMDq5a
2v7PnQAQ9IQyuf6HtRRx763Xv5L+nqV1MTJolz/OooUx6dpQrrQTbiov8ywN4eO6
f30PvhkmqibB4eRGUiUk5sPdnT8dd6J2KbKpEN1/Qod55+D3k2nBYFIr8+EboFmI
825BDcDrj+BrdBlQmDfoPFm7i1TY9B+W4hkUz1D7Cgo8da3TY2dB/ZeMhMZEs8St
8wQh2yQa1pkYWSJFFuwmCo5sIfYp6ySeYKRQWJF2VU5ggxlHnbB0WEfOpGXX10z5
nFBZEGrUNa2+jb65SIb7vUxYuDaSj8ZmbMfekQzTCYwohDbRfmw/rflz/JpdGNwC
yHFitL6UuuKFe79ut8AEY4HCfzGdAiD/2/bugC4+gWnMnmzvjNB3pJSVcYtl0KTK
W6NYPoDSelaMiXE4nnZDZmP/iTRoswmQv0UtmeLy59/Hs9HT4wOMAR9Az26N6RPx
WcvkmcJuMCRHjbUQvgtxtpjWcvA+91P0OTcHi0+QRd+jx4A1wL9R2RalNj0UfDwI
x6H+AcImvguYYJ/jQYgDp8vDUzBUGf2Oj9hXNhr1aeCSQPzV24lxWAOMeSEw+Lb2
6JPYx8diQhMALdEkpSf5MtQo15eA0UVHfpb6QGASN8QWsrtY9v9lieRYVuZXCwbx
nVh8uVrkWGCX7AbB/Wvgn2cIXrkrP0mSpIBUhxmSqTsrtIaQKZi2svY3JTzwn188
BZzfzVMBfd9R/Hs3ZesBiYRagpx0NJmv0JuYfAm4XyMelLLshgse5f/STwJsfOlQ
t+MIqvyP77U13pscHi1ZRTenF+1JCqH+tz7HoyXW5QZPrCuYtulheA9lhR/XFCpA
Y+IamxxWJYj75i4UJoBr1QVRdjPncrd4Bpt3fYH5e93ylvhKx+xO+8tZrqowwN1O
asm1FutXUlPar+P75AR+euMWgGGL02lXgMg8600kzvJw31rYgP5l/5ld5X/6Jb1u
leoUlRUTAkUM3+OZ8atBaaF8gxPzRhMi0zgGeQsgzp/PiXTgwbjHEnim87RedReo
5NfOEESKKJL8J/u2r/OEj9bfshTnlsgdQ8BvJItSMIHXePD+fa3JcnOuqihJ6/vD
l4HSdTzPEWJV/dsmurLi18CmtzUPDxr+tWxCq4FNdGrdag8kqT6zdMdsqtSPIwZX
NTODCjdqxRASgf+YzQpBLu1plM7oJv08hlbxXkBe2Y10MMkJ1BX3ASsNQn+b0inM
+pZ/tq0Urb+I54Kde1F2ZoFJgJyuMszhdpdDyuLh4EQnMYiVyLCymzgWgr+cUJ8Z
X0Z2wS+3K4LzEl/XW0gMaBmqNAWskyId66PtJtpZdpBRkYbgqf8rkZ4kBPRZR3F5
KzhEt5i14yy5AG1u8t/MxFGq4Wu4sG2aHcRSF+6OxlQuVy6N+XE/dwEOrywcY90g
bd2wDE3EjpyzrWu9kGRvUw0WHjkuEI7hqqce7wpG5aUS6+iSwv3Au3WuqkJlgA2o
RBms9QWOMhW/btjuI4RiX6aNP3jBfwNxJ7QP7PP91MA+KyZ5nLu6SPfzQeCbbhSO
8T+WFYGuVsGWrczzJQu77gUSy+Gjea3IiD6k4dmDEDKRvSrNifCaSRUzYfj67hTN
ZQGvlWaJGJw3BF4DN/bS0FDn5zqD7fww0M86RdFtKeTqNURMQsDLsORgdCn4Votd
ZXIv2cleLi8PDrpSczywkeOPHaeBA43vFso7i6fK2I75mqtecm0rDim0K014uPpQ
QgTF/k6lZ7CuJqXRiFT0B/ynK2Q1MZchbHKkjPQqydZhxHeJT8gBprF1B0gAcG/a
OROuuxR34e+fEyRRHlNY+SjLfrccRdrizeAYcVBEPh/ajUEmuH0c1HX1hqsL5/Je
J1GuW9x2NWpl7JGQyKzvHY/AGKxB2xKFROB7bzmkKgg9Nanxl3LueiRcBrmyv1yH
Yvo/Arrmafau59InIvWc11b3PiG0KHuD+gPLYWU3d4j8DzrREcF91VK/WOaEXaDv
et4Mgh6GPQRpfuZsBCCABmR6QBI3fSIvOSb+Smh1Y3T/ez5qWWnwcJTIRfr6MiI4
Wn4Gi0YiEfWpswJOP/3IJ2VbYpsKfawznASb1bKDPVif9voQN1NUokss3H9lr9RD
y9u/2xzLbINEXtgDXGEK7WRrcgF0VdL44IoKEfzWu8bsfhpXJKDKg2e8Sw0eIGHk
Kt6W8k/itePi6E2kqvQd9675pchMVOAreC7KdeEgJzn01iTK1c/5PSVG3Cv4/wSA
vNrE4JFOdDmeYbNOQwA6sOGLt4Y0dRGSv/O9TDr991s5Pi5Vj28Z6Ygvx6vm5DCQ
Jq30hJQhwbs56D2jkCGSiQy/q1rvP/ZaYKp7dWK59n8AVyuaxIutE+9CfNqMHUWo
sjyxBfJ2yMkZHsCVMQDeZxRBA+Ht5LwJty0+a+auH87OtxvRwNB7/OM56iQ8raif
VpCCYdz21S58n8Ltl2xd2+zjcx+eWt/Z+tuKJ3lruv9RuJJih3y3gjQe6F7tWIn7
8VtTjKHTN0qNEwgGON4MZ3oI6lVMHcfh7KCDQMUP0M4K0yJCJ/VpnfNIEeEWhjFa
I0ZzYzemH9hgaZSkZar7tqFW6CF2RBwAdH1lTcTxmd6QukU4tEpu3Cxn0spNZcIH
xGlTZCgdOheXbrNuDvprglBrcYT7wAmP02xcVClhvQhSfPMTFhXtFPTvIjRiktGP
3XZG0dFHV7Be1kRupvh/U+sOnvhZXdqNVYG5z52zHwp3T1Rnux5BCCflbZF+0xKQ
b7SDPj5VNvp7Px2tC3rNq5DsuJns2Sh+8IFc401Vp/bHdrbwz+Yf0gTjsoOoPUVp
mVmqm/amJg1bPpkq0AtfsCUmo7dtWDgIoAjAXUhqKXXEAXYsoorigsLCXUdl8Tka
ik1ZUQQUWJdMrf+3/dlVs4K43B8hQi9znU03HJoF267xmZwbZLcVoNhOG7UPO20m
GcEDeF6kqYZQ1jVFd9v7E6bDY/JC2TC8wlUmRXOZpD+RHvXEoNyis3kU1paUbe/H
42ax4xW5ahAHlRq4SiVb7ILHYv7vUfeOM8EgHiOj66i94T3jy1kB/vIjP9j6mV2N
T96OyaFBdXJgmO5ha2rzc98sxsbSQivwmjUNLij668TvEcvAGdHrGvV2SAaJQLUt
KHsdgA/FldmJjinWox9xJs+3CTHozUASLep3SQVQ7NG6KPf/s9vfL1hHl/5geS7B
EKmWkBO6tR4qrQkANPRmWhbeLEvooGDdWp0X1JFrEv+bgyIfS+TOwX5IPPwqUC6M
o0oVSoR/tn1iOlUGWI/loagpWHX3hWeJ3OkjzFgGtnN+S5aEP6HRJ9DR2SO5Wt04
6LXLamJiqebv4tme6Q2g5eFDQ0ARTW39aKHdu/d5oIV6M744/Tm8cYudwaV3lUtM
LH8dahSUCylj1t3O+o+vpV795ovhum/cQQkHO90m6adBGZ484A+AYX9O3+1n4GTr
6yD+le1XgRgKvNEBD2FjxsrEXIAvsXmrjfsPTyLaq5fJogDf1pCd2IYoFIj90L+W
5Gphu1m++/bycl0seJCz11BJisbflsn2eWgDXeLIumw0YJKJJwXAZnnZg6wrOXFM
oZjRXPwMJ521YKP/2odjXywPmjqTz/GHiOZRYGuX+pRCoYhaB+23BgRcsSWKoit3
3vgwEaqTrCb1Otcy6Ws0fPWGWbDnPiBPPzL2BpYuJZdA6jLggaliVGS6+tJKwIBw
C1+lvmK2z0yOEf8oHj+R9lRKVHBUMvsry7cnTkqnxcXAj/rJ8wKMyLL5XS1Zw4eP
OCuXApPewW8F6YOw56/G8YKfjLhhescRoOzciIgrmaNVK+6bhnlZQVdWwlJQE2qI
61yXgt94SjDJ6jJp0bbfw2uWXIFrXZu/i6Ke00yfEBIMrhHAHj3hLy6gfi8aMR0H
f4ex+807TJAcmQXz0X8zxVU/GA3E+uZf1csBXMzk/jqF21F3K1c0PrPv9csvHHow
7QbxE5Yd87tmoy+9AHtapf0USilpRTQiZiERjro4jgcAzOwFtFJ2y2NND2z7+G+H
VNqD9LilPEa5biJV2hj8RK+d+FCzTp7Eh9meFQbDjwqYoYM8U3uAQuAJ613YE+uC
sfKviSUqfq9A897lmoF/ZJjZGdRqzbea4C92gwpI5/QH3VkUF1TVpb6AMu5afXhL
Io/COrer/PBPZMHkWSjNWqmB7PwdyoHsyuQrECDJewp6BTuBGhYcmXm1/6y/HQip
v0w4R2EKg1ywkRHlOXS16rIk6wtsgN1vBnsIfoBiIhvaVf+SKxfJKFVibZGJ+ACe
B1jZYwaIjo13w3z8Yiw++0obVBvmtMM9LHM2Pb+MlZqMwgEGdIASwRaNOIn0rJgD
LkF3dAgwjE4hJ7INuB0BIGSMbYXSsbDyEp9C8oUW/a67VBNqnS0pbYtFs9/rgUXS
k6ndMQtL29kz+PGKs7HxIv8JNe6JKQVvHRbYQxiIhn6Zgv3KR1r7jUtyxWf9gAwn
u4JUHkQx+iDLWtQJVWlG73i1hHbyZ1B5kCCTWohGNi35LA6SqcFOJqT4GKhz9Bnz
FfC/zNw2vekHH6PrnVrN43lRBft9XG8s6Ig0u5tQtKXWHRe8dmWklbfZlUDNj8pz
lNrvBLc+2DPr9h/mm7jXVPFplyJwal+1+iX2hZWMgE7KkUjMuIQHHZWMBHx4AQdV
IS8DGhXAOFSzNTGs4V/89w9wBh2Gkur/KLOCcL21L1CksnS64UPnQh+tDIofxb5G
reYfttWs4Rhee7v58RtQa21EEMQK8B402226JMZ1mqJI0FKZ5bZ3ta4LBn2BqpSC
++OKENbn3EhycBzg/+4V0r6TzH90i2Gl2lJ0YmMxupfTYc+xjprORJHkA9D9r+Ov
I9dYR74+T3peRKU+tET443d5xxUaEOBWcvrlmyMAl1isgwjtvOBQRQciy6pdb8iC
uNKhzJf6Fhwlmd3Z5tMK8Gs4jExFpslu7qcUgp4hzBYLyE5jLesB/GRjDGvvdC1J
Tvyyj1W4g4Q9X7qBtrpoKm4CyA3uU42W0DKBTdTnG51iXXgTCv3TqlTuc7pM4CRb
I73zkg4/YLdIsfcQL9aLA692XCqj+YlTayf+NzsSeDYshAQ43MRKlL7C9CQMfKz5
JkyYlUNOQIg+OuZHX2J/uqyFYkwsQ6IBB45FicoMVpaA4Ouhlyw54nHZD7/KBM9c
T1UaLNooBAxFYa8FMjj5Ec0c2X6TlncZYcs9YQtfbooUsoOAtiNXel52T5fn+fVn
PDgpjSoaX+Uov+Ed0I7lyjyGZkojl5fIRCg8IRw+vMePBESRh/tuUad48qySPpH6
YBomLpq/4I4zYmqAsk1nRqXLhNjViQGj0fAusGYomLcuo4xlaefkdKQ2+6SlPYkU
qi1RexTS3DM8IM7zjzTRq6xnPS3CWENTXvGzKuCHsaA/8yxTU1ha2XVJTmzIQjoR
fFJk9Zk88Kt6gGS/V483kCc6Iq8NKwmi2x2j/QLRKIuBsImhFFCjgd8BVNYg+XhI
cE6zd27789lxVjPQ5iqYLTmGfLZwwSK3mk9IFUmA3zITwXnJE1u3C6Lg/sjsZVBG
J2NNFgb8ZuuDad3u0Zuhll39G3VKCMv+VWyYMHqb45bYhzynOZec4JDsBueiF7YA
eKejqsSaGiUWu0A68X4KWBmK91s0m2W77KOWv8RmsbZxs/DqFW/dNo/xSnfhlglc
MvLzP1z6jUkbFzK8UJPlrknqIE3VkqsauX5yQiyPVllNbeydpzhPjHKXaaLZXYF0
JwIFRu9dKeGnTxVjG0ADd5asgjwo7AF0vqxamjCP6YRWX2f+XuiUzqvatNM2sxYn
Wxmh90Mc5JhS7N4CM8QfDhvizS4W02bGeZPYO6BK3gHVD54eddnI+xADQ4rc5TR1
njI5ppuABvmvK5UQB15Z0PEvRBq2X1f4kzORukcCs+kPURE++0jLiD1K5up1SseF
67RbAB/vegniWkAoqA5XA2dDQlasZFAilk2agoLPSuk7MnlfMvbDMKU1yBFIxyV/
w92xT6UZc4pUqTth+UrJHym+tZGJl5wX7Zsu4TbDK20Xs6Eb27TUcJfL5dPClwY4
RL7INInCKXGc1IF+KYXtW+DcVrngmQDlWie7NOiQ6pvJv+MOezxuD+rJsjAuw9sZ
UQofYiTeW+K+C50i+D7zhGfdn8TZvya65srjNVjqQLOD/NQZgwnSY+g1Nzq+jeNm
NainIyGZmjOaYngvtN553ZJJmQs2fI8Zc7UNst7HIPGrIvu2CNpKAi96DspJu5XX
iIY0wvRPyrge/IiZIVia/CeuiZ6uJb2yqP+X8cxLTfOhh+ugqXroV6jWVFBIvOeH
9OeH7WbhOUSeJ2qy7eOobClbwc8GPVwzOUNoKjpVdviDzhBsZTi/9GJDWgej34K5
AJ8wkeS3TudixSlSBE3EPVS8+tKLsn2EW9qaNEJINmnt065uU1XXO29xMvPtuRek
umRQuCtS+XFC657LvFzm5N3GAaeh0t5gOBtEhZB2cD6k0FFoT9aAW6G/HLFj2Z9U
7W2EH+I5KXkoYvKabrQKWUzTVEm4CpDfm4dscMRG0Fbs/8247GUWoum7MQ/2x2/N
8bmL4mvHRHiCVOMt6mgG+gmj587Pkw5oEgIOCvivt0Vwoz7RRM+W6fkYu2IkWR2I
g21eA1GGEJfxpMwxJKg8XpsgoiQ2i2l01Pv/AGvEjtRSjaOfCtSiC5ZL43f3r9fK
Zvy8FRI0lK4XavNl8IAWbkWMD7Hjmw5e627VRFiGvdaOaOERfshjxJto5pG6FUU1
1hwX5L7dHM0tZfCQ/sGdmQOI4iS89PwdjHbpVs4oF0zrfdsLE56n+BBJrYKdanmx
dJqAriagax5VnZPt+PKlQs+1N1yTNwqmpHCDrJsmTyWyOZdeEVAtZwEpKz5Z4DDV
MuHK3uQAgtT/gJxcwZnatXwKsO1wdgzdJbHznwtSdT6KvFrwYGHXkDtGFSzWI1PE
rgGoPMm7WMtLhrFYApaXdLbvr5Cl2TrV6RZ8a6aoLLjrEAoXoZVqpw1asIGaEss3
N+aZCEb09RBwWnfUZKzgLRwojBbILNytCfZUQ8fqbD98kOodNTv5HedVlyK2inC/
4+azs8FMBm408U3aNRzm5fPkKcQLkyUjp9C8w2rYZDpDJ92CYl4SQixZsk8aL86H
DsSwNIxcMPVcNQ9P9IyFO4MLkrIct/x0BQyFdqTPheDh/wLbN/cw9o4VDoE4CZSN
ZAl4yvcQlT9M0Z435WHCxNvbBEF2QttDY+PirqJUM8I/TncvEw8QbGs4xDeEynx3
IcFeYJLhSdSbvErt6NABdnxp3oHZg8RbuPfqanMbAEBa6hnQCyjhr6B79O0XHwi+
AV+ah3EnfsNo7xX0lLerzwAE8GOflW1sjJC+kAUbcjDn3BOGiG+SjeiSCssPKdhF
zCwXpRfdVk4g2dZp1Enzt8AWaKAoF+hJGjkYTkLhlIlS5GmnRSRITQcv0osCVMxn
z1df947ZIZ5Zt5Ja2yHEpeXKS2kRN0sKesq5H+0CKCuwDo5zzizmIzXlFqNNb3Dt
gd4eFvvzcPCfvK26fR2jzRP+IAygK4FzVTDLqQZVEurURLdU9mPIgD6m2ExX6le5
s6rvKj6gMYX1sNH6tCOn/VrFu+kjOY1AciCPdueTJWGuesbU3fplHlsJ98loRl1n
UMHzlEEbQJDJ00zQloy3Jm9mwTgUfDJmHW3BZo9KWhlHT0tgj/WuxpZ8JFgStxN/
9kHNWZ5OcsPopfbC9J6yuHzA4cWZTpDLslcM5K1trmDCYLT0raYcGrjKF/CMy+zL
JxJqhYEo4KUON/vs988DIePgaDtGf982cpv+K/U0OVDI1aaU+Z6MgVbsoryKh+4j
Qtzq5LRePF6hIyduJaBRzg88D4lO5moww7MXzETf9GXioBP8Ywngk1IWcXV5Uvbt
KI3/npPLlA/ZDlSjz9QkM9mG7mL3svPeNj0c3jl2+PQ19cn/KDkWvtbPcaARZPpM
sNZo/Oq5xSpXVcgLav3rbh4h2jxVv4WwRd5GvQb6RuSrZ2Z90QI8qCp8S9WjaSzq
8GlS2wKFwH758KPm1T1OQ6Wks75BN/4tMCRmIztznYvR6c/Wk5kMWiS5OrWmISD2
vAAx1y08gocBljedkgkDrolKA+JkwTbw0IA6+cxCsLAzqMQCOj/FEOiknWtd9Klt
k7anR7L+xZSynTB1He6V2w6omwchef1gS0Fa7Nfq8ANfaHiyUSbgnwH4xZgw5cjv
gSQ2pPIlacNOWrDFNuic+yRkJYDPvpogoZd/qrujZvxdmQdTaxjIJuFn/a8itNrR
Jsc29J8uWyNcC5Futp4sOgSowEjgnqulSHndjM3uEIOh4Ux+KCEEF9NWgDQPO/94
KBsUCU3riP5ubSIQfhQdGXSvFKoLTlGdDBWNr3JY5HIN0fQbt31oJgrqiF+cxdXL
doLsOZJGs5hT9H+RuZHmc/4P+c9C+2ZsMhuDxqEsWtEW1HVbvEhUAvKpMXZ9c2dT
pBltuiiqYOkEG8lVwci0x/mFPejpP9iHjiSN5xxM2QRiowJCmXpPF/cZBm0az9GN
SGau4NeyPRJdXCTeDyaglI0cD7wsJzFHmXtu5aQExR1pa2Zb0GRJy4YhxVNTS7Xn
lsgWjog4XvYDQxOVJnHnVytJVZd4PnngDZUTfHst3NOFc5SzJ/mm7CzBAVlvpAsr
5ofqrJNt2+TJd4qFVh+pIdPhGxg07jVlgDbQpVy6wID14dk08eCKANLnqNxqNt+b
Vqsf2DX5MKq2jbm05Uz9oO7JhNrzY0F1wYfLXzDjnoZad+v+eRgGBwR0Zj+w5f46
NGyi1qIOeqVH2tUfl5EaEHTQcq/HzDmD9At1ABXORNbQzDZXcLK5/mVMcciqq170
irxzU0DSiXmMauNCCC5gMWQsCRmL9KBV+8qSf0mPlbntUXJwzbo0f+QHiw8BR7V+
XR5iCtNGbK5fZcWqWFVfC30QKuSEinptYqVLln8n6dUfCk2l6KxSIeKEYq5nRhOH
PsFaHE/wY/FVuUrn/TOGpA07rIFpnZW0TzhHqY4+3iGRp38oOwx33lUv7UzxDRDr
6XSzYu29GwqhBYbz+e0xyeOqA3sR/+oTkBdf8WZQ6NOBS2DtnwDWWkZ9UatXUXoO
2QTX1Xkq9Fhb2bs7Q5LEPdjgyKQmA4Z33OHfWXvjUnmCJHXkZsZO+4qmfoDylAMS
ZPgMVujLPNSqSrHEoGKSnF++2nJMN+GSw/4cJPOJiuLJudatagowRRi5TzZNiArj
+r3YasGZJAb8uQS1c7UU9qitr8iixaMyaqTUhGSPBj5ClsL8a/ztnelkahXd+eOG
xYD+8aeqBP4OMlaeVmsej4E9rd/uqqBTOA8fJCmsiRhNtyMn5aL3+fa+XXm7qViy
DSeCgLdoopMZZ+Phy5zfEokEyuNcqyOoINv7kYt39F61hqb6v0k++gYfs0bvttU1
MDy5IuuFh+1CUfO4oIhr1ra5YtnAVMIihbRRWBa39V7D5K3ZLvmCzeq7SwURr0zJ
cuPBDyrrstBJ1G/s9iDHPj2wzkv2JpH9SebozATgQ8tYBgB6N/8zQCO7hYxTXHl/
Gu0nIqJ5v7gtjIKhDrLTV7Ye+B7T8ZiN6uYpYJF/WLEp+g1nk2FvFF1MRkHcnvPP
Lsw/9d+Ja7UgHMkaH38PqSoDvJpvFUCS8455BCk6s6+M5j87kUTTCiw7LlFGOWMD
FzUEeqXRzrUJX7ipdSrhKoSCMfUTMM4KWabClmcdc1rAUmJs3j46xMY2o/d/LgNe
rvCGyVyE9zk7Tm1FJEKkb/aZ4uzFXPZCmJtx8BwO0j5FddsWusgnV1vJ8j79fLOA
GhLzseoprclwn/PZjkcTO1ZzeBGyzq8iO3wnbw4XyPTO3enl6+nD09/WymrO/tsp
a6DvwDBW2GUDtEXhQEhszE1Sfo/LSpMHbNdCVYxvOeSxW6LOo3wLZNzu6w6aPm12
kuY56TNbMDUNK20YBU7J822KjO5VGNjQwhYIu+LJbIv9yIjj6Oy08guByKgRGYpi
qpMatqxbue1BPricTHwVk9bLNSrTas/jOhmFHJDNfBNVbcwm40WqsQKaQKewmOp4
t68XTD8MTWk125sERl1scpz4rVtlle4gHmSMpbPJYIvtD2ZbSWLXMdto0NYLuncl
XVUWUk9BOy+FcAyQkrg674XurYnw5qNQEe0w3Y+FYL47yw/0TmHY41vm7rWPa2cX
vzQThz5x4tlYswSSD0nNQ365JTFqXwOpkwfIyCd5bwX0DdDlJR0UoJ22C3JpTg3V
5uxfMmVS31YJHea5wDnLBs7IERsxNw0+6tBEQcMq3tE7p8IkkzUPCKUfCEVmDyYF
vmdvx2H2f8erc1oiNsDFEJSGu7R0Z2veqH2j9FbSTEdo7biJLtsJTOV3UthdomAy
k2FRNf4+hN2gLPT7Eln/LAHuVxLKeoenTJ/FQAzMEUugZ2l5v7sBopwydqP/KKqe
uVrh8PDl0C1Q3v/go7H3gMzEz0x4aPv7VEyCe/adfYIYapMFlTjoGPzYo3Xu1CmP
kg18UR3OoYIPjxnIHdSAqXibe7AbowezzQHZ68secfSCZpbnRQi+evbnCkCoGnNK
9uBgmsd2NWn7dKVcaeJRXYvi5L1Ah9gNzTP0Sc6HdvXDsE3DlsLC3CfOYfbw4WYD
silBJ+pkG6CxtNFpgutAekjwBuvHdL56wOH2X5LD0kM3y/82IeO0D5Ki0yV8KNPm
jZALOGC+xEgbwm7ULNO2AB7+VqkIolfNznz6u98Fjc66NBAK2Yjl1y5z3HHScTAT
iO3pX8uKtR9NRA2bU0hG+wK7zz21TWBg2xkkYAcD18xmpFuZVzpwGVnZafdL0whG
RWMUVPE3sT8fl/5lEadad+MXnAvA7s+vyb8bqF8N0DrdTbl7SccaZVewEwfAno5X
1ZAq1h2RTDyFoFqxkJaXiRl9xUIZgQIu2t0x+yU+Cofcgw+YRWFle/DrTZdu4LxK
d0nC13O0pSSQmEATZebSqGlJxSUl4RuIEJiQ3l6E0eCyBrr52zsPbeikXdn+HAIh
aTZZsH/Zw9q+2xvOVHK5w0Y92XlsSHFwJj0L02qP+2ZNkYttoPu7DvipqfSNfJ1I
PdVrLapkQPzZ6iWPeHmrqMWBwcd6BrmIO7uwUb+6KkATro8Wj+RMW57A6KFEXltv
e9TisvGztSOyUVqJOFPD0q6SK+tDrOJaHWV3sSOboajujIfmtNCGtJEdEirqxKRU
lWMEH4LjSAyTl0Hnf36mDJBtIXbFx5wOHKMejyho9erzWc6N2nU/ZYnVvtVM8SNg
8t8tm0X4wsuAsm5kVMi5+eT718UzjmEwGHw1csr+qjID1BjSbiVOqav+TXmsJjNg
zznMZ2qCxDo4PXknV3My2mRCfpcI8uWLkB7JZBbN4FACpKkFHxP29xiiT84EH+sy
hxz71DE759Ab7DNR/Dz7XFmzp64JEHkT/9/APzG4eUJrmP79akkjSf1gIKQHAlWP
lDxVs9lBdlUGsEYMmis+7qRUpeFEbVwlQRV1lVjw1p+XwJFjesAyzjGwxuSHe2/f
PRTbEo4vTvWEb7tsCdeWbkmzqs6Qn6Sef+CKWln9ffcoOGUy+lkOy1z3QA9uNKyh
yf1iqTW6bWX1mBMuIKpjsRLpqwVnqB2ieY5ZdZERuCAVOKk6NktIsA+1MWcKf/Gi
y4Wp+tOA6DZ2ZUoVM5G5oMX+YdQvqX0PD15jfIspXjCn+I7RoVlDxjneD9SYJ1cH
kUuFelayCChhB+Wax7gRjF5+c47Bq80zCwS85ww6Pu0hZKpwH1h+d1fy91Wl2ZL5
R+nz5EwiITcyDCXwpy9JUSd05mMkhFxtSYSmMxhE1XNeSO0qRyr+geRpyDF7MZgd
sLD4vQFrNVxQH6p/WoplxlbvO4XW9zuI09b5b797EkgLpxZNx4QQZxJd6sIbrnrD
hF0h0TiS9CrZqJShS8Zu9+OdlkLmRtJt/6m4yy2KtlBL8Uggz4RunLZHTcBImttz
IgaLjKNFOVQ6VXV/HpocG7DT4szC7Dxk8Nm2qU5VNF8dlFwA0iBhJgQLY6xbap0b
XhvSezCmi1gbTQbbUGKBDxK/wLa51y1zYBwj5kPu3+t7mP6rG4XjuGDNto3I/qBP
7qub10UeFXcjWZhmJrrtK2KdexckY2ttMxtq3XeB9BQZwJfS3SBktQEb8vrBbjYl
Q891IvqTsMfxOZprs8p4N9bW191tExlC5gdYVkr35Wxl4Kl1HZT2J32rQ18Oq+Os
FSsNssCU8ox6AwitTUg8zNr9KQQHF359BCIewVPb+c3fNN3cXDOF2QwdvqRNpGIt
QwVPMcv4p4F8Q1647koeKAMalfw5PCwXMh5ETkPDZsITvh8YmcWFx+zPoMq8QtSU
VczKyN0OMLd0ZA8bmjnbiBC2qJf3hv4wugacjxo7w8I+aemb68EwIkKY5HhZKuvB
+LJI6e1hdSkkbtRxstSnjaiXCV1ijYUcdc15W9ieE29HtFDAZ8YIrdnJekPwZLjz
R0//u6JqpC1znrQ6UdPAcklHMIivwy3gL31F9NR9BrLpN6Swn11/UyK+zQ7Si8+k
ivrrXfSL3K2l9Ft/a9GF8W6786NqHsocL7YoQ6H4JixenjQTrNRpfachqxx6uod0
2XiF62xLL2+feFV7xLq6c5S5JR44mIJKC/oPnOsGqXRhuVlRadyHFlAR0o81YHO1
EqC5ac7yA+15iBaSrNATS2u9AA/rGydShiNQciu9G8LlrhuHXQ427M7WS80xSVBz
mhGhFBGZLSXr6icCAp6oGuIs6nxe0Ks2I2f5WlxcgfLww4zF2GI9Tje5HNPUdU07
pep5bqoHNvlxylm/s29PpiNfZiyMOPbQkuOZ8GWI2HDor5wtHneel6DlVu1cYspo
uEUeYYVwLqXMWWT36L+EVybun5LWfaG+O14Q67ssRrgHNBGDI+xIBrllkbaeN7Jc
T/6nkmg3tfLE6Q9V0ZYHduydk5iMXk+CXoWmiTZeBd8K0O9Dfw+7ag76or7H6JqH
Id+6gwxp2DdaHdh8eNTs+VcvGOXVsK4/ICgMq7J4CmGFiSZavnKNM1HZDLs0mweE
fwemjkQG76yUgO58hEjvFDT3q4hk2hP6fm+jf2U0SNCUjDnDl6nMkD9fzFOuAtYp
+EclcpTaAdb9D6ipOWkXKF9+9itYxfvUDySXTU3j41I012gpmeR9eBhxvT/1Zt76
MpvC2nLEkbpI3kX+qYYPB2myYj2p+UfpzOWRuPMr/gs/FD91JxOUhuKyLnHqkMRu
T0IAS87DJTLGAz3vaW+uDtFbrVoG5xo6vBGwM03IgQoZSoXQkXPsgNonvExNnrq3
dgJkYnp2EDyuc+lsarYCaD9+dZVEt1A/UQZDfkAKuhr63hkIhWiSDFWrli4zcY03
gT/y1NduCBU053l3TkPo81kibBVkDr8aalRHMe41QBGLw/xqa2DARu6UzJt41JRm
J+RLAqD9RCiT1artLgnlmQH/UaAbkb3xy4O3IvZQ8pBub7cyviG4TrWe5lqmzFwt
gfhv+l4k9O6gBWvoPNH89pmB7t31ef9Hv6d1H4DTzbuPlvRNscuWIHFqYvHhn6eX
b++vIztxg4iPLkWr0CoS5GTGlL/rRm1zjH6lfxP3cVDDqJIgg1ToMgBytniyXXCS
EV5AVjNzY3WqvGiFbhFYCBuQt5OwHndcItL4GxVQzvIGsmTqsO7C/ntWyD2t69HT
4W1rXvS+SQp/K74efpZCaYhWK/wvfHCP8kGzrzXuPvlSDXmEsFR8ZnWyqyOUHpFW
bQU94oMxPzE/VPwsOagOFPdqbD0DuB/56PE6wrIMESnDWCwt14wlcY0aTFC3gRyn
sj7iNMtiArApP4wVcw2Mvnp+wNiu3aZGq1/wU4JmlVSEpfxnDXopHvj9ooZjUKRP
fv7TyiA0uL0LTJ8F/1W1TeQ2gV/YU1ToLtshMStBnkZ731DZSeZ+lb51wZzAWiPt
Ybk2t6yWqb4XNQjtwlJtoLMq/JQRlLuQUxRNx7pZKn4FO/FDlBXBBKQ0odo9Rnmd
ImB5PSztnbFcdzEWMVs8YLI/EMeHA2ZDc6UTUcoBKgbR4DVTTagw7ubwDaTLdc8Y
RDzsmVoPc+60AjZZ6GXjT5SUpDjNL4xAvWxJUxFRhlAoL0cVTztbi8bQnirCfxTI
bIP4rS24yKB526VUx+C+GsbEFHqA2R5y+9HbEMEf8kO3GQhxKShV47TBoU1Uc2om
zAIBOC/6CGBhBzHCv2zL4mGarZhKG0xTkw0f7IwFOOK02lp4B9xDySRfGJtVn4+W
aR7+M3UeEVx1nZ2AyCbp7risBcFo+rgEXw1ocUpJg6lSEdiYSyY7+sXDxqKpaRJS
GbL3Gm+9dHuWH4gkp5sUMA3IKrcQ6bHBnw5vVXjc69STwmtC0HdMfGOaXmBzUYuR
nB7x4YakfmRCXgBNuLLFVjH3Dbjz1BnWa6bbw6pI0i9BSzYS8qI88zdBOfi/24I3
df4344bWzV5D3YXBAnvS9JNqxptp5rrJxewytrMTGthDKHtNQOPSrTmER8Ll9gKv
wWomRl3hZbSpNj6dJPxpos/unFJ2djv7CDafT9Rb3js9igBOnOc+IpvrIYlqvipw
zUzNB//noR0rrWo5CK/tFGQIjVCQt1s8qjaiPkLLotSWcGiT7tBEif17dRr5taX9
OOakhU2M1Zd3q46LjQTO5mkwskR30H6c6x16ZKSHOpgbaSD52+az+Dfx9tgFK79f
xhnXVjG7meruQjKbcBJdYUK6hW7zLTfhyZ3XtdjyxF+HntRWYHpOn+9t56Y7eOk/
NqNZaIAV8XvAXZ0LUnCwja2AG1XhLqtE+aPOFYWbGFFIQJIBUaEUnap+s3cc6tEu
phM3CL23p30vZpqrPZKfWOEDvKLL99O6HTQsAVOSMrMGKSVgbyQ2eZ48SN991b8H
5/9epV5cqaKgKl2cNiZfbeD1NfWfHu1246YvMPaFOSMQqDyC5/4qow5bXIKVOq97
IEwXP5/z4/ocEpQuW5suU+a7ug5/fz2etgExNQ9E51Gt4ycTpcPyoDM/wLkAECgQ
nZvwGtE+O+DebnPSQaNksz6XtShez4mKvrqhfRsxK5b26CgOrh+dOFJOzDQtcUh/
ESFqOmVnBfkfTiaC92DP8MuZND6wo3iVCWB/68WLdND8aSHMWj/r0dDTO4s0KV91
lnkNC3GC87pPipuLSbd76ZTNg+y88gI4qdPQ+eOqcvU+TnQwd91QyOIgLxdKIgwd
xF6XAMeMB6RHCzOhAyjD9jPvbJhEQ2Znpwnm+CsBx40su1KeXfRcnpl6qm4PJfuK
Rs3Mg3Hvycn7OF6GusX9H7U5To+XyCXfzDa8J/XWbSbjr3oYe6lwQgvkzf8Trged
Kf7tZHEShvA7hkkdwZpevarlxrBQeM+AZjbL/P4WiXP2yc4YBYDzV1qHubJeb5xu
KWPbSB89UajjDmovl0DzMrqCSEYFroC6O3xqK8yG4AV7WkigPSTnhaYjGvDWYnnk
BhyO4iDUGayxpl75XCp7OcuyrlfIJ15EAESxt3YEbK+hcic3BvkaWLrno49OxZje
BCYanjGoA00WpEABbtodvEK49l0evisPHmh15PYfq0YCi/SVl9ai4O6H/Ldpm6e9
Vwohu+pFuOrm6k0kxHEApf2ZHS5w9xo0YAjHN3kwaZ986MDEoVXugud+0wDKxhUM
D7EUowYLN2OYzhdB1rGyuLwRIlgGmdA2YjFy7POxE1C5iQOH1aNKyMapn/C8vQnD
Nn+CxAe6fnvZ3Q2ARq3Yi4hjM+iIHVdY/oZ1P51nYfr0m6wETPchePQ5g/mIUs/s
c6d6VJliVhYHuJmjbhR1ev4flShn9M7nx3yZFb0aoaERtnZENSFpc9VGmM/TxRVD
5/25GWZ6hjj2nDynQ8e5L3R6s8A0NgvUJT5TFrySyfxMoo7WPp0JldZCBnSncj9x
E5zM62O0wU7Xju1KdvcNdXM3PaCmGCOrmys0qnqGTIkx1v3EcSvnvM2Q71PDGA+1
OwI6grS6dDCJTFA1JJYAqc5eGx7TpDyEIWK4tq6cve6LmaoNGvaShMhim3T0eqe1
VjpIlR/awEgdMRqmiM/xrNL2LJn70xoUzBubt5eFS8fja8y49nQeyOLbSatIC0wn
8lXHJjMC3a6+6Kd5bpMSZJudVXVfKJbVroOpcW9PdFqJesjuuHI6f3Dh9gbKGgKr
moA2kmPU6/mjqwAjzVPuvBK6bcyc4cIaSBDSACyjVvdi5raSIfh2y3HpcxNCc6pF
VCBScOFOSjlFY/wjpLCwSZMss1f5TOaJSYC0Z+6B1aadIi3TWmbpiP5tefHpqfMg
GQW7+zopRA+zl+dN467/zBDWjupFmfzBG0pIulyv9XIc8TY/beJxx4pZVPJkqzqZ
otpl5EZe4YTw6Xpbp9MjJGxUTPjSrJA+hV2AE5Puo9EVnr1Eaz65JtADSR/GSOOm
DTdKM0pb5o1VdMYqWEuzzZIdNzA57tWQSF4+tL/NDwCvSWexh5KcyTpQ/CNOUPA6
WoKnHh/BKlbJ23Caf5LqVsaXshx7NAHq9h+M34/VP4GM6BAr4dNMgCAwD9u9XFzT
Opu0+FZ9ryq7CX9IfQEqsBvW3WHuqxB/FAcorSUgJQahRg6KISXGEifIGzf7ILHE
WXC9MvXpnGQUVXPjHKi2FKIIhSKV4mHCVqdupgvsNwMfXL0nZhxdxYAEKVtuCP7b
6GN3sPBE9s3sLpW8XtiRXJBqTUPHdKGoPO33Pl1yFtPhzlDiJ/pOILKh/XAzOTAd
f0uFg7wDGU4flxaOpPfgXO3OSYhNfU/MuNux1GHjFilt56pS8ZoX+TSmJSJlft3s
QKjY+gmtxXuxqa8asaNPaaCVoXEdyhR8WVMPr4AvvKHJJj4bxL+C9ZTdMiFccu6s
Ava5iBWIQbuh1kUgGMi82DB58u8x9sEF6k5z4hUVp3EVYQQBeuFGP79bHorsGSFy
qSq3CxrGOHzZKjE/9FpNBtIw8jYujK2OTHFkUZnhrh3G4hRSOoJaDu0hXftTvNVK
wSzm4m7CiWrcd24P/RROpvCBAu6fmfFMviw+TGUQPg+qeOtMF8/cKA9F9CpR4eMz
eAAgMyDMEM1xwiKSORXFR7OmEPbJ5HP3xPwyAXBp6erQPTT5BR+pyj8R7/pJLAvz
/ziCQ09uwwDv4cVuEqMQgGwvjADU+h43qbGnwjROgiGDRXNj2XjsfInGM0b4OGpg
B5g19G99VlNRo7cbikXjVDizJcGIWYCXo8yBBCKdUGzBvgO3rDLCO8B+t1tZaNHU
l7gR0vWuxlkJ9qm4vG2jLNTloVKl4PQUhxAQygHc9xKHuVA/kOVAC9e2wpMK6mdK
8UxvuNbXriocuw5JcwIpFRSz/C+i4JqJyjwm73ENWZOyzNfQq5jDWkV4567vsVIa
ankSM5OEaJwlY4Qqpvpn0fm9vq4HS5HzMCBHg84u/Zpu5Y/dEDI9Zu3OiduFcPlh
lJWY6vEIk+UEH9RWEtC/sMovx/dvR+RTigFf8UVrrIyWaZMp75puLJW5XuWWltk2
nY3rgGzBeqq2bp1gIb3b6kwW8lq1M5nXbb9lssxfEswqMdt53jMuTJjJyd4bfYAj
EG9sJXrCpgHJCjI+D37VCaPTLbvxrQU0meLKZ8pjl9mwhOiNAEsDhVRzmC1PNyeD
JisWuIY+HgpP4gsgV8ToBwQ2E+xfw42TdgQPK86nxsi2DKZzi3itojjjbSXN2VRZ
5ROo3/qDRXu+stPVL+fW5niTyrZZUBIigDJI3copv3yiXgbqkiiJMeEp39wwkTZ0
Yz7IE6fCM7xQAnctg0sAc/lWxRUYQvAbZ2ocKTdYUZU5VhAQ6rMHiEzS4dQ//19n
65Aw6vfHwE2oOmQ2KjGW2kEq3rGXcnqxZndgGtY7TddlJPk3ZWC9A0oQ7LvZoyuk
iiG+w18zOXFJTDNc5owEqpeXnxPgEtFXP/2TNKSFtd68hdiogLQvZ2aYhRc2L9Xj
vmcKvxHw3P1NGym8ihWVl+vS7yqp8RPrHYxdQ6wmG0fNsGBU6NdUTVf/VygbPDRe
QidoLdE2Qqbo2NeeBoWpAilCebP9Skr/nIy288njmT8d214K/ANN3dbnHIHjI0Wk
j47NE/3j/Jy1b/otpCZ7uxjieOAGokLzyNpE/i6MvmvO2RStcQe+ixY9Q3K013hk
BR8Gwt0G6TE6pXeGFOYyjhJpYSaecgE8tMqow2g8515Qf9950/KEqb39kJYc1xnn
zgb75YZUtDUM7+ZX11TcuUGNQABQEtI6wYu3MwmDsAmllET+ZifWn356GuVnuAqY
LPU0hCPQX7aLWc5C0DlDZjRDjYp266W+GiIcRh0bb08J7gJricYySb8aJvQRBTVM
WjBSd2o1YK4uGkw7e7AVhLALJ9pn/5YFSs1HT3mSlwnqaRO3fuPIWUuXtoKdnsYZ
MCGh5LRRKfcVfGZDHpI1RRfHwor0botSRfBu5M/Mi0Pgz01YlogngTlQ/4J3EHGD
V2hF3ueJjNntBgc2W0m3R65Bv/9zUoWvMDaUhwPAZB9tvZh1BZo0cijbHVvmV2hS
r5D0rcBPhANmmPudXW17bmodaYoDneYc3qmy/3+Lui4R+1VtEpCtfigQyVYuMqM4
gaRKxfvmhOIMexe3tmcecbeYYsw7RZ+Nf37uUwihRdK3HDxbsmO/K/id65DIeQIz
8mGlNWTvHCQhTuu3mjT4D+MZCdrxedl+S+XR+fOJ8hJ2t3PxJkYp8VDIfNaKViYT
4Rzngkd8Vg9bZb5BO/CipFoMZQM73kvCeO69cOg0R+6IVmQ6PIhTeu/ZF+Jkt0or
GgfyFIIlTDh8he5UcEnfqcz7YfNk8jfNSFu+s2zVqCpKegxRdhAggTEGZ4QsOx8m
XAKnOQP5LTJKEML18pn+lR2HFv7GWJkstGWVydQocT+SdAAaTCCu+7jCUF/LTEsU
B6u64EZ4tHBHDaWkWDwBu9g8lkvzGxPx6TEDs/1fk9D6qP73Km29x7VH0IJD9xbA
pz0h60L4cZ6913N/BbedbUoSFIpoYw2jjv7DqrDwNT0O21CMWBaS75CE24WCdooI
I2JjJlezLai2FF1S1HQ83xJs6KXFoHPVHkvmBGEztvOhIn6ZtH67+wZZtxk9/702
6OER2Z6S7lZdUaFMK0Z6JAn2uC1KwA58iPfiuAYJWc6GgXWerCx9feGXPrlG7E/M
4MbZYCVXxQ72E7RTHJ4xy4/3AJ4uxvzMEFv7zPx4hAb9PcalzF/M5HWI/Mmfd6S4
XZyUwr2WosqP3eC8wjogUUc20GL3SKh9028KcvdI47xQB38GTsYvW2y2pbkziZdo
+H25XTv5DDL6nzgk4jkOSdPRa0xdvD0WN4xkkLJR4B1aP3OxywSPO3IMly/fxK3e
WgcVQeW/9Ol40H2l834KPKvl03Ag7jOAB5koeygmpSGY+Z4Mmyfq4Fjx5zYXnDwp
ET/U3w5cd2CueiGhUDUaulS+Hp3EMR2njsj8SX9Cwk5CYVKJRmgltOtzQrQwtQ8W
mvDe9JUaqt84FJdvPq1N/IDbOBHJ1UiJMkOG2UFbC9q6NQa5fNkOu9Oy9KLF43Yt
2TXJJyK+PLb6BsywJ2FkVFuJMZuTvPpBl8f9LPIdFuG1rzrNax166mTp3vhF9kos
vvS+d3Jbk9T+CD1d/komQoELjiUCL3Jepklwp7lEhT6IG8L33YH5hrliUsbSsCEQ
gzu4/Lis+3vLxuXXgXv0PEsi1mDZPh6Syo3tzlm3xoO4U9YN88hUtHYso8CJCcpM
F5R8lrWeLfyqgVulNmDiiildZOl5ibagBZR3rxt9o0P1+w0Gi/BSzp/WGa16Tyfe
pFyk5KWZbrsO5eVQl4ui0cI0F7ATwyacUqk6PoGBLVMmXrfI3yW5csfCXmnaswlo
ZFTF0JRtNwf98AdUV2pczWynDEcYTrYXdMvsYlp/blT8PGt8y++jf4ub+lltltih
bB5I0gyWrlTQmAGwM/C7pWXl4Ycn6/iYpSajKvgTktM12HkUaF6FIpEYS+6U+qTm
sAgnJwBOT2yf16XVxAdnOXFCjwhfx1wgIuUGwRk/s7WMwD87eb8kJC3o4sLzA5qj
30dP4bL+d21qAr9NtJD1B5NM+Ajh+2Jix15jKZqOUCn/jfI9d7q3qi8oUszUHA89
y1P8g3UBLXg3V3eGdlP0/pnJ7Q47Y8ZKnsNlJfntbeZ3BHC/GnJbBwdoDagrs6D/
sUyNrbagp6v2nxSMlG4fpgtahHJgZLrzcBYBUmox0mq6zqbeK2Lt9akmykjWdobb
h7ztaK/wWaW0m1FZK+U9BgmYEgwoVV67d1i/lkArqMgfCto/FTRhxQVDqFnREkOa
RGphi8hZv8tj/BpCrsm6bbZs4vsferlNzw/PYzxBX33pQLGMzrwRQwjCWQBR3hkz
BDNBrC/ttzFES+Knwl1HdflAPe5eB+I0cyKEInEsBOc/bOn7BIJOeXXBJ6L4kDpe
HxR0+8FZCDELO0SBW+sN2bfI6LlOjShMyqVKw6ltFaHFkZniig9O5LubRxIo3wbX
i0WBj3KK77OmgkUijIBeV5Kquuh2sxCizKRaLvHHPVAHR5amKPfTI1+t8c5HlEvG
8BOfl2Oa3N8boOU7mEhE/f9oNDLjIXAvspqfwQbECtzBxfxhaqAwYfRn82F+8bZ3
XC2PXhdoHm6ennU/IogFMgELm98/UADoMEHJe7oTo5mSyGGgtFDi8juIfwDYxUJL
AOtDTAVwcQmdVgwaZs9gHWjCgwUCT30zdZKUVaO9T7wS0qVC6m9b4mr8sPYMT9/L
1u1Wv+LeucNx+sZBkDG8H1hJgq2TzC6y4gMlAnBebrJwaFZqmbDJzg2BVyuPMRJP
zxyyzIiRWzBS62kdLZaOzYesi2oAiD6hz4wsLki4RmDGRgRSG/j9NpKYIB6TOhVS
QZZcsAM6kfTr4IPjREcaR2RpI8UEHA5MEopugyQguggj8eoOKq41aOCc6HN98pwC
T2MnMRBbkfmrgLU+97yctXVbENKgCsA7ovVuNJSSaEDW455XBet3j4rMuVCqxOuP
QPpzSh+ZZqCKbo+0OvYVq+ZtOWDKZgo4Q0QoUiagXUg5Uige28NqipN526mNMEC7
vvzfl1frUJsdE7MTHujznrrFVqTPAtFJvngd+f8tyx4lSDWvdPwC3Kks14FV67Q5
hd3oIP3bXH5Wjpo9ND6uIJCT3U6U315kz2udgAvQHl5HFJHG6k/AP5oFTYb1GKby
xXxzyVqD/RhaV2sW67JQy3biPKcu2/IpMw8kui/vvZmU705EGEwvktmy7zExswIb
v83jZuklf32u6vQvKF36JlFcJzr4PwGap87UzSrk1Mp+emv74r39UQSvoUzsuJEX
rGF+l4KrbwY2ML+DzePqAOPtJkCLxddBdvxXmUNPVSR7bnhFQDFk/IrGkitCNHWC
fmz2HNgImB/GGMAxFv2eCc0N0G+cHzCmCuiSaMvxlde49Km+DkUnv/h7TXeeiIko
QpaQELJKapOu6Jpl8qIBUitT5qi5ayIpR1R1Y1Qs+9JeuNTJkg3y3zJtPH0yLOkQ
c8zPznZbP6B8tBK6cbVzY5CRjSs5s2bUEX6Sidwbt7fy/5zzRys8YY+6pY/r/tbO
G1pX/mSmKmFl8rH93h1UKq4V7fs5IAPWb5Ia6oBavr92RSN22E8lGuhD4dGL8r93
dzBlD0010/aXVzFxlNOiwQHZKiG/ineiygVgKAmZrggAo1oqjaDx3KM3C7NQjUYq
kIZ32sxhlolo5+0Kw9Zn4Deh5CMtaYba4x7FTPzc/UQxoUNsrTeAwYhIuXzI2pbk
L2zsgfY353gWVRSAuUSfpmmQcRY+HlewLZLRfN4oEByI8Zhw7BqY4tx2tTvl/3aD
v6mFS/rEmLt+0WF6g2C+Ygf5WvwPq6K4QGCS+eZvh5MbOXy6bXt03GRQxhuWm0/E
0N31jCkUvicRI3n/c2m2okFUqzTLlH3lU6CoBY0xK6AX4Kzy2rbI+2e0XTukXW+Z
9Vd/jHQohIMJgYP/3zm++BZYt405a4E48ni7YgT4plDZvcdU0bRDk5SedpHP4ij6
ggy2Z/Ijc8fsFS4Bpe7sgR4mZnEXshexzkjGhzzMxS1Cbi2kDorvNJBSV/ZZdOsU
C7TiSpLPpyonTQpwrI6msLuG8TvA09Lnaosg747+euA8m5YUdgSa6fUyKBXQ/NeH
fxew85Jzf0keksNI4tDRtHlfgvP//8FLsXWa3INVGIE2n9/CFnZU12prV3EIYdN5
XXmVg/N8ox1G8zUtWhRQ7ulBg+6Km5pQ31Nb6O5Dg+RrBpO6FX/b/DkTgSI3a1JF
hUEtIQ9+YUGsxIJ8H86tgDu+qmUM6F6adtjdhGvOq3W1XG0hayvDHq8Kti9mqgIA
h/VwfdJRhTohFQIYqfF2Jd6PfuKsoYZonSbYGKWWrBhd5tHTFGShTxdCNXmrClAZ
AkBH15XFGvjEk4PBBLyJVEuus58wbN7El4GMtDmMfbZkivG2TZ0Q8D/oYVJPZjh/
nUEeCjKjK3amFs5xam1ZVjCEzja0HzcfJMA0tbiNCW4+REXqM9SRzYCHtPzEmmNG
THBb0GSY1q7sknCfbMOC5knMCaDwGr9svvxjzWn0elYdELRC6nPw/0kgVuVybrQz
6XTbUJ4wtHFh3MTSKecDosdN5F5JrgvsrFWmU4t92ytJcS4vqGugBsvFj/V1FDsr
LRyso2urvgN/6qPH9J3s2h6Nhezxcnakcs6XpHn5C7CAkFyOuxLkj0o6Z78m1YRI
kLNmSbBkVKeEBRZHQyDSwK7o02YHF+gcNgMzVjnQLW9w8zEq72LJ5nvP9M3RfE3Q
+gPKgP7xuPgEkf9Unp7dAIQrSey27sMB3n8bMtBuIiqk4NmwEwzugVWXUchdc6Bi
WC9xRMc43cdqLmPdJ3pm7dM0VY5e/FP9ti/4kkTJm+JF8qBCEQM3pT1wMvkqvOhB
uzbi2CBxt3G7P/qeJrcoQHA39LLKHzoP/gXGhcydTMjQ7+/yNGX44/Z1Cq04DY4F
glk+fN1pzGC4J+g2pzGaMKZKMwnf9pOVEogAYtebsWsDSZ5Z1elJFwVrEDLLfvUa
+9OTrUkQMyibhbpjQXYg+EVU63/dXoE9sLmrP4D4SbBoOPAYtPyz/QJCPrwkB4+d
Z69LmtwLa+f8EMU0ZDWP06FAi3Op9jlOoElmVMvGQ4plsqWJj+hH6xOdNHC9DpLh
nIec9rpkDrZPPzqcdrYQNs5ypNVMcJcNGJCsf1dg7eYx1FYr9Olk/xheM9C+4y1u
7XVGyJgg81g28VSNzI6i6TyFnKeew8Ehcu5qfQFgSQBbEHPYw5mf4n+aRcy/nsea
fQjVlhvwl/HmyrAJKR7cZzvlT2KazNXMYc4ob/UTnne7UdIeZhdjNzo+Yx7vh1p6
E/qPoEgrRGWESqLnXU7y1Tq4IgSkkoxN0dfjShQ0H+ooKknqCFaDsiMozVW/ia6V
+Ytq5UlI0Yjw+svNrgKiTTMEnIoNuq5L153E22I1xxBO/tYTqfOXWH99zCh0X139
LLDGUlD2ehrr17xjWjVh0EGt1ZSBmNJomeiKJwnrntHqFoQ8tnqndIkdkf4Y6+UQ
9/2Ago+K064REG1ue+iDCcm3yGf1Mn07MM8wvSxgUvUsGqXebiURPwywsFV8bkPK
rI8eHJUWxmHeA9452AvFde/sq/Tss1aoFx2FbCMEUcEKhSYXNHBdxElrXd3jKO24
AUw8zvO+0mxJe8GmxBjNLSIYco2vVbcsDqVR2gtT6IPYndgNODyrJRJG4l5qmGYV
FilgGBu9GWVCvRUpnAuNBwTDKlBbSto6fn5hi1wSDX1mvFYplEvpS62VqGbgszKx
iUbdQjV7orEPNbHjD/v/eDlhMyr1eCLA6LXZwu+4gdFDz9VlnGOmhQcoc2waAXq0
MthkX5n/3eaC7usJ+eABSXfF41o3mtQ8IQ8wQcVYBMDAR0nKAZLMjy5GDogpUQ4l
JIN2tf/cGNWcYJYbJpA5CK56jHGBy1GiuO8h1Qm7PPWX+cB9mRpS2sfh54UDoo2X
bSB4G85ksN2jhuJu98NSOGcbeQNvtmDaAMZ5r/ePiurdB8V8J7MGfWAOcqEwq6jP
1RjbZ91PvkBrHTxLXnvLRn1uaO4mKgLK3jgF0sLMSxVlZjBRsc0wNo7Wdqzk0pmk
pwObMZrJzHmg2yFijmjsX5OQVRXsTgJnQvZOF775NrqgHHxBbBBUH7mktnsbcUEk
jkBa4yNBpeuHKpPG/tMWYqQJW6e/A+lGVb1pnVJi1ETGQuD4uhy/NCRqPHFMX9wq
daL/BOUHwN7Dn8P/2fKIdfU6GFZsIZnQ5RDa/NGNKAjgFj8KxMC7OgJpQtIrgXcK
i7k3F/sgzQMBNzz5owwidsdy5bFW9jKUBB9MJY448+PxjRH2C9Lkg3bSMxIWVLzj
+Puq4xC3tlSSXFr2pQAleLPIxn3/5LvVYeV8JaBMfdPp2sM0BLlvD5XK4PJBwHM2
IFpN7+ppEpagCXkQIO4G3Y79Sb7jGeGST/Zkxekqnl1TguuUw2wpv7oi747nQ+8a
XQidVC9Ct8VM7l9MEtndjqUBixkrX3wVVMQT1l6NCtG2IVCp2eO8Nb50iV99TK64
p1Z8q57W97sFIJ7Fq0M1IxzmVPp35Zx5mCZQx5rH/9mnWecduVTORKw2UqeLMdV3
2SUW4zGw4bvfO46bBrkYEFbPvOV78PqneIJCJaqlzHSpC/B6h4978O324ELRoYuR
Vnvvm71YA3YE4OYzcqc0SiBgb+tKpdOFy24XGQL1rCi5R7lN7jUyVKd6ujWVNCCe
3zjaXX/QZlmAnvzYL0Pwh/bRg8FTkFHcOyJKgPwWIwGHCTljgoo1HO3y0fJ+xE1g
GaAeDe4N60cCsau0pNSzrEsWqiLwF9RDCo4wHleGdUmuEJMoUtd4/kv+zLbbPCfR
a2l167KxEgcC5PR0z9GzdIPGiNYUhiZ9bRpyqLyrNa8ddzJkr/6sqeTrS4rQOInc
6h5f28G7PnLb3znnrJa3Xz8BzgaZXUIT+HqsT/utWrcq2CBh39GM1Go9TQXSLyn9
dYOE5q9tT4E7b6GrECk+drFStVq2HWbt+HkWuoAuAV8X0WgOGdJvyUaCtt62FB1w
FXicuKOjOhs724RymtL+6EUyxTwg8zRxGh0Vf2kvsJ1BNFDoi9KVie+3FBGeOOqN
D1FHv6/L0kJF7N61tvsPJg0YoI1/+CnJgWVXkQIQOkBPm3xrGrSLYIgvs4q3Tjra
1euT5Uc1ZcwgP35KX9QRcXM2aOu1M1gFZlDlYd6Gik0X6szq+qIiWEXmCwg66+7G
x0yTWPZ+IpRaQ2PN78ZKVgSTU0/A5Fg6++GyfqhRR1unv4joxWfGUQlRz3JFRQwe
r8dvUAB/oMDs5K0B5rMmhkBSmLkUXjIDl9o7YeEFVbhVpP7P5VObbIRrWUdMNRwp
seArteiVlTR1qFMCDukcOy4hY98M36ZnevAF8zFUR5sTMGNitGAuTwYPTp5wLxid
vPCaxEvb58zgr5iyyKpu02GRWsV2ee4PDmnJk158ofqiHZ+k39r64X8uFosRPCex
UtgQKdd4bTUUBZEdadsV18KNYuOclOU1b9oqBUUTsjU8xqb3Me++3yBaQD6GPKT3
vrgMw9AY4mF9jfhIyzu31gw5G2S203zcmevraraQPkUeiLv3C9NXwFBLK0qQgf6D
GhtKwEGdCZTxjeBf4woG0QhJlp3UsbaORAw3SuGFyuUmjnW67Fe59mK6MhEpYtEh
6iDzWWXi8fClVuMwnUkUlApmsJ7EfGCMGPNSJT7m4qAByyH/5uvOt1p3g22nK3lt
ijnFsfymfwHv34UYrGiZQkb62RFoXhbFZG9Qt+FfheZxsR6Cbz+jIvAGFFcen9LZ
VU17GH5kD/3buCbiQ1RVmNXxvCN5YKeuNQnO5bLXF8qBvL0HaTPrHevzFr7DMqpl
xf5QKHGB/hGQReAp3GblRuuLLqKvRoxY+8m2iNNPq8MXrk4TI5O9fgHp2e810Tx9
FK6Cd9DUEt0SZAzmaZRQ3YbcTtnNKTiIhl46kcpg77vM5mwkW6T6Re78beG9g1v0
mhXqMOOiSZMc5exIHZzqdwASNFHoh7S2WDoUZmbm5rWbnPar070W3KD8euTev8/u
J1rDC/vcsYg7oWxxq0W7o3ELQlDL2IdZ/YAWE3zXRjtShcXXF5PwRfJtHn3lvwF0
8Lt3uNNynHTn67ROq2aq1IFC/3hcIic9sfOInhn1MJfBA1Fr6/CAXSWEMAXEv9rw
geSNIb4paWO1Kc+3O0f0kycAa93eaa7GGmGkVSdqMJiCGkiEqfu3a9h4XSzikO6W
L1sHK2BN9JRU/LzPj4dk4mc4raWEMem8k0qBRGUC3ijE8w4FmnWCBr03f9MpURc7
HtyOQB7BtIxSrzJenb/MEuQFfnnb4tq/4JpLyaqGQTxhIvT466yNubzVjt6sSwSG
mNQSfSw6NOZt4o5Lb/kD6M3n7hASr8vxUl/tgMc/on7ZaFeCfsRhBuvVLBTmBJBi
karU1h/j8vrfFwCpAkP3PzaezCmDdw04JlVqeK3naCkKwCTbF4XlSNf5lg6IBnbB
4FgPo8umrkGDvCZuBkWgTIoPZgZLX/yj9MSG76JlcTV8KNJQ+Dj6ZMfahVk7aOj6
lsP93T//zoalor1VBCBzspzMJw3V525i8xsN6+JszBYdtH6T/anCgJChxRsjHLjB
jf5qWnu693rehmWn4hhR1kFxzziHNv8BdsDWFaknm7Ut+OqlxGQwhTFLBepddimG
1EAGsmzFlO+1sW+TkjwgeYBlid7Vx9Xha+acPCLIEDHjyWPtfgRCl4x1L01yNeEn
7UXrcjhuLFblag29n17XIaTbwbJxijAgFMqvAcio5iwM3oadn3Rj91DTEdVK7GOg
Ft0EAhhz9vgpvbue2UA3m+T7YF7DoQ2hmUom89V9DDT/haVAl5t9RHLLWLoEricq
L8Tnm5PJ+4D4ZkWHHu/4+6PNYh45eD+xBigXhUnJEAUoxX4bJ/JO6lW0acutvWmp
qps4UA1YpB4TZOe1939jOatqlF43o4oBpAMQ39jOWsCw2uKsr6o7wliygsUl03b8
Ahr/WY3bOXnYdBJV6Lm4FDbEuFEGAjdyMVNNqqZWWhpmUtsfUc+EpuxIDDRCyFwM
NUldFHliWmsWH5wNNTTpXZogDWBDGhQ4g4Ty3CKHIHI08uX+N2mo/TVnGfxJos7w
iF7F51GCXoLDwErefNXkH65jQ/8cAugVLQsVPwkrs6qUvyx45gApD/0mN6S+dBaD
GTDfuhzkyAQbK1aI00Sm1gxdUlC/hfsX5xNMUghWlHUVvkpPJMzjBksg5OA5YPvo
L+ju7BpQAUuLKRPZEia+MP8l9UOMctVFbvanHs0+gRPRTLx2/49Kl99UWWUQELE5
Z8veyNvCZZ+TGOG2z1i+5Vhpkjor/jSQVcFx6JjF3VgX/wvOeaZd8HxA3xZr9H2n
XkQ3oTQ4kBk4qozG+ZUk7tSUBfx3fQ/9XCqERrvwIvYfXxXcvPN9qASigx64LNc6
cnpdRtXACgil+qQStb4O765ruD4ZUoMR9DC6ca18YMBbGZdZu7/SrGfsu/JpAhNc
ab4tY3ZW00zN8hrm/r0xDg+vofaYadFa/a7NZtwUzaXd1RV7vHY8sQokNKbNp6oT
nnMP37l+nyKq2PeEQB1C5BKcfxlXDgAPx+LV31K7q/KiaEJXqcp2thYv2GBuoTmR
6vOyFrlvZCc4YqAK8XHkGMVcXc0OXhopoSBUipvD/WK4DRMfcyV2jI4w/NFUjV5H
7dxobMm+qLeyGlUcPF5o0gHJun6JG/1wMdZO+Cx8IiI/fffhfvCMWvu7C/bE2fRk
+v29ifcYuUGSOWL14cEjW0Ri8tY4NRXNXclb2HTusC36bwYNnfFzllPw/LDtFUnI
L+CL3SiomWoylQRw2vcnpImE9KVOoxUGRwxMHEHLL/MNNFlwlMlgrk7ujU1WijMl
Ivu5+0Q/tKaa762F97snb0Iu0d+b+ZntH4BnML+WQUZb1+5eP+l9kWDiVGbcE639
UDa/RsslLxVvXMuF9s66IIFRMTcc/5wwUzcWwSFkWAN3a4fW2g6E3eTr1sj5IetT
DV4233EMuUBok/3ER4Qd27ZmBJE7PMS3RBuGDLI6AIre0IEFqII9gx08l88zS9B6
gEKJ8ZMmpupZMUFzT0lM8qU+dvJ54m9ZiDxApLXdhTcHTFB5iM7IKSN0MfnWXxxW
q5EzLuX5HSigX+BdFO/n+1tp8bc1ue91KFNgbA6HPTLZN0yGogizobsmd6xpDj3P
2oFSPKyLjqe3hK818uNarYxSateF0I9obia1pSA1ipF3RCPVqoHhvRf3TPBRPSwS
csHpvWGVhvbgSVPMU+Y2uJf4/xB1AdlPByD+Oo4sevq8zhs3TcXAWckjLn+B/civ
Ir6mgTOJ2ePXFlAbR4NENgYx4bQIsRe1zgfABhSIhHiPQ8H3eX0AYnh7inEFWZsb
rrLitKZ1Tfj61Z6aDxam/dy/G8rJ+haCZjucLJnGuk0Md5GqjiUNQhlehsfmiern
G49qNbsQGwlL0HnMf6mdOiUxKfdzIKPgTFRuND7PA4A2PQwYHQNJnc9+Rfdl2NAv
Hk7UeMTuaglet6MiIlEcKNT5DuS1ogJu0QJ0STLcU6bsu6Qa/3DYU4UkeG3ZkJ55
9ROmv2G+/6BQWVVz3RXUzhkr+pkmL9j0tPQ+xIL6G9dLMdZfSl2S6jVabVWCkH9b
tzvmniy/BbBcQuj88yHSfYDJwHNG5hmAzvcvXeUG4TCW0driL0vIT830axKsXNPJ
ccMVD3LmLJJ2JmKkQG00Ti5tIH8/xXSM+zxmcP5lXy9OPAGPmRDrVHRO0mjJ86BS
33pv1VHzu3hVO7RpGrAQ5a7hpAktpZfjues6lZgh8Sh3dKtOLB+rEQnkVPLictJT
XJf+rcAgQwrWiisTxku8K8EznLymn2CKGyhbxiPfG57090o3Zl8OI73gJ0DirnSt
qrDjdnuocuIRYsNkPi1vo+p4PZOy6bHQ2p62uBaM8/QiPEI+dppL5rQfdK59gbND
6UVJALrb4Oa3Oh94TRkyQOc/T0ErvXzTsVI+jl2RxsYdjxujI5ZIkDo/kgGLJykj
7PC3F2mEWc8rcYGKKt+VqElXrLO7MCcPeByZe4U7aKBuPNebYD7OUc/1Sf3NGDik
O1vpTf+0z9u081cruDxwudt27OucoKKJI/BZMuFywLYmm6CoJon8ZWC4yQmhhO6/
x9ylZCrvHXgqakF9roRGa/jXFhbcFZTD16mMGX2LpED3lrxEsNuIP9JgWh8TTQgz
Dam1vs2aWzt6KYwRo8gXws6D2U4v77icr613I+WrT1dhBLvwtYDouc18d+5SqUoX
/oo7qRGaaGiTil6iYEccpp266ewGrf2hKm2RSkpKWj5j3Bui8stR//sFdBlsbn35
t9VT1KDJ9DrlsOz0Ze8/ldpD5WqjXDK3yKh9FmS3w85JQ1BgUG6/dWF1mMY4gIC6
CPnpxMFDe0UrRur9vyhxSBq1AV4MCNGr0mmBl5OW4ByB9GfdlhRONpCPeKUEDv6z
j5lGMR2cDWiG3X5zdxPq67l6eyYVetVRlCqSKeDozawwNB+jOV7O/t4J56fs4eXM
fLXyk+ZW6XCc8FpxFLPQUNgcmezAPws3PAc6DzSsclOdgj+W4paUkFK2K9k4PdGK
QEZ30tbDYnB9uBqeaLPVB+Q0tSps0AzQHs5KsvSGsdg6fApE3WZUojr3MiKFE0Bh
gFMn3u2fOKEPBKEWwrQ7LtU6gy1wx3QpdySzBeEJnBESTpEMWvvGKgrxWhbOXcqv
7dxSsztyAWwz6XmBe8yz/eq3gU5p29+0vxFW5YhxO8byczEcJ/8qzQoHMme2EH9c
cQeN1cYobD9F6NMgIi8+7XUCU3KnTTuS97Qc/6Jxehg8ugd97Ge9KEJUnA0blp0Z
hvDe7zaO3R7lBA6WqnAIaU//IDBrj2/z/dJO1i0FZ+0WEy0eAnRW++q3CI1LvxcV
P6Gdfndsi/iFlPAMuyJbeP5lMObOJgrj1ob+yg/MCqB4uLZ9imfnWHg1AkwXUHIJ
vnkT4pQ0QsjJLRv0w3fWDpMYnwPJa+GQ0lIjdh+ynUlsFt4dW1cA7/3VkrYQezwf
RUC/ecQJx49XeEBoaQ4SFygAL+NcAJxgy2xuhkBj4TXWYkYP/7dofjMVN90I1xQP
SjDGqhIGy4nJkxrLOVb8OohsCDfU8CMDBBMa5KeNENip4Co3bSS2V0OtNXh3y08T
wjQjIef15v3dZjECLUUC2dMrgJWrdMVUo6PNYx58e/2iGH9vpx+OONLK7jz5+HMG
5ZpaRD9f+lh2EVQJawL0D2TSnMey8lrn+Bu8eSrEKixSvrU51fZG+kMj6XoK1dL9
RfmBicJFiO0NHi3FOuGVz2mD2oxIQwcmqlgekMYEKaWnbCCaAa3fqG7g5Eh+A1VN
YFVtvh8kKaSPNTY1Ugfwp6L5gagCMHRTmDZg+jhjyN0eycrw1tY+p8FaWsIxilwg
AUlldIfZlvG7Ct+CF+NagBCvQSV/JkzYHFJRX3Dg7CIzcuxLvbsVlumVJWYk36yt
/s4VUaxs6YNZ9W3WQz+9Rnb8m+YoJjQd02fOC1DHsSAJawUIcRtKnSlKo8RYktfR
7GHzqYSEoRGpnvS7f+fH+pbDh3aqb14kVU8whpgrRyjiN/Y9mjhGkiECcnLpmKc0
ekuoW4WZQPF2QKLfTSeDZDHNnf21pivUh0pcKzEw7Cd6+S9jHGVz+T/gjkFXEiNb
USTkR+OlWhTEmG5gSCBRoJ9628mz2t28bDWpPNNmW+doW42WLIWZRP3i1mZI1PsE
bcfbM82PwW4aq34C1xsmNQhL/vDs8lnWueSh7s6bXWBU4IU+uwtFXZKZnPt82XuG
RnwF/+tim+K2IHUQYk0fjSuINjnEb4YVCuRfynXtK1op+J2Z5zgiQYiFbsbBBPqu
69yyxEBZAbKU91DwCtuRxMfg11iDt1lj/DoMpud8m0DBQ4kPVeHUNaHPiuc06n5V
qlQGeqUBr6ip4zApsZ7bXdwxHh/qbkU49jKIkmwejsn8QW2GVggvYt1znc5V0l4q
zqnwuHAOaJggNgMReJMH0vSkFy4E19Ws2jtPHPUAfMJ9GNViUXYCzK+Jk1eBz0Z7
kGsTZQT8dr9D8KNAK/VosJwg420kQk3IcZJ5q8YvPuJ0PYSTMWIoxDOA52nriZOY
YKn9BP/zX7X36w34IUPW1iq8TW/LZL8CNoZAnQxtnodBSlF6yVq7cT5Oh8ml4yBJ
wpGBTB9kLd6uQ46NUx7+yL3Rs8ycll4sNE82DDw8XAH8Sw9mvZq0rS4TgRwpjVu6
3jc4T1srrSePjmJl1fHuqCmDvNj5j1TcY+c3YloTo2YSf3G7I8qQpPRHBx1VX1yN
LdpIIsqoJRJzt9HytFjdLpkagEvls5Rxy6LLa/50XDC9meRwA7c1/+QnMDTHPXi/
23kMSuXPZontrZn8ocrec2cda72u6PgDcQHDSiULgx31OFBbgc7LcKcTP4/+8M1o
HtOCT6QNolF/rKG64iT7IuYevqb4IEK/GslDJ1ImH7WD4P7007WDIw3j6LCQKLO1
CcHvGKo8cDtqke5WjiqAxA8enH80wohBs5O9U8TUhPjobEE4YJumwdWWtjB8ZWNJ
GYP+6/EM6AWv3oqkkAEmEiCCnNfCY8CZCD7LlTw+nk1iLEQqv03dIna+pzXhR/52
jSPSrl4CBo7eE3TLnJDZgZRafqwrvw0l9QJQQCqf6cSXDvRcfNwHHf7ftULFpk7f
5OYHvQQyzMd+rauBf7Z5NMlgDMWV3vdAdqakQVqZaueJrCsq3NHdnhbbkuUO4k2A
W4pPib29XSWRzpXT+JjWizmz8JFwXyDutiIXIBTIAmw4oTuXF21welXjIvUGGhaA
Utzh+FV+XHoJlz98VS9q5aEBamjxdruZUSqSeG+N3hyjwqbvgfb00SuF5WciP5uC
Vok24sct5y06DgnwCDGuoHtiXvUuxaJjMOCwcvCnUmyvADjE9fKQXMSL+3xDHTzV
5ChVNJiCKFzqbUP5g12zRyE9V4o8/v2QCrcl80gv9ui4T2QMvmEHPIvAycxFHall
JKcn6l4M1CcG5HAj0kMdIBzg5V76uQCjcmaBKKA6MlGYAZJLyI0JdBtBBhq239lJ
n0FOv/5wGcnDcemqdBGULS8HMsfUMKJQ8RMNGD8JLjZf3g7b19PDBo2u9zo86ujy
0HzkUqA3dFUWnV6oMXCGryWHvmJUca7rYXObt5SwosA67LZtXL+PYqCjkWy9RYYX
C/iZG9WS2ZeCAtIzF7qG4MTfnDUnBjAcyjmRzBxQ+48GIz7IfHz2COTs73DuDNGe
kyehG4h86A6Aa62UvZctHcUlbzMWMvmS3aWRXzDvBW+930TiD5W+QbBUdtjBbjZf
r4tjZHHjgIh4Epn0lmGjG9r7U/7luzV7EsGBwXBocyUAjq9HIjlTNPqgn5KNcEnK
6WuzDfl2LQjLVPkg+/5ErjC7Jyrza9pzIdr4DguDuJtOn0IPT+9QRJAwpyg44qf6
xmEpmCCvV38TcjZ/zHH/A4qXG8NLqYnGRj3N7wrnFRbhEijoVUZK0RXZia8KoMcJ
MwlWmTXjNjQ6Kl1G6DNGG8cGdkvOGo5zfbsIXCGyku9dYehf6bnR/SAKDt8f2oSx
0l9nOEVMyGJL9L/8XHbPgnHYXEOLOV84RSrPdydygwX+ZcbGvTi1rxDPCvx8qqjv
ksA1vw/sH+CPbc0dNsnXAwNm4FV4iXgRFyOca1DDlUQkqgG2dWxapO0/RCk1XUgB
ruvc1iU1JU8vZ3lucMhOjvv3NfgSRy/teopTNnwzXWtQQ5ZpiOM2JPsBT0rEcaeu
JJJkmTQWOywG0+TM9uVRW2VMhDMeHNZAhs5nEIyq2HCJ9xDZU8PkGxX9Wfq5hx3e
zMZCEe2WNIdAPV1fTkLsCLUqan9eH33YVNPEFVigpLPAX7x0/1JmvDyijbDXLzCn
8Bql8AOwOrSnfQfoPGKidNvBWXr546uOh0UCZftCEzdYrI18sMfI1FUqTq2kK+4e
IDj38M/mqROyEJMT5TbAQcVDqy/t/O50/pP2FSXeKNqyXFO8L9E2M13BtqH/m1Pb
oQFkebz/+NZ1tOPsmaVCN5av3UBJ7k1jJy7rOSLdR0uNkx9cBAzzICB3WAzczO5S
3oYbitawMgfYLIksNgRQg+e3BI6B1sLgIbCpW/haDHALTIflL8Rrk2btKkSE+Wc4
8ak+gL6jpln5XGQqD8n8l5jGVDnnqBcjXCOuDAoPaXleozXHITwm+bISCeqTOmK4
gF41fhSU+3I2Njjq6x0IqqVlqePiNVYWDc0/wljeNwp853mCuyby2q34Kpyh5Tzl
RNBDGiwLlCEgwp9JgeE2lL9dXmQciyidgYmRw4HGjTIJ2hHhIzEeeDC+Jw1avgRO
i4NQSCHkB+NKiY+0cst/mdVqT0Tl933NpvsmkQhDupnVuBaGqoKoLoCR9UdAoxky
aMz7RNvGrilVpLl+3++/L19DFlCBtVy2tfbzvnn0BelVETSgqnpkDpHoj5A1USgB
RyPrEBZT6kgbL3HIZPk3rWPD5OC4V+juK9cg9EFQZRKJR6yMT2GDcUB6+/KcAUbx
tBY9EOJnakZURtwp3PYKFIUEJSvfroz/dN1sYKZSiB7pgd1VCj+eowso1e1yuujW
IqUlNh9R+KxTUyLZ1ht5ZklZ5qXR2JOA7jWao7qMT4AG8nubZ8uNvl3S/LtyNbPB
JhJ8V93RebfiDUtr0WCmUywVE31+J1sXKFTvKDtQUpcgJ9ykYCFZ+As8f2MuWtqk
eToT2qb59gN5rA0CIVDoGxPPDOdIX3OxEyYaKq8Qr29GPBrIKvIu9GdNMjkdgbqE
DeYbGtx8sSBbDyqAMV3RwLpkbt+8LOp+9IK7ItVOFr7UtfdkY13vOZK/W063zCNT
fsqhEj3H7RynMVX99tPVnRpqyNmZkWIFCMzseaT2tcUfW5S4P284rmwMtgOKG0Mb
zRFp5y0Joot0x8jvbnQW4FbJppZgCed1sgX+Z4jGXJW1+jONDHaWCjKTyoaAlFJj
QlzbS4qIU0X2fyVYxujqlVmpKBLlwKFbUYiVjFYCDQ4gYXI61fBvEbiMVcOe4r6z
b7KHwkMyctzg9cpRixS3FJt9taW4se2ri4zhk1cnk3XH9YehrdHeYpxERO/MQT58
SyVATbJhOlN1ZYLrqk3ZyDuA13LKRi3L59OpRclkVWZ7SPCJcnMb4HZ6Omm0v0mp
hwHsHnZZw6Xccx7NKH97DqO9rWi5aiXNztBOfNbAo+UFykwcGbL3S9FAkPi8umpD
eaTe45lL8tJunQ7ad7p5h3/schyYhouFrCtogjOWZ5j6rzTBhIDc0p+Qu9aFtEO4
3ekqFpqXETVqrp4nGci7ECScRrasDBfdmxRdmrfuuLGbIugHH2euRpRZuajqRBWv
8pBGLFIlHnEEOZzCkf6V1LbZVWKjGjuF8OYU3GQSPoLmrNmIzugFsYntbKqsHJ01
2XTX3j62heDIYxTaCOJyy1OvkmIslMC94Kp9VPgBfUxHEyG4sv5NfAYmOJNdAWVx
R0GX4pF2jnVSgV4+kN5nvIG8BdZGPbeaFzlrkZa+0aY393NBb/nBc7Xl16vf7DrO
qOsG/9g3T8OjtoUGnH56ktjTRw4vB4UnbUjFozuRKkS89Ik7/vRcAFErW0dFCEaF
k9p+F/zsujzkZbsguJII5ya5nl6H6RRTuUx6dJKtk0gQD6fC6pXRZZQ/phacAd9q
wpH4KaOpe6vZ3GAn+bNA5EV7qGlmRkF/9lvjrRc3R2J+WsJksGVPGRKxw//Is7aO
v87uY+ZLQVWa9Jb0EXeAOfJPTir5ric93ne639goeESZDpPi9Mlity52bsTGW+0q
6yTg3r+op79Ke7rzSabIRFoilBSm57lWLDJuYKWmrtrdSatcPq1gs9z6YslYwAzt
rYPLC3fYXScSalI7onXI5eAp1fTaGHOF0C++DyeaawHTWDHvEuf2HC7Dsk6uCE+h
VtiOl/BH9b1eU9HSuEn9Xow9Gfq61rsCxuQWL90KncyTXw8ERn+D1rjv1W8ey2Z1
sGv4hym59gyHGtWH5fn3O1SfvaVNRZt/edt1ysoEDIOtRkR/pho2lQr+u8ijfWA2
VLj+X9PwPWKkbxYDKkZFbsPqBe/1zbk60igEfgnCzMHbJ5xuSt7c/5uDZVNIKc9e
yMt6E9C6VH4XlN9hYiQNvrGjooyL/5KwYeG4LD4YaufdBmODacO8e1ufjQbM6oWd
yWfbyPuJ6ZfvKGVpysmm8fDmVZ9QwIn4Y6/cWu0pRGKJbSGWTmBIs67JpuLlDGdC
l3Ls9e1uh6cUJDDnsfn7l5hTMUchL8GcRsbABaBvZCnrdUyz2jkq3E6PmOljfjp3
Z4Qfg9xJNy9MYAq/oybIdKm87KJja5+WLnM+9dQEWQdebeuIwAoRCtNjsCn5ZJs5
PinqeXdrOGoQklkp0yorjsEz8krUsQFq39EM+Oj4oL9cgwsvQskVpJN2KBN5yRE/
eaMhApJtup01yVl8ntfT5lpgF+QVDxutUqzSibSk/ZNRSK5dIxUkMg22X9WpLHNo
gJhwsu/hY1OKsPTj2CQKc558mgKnA42T02mI/eSleIdsd5seoK/4LNnllLIMuW3Y
jISn+rtC6YbC5g94s3RzdPDHX7ctV69NiPUKSILvFw9YHtbKh0i1pYI9b3jh/QMr
s/lfa//gf53/ujVKzoLwfyD1XnFM9FUrKaLKki7ujAcqaxT8YhANi8uUWwoP7NDC
YegSvNnyJWPuXIhbWP7DN8484kW8vFe4TlR7J8lEjGin2LWGXsW1FbXfIIjKumbA
fFhiT5myinw6c2I4K+5rpXTK9yR46lMvqQDGJLxr6TFNPjOUZI8BD7+l8YNR3ryv
0YRDorTeB8xqnzDtRdQlC5jbeHl6treM5eIfsLjp/Pi/9OI6Teqn2KaGMAsmpuZp
MeUQL5k03OdHuPv9QxvLCwgc7rNyBKToI8E/+fyfDsFKYgb3BHdiBdY8YqckqBA1
42ISb+caPggQPHMjFkWLOgygLpuvykfmb8LPC0dK0ynxCFNE/VL4Wvglh0jFWqmO
Jmky5HmQGQRRsvpqjA78NqmZ/bImbp7rw30XKbtDc416PMN11VKiZmsEdU4acgG4
dRQ82A57ChkWfD/Si8HsAQ11SuUaXkam+YM8wmOxfwfnZ1rwB0+ar/3KUdKCgcA5
T8KM0JZvaIZP9ksuwfsLUjt2VF7TakzBf6r5Xw9Zqqgamx+Dn+nPla4CsuV8MUN5
R0ckDhxrsd2nHo/QqUycVqgzQQDXuNtQBgk6R087mclLg0Z6QvloZ0c9oe1nz9Wb
csZN8FFCW8XoQDhAZpLYMqmGrrmRTFFzqcKV4oEoyg3DMQhCdnXflFWGu31sSPZR
C4EGdkq9IHWDrcq8ek6A+QKN45WRP555yj5A8KDQ7pFTwN+4uAKwQqhkhGeDaN0w
KFZRaTJIxAhh6m25fL4soRWSF8/nGWhIMxggqJw/9YDYZsSorE+SymFNhAEFQeG9
lL+9rf2NKKcf2ASAM/I8Bh+V0z1A0DpstIGq4q3lDoxA/2SRL6v+uazmJh1Yfjga
iJvyDZFogoatFMkG51tZd0aTwPgS02+uSG97bhyeaRQA/NXH2owQdtGzyhigXCHT
c/ClDj9W12izAqfueS+2AnkNFqRSFMTxzWXG2TqXpLB3rQt8YWC8d/RfOx0RYOid
tPVSeJ5Cu8jQZaIQUXMXAdACkBw+Um7lNgAc9/wL+2pqqAT5zyQcIuaTkKUgGpIT
KNlBNOxxVTm9lAe6mjeyTluI3iaKQDxYTHh9Zepz9xhSXp5g6XiIuU7ZK5dQ7HsO
Q76zYMcZKDnhoX6K0DArVeoF1fM6JLqQRhfR+5tEIxe4eitZ6MIVp/sREKdeXXc/
Iq2vEy41rmCTVupjesYuw8JRZxfpVfb6ZyCHtp+HPNVMonmGLu7DYRG7yPpbCDSN
pkJ4uewuVDu5oEApD+KqT9j1wovrVSAsnVcK68qSX1piF7QqGDpsh1fypHwC8g75
ZZL8hoiFfbdlqQoUQqozcs4VPwyrb8StjjM0152b2BqlweJAnocI7mTMVgXrWaLs
UcIyyNP3gn1NSxvWBOIe3Eu08KGU/Etmq0sfNSQ9yM6hxuxTS9uT6C3w35RVdl1u
E0jxSbSlwLtoqLzvGDCHOnmZQo/yblK/CtMPqIzApGiXaMBxmJ6DEbEd3HMO45qf
WrSbvjJ7ByqcntRkLx1ImisrIlZ0Ev7tdSj9l2p4ylrGDalGqpAIaLQUvNns0dg3
+SvogvPAcIfvTVwx3mhFb5tlKeCFGJTB7LYWpP+DanTYlJk/hKdgGh8cMrJnvW96
3HqhuRaBeZ2KOwK9wJNIzjOsFOGH0psFZtryY8aSKgup50S/wPvUs3jNfBfHalHi
QYlFRi7oWZ9iKRRN462iJFDstxVzIMkqqmIovHIqikBZlLtMo2eSyK7nOInc9sRI
FWx7VZYawr1mpnqoFgpdW6C4V4HorcUQBdUxK2G7PYuqb+QswSE0RnLu6+Uc947O
6Wri1yMgounmt9r+HjIDcX3S3F3rWFy7BWcna5BXsoYfEJao0j7+d/pQF9Rk4vyA
aQ9D47V1dKcktLdyEei2Obepi3aBjO8Azb2nPM78GaRJYAX4Px6CtftWkoCm0wbW
ZtcMSJ47kLMXb+AVQ7A7X2Vrzk853G0Ng1jHQWZIJoQT5CkjmUMvesN4uQprUUeB
3DLQb2QqA9lvh25cBP9cfx24v5DQD+Xb68gpEIKGV2TfXiaA0eCYUzQrXGGiyMBw
t93BE+HA/VlunQbfU0S6dMxaX0m4vL/wVHxNzjRxjAvuSFg78Wukxmzrw1nOpkRd
CZLJHpOPzSvz7C/WCm2I0tFN+B1uY6pKwDxX5DSqKIT2oXS9LoXZ7DRemAvz07F7
85Jg4zps4k3rpHBfGfk85XgS4/MHUW00YSo0WE7ut+HNOHXUa/fnZtf6Kd1TAz/G
Q1DDDQSzbl1BK/9XFmG9JIZ1yHjBWeIozKk4wVKaZ5cqIMc0JaP+7tOHA1oGUi2b
Whg5XfNNeTljRPzMgyUQ5t2ixTMDzve5lQFWbd5kH6iQHd6ukjcAvjz6d25ayBFT
5Fain80xZpTpwWf1o/hkPJ2FzN294hAaj79MYjildW++87KOUtLBkxnGxZ0qU18t
O3ot16VBNXd7V0Mnhj7jEJbz5jH3SCAfc2dJAGvbSOVz9OKz1C4AFhJP68QXPjat
mOt5Exwf4iJMXgNpkYWn9yLWUbn7NK0Zfo/I5gLfvSrh9le1feXMffCxTJSlKac7
7VHvQ28kyW9oxNiQJS2+T5x4B+KV/mgFCJ1nTAIHtXH5Bkh/ecfJxS/xW1iZfVBe
wWs5DxcRrpq0SXqO7E5binraZ7cUUUgRfzwzpMVB69NOcbwxjC3b9zsvD4kNivf1
RfFvIeZgHWDh9LKp5haQtLwXW1B8GXFCZs0iBN/KLM5aSs1fl8+Clx6WQDjAAHP7
6xYNKP8nDeqKnqmLm+JKY9mPOpXZ3vNxuyuftBHQAWVj5J57kvoEhv7LEVo1/3yL
C1AQK6QPKlIH7NeUlHaMj664LYCekAUjSgiYBFLtwQr8dedFHmKGP0BoUJ8QuY/e
PbK6KhJpEN+ZXwN9yyEP1hM2ClRvcSLzbrYlTjVqLNrM+dIS2W8w0iPSc7tNMOCs
O7eNMR++jA7KG6cTKjLXWkj4fW0xKb8duWUdhJ4Y5VG2MZHbt4y34PPudTu5OVVY
+zwgbdyktjcz9eHOy+2DBdfeq6ipSZ/N2fVOnpDhFnvb5ojAvUkvAx6rTYx57+b2
DKTtWzDG07a0QpEZ3CBgA33+G7z//PLYl7CaCqxVjZJNhdWY50ZuBUqtEibYSsbN
8kaWzscppkZWkcyABVtE4nEKsgmVZyDygZ6qMt2e94zG8GcE84olqek0w62u2N/c
oCIOB/j1cQIQ0p14IQesrw2wX8E72AArQl7YHVzggHu7CSVZgS1SuwDpqISTIdnR
61x0pnlUiGaHoMXomsBIwDkVKiNIfprBCckq8qDiqs2UGQK5gCdaudviOlpJ3Ids
gkqXYfiZ4mrH03nHGqHKW8MiaJcgTJDZ3/US/BU+rEsLbY0s5A48WUiLfX3G6JRh
9IxMuLC7EIyUzrkSU2TbzjBVE7ergVqs3xVbKp8QTCZyxaSua4Hvg7B+860m75DE
4codLE/ayso4we7Y+I7LsqlB9kkV+SmtLnQ8xxPZXnARw+OVj5xzhn47ShNeVoMs
09FLuw1SYgnlUL97mW7A49kRdEPUtXE6OkcK2vOHD58lZRpEHonH0KRntv1tOuYf
ufD+e733LYBXDqj9kU3WXt8lEdtCMWIuGEU1qxHsWv4uw+sLzL9U1K70fkmi2lia
5HrsnR+FItMlXd533MaLXs3tvM8tT/BNWtndkaVeZNv9w2gs0HnFc//r4kdk6cFM
yX+V6Vq6FtEmJfpTLOsZwFyp5Nr2aJ7C2wZ+HNeerfzZ4diGZeFGhuZlWLop1qCS
VufwdBRFbuGdeLHY2zcOmPT9hfRoA1XSbtmYS/wfzXAWDNi67ljJlmiD5X7XnR3c
mCtady6RIZe2bUuDwHVjrIp1M5uh8mXropO+zFsw6s+Nho99Aj9vYEuzSnU1sf5G
xLDxMWoTTONhNJMRqsmsQvuswjgy3kMMig6NFGT+PwweEDf4k1gDf6Sep1YmkNzt
EnjxwFOlxnWlKlr+liOqYJVaFD9GQoFfTiP0ScQBPpC0K2HZTgp2GsyIEiMFA/6C
UYd5i2V/AeyTQjaCgARXHf4QIB1NFaCHB5MTe9Rw2bUzAyYop4aBt87AyjHBeako
fhX1bQ+cR41C3lT6/MNIvn5shpLlwVtv0EemXtkL6BQkoM5aiH5c2LLSlOs5mrM+
zs/hwakpuwfQs3mwehEbND2eEV1lhL7d7hIfEZSkH0WPnADA9q3oSpvyn00FFAQh
ppsx6KGj8Jt7tYwAwAhwBMW4uHrai86tSE2lnFZ94I2CfVeNNDVLSRViZI7DaQt/
i7jAIptKzwgCtIMAT6nqkLvq+E5rbrkVFFXvvnHelIQ3JuU1dHUdV8hJJ1+YYFGj
N/uuY5VHuCTKFgZ6DgeZskdVMcZSma5DxRNcv9Wax1/erX4yNU2fQ8sT6BI0kTve
jSmwY48V0KT71Bj9Voi5jXXsfh3pR6Yz6PaI1tusbvw8lgiR0vrjqA0fLT14HFJv
NR8W2cidLZzl9PjFLHJa8/EGe6oeq6/N/HQbZd4/HcJDn+d1SnrgB6gMCTqDiq4s
63mbUf8nFxcuN1KGUvzEMDkqxC3iPz002qOi51kPt9bujJpKdYbb74UULlEmstbH
JSCGRD5+NWV92512x9AhYineyqTqvpBd/nkXPaon4QWr/KToHS+HgGP9eoqdO+vO
xHLtbdpFqAKbUz35JI1GUWUOirVD6OqVIcrrxh/rftseg/RGYY9MkOz1lrsIjWKz
IL1IWZtHqoiG7GVAYIMY7mL3sMforkdaZWJMERZclNC46zmpjBvY7th9UzL+yk53
eZ55MGq5XYtFP8kHzykmkTcjG7Gwel0iC30wuiP9qgeNJhTXIFQtOlHarokddujb
laqfPS5rtGtzQi4F8krTHgy8o4f8t4ogntY0Tt9T/ApBihDS5GEzriIPe+innev9
Bno0s+dN4u2KPjG44jdRtE3JIt5LGLfD20DJ61yMNsrfxdyS2Qw28kNkro64+Jxu
bzs4s0Zv7s89rAjoO7uHWinhPGv+knT3UGmrL3l7Yg38V9kq3R43m6epd1LxPqrd
ZgH1ivgMhtLqBNaPCVvdGWFuPc2RpOAFPCwxjmxzodx+NpNUcUz9GZHocWqWhFOM
10RWUxjgR4xEnPqvBkkGVXGCZxn3F44E5ZB8brHcDVrng2YJqqEjhPkE+I04rZR4
rpljcFfOITgLFVo0JIt4YVjgo0zAHQvL+lCmqVW5Mb0ytj7L4MvrKADlmjwkHX49
IjSYqmsJTsGzxlY4JFx/cuahAMpro/FJR0NdNnpCn9WZXSwwrJv4Pmx/QHccdKm0
nqNYQfzilM8wQ1R06LljEgvmG3+MIKOIzi+MsuRDQWqqn32ok5dDUkppGai94tqY
WeJFsigUdI+IwPH6t5ofaYXez4vihjkQOf1ZZpgcCa8AEfZBEFDQtc2G9sRgS7x6
bIGh3B06JREezMuwOdQYOtns4wcRliDLwrMX8cKIswqLPgT/A1QTod48TgQ380Cw
ycd0s3iklgCUTgTB1kDtBTX6DhX8P8+DIvQSAAHlfnbHE5Z7zsSveZgQiVu1GfC4
jO/nj5Wgbt8MHZlnHGbHFNpOjWkQNxO+Ggd2fz+VaGgrefWu/81uD21K6fHulaxn
iDdj2yyiBuaq48fB/0wvzK9shjBiitSKRQQI2Tzf19NK/OOujrkdXzrOE2OgW3oE
UfbL90Oty/N9lODssCHLYRyF7xNElnKnAXv5Y4FcmRple6oZz+dlgCvLg4gM0AvZ
7gWc+dvYW0+ZB5y5qMxRhSqVwLh9StRiYCPBRUjwkg3wyODP+P7i23FsExVHSYeL
05Sf1D53u7FHewOHYtMItET4uAgyk0dW7vIta1JskmFIi9soJLuj++eAkG9QyomA
/kbqvHcNg/7FWsOQB8YCjqnNvLklAwufVdC4PMujxE+TbasbkwbzQgdiRc+5NFeb
4uo7BJwPTNwIihaW7MG4eY6qUeoMoDCFrDRknK+ScxNYgz6vCJfCkVO3K43OlVej
KrNffiPrOpn6gtIDexkgTajr/GU3bYvzS7lLlRj3Z0mwC5MRg1DzjWyzJ0WKZ2cJ
9ZhFNkMc60LHY7583OzsknkwcM9YrlO3gJzPTRCH+soa6Zkw7A9EvyYSTC6Y50Di
AlIzaUMbMlBthhgJIuSmdzGs3yCB+KYdUYPOHgEikzygVjQTdd29TB1Oqjkmlhc2
pwuB9uSFvpyJAxc4soyft4cgBtvz32ntSsIu6NlZ1e3vjkLnCWttaO54vrAQHHWQ
47OCqxWsFDyyPALVHzwkf/H3urp7BlZ3PHTs2vqVs+BKbnm0Cx1QeHHtzSP/hre2
Lq6IMoSNSimtUa6RgBE7GB8AHJ7YMg7uuzUYsT5KUjlBkyDmHufIoxq+RITHdsOA
wplvfqcT9W7bzeAS9Fu3C+HU2b7UGg7aVW/GPjRY4eUk9I1dPCqU6TYKDvFvI3+Q
zfpOPf0AJVolvqlKC70DLQmZEYPOP0YNTQKnNG08VMtOILGMi/8gPyFpFL+EWOMv
UDAe/XBN99fm0fGZAvQuS+LG8YZIJsvmmyxPVbP3JKkOV7obdAXm+aqfkn9qAgx/
K3sikuQOiTl67RwDRmXmdzQi6mneGRNJCWsJmxc+h6Dke7VBeLR64auNwJwNRCWa
ekVIB1Mu6PuJCgJAobMvwh4p2Q6TYWboOjsp/ZrYY9QC/fbfSrEwuQCg8Lx+pSQz
omFSkTdKKBvcXIVWmhJU6Z60iVcgvN6IskPppx4UGSeiq7ra3sSGdDAJDvJYMd4Q
4QLR7E31ZWlS9BdaXAgh4Lb2fx4TQooPnp0JJUjVbEPLpL6lOjBAOXCGi7xyfVup
PEA+eYwdwitt1RXUI6F1x2c2q9fiyVeJLH5rPPFpIPT6Wtm8o5xbEkqmwf8TiO5v
GhI0jXy+E7DrWsIih1OhzA4+c6CbkOON6sMiEk6uBScnzHzrNyafigsjgvbjWk/R
INquCpH7HVXR1+P836mSZ5ITEKg6teM8r9vL4+3Athh9XivoEE66MaFK4Eg/Hwsa
XPYtgmazdCAiRSwU/d0ERrCxmL3Q3eypW4Wx+L0w2XOlicBxo0Umt739I6IgW3gV
MDy8K3+wFnRLPn4Mh8LcI8jrS3TMETpQqafkFilKZ032QsTqrKfgvK7KRy2Ip0XA
pkamZbA6bdkyo0L+r6RotHTfRXa3buAgG4sC+Tv8R3Fx4LR10IeGSPx1+3rMbmU3
NgT5v9wtklUyuwItKuAay+0M1yi6/Db+DfVGreZgv9IiO23ZVynx40FF71g+xgEb
g8RWsItK4Noe05CZ5U36KcCt0GtbUEqP1HYalU8BodOWx4ddZIIASnlYi6gFgFrK
a2k1yUYBYfTtUfpdW0IY8W6fJnlJ8zwOxGpnZC/j6OEH4/tenhLq38xkjMFO0TO9
2bgWtFgEQBYErYO8iFm6/Xpe8PvuwMc6k4nBAFmaeiIzGTHTVjJTGnwIr6n0s6KA
pRir21wDkQpRM/JvCZcfGnWYyz+/C1F5iOz4St6eWnzJ2liPI6J3iCGlTKQ2z/1w
sfNcDTquVRToaLHq7I761X6+vrZwPKSNA0DdTSfubMJNZtCX3XxUc+460LNYR6Lk
y6LYEkkZ0D6BOZOP7rHPBs9idYhmPqosxpf/eVxsABn+uKvNpZI4yPOA1RqL4cNx
lWhGArV5aujDkNu4buf6l4IrLVZm74kvelBjgSpbm7d5+gmZOkR/6m/HIBwkY9WC
hCvQEzDyVm2JRlzIEWCWxLwg6HIm7A60EGsqT8g8/UWFOXspbNih5sxflnXHX+Nm
rt1wFM1LgbqtEpdRrea/JQHm1LjQHkYgGw10hHjoeckWP+KxDNQRlh9JjlPbP8AD
CX0haNiCMDiLr5inQ9wDS/87mKmnuChucxHHv9t5IsV+LT66PQRe5bGw6lWV9sKw
M6MQqyMTfmlISr53lJ5fUS0Ena/+yWd/uWtUuRp6/QWeJj5Ip0pC4of18ji83NWQ
GtiFDt9OCtuW0IjBkio2loKZNWncwBuXiZntTOBvWXVx94SWrIN46iZT4+lst4hc
KB/nmxWDlLgqakViu/zmXzMZ3+Rj2yc+nQS9RW2yylY80+FPDnW4KOHBE9oa8KhZ
3IQ/yybFAs/GVtZ9NnLMk/hE++sNgvZ6aemj3uVIHg55hdAgTlVy+i1uM7GZil46
4l4EqZ2HjNiDzlegUBJlPa6X9S3Op9lm0S9RqTEuLKzoUpsGuPRO50a7m+XzgVMH
Oedycrd1dwzLuQbszzQNfN6ecxRe1DprtwyMhzMvNWHIIVWq+mpU0NHANeOaUCvx
Y0/z60Q1so59uxZHol0G2Zdl5Efz22x9QCt7cFCh/0i3hQETqECXx75C2Jw1vjDH
2lY22wLrgFklmhiyVwRnvPq4DKKXHz7rJgwyZe9suFRgUfRgdLBjB6kuGUL8l4Gf
AsMs9tdkpCli5Jr+NWd5c2FM+OmMbJyFstTpNzVDVvXm6NnXC1GRYPlEirFS6+ci
svmS4cKJ0y9PFKe+kijNJUfGZvoG+asLidEoZHh+3VEjpfnDl28EePT6zZbHReci
OFewCu7iG7tToc+NG5arXiahwfqWGb6nG4+gCO0tR1vBrlJtggDwbSTXaDnYlou+
4e9dSTOQoohzUAgUzpS+F3xYLwfDf2NGvtozyh4EqjBkaAb/czZvMohFAM1EhPcr
J+rVnbQbgIh3eeizahz0YP96IlNFrLvP7KKisvacRhJfYh04XkLi/aTD9fK3Gwgw
R61QdFUp8RPetuDjQFwpKV1aYaj4hacvCCW8Gb2mXzrM9341o8dpZr4VoMItGAud
Lwtzn1m4l9xUzoRwHXXwQCeqvrLHLeB2FdLyB2Jbr1/dgo/B0KPgokyqNBj1Y/jm
fXmoYtF6oTM2Ms/o7EpSygTHzx9BPo6tkpMmpd2o4sULxZXLmGwWMC6J742bDj3l
8a4HMxvGuxO8mXnMm17SthmfYCNTXiSc+t1ckFWMTBdWtVG2zG0xr6ivOipPBUuS
C6nNAkGcJ1D1//hXF4BgxJZWNzIZf7NPN73Zz6BsxHrSS3vD8nqmkiYXsZgSWGJy
x9wHf0SZjP+hdedlNTIT6XMcjrEcYe4rQ2JfB3wUgR8MyEzwXDB16xZnVRj8+pAh
tCRe6tG34nGop4gh+zl4+K1pBv/bkwRhX1yc7dpX7t5qwcEnNSeaU04GXXXo/+Hf
/XZukdm9+9wSJlINGm67nAhor9epN8KD5v62DK9C0Dk2XJQByR86NQJ1Zvrcn6qi
z2sJoUU4571ow9+ccsP9+AEBQUL0A9+lMDw8MLI434u/XmEGDqgT5ksXS6YIcWf6
v6QPXFoQ1xB3n/iY3OrqLrex3h0Y1dUdOazChCjBJWEMJsm+WkxczemqXUwcuT0r
mp5XXrjICKCzXXsjjxlG9SFscbzpuxpQRs4CfP2SvTvFw/FHO/To3xXwWGMqGTUL
GtzD0gvGeDEfW3ppYC9UG1Cq1gbrEJNWv0WCgB7NftypT8nxtAhJ8EyVuknwtYaZ
gTPioa5WsFLRyuG7S7+4ERSA0sOIZ4EAhYiHMombVApF4rUHW2fTO6f3Mxova2KW
UJH+3h5iT7GmJkmumO0BNwo0uoy8HZc1wN+Imc4+vO7/yBQeoKf11bvCQ1anRrOf
xjvt/HB9XDSmY84LhC2kNEI9AauMEUEpLZcsX42cbT38ZLCI0zdgJ0XFWQ1qzkn7
vQHC+/9wTHggaD1b1vcitOu55/Nr529jydfJXHDYHNu99lOy7aq6Qpq8/XOllCvH
/tnsJljeF3Duz/hBUfG+yCksmPH+taKINZqi2Wj7cNmhgRxubmn3h6t6Nm3UM9/+
y27QC9ETlS3yUszB/7YWbBoKJSZoshLt/8rB5zyYPpMakhk4ozx3zg0V7OEeL4pb
YmQnknLFIAbWYpME9RcrptVJ40MBLb1Pc3sYc+uuO3jQF6cXyOoSi3fKAviV3dSk
Q4HdWrk2bNAc32DFsRjdQgNCOJXOipRPPyvoOHYV1sfmNAquiNG/vLWxq9Tj/QJR
Vb00c9G/fxY4MyjEjDIKcU8Lrn01t/5+pLV3gnJihPDdTQR21WADCAJVBCv/alvZ
SxBcEv0UXX01d54H3FY5r08xPpZYHyj1NV2sBhGxU4Q/FDKuH/NYVKMw2Zfbk56B
LYxDKqEBG6MEE6oMriaxKh3aielAYZOHNvIkcoEd8Rl1E/DZsw+qVhZ7GOg9+CqI
8mrvnv/pq7bk1KO7s25uOTuGd1XAZvlAJVvqc3DiEbbP3ak3FfurT/lQfSfwpxYA
dRu8EgmSPV5JpjgUfMTkbWzxlJKqDrR1YIuYYeem/8Kkq/BAoXGY78U2cwYmoyCu
gE+LkeBSUL0Q76zG5Kgw0hc+LCkFqP1WJl//tH5w9xuaOAMqTQ+BQIhk+Rx5eArr
XRhcDY/uitaupgMatzDA3YSDsA8hByl+GDo2sdf2jnxHfS4VUNWkt+51gPGnYAeN
WleKkTDHKH9nm9pLcCNpXvCCgXESG/Qr2EljYroGoGJ0U3/ps75xXvWcStX+rEp+
Wuk45ZtBB/wsvvPz0BhuXzvLAdozzYj12PFGNGhB9z5xL5DBzL6DjWXOcDXkroaZ
5yaE6yLDWsnCpuGIFfqGVnY+iS+gV2yBmj+noYXcSc8ytWWjx8FWiaBH0T2q/i/A
pFmbgIgGOKJ5bVk7wbuU9b57HZgi0olroIlPY8YTzqTm+KVf4HTP908GxIqD4Has
Adx+fjSIUSbERq53JejcHtiwphdPBGbEPTX8zGDEyqth7dBJmiBqyeqYBClw3lN6
H2YpYLYALxQ7qppPHHG/6hsI0qMq4mG6ytLWFSNKt48xRCLwgUzfEJvyK25jsXpp
Yf8eX5glcUgp3rhjfabZWpaExFeLyV1GjM91oZHKf9gsHUzqraJCyM/LmbXkZamZ
Unniu2SYbh1fxW0CLY4noIPi6dN+E72pPYk+JKl1nQge3vMM9M4fY4cupNs+jvxp
d1B4Edu/d3S5RsTfuuaDQ3f1FfO1C8cU/JqkVvw3SAxfzob2006R6Blezousz37s
TW7ek/jcfDx9juEuErZqBusgVVooQSudwFGu12vmqOMCpSfB/eLNJmqbQfnKz1IS
EHu5cR9aq5Mre/S1pVO+UkU4N+Q03UKZR+2u8CyPF1nOGDs4dMrT5kIBFuJNOgC9
aM5QmDXoj3A1fEyTeg5Uj9Z1N0HbY5iy4A6id4LLLKpvJpd2WWfSHHNbmTh7tbEe
K+jLB9g+SLZ2DIMlneGDjrRKfbMUX2I1Z3OGZrrS+b58e6BUT+SzAmkhmYWVyw3o
J8tp/+LtIdGsBOSh64m4trSKMuzPT3gjtglJrzO9ghIucGm4uzPfsbRQKpXRNizm
HQqHCaw16WclmCEDtKuXucprUVzgrU/2wpaGzzP6GOnzbVGeVJ5iTahw/Sl4vTKQ
1dqrOcP047Iy3GaM+88Cm60xX1sqaJ/QkXotN2f5CLoyV/KOYikCc7RPQXdViwJM
fHXCHNrorr7sFlTzB7YOwRbtjbtGLuOI560KeF7Nd4nf/bIjvTb1g+uT++x+5zwP
L40TyRbB5mhTdnSpqzYiVxUwSliYWLe0NQsQ6cYOm4w4mGlWvqW9NH2vMVgftZwg
sqowNZZL2l+ldC0fO3X6PZ7gJbZxK/otJL9ofGRGUgb+CTtcG5rqux1XvX7ji58D
rlbLcAmkCNiDq745AqisDjg+hgHYyQreokry/5YAyT/Bk68OJCQXSr1RBdlzdPJl
Fgx0UZmFYC8DNV1+7oXltVgOBCrTp6xAeI3oYQ2LA6T4oHFSOFUfVdckAdgDmg4I
KYsakChSCOsnubaa4OpDePJvTtZnMAv1z3p7dLCs6DxqqCymEnp/onByWnlCdBLE
GFAg4iCwVfmxIZ9RigUSSm2rYkqliPGHLY9SbBbAQNXmlip/0V5G73LJskZ01gJz
u9cPJXRs1q36FhC8RtSNEfUr4j+l5OyHf2LglsuTP3GpCOvxEDqg+lkvo7TmQuva
dnNDQCty0eCzvw5NDD4XmfnH/KPJa0qXCdEVkAVjGPgKW31mi92hjFhnMb1fwWhp
lWMx5vxcbrIC/TIWeubgqeNCOKvUs+bJRjsGxJQjFZT6R+HWZVxyaf1VtC4fcaxR
hVrWgtG3bo6Wgn8764gfXqTFegaS6+/gl8UfqhPhi+ArRBtVTXYr16zJa1Iy3KYo
xaOJT+EbQyx/KAx5djaVoc93J/hIabon+3ibLUyqDJRM1rZx56XDaCTfNSF/H+YW
fM8F/MgkrYh1RXUpUef6oLhTDtG71KPsrPiRdV8f55NFd03gckoMIcZ3sGL70+Vo
wvuRiFzmFX7wqi60kKIJZW7nEcgwzzK7FCsi0b8T/SY6M0DE0vZcflxaImkc/KI1
IDBymK6zUwZHev6eimH70496OqmlwFpCPtWq9Y1I62inyZqBXursz68pzk/E+05d
X9izKm2KEyucVOY257tarFFN61Xy0Wqwx9Y7CJqjr0vnpoYT0w7jBTbsXt9uLrnc
+1JIkERoba6ROLQWxVDHXZcQx976INH8Kq/Bnj1JobiAV/g1EYQPkdpeGbmLGHOa
w562s1abemOkIIOvnKnU9tbbzKZPbIN6zQMN4lvq8r0T/GNyoKBiAEGq/Y70WMda
6MFMze/8Vjt/jYbHue8toGY34lEWgI0l5eeV2nJzexPGzNVxdbokO4q+Gzqv2ell
aWYM3whloRTlQcp0A+GFhhCuOm/k8NP/J1pbugmFWe4nB2A9XA44O0rGymbKxNKG
vWFLR5+EyucHrY1IRcLYMxsc3I9Fbv2h0rsQyaeVTGFC00ggadXKxegBnxbyV/9x
wbf4DZoaK4LPMHTptELFayOEVu83gXFNgeCIqu4StVCpihu+9OxZ6KSaUpTRTvW1
cead6hDp2M66Pt+dFF6n97HRykOcLm39Jkx7yTjigumwQVbWx7nEm1mls12yehi/
X4HNKDGWGha3dtEvuTj/WbEd9zTKKOc1g6Rd1j4/3xZWqwU4iNBAm6x9TesaijRk
JIsEuS/DMm/MFoWxRwA+pktj3Ei5UJYpIeG5qn5mTVzQEXOowupvJBbK1x5rNZ7d
n+HajvkY8WReDVB4/INxIkK4R1OLgZr3KF8fjbI9MdppIo3ZgDqNsDhdN5IFi/4z
S5Kwai7dwlFdU5aA2VnAWPd/n/NwM1OewjNJOmyYm8tHa7cTTa0lLa6qPe8unwjt
jB6mrxaYSPJhbufR29dxabG/+ZV2mRIfJwWsWzu2HDM2ev0VJAgOipFoDcSRobUq
SYGnp4DP1ujoTSQRVtgXx0kHcPJQMC16EiKUyi2YycI9XGuk6zwGsHUjKpEivVkz
Dy5Ucpc6fj86G5eFbaVQNV5lVCljnAfawul5W4snUshNfDPJHlkbcVgNQkjMZU8F
yXFZh3LBgN4Surn92qO6spjwVk8a6Pwh88E20retqaeC21eXwMLWHH8vKxWN0/VQ
n519FaGHYHDlBvWtm7rMep1C2/vdwdwBAdRJSGlnhtW2KPAQXhCd7lgsDs7vhAik
073XUOZqRFw7oASH+UfQlQrUBjzECMM4gRj2Jf7rvK+BqVvb6l0R0t0yGUunjfmk
pWZGACjXyyjvaQHXI5vJmqSGV7Jrt8+x+v/BoboVRSIjlgbm9+jVAtICigGxei/Y
hPbaLWEahXuOmI4ILAGQkyZ36edp/3FBvKwtTiAiNO4WI42ocwRhaAkpXomdELYY
5jkYmv8KhtxSKl1WHD05VXO1ETVK4n6aFi8KX5XTV4DWxfe21up5rxnEcfGnLT+r
i7VlFCSfBSUXY/yzHyrnQpCuX5Ru9KhgBnXR8WsDc/n81+ByXk2QXehr0r14Zqlq
BtP926P49W6kQ6q2j4ZjVKtpKvYzNUlxeIHV/IoUa2QWP25jl0WgFGwm+RXS8WsA
JxkwdlytDsMSDdEeFRI6MvMwvsrwpoUmbxC6G1LY30oMigg05nXuGtxejWbOTNi0
9z5o2TUy2p7Xu32tBOAQ+LrTSGnrE/8aW7b0A3yrGmClZFftAY00MUzeX2T1+aJm
wZomrILQfZ+2kV5ZZUvg8cJkXXKJCUMZmc68jizDUX/0HROPXhQb4yb8GJhh8x8J
5MSVyPdD/Z6p52zRZ58Qn2kAY52Nfdp47Qlb+z9q1IIfj+uDre4mvSBxojsg4C4T
WEIItYrcUe5VWvsTIwp54Vd8Ne95DmODP5pO6bMGu0lSX2oodySPHFZgNEykf90h
QDpWlbxU7WyPxLapMNoKsJOHAToeLIfMtiKe1N+hd6yB8WcHWxGyXsUdFVMtIL/U
DHPsqdFGJPEi3LJsT4YtcYc2H9fcCYlPwmoasD+PzaSnW9ANanJ4kgFhdkJfWmEn
RVzwEZQE1gpli5B+0jz5LsryVdQUnmyv1dgmaJJFzTlZTMmgx7LS8TlQKmepWhWz
MJqjOmWEqpam8f4T6C9IKaBot4GUXzwX7JN74s/zYJkLwaw9sDeLIvDRR8I14QhH
vC8JUXmWKhyNKOltYz57KaBXZ00ieR90htU53igqf2NOJuTz9tJ4Je7os67ZK4/K
ZCh5JEspr1UGAgSMsCQdSflRBCFHA/vMHvUgxO1WmG/maNMIRODnLOwf1M9SS/bO
3DUSf+PD4yBK35B0PUtWxbDfB678SUo2v8PcVuhVlR0XifGbFurPnnd/4uRJFKvh
8m0IqoQMb2UPlsRZWLI0P2loMimIzkNk6LpFz7gLrIdlGGe+jfL6/9nQbtX2nupj
V8PimsO40q5KPJir0qx40LUPMeuId0RNxQ927vLQ3dBvTLN5uAhjnFWLK0UdvEjS
dvDvTrcdR3pGn3kQpIyRDoSdi2q/YhKUXYqOkY4+w6LI3dl9+dNiSU828NDld7bP
vIinAI476yVbmfMOja2SMcuhuY+E6mgEwh9BZXbqSNk7TO76uLpxEefu93R7mr7r
PLxIjHwJ60e/KW/mrRvt1yqsV9XiX39EihOXSxy67a057k+KqcgjEXE9LVrqeWec
7006th/S3ZmtubhJIte6DOaVfk7988rArOepORbsHkd3ebk7QrBfifxMIzu/OGG6
g1Hs42ZyFrm18gU6/EOY59yVcRXCTaRIzargpcyIydi5oyUghiR02uvax1dzZsyC
5YP03HbnkV4/hvnbLXT6CmQDISRwhQAvguuBKmV2nOnuT2/hy0jhnS7S6T6hujCI
Kr4ThDtaytLbdimBi7zZODLkiCYNAFY+fz/LH9MxP/m7TtQ5ptItaaSvEGeOauss
x0nNy7N845C6rHjz80P5/C0Pwmbkzlwih8VHBrexfW/01iadqB9JNwjhx56nYqqw
hK4U/xO9sUwObf4Ci0HwaynwubzQMkaqkkvNrwDoNLLA45iJE1bGoyupSDTzxnLn
D++IB3qwtch42UMrGnak35VuhQJCUTsBmjiW87yRXj1ovilJGpMyV4MNMLsMsoB8
yOHNMElhx6qNGz8c5N44vUyKuyzQmEBMnyfFtoXs4njjrBgLANboc2Q9GKYIfxLF
4Ccjw1HZPiqDBeQA99zfYgKEDD8RouhBAIGY/mFPnioGHdVrn7mr4td2sfLs4wNj
N+t9mxVicy2yZU/AdmK3UVrpxzEtks6jByEUncTx22+Gl1e8ibyZErJYx2rVrLNO
9QP8sGadSGib75HEnlMjdZBaybT0LzVhPzH8nJMHcHaUBVAnPqPbdGdJr4zzRXKc
WgxHR0U7ItB4lQ1xua614kerUHNdiMUg7ugrsAfPNExT1NYygkvd/hPP6deTjDiL
ZNC+HZgBoUrOlZq8/Ofhl40IszySKiGqIiSv2ZPKF2Hm9o8fjb7kvIXo5+bgJW2p
Uu8m50dKb2QspTGWljLwOF9A3/fL5e7uQlnkptpxF85xfoT/InhtaJwy87668jqq
ZyT0tsjBAe5thwIxp5REjv/NJdjXqbZNNzEy1UyZ25wc95y/OnsH+ec+pzVXpBEc
ZlvZgkWO1Gsef7rgLb3qDukt1PJUKyUwX0JygRCqJ9tb+3HHfHD919/ASO0sQ8ko
qA2nOXsCWwEExsc+MkmUi/AWky93nWpz2xDxl5X47tsxaY68RoorLjHbbBWkkftA
IGBFA8s2aXYahMfJfN86w+d8PeKp6ULdyjh7fMWloI6qsO9QVj6iwAC04vw4j44y
rZsyHXSf96GgTSQ2QRn7T3/amAFZMui4t9xdjuPQZLLzcLOUGgUa9pp1ttlEfBL7
RpP2pvs4tS6eVpe81/srxWJJc8T1VM91ZM7hglbqC+86As7wLLc141/Qn82herSm
vI1V6rel87OZYsRe8d1/3T+RWZr+jKmBcvNA3hRkw+PSTkQY7gvN49zVYJHTyQBJ
jcXFS3RBNqSeiT9S527ZUtANcyS0QnsqKPszXTqkpnIp9qonng6WmyflQ0el3eSu
NVZExepQLpM/0DrMg5NaLSSrR7uTPhPiJCfsY0bzK0IvNUQu46ZIPJ/i9lqqZLU/
tB2qKo1Vu8iGK0CiUhQx+HkuhFiw4XDhSupyO5wSV9gOj6+JBRba6v/xmWjG0Bl9
sRBcDoP90YhwO0CMLuKBdZ6KEwo0CXFDolBzamTegZo12zsQ04kk5BseVI1R8oGU
7iNEpBo2oOEHGIWRFkKW4BtUxYhzBshh5HsMmVj7YzJhxHm/Qsie5BHALY7RTsDD
nkzjOqCygu3MQpsqBwk+mqtLo98qgaKN7erON7YDcl5i8BeCUwxyN3UEWS1SpMpb
0/JBJ9clTksr4w79EDLB0RZXdl5wXwPuFsmS+b4OeMrl6PazDMlkuDpKrtfPfHqq
j5YDQjSJxoW9yQh6SIZ+nLAByM82PGpvQzQV843a1kXiMeHdxVKjK7zp/7UmVP2s
C/0ClQrsWF68UNRRyrvaaAGEWoowvCHJ3zxUwcMaIBuGnsvqFOmDVmnegBhoTlRk
C8tmSZxCD/Mo4oStJRf5lH0ptSBRbI7r1t7ft1ASY/+S8pEkimZAb2RBoH4TdRKf
4sz46AHR/0SaGGl8hfg3bDkOCwBuBaXtg7CH5K2QjZC9HP8RUUdNxzREm3V3NYbI
UlgyGgYQ65fCU4nKlV401W1ndLMdGhV25ipKaZRTK94Hx75SMA6Ok1NxO6F9YC18
A0rqAQbSa1oPFxxC+eXwuXkttlLM/hX4VFjXRaIWQIn+zVQnR9Ofecyq0vE5HCsv
qx4cmVScZT2GFaiCrARVmKwwzVOZkEHbpCWmJ+0U8vSZKIWbyqfJCusMT7YCiJS8
gXTu0k9r5f6wu6X8sJqsZmodUmQf5Mor2tbVrfMxqHVYyUhIjayYsT0BTsOcwKfh
sI0Ga1NPJpmZy3SCmXVdvcoqtSypwiLrmvnzlEb4jNAa+8BQiUgQVhxHFT8eswJP
XfWOJiqidgyhyKXABHrmM/3y+Vlb43cHekHXWofqMhzwFoVyoivSX/TEOSfD47Vo
UMjZQU1TiJeIutCZ5asnGCDBJxeESvLhtQSFKcMwu9WTWsELobMCpii42vR+ONn8
atCI3TtE3HDUxL2/7tPLH9RO5uhpavKOHSOE68WgJGYyFiEj5L8YzXLJ+9XXnexe
6eJWRKl7RDDPlPzQNh4AFG1b7/kofXA7EioldHsjtlMeSqWgAiD78UsObSzjOJwM
SFfhFWGOY5PSkj2Dpeex7U6tM+UYB3gPR55ppkuwGmhCfbSp+L6rG82kOKzoUV59
CRHAXtRxfhxqIDp2hip4Tbhk6uoSw3m4gkyo4PVRvgbaOqhIi878YUHCMLGjnn8O
6UD7B6I4yTB0JachuX3YdlJg0RM+mff5UTxq7U+5ZTdCEAWvPrwHn7AgAzofNymI
ntEbkvzcE9L5kCB838ylCJKTPNOmtzPYjEh3Tf76ZjRm0ou1R1V6XjqZqaWp3dE8
33RiDbrm71yMxdkIY4IvryQ2jaAD9ANU+pBHhEPvtm0dW2936+rRx0x/MybFoB4i
pkoGA9j6gD8FYpOoJTghtvhIm4tK4XtSel+Bp96YA8Nt5Ue+3vSeQIfM0rxGHblS
tjghnMtNzLRLlPXzqKR51EklMB2g4jo72X0buMB35GKOUc31J6j0Ryh6cf1XXk/S
0PEGl+zF7VlCu8S9pmBGIizUBT/uEOHFnEl5JRz23cDsYojtzRHTg9HT8U7OcAnO
HciOzXI8/BJro8svSnnYpoBE9+pc2D30+onWunr3kgGNxoYKkOYgBNmj4qtPk1mo
Zphtskp2vJs0t+jAVEwxHjbO3rFu5SW8TiZM7o1OY+rsyXILrXn/+1ndIgLoc+fX
LBuwsl9/WPZXKx5U30CNtFsB1aiKdDYbLYn5ryP6M4XTvJNc7LNypcjXKZTKxMNv
Q3ReyPWhhghFF7jNdteSXHLCr703oHpqtZ1Es5QBVA3zuCksGidEH5tUjmP6nB7l
GWFLyCEOt2vKYStrtoW2p0844DwUp4tk2JwTGDYgay1wMph3vAuJtoqclzG/8CYV
fR0UYZZZe0URDMSDMyIZIJP4pVgl1BVeRI66Pdgujr7vPxRD2/dKOZPq6b9XtL8t
vlIrO0VyTTlEmfUjPaQeZoXaXjGv7k7IVBWSH0zwi6zGyop6OV3iCocQlvnu6AEG
/aaPOyTbCba9FRHBzXh54LEh2S4t8AB8fZ7ENIgVdYRqBZXHDAxWcBf4ZQ6i2w2o
7crnO0MnUmuU2nO1IoC/2o4R345OvE9ekH5X/Gmq58oLDHy+qy5auSP0s7h8HtDQ
+YlxhmpyXhkenGd1yO3nbiw2DAO4h/SEh50J6j5J11fpfDF5cFR/zhS4COXXIXxu
0Qwli0/Y34rcCVxIIpS9MZDSlemwUyPaMtSmhWyr093fKhkKZ5Axrv0c6crEE/AO
oUeWkkhrb9rkcPRQmGEGXTLSQCKfMHhtXlT2FEnQEWM3XIxMs8j9ahAH3VU438O5
EbtCNE+1auTRtpsmhFUd/RK2DPl/nPx2izUlfAnJbHkqay1i4WkvYs2KKI2oHYQf
cMquPA5G4e4Q/ZdBvAerwHTOiLv1UqgnplWc7MPVw7ZYRIur9jg0MT0GdnGDyMK5
+b6jwdxDea7oYfYIPSe4a67g21xbqg7k+D08mUDleDh8ACluoRSYo6esTw80kT4+
GzKHtTYu3x5Nvi4gyIQ3EfFk22rhFdg26kt+YhZ1xJmK8ulAuEQlvbTA+obItzp/
WM0Ng0+VLPpYfJ2niTkMC6mhjYySTU35MzPGB61HPNBNhzn8X9HK/ctET4SH3o1A
zRYa4jC4kkN9l3HNM8IgCFhtMXu0Tct39mm0JF0X2R/nwf0gNlm81q9rIBj0Qkig
4WtjZBCsWerKPQHMfYNFQBpiLxQi9nNr6p/E+gcO5f0GHN7ekRKxb2FRaTEyLVK1
dMNSu2c6qS8O9aW+vR4Uf7Y9DEjxCuAzvuYC8zf1mwBIgA7CFGQ0d4PbaWVaxxXc
vNOGQ/HjbZnuFT4hi7I470+oFfttvd8Q+QRndO4uA137iFNMDRT27ELdG3+Du9Ys
2MbPIsMhOEQ0u7devWLXEsXw/yj4cQvlLtJbwPBcowkZZ6VTB+a7H+UFiwPYhfw3
9/OVHYCIbTqr+KuCi7xfXp+cofPCq/1VIL7/RGGG7+jHb5EcQE8OSllVfLeeLNyp
VyuCLm7Gnnsu4u1/8Q7A4BlNfy78iDmD41yMadT2xZvE32AZKvrORMaVpLSaDMe6
v14tXOGHKHkAwVLU/Bs+ChZo87BsXyNLGs1lBXD1bwplR45OIlXbs5B+ppYnFaM2
KJpbmrOgO/L/e05Lu2Ln5iu5xpgU9m6wM/Wd7cWvPkj/ywkyH6o08xWM77wTvH7u
lx3fU+W2gSZRYcz4xlgUnNUS9D2TyUQ8ggaqA5TYqc2VY8ynFPaEJ600cnvsAHXT
z5kpYK2LiPHZsZsXuC/hYC7QIm88w5r+3aw1PQvPsrDbQLdu6cOFpFBFe9FkzBWZ
QTYXos5o6mkix9dOOSA+CV1fS9ni6wy6xZHG/xomqjlPjxSTnFKRHc5AzEu367fU
S0OGdDXh/s+TgmUZTsRiwVI9uQK+2awUth5lcFOim+jnJ3udRGGpgNyOWU0RG4Qh
r6NdInFMOByxlAWv9qDp+tfXZW/5bzwGQQBWa9+4ABCsa0kW87qijaft5YYQkyMg
SYBb1Qz9/dNKwRwuIq0X+tQ2qO52hggYY0Tm81riNkwq9TFg1opykSGSOSCEBRAF
YlXaKEFIcECdHjLYekiJFuqQwcm8J2YVj44KGPrWIdRjsnbmvaxka92r8EyNhFlL
HKEy2KrgP4353WxfQODHxSSa9Li/nzoEFXi1gWptWPnhfD+ifiMrAUwQplXGFCl7
SB7vlFnAjC0nkWZP9jx3dpLiJfYFKdzeSCHC9yTK76Ub9yfrxvjSjTJp0gWEkj3f
lj7SE6Eb5bwcX7nRz4EP6nlPu6M3/ivF2F6h1s8yXm2/OFNxbnuFKTtBzGJHD9NW
LWx0NvebKMdTLlgMnvWtoxxXGBTVjXmP7OrlJ35ML8rRFKJmTPW14Z3BlAGQguJJ
ko4gPXdh+ASGGms/Z5P0Cng78X8vCnE4qopQwBqw1C5SV4t7h6/6hQWSkXlBg99p
y0vE4nO/BG6cmrgS4A6Rq/BH/tQwlhWg2cHEUjs6Vo1EBkN7AO1/YlJ3/LqpVd34
oQNzT5r0/pui+Xck8T+u1dOq3sYYt8xW6awqzsPWEx+rH+xHHy0FHvXjhknzul9c
iy2wC5dkYjdGpXcbSymUiWHdEG1Lpx0zt+p0wh2hLaArdqAv0hDVqVSB733FCSkK
vbudriDrZP1BQD7JZNZ4TzSeHvHC2uMs0IsxhOA/1DcNh4bq/3yLvlceeGwOPlEb
dKB19zYscaSwXRogASv2+csd7Zc8t6vBYK5QdmGJJFIYVAqB7GewLbVM4ghc7bmz
Pl0nPGzIhlKmKUp0k2hgowcP5IEbWvFXyBb0do4SiXtxN0iByhWGcjWOR6IKUxwN
pagH3TjUTqkR2NDlilAGn8od81dFRCjKrgMyS3hTSindtgFrEFqi6E/Jm0PAUNBT
mIj0O/bD+L+S1rnLP3L9+1UZ3XyZNqAbwTMz/3+mrsggJA6yoaCTQ5IyAZ3Iw5HT
v9gRrELwApI7bL2u5UYwzEnfizmx565UNUmMhYUeFqSva88nALlBE0mrOmgnwAGy
EFcnkrGH3GQGZmdqH7W6TiPu0MkiG5yN4TXnUn9uupY1grQi5sUsFlXURSNBQxlN
6k31wa6Aer7OeGGiMTe4sQxcWKYrZ4vF9s9Cb/l/BtCjw12G0x5Nl0FElHW7q7S7
oM4b+Ci6hTiKLh7FSDUBlEvaGT0dpdVuNshgMyPso7CaowNDxDzSCiSlnrky7KUf
tuOaTeu9DPQTucTMmWfJEVVhgp+afqtLvAoJJGJ2+9UKdtgQQdH8hdVGyWp9onSO
ab8RRrjXSDbQY5aOQywsvOyxPASmfBmO9AWhBaRscGr/Rpni/JJvVSrp57hFjgeF
7SuTY8Fmg+m3+RRNFYpbyvBvhT5hv5prVfMcpCP03BePU+Bglxgj5ug2EAsHQjGo
5MrIxnYSdWUDkIqKvkFH4q98N6Y71yT4jRsuEd1x5ERm2bf/RMUJC9bTeThe+qRf
WfGf5TxzyrnMIoyRrwV2YcWG7M2/QaBYNtkIJAyUOXR2ZYxF8yBHIOBKhPLmMYoc
nNuAykygM8/Xs9ed2MHHRcbDTu/3Z6Ymq9a36G699Dzan4eWmghV17iu/P35l/t1
ZUGpvOCnXGJTn3nSexniYuYbzOUDNO3M6M6aVQaQmhr0pytlGy5fQkd0mo/N120e
4VvncBVkf82RCo5MN8w13GdjyczwizonnBjydkX1VPbySKovCrKJk++8frvA8lM4
471YIDKNjt6ojV4kI6yfjmu4z7hHDdGEUAMivsqRerQbU3loGkWdgNXI+2GuIphA
QWE3knHhU70J9BE0ZVixr824CFal/bwdrDDEHVFUUS43za8zeAwfsR7fQozTlG2W
zPpaXNwHvnW99GU1+TKcbBgqJsoMNDkq4bjm60et/txUgsyAVWC1AImc/jJcW1/X
XtK41DpHXYbpxmbQ4n+Up3fDYIPbPBYGptrMYe9ecqPA7a82jK0ak/PcznYenl/S
J3Q2Q6Jarqis30Z2VhS+fHeYXjinRUIptRETFWsBG9gFw6W9bMHQudZTthrorRKM
gvgPfAU6SvBtEYnxYXIP9nOMn4oO+WiL+ndv+GiiBfIrW1kdXbZ45GtKZpqNDdyb
0MA8dh7d6G1DeykDXqmbY5iRhNE/Nt/g2jKRP1i0qvMGzpEJlQ1yKV8q1AbXWaRc
itkDBtmlAbFhFitjAdx+KqVWZlGLnrp21Gz+PA5Pbptr50r2EDaZrM/ytbIuOJXd
D2SOM+ZdadX29xYWYXgq4VoahiBB5l7gh0NgGaCMuUnEKhi3vPc1Ade4JasadVEb
0y2j+MuhIhCVBy1NvHnphSatmWnDvYYFaKQ+Ntj6len4BtqjibVFoTk3NeevmLxc
5TF8U4s5ICJWJjMARKr/IhG+KpJc0RxXLjpbLV6dL5+ZRB7iikXTXsq77WeMF7mR
40Gy2ko5NBUPFc71uRgZt5KQgeSUudTx+CAL8prKiVPCtjZ2SdPthH7LIK4AfiFc
HXD1efVGuM+OAKoszD869xjwrMJIWflKoK2sPTl4K80mYI9EzVTxiUhHR7hB5ctA
/2kYoVylvyuCuPUpIyukmxeveR5ZsIhHvueigComXkwPSYnJD3E2ghVPf0mM4upJ
8KqOG/ufAxKNlgfJIscCNSI1QTjkZj2HGcRGd+ihD1oGzBZJfZgwMEV7i6M5G2T0
N0o1Czqpx2ju5drX4VIJPyUjmHttyFhPCnnkg2phN+Gq5h7RG3LA6RKaxlxPJOrB
1qaPrahJeDRtsV3eKzGlvfeMGrC6fz/I7TLJvGMN0DklhZs6ZC/ZMvvdY5fBoEAq
wC3cRJGE7FadYdbemiBTzVqF2p6np+UvZsh+GfwV/zqqAoTH1Zf0XL47V+3ABJCy
OLuzaW1UZ7NssXsggPWgCkFjL+yzvQagCIBppq6c3lvH14BolOFg7vpgj4X6cOao
V48vb4XWraP4l1IqKuFd3e2aDlWgIhampDWZ91F8gKTmSlSXEU1+eXiWPmw7mzBe
wHnK9Hco/3a9zvD+ywmNfhLMZbx4z/SQCOiVYVbwDoRb88KV3iZmCTNO6S0ydO3b
Sy3PmD8AXkzY5XL+9SM40XMkvwNPpU5hDGKOWp6s38Nt2WHnJO8E0a8TlaGvfzGt
t0kQcgh40Xjj7+DgzkLWzFYLLyrBsx07jjHDHSC/D9GDxaEyEnbilToYRBLi+j9v
tAd55SJg4pau8NIsAm6bTSwQNIzaoYNBepIjQUC+mZE2djPWzzAKCOg58sV9pBlN
p4U0mouvMJOl7eIRYRRfoiNVUmIAR4p7/szpAVBQtLDdKKAJVPva9H13RC859Vyp
blEb2BzrG3r4+fGMSkhrgstOmRZ6QZ2YYhfZg2/EbH5dd5nzt+2JHugScnBHIYUx
FiTrMaya2BiRp6WsqvKqY087P2e/ZipdHm/iuk22scBWZGb3vtDqh1zlRLfjNzPB
S0EZpEizTM7PCIsy27KZFUrNCA8bxZnHiO+4kpeJAT9ZtXFY0EBtL+0xBiKihQBn
G2MQo6ahJyUD0G4321FRcasSWxL0KL21bDAgOmYnFD7z4PnnWKv9tg/22fZ62ec+
GBbIZ+NQblougHrAvQ1fhuQUmzflYaplJjf4UWVjSHZdRbE+07AJsiH/nueb84Ou
WYC9KXkElWZnXleehFNu8w2C9rkUQdJtcuVQhekGVcaz8mn+L/tqzkgxau/rdI5u
BqSL5bEEaVJ9zquppa9w6xrzjr6jI3dMIG7GEcn7riSEtu8KDLV+rDcTRTrAcS2x
NHsZ/5cMr8+RJI+/vMIjku1Q6mbk8W0U/46TfIjnIyl/2KYCAO+nUFt8w7den60t
FgBlvB+nv8BeEcMfAL4sHFThnktFDBur0QOGdnPNfouaKTUnzQzLhNP2IDHXRyIm
gBprlJaEDIL89rUSp7f+QhwE/+O7TQgCHgOl37EhTpZNNfylC9qLfxMn42R0H9/s
wGkCgUgS946nrYb0WndAIjo3oqjuJpvvfPY2C7EdckxUTjBiJk084If+6dB/CZnW
YAEAZsNVgT2H2iaLgSr1CDqQam6IS7L253seWrMks39S9qXPENs9vqyjyb0ZTp5/
vISCnCSZAwiSlhqkC5DYlta0+oKW1l7zYl/A8RYYQTfxybiXhJD6UgTKfP0Zfy+o
+MtkI87bEYKy9EdcO6kBsU4zdpuyU+/BZva42ppVTeieOewtU+yo0qQls6V3IJCH
14N2kPmODUVaNUs1k+xFSgtJLkE7mVmoY676bnLZnXMFDJLOhOwPttdHdg4kP3vO
GtMHO1BkuzQ6xZsX6WTTBnxwRvkjqM0DmMrkf6X7cY+zof5Zb6J+wEPr5aBGVLLw
cEDjs1KIbBUtpFVUqqqSb4870nULn9yQARGGzLEI17FUG8+0AC4fmREOICQkuRSO
YxwtMwqt/Lac8QRS00g1kskGaqnr+WIivOQVvKG4bIp7dO4Xa6i4jJ48Ktrh0GAu
0WjyndaKHGWb77xOempCU4fq01vJlbvoi99puGByCexfbvr1BLbOKE8OEWLA9FhM
zHxuMSfLFvfAU00kc3aqB6o8TYuOUdcZiR+6WjbJK/ry/7n8XyT97gI+lJYg09WP
yr1GJzyR2S/qahk8NuSE++AZhdpZWFd3M8uFJjStABtszP2sOXQo0hcz8JWTdTim
9h+EgAJ3qoyM2CW2R4GlFt9+kXIWQtJdnwntDiwe3vkS2IZSRQ0H6ShclNNmtvuN
glFSo7zJfok7yLqc0zw02trN4AYQP6jVxVLjWyRSL96l2girsrqQmIDApIgOJrff
VZYPzBM9kGcJwwH4JPrRdgjCVhYjj0biGjE7/D52XE6ZhFVUJXKtcUUasni4T5Qm
PIzhXa/99ioojUmCrbcydt23w+AvPNrDHnfqvth4EpWh9h5ahQupkgY1a7Z68u6J
bPIV+XsWGWoNG1GwSzFeMZ6S9HNnPT6/tyfvOUAzCUKiJg/Db9il60/4x0DHqwl/
RECRMk5J/CLX0NInnZpc1+MBk9aZO7feR8qEeiBALMsZ6njj2mkgZ0tRohCf3uns
1hjree4PHwenltKsfEnaij8XofujDPKfTKVKs3g+1rT/7wIh1mOTuc2GrYrlnhrd
182PHYVQERPR+1Ik+MdOPRJxM2XwN2RV5J6sLmFxsxfs4mHgMNiV3YQR/KlNHNnB
Qhapj8P/4fIXkGbf0IdCvONUkXQf14uFNT9WfR4N3PLfKOCINXnpLT81N0Yssxf9
kW6WU15MegJJkvgwdr1qjr+oJrQ6RJSabbxckDh98zP2ttoVm5/SlGaz7zT0wRkC
0QxWzyljLJrsHFT4nXjZWRSGmPTOsebfwO0OfCDgHJTk9mZH2u219dnD/5NPH95E
JYz5JO6P3DS6n6nTDdAFPaGgaMDT4xNdPK6J/p+KrslWxawxMnVBMl4SHawYxdaB
Qb+TX8xmDe2oLMG8abCXXzW8qFSfGjHxIHhj6OE0mnAT7+Nqm18HcIfzA2PYbidr
EimsrNKcUtLjNpcZy3i7goElnQ0gJiFP79NnvbZ4V35jrK0yMuvTgaYqeGdTEKoF
3AMFbqyJvRku+mX4KXOut7+i05+iQ4KoICZKBTm8GmyFyUewq7xJWP7SJKd9y89q
F5/YcY1lbvxluX+GUQhfC0EctdB60s6NyypLaaWVy36Bhcajw8+uvqrw/kYQFVrR
XqPqPf203U4jQCR9ewEsim5YBAtkaUkh1wCa2N6BcNGbPnBJJhMzb0vxknMMXeVj
lnHyfonk8vLVznlGhnuCRwJG1opWrQUL+yHiuvW/ZtAQSocHNnhSgcsqa8pqXkzE
xhHPSgTpSs6umrYpKp0YFTOZWr2mOGhY6EU5onBWTSsWcbOGKnUTklcZS/dT3839
4/Pryo4w+FX88lJZIiRCXotCBI9eK35UbL/IcUONWmTRE/Hj38zKcpaSLqLG2kXH
qUutXl7i+9x/ju9e6y5Y1lOO9dUZPlGioXempdHqlMq8PvgG9BHUozzQGmFJsIir
rkUkILovx5x1kfONqsxv+wRGVI2y4FFsteHggXCHydJybSBmq+eeLvlcHCbnsbK9
WSLMSaBu4fOOm2Ly8wWBh3z56gQlzvXw5/gJi7CIpPWM4NXEV+reQejkga+P6Z9E
ykFytxNHKd66UAhIJrz4G4ZygfEWJHVO5/38kPFnEXWQCe3AgC2Q/nOx8akJCtXf
r5rhDAb//NjoF5Aov7n+O/HN/7nopVvsJhbfVP/oprDXftMqm1C4QsGjMf4O4fsA
/kXEbVFJ+LwKveUD/go9e+sOZ5OOy+d/CUID3LLyOUAGlvZdAIJEnySe8ON2tAYx
hF2/r6RpZHPH94S7+OsxQADeTKGtGzZcjGHXPfvVAAyzkWbZnKhzXUReENUOiCZu
Evtsl1ycXYJmTb7YJ3fcywD0DFGB6TZ6Wq7rdKTqMGPcT8L+cOCdPikQrum0HLIZ
lFQTeCXqEx44arsL5YgF2G8cNII5l4yKXU7LE82FnFhUrKpuLNj41SOXI3294tC5
2tGhXnUgt9HL67+DQ/Hvyo60xAArDpmnyRKuh7v8NLi1P4XFgBhZO5PWGXMt6I0U
aJkwFJQNQnOwcGbTDQn7bltW5wgUieNCitbV+cQxkEpP57we/ir50Ymsp2xYkxCZ
fxWkqUx9ik+I3DSVozJ+9jc/zaxtafjaS2Ffnz0RrrSqTj9RLN0oia0cShZqRpQL
9659Ll3vcQI8BkcjPNzQIhIfqlJiH4IVZ3oozwEC9XeIV468+T8MfX+zVyy2dQvI
B5FZEcc49dL0XsBzvnOSJ76mwdgup4891z2ELmt3ysbV8KwWhl5jQMr1lMLADhD3
iH+QSwZPIOqr2M5ysJ83Hvxy2XH9LrerIVnGuypLm2UTwR9HcsPe+Ycd7rVOFi2m
rgAiWTzeG6Gp8V0Je5yWcg+UNGDbczwhqRlSMoTKmDRMYyEI6ehNOtLdLchMEC1O
vKM3IS5bWfN+SiJflcECt4d9aiDTkMiIsu5Y2XfYGKuphZjHLmhrIMgMZGVpbw0A
oGgbmHM6TrMrC1XQTOwyu2CV9SIF4WaORoz3eC+kG+hTqVnkI4XV/QLv/GNqqMCV
nUyWrmEmo2Ybnl9v90A1xJ8FRNDFnJDYollUYmdxldZMJRY1dF0iO3fs0xV5Aq7z
/EzVJdg/3LoJVhZtD+tZ9gc8yLvqtnlS3rc1cO2MzYSyEiuyKkVi0ZMjlfgI6CCA
ytMLnN00gbQsHInIr6CBV6DM5Erliq7QSd/VhdEf9WIDGfbDAR5eceUwPOwLkWnc
hMqbE9D4SV4caJcYUSJTe7Qium4ebfT5hvh6hodFuK3/cZ7f0NOq5QOmmuuygK7Z
BwDgHheyDmWdYc9bclahylhezEt2HTJClURocSHyLQtH9aWrlxMiCgFIRuChX9e6
fb07m1RdGtGg3Jl6WOtNUv+41QkOkzojeh7LeuUhasZqtq8k0vS0QQz7R3afOM6w
BAJsGy2yi4k9c8o52Ee+VxEMnlBHGFxxDDgQhqgjvPV2EtiOXtRNkI+g/f+g9cgc
CPT/kCE7hXrOa9BuL17NzPS+BW7ApKMZNPgBI863sQ3DqqnRdyXqIydWKhSPTbXL
ZpV62BUeJTykZKmop7Mwt887E0GV2n/DoiXvrA87+Az3Sv7b+xTwVVQfFUZz54jM
e0VZuB8HhAJxvmJFaihsTRwvpbZxifbBshXIs7KDx2TY2+QvFwX6GccdjtjUriMs
KuYS6FN8ydD7ueViXG5tCggFBrtWNsy1pVluM2t0qgp7dYYNgV35lZ99+1QMvZmv
AKwp0OVrG82DQ174wxeNNDjzmLOanhJI7TuewetqbW/PW64/tFYJNbj5XQ33IrBq
CzyPq4Zn0Xdyhr0EyL22jtM40JTNL1ctUCOVnOlXd97ZgHmRqPAhEZi7DpX4yryp
sXDJdXndjulFbIbW8/hgcYDmuLCU7c8nKpOFL67Y0tFKxtXw1hUqy203wH8AzSHk
74BoSAdGcXKvs/7CTBxMmToXGjSelLb6tTVlOsI2c+mQrO0KFqtuqzT42cl9rxbE
ob6nfh0BezSPyUw9cGbm7BS84A+/MEWBwNt8nkR2ZQ1/GmD3TrospZrtzwcQhQaE
qUV46v3rxeVK+0bGB0pOYv4FBI/ckMHoK2xgmic7damzLtl0PPVI8Vgvd2EXSFif
3sm2r6olul9wZTajzfsfxcVBO8WeyLhFjW4PVVMUqtGlFQ7ENrarj7EEsYLPG6w+
QTBKxbxcIpdKNZv0UaiHowu9X5bmPVTsoqFpIqVhvvoROMk/DChOXjY9wii6rh4T
kZ2m+t0IqvAIiKIItUaIgzAj5JgmkF75dVSFb3XHee86HEK0MaXHJILKpBtSxt1E
znk55P/ee0x5AxF3PWCaXG0BVU+nNUnaj9eVDacucBknpL7kHH9zqXKkD1npUKOu
A3kVNCD+rTk8r+91wJ8jSQD5YRcikoGN6ErixItCbe6OJrufcZ3eysDXAFnr8b6f
5antWgGrV7AwCx22TleNW1a7kjigIpkG3wYzkQsGBt60c+rkTmO4Kc14BZ8E/w75
enWxO2StkPa3jbuv4NOL2etorG+qU1J3/+sUD0l27TZuqr1c3KM3FX11YGhwxS89
fjZMYYN0jv+72BUscd+GDMqWXH+1i3GPkdlVsC+ZfoCHGJpgBF6dCZA7VAi/qtxA
LSxmO5x6e3ntb8ZxaPM4zdhmh6IBBEagOHsTBH2a8Wp4hCZD/IhRAN4eNyKtzfJ7
b0Z34Z7Ah8Yvv7WHznMsrCVVMIEDhzU6272TZRbhZ0j9vhM1cqNymTRno3FD2dsD
WuHcreGRw4+U03kxn428uKwh7Gqk/rvnzdU84lhZXbYCv7+vz+go/T2QIHNXcXQF
DtNNm6hYXcOP9GJ83XJpKq97UQg9NBdbXnpeHEzY7Apnf71PtBT+VxcJfSdF5jc8
HRKNhS2Rpe69n9pshHx+o5TpjlikPMqUWfQxSGS5RJlZZieipytQEVNGXw0wfwBH
Y1JWD9bENLBpsfplDslP7iryWY1LtTWNs5boeRKGEjIOcbV5WW8qFxamIfhF2Bi5
VhaJX1f2ecfsm9S8rgnUSrifH/AcTsH9+M8qNAqXXhf/xAGMKv98tJZefDfRXM58
7wqKazYToA4/N4CFlf+nHBXBvFcdMMuaSikIWpC5lDagqCO4n8a8o5Ma1m+V/0Nf
gqQMWSci23+vKVGiQPd8GjVb9Nt3a7QZw4s+rCAcrH2oP4umHSH7erzUedwN/Csk
HLd7gI8/u0vtAoGPbqmJ619FPstxcANmK0N1zt4JfFS6AwlRF1pdZHjpFPrrR+sj
8Bb8z9gmG16rCKWU17fb8oPdOqA6V7myGccNYH2wcx+wzGg5o3OdpOQg1KvQ/FPA
HmSozaSkFtna2Jf3g6aQuBqAsl6o6JuuagzqgqJmByiqHrevl3/T2tj+Lge9uSzy
LfQuakwPKu0SjJJZfbYnTKsFiOGk9lcLjWpLh4T/9Qwxdq1aXo7PcSC+qiBD0j5e
AoqjcO+ymdpu7Nzr/+UEcnkhVTt1E/nFQy+kQdzx//V6Vk0qTuozRy7mpPnKLN6N
wNcrr1eY+szrDPmchGT1TJe0kyvRbpD5F66xy+H040Af0fHDeK0tpcq5ORTt3YD8
28vGUykxgWEX8ofIeLumbtIVaMshUYv8/mJn0dpWK3txyuOo1ul+j5pWIspO44GM
whtCrxhcFC41rR7BYCtp2+priNT3jnbfOpiHLjrMUBp5j6QnxHOvu36jlmmRa3pX
U95/dDp1AiFjPv63EX+jiMmapXkrYzBO6CqxJI8dTPUvQakwD+BOpUMHtm1jDLTc
8ipdgakz5Ohwff8Ft5wDTgdn8BCKeYoTzXenNs1fdJPTEiyOb/ZCvQ5MkadMAmAW
i+5d0vfjP4ZrlxZ6qAoVnHU+M72nmV6KOOGQTedSO+jwWNmsu3XTk4HFWYr2x4gr
LBsHylHmFtXd4gZ8/URGnJkTuCIBgnOf4rurVRfp3OTnq9XM6LiBAIj7Z9UeNz/w
HBPJ4uHxsvYx6jBR8NOo/4XpGHhWP6ZKYWpkSas0YDHpxvjd/UNGy+fobUjonnVJ
Y2//0sMoJGKUI6qbX08NEKiCoHI5lpgRYUSamDJ5kEtzm68S350/1IOWuQr7AkwH
YNsVoUZureJGtdM5pz841E7dC3IsMIbhA8F3Qf/7jswb8MjwU+VZIP7gDvkOpf7a
QJ22dCOEQLcvhimhJu2+6RPMPBVaI5LjYOfSf+DUbgqdwV75+T1bQWzosOS95MQZ
QVFYuQHhva146K54ViN8Jx4+t6Z4idkIYrUnEt9PziXidLsKtD71GoLk+tN6tedh
ffnBS23Z5q6REAvc/WyS6XeTfN46s1P6n7xhZp9fcfCWXXaa1hpuLaUa1DBHXCkQ
OHXxX2AK3auaXghEDNZdyrbFHcPaSn6dYwWtKA6HEUpXnWAcIOZZSVRaqLBaMDNq
m1AHUGAKFurROY5AwU9eUaZZf2K4F+9CL6SaX09m89bhrUCZNPPRwwlJBlumKASX
akCWt804s5uWtKLsDh6Ng3fS+E+QjOFQ2taeryBj9Cp27O7xZhORwREBxPJq47Dm
z+j3gJGOMs6tNOU24oZqbVuX33ouPZ6li2l/p/G1nAiYos32aqQW5Niojk7eSECY
XquqykxOuEZ7TDT09V0XOFiHaS+KXBGX3Wo4vgdaQbcNj0k2WUJqmLLgXJXOGaoK
GEPnMvbfAyFdzAUI+lrpboPLxoJC3JDA6q1sA17S8UrN3Blg//Dt8bd1cz718M6N
jyX6oEhasjZRKGl2B55ftbej003Slib4CVN+Dns5vX1t8dfVt4vUfvjYvj2Ifu0u
yu//UOsRgfwxV3aNAsdJFA2ghQOodIFAhLNrxMgMToOuSFI/taFHQQg5JObLsKF+
1utzqz/QPabJ+miwslKHe6OgiLu0t5H16ZT7Ot/QBZra8SzVC5Qu0P6kK/6EX8pi
mC14VHeQxruwXWDXgwOqOhezmBOXDJs9DZv1NToes4uzsO69lUOIC78SJBHvnQxF
ghqqYcztAcZWjSxnppqugdMRPVM8LisFI6TnoqGBekCQ39heWwTIvfBqInhU3HN/
Iv2ie7sCU2rH6vdt/gMTXVr00n27EL2QyNtOqn8KCKPZGeQLj5BMtzWptLNJyUDl
PilHbYOH6FwhbdOduXRQwjQGh/Xi8TA06f6nNfgW6U3g0dRzCT9V5YYJAK5Eowhz
A/yJINMPq5tAHcdJAeBiV0/JMC4MeS5fZZiGR5jXHSX901Cihlecmfwkd/YJqQGB
O3w6skCJOrmZQMcPhQk9Lzyu3+wo4eQd+8m8WGjY9b1VrDqGgRq4wj9gWhKW8mwc
uVMA7FDeRuoH84ygJKLW5F/PNfRmfFhYHg+RxY8h5sL1iXJWedg9EXtXhf0B6e7E
KkdwI2pqMFDgFY2goswdCMaLkEnSRhqBEejIOCqRVYENawA+ykZ9tDVwlRKRq9xA
8KStDbIix6hcOJTiKeHV07LUaqWFwXI+vspuFammNZmyQCJ3/iOqcE9bvrYzZ229
wPsW2Lfmw5uYsmf32XqobTlzOnugNBPV9KzPoAzraOupG8HH3eQ46xLUznlIG6lb
RsUqDgBC9g/4nGn8LIpppT6ZxToiJqGu8p2FjbKMHL3Ctd4Zo5d4e2oMzIw2ttF7
Rm+rpZItE6Mqn91CVE7mno3DhTG7QCNSnKkJwqHfc2I7tCkoTeQtpXqXOg0JYVWM
FzyPg6NC2YxTpjbEzP8wG/UvYzVP0WyeSax3HWFP8O7q82Rfftt4TFNz13ZVfVoX
SthcnSdPeyH1TbwQgWgT2zEowGR2WovJALw3aMz9xE+2EtuQn3pqcE8QEfn5NkPO
qoOHLGDbYjOiC8k84sqbQf+bRKjKjlhd1gParYgg6vK5dntv/HA+9ND7twuyuJB2
lnRiMi62+PHZLf/F1Ou3X4bKlPKD/5ivVFVlbtNXocqaeHD2TTTl/UQ7EOIU3v7H
Mn/Wqw6a94HVRe6d1L/Q9Zd5qcvvySUBggT5fGRwUGAuDbQcrFmzCFrloiNQHjA+
ql+6eUCKYfOvKn/PpyxzRpNctss7OR/GiU+Rw7XCN1ztR6ct5Adthh3MfAquw+8O
AR72L76Rx+ZBWpGlhxD/La1TUnvjEKAlWx4JBCKCbK7zAmUE6nQ+36TFM9ZVZpgU
qANAPfIgD71X7FI6Cxi8bScm/sKl8oQfDcDI5Fu6weF/34HjMbcWnt/M9F102GrJ
8+sno/R8m+/jQLbIvIOAPnahlcFJGPiyXGMzlfoP7y+VUnYA4WXDJyAsuULLIFxF
ecxdpDWutWj6gNX1gUAX6pEI7ZJXsMPJNJbDqacX5SB1hlfjWfH7DAyKOo1/tAT+
Rki66b1RdDm8lDTevfXdV+sxpRmB6afXuIcQUWAeXY5SBrEW2IVjLMYl9YwuwQAz
Y8gVb8xs3f3D60sXB6TNmIkh8go9npjao5uRpsFQkk4qTVucEd0WSgrfZJZEOdgU
W70Do+sirvSnBHAwAebwJeCvWzmUh5fGPm2tTOqGES9+jrZ7aVHaWh5AE+y+VlIX
q90cJvV03gCmAov2uxnnxgBSkqF2QJCVF7DYCcQ6GPCaOzsj6ePMSwnvAX9FuyLW
92DIMu97SaXNP+CWb65DqlmS0x4St7T37p+WS7lY19hC6+up4xjCjLkZa3kyVKfA
O1Yn/268mH5cUEociNvf1PFRhUQOROTJZuG/0ndS7mYt4o4PTnNP1iz+fDMVF+jQ
L8JE/CEq8pRiP/wbOe5NEUnlqk+Razo8m6+CcHqZWrV6EOhO0VRUysgQ0at8H1ax
xnYU1dADIODEKt4RWydKNtNtbHZkcdqbN9OZy6fF0mjZKP0FIYBrV+FKSlb2ydem
3fe14tf7UugTyQNIxF9utMblJkDxBHzdzvA9peokPdmQxx3mQ2Rw3tIUUY+Bc9n2
F4PQWgk5evJ8BmurL/NPcXGto3iPtV/P6St2IeI4Qd2cHBARj22KsRhDYBm1Izkr
tJlLzHBfM5mDRqwUe22fsyiyqCkz8LQXfS3pR32Di0hmIfWE0j/m2Ov7fKjYtw9R
mA8o8s79ZuwP94DZyg5zwlnK6Pnln8tGEpmujTgXklNFHU4RC24428uO3JwKJHTT
8vqvHc57uP5XZ1X0xrG0mbMe5TZytmJi0pfbxpeEnGKH6RW8fp6PTEGSdwq8EwLg
PiFgsmCyYJZFA55EPheuF6DRnDmzVyaT2jv08QelWfeZFF78tQW0Bt2rapQr/lL0
PKBKVlMwrjMQFcWiTixiASWexw9vOfX63S5K0+6NGjZA8Sbj/2cqT5o+1BsAMpZ7
KL4B+D9xEXbXGi9cLOewVuCaoFg9kk8DReRNyS2uIMPQKD1PhUFEmu9bCxgjo5YR
rrbV6eejqxVj4BQ7e00aJwZ1/sbRdxif4uef1FbKchsShqDUJ5Fh04HlLiEWA+bq
coLpvutcO9f5xnpcHGC7GHqblKlYQPvSXSS9prmEIPDQgSDyFaD/R23Ov2KMawqd
nCjzCaXI+46wKQkXdn5VgtjJaB53umnnA0SIrd1HfXt0bUWvKHkG0JZ+a91p59SA
AzZXqAi0sElEeBvTlvAy8TT9gnLeyauQwgxoRARyUVvE9T10FPd6Crdv6YwB4LGy
naKzxBbGOfbJ0IfOc2Njg0+GMtLqc8eWh4eQFhcTP7HUifR1QakEZi87gQT5Y0f4
kxdikmn86F2sLwSEqqgl5SUL4LmNIVPxh9dybV74QfuL2yw6wxyb/3EE6d2OZTkI
ceEBGKe7sEqy+nvsQPKYBinKTSUoR0ex/tLjeWjEF3Dn6aMhF4pXr1e0p5rBb1Bw
KdlNoE6bqtuiFiyyyeMw5peFwtoHuk71jit6acKFF/2u1lErwohgeZXN1R881YSR
RO6ThJsy0SZtwQuEwI9OVYQ0DOKwKHYAqfwb8kmFCJ+GxCQWTLL6sND+hnbgM/sL
4Je7WOl082sBeaO+Keba6XU1r3K6sF5DBwrcsm9ODNdF5THJxgBCcUATFGcqsyDE
P/SKmm7BSscMWNwPVOiKjhwVqow6xHsnfY5jX+9mxR+nRipUlG6RSayIVKyCgSyZ
3SrbS1YssF8IkstQjY84cRf3Y0ltDk72Gby2HC7SRON7GAkiYw5ihTBmYwIZru+Q
G8BnbwAL0b5tI+dGyiTTM/bZuKNLtCJ0bsrrr6EwVHC0cmiWt0fS4U58QXZWmTsU
whhwP3sCbzx+GOz4+caEiFGPFUr0TGqY4RuGwHjjJZj2jPVVpgwv4NQrefhqPXSF
4gl8P9X89Luz49mYnebTT+BKBqmO3qSBkiMs64IkZjXcSkL+rdsCSYtQ5tqHjYf+
rCVkraqd/4uxnD0/VQEqCIDukWTA02rE6cSo1zXEs1x+WdonQxWO4dgVRgr3cmMm
pjg1y+Dq0z1oNl3w/O+7iwcwqLVM83fxGV1JRiolGjfpqLScrCiivRsCMPkzbIxP
GyDbYN+0ehSSrZhG1ER5W0SGDJ00Dguf0rvCpVbtIjKh+waLXxdOiNDfUNPtNi2i
t1QWzmMX/ErrALUxkJ2kcIyqcS34uArMeNQCw7eytSr5LvtECUQ5lYL5Q5KaKHq4
7WxFWURlYP4ekz8/G4dJQFy+6KoaArs12kLAdWTHQO706WpprYRbXxMlZhHapqkO
OukEfVXnrOQ0fJX+q20YpTNsVgHHqmJxEENsWLQbgYQfVm2edN1fOk4j1n66AAew
jseY4zyMx0CqVZfS96hymVLQXsKdNR3A8BGqAnSDfWNMWYwml2K3StHY7k7WshGe
8DbXj3a/pLEVYXqZMuaOpfeX0g0dert+63Ie14dd24TWJrlI3vUHkhs0Hd5kk31z
qZnNwKU1xADr0IPkJ9EWo1OVbQpfu/pyrAgcbPkawzUC4Kc7GmzQ5JOZsNjVZDlC
HcYZJBImMSx06n6GViHUoX48cCPStvt4u8jyq4BOF1cnWQw7PR2kHInlA6nJzsNu
weWLkOVHILVOwgTVQQRnkECnouheIgm5AQlw9UTStH0C+rntzcTXg0dI/LzdIpkP
oziizxOf8ZqgLZqC7j8X4nwI1LVOm1ydGEh5q0oUslPGwdfB5sHFVyLozyPMaogh
wpCPiHRNVCY/ONmTI7+JivnwPVfEH8BmkXTUfj7sX5YFR9ExAG5/I67MxtJrrf11
KcSh5d0GXvfJzM6cBYd1WGH10FNnn0EqpiOqbTgJ7HIDU+8rlz8tuyIdZ7plWNZE
5hltYn+++YLl5h56xJL+vcZZd9cS+AIQT/SXz/NzgqEIhs6vUFCE4PTkC5zoNBBh
8YVIwIwPwYELrPMCY3PbwYCB7bMDU2yIX/j7+5/9F/3Lkdzpc9c8uS0Hsdt+bvf1
8N04p5kCPxlo+QG/gIlohFyI6BuhZSnIGGYqzr4oKih3sLecvv+p417M8KOWUyTb
rNVYEQ468SJAK8h93T3PyXD5D+gmt+9ejidlQ5HXd5XL65Wgjbv3zim8E3UuW/16
uAFV2Cno9g1fNbcZJasNXqCrjrW1QN41AnREZMy40kzHnWJZwp93wzW6UmILkR4I
/T2h1GxijqXI7u45OY2PrKalWerWSAOx4kDPj6q+kx0tarEifzCeHAK5MmJ+LGka
Pr08z0aryt+1T+IGMENSJ93nkB+mQOAvaDu2mZi3UlB//WPEjKhrFwuohDPe0sWX
qsBGtU8ED73FIvnifTwOCpjofM4qjFVk9yP0gNx+c2VuzfTPbSff6YFbAJLKubBs
8VWlk9ZGwczEIb/bE3xI8s7zeuX98KhvQadBJVtsmoEDkyAEJ3te1QFjzSWm+C4f
psAg2Vy7Jb0YQaZBiLN13X3KnMPdeFDlBk4ITfAqjego13RNJ2Cn+7jLLRzvZlIi
uT7K/eqsYMyU0JJStXoFoLP6FFUyuGlDO1fKevB3KjrRCSWWyPMTIJIfSVMBYUnf
20ezc3Y2We28aLuHQAutLzH/ZTy8RsuKeht0wHSWzds66fjj4DoxfYhBmPTTP2B6
K8h6Il2332uzTzGpAVHvz1Ua6G42CiFnxlVjMwQmxT9C5kr5gqQEDvL1sQRecyPv
/chOh3jTdeibF2t65UlwCJvZcBP/dfjmXRa3ocoJb7wb3SFbplmhNJOmHOBvUH+L
nPaRnQvWHDqor2l9nJ+b1ZwwuS9czICFAJ6OImL+uJfQ09Gar7zFGjh32qpE3CQn
5LYGKS6GEBg3zlZtxrRvzvU8xwWvTYSQv1w4bvE7/v0UzkiSRpAJ2PETQiS0i4ox
KmRTFCOpW/tV5TVnGB+yoLj2BdBGAfl5om5GQK328nLGoGltbEXYkmiIpxFhqIgX
p/M4uW+imKZ+rt831wMwo/LVlHImWsaTVHcGECZOG/Vbmf2zmCzXZO46U3VyrMKk
krh5DvD853OHWErIbTQS6FSs8Fble8f+nwms8nmOQs0pDo7p+to+DW359cMvej8f
wRDhComIm6fbmM15RtrP6DdtLmCEsOPKHRxKt11CIXa9DxexJuts9jCrlSyxIId8
hx9jrt/QCEdIN5ektKoC4KqcpgtvPipeUTAYYY9YvhYXfS+RKypG22uaWNIxNRkR
rkG8k6Yu4GblyC4uYPZsiqyYIFXVxzGAWYajEP+QL6TpmOI78mc0gRcLcNfOJr+2
1/u5/V5CEVDjgXegFG+Vq8IeKIxNLaRn0hrwU3a4b9QT//aSTM0HUZnDEwMIXTTD
KlQywLsCIQ04ialMpMjOe3+OCRDzriKy1AkYvy5sfKlrYX7pNlDG7Rq/xWig0hy3
oCxiRw50NTbsfJTTTQCWQ03lybi7BF7D7r7mJhDVWcSG7pnnOffhx+5mdN9j+M/5
LX+jIRJuV1BPskokAhYcVFxdYZGdp8xE16JIo7QFb3iykrGuw1MVhC8YJa4pdkOp
5+/C5sU9xBZB012Siq7bCAaNGKO7YrGBRtrSOvlsJgDLqva/1Ct/nwcyRzYiJVPT
wq2XkhhWyI6eKOIkfJnOI3DU0dBDF0xEym5iJbI97SSV8Wf4xPlmOrfg8LDm3z1E
FM9Y/RBR2HTGiEXVct+RfSv7eF1V2tduOKha/W7kzQEsBDeF3levkogGnn7PMejm
sAXxLSZhbFOEuNuAhWoSPmOOhl6GobHgxNEJsaRsjuk2LxCgHbkVoGaxZNZeAGlO
4DnZdn5COtYKEskvvwtIRkmr6si7TOdXuOO9cKSohpIXv8e5QVbIYUOmo/gsu0ki
BN7babfe6g7GiMONAGnBXYVyTE17aMRJJ7TZWl1zaAtWFByqPj/rALIWFB62JKcG
JhZHpBpV8N3lIBkF2ksN6Kk6pD05v9Pn+/iR9TeqT4dI3j32I658w32t7xOzI48T
31v11cVnR0RBTRDPAIslGQsgStH7uEY+sZuzf9AeJxkkP5o0FTUh5GLWMxRgNXF5
GR6GfS9SmUg8Qn+gkkwxwzQ4UEMfwz8T92xES2boJ4dkwg94TFgxMm0/HbDFcBJs
vCd/YU4t7ureoo/yX0sPyS4zpaJRiZuPO4ZYhZrx/KMODp8ZhnxRwSGFZ/aD1aj6
NRh24vtu8lYQuRNN5sV7TIux7Wc/tkt4GbZqkXvqfJGHbL4F7/9Wfl+AhlN6Fsrx
sVchjaGbutOUTBsqNeNxupp/AzeGLtNAr24aHeJEjMoDBbs0W7GHlFJ1XxKij7ny
e+R01c3GQMN9nMwjTuc9EsibE/f+9Gx8kmaTbNCJmELMJJn5lScH9prsIn9lOQPF
C/T0OVKR3IsyZ6WlchOeul6P+jJqyVsczAwfJuSNEWU66SDJZGw2Xs2BZKZcVaEG
ABSN6Kl+p5ZCZY+WU5/xiCA4+UB1Ij8lbFYkqeR5KgkKPKxdNQmpNVz5nDJobzXF
5gGp9MET9S3q74huWWxsD1v1oleftEymrlBMGj2WefBCPyxghliX22YwyeG5x/dd
JCPY2cddHxS1I82Fr235W1xIUHEONYN+raykSCpLD0o33WzneoqWqIuK1gDFF6CY
PWuofGGr2c1JYJf3ZL1zWLY8hkwSnG/nVBVnRpSAg21iVGj8oJby6zNRbLD5y8rw
tetSl12kEc4E2YlBS2uz2CVXkPo2vVkjPwT+Tbe8JpQBhEPt6q2f6qvDofiYtdBu
6t2+7ozfEpPLOoJknHz2wNd9sqfZYTiginQYJwvrplKUyIbPuGlwzt4hKfYGbnN0
mbsv5TFJufu2ApsCdD1SL26LHEmomuv3WjWpTB7GT9t1CORzhujvDXFrxzr06vua
8REqUEQ6dVtIz9mt3HfGEFinMVwKzv/qEiMwYAvrOFJduyMBBShnQgdVszfI1qlq
3OmNbjOWF1DhMO51EQG+nNbKkdrwdryY3XqkX1NbhuUUSkgt/QqEZn2adQvt8+lk
ceBwieviXOI55h3sEv+gZjST8tgeZNofDMQV4IXL9DYCkNuKloIVPGgIZHpVxf6A
HGHatyzgAQbocZfMa9Cy9dBmi7edB8wTt6HCUH9MbCu3dWiBSRlAu3INbtTW2+9I
nmhEG8lZmVqm0yFr3+q7vngLU9vk4JjjFWkM2r3ZOnfM/qkDoS5jXRKfuYSH3b5z
+MRCn4lwXb9/+aGMIlo8UX0SpHj48oyC0fHPxi1+OhY+dCkG3RjxFnhdsyONbVx+
POSKCHfVdD3HKmGyDY79UgrsorjDPs1ySHycsvnxztEg90AWbr5xeaRHrixS4gMa
ObGqATHhWpJ3D/hSIw+4i3P57FtSEE0YRnSMarxoPMLQkQjCBXd294moJZEO5Y5y
dQISdQVjTdD+estBt5kTi/41M/S5YHNUCYqLCuzF+GPAnXoTTXEB7YFmx5ogqGSS
wuBuAfn94x6/5mZ0808S+MguZcvHmxMnQ+9+Ys6lvPg69ZfJsIiHW5NZ+ffyRWap
/Wo6wjwqwdPeKEf3ni2Q8GRGgoYvJlW2/yHLwenRNtsqELP2UsGNTdLSmpURvrKe
367IOMLhhBz/ITePqqqlIMPQcNCQaCJm2fKbCHlOrGRi/YNlqbbP+VgGjNJgb19g
jw149ehkBdAjyCUkF7CbVc93lJcfjz/Q74GSzv+1HCyIiAAexn/Pp8rurzvBY1Vu
AT17vTd1dGvodLiFcgFGKZ1VMuSlw5iV/7TDeDNguvHlHyJadRvwNygm0LXZTSaJ
PbTBXaDhSH7gw14yYOcqmr4Lw6w+xyiJzGWLiabvp2WwhLFhYOSDeh60NBdwy32Q
M+K0hg5YRU+HX1j/EPD6Y9gxGN36RtDNJMSBXhDWLeW9Ol46R2u4CUIFmD0JoPsP
Us/Zd0Ma6+gnyL7b8FR6pCMJXu/iC73qmbVu6UV5UKIfLO+mEOacBHW6QjTaiOoF
chRy8sfT+APg8AzeDESvz8Nyh9SlDEuXEFVHnE78oNqajDO1rRZYd907/wSXUx+u
zpkuzMHkOlaaxc6ahyJXb03urbVnX+gpwZz+Qjn4xYhHeEWyT+X6f+FuPbIOLfMz
tSqQKCXftQcU350TBQMkpV+lNC5q5WOfPhlW5kjhm2ZT939b4tWY4dKi2CBJxBni
QkrMd0AZArWNjvV6EO+QLnSkeRy6cCjw2RjwlkGXCAxT2Asy3oV5QwFWXrfzwr8G
owBpfnhac7zAE2FqjoUINL6IwU0BizIHM5fZj4mG10hvKgWllKId7YAiTcdpE2wQ
GwZPqFwQ47qtRx+ucugc1FI71pP8Zy21ea6RB4BaUFfVegIgv9dyQEhSahbYpml8
30pBfBb8tXWG73EI1Ikzolx1wXodK3GLCjndAusb7jM41l3LGcTCQWzm4GdjM4rs
pxip1ddlZoLK9NWJyCsE6a0oEZU4BMg+Y8FcuGUH5+DZ13JRb4mLBZHCzhMYKmhd
+UjMW121+PTJa9G4y8PLh2jiTWPgEeOAgobZTeppmSicQiVP7QTY6PFfr/BqfaKP
9GNf/1wnVLtuMSqeSdOFRdXTYSG5F/jbp9OX0dTdO5h83xT/GmEH18U5EsiVuxSq
8YwzPntZFt04UNmAIogvEYfmCPClN/6qvK67QDVXBC/S2tboUwXbCpb9nZ/2hJE9
1qeBcsqgRwIXUMzYr08Zu2xMwmf1e27ZfP2QmqEowFoftephvNi1njUyDmEKQM+f
dzIG3T5cchpDM3JjQ8B4EncNxAmkljdg2Uba23fiIz7Pc1VcIYFIu1D/4BTDJLrp
+8gr7kNpGus5vWAJKH979nvovIAOcQ5gpc9sCsi78geLNs//xSY8fkFbsj59opS2
ettGLmHsD4M5nluWJhcswNeNFsjRanJxul6a1No619e4GkTkWgd+xpT2bB5diaZ3
4dwfr2/GeP1g8ONpaFw0fuMsGI5uBTlV+y3cElWHrZpuZkLtSwqz0p3RddGGM0yt
+/l8F47FtHkGMZ1u1QzyDGVGDl4Eli/1Ej+L/uZ2qd4KsIEQBM8BiMKSxrqVNCcY
1NVsqihSVQfhIY/okIP3Pooi5iG/1uTXQzQ1FqkOx19nkvbN+wjMDnbTV1ME1X8g
HxKMGfEmNVnrLJtV7DiFxVs6SjqYC/OAcHXbdtRgOgvE5rUHo+MEcbON6xdaF5/I
lLBqis2EImPHuxk2CY5lEAnHsKarJdpduVIpjWnUA57moS0MZTprki8dQQqHM2j/
zqDp4gVjitR3BdM7BZfZe7vO9P2F64T6cINmp2vg3UnB7Vbtc3zuPQuOWAyutRT3
L4BS+9SRMb5Md2Rzo3OOu3w+lfIuW3YEoW4vrzSBG+Kv9M09zLe6YdgRJjXaxg9o
Cya3shzIOZaRdhTl8UKFYRSRVdvQ0fmCuArI4yUJC8fHmAExH+N1Kd8WSdTmZLgO
7POZe3SHAzHtoFH0NVDIsiWczz968/jVa0yEe3sFqERWA0xbkcu8LyUAN1wzcjr+
3gsRijOYUwf7QkL0TK5A2BStluJbenMt0Hsip60zhhlGQX9lxdz/8OoDjA5xfiyc
4tgCKEKpnScXQ+XROf4pN2UGh1mnH9uj+TdcCKGowChNhf5JVsmoHEI++y7dqrZ4
Hh4O0O3G8gGKGpn9GInCuCqiRuRZmp+BtLaG9T+4eZofYP4HjrDMI+uvHMyBTHD5
HOgob5t1CPTH+JUGByZQClIpoJGIyCk+3qG6K/4ApSXmvxHJrXi5gijfU9gJ+L9Q
pQyvoxFqWpDpWmjRPEmRhzJAWfPHURQgG6ymJOceJCgDkgIHVwl1F86evAL1OahI
LkR+/+EyoGjiMAP32tUjIiT2G1mrsjjltwQiWSDz1mfPQqm/h/E+Jb2KgaMZUVT1
McvmesgF06PSKlqDAJVJHyytrQMoweocf5cuFyMjaldeqp25V1Yn4snH6ohjj8+5
l6AhBCuaRvVyRR6IcYd5SAmvgD2f4R59JaVR0A3FJYi/nMk0P4c9C+Yn20S6HULC
+DdNvP9kyQaYeVJOsyVLOW1pF0u5IODaVUiarr9tNL68kj4PXSTMPkpwNJvaJFq5
OEtcTMy1kQyqxrI6Yj6/HtdoSrCiMe01MunhZqp2adt1tZey9xIAZSEKKC0LKghJ
89+5TnGqcsKeC++qnpk298DCJg5aFxqIq1nuZzCUkOiKb3EVilYG0iiRawWg0P72
Ze22HWInvztwXH6EGQ98e279nnqXMZ+KLeD6XAbEwkpJr7X0Pa2zj47UxOgX5E6C
D8/xdu003hnWHaRpmlDQPLk6tJVw2v40uVay7cu5ZHcYqgnxyd4/zeTSIbkaZFHU
2ycGzd+6li8BnemR983p/BOSEeDaQSmnYnGfZvhnF7j5SW/FAKVLZXB+AIUW0BOr
wcwaE/P7se/myRWcJp1wITT4MGyUgrHqefPv/ysGLD3FediVcK0BtTJH2cpvlgHa
UJh0fCs8HgtkE24KIGt2GAvf0E8/4DdjCgRd1o8bewPbV4er7YGQKLC34kDg3IaQ
rl+ETGv4uLlQ8m8Vse1TDLAM30f2Z1nhfMxGpZkIcDauTFqWHk1HmN0CNJVFETnD
Kt9l79wjlpRJW0HiIecMw84pGZjSyuIg7go5RuIK1Q5SPQJAZ/cZjDdcUWGqKo29
aVCcnPDoxflUdbmRHdxecVwxJ+idsaYGyLgb11r67l8NCdUYs71LQzQ37kARgNzk
YFQWD519YzKFWnCVb0ZN5IRAhTZeDnoyP+1UwehYTsZDHdFPWu+8llF/Y326apC5
yyRL0IHQASupxfJKbeS72kDG8BYNiZh/7RM9k2pO51s51bRt/+HeY7LRWZRAwlGC
aw5iolNXIRh83yawjn41VHBKYhfaJSBTpix8nddxKExS0kpMjl+4u7T0olL9ICJA
2qHGmvvtvulSYgjDg4/Bt69c7Dt/olckqxedTWvksWFSxTxTpU3sTq81KFJDE2Ay
yPXNPuFtZAfIhe5ZnE+2CXmC4bva6WU8fLD2SJPDBqf/vrKO6Xb6WCKMgwiafBur
NCDFDr1w5x7U16pFWn1oYGjzoKQDz1Ohl22u3MBXQJpw16hkZrnH7lRtGVX+s5o8
a12xdbFOuin6BxpMXpjl/edqH6BrlN0xbv/KRPYbd6r/wxCoMjDOc6FecRJxATo2
gGLJGgzQgWhyOHqeT4+ttk0wtmcOXiPsNK3/G8VT9al9TVzTN/5SQm2Yd10huwA8
EKn/CB5PNKJGAB/JRCc4KanFUdBnvt0yu3tkCmwsQ8GyahAo/N8B3b/29AY8Jcnl
nPDH8ZAiMoDzzQxCj8bf4oB2iA2X+p+ArMd951E/ogU18uAlHq/Lbvy/cmT04rgy
FJz3FmoqGXwohpq6VK4j7j9EvHWralEhGg8YHfJkYakOHs4F5li4m2Ra/RjiZfwf
KgvkAAlyvnbJ//A0VRiPyz4N4LcQPvGET9NloBvK1OXPGigMLsSKvBAzPbJjHG6A
wVh/bxHAcwDL7/ZNEdU15ohTewH1R+EHdGol4YY4cqw/NpYBQyi8UBcehDIx3wqL
srTyLAn4kuNKIM8XhRbqdI7kV+X1Q+pbLhShoyOnlmlZQ9vE97/7fu5eO+YlsQtr
d1zhL+GKZRJJcL+fNd0a+nd0XDHl7AIJMRtWjSMWbQsIgR/s8LhNzhPO4/Ddg7yS
quHgHFR/Pti7C2aMzTwUExoLyY+ID7u771toERKBXqSn4lIVpuWAhfVOEsN7DL/F
8KLhWs+j9JyV2/bx9DR3nFuYLrdIvkhyjRR8pmUjC5Q+4UWUuaoK278hDmAKKx/Y
XLkQw0CI2EkKEzWvMrVFyj9NhWAMMkcfdmtsLr9DY0oXfX/HlrsWy8X7BfcJDlAp
Cjcqf/hH9l0ggQD5XLrlPl9mM/5MYfJGEnoAzjyjRaaDOmD1b/1toGXeX6dptOh6
VkZmpJCLZ2Ktoqkn9Vvx2CoAFjSa9BiwZ2KLWCfYTh3jkH+Sy2b0ZH2wvkruDysP
vNEp4BQigE9kKDlcmwsVvtB17sm2RwBPrPw14b1vPKKvrcR7gvSW/SygL/12baiT
XLHBZ43kguRIECpqGaGhtK1piiiMAtab9RLrtnUtYGDDthMCU3d2NE4az/MowvdC
N1srEhBaC0wXyubybocu70PkqgjlwDJKdCIuZRu8EyRA43E2CQw32K019yOA32cN
L9FXoSyKkE9D3c7qdqPm0X61pNqvZBZ+w8Jk42G9UI1TfxMyxLq6MZyvcUwvqR6S
OedJLJnKeCsTuJsVOxXqtWK1UzQwUKDkr+CtnnyUacNKkwY111sZCk133xs+0IEt
5dd6roIGq0mtqLsJGZgN1YHXlhcea6n+JAlqvOtT+2BVOwrdQ2WlWaFm6cQL/pWS
IYCyE/bM5ilNgS0PDvlNTIO6sRcfRtaWFLB1XBHX5gzf5p9d3JKt+S5YIhJMI1cs
KDaxVmHCOAg17cA94vS+V8RmgEWzoGE3hDYhujzMBBZdHUb0dqiXwLgd+tDiyHvo
dWLaj2zWZHyoD5AeagD2Fcr0h5G+qBFJ2w8qUGqIqyCj+oqVMrMNPtHegGh9CT3B
xr0KUUAex5EVqx0WucnFxHk4RPQVsFFyBJ9QU3x8C/U3d9ysmuEzAd1MCk6VLvHH
2ZzsRr/6CZYvCC8SVWYgWMNvwuuY+2DTe2+7Uqe10gpus/ZB/TpalIPc9unqR5Ou
pVMxAdwd7VxJ8ESGYSLf0PUUTBRh2gjgSDd3zIh3XwgBsbxoKx/fyL7fAcBahbgI
HEqeTLMfHL0dVX3YlziSZbUx+NZuI2w/iUmlm/LIFOx4ufrNAzeYxz8cU8uWBBEO
QNbI/EZf2u1+6k2ZOJZrp/4JRP5V58z6+fg+TS88yMUTiQUx1TsJhH3JHIDe6/S2
0tmolDrjdA2aCAOeejh0GfnACa0Vx/iRWh9UPmAezK/REuq154j7/nlSqAVfpLEv
ed7lGNDw0toQKlZ1yHlxq/gf40E4wtQFBmQFEOuw3yD0BIgEr5+EfmMXS878Ogmd
5oeyJJZK3P5Yg2xTJ60TTH3SqcLng8VXfoM9X8ow4oLxfOFg02AwmQLhbnTF7O6x
lDO03T2IDjQ2SiQwf9RhQCIxcOPTerozWYe04ZbkDFcPUTKoL0pzyqUXpKGqAUFl
RNHufhb0fa+/zeD0s2ukWoTpIimqPiO6DwK8o19AIQ4sa3+nE0JxQzZvvQMdoWQV
pnXZpl95V9QDpd8xyx5pnRA4OwpM3gY7wYG/SPj+he1pGYCYBfBCA9bfVW5tDqH/
oE1NoKs+s1jAX/Q8wTwMniSosH7qwPd3wpRwAe7wo7preDntUvxT0ULLRE2ILaLl
JDen9888A2BmZ+aElJcuZED/wzyEXxkVKVQj3aKERjSu0eM6dD63/wE1l8U6hxCr
v4/3UUAsWLtVaHIaWXdiLSi4/V72RpNjeLVpDTq8IQuDW/BIgRlmnCN4jduniwrS
rXZ3Lk5rMeWBy2R4zmTw6ITdRdIB/6+VSvkV7TUNA6dm/b+LhGK/KgkTiiRDyfV/
lzL3DEkBQIKodpICLzXvFq4b0pJDnX5GztV8Wwjje2w0fCdWeyEv0cHdUTYBRGy0
ui4Q+uWaBjT0V1QvUCzVOtq/ws0CgcU6O+T1uryuPMOogR6PDterL2wh2704BRWZ
S7QZLADn7huExGtegsUZwTn3YkFUV5WgG1ryuCgozSpMHJotKcpsCagVfF+avS6v
jmpBHv7g29/wN3HWiJrBi1U8HPZLJQK6T8pXW0VmuDCl4cywrAVPsDOSxcmpoJVM
VjoOw7K5DNV5qAUR1Ymn9GlGB6BonHu8YGOAdfKRuYsVobfGwrdVLOZ5yhz2mKsb
+NUrmAgfYpHdig/jOK6uJzXy8fbS0rmgLj5WXFCacyHxjAqJnSWgMR6BfwY9YIMn
Uf+zV14jyS2NfRW/slz7zJgBiQSioJviEIZJFqkFCNQP/ZU2MmZCiBGrj2tk54L+
gDhHNB2vJbVLujZv70LxtYQyv4PaSaomowO1skmN/O3tVHvTzPizy1Ay1uN7A5MQ
jKRyrmzfcGn03KQWb4rVWDO6I3ERhukwbG4Jd0zfZeMUeq8QVXxAMQ2UfvJJhp6f
JkJDZZLn8d8YYPytIQOVCA3E7DZJGp4+CBjQ++rmwXUtixPxgvHpUdkBfq9BNkK5
V0IgN5fSfp31qlw+JtRb5srf8bzaduXiTtRZKWnobQM6MbtZmnzxdnaKZNBI2jtV
uvKOrHCJAIOXpKmQA1yKjcESLCUFnjnSqRtY4Qn3eKwuKZnB+1uGaJgICcCyk1ug
uhqTIy9nQZhPtmusl9YkHLZCLqg8lodo1NNxcglyDzW5XSueXwkizslR+D6fTQCX
Grsh0PV8Pvf7i4ZiXcvOb9EzCTan3fyNklcbVFoV+vMqKZrWEWTJzB659lXgE9dV
EDzT1HhMmXql4O45Djv39UlCG1z9WVztj04zoZbptPRzinkbVPYFb6gyu7KNT41b
RN96SadRRJKLQn+OmZW9HkN3hqY7g++cnmbyHJplNSa7h84EOomtH+LEE2CPux9K
wC9Jv7IGCJcg0UL4CYucyp4Bt0G/sGZZ2bqCABBkZTjwtxSGxUZNCGxQov2SK4Os
Jrw/32KCaIGQ9Lf2ot0rjCte1DpNfikLm1GD2vk5Oyq9GTb3HfbVRkfNOQt8Lq6h
R11B07uP1+ncZZa2snmer6Jgb+fdiSkz35r4NqpfJKidsUbBUCtCaOAzQArmBTxb
YeTbmynXNtuol0D6kL206pRzmuADaw2WrmcO1iezJzdY+/0OEQhHE4FMEGiAndNW
M20YPEsJADu/0gYjkFgsJSHdS+TzXIJ27IYEkyP4H75fUzPzLGeVmBCodq8+EBUX
QhIOOpo3wmdnHaQCVlkgIVGOyFrLYZ+ZkkZA7exoRGDVSqBZIKvCsLOef2ba73Oz
uHRorYdaFkJexfZRYj26CueJXAGfVDNB9rV+DD4REaIbJNHdzHhkLN0Zq8S5+zCm
aoRpZiwDzIp6ISjcBmS8WMbbZSu7z6gGbxXSk9r2jqJLrf0FV9aN8S1Dm+krem2/
zVRXhd8TG+dQYUnzdujuubpXA0P2k3tR1zEQ+olbYDC0EQ72RIXUU4CgWIVnYAzY
xe1tIhEDh3x/BzmGyjjHtpjRdoNL2vZ6fpMoNnWyjg5zerCQVux7r6gaioelps1F
7Ig8VeYgm6WIrQPiLf/5/Sfm5aJq0jLfwqmI1RqbpHdj2hAnIfF7A6a7WbzzvQA+
qNn7vCrcdf++qQUV6pBiiqkYfHnoFZ2TlL6BUEO9eyKA9W4riRpFXOhXmgwdzMHY
V2N23q8wk4z+BSU/O9owKIrd6kwl+7dBTtmFXKUHTdUiwynFePreqRMAfSMRhrsm
6aLTK64boXc6LE6hUToZUcYamSal6hHC5133HQ+bhXMtKnTHNwQLZnCCizRGHCt6
kjaYsMGC5pj5wvXBE94hezBChszd4ypJj/LXfpGKg66e0YtUKJNgdhShRNKKhWoS
BQ1vKSutW9EW84JJSKQZmBLOScWvdiOWAs3fcnirpoSWrAjn+CCtrNpd8r8y6CCi
xMA+PbjJhg8rko7yL5vcmttxtBaJWhRYQHw/9lxD4OZnfkWxVDJMtlPCK49EUDJA
ppbreUIZF18JvSOQil784bIHkbBLIvbSoLPmSrw+vpna9+g+yAHZky9wuHwGjXnK
6zkln+ODGy2NtctCraRGU7izwcjrNfUpt9S+slS/GsG2JPCqm/xdmPi+M0i29mJV
JcXjjaKwWLIUD2s9msOEb+UuEuoZb5ihPmptcb0aO9LhN95u2OwlDucO5TGd6COY
dqE5IuFHzL7dZsl2ezFDmPc5BFQjFN++ZHJY21Ny6M9CBqd4EpVXIPBpskdeUf9d
pnsd6UY5jCD+pRLYY20xo2Y2WKk4FMl9BXw7SBPPANfnadq1ezQYUvmlUILZdcM8
TDnPKdF5EzxSt+elkoTBesa/YcyYYn0ne1l64uB5gHBBNzBc7QYXN7szGczM3x2R
UbJ3OgyH6mWNTUAFZptd9UME1x8Nq1rotAe0CzLVdBOhE7CgGsbKyNh6rOEzo81J
K2hXGEjBbw+sjukNx83qhwL+RyVnzYne9G6YPcald4F/6mQXSb8LeTpUlakAQ/1R
1Me2u16Qgo3wbiR5fcJYJ0xBWmDW6BFktdq6i8wupSUJkKGeH6QAqrH9f3d5Lw3g
0gwcXtOW8PKm7mawQDpsDEqMfWPpH08K/EibzBHVk2fXK6XCN6LOCkuiDbdv49aY
MkoK7nG8Kuw5xN/M7o+ljMI6FyhK0lhGYp0LkVS+X2yoptlSOEBOKUX2QfigQh9W
8ZyF1ZknGqU9A6fS4GzpuV7mtZF4N7FjIxRMMLz+rb2rbU4VCIRxEfXDSCQiyIr8
45UCUzfB4voMYKAWS5yWhdsaQjbxPCZK8zhoZoYtJ4YaGKm9g3QWPkIgnotSt2vt
H3SBllp33YnxRLrILRgnkycpLUiBi0FjzL+4HzQBWwyxXHy16LzgJB/OSFESIJXd
75PUaZ1+Q0ADca1T0gpm2JkP1D/u4Gj9tTlYXJLuGhVOXk+qZlQS0T40IfTOgQA/
ax85RrXopeLVwn9b81y+ouck0Oj96Gf/nOne7BXYgKyB/S8itEDTDN8Xdf6MLI16
SiJZiax9yp7C1bFCohzoYbQIEZvuhtTX304yYLdzIrBmgVN0ihT2k2jEZQIQNxqN
CoK19EfqLAVspsffzduUjyhdyn/NkspH5lqgzQKKy8DJLdR1Wc36OGWeA19fUlh4
rxNCmvqC+TrfXjtuogV9yHY/ggv+fEjzbOFULtSiMvdwU6nnm9L8MkEu4V9Nicdk
D6945OZLF/psKsV9ChWb8Y2DqbgRi8XENn3yPqYCRSAvFiW1PsN58MOgEd0TkB+c
k39SGvnEOG77/PvqZ+xnbUpQEDox/9jJUWLw4Vip6MHdTdkM1NzDD6EPZbq6zqU7
5wNuwB2b/w50KeWbjQt1qAFGdbNiBwR78+ULS/zcp2GeTokVzoq9Ep8HcQEK3F0Z
/6iN/xSlKX52bs1i4u7yfU0s866h1vCKgnBD8MDg7HK3/4XFKIbR24qFX0wtzj6L
QGPPA6XstdG8XHvzhtsYNSq/ZqrYoKfD0KnZ/MGNutgr7dU7/l0a4JagjhKAeUS3
mXYFHmV3Dwx2Aw7bloL7P93d9amiLu+8QfjbeOEyN5O6xxUX7ItF9M3WWn0FjzIz
23rLZl0N3eKPDVXbAn5Etwmp/GpJuxGL8r2Ykm36gP5rQtAQO4MT9+r77vRRmZOl
nGg8o/p8sbkeOpZZ5nw4paAJmcMYH+J32l/uNPd/SYyWZZlwhGYWRFOj2g9Zlo5l
zBBNsqlw4EvNBLeFIYONIreU6iwzqg4ZyCDZ5LblhXyDNrihQ0hkBeoFZCoImEPP
Ryg+QUg/40BU982kx9f7RVSFq67UUdAic3xj6FiOUg6I3Uzqcm0W881j0i+1tnuc
bZpXgxEgbIWiuDih1rw1KQcIyslGj1SrVVcQjel4OYeqlF78mVuLo8CIWGcCQpkA
UA1SIYGlYNBlcbloYo5YX7dSKvbG5VajAeCISjRjOG+oy1kp7wNnO5d688uCXT3i
znQIHqP4wCPX3EMARzlHz/UZgjx6BRJAnTblqooiuU06xuJf7I1bGpjiDMgHBmAh
7v51PjjsN/guShPQQeccMM6DD3h0PBZxGNKJAGS4OOborH5f4jq206xUqYgfVLqz
sSo0B5u4iOVq6Z9vh08+83O9Nl1kUeEC6fSBFluRxaQWB+5dA0VyJxrRKC/zk4dC
RReCOwgMk365lInV81ByEX/Nqm9fU1vPFLZA4PvaqkLOnvF43yqwaav26S6gjDFs
36F0wlz8Zc0Oo+X7ig1+xt2x1miTOR+dSIvU4SIPpbQ3GWwLsaJAQ/tYkM5vD3/V
A9Is1ko2e+gyuL3IcX1xP6jBQLYpi4Ep/znj2smmILMuisjr9eBUeNi7xdojqD4k
xP1UW5xD5vxlsR9nazphISaI1+F22Q8xfMrdXMcKpPh8GOysmi201fSIw+CR2w6L
a/WXTliG0kw2p+gIo6Y1ssHbLPGMDuaK2s6U3EjncLuGCXwpDf+GyBfJUWN5+I+A
PO9InKgUH4TLs5R+xXdZR8f1Hwr/WbhZW1p/Vk0GVSpyfba/lBUiS4L7jKk7V6O3
gCCYZevsG1YDLKf0tU+/vkOF7vtKMUMaHM5C/9gQf75CMtEZXZ5i/c6+00vK7C6M
0DJtfUT05FAg5FMCHzPnncQ0OOj9O0QuNXIfUFG6oZG8wPmIhQtBG/ORVBbGJGhk
+21sBD6+RJxKUSeQ3iGtZ59HTCjaRN3UF2YCX2L9WZuUnTm6cvYwoIkgODCQ3hyS
cp+WjgdTa4s7WjU+Soty5wdhUFrQ8V98QOy9tzjf7Gjl7gfhNZ3G9k4dVfqfvcng
JBEgGV6P4UvFfiVG0ApFR+2DMcT5GGTOVKx5HA5s18fkqVOB8kVUwFOp+N+1R7yL
NGAA5M3nZgz8aM7pE8PyO6aceqMs5HduxDWPZ/6NCcpTE/0E1LqzGJBkWVFHCDsy
a4FPfOlSwQLCMKiXCxOqRnUBrrVaeC1tCmRLiSAVG8m4q0qTcOyE/zD2L1UChcqj
A0CdTJtvoDqeni95CbkKuyhixN6jmjHyxTTuNuQEITqgzKlF2AlIKE9TGEkDoQHi
wGDQdIVtleWXvh7r+TnG4UhoT7ev6f3ATb6f46TElkksXEWM9DG3rMQQ5tQHFflg
cyHPO/u5mVtNr5Gw4DWUBx+LGB/0z9ReUUWjrLKV6zDrSTz44lJ3FMsGbuGrhlvE
FbAWbN1L8i1I2ZP+e+YviX8FLr3SynnUR0kB7k3UQpKlO/XkfKfd3x7hJkDKPmwL
Vo1JFXGey9xQ/7rAESTFcuLcdC/n6YlVdslm6PZpt5k2POQRxiUIuo/TndfEmXk2
UQAMPChMCe6oUDLjixZBNtkW+z+T+hLzRMYjVltkmAkF86vUsHJuj84T4tfVRf1h
c2klnnipcAK/DmHLHGImoc3SK1wU/0Lfca5w4+AiCxDSCdmfeC8ITwKlOD5o2OtT
MmW22B8wDCqNWCuQRSih1y5ry+jacszkXxhguStASF3P33bqALcATk5cOXrRBtR9
FouOkT+WoNQnUTj/OeROUqkAbdEtWwOCQOcCsycdgK4XWpGoqpo8hPIuzG2kfodf
f/k4mZgOO7mtNlsZ+JDuj3xgJhmhJY1sbbOdgBWzV0QccAS4hVvh3JYVFIeAPxpo
6f/Y980lwTf71F7dSFAuda7y/BHsBmrywfBRTfK+Ay0QfLHvFvM1ilM2ztuHzWKv
+T0SoC6KdZUzY4VBuEQByrEkGxpPenNXJACEOjoBIaGxZxqAv8wt0vdKRW+YOPCz
KjenAOzpr8is+jXdM/mhdsi6W1LGfbZpCGXHQMrADHCzGLQSJ573OmZH9jG+ra4U
aWFfrYBJDISpfoZoMdnLD4FD04diF9BhIKz4ybxsVUeOtg0lLtpmzUuIzt5KGO3W
//7oKSMPdOah+gRTFlYOk1ON2CvuWpY6DHZ8ItrldaZX0v2mDzlvRwpOMClbwZBy
gHtgtIr0iwrcU6cjhzQyT3yVJZhGCoGt45pHrpaRn42MsslrGaH7Np3MdtQIN8mb
H9MAEZh3LniOC05GAgV7L6VYcdLkdIzw52AwAZmvo4ymc8VeDxtSsm32KWV8BALa
qIMff9VfpjPJgblDr8f8eVhlepeWJkCTvWXF4sPy5/5MFK8+XyIuNbg72pBm71eO
e7cS5LyHwZzXIOqoSn5CWtmo1oLAb+Tq2q0At/ABoiqgMQrBOiTt+3rGuGCmy4mV
zVpNGflOA3meDjQeEyleEPQ7eLP5/Qhp9qi/1J3iazH4xJKix3QEx1Irx4ffJZs4
rh7Ryku8ceAo7kbsqcHJfOcPJQ4tGjetE+ZHeXsXwZUE+gCPBX7iQeY3wCyDG0qO
QWAQ1cTo/SagmwBA761tXHkpjxkeC1KxoFSgYNk598TZ72MWC9a+LtCq1sh41Vc0
RVajLmg81ydLeKtC2Jd/CUKY1Kvj1dxT9L0LEA5TPW0SXEk2GQQugcflFPmyIFRQ
BbwckBXmEQclyU1qH5dKRyszDqVGP2dSF+m33WPUACI9G881mq3aLN+uJ3oyDmSa
/2Ykp4HAsxg1Z6i7au+MeJDEP8RoSXC9a2uUkOdT2uQknUeQAOcJ55j/r6edFcQ9
W5rOR7eqyGc1xAUJFwImEfPuT7UHKt9kUMIAN0+az4c+leGXkbHLBjO8nMxMHpGY
u455Wuo5LgL5ME20tThYr97qxpPC94zDpfZVoyBruvY16++in/vimRkfa6DNt1xe
vXHnHvsKvQVjdLOLUCHCdli2bsX07ah8sOYzJs/fgTmQRhYmpkl5YVzteuNkjyr/
rNUd10xRN/ZBBQmeKhzdiDJ6Yf48PNvq5Fp8LEq9wFSUKB5YKVaL7gXmqKXya+E3
DK1fWzvsMZ1szz+K0cmWSkr78Tzvls5FzL41rB9Nn/TfbFwDPAwCAIvj/rfAiFqX
U4Ve+dKn+xj0d54uyyFG4geOvUBltnCGkDe64yEI67vzTBB44wDwbtsbGJtHLxY/
ExHS/sJJF/Bny26m/dyV78NlPGUFvELW1aO+C75Ud/+2yFlw48B/uq0uuryKM5Cn
lbi3njkg/5KajKiFcgvgQp2wjANsXdDUPUtdNyQtyTHt0WsQ8IqMlIDq5YPzx++G
+eZhS4+MzMt1u2a6mqS240CWiwbif4XaSObseo6QALjwgtgtJKGdeycU7rOWBC6w
oOKrDWiFYw2XAdcgi6ZgatG5OVADM9cr/61e/tSVuTgK+KyGyG0agUwJxJG8hZVr
kHR3WCLqqy0peO7p9CmexT0lUHaoUXfg5L5TXXy4RztrKzP9fkDLEzl8rtTinQNa
WAxyuc2POO+FHM74VyDURvlG92Wwc05XlrBEhz1tqS1DU1DYUAItJNyh2prD4n+6
dn45GZeTlrcvpZYkZJCjBiw2evOctstdZY9zikk2MYRrWyJl8qUbonNP5eCTha70
fRw/t9kO/LKMyL4nMU2pc9qqQRVzBvmW+SYcpwmlJy1wJr2wQG/2HK8MZ3TRtBTA
hEV5E9kGBXOoLGMZKTGH2S5ZivqEyc6y9sEqgiIdur9eIoVg1WSLi7ax9Z4c2WKb
gxgi/ffrYwXGn9OM/eNsOLDjqeTo5AEnVbi1sAle6ILXjLHOpBVZLj4mRp/LYJ08
h2XCY4OPMFfHIepjFWXPV9ZQfVtUyA02AKRoSFe68344GQ/sAzRH0ArkZvL7gstK
hkF0stK5d4a574j8BsBeE5cPYjztAFnpVN36iWr3Oyq4dES3FzM2eLZn6PBpbGTK
5urMOujD9l64175ndA5o/A4xVZb94x7U4n+cYK/spzlJ2UUspMuVqEELrEvCApeQ
EAwXqZZv/FAzlJ4vsVQmuv53Gvn98BUDLEMnwQo4FFANuuPvgKq0wQmT84RBwlb5
35m59i5OrorWAMKv797TNQQI0aw2r7Yn/3o7eR0z2NIpIAjTlkIUE3ziMgSnnubh
kq/URG7zO0mPwOhHD7UNvNqaxXcV3rIsUOxIIrMen9Ul1LGDFBnwvNJDX7QVzPEm
Xj/wJ4uXKJ0Xk5RSks8VqT+1L8nWBicU21BUVdkGCcaFsDN9xIVvrESHvpqcDXB7
1rGoLUWAgGY2vqe/AgMD4u5o+k03SstJ+yHDBkrzCcGhpWHueaZk+Gos2e1ywSV7
k7fJnzD5/Vs5ofVw3v78pO6u/ENgANa7OhdFQapsWN/pvpt6yCMba4EBU5tBjHuC
Pe8ikx0v1gJ5pYomOrwraatpB8Kq4LuKI9Fdkl9mWfvBhInhZyDnkGM9lkHU09F5
JzIkOlncUaZpTnKmyohLtNF0T9QuR8LY5nvetF4FzpuQxlk9wx1IBtI0jKYmO8Xa
Wod0/1nAJQTGYFxhYpFptrgvCLXyaUzAOZDus18WuehHcbHs/sIG2JTJ1t27oBjq
kXi0KQy751USSwzsZ5GmaOcKQsOyH5R66X0+kgbK9/PNuObl7dDBeI8cOx830vMu
mOx5222WVY86BhBKKjCHz3VfVReUi5mjCO9lUqIoVK7jFlMRW9kq3ta67Qf6pElc
2hcVBfugFseNqapmVZSbdjxGuFm7GaVk6ZxMnvJBEjNU39cy62IfSlQ/C2tRWHw9
tB4nqqhVRtk4lCFzDjZI93SLyQoYK5IHmFsnjt96Pqfeog4gaGHjToMlIuKpcEbf
oVVyJN8mG5vXibdZZmWP6+YBhbKyxKKOkqmc4KFkV837A9fMKHPB62a6Vo1ELXQr
JBfI/phogH7Hve0n3AUvP/DY7pzUXDg1Jla7QSx1WKJVgxf9ccbBJ/scKnczaBeC
lOFl4wh7L1iiOoZVtnIOHzrEgiWe+YNmX1zi2WjO6dgQ1rWiRok8WTCPy3aiYWh4
noaBmjaJe3QK2rPC6GTwXRxnYtTR+jyt74GXt4V/77I0IBv9225Ulq6Qyt0Bu1ax
JjorPNqZdYeIq3nef9yVK3h4aPYQDeoxZGd/oWGRYchg/TDIED5pMJ/V8WIeqcjD
MOusN0BIOxs85kk6kBVE0WmXaA11FkHeOMzu0BpSSjFV4ASNwbeagQhkxiH3T561
IlhJLV+uwuaWpB7U0VP4Xy02tM5tYX59hZIEOLkbab5Y5MeK2wa5I6+kmA/RCmee
Rkx1gpsEjatUnz6EAgWtsfnEaeEMCRrinn8GJYVL5G/LQ97dEpm4YEcay61JcKvr
d5tySqGYke7GyAHyz2J9Fe8UiGWVqBIJlyfYSjecoQv9aOOGUg4kow8VD1/DTM6E
bVomOo8sVABPWXPIqRqsrgZejxVJBpUQSd/0/dIIuFSiKvvUv5AaNBVFSg0jLOXL
52Dk0lDcd5g3WBsLphKnfP/TTu7LHFzin17M/DlvLaEKJdZhnjDKiQqvAodLfaa3
xnYDNfwfEuQYBPpVU86ykU+Y5gKXF8WihChjoTL1+DU7eODVaigWruSGzw52MGGP
wMb7ngJWTkptzfcKeSBdPKXwCWuzuBmDcSDNW6m4WiYSKZHHBewXN+KH/V6TKHOC
mS9IkrmGkiqqyX6mpjihCnxhmL3xIfCZw87SJZgSOTj58r/674lRO7iyD8FNV63f
HDG1iFp0HBWcAeWt+4uRZGUa6L/udoA5CcJlpZsR6q0ZqPizCclzpxlSLDx4GiWU
PG6NKVtJuAsY70QCjQMlPN5MRo4QGqmuJBzFWZd5ByfHiUDwaQVM0VFfkvMNhg2Z
JBEvziuem9AWwx4q/h9wbgd+6fYu6Z5Ru3K25xbk6EyamI0xhvbuYigNVNm+81gv
IgABousuJz4x3cTC4KuCXh/jzEo/cWjkLIsoDMokmWTE0WKvmRuzKpx1Jld+trF9
vHdhzaB4+t88AQIvlizQso7Oa+Tn+f10fF2iVaD/L/tu3gcMtjhU7hHOUdQ9m5PN
Pzty4d6MJud9OjqjkkRtGd+HQrbVlkfq/VvHb4Q4mW5MNCx4aCwrTaWpHQw5R9DW
L7fuHq93XXWeZXFDAmO8QQCdrJEZf9oM/gHmyViKyPCQ9vLHINoOEoeV8ODF+RaO
Mbg8HlCbD+H/NC5i9kF48Yx/2DBD4Gkg3H/cPe8DJn+N/D+0ibakZ/u8y7JlV0DZ
CsxNdgb3FzcOv1WhfplFzC6mtvW31GPasdYt2Zv3Pqz5eyVRF8mKSeBJoZLObFq3
9Hlu1ju5+2cQPO/d8reKc+8qNrJLCuS9B3UqLi4OTJolOzuPUTuoLBC3SA/ZvPjj
FQLPiqReDzQ1CNo+3Yp4YkflJXsM50imoJ+HA9QcNqJOPWAOwFXMh9T5yoHhX6XD
d/uxpLlmyuWo0TtmtTJCN8zfwUlBK2RclTKLVHYTHCypBZ6FYE2r5muwO8stVQta
RdGV9Co2mu86Q/Z7g3Sx/80X4dk+YJi7x5p8DYZHKtUWHE1GfQz1v3v5LS46GmpV
l+OVLHrfhRJ9fi0rQ12s6DZrSbODJ2J4VyWi8/RQOK6g5yDDEfTwdqnXcYwEWG//
jhc/CH+64iuC5f8QhvvGNSVglyk2ImKHrP6XvYzj3bV5kZh8Dmr2PiX/TbE9X0tS
NLL8sIvaSULp0gdnteokidLquMNcmDXEfvT2FRASSCi+rPZG/9t1k9Iy8inunJ8u
CyOdqW2ZbvdFKX5fiQw5w8UHClH+4xRpt+V0f6qB03YDrMM0Ws7/1wKxhBB4lvOU
u9LDAaq6pi5/zDGwgw59f/jnKRkF/rS2SSjIQx5Y3P2CrVhFvA6/+nNvWUORAvWG
dWUDrvQozUdknsQeUoRcobqQPRWHdOu9iTlzAJKFI/XSUzl3EWqnGWL0IsW2jZd6
QEgtsb4Crfn/vLXsgU6uJX1/Fol3WK/H0OhVoo4XDoKFYdycyggJAuTIXN3M35AJ
DhgFmEQNDrinnE3z9F2KL4WqrvCusx51c5J/TbcLiiuyTYzKYSZZZ+Icj6ScVPK2
7s6cjxcj+cMSpMn8lkoJ9rCuBdPRLDYCTkqPDbCiBABnPqCHgZDBDtE8FUXecPYp
L1v0st1ZQ+dUhQJpbPl+kS3mDguEJW0uEHtmr4ECu38zLw8ENsBNQ1MqNk2GCV6y
N0NOwE2jZG2fKtcrViDJGhtmTeqUz9o+KO8MdgKxPWvzB4oJ+blNBuLrolJolKSW
bclg9ra/4bajnpbHbLoKz3sA2F9+hQHIkoxiBhW9YWwp9xNVsJgHwlfOtLssPxg4
qtxMunjQ2HDegyuEBKRtgET7qArwwMe9zEQ06/Anid6e9qE3mFGGrQ0G+A+Uu/c6
pfrGOLLYqgrNS4Nby5uIBSZborbgb4uJOlAAGJaX8sfZdmwnTylYgwMXqFhsMTl9
cocFnlo+o6l0IeY3LWMJfWUgR/tR2XYAEWLmwpLKJjofXbRBtupR9vefz+N7uK79
3pXvMEbsdv9ZcFGAmSc5wYH6zjqEiLStp4RmHaMLiAMqf+hVR2cOEWKm71G09Yni
29dRu9kgWGuHCJivN5/UMOvsMHekpdm3bskz9Ud8QSrD042IDop/9vO9WmYO2g7a
MEYmBFIzCsYe761kjH0bd7BcnqINGOpPW+ZebK1DDovxe/qFB1XgR+U/GTOj/wFn
vHC0dUfLWjPV12ufBjpoJukV3KGrr25p2C8rE0hgsabuUCN8KPrCQCfiNx44M+K8
CEaVFPsuNGBwYTfLO5yk+p//IBfGhdX0dQxssT8KvQj0Lp/LGhhPhzUPYUFIHsMO
++EtMfmq4k4LjTPkwR4VTUvQ3efJne4ERMyRtIyoc4goWyiTdyoW5UV9Cg8Mi87H
LbY04PJu7Wnpa+ho+nl2CeYtzOK2uXxrMhXnfbdiHzzlqkdqkOwz8EZJdULpc9d3
yGh2jyAuuq4K1K1LTukUrMF4Yrup8asGOWPX3Bw3sZV1LoJHgw3Wq55SMXSPXwtR
iBQYAqz46vwOn8hqFFsTm86Qi8bF/OgGrpSCyxirvWxoB6baB1s7rHH+PF8Go+sj
mSXE4yIbJFSGPPLqnKE3fFfSDAClVWqOMN5UPOPoZxSI/80pP+C+AjssEeqIn9p5
wvmXawFmHLdbyeGfT2qgWPxwKKewNB/Ut7DB7Dqa+OkrWuUuIdNt7eaUDp5lpxwh
QJAiVEcDOehnZF/5elmo1jcO7aZMHT1UCJqrl0qpYGlWoC2bcG+txCQF8x+Wc8Ri
abA/zC5dLW3SaikzejFgVV5oWteytWjGGZzhwZyFoH75cbRT3AIH17YnRiaqVORG
HLotipsKx4u4RYu8OdlXz8xlRxDDLNBYfe6lYGP7thPkwWeRPoJxnISf3BKbY6Gb
1p4JOrfTGNRuzpnKuYO7GLnsKEfK9ltK1P7adNUmffLuByxFjhcfNj8zhFNHjhBY
IKXqq1PvlMRhmOcj1EQFMuqk6su3h3BeCva2TRsnfHag1yb5xb8HtZY/g25ef/Lv
teB73Bb68XCeIYp5YkDufDKA/WySadi5FF41VbmENGyXZ/WL65CkHgpKyQ4IpbEU
6w+b7sZck6jwLv6gDG3Jds1pLy4M221169YsUJUeAAPIiFrAUtHKIca0u0QVTQZS
HS+Bb0V5DTeVZFmigPvbYtsBRsewHt/GdpP1dFvN1sw86ma/IGnINXuLpA7QXnw1
3GFDB5HHy+I3+NBaM+5XVx1WfjOhlRKR8DLsqUrvZgYnBoz6s5STRD/dXC4s9I0i
oZWf7X5o1wuOPFYEp7RPBxCE37kjzlheMWQGJtqNcAHJSdbfWyzIOUcqHG7505O7
E0nptIDCxBa2KEhpoQsE6Q3X0meUYErlEPOi5tRGnWMrwITkVGMwQz5PxxhSnZ9R
13ZWbhobl94XV/8pjqMoc5EiJZzuFu6o18oO0uL59/brV5Fq104dZy98FzzZWfN1
5q494iDhggsew13iSbPR5xv+DP/K3XsfI7JTWhgQhkE+GxaagDbyEOJayy0xiWUt
iIek4QDqJHMRYyjbev9K04EfxHt6V6wyJsWhseRlUp/xpv0t4alhBVBK87HSs54X
5M6CsO6BICfKm0xADTisfx28t7fIZUKF5OATxfm37c+ZKJ1szFHQenACgbbdc25D
ewMn17godNSiG3b061frW37X+ddeBl6gXY0m2SF6fmdN3PPUJK5Mb2xN+yYVJ2ol
0ljZmPn4tsHCzEjjr7fKgQ9udt2xWcXpUFmAFmrOFW+O/TCw8oNdSU45rMjxdKsY
zGqByFWhG4ULyJwsMijisB+p7A7TTvp0l+db5r+saoqoPIIwXUpuPts1gBUInCMc
ySsAjEzS63Pd0z2iB5MtS1yBKcg6mYb6zyjrjmpL3G0v7SStlXS3G9EDLciuH8sL
eIBiEec9uONSFV9+TFcwzWCbgnuXRrss8j1xQC+K6BTeY3bfwznvvYG2Zy0pSmET
eXzoFQ39l+x/trJwyfmrEt2l1QBXD9nwmhWojayQNxSPv6lAdNeu+oYlrU+YYyYW
jXT5XA5WyfXHsJTYXY7q3sRN/J0AK4V5n3PVT+p28vvMWPNsYOSHWRJtXaFJ0Hie
iuEgNpVh+cf4cmNNT6tg9S7OJhZ7+d9XBTfd4R9EOKgMbWEIZ9WEpu7lSz8ZI+NJ
muOHMTL+uF6EDbpJ7yHBpuk9wKCbAwIzZs2daPO+sISwAfiwpnuEtg9E/7ZmgUDi
ZhiRetHiIz1isfWZYZGnbtxmWl3Loi6UcXf3LBbrsadeMuFG+UY+kg362/7W5UFQ
ZOY9Imd3scn02nKDB5lDAoobwuVTZrDJ55vSQYw26SqdvwIJrrY/YmXxjO+OmdKM
7tlRlIWoydu6lyHyG1MPDUdxzGHlRMVhr5jjD2QxMEbzaQmmjxsV7BQaTJlVLNq/
k3Gs6nY0ZSZgsV7IpuhF69Bbpi347YDNk0NzTlOUj974nv9T6pzZMl6zzdgPYYPw
C1GlAcgt6nas0JHaYh8ZyxKrJ7lIu0jNq/XVMLz4lYuIhMf0hmQdV9wS8q6xswJ+
3UXIxyiWi/D+ULMplwtMAjEL9KlOHedySeboUSavITbAF+xADGAQ9CCiTRvcYHZJ
aV7q6pFsldGWIeyyLl5T0+kR3yUBanzUdeadgOCYUuMQBLOsz0wMmbsfxlu2B89o
ZCpF8jkpm73eAVnTu1x/qO2XBt89M24aQYURP6/1rG+nfiHu8EJ75WZzVHvd9dgy
QhcH5REbKl54dI39n7ckhxHh5uRu96P5WCG9Kr/8ay8glzFQABjreUdRhxN8k/c3
s7JwTxPi0Ad3mfucPuszb4txUFr7QzGjGgNsosv4wbSk6G+aUAWeQ2hiKRD/LoZS
/IpxFzNTJU9OmiPRhaF9hai6ZxqBJ+J9BTI2xBcqRFgQGjQPVdQZj70Xg85Dzmv4
7kt5s5h+6tcDlMyR8CzJy2sLrxAEAnJIpz1qdVYmY/uJNApmKmaaSjIUnXsAztFV
q5E9hClsLKopGE0hqTt4bSC0NSU5YxxIhd5vGXyuUnRmhKGY9ltn95gHXsd73B9a
se8a9tCSAv9+Q0/hBkJYVTePY91M011R5mbAoStjOk7iDuFxGWhpMKjmGMDOb7LX
uqXOCpSWTpGeY1a1Zn/fe6OR1qnBhtzHLuk11oMvvZwMlMm20xws0yf+vhHyOZ65
zXwwGZ6qwxl+EJdr+O5xJzq4Adf0Oij3eGok42We2CFEHwGskUBSW/8wzBaU+B1O
OZT3pyr3z6+mXx7k5T7Zs3+6fam0VLW4gbmt8CbGMc235wvCgqVzBWLft7Ztrp5M
6dW1UY5NI+Zf09en5EDg9YdRdyCHx7kLkqEqGuTWIdpY6xNgha4XyHomMUCG3cWv
mOEf4RPXBYthPnaWRpREm+p27p4ClKNno/ylFNwzxNxiiHP3NL4GEPWM3qw39Vlv
idR6EiskvT5OjYxWyaXxoCEcNhuKJZ8GQ6qcrMVjCVvjv1P4mtGvM1rmAMUmhUCE
ZLo6zH+FHP4CNQqa2xmzQMNdqXhr4Q0+6ayu/M1zIPNBR4WLBY8ki5Hr5Q2cE1ua
aLRVpMhuRLXHu9AfP5vrw7//rEueNqVqq2FMiFL03OJ1y50zDgHcFUXdoSpxx7eq
jXogs1roUoW/JtfAqHeI4mE7/KWf3kZHXe7ZUeNqUr5tJL3dGO7S6ZOfyOSbxfaT
XTMd7u9jQWUhycYBd7kv8R2pk46hGQ4us7gCV3yCeinhVAoSUMILZT9onfI6Ovo6
Lh5KeslxqOrg0XuyLlUVupbIkdmhyQ4/PbnQulYn7xCk0qRAEPitKf7QYR7VFHAo
PhgjDV3yikNYt3G9EJup6Pl/GjTOH/3KmRrIiscy0aq8dC6Bh2N4BVjz4eSMVsUj
3qOUFUVwzCVHHJYr/NIxAytVE/57ucrAntKldUB/xZri1po1YCIkfuuaAXzqdDH0
v6K1exgM1lo5Y4BPULF3unfr0PGXglpncCJcyE2JZrJqZ1fgTqrhujIy4p6mtZgH
CtAmrb8l4DmuXshdftDxFebUSQK+nSOSJlGqjYYpSumYs4JoefM6STfV+gvAf8y8
HPY+AZy44FyAN0/bbF0hB1QWXWUkIoPXg8C+MRuXQ8hFeWB7WdJweKG/RFlh+2+Z
juJwlFA1B/vYHZWg7/0kBrNHAGaLpEKYNZS1LK9BWu38KToiyMZnf6KZDlSxnkyR
N3Tf5E0Ipy+QFavHI+PiiYCc+H5HNwH+uEoqYW7xii/f/btP6As32MzhWzM/sSlY
zjFbR4BMCBEmXpmXMPxWNSbFaebu9WdT4Bw3o8Rc5nFM3EPtC8Z28v7Y9o2Vb3rC
Gexne5dwlj6uxfHM+rqF74UpSPHqLNTpxG3k4KLrDCMqL2W3gvtOs9s/ofn8fWAV
lyUunWvgNUsB5zluY00nEXLdXrxLIW9mYXE0iyfLEcOg3VuWZGQjvg89//m1CLao
SCxyGnZghw6HvA6KeV8A50y5qCHFFBZpEIwbdGFdnyE8nMpIBiGnOEnqjwU8Ypy/
ugyJ4qZG/iwzvZ5bqZt7J8EBuP7AZKNG21YxVH6f+eMehxXKs92hukUfIRXxLzq1
b1Olt3/s5toJYUX3K19p+O/tjHDseDM+yxAkbk7PqH5R/+joH3KwTvX5cKZyyD/y
klLi2dftDfbZ7HvWz2ZLGu5pCnkr/VkRdwmT3b019ZaZquTnwsTulyqGvo2wAt6b
E2Y1Ai4jXRgsXMVkNKUFyR6f1EVna67guyXPMJ/TDQIoa+oA2+3EJgndlSSSDeid
bW/5cz1DJ4AadWTuCt03NV2NTmgOV3c/FijXOylXnl+uL1Y4rYFJzf6EvFL1Za+e
AQ4mrZg3u4V0g3GBG0/JQ2Zd/vKt1U7TMFrQfbOJF9m8BJSPKqzQA83MiKeVJN4l
27EhOA2sFedG/QF8NUeVOxNHh3DbH5ULQ54OH8DpDsHs7XnrOIx1qtliDCw98+VF
8v9faOiOjS9uXGRdcAHI3YOyDRHaQUo9e61IcJV7oLLPGoC9JwslWTaCJgIY/Fcn
a25eyTb5egd2xlLNIdB56AQJhGR6jXjTpiVcHLUUDqcKRpsDiZErCaPgGL9Z5hU9
H3y8Oqy6ZaLYeheqxiqAYyFsbCkj/ZplO7bu0msSXJfjQfuIK3HVxCuw+mk/E6mx
zII0MVBpfqFor7dM/5qe1CH//rHYU0ZUuaGypxa0WxEkB/fdihocMD19mw2uUbYo
MeIqQ6UwuhbUhLLTCkFrQcipYx+wChEqjfkVVvdMFkYoI0hAJEl/oI1niaXYHoKE
a/UwqMu4O5ujYgX627WoUa3k22a69dm1tNZ2l4QZsyyX7qiPQhZhYJMnbo2+DQoe
TQDCpg1Nwd5XWSV6WkTLZ57q/QU2EH4xnaxxqWHoh3dIwkf4FonE5FjGoHSPm/G/
97te8Ssswj02SqZCDh8WWtnRTkSpKy6BB31zyAesRw/KAG7bZnZmR9A2XCQTxFN4
jW65oa8uy1RVWGnJF7VlGeqXDh3kcb5//tYPXw6Uuze/lrX/DK744D7HtyhJUrqq
Eg+cYUdl1qEfnNx2hrSXzjp/baSA9PvUIM0q5z3B9w6QJ/iYNLvOTcmNbVeBDCgI
K3CpX1CjDefPwglKTaq414XiNTEfz+qxUB2KD2bR/ole4eQQRIs444z+t0yLvMAL
Iu9/BJUUDdpCYDdTFCVBpFCOTgU4VlwT7hE4+N2gjhRpS8mT7rzXHW2rbCi9oBeR
GQbL3UYIOfr9DaxDTpmqA8RSkulKS37B4Pz8YIDVC4UzQEGXZ24ZR60enGWvqcGw
QRzUSqMPyEEqe9JwWgJS4ZSDbFT/o+JvFUmArEYZW6MK0WtQaZouUc5KrDzAz/1v
PRyJlpr++k8WoqKAbX2kynhmNd2McuREIFF6G4TDs2W6Ij0FVZcp1Zzbpc4pQ5C0
DqtBkUNh2xqp3Ed5p/WGmuBOzj9hmPPvZpane8eMsjff6GmGJEYBevooruOxUuWe
Er9d2lxlOYm0IMefj53fody0S6gsXog2X5qADHoCDI4/OtFN5FsFOcR9+AfXXG9i
HySzfFVdgUjBWO81NLKSD0+Abb6vERcHOvqCfRZR6lg7xCGjqlaJwzkhAVLd1zT6
1WAKZbwewHEzWwBJ2nHSdVHa1a5mC5uEZRpzIoxO0h32PDAtNJMrRrU5a3G9Z18E
Xk7n0lDO2LXcVL/eeOVwcRKO+vuvyeUPmc3UPtJbCwqXurbuRu6GF56ONifaG97q
kkqurRpJJnuA32FJ9qO+PhzF12FFGAtpcJOA6j8l8zqSszo5OuYGiDR0RW7Ij3hu
bVEzoZ1JeShd/IKJOZU9rl9iJB+qRdvx6wUV80o9sM+vQrJJuxA41zZ9dVeWNaOk
DTebC1ypOWMXqNPhLZxVtuIMxu8PJ7jDsxgxVsOxUto4OgvIAAcWl1N3kaYkQGH+
iYsND19FmB/cttZh1LFihwx/TRGGvYaktIan6vZ+1qZQL0AKvcR+AJaMKUBpSMEb
wWi6cyiUxNLQe4eDJ5+gqV5cK+XTTvE8KdPaJGkSypuShQh5Wl+Zn8odynxANmbx
IGJzMwirH7z1afTuBiSmY1tmLJeVNiHLn1c3aBr/OFqJMq0OYkBK8DceNFuo3AmP
C32+2RK6c2zi1yjIriTNGbgaExu2UrIrFwwIMRJZbOqezoopbSSL1nKI/C6L9KdS
lGcVZLWGl/aX4uBU0FL/PALZvIHcLkB647BJyffWrZS6zaBsw4zQUfkVUsuHQn6T
88tb0mPzGZyFP6kDIi5Y5eyGkQEQughmdd5QgQgIiLwcs6kDgeuPVg3nEb9/+eGO
Sf+/XcmFMrjTv1Rr9nxBIvnGgkc3mgB6DemENzff77gYrwdtf89ljFQ42w9TOVNB
qO2CCJyzerb3kulhVV9RffsGW2+fu0pCoTNL/i5UWPlj/yvbB8VH9b3NOuryXrEV
lG/QZQKmm5xAaTKGwy+LhmuNGpO2QiOlBrb+Tyk8Bz7fLoyTLnBWfwBosLasUPHY
c1SKOB23uPxQGEJiTUzRdaQRDRm+86TzWtboZ749jQpN8CXGjjRd58CHDxAEjWP6
mbpgPDxGUf5BPs2YLPwVKMUYwYpF7UgbeyMNSXD71AklK/uCAULu+/Cyy1r2rWw5
xsdLI3A8kVA60y6PzRk2CZvPoM1Kbcfgm8ZnTJCFeEFp1hmFjopp1JhfEoBSge5r
AiOAhYqR882U1bMj6L35NyW+4wa0GE+IfUMoyJCnl+888ccFeK1cVL5gqI+mMhHh
kwN/r84ZEfhneq3GHAK0n6/Ajqo5bufKWp2nnJ1D2cFsBQa5mkWVKpaScz3b9/py
jKL7gJAj9ZnMrQ2GueFSSd+OHKt+HhaEecJmEG/8cdWts1rB6UCIPUeoDqw6NI9k
c6vMtUKpy8oVdKm1X/bVn5m/lt8mxfm0SuIsh585XSdeweE1ryhYK/l0SU0Xj3nW
K58E7T2Sr96eWbWSZ2G0TVOPo/VeIXvnZCZmKDCtLp1e2a71rIesgSSL3Af06rpv
zWX0prVOC9wA6o6aZ+WsNyAGiKaYFcZKS/MSZsvyw8q2SWBhKvB9uNwwnW229UzG
jWN4NmD1+/MXWF3656GOSPQDQwZFZfnPF548aDzyeNzC8F469YwkB5fUaHyIGKLt
0D1JatH6tzshVl3bdsXyzJ9is9w1w1Cpd/ZTdEnrmAk0FgNgIFapCXOs+Jy6xaPm
mLGd0Gfhz5RPSlQAAZ482KUJOtPPSy4+4dbJEc1mImNmiMTLo51Fj6r2XuqoYI5o
ppPAojVvQdAtzJUEIRrdFvytECaRXFYFmCRNv9NqjRJyLeVnqCF+0OgabKFEZntH
YO1JHp4M2r1leFjKl2B8chx6stml4Waqkj/uGdicOw4YK9MN0eiLd/q82Qx0aYgB
sBMGwM4+j7yaH3+3o8OLm2HeMuh8xI+TYlcoPQNViqPLzNfEhf0pp7vGE6olejTY
aVjtUmKFBnb0742QXaRG5sAz65AxTVj7hkBn8A3ZoCT+2JTuHNhltqn7A7Y0YrwI
FFkzzdvc3aFu3kF3s48ZN9v/c8Bz9kzsXN+zbXqUFUa6Zq0IAtaYBzwyJ19qUyXP
KSp2FeBUjJbMR1d5emmFbsypcEmaXfv5zsU3I72Sb3mNjp3NZ1+INfelw1uaX6yh
7fBmGrUNdadA5cKgUBLEZA47s2QWmtywfKU2Hh6Gbq82H87IMUSX02gZLmhOR0mM
7G/4KhzruR/ntSmaod3fVtlu2RSL+SZSwfBZTcDLjbZpsEDVvRqa7XjQXrGxaHPa
u8CD3hL0tUhglPIOG2MNtKihHtZ5Y+Hh/calkKipYh9b7ZmLEACUEPL/12kYFRHA
bsVsr9nFdaSyDRnOQvaXqVjcorZIwuAIwuigXxA2lY25p32tg3xjKzkns//hXy0l
31R2znmQ+3YOMGAkZumUe1bzgZ1O1VdhtVQHtVAhkiueGQsmTH9Vl+XG2oWKOmpV
SVjcw7LctF9WDoAwsKcW2fuipaoLXCsY+EtBIqstZLtQhEd+5nwqhFTC14/HBP+k
4dlhR0ltNqmU+hVMIM+SO/BUJ7UX0bFQaadesmP65L5u4C6HnLk3vI45XiO6/63X
6T2c0eaWYETD0oejtjNcsqZ3l6K6qK+MJNPOOfbHSuEP9kq4dnboWFkLd/ttYzCc
K07gihPDbw8ZmbMhtsoLHRpvkA+92+iAHFWNqlQO3tekhqyFA1B1XP61EBeumDZp
wkaoU6ezp7Je5fmdY7rfl1+ufosMVqRTwR1VtOg3zpXyJvsQXQLS8nAb6bH0fkNU
oN8n9fTJfzSDdh+gvVy0ks4Gj4AdMvz8GqwPtcsDDo/3mVW51sL3MveHTM5fG9BI
7sTWSb0e8vW7XuBu5vgf4HcwtR67wdPuik8En4iNPEYK25b4wFCFxw33lHtGHNeh
kwgAFMCjIc/1oOxv70kgAlrQ78xkkLqTy9ARCqBovKcIQz5Q18w+fKcw6AzJ4FnJ
iYrUL6EdpHI7VLutCVDQLWoVkbs5MWG+ThiJXjjPOwDK7KQK2XK2S5TUL+3nZcXl
ZA8S6nN9shMOYc3CDsIP0Jp5ppUTJYOzuIFfZ61NsFn8PXfrGtpI7zmdb/I+vTEv
WeJKowkQ5hGwzZ6CtEw2Y04fjdlSaTZjBbHHNYP5xSfWuJ6hX4ZEWc7xIoaq07mj
cSIiUrNNZc6iAwvIOY9LLI/kC2B4/2l4OGwjLSQOeU69mox3digJWdeU9SrnlJ8x
H6XUNUAu/fu/bcVdUc6MTVr1JgSSwtRnaqes+i8x0/IaZCFL4vliIPI3BZBzWGPk
mJ5oXpt0Q4RFwFXfmCMVMuArpAO5NewL31elabreywqb4JrTw51QFOUrGH5qSiUx
/fl9NEQTj6obc0haErWfUh5tlgaPq8QWMnqZgP0g7WcyH6Bjzf9D4YdfA4qbirCw
U/S3KQGB7uMCRJTr///tFD2IUVAbceBj/XSw9+bC94O+RbPM1DykaICDJsVXmlFn
N/nR0JarirE58peMRa4tGIzGaxYCjzocHZ7ajKr8J/OM6R0lDd0aeFHIIcqVrp8v
tNtxLkGuGC7CWhMiUkylwP+XOjFLA4T5NpKX6zctw9x5riV8F4gI2Lme3dEqYClz
SgIbu4GRA6cJotZYfOnnqJeM5XAb7NjtgIJp2AfgX1XPeo/W4+mvgG5UjPUL3gdh
FZbBsB7AO2wzN/eUMByFKTqTPKLhUOYKsbNXW2HYeCYkpufS1wyv1ePdVMelZ5S/
c7KRLZg9v52iuM2JVY4kLAKasJn9WA2ZzQ0qIQbM7HOxy9yrHzCzhWjGbZVzVTiX
Kkr4mpgR7m1C8sWYlmoVbhOt+0ZZzACUEVo8KvBl4yKmp5U287i7z0FGYUbwuyu9
WhAnCtP/r/7kO9LNkHa/krOqTpkX0LGILjGoaUbl4VQi61R+hlk6cpHd6hXyaAQ9
ouDqO/18EyFeaxNL6C5zjr627jAB6vXnfpdVRf2kIA2mXftb+qko8jfEOxXiGXca
QnsGxf8N2VOcK0YrDMeMxtH0Cza5kUSAn8QrTzUxNjIYtmykCiLZkjP8XiO3XYMt
hHDn20qAh2OeNeXUr96rdK+Iucbskbl2GCGgg+cbQ68ykB6tPN3Epp73ebb4hOJC
oBCq9O68/PLMwnJbmJZIZCfQ8VbEwUuu+m/L2fB8238ZdbM+eHthnwhWarjYTRND
L9ABFowZK9K4o9h0NWwyfJ6GbuxjO67BcWpWAyt5Ie/vxIVqC+4O9C5No+O0h19n
nYB4qtKIMtjfqOi9jz6Ae3tb8gocpRHRluoH+l3yhtiXoBL4v6dCjP8FYF6aFZrL
+ZRBK3HhdPtM/oIikpQxGKikpY6l/7T33gsXmrs10L8Yo7/8Mq2Z2A7z+lddNztq
TuBGbQprFXhKNyAez5fXYHCQEqyslN44exQULRs04bvW99PzjeKLJTy6wDK9cktW
rGKn9LCCgdK0zED6xNua8j43GuGiPBtOCbfGTEVeMM2+3PHAoToXs40Z5JQaKhJo
kcp7JLgUsdgG43BnK18QwhA2Wag24u2zS19+MxHXBudOuC0oDxouGH/ENWDcre9s
g0zJWWpA3PB8mUgmFyo1yIBokhRfTZXqksGU296T4kzGffJpz7LJohcHuzO2Xscg
R8yOu2LJdBvUPaXKwssKUTcbEzTXj6ZEzfIvBVWk9Mw5wUDfGzQ3FLwg5rb0Ga+M
LgVg7g7vtF+cTITSC9toe17EhwNEX97tpAFDwCESRedOllh0UePauVvYQPicsyAg
5M7Vaq3WdCaBO16DzkP56bCaW1aVftZ3lLL78UCApeeCZepYSm3dJ6pY/GxPljm/
kPDAxeMiXURPeWa2S53DcV30XdjTjhBC0+KpDoyKOWhoHkNPnWgl+NzK3gzIPsV3
3GU5vuyFiO575BdsU+iIr8VS2eizJE7DtXxWcVuZARh7GSbkUmr1wEgybPktL4sA
HcKMgPZr8sp7ATX9IrwaKHtoTfzYhvGPgxz//LwJ/IbaPzjGKx7o/jWZyoF0Upo9
xXKp/KWvHtTzfEPmtwyh2oT3jJ8EfZvxZvykZFDW1P3iwfbw2480f3u+FpGgGJ4t
oEBawElPK7L7UOF7RZVLjl/J8ONeyUaM9CL6UowEEQM80P0lDTNu12zbl11PtEc5
iTTADVVZzEYIlqwfnCkILVgzPaFJSJgDyq0oVucnLqUSr7a6/pMQgstWvcj9pirA
1+YulP1uU9ajve3IsX+qj4V9Gew9dnhlPHU3mCg6eVqezdloQKqw6RVvouFcELw8
VKGxtLDne/nM/CBQUQ+/4YYXHPkhXMcCG1q5wyDVCMPq6h06DJ9w8LAgifjtYmpu
LxcFWg9aq+E3aoJ7xIavsaA0xiJAmdVGYmX62+4D24YxtvZKNhY48Mf0bLHNbsnZ
h7eK+Lxlg6RA2by4NeYURxA/kFZGRfFFSWpGmxGAnFhSKR56/CSfue81CvDqRj/D
LuWw2hdGroJmjDVJSUWvKhSALFOwQKVMzKBR54EWo+KVyGLjYCwdZ9esFfHpYaIm
1KJnNJPMWJojvEyuhgxL/vpjztBDox2ncnf26Qh6Ai+DSBpi5TbghE7uGjnWet4b
x12JNs94CUfpW4S2n4mGwrRmnk8SbylBtrupvItcm7kfxep8bayqi3V1rvZw6z7h
N1RhYrHyOmi9mq0sOzTfBjaKeVlT/gj5PfNXEXPI0uai7ky092HxILEWh1LrRGiY
WjLylIew8mET27htFC68IqA4HxP0003dp9aMmzPPBu/6ZGx90ZE917aV+jOepg53
kP7WAzaRIo4Ti2wLBMJqsdZIuSGtr/YAbg7ia8e7g1Rw1EvubrhLh/F4Ft2eewkS
NcEZG7IMfcQtctxjdb9d3BoSLxsRSuvPXZGdp0akrClNgSnzoROBL/ShZxIOxp2F
87iR6zOaTajz8/fMcF/uLNHEEfR1YGDtoYTjx7wgAq2Huv+NTM4vhvp+M8J1Oe/i
eDLekylAGZumeddaNAhzc9mvWFXiX1cHCzck3ruxl/gzi0MQ2e0IFk0RG8ocb/ZQ
5zQe+yCfYg8n5M/mFEOLj4TyQqH0JHe+Kx1VzZgkFueIBoaJsxjCPDkqisgMtIfZ
xYvopgnYblI+8cqqLjkWnNBikpcRCxOOkH3WTuOd5E9MP+3KvBCi1Rg2DIp+w8aJ
0iuT1sWP4AjCIJyoQUoFIiHkh/QoKFmtctakEws25uQQDL+f+gDRTxSgG/1wQhzd
sRDv+5hG8XDUj1Eu9aDEvm2Excbd91JanUENCVnEtoS/AYDIhJLt5ro22N5c5SSE
AymRz6pfWsmtxHMJltYlbRIv1yrQeiQEY6/od6rvAXOU/hUEI3B/Nj3O+YqB68LI
8yH28f7e4tcj2jHeecq6T4kuK1sD3KVgC9+th7cB7yl+GmYwHyDivcTTV4xxdzXT
/Qd+J2HzUAiMdMOMM8jsj5tbjVayDBTy01ZzC8fFrHGkR8+TNTU2BOg1z5x+wdRm
uYN73WLByv44Na0pUw56myPAECA435JAcRzTyHLRCfY+znf1QfQrZtEFfpS8I3Uj
BJGI0aVsjyw97rRa2oNxzdrveGHz6dzCGzDylPHQ8AFhX2SGPEJUNOJTpXl+2Dmr
6145vrOfBPJgZHhLpMEEdlyskznxao0RwvXKFstIEFboTq/Lnr4aob6JOLD6Qhae
JUEU6AdY3qL3H2ewlXrTCrbvQ76vXuvRxlHuQlNhYGtfRF34vbiX0fksAYFn72IW
aSsNW8U8vO3aZlMu6FbBph0ffoG3/u+xV82d2Z5T44DXT4QFTG6SpuQPVdklgLto
tVizUi+PyTEjxh9JnHznKLm7hRlhEzhusS0efwlHRltzRNNEza4ZmmxnT8XuKqfM
rKhio5GYe58GYLXu569eY0eHflIRl6Pg8kWvWGZufndFLEAjSd2NdzAg16NLAB5+
U3ekPXXbKdD06OEr0bk+BWE/UuZFFHSmAXIo0sqcNsyflQ6WPHPCyieLQ0DXhHsO
39ixDAkJEqRS7d8tFITQputT7mqaLQDS+BhTRjRvGFT+QqHnRJlij52lcgLWXhO5
YHgcKhpcHQXU8Jkj+RQwqR3aRBxzd66x+Ws7oypLQNVHnAqrhtM2hiBaArpn+BOL
cXMGlkmb8H12PI/g0Xnus51reA2xo5hItcivaoJnjlaE2NcQBA04G0a4FvM+1GHl
wp+QGSmvKh4HfDAJ1fFrE3NlnOkpXPwM+g8j9JhovZI/FGPi4BXjT+bVDG9v5QTX
F9HyLKislGJyZjxlHAn/jrdP7kPH6gATLBZjDXQxJM2ozVg8Vh33tnA9mHk2LhS7
hO3bDoKF8glMrXDklWkEF7rSaBlDjRimUcBuZahGB9sm6qwIkR+o6Epj6uFQ5b8u
N5buWfHxXem8FsamG2+4neGMTEYXRpETL2z6V9ZXszJXCRL6n96ySLHw/n0SccSD
ScJGQUOyr2Ut9mO03DXWPSDsZvxBNPAevPQF6mpG9JOxGitJDVNd5JxlXZqt5Kek
4+G2FRUhRs+TAh0i4EuOUlUx9TndrUtiGnSJiGPrd0aChthAa5omePdLIRrlbb0c
wyA3hO8FtmXz1ZwhSDvWBuQ9mzr46HPXyLmnNhAFRPmKP+blJd3/RkCJ3rLpMCiw
NqZdn4x3S0daRKaEzpv13srI79yHfynQqaf0FwSw495GPT/VpZOfSh/+IQAiDTBu
r4BG9n2Mu/bEXhsjf/z0Ag8MjlRWdkEMlqxl0Zm2qSwjv4osiDHa6SAKVHmYKRYi
UjggcgUWUzzv6jfCVFw5juyKDTxqk/Ihd00gou1qZHLFw9dnfSD7Xbv09gF7Kh9Q
mkwYbl+Zpzn54+Gr19r1bKzcDGqCN039KeDDWg/9EgClvMkGw7dewJdcLTNzPmMU
gh/aIvCt0UuydaYSUljhgv5M9kMO+FvNlWlupoJde2OJGRO83xgVckprT7Lw3VQn
N76V2OpjhmWOIuH+7wIK9xdKSVnJQgG9mrma44VMVweP3MUCJKPTeGW4Ci0DNLKU
2m+2DfhNDQaFtuJ35VBOu0hAeuqaCuvf3AYkDokvSlGXHJ2V6ygb7Pe9/hV73E7o
CYoyDHVvVtWg7IxAgijMwWcYItZ7OV0sVzc5RN6i3rl2Jh+Ywgde5c4otz3fOXgW
7e+vqfcV9boxPEp9RWfkiC5pu2++f76PJ63DSLgzktoPa4rW1S4LMyHYa0d3hLxa
vj3DkmFSxoBMHBrGugeA5WWtph4r//sytAF7B1uZ+qCkQo/fHKaLceyXEHXeJHto
GWrQxeTIroWCEGkMcL3EFsRZT2rBUbweQRiolqOBujvQCrty2pEmpmj+uVwpXrwc
W+idmqjwGHVVIGUBOWg2I+BkCy20Q3zAS76vUG1FvNQ0H2wW3WDA/gWiQPXg5a+0
dSeAmlmYbILuo9hwFLBSnGVV8BzVJ1NX8/lzbNu9R0csOjvKUjYje7gIH4gzF/1J
rSpz00zLUnkriKA0QemnkdgGa48IaYFrI/f6uOiU6m1SfF8JNHGtMQ2hEqQXjmI0
KZ/9YDJ0hg2Wbd7mhoRPM4O90WPW6dCKv1pz6YUW7U00SAlF+e+m8VX8B4S7ivP+
he2BmH1TxteHbzEbWsw5S0t7q0ju43Uju6GZgFdMBZqbat4UOZ9x0Y/kKbl/V6LX
s0Mpy5abiWciTYfJLZt62d0sAFznytArhkaGTGZ2qV8trGS8lGx9c9M9hJ4iezt+
kECOQjvBlvcBxKLdwvssLPfrWYTWzr1cyroeRf9REoyFnqK202cKiLJxf8FgWSzM
NTZUmMOPC5rPryibnNFYEJnbL5+o4ueTfieVwQDAGr3gM35rw4aOgRK4lT3AgXp0
ib9og88Jr70t6cUjhoSEBgwciVmGrF/TIZjzAbn9suxw2GopOv0gNfFK/X2BSIZR
36k1c5AmtM+sHgwMCJ1De7ca/mIzcNiM1buwbpQSQJeUxsW71LNpHW75/sAdvJyK
bLFBOhIQ2sFzSSBBD0RX0yIAHkGQaKm19bjKlF5lr7lUqZO8SoVBuM+D6HhheXk9
bogYJQJ0ipPK1eyLj54ZjL/qKvvXw1OhCMsoROPqnmH27GBVJG5HXmiabXhguvct
dJ5UbVRMVfwQeFyJox3qc5Bd7fUpq08N/5OodsM5csgz8GpfqQwl5SRF2THoWlTM
t0O/sXhhvEb7YjrBwQdfUKkfO06dKbig1hFJcW8QzFNICHNmYd8EPgXcqlJcsSh5
hv/bfwBJFptGA/bmDKi0GIpp/q+LUgtcztKHKkPkAdk4vRcNfqM1JAryENjVYpw7
o0mkn3Gje1z2lJE/5WkZ8Ad0H1Ig2paWe8ydQ3SQhX0e8WdUwstAYMoAgiwJOecx
emwJsbiJ7suhg1pX5oetSY6FT7N49wCgnpuxOtQuLajegAkfRoZdXmScL3tycPCA
7Pusx/dINwtFyhn4ZpPq7UIBxstbxqC+HFm+aSxh1FMb0NF+kEPr/isueSKJSDH9
fUcXQQEkFTBt81YwLgM8zUIs0BpRX5tphMLW5p7SDluLTDOrWaIoYU/D0MKJlgLB
M5uLavjXemhGeGM9UagP/FNO3lizN5VmhgzmjrOTAuYhCV7nair7ZUqGWtBf5COJ
sUUGRkPEb91RezHOZx7tzr4ZEoRuihuZFaFA+H+WEbhzvlZ8IAKR7pQbtX45mssh
7NwffYBBgYpkCct/jqPLuSFPJGFjTDjfGsJsU6zHeNBdmOuuBoCsr16/X+EDkGuc
fBKdTPZIUogq+rIovKhXNIuwUz/3qWzRgXHf/0EfrrpIXnKSck/nDTQ2GT5z6sAX
dGMB+B6AJdIjDT9k4/3HBPm3NaeJPrWs9BEnS1DNDObnhFyUi1l3mg2HjcOQr7qO
/CjbgSXxmu20SIUtbVteWwE8wiBSlGggRrkihVdMoHXUKgG8WvHud9vT5ozXsyv8
gzGuQG407UzXH9drJn7+NxjtvXbCeFmk1fYOvnAa6Gd0LNBJHYCc0cnjjvWEAwA8
AEdsN47LQxKiURxLPATVCpUHcozy3NPeyex0wsrhF5NPGbdcdJD+/ebVIo4A6kxn
NgJfQRN5DYWEdSK1dCl8UGGwwI/usHrgqJKKAbqIQ+iTZ08jece8GGEbWEXgR9K9
k5WZjJm3irb9DiKUUUyes/pqOThMuZC0zbmFwqxwrlgvagGYwSFEFZ1JOCj0snjw
Gp31l2PDimHufrQnjO29GlZxY1UzMbig/Nzjj0CvxVWm5/zIJdNLwRUxT/yzCqxg
wm8MhJondelmVdPa5Mkg+M8qYZx7bz4+z1fpw9An1Kq8pRtnL1+29ICqF0rUeleY
B1Vu+MRSVcx0IafKdXASiGcSrH+yihQlLOvbnzDS9tyUpbKPXs/2DpDeMvRzJDFJ
2RWkYcqNBMdEn6rufRQW+yM+91s2XQy9aZ6iPQDF0j1ETxZ6459TMBpCeEGmhObW
H2RZFNKBl9ddFiaYyUBl6iOAs8zsoSb1lg66l9bMNzjZFvXbkDyS7X3MbNMD/1Cn
MsTkgqkKmsQyukNI7CWJXJFS7IIormQpxw7nJkht8tCSCapDZgu9Hncod/UvvZ7d
HzScGzbJuc5LCW60kvgXwhWztJxEs+f8J/n4xWU6XmB34qwjT61zobhsSXFI7dTQ
QHw2fdFbwIdBLeTWkFEFpZR3vaNoWz2D+PeB039DWZ3XFmvYvb7eipw9Gq8d6CVt
18whxz44PqkNisipqI4F2n/ZZjlQ7oaV2XPBs2pXzh+ZH179EV9+RfMnKjOtow1+
eo2KE29s9zdYqtu1JFZajY/YAHqiIMYmdaW4ibkogjxITwO/x+XcEFKiRGUYcwAM
SHVb8tABv/rqN+2SjNzc6xqMvPOgTOEu8A8WTMDOU+HCBldYtXN5hS3Z/ijleKfV
0FKVQofHKT31YnB3ylJEumeU0jm/0/RVcf/v3FvCe6gdpqbYX23ovNdD8hb6yk3/
Dc6ofrXtJZ66brm95DjIl88/nzhH7YvWYbUniz1t1SnFO9yvtnrquy/UvgnIH+N7
sVoly1fKRr5ovz2SAABSmxXZMNezbJ+19m/DQjOJBPm7pSJdbIhvoBYAu23hMU7I
xHFm18TKH7t/eWuAbgNJF6Myqf6AkeNnrjo2jTTAYuXsjW6g9qPIUi/tOLPvXH66
8/nTzDNH+w8alWn+D+nx41cSPaCdJwanK8WKgExi3VmUHkjmAPa2eHm64C+o9pFV
3DKfMU8fxru2wmv2i9C14R9cOleXc+D7hk98iMPs0oXVF+lF5V4q/sOIXRpl1UZa
keTJRVJYgT0Bh0Eh+jqY9IoWqFwsiE/1AcWxT1H59DOkZ6HY2zrSxkcTdNT9h+Td
DGHk3pBRuQplaANLk3inzt7u2Wameznp3B3giiJmqbXv8hJKJQAycvdJIDpsKoAP
r2ee/j6P4pYwDJpuTYp4AS6p0Q1JmIFJ3aFlLprfeJ+XODr/n6ikjtStQLRJ+Dx+
sIbmnzqa2y/L8PkkL4bwNWF5kw4xVTfrD9qdyvckKDekzml33wDGKEP7gf/vLII+
foyJ52FPZ2L2Tjt0mAExKJsfK944wltKZxUHCvEsCayfLrvSjzqMfTY6AYAmtl5P
2GMY+twCN+oI9jyhRtVaQ2zzqTiQ7RrWWBAmOcTm+gjGsamZDCg+yRVJmVJRvdvR
wW3cE4LQ56f5RiRKOzOA6oNMxfpsXoUjJ2GYySPYIbf8grYbjuYfLUSUMl1Emh0Y
VIs46zfo7YJukcPqWrJlvjvhzO6nEO0LT12Y4h2wJ9hOOKEjDp0YGjdu0UkbA5/0
hdpG7EVJQiTVlgmS4oj6cotp98dj8Y29s2OcC/E2racp/xi5zzumbB96/cl+CjxU
BeQRj4PXo6D+mgGlxXyoDfB5mcHpjUtvGX++Y6glmGesik42MiMD2n9VCpK3aFrj
hxtRNDEd9jO7nHlJeuiw3T+hehS7DkNM3nR8f0o2yKOPvKV9LRgevwkPAxh/Wtmi
QY86aYSWtN336X1Di8M6TBg/21m5o0W67TaAyuQvYkBOjrOFNe7KvU7KckLvHt9h
reivOWDuUBMegGfR4fUxmNCuxDErogY0fZp1G8Q0jIRrZQF6p5RBvBGceZQAy5Ze
S9DClL6lWltPSy2PNx8Ppc2z1qV69IabGN2dPQZhljuK8bEKtCfrCpvRl/eKaFNY
N7TSSi73OF7aTX9xrdl/MdUHNK8OYmkCm7TOKfhHnjveGKa6P04x1zStrIyJkgEa
fbNUYd0knoUT6ItRAoD8PMYFVptT2MSeTlBZVyvt3BM1L7CwPqM1rYT4o+Iz19FW
JuF5fN0gcW6d/j0Q8LMHKIAOHBKprNQZgZ9Ccd471mSd4EHF86B/QuLvucbkri+S
X+AXVopETzLTplMUqZZwPUkH544reTdEIsCKkYVXv9MS0tZLaO/2smxOnTh5gV2s
s32ECX48sEC57J4ez6RAi8/MA3+nCl6GiUkj4+l3bmq+juAbZssCRQknNWf7mpLj
Lw85KKXPetohvf6ByAwsCHhYHkDLHXzfNfjzRRu8njpi8jvGeAfzNVKy1znWTR9s
4L7Jf42T65QHvlX32fRB1m8L59gyWoRd9csJVRfejYGoFhZOQ8C7gc/ygu/Hhhcx
/IlRdY9agxLJ6T6Xh7H3vlCY3ZHfA4WdHnaHkhppyd9RDCVTHIfcKESZOL7CiY5k
jqnKYD3dMIEHOOY8jRa30ypNv2DWlyUe7eF8TOp+UxiXkHBPI9lqR30wvCb/eXqI
lLMMRjLK568nGJjwIWhR6XVHMYxOPAxDJJeI0uCugqHgMTjdXMsXhzQj8osptSOU
swMk185U/+7+1s9uHzZjABk89shYrK5OmWTUY9otqng//b00jGOcEabZJbAD6oDh
RZkh+hFlnHPbZWDMP3TDRFxtyrz3Y6Ptn0zt34jn6B9Vilh7qhqFvFondPp0xwcC
fGSyf/efihPf/qaP7SJQHTkBFEDvhfuvx8woezFH5q6Q3HOsKtsfYeqFuaVjdP3N
XlOoJ8hACxBHUSmTWer6IYz76WzKR/qB+th6BIN6qcE3TrdCKOkF4qfE7eHdjMK0
G2J8t0zrpTcO0hZ83yAeRgCvbZlZKQfaAyG84D07OD/uoj4bZ+xBWt+2ecyQI3FZ
/NVaFvSwJfdezanbdz4oH2nfPoCdiBSiBCqAXeXkcbyRZO0xmcK+EiYhKFcEchTH
z9xa8iRWZG6Py086+93uab1lQEx47/Epx/XNvYK3pvtW7JpWNX7wk6bOFT/W0um3
R7seIR2Iud4jbgOcykgVUQVNrkCOrMtqJUyiVmo7KshukRP7nY7Y70InNFFeEQyZ
D4i/whpUpaSN6sv1Re34pSboxVhtzGs1SkfAV6Im/epH85999fBl3gp4Xhtjkkux
VLXHX6OYDxHmJzhiJbZ2zugwGS1qIUFh4VK/i4/JOxJ3VABOvp7oWaIFW1VTlrwq
V+Xql52wW67VNhpeJlVOa/ahZd0Yx3KV/AVabZUdcNjiGS1UINRaNapXcVLAPFO9
ghIBwuiGnGTvZPX4grCjCWrjz7mN+PC+q2YKNADTCIckyk2kr8RktuwCXGqi7c+1
zCmfOXC1mS0E2foUd3+eNhrXNVR3Svynh/ZT9mwSjtKeE9lqo3VonOadHU5HBVcw
/jNFI2FMKDFrlkHpf2EktUt0SIR2LINByz9IzYI3+du2xM5+yX0myG0tyZMoJa66
ceO93qHLUiXBExoaUmBRTHP4mOFZuKMzRbicSaK96eMlVCELDhVvkSY+JPJEw58P
MjCW+mRt8uXQtcphT7FcXWR17cDwZcLX16uMzO+0MaGKco69ju0kKiYkDaURZicw
HbJX3/YSqcwwawGIz0aMY1lZ1UfePMFT/4P8BaFzfovN1ArEnYT5IWqBOE0OIAU7
1x02piSIoGrAlDHNg8yFmblEEEqUCgRhyZmZfdEc7Gn2zwOW/fVx43cXXFygibGe
rhcxvO+YC06xZP4C/FvGi6n9X6QOWp/S23q1tf5uum/elF3/swtvlyLnFHGHoWDn
Ns3O9rJXzCOTjOGGoCuJ585WOJXPEmpFNaSapBL1zO7fhpkX4oUnOihEUM/CeMmJ
y2WDjXPncVXU5PFrUh1Ja3BH87uymSg69hcJl1Sk1yEcQOns1U6x8QI2KxJ8B6fs
rUA1f9ZrDWrSxijdKi7uVG3ykmV5qPOysVLtOp8lmoYFdWqVR8HNB9+SIUU49aCI
3+Y+MeCxCEzPfBvdYvaVpJ2VjA54AmVlqKDAIGc99VLRjKw8XNUyWUGZWITTmSSJ
py+qrYubcPgvnM1Nm2nvYTxvY8Tgg/oJFJSMiF6FmeOjMC1HcqF0IxcqaXTryPs/
dQ3F0TrqQdyMXII3dS3dIkjNDPWhLZMJvIPwf2iTmuCKMKt49mrAV456r+B3k3am
vIuKiPGLtkioYoyCczzNd3goeKfz/qvtvICp+4mGuElH1TGOeg/robFqSbzjZ9s5
rK93quUDCyamqiWlTd/3F0BYIyPWTG/6DrAww0sRHkoeXbrWSdM21QdwG35AI2kn
5qAn5ouVxSPXREh6IrMYvbNMu7m60Ki4zWpEy8HJkhdhGobn5dg+ZhpE4Lj2dhpu
UKipFRPTd2LJ8NBuvPbvxcd5ndbSMijtBUjOOHH20nZKIKlc1xcEuozJL5dvN4Ad
XztR5VsreYST4Jb4rnP3QbQiz8KrWA8mcxenftnzOGhksv6eP6Sgb52Q2nA4XmFf
FDZDqgydud9q97cQkYi1lvqFok82qrfzNu7O/+gIW2qYgMlg34vwBBoB/kV+8S6Z
m2WDn5pwXJndHtuqI2KRqF2hvs3r6hefPWk6xJ94qhdFTgmQayTaKlrQXelPpvJy
vt/4r/MHnUnbECIwMLBe9GLEGh5FmoJa0WvOWuN5GTaBz3UUsj0unp5fYHvV/eCJ
/WHd93OQA6S7PdMzf5Uli2C7+MGDoYpNTghN/fT58Wjy8/5uMjQu6VzcGnkHswHt
efyIMNnEmhWjdHWlVBHxn/uIlacz3dxPON/y/RbcofHsLORKQwnu8Ax4AALbkSot
sMehCZAM7dY0B1blcpWCNI6xykcejioXh84y/ToW09svTTxtilm+pzzNc+1+3YHc
OHf2/5DQOwwq7qzhOfD+a8+JJeNb74JSA7QjrIqTtJaMVbE5wOKwgtBf2VD67eBJ
sU8ID/4psX18B5SQAOTS6usTRyjbE+sVDx/GCLFYEFLtXX01KNtAKUIkWs6c1CYR
NdVZQSOXT2MFVVlZTUP2wbweuTnXzlrHpQUmRFhvNRT/l8On4y/TJ18AO5mvvHPN
CWuZtG8sMJRXGok8sST8LpmJT1ReoSXmY2Af70FPlDpmqPotPsunE7bN5/VezbcU
ZYYbMH56DJkPzIPQ50OGLSFXWuky3MlfmlnLyMgFaYWcNx7/KAt1ljnOneS22OPC
g81GRhlN1aFlzp31brLbXwTA8oMLGbCb38RKBaVS3xXi7Tf9YUQPqE6/6R75nI4p
OxmEyUOfl5PvHn9WdXQL6clDYbjSEvdWfynq7EnLGASYjcPHCTlc/3b+9irMseiM
TX38yBIy8bjTjfCOfBzdHSOiD/rIBZ1vLo8HZ2BFhhX9fiBfzGjHbUle5HARsv3e
ajA9BFJYFnNh3rvfHYKOWy1QYifpygKCBkC9blaMpG+MNg+7MQzAXbiRy4GJ0tCM
HhLdMeA8Zq7aDrBSZECfqbrTMAaKlgGTj8jMTekHvFY1eiPX40dxm9cP4U36xYNe
h9mg3werBKr1ckTkpKqw6RVDRdKWON4/GkBpr2Zci52Dr9EDECNUOPMBEj9LBTZs
kZw4jJi6bueQ/IJQLfcuA+dVpVaHFXMjmgW2cLFg8mg1+iCgvVzvM34ld0q4qQS5
QgBBabnHUXTSh/pHDyokxuFqwPjTI7VZ5u2otrMwT9OK3EqhDwt9RYZ1FiPyFbaG
riJ7ndZ6g1BF72avEm1S7RJx3SCow6qfCpDHwWYofBVpGh+mweUAP5gWMoGgytXp
IEZmzIAOsQ6J1tmLEGdtJ9N/OR1lQY+cbSTgUCMYq290Wc9g4Z4oNQIw4ecARwoN
6Rxy0GxlQu7d6J5eoIs7diLY2Gk68Z/izOPudfVLfz6VRTgcXNa7vynslbqfd95Y
Xk7ptuvQM86FgTMZeE2WYVzCY3o1zYKyZoOhbBYb4s0pj2dzOmld7dcEPRYRqV2m
W66c3RWLRbMxolOqBqIXacJ31GFei3WYt+H133Dx/mWoAqAwn1WCSnkB/XcaIlTy
fGhiD1OauLnCkM046JePa9XM7LgFLpApsBhw91x9l2r4TiWXOLsyn+1Ivq0VFC/t
GrToatN9foxN9CHFRI5EN8lv1fhhQBuxK0BfHIteEs5VgqoJ+KNpmDUrq3Amfzr3
TzAelgBLn9IpLX8aRa51TOKI24ldQlA7Qhy0fB8D3x48Hqog517c9kxU6YfHPa+L
gorfZuCw+sgZ42AvRkieCFiVPiFxZPZoQowaQCid9wJZyDY5fuxFu3KELmXnHWsj
7UB2wirKdxw632sa2S6o4VzBUKYiom6LARbmIo4TwKoadGXOxL/zE9CqLD0WQ1/h
46JupTaNWIH86EzOGuApRHJffBFtdKiIxFeEn09aYodPkk7Ju6RRnRMO/Wv4iNTf
XKqgahlj35P5MNXwWIZuf6mZfh3w8UrAsQ84YMBZcte6RME4HyQ8FJETjFnRFXQp
gVNKFsxTscKhcdsUueOojcp1Q+PUiUwpEhwM2yj9065PVVEJz5mJQzi67QU0DkdS
vFrZ340SbpOLp7rDJFS6FRTFeuDIQxpQ3OU/c6t//yyJK8hyNubjBfhjUSOTx1RH
xUgsHfK/VGP9p8M2GFgBInx0H1d4NjbpY0yrysftQyBBhkzGKHiYkr10B5KTOSq3
bCCxloaIkwqUodP/AG8V6sLYGx6NxcMrsiF1UalvC4mzcIiXSWRxdsKIepxO82Tz
aJc/EyqX1Ldfxc3fkyuM4kZVidjTYjBG68dRJBr/VxAbIZZZE4c9dLWEGXXNakHC
B2qQw7iWBpk+7sMxm+Q3SkqRBHL88Us+cnIeskoU4IjWHGthJMQTZAsvn5j0SorQ
eS25ZLMNFHwGDTf6MuJqpe3sZI6oIGH3RJ7c/ZC7NEGV9XX2wOi+AeFRA1dP1wsZ
nlWH8/YmrLBMk7JL/bLCttKLo9HefgTLjtaGr7QUiDANM2zk57h+rwusZ9FHLM50
H8nqNNQava/wiYR92j2I9zEipeHNV2OExTtxHekBkNOMe1LXS6oxrUg/GZbWlY2H
qzzhUxEfx2bCmr2/Yiw04vpuvxCfawrCFXHbEOJ7xRx5UNI8S6W3sq8TmuASKASO
tj7xXdKhpK6sSq1U9gIHNppbhEDqXSAeqgJJEQNSNzD4estaZYMNkAy0lP+ibZph
a0E4dVOVedQITuIaQo2+G37R0Eci00yRgxU1zAS9sILXtWPB6PSrNWLXwO8dtfL1
n0ai6hlm+CFjU6UmpRawxUj4MhcwHA7QxTy27a8NzX5tQe2gRFXEPCU4hORYgsUC
5NpyjcyAbVovJUYc72VSa4sV21voM3VwdJfKdlRvckqdyLUDI3/TqL3BzQocvhxV
TjLP4zcmDb2Z/+YLMZp0F7ddJfLEbbE3PHFrScwDX3nd0AbzxknREeyQOVPYYKJi
y+odENK2x9+VBgMIce7sm4PLF45eGoXbnSRhTFCPczUU4NqVgroo7KtRYKTwwYkC
Eb9ukr21NDmT3nFawbHjpxdV4p4+GPD9Q5I+4kfvzJIO3BxEWRF6ACrUCoxGsSgj
GxRBayFvvlWHKWPyDT5Mu1sxJBR3QccgrF2FlGdTqC1mtl8wpcuy/iSfyim5c0/v
+Eoc3fBarcTWULmBq3w40OO+xWvzcMkLQLeeLTxUFVO//KEyrUvEXkraxugz1hps
XlpwraXllr2wj/Rk5gyO8K91uTjgyie/W4+dwExczzPDfQzNhmVotXJ1Trmuo5Rf
Cnmf2wvaoLxGipVJT5qzQZPWcM7XrJt7mtyyv4AxGriRQVSMmvs8DcdL2mPe2/wl
yU/342te81Y7pY9rz0RpiZVLh8XBooz41lmOC6WU4WFRLAGQVHV7fSlzDwQ9AgAC
/0MXL9aFyyyRj7BfFFIDVJlygKHEVZ8hYzvhhu1PGJ8cEVt4wqVwoCo4RfZcLsrr
Ck/0XBT84kGVSrnTjQ8E4d3rYJ3qBVoUPJYpkiP2uvg7ewWj4bn3z9JC2bi50Z5f
HvHsVP4qBvssSVJoewe6hriOUAMOJkm8nhhHb3yh/7rEQkS26LEY8WWtuw00BnWm
0C0hahTDVkZ/taU8vZWSjdtGY1q8IGrPWDFmEb6X+ZA02ctpTL+d3NMqVbg7DzIf
2iWZZF3tGsfynAkGuFsRE6vseE+uBMYE5/vfQXh68bEZ7nJagfcqPtvM6hYh4vw5
CKFl5SbqVvcXL6sFRnRxxNRttZxW07KZDtpZwMaO6NRWcBjh/kuWu+wrLZLQEVdV
XjaL0nINVREUd+P6/+/chlTTmJUcTHHCroWf+odmNoJBpRxuWWS31Bc1A8FneWiV
MOqJtD2jKslCeH9E7fHvm04qgqQ/WrfHzgx1D99uHXHr89qebgTzm79y9XP6U0Gr
W95vzoBOaGqAJ4y2sQ1IcrK7caKjIOOHPzvSGD5ShwCDkwPssIyW6EPpoDkztXsZ
qS+jBx+XodCml8o2DC3Dfbc+4lE+AgJ1W3zyqmH/ZM5gQJob4miDMBlVOMnS9Ckc
lGNBHx+Pgqqxo35FKPFrDBR5eoHso8t7UF3vr7jXwmRxciGTC1ELltgaWwyHFTnk
7YbDf3LnHsdlvmxqWsyFdRTSV+R2DtwmToFe9MAlg4ipRBgruDu49O1UDaJrX+eF
q9V8Ia9KmYaOvkLK6WQ59Av+3dGXKTv1lCWLenYi9CFX9bNvPAyKMkZn8xj/VsSz
LuNN/zxwnUfmC/MkKzvbXCbhkrwssWysZa6We7JRnDVhof7uX3C7W9rndhZU/3C/
1kjgx8+cL9oTW9efm9DzaQ5SDVXqj1IORWC1zF2Pn9Ul+FHRe9n44ipEMItkf7TK
lHfkGq7pFMi6uO2atCAN9nCnRJgw+cbYUHNYv2YPlrFY6oHTUotFG72kSi6vkRMA
m4nU9N5yz35MSzw3MU3E0g5GGhyKDw0Cinq/cnSSOk6CsII7u+LlgFnb8fbWwJXk
dlXQXJj/AVs/azkWesnStigdFXZ38qHag/weCqdu26Ju5eeIxJ9aolbCtWtjKBYO
QokNmAz+NNc+EkN/QYHYomyh4QwjrTQuYARmuI3v7/ZBZPzrVRStyR4BqM8vSwPv
dL7HxYdCoBXelycEmzqEgcZZlRbGY4uvX5PBSR+4Fp5bHHZYAST2uK8zKsrxJM99
nYd32oHU1RWTz1SmCobamrksBgvWTQGL1lKiQG+4thSOi2B+5d3zZPqGiOc83OnW
q4th+T7wu71/mfrrgXWMcRuWI8uvLtz3oUPU9ABQv00Lfg+FrWT0TQhFjwcSOAuU
tJWJ7r505TXEdWNHmmDKVPYXyU8FoO/DrIOPvRs74lTZMauGhnyqM27Mpfk8cGUB
j521IlK3p2ybBKhjqS/39pCnd1RCqXKZIKd2t0G6cy7/fvN+LJsT/+uFV6Er8Qf+
aeQ6FIJaYx85ZU505yFyq7iaWewk68UUzG3aZM4l7CtzVTjNtr4dT7xuFhTGXDu9
mpCF88eEu+tAM429i7kzZKgJE17R6x38Luhacv6vFEVrl4+1EiEXpbB6KZXJbT3q
zgz3b07p9YzHeBBiQlbPl6OsSFzynBY+kDlKeuknfAPtihVeIKG/hKPSBzjAwIBA
wMwJ02q36gNp51VfmVSU7UQs4XfAwdIyJsrn7RSdMPhbemxefpAXb4T5hHQ+4JN2
ZUQuNgsA/W6A/E+e/u5ONzDWx+qT2qpC30xwLaY3S2LnSZ0jaaa9onr6bzEs7b96
FVkQP8HgCw7uGNqHRsY2Pz+uAkI4j8umXDfmxcklkLdlf7ZOUx1koOxwFU5snLkN
EfWt8UHdWcKnAGxkt64Byy3byQuGHOXFoZXG3nr07Nb08A3OdOS3TByhhD64ZI30
1k8F5KpexzW3Duu3ABZVJwkz3kacpyzMVsxg3Q6n3OOPO5an/s6/VUOhlVEF+imc
cq9M25ZMvwR7lx7DXigf4VuFem5b6uZMFwFojKS2NRwucN1OPgUy4pzYK+OFYEwq
ahnwFeTtxen7xC4DzMM594vOwu22p4KvW5gEjc/quTZEgvMf7sPLO5VOWwoo5qxs
eOWxilwwSrUHvpYawcsjYSYuPC5//gUeqxXnVDVBP4qrbJxR0z2a34+iz1XwxHWg
YXZOBZi7c1cTFO8B0Mq9JHoL8KDWIB21nsuAb4LMD70LYyV9Zpi4NVsovgPQLOa4
wgWPN7c438xr8FYXK4uBIzajw5iw2JoChqHCTnkfo1SM/+Pe6g+Zozi2Li1k0OFD
LWy1SZtgqZZy94sCdH/78vpbdqcHujFaisc3qqhx143eBlVaLk++7Kl74J1kjMU/
YJIIChu3M60i5dO6l57qB+q2OHqFt0jjXC7l93U2TiG/OhaRVZxGMzoucH/7HtsT
kTwnPNZav6Hj6nzQ/rT5qcXMXdaT4iGKEJrsSxJqGuPcjqsJuamr2kqaucFdi/Sd
n6JV6mM7i6WNZnNf1Z673kSrBCo6HB3m7LsGGIExZTU0556I/oUCR5ojqMwsbyun
8iQjQlHhR+VTnMthzWbW8WFnt4hhF+bQWw4tWTXhfF5dzUE6KpWcYHPBlbbj8TSo
qkYeF7YaXBweDVglsCyb0fEkEyll7ZrUiwIWgcI4A5K4B2m7jSvYlg/9SQesuHd1
AfmGlOYX90L5x2gDQs6nQByueRFUO9PgKSa4628avZi23F/0XXqfX4tYEPzROsT8
7tLSbw9v97E4EZDlRunlAyNqTdWV4IL0k0fPGgvs0AwX45JqnjTAmBPtaEOVDoU0
Gk8lY2bBJmlVMWZkDwcKgad4EsMtKsG90Z9x9a43rSKXFMkbJazH656lqDKSPEN0
pVIDFEh5OL6xrwWuHdO/YTafhLOPvvWze5oHI2vy/eJLmUPDkLbyu5+lE6d1eDru
2MdmDlebFITDiP/em82TSo5N0rayflZ3uHWCaYDuxa2lGjZD+efD24dddNHhaQvJ
tomH0hnmtiEDRuBOewnP0d2VxNUt+f3vP2iV2qmrGFy/c00sPSv6VN6dDDXP+qLM
YqOZjYn1LAap01vamiCeBdzURYjrvuFe/AoHHxg2zKIvTtXAQ5fnNgYlApRQh4Ha
bsP9xellxiTsbf6PGZTeqkGrLkxyRziWMiu9p3vRV0if25+I3ub/bjJij42QCRbb
FfZGZDU2Z4IVR1fkBWy8oVzs6o4LP+H+D4X7Q7X8QThMQHRuWHnAcNAjGEwlLLbs
m+KdzGgoGmKA/CG4OH+aqc2Zk6B3x2y7x383+dUz3s1pJBatqqUnNHO30vhPlp9x
WIwVFquvxNoPdC5WSQnFMKGyntYgOQ0t5zsJxuexh9kHFJvzPA0TTxclt3iHFKqD
5xyjGQnhPY35kuToN93AYYP3FBbmdw2A7Yg7IffrOQvrRrOG1Y+PbvzihtaOooC4
fe7A/XL8vQ5bmLDcYtJMFe+cfvqH0aIBm43PgZfLIYJ9nohrpbUhYrKdBz+HdAEa
Z+LHIbgYeHKNVNTmtvOyhSmC/6+Ff2eLNK4ToPO7Q5yhlUcHYqjdDAkJe2QN2bMV
xq19ypK0ocubglTgp6GlIaou4tOFYrJU88/HuK2hMhJfsADMLf+8UaQmEq9et1Kr
WaChB1WBQQpyNOM2hOGKLwKr3oZzy8Zy8+Kmv4r/K7APgdkFsDRImZ3+q+cFdjbq
yPVVeEUhqDdQ+Ar70Fh3KSNnBBMWmCv2CGEBpON611TJjs5pu3hzyUm0UW+Mm1Wy
QFMIHCSor3Q5wsniBl3haa2sZyp9EWVWYeQ3Fm6ZQYo0tjn9PWnHON51fzdjFipW
RE+sQpibpVqTXvOm0LVL8o4guEwgsoBBZusDqt7UsUQz0zCVVG2LqWodh2u04+Sn
ONh5UL6Ug9sQhq9WYyiHnfWIMWnWtG4xrQEdpTREDnOqWHuKm+b/y4oSLP/+WCAU
T4bw+6uW8rjQo8LsrnLri6v12SSiz2VyRnMDSZp1P4+5zK9FmntfQjbShgcZ+ZuF
q6KbaUsvouN4W4ZbIBkgbNZiZ0r7aS4+E5JC7SSPrdoUv4A31DZ5Ir+QDEo5ZCmI
JCGEowJ4UjXHZa/EvhiVpsnE+0UHk5RcXhC7uDNZmn4nGO/2BgKYsZVIltAftTFi
tjlB3/rOJVZNIaElXbQ75iBD0m9AiNYoj7uaLiRijm/0niMEXY7JakM3/W1EN7aH
vYl7LKMrYrMMyR+7rVY0sEC/jiwShDBIiCkznpdybJCL4NyL7ZHIldo0X8G1dUvI
ujLlMOJpPEremHKU/OTyNAePSzubme11F46KsJnn5QB6XbDKVvVg2dpG9oMuSe+P
Q97OSBNahsKeb1HftyiME6efqt88edobVlylP9zuT3A0EHHzc03IYaSn6fZxGq85
ZM/ntP6YQz2FzglR3dK1r5/ZzHBjbtGUPIeeAKuyI95Hw0kqgCg4y39s/VWd85nn
hkolrSsPl4qOM6DnpQSf/GOkd+Ts3nNgDNB3ZHIIUFtsKGoTPIP1uUbrY83OhLCP
laSA1Q7ML6o3H2cREK7t0utb/BxeNDBHXBQkrVolNO+UurSHj+VKiGbXlYxLXrNo
fmAIwWzwNmEBe1Eb6UPe1RaalAv5Nt8x/3mVVEwKGnXHOW5FV55y7Z9Nt6uMfe0d
s4c1olhABhppDE7+HOMXAfHhzjW3FTCq1vCrti/zaUA//SxxA4nRTE+IGDAvxCMx
dAqZv1uzJMY7yquwi44sWyF89RgHq2pH6mnWX98H5SAhyNSgWLH0rqZelpJrN/eC
/ZCwus4X/pLlKZU3hL0bpz/d0cIVDNqtSMSDII0LMmSvf65YGXBe1DWQ0cHINw5q
2bbsIuWNONwBXIjoRDviMZJy1jHrR+KolZhOWwakLq1q2b67mGSuB9yC2hnK1Cuw
RF1UrtCjlQw77dZ6XoyT0fI4OTXtRgXdn9pJN3KVqxnkrcY7Rgx8IuECymKhdRvd
83ndRkyfMeqdsvkVJLNuKx/fqQImG60gO4WHQt2DmHrGI+d10ODOjsSr0DfK2z0q
tneRmOZE/ys3J76fa6k3h/sEQnIuuK2PS/NSOGHRDjBmrnu5euj0EGJZ8rOxH47+
ziSicelQMxLf5RSXxoiLcR432wXGCntFsLv4oZ2HVe4stc6O9DMMb/ZrWVmS/v2P
CYcQMvEInFu4uFHAaxIZoqnwXwNiGrUgOlTwytrHnsqhfqK4A11C7Bf6YBv8e2r/
8tUK4H5kBRB9CNk8RHMb75ceVxD/7dA92fDPt4Rp/9pp0ix23LUEaoQNQUUkesr/
XH8CJSZPm2Ndm/LypO7SF7tUVKduacYDv08aXnc9xuVIhauYfSUTS75boOOdQIdt
F7+YuR7ZIvKF52aWDzWwrJIoFqfBDvx15LgCKX8lpf2m+OHQskumTyy+Bfkqj6x5
8VDTFWbsbwxdlZ9se8bWRw5cJm5sxhvrSFswI+H6hpx0jj+u1Lm6uomuA91ThRhI
OkaUs0gfaNNIbdp0+QrPmIUO0JMA5k8b/Evq8i+LX1iSDXQh616kf3xJHIjNwVf3
nP7e1Kx6Hst8D/yRYcmmSjmOn2OMg8KWzsRZxHpxPu1kFi0xt61mdkD3bIfkmZ8M
Xe5/Y8tzyArc1Iab8TuM3orJhdc59s5E8o6EU6PFABemjP2YMJipQ8bplDmM6Sx6
PtBjKSN0BJdjtE8Ii5wF/4DXKrFHJlf07CYasMqmGQP2N928+ilck1GaacOZ7eEf
Ecgx1D7XLa0ik64wBYM2aJ3UuvMk33M4iRbOPq/1sooppCy/GjPovrhmtigHFSaz
vU3ALgPsfB43MzihGXJiQ+wWrGU+4BnV3A4pZfb7bMf/ADY/4W4Zu3W7XbfqaCeW
aZqiIkxfbys+TEQxFT8ypbGlX+3bZExQ4GqUUz8foqbdfHatuuuSrHPI9KxcpIJG
Z3/4Do6BX6W7yieXpPhUqfbcim1KuEtM/cC2RQXwFOSDQBere/BruhWQrNF/qI9k
BEdfV1Z8w1zMhvA7e/rdE5h7ebfxLZXB4SFdaR98i+pumHpMeEgTkMAY2FOwTiWo
6v1CPLygouxdbFBKyH7KBSkYoo6dl697Myjk0spfQ1pc9DGkeUKvZV7+uc/rnmwj
a1mkgXbpfabmN4VnHmuhLcR8ODqYEB1r6a+h06uGSh+4UUs3CKqr3mRx5UDMduYc
TkrSQrWE5GE6SxnhyQvz7nbhTxjwW8UbunJ/TXRRBwlV+n8I+yUkIwu4Yv1hc5yk
tSjTRUlLOLYXQgsvllK/RXQnOWZT0gHm89V1UMu1VLoLFgbZ3VWOiMCxgraVwg6z
HzzkWENa3mFIeZXxctfSPc2kK9QRhCC7yTk/l2sGE6M+WPPQKtab/o/3pFu9i8aq
uH5Axv621bEw3djnObg4Tc18NQtuRM03hs082NHl1gs6FS26NLCvmSrWAuQoZ+n6
Eh1FiJV0vSp/jFfQbuAkNYVQ6g6jruEuIsN191lUHvNJyMiW1IQNepd4Eu/nKBFp
zlEofJ2/QJTTaWlnyshfjY1793wySMPsWjvCJsCbIBeizt0StYyUG+8vbTyo6i7h
KNXvfmF+nf2lxNk3wjMDZGmtBqazGPu6lMdKj+tH0MdlRvgCLw1kIXhtsCgWFHbp
KyuB1bvZp/kV0M0k8un3Qg3aZfrwTNWY5TTHrIN9Ng9YlFu/Uxjj2A7HLPU+WcLm
jZGQYdvmxuopwPP6dfe9zpXqKrbCzG8bGF73lWFQLkM1pcYlzZBqTbxvn2OgzQ0C
HjeH/FyJY6P2QUdCX0hwSaErWtJQL2hSZECL68dTzwWXCHFt9K8ogMgvC4TYaMET
nk5RbacLOLAOgfeq19e3HuqLgvVgEd46Ne+jZ/7d0bcfGuoljyi0HeqPw+EvF3Sr
465DzZgtvl0ofz25r9vmCBim8zyh0m+gBwFR0rNXOhW142ZLBqkg/ZbCSsvj70xp
mnBoLSAf/EbLtPPLzsXXDjqQHzTe9YQUMp9IO0iSFJgHUpN3dGgMfSbxhYh8CCry
uttnYi4+5Rt8lwjcf5ww6gdYJ0q17ySiDnyZJGIdrRqjWT74siKi2QZTbIpz4WQz
6HSgsjptFeSb0GOssAFSG7YrL9vnX6ejQJ5E0YqSukIHyaDlq7SslQiOA7y21gbX
YYybSdZ8JkghbG/KbqIkTpUrk1LMObcTUlysxte/Sbrra8fq4LkXF5Z3r326+PqT
g6Piafx7kSgkWcA2pidiMFqyDfc8o5vljaz5d7hN4nIL3mB/9AYCjEYfokXsNwoC
0Hs5eFseZmQjlsKC7jPCppARrILJwuqkJSkzjzTR4rHRM2GAlf568diQLheW8jaV
rR02ZMuMBsIBVBIxqbFswNfGiutBa84qa4BXbWqeC89hU+TqeNhKCo9eh5TZhNZ3
mYCZBGWmkK8t8cfUoZ9nzWR/aLpkkUF+LI84csfBGIBpF+vVoSl5QRZVILnISAYb
zv5v4DggP7y6844c7N8Uncv7nZj/Ydfdvj7ustFUmsDLIktCQu8ByLtBdAt+JyER
z06NAwj+wSMkfUoMueseXfIoGLNuUnazDb+mne8dYaFjmfE2rbW60KhwEspUsqDT
BEs3b7FebZUpj4XxhqkpRe9nNaLXPO4b1xQCOPWL5USczgq/Mk6kibM1m/RS9Kbp
gDDnNda1nAEC1voyHUjzmDdz84E3grsq2Fl50lHF/KP7b2uF711Z/8+EFbB8GrzI
oYCrvd9bRs3Ah24XEjRzmeOP3sR6ugPDuHFPaReMoP1TM7p7sSbTk1eg+BiY4mH3
LcGDuAYXcL0UmPm17rod8P+GIWqxu0clZsB3GGQjelX4+j++Y4aXgHFvNiBvtrTV
u1/13xm5ieh/FvQNic9vDHjUpX3GLlwS7ytA8KB8E1xqrmeg6/J+E+c/WGLcW1pf
nZSvy79UroJcVXkyMnuGfGJrBbualuHkHrfVYPLax7wABdR85ReMpC5huD0WSPU5
MBUB2H+6yK1hIzTa1pvI51YjJRkRSYr4FnJ6x7RZNmVyD/nTsvLYWCmU2Rouj5m+
uO2KkAlBF4/ulSgZTdFWhq6is34JmeF00Sa7SS99kj5ySGK4KM6z1YJANhnPZtcU
WuaDGOc9lvqXJh9xMURaay5xF+lE8AkFIgWG29VKsXqCgwNKMM2vJanBNmflpbSK
Rn1G1r9cN3uJrtFA+DHKlMzCMi+xKyBs25BgW3eOSzTey3Bto4x1Rd9pLpMkYj0p
iBleyA6bsTzl1eazxKRb14Zr439ut1YuN2nkhSevFLXmCPlDeDfFv6ud9LwkJKls
6BSMg9jbKa7VPJM1+6InBIbHdBJ7Bd/bcS7jUt02SI9Ya5lEir3SHOLkhkoe3hyz
ulXkR++tOWfjy51YHMSV48GCIQGsJSR2ivi+HTmmKt53PYcshLUuSI9qB5Lj/fZu
1woEV0cgIO0hugLQzkoKESsJoMPSEBFHsHCGQ4Y4zNslBWyFTmc8vueFwTPclqbT
v2fOoVq0pVCundXOCF7jMwBq2tT6Qz2T8jIWlyBKQyhtWHRr01Ri3PVDXvjq0bgF
+8MCD9sgxtefLdAuMRAp83Yqrkg5puCdSeZpPACm4Ulj2gXozbkiBwoT/kjz8DZN
nvrYiD3appyE0LHHlhDy+sYMjj3PlMHVERNtUlX2NKbRGAvkUPIlMl6GLxDw8kta
jtJKwzdvuii2H/MHWQzlaJGzhDv8Zx3DKnti9dQWDOTufseSEtTztvforyLXw/7o
4A3H4eI/9VQl3SjSvYlI3XNqDY6fp2xQ5Mj2cN8T8xxUwBn6GU1OBSEs2qdkxzIx
2dWoFQbgThFqCGh8C/DLPCi2zfI4/i+TnEfmZvPcBUm8uCfKsGrQNnhi/1p32ybM
HfdTa61J1nJGRn8vx5PyMQdMHwrIPJC0lku4IxvkFgFw7ndQd/8yi89fuhEFPnpn
nhiP8d7cMtoUYsIAUACzmiSjLMyln0Dyp7fAtojRBGBQb3HHz8Jk0YooRR1AMQqV
k65RvbeFQY4n3Nh2BQNcGCirCxzKqiS0ojJUcGXzoKrytrhrSEJRBdyvcxFmThHf
fhdOduc9AkT+WoGuisr9zc2DZ6IscFtoNUYlK1o9zP6hqS3AHMUdggvMOEk/RE7J
WO7LEe/yXsCu1XRARS9CwzISBQWCKVC3kVl3fv2gQQDhUfeJLP8euICX2Gr6btvQ
1NE0RObEQeNC/xcay0YOuwm58IiI+NHXXX18forVLxVYeSSBQoGBPM8oDaKdW6G7
JwtA+v83AbNPqMW+k4DbUf6RRHSrQeK6gW9u2dCGj4O73sUmhLcUC0l4POdcasGd
5BWzCuWATtf86UlaH1B/bpAFqLAvWmIrApv1xKWY7oMNFNSnXufVIP+1ER3r2jJY
WPnCx2yj2j2BA5R/zvuiT7JvFUSW50GOxmYaNFtPpD0j7yHvhYdjVKM8EIm04eZi
tIzBS2lZd3d58XU7kSNl0ASpjV8GmNNNG6/g/MEXmBepe+dWo7c68t/l0B7gM9ge
nlLjTVCJHGJplUTJc7eNk8JdRdT2Jns+cHnncOSsq0aG5PzbIkuiiW84DwS6Uv4i
DrDkQsM344wP7CBrJ5ZZp9jAesH4kw1JsRauXhYrw9lNctMDYAZz//dpt77fb7W+
u6OM845o/V6K0vMjKob1NaCveC9U2ahFMOS/VOagE91KCUn7L0itHMTcaXxf5P9Z
OZ+Y6SW/dCigc7+W8/rxbVX22AgdQ/XsV/tAVEVhTrTJEDd0/4QMGrkqePayjurg
IreRc35oRRNxYDjCp9hAsjtPFsCvJoL7qITzgWIR9n36aqxiSvgdODS+pZJbzp3c
G52Y47XhiTtPDs1w+3uHZVYS4Dy8fmBRo7hbCCJwvIcu6w4GZbDAd12hxMUnZjHf
xuIjMSDcCH5hM1nGiztHOACNL4p2CFk5stIy+zbwyIRakDBGYYb8gZ2pA6V/BGx2
7M0q5je/Y9Xn/1HBLQsjSoolcpgx7J8IzdV+ZVY3f9UibvrNrKCbVKjLO5tHfJne
bARm9Ez7gxsbHQ5fYEC4pHipzGhSk125QJT0FbwqSUFqJ/Bixaw/5zkaUztWfcmh
zg2NQGvCJyv5wm7oWM9BZxrk4Po50snUgjRhF96ey9ruVfRCIkQoCJeR03OoR+xc
tFbXph4QDYjxK2GgcAHUufnxwhbcWQZeKZDMSuyFUAliDleYH5IJxEUMtzLU9Gcm
6KthhFjJ+4LAVb+1w8D3SnwUKKJcLrjrM1MrMcilm5hURnpEmO7/1GBy+cGF/8Ol
erPbrOUdff25vfPaKIFmFhexZD7ul7AkpAGCuCWZbLZKLxOZXUtdEeAnc7fwsywJ
bgi0prGsxKed7vd+BDTYVEOX0wJDfdrZusSPW4/02DeejBcT7LOBBleYZM4jGTUV
GcTs0BhKbIwpg+vOAlK1X/TneLUDPVWqYYYON4dAe9eRzDq9YHvY51n+axObMpby
mzMxGg3LY1MF0KQOYbsbm0Sm926+0cPyOhV4jE5kEy79fwxNc6Nz3ulKAkWBufH+
foi5hocyHZGCdH2UtG0oTHAAbVMQo+IyZWWFxAZe+Vuf8cWq9kLOxDtsO2DYVa6u
2O+LxQmi30ZFDrLUVywXXTGBE+Way+sBWUCT7LlEtEC5RqrDdWO5QcWEipBetLi9
yckrTw8g7MnNkOh+APCww8967IxqA5Obr9S7LLVoyGRl6xnsVoVQQdwRJRpaMCE0
TYY1iXlyH0tr3nPQwH2edAEe638YWV28FrrsKNJMyZG706hNR75TvgA4IBsz5cYf
MBaATzhr8qZnX03BTaOT2sAXeiC9cQ09VYJV/gfxEwTedfS77bca3Yvs/2TaNfCi
DHbvCRI/m7ssUkgNu9aIvSsuDxWJ+RzIp17XOxF3GGsrsQj2byhRZb1O9xz9uG8M
ZQR1BuDl1ZyU8LKQI1X0+PydEzekg0aIBSSG0UR2fQBkBY9ukan3f1zZ/NoHkmJg
dqvg+6dyK7gdDaxL0p/UB4+vqinwyJEfHB2bOVDQMqqr/1uGikUqu7369StO/FgR
gsOIY2o2JKQLc+OYKEkNcmGu3g/rdBRYSlh7+hz0LR3lqD7etzVlDOeePKw3X8Xs
tIP50iif/r82dYmNdUUIt7WDl/L2kBvtWFkQi0nMwetDqGIW6uOV0x5T2JTR1QRS
LX+vRDAZaWeOdQZnc2JRx3VKBPuzgZe19XRYRicuBXCYLJFDbWkXXI3Fz6zgeEVv
6loIo4P0oNiajD0bakHKU77KKLjWui/7Stl77AP3t5G4C3nTRbxkbA/iuzXCFnDA
D87Ndi0A5Gu7cvZlAebUbT5IzUY7akTmOltvec3TyxVS2ON9SNf7FOETAQUyCxk0
WX/wgBQQy/MC2mfRjF/4RbkP07AaZUiLVcMvPrb9aVcHv3ewN27FXV/GP6h+827c
MmXy+TIedozJ8KKOyaa81TQlD+lXB9PHdGdcGYnDLjdrgZmfIPJQXlOOLgaLh06f
LRkh0M1QnQKwLklizqueAmPvzNA1LNpieOheZymsDex01c4yRhSXz5WbW+x6FnGg
oQKgJiAGLMScnHNTOQyvfBsAjiNpuvQjRgHZQyHKt8bBxgoUhq4bob8kk2fgSfD6
wDifq/5lDoPd0pqkIEs+30GpK2E41oCb54SbWzLBwul7qSZ0KgePvZmfPoEXMLSs
oihIr4xO3k77Uo+sZkCGRaQxiRFvccJtjckJbMyklmo1DW16val5SB9CLqtnwR8X
uJ55VlZvRvhzTjdpSOGlB8ZWcanGIwfqKZlVUOz0gjP81/mrmS3QX0Ak26Q1PxQV
dTeOpphc1vBKpBqhX7l1VgPjhEplLLNwwq+5Mkm5NQ2u6D3fb27EG/t1Lu2wMhuf
VBFgsIeQ/QVYyh5dOA8vluDa7iHZQImjni7nV8HBU05zQ4A3cqqrhsRWIEBXZ4fc
z2rp6E/kjs0sXiozpgdrMhP5KOZn+fNXsCxCe+qcAhlPzOkC2YD8jzCnpPiTfWlm
NAxAfCH44Dc3gOEwOTm+R6ukZP6NmnagRgsqBBoMzxcM+pSo0BObP8svzgWySnDq
bKjWcz2D1lalmzOVr5cbrV4+4X1/7QxSHiyq8T+JKi3MUgdR3nmW65E4rs4JG++n
WdeFU7LwOdk0gWEai5AQM3+zn+2aMZ03L5RdbX+xaXIMt2DR1/Ln0xKbifJOMFib
QGMa7uzz7f6/WwQAy3AGrWybKaLgA1nfUijGTLKWPsoUxdUkTAC/lTbfxWpB90et
mqm7CLWSKH2r5li26i8AAfEB0I2mGAu7wTCYoRmSuYWZV2A3RhAzYhoNwKrmCWGE
GKhQePlkzj4YKZOhnCDLB1ubjPyXH43yD6EVGYLFEdfcISnrLscZwJkTQq5YbPNY
79pyv7Osq4P71q3xRwiN5w2hhvmuFmgxYMwBvi585gNcv+S/U/T6yaUJLByTS+mg
L33k50nSluCnwbqX2F6XiWJ1Zvn98qo7aO54GlaY0X/rmpj4kehUlM5w6XFw4p2o
QdQqDm83joMtcQISO1asJFR+MbIOwETqX5SgM4WS/ltElHRHjicyZzxQ27GBGkJO
TyAJajTg3svX1ESQ1hkNFoEx+PM5EpRaBnuoLV88W+/fDN6QWf5Bkge3vJ0iP0sr
IOSI4lXHilch7vTstu6l7zmCrLjgaSRzQhNULCrxAVo9ETdav9f7WvBPT3IednRZ
zpyceVcS7rOi5fs/c9IOGFVKPsrehfR+0TPOPqyCyyN7csupuKvWgQ2BNa1P4YLQ
t0dwEGFTTgdxq+/Uetw4JfCV3XyXfuXOVw5/Xe6O87aoKMcwOgZtuou0+L/ze4Zl
QqS2K23tEp2p8rFOVIXN/lkYgouwMuQjvpSe5TLdN/NJV8d6JAFGElOJ+BsTErjW
kX6B5z2Bi7WwXwDKSfWEc9BFcXT3SmMMWIgl/0b7PPoshj4U8YxiSkVK44NWzFm+
IJLF3/ZkrwH88mGsmuNHxKLfpdMd3RbVMEWDXAasrPcX6UMk7EIoaWtpmgTBFGjR
DH04VR/D/fL+huYLT8tFx2gmspCUJIUDOTPvYTl5lhZBplDQHOF6U4R64LI9If4L
694RaTMms4wem8/AbKng08bjMsvtxoghu33rvicZdPP/zBMxSqEzm66f1IOPRQcb
PufCbGHo+hZyUSPOivdv5D6N3ULfLSCeH1h7HZ4vjLVKfG+coDdFBNGu1atWaiRX
5xp7QN8ffQRxONxksgdIG5pNGi1ZlfFAhl+v1nDdfBfqmk0GluwgOnFSbEXqY7vZ
c7kqHOCg/gkUVvZdhVCIosh7wTyZ789xhZgczHB3TJ7U57jVgb32iTvJTKUr5mKN
3gPieLqG+L0Trv8RbxZnl7ajvrR7Va/+qzamZl/7MfzQGkaE9WJ8wG7TF5+yFJ7e
jlizkeNcaW14NKqUZH/mHuE8sjsuwoZp0j+BwXYXB91+YoUYSG4CmbzSejpvNSDR
YkCNjkF/w9hbQebh/lCLxkNO22wcczKzzXl6FT//WKaNG+PR0o4UGJJkXtIwJZbK
wL2KYD8jYIvksEgw5VIPLxaZs4Lkct7SBCCiD1UZsHjMAyM13hN4WbyakuLtfofn
WgTqxaPej7xs7BhsyiwpMU1a73w/+bGgIf1pd/dOpiUkv23hfFrOqXoMr67tfblY
4RyQHDqORXOXsR9wLUtVCErVGCEVo7rT1yL4/P4jArkQaF72n7AnKu/2MBaieNhw
QSKawRHaofjwGCpIdCh0/sXv408Inkqm5lQZeokbtBF8mOUuNlJxS87SBP1GjvJx
z0QyDdidyMRzV4yFxQ4fTGgFDqXixUHFM2APoU/lfIcrEb63VGlz31gdVxHF9faU
q6SdRC6KyCzkJ3PExfJP7lGqiJPwLlDTfhCGiyCtwPVtWaccQYMdckLsW67qQ4JN
sIMiouyrFTEIo2+Q1TXPXQEcHH25Xe+P86tHla6znHjmdrL3OcXmOx9qAoDIk6iM
z1e0/sz55CanQLdg9yzE8RJe6FJFkVXGuql3lcIKoVQVinNwCLwNRudehuJz3dA+
Y0TY6Pwt/ze9mC2UFvxLJdtmuVQfEWXxPQQHGdcvvhabIQwCx9iHiELXoKE2cPbh
WUauwHuh9N/Uad+ktXpxL1HeE8yNmbZPqmnDMrafxdHpJyImw2mmoESLdWmTFI3F
27/6MUSL8sm6c/BAfsSaz6uKR2qBEjDhdUUYqK3OjK8kS9zX2NC/8zL8OfiIu3V6
rjz9MKfe31sDvXe5yRjIPfUoHpZTWcU+mBoD01de0HwhqlL38nNDzhs7unj4NZrz
T2Rv8DaIqJeZGWSBp8eAY+RCmrUCF5k5AmLLNxyJWrUKrgNUn7UsxA+PIvIls7pC
NS7I6gFv9dk0F/jYryUOobE7DlCuan4ttUDTA6Xv1oKHwoELUDyP4rCryE1V4Gu3
OQhi5E6MUp7Ki9qyxXkC3xlQUczTSrbE992mdTdXacZwhaZZeiI9CYXfwN0XciGM
ReCB3b33cugF6BadY20cFh2o9yW+F7nDU1kNFO2Lcap5Q3H3uf94YTDghvDYLpCy
YONQFz0r2ZdnbmCXXd9IgRp0WrbEJJrKLxGwzY9WwxXe3zuX7XdqnFxtozXF1K4X
Hfy1Ph4GOSCxPRDFEIkROI+gUijbe/ZgzsZ9/fQiXdnWztA1eNIeHrKlLTIUN9BJ
r3zvR1W+gjvGvfjug0jyRZTH1qJGEoM6paYbLktf6se3h7jsSsnxgfX/meACD3Av
DU2Vjm6l+x3K0RXIP6tD8Ae5/8IqEOPfu28hbfObt9J2QgdVsL4aKvNYJFzAnNaX
PUVdqbUkvyPZBmneb0N3w8BCFCWxM8jhvMnDCug8bPlm8YN2MV8/Jzs7RZbR7ACq
Wb/araBh9YaZOn635h9ZOpsDs9BGkx/utKDRNKifpn+2ktCVB7ub8sVrcMOYvtIs
eQB0Ra7GcLOycPV4XebckA9oKwGqzoqu/NU3HGwmTm35owKLWSFQmwvwwbUMErlD
29xr1liDL6pFI9cRhKgFZ21QXYCcNCGLqLy7Rzx9m39O53tIUgQWuOIIE3ZLWkhv
ZEogjASHGFi1zSBLsaDMC4PnP0sI49HXOPcWfU6ypqZYrNMzBsFm6X/M7Z/O6jFz
TC0FXhlxrsu07/bSJFw2gUT8fjnIs50f6fW+itdRM0mpr62Cgwe/FvgTXQYAAhOT
rnAG/fYbkqaJctUPBwhPi4nV58QEESmfQ212EQY0awfYd71D7k+ShlxOzxaLHPQX
HIonlGQnfSbBreYGVxqj3lb9cSNTQWWJLZdBAiP3OHlIXG4VUBNgV9ZrnS2dIbme
UGfK6hNtc6WnHREz988/CAkFNVvQznBALiUv6aSyj9U3kWNF2Uqejl93tec8/pNp
EzBPOa9n9FLBlNYhYL3RRaf0+mdjfcdn3btujkO7pxx5GK2nkXRfGEDWzAPpXXAu
0mPB3sOYzYuDVzNn/ISKWdrn/eT/f0U19zz2s+ZO+3n5IDpWfjo1LNeW4iiMRWLR
pSIBGUyHxzX/AtAb+BC/Csjx7S2an4yNgt9vzxCVBdM4EAF3H8njnhVbkD8AOOB7
tcDL4KI0q8Vi2VGJ7gHNcP4SUgGlb7g3e3BHA5CmY5nhMenoq51SCJewDGRxfXev
XdRjuXL3oEM9i678A0k8mll1Szks9F3eKePys0bT/T0/iS95+yQN4hdKPvxP3yJi
KL2LL//MjZF5uPWt1HG08yoz70vnGj7CJoGTXPFIGeaLwnjZzmaReyp7072mudMQ
l9nTAO0clyxm2LEDOZnyaBrkbcOYMkWRk2kJOiRa3CcAj6zrYBlch6SyoOYGreu0
do79W+cJLtWYBRoURxLteWvrU68HD0sr7DczX7imWB9Jk4bUw578ehP5JIA5qEWJ
ISN+tGfiB4IE3eWwtWpbOY/pLDvOgrlW9PkTA9K0mEvahW+JV+Ot5VJL63leRjLN
UINWE3OevD70NAEexjmn+HgeNW1BEorSOq9C9E+I85vshhyyRh45WBpzOXNIsCcv
XArInjv8DTc1ENO8lXN8rGLfpY+5EJKRKhWx1omdTRN3nzARM0O6S8hop3Y2TOt6
o7BqEAs7PukWmfMQU3dswhSSN89ERgjBSWTSpC4K9B6ik7Uc/ALuIpzAx4haYerQ
KABzdJlR1yPOvh0t1GTk7WtNU9N0i/HdF1sdclLXLskWBiCg58bwrNtpu30OahEl
QLbnKec+x0/KesqWate0DC68uVAcPrVHxXSck1fiv6ubpJKy4OfgJVyaJMt0c+At
SGD4OwfAgXKM716l2mDSqvFLHN68u+VlAmzR88jrG6mvyUaph4vTB0FNQJaeDcqK
TpUb5TcySKe+Zx0kITLls6AIsQuHUtQ+ASgCy/bfesfd1Cf8hB6Sec6nxmAIFTha
OVt0oWxvzqvwhWlSwTSYjyBlhHxDCEM5G2gOmTR4aPAUjmgKl/6K0rf4sr9i6LLO
M3DOJwh4xsnPNl96Ym6cYnhBGZjMMk4Gdj04m4acJyd02MXuetc9pVsHo+JGlLHc
jHPZpJbNVmKgEgxqFbSgSFGYikL6BMdwIZgzOfEOH6Qvx/eJ3upPrrP92ElV4+ih
24vok6ZWe9SuTSZNLkHUJFr/i5jnrI52l7cqdHyRcJKWGLHdWVXB4vo5sbL8er06
0HlUoORSyo0ij6pCZz42k1w3wY19YM8A2AVqPZtpXD+hbo6XLZfvJUjC7GFZZo+X
7JQMz7a9BV7MQIO/iOjF5MMjjjhRleps8LkOmkp7RQXeRmvOFnhJtrkYg/GgvINE
F6Wr85X9mi8bA+XiZg1Q5eC+ins9nC1yI0eOBtOBtp/kuxIh+YiBrR8nOXSgD3ME
PaNBCH1Swh/qtk1NQ/iOP3IEcgpEsfv/q4Gb/2G9HffSKYIwWfwF22mXXVMw4qdK
blnVV/Fppad6TPT5CCdtIn6iII54eEcMuCYsGQIDmwkcSniUFqMUOE1qY1GUZrm5
zLRqk7FimARKHjlEtq5GPxnAcZmm2uYswGxSB2QuR63Mu0qCQGA/hi0vs8sHkkE8
D3m5mPoEP71jNVYP8aWE5/RqIQWkIhmU1FJZbm+ijos0ZrjZLb4fN5QWvi6R9JEv
8voZPLKN2Lvl0yvoHwqC9caltLWmTMmLGTI5xcuJaUU0Q6X4DH8X3EhpNLdA3Vtj
55DFDbmLwji/dUGE2zMpTRPRhnKHnzoqarGicPec9OjFcuwJIBe0uvq4BYW5NVdA
IAyuXRjJWVGGOtu4p0mtt5QRo5Rm9pEu13Wans1EO/uRQkSUORPywyeC/9z0U5H+
KKbJmkbsQy8/3CA42dJtMWtTdo5miHO3K927KCs7m1bw/WRqgjYCOXlcTc3onwDq
oC5k2ztSov26WsYg/QVKBiMXgcs1PrEdSiQMSoPCyTRRoPmXCzWA0XdCLijLKpVA
vVUMejh0MDnr1jS47a+7N5rL8x179BpiFHf6CRHK5o9Ou915EhUu79R4mRVrB+yV
a3xkQutMNQ4qHvTTix4U/xtkqVFXNtvKR8P8LzbRbdk37r0xVaj9OKVoydMcTT/w
SN7nYmrTBpjl/PcAU0W9P47MHzXwv9p5pTPbPhn+pJGxsvvxazoXlMp8Y1KKzIbo
BA69PywrolFwpOUzjxOiJwRaABt/EeqAGp1DN2M2UlxpW+H2RAbbUeJoRpEvMIFy
nYs41AlTg0akEK1fszH75Bl0Jn1pcSRsGJjIYa+o8+4dQVPj0BPQvOBe1LwQsh8x
Iwt8Jp8JWOfhrFZnY323Q14bXvnHJRBUfOsQWy26q5lqCyJ5WIjob3OzkBCMtc4/
RBGnyS+7nGnhCb8ht7EfmjzxaXK4Mr3jjqVSrJeOxTpPqxTeBnez39uFYfMwucMW
4n7bn6aqvLp7xssQj9EkBNN9avxtYolwBDptWzTH59Gg0pikb+Jkmq8HILnnzGJy
dfiPVZ3smhVb+eunHgDcSBky0EBApWPAjr5zeSyugvjFUgtrDU1o5wIIhv6UL8B7
dsmjSiGoXDwTDL980ZOXOXEOvqp7P4ccXrK5y3ugcChY3Cn87lGeMsj/JorTlGUV
ONLrUjrS/8uPEcIU3doLBQeSGiLF+F1e5yiFz7Ju1ROTUii1ANPB5sSVr6bpDa44
BbpQwjYkdEzDS96yPl+oZZmQ6zYwx7Aj1e6UNXOQowNQzNS3TMuFdCtWGvZWOZeS
gSN4HrxSNPm7JNUSl5NcrYtYtwm3Tti7OlTrfjlj0V+fLtJBdClOgnDdOdVP73F6
lOSQeLZLbb02yZ7ji6/aQzH2VC6ViaJoDnS+E7ga81utmy63Z0halYUW4V8bh9fk
MOXvEjaqZN9i3ItfrCFLMJ7bZhmLBjAivMKL9d/oG8+Kl1YhIrApR8TFF7rADHMt
OywzPcNfW99NMtmROC4WkUHIQ+WlrJkI9zn1MfM2jNcjyOzaTXaDAiVNJUi/v83M
PjKoEjPmoLVzfFokupBELe5E7KuVDAh+qZNPFT2BgZOmh1M7voCFfOrCYZ4+4ZAb
fF9e3FBg9ERzX1EDmh2LZqQwE6wAX4FUzk2W3LUKkxu2DQu+2WHtN2x2DXH8OUUk
jYs2F6+2JRdyUTOwNdBWtjuh7j/tsV/yWsYKHIRQeqTL1JmyVZX0Pw1T76NjuF0u
vzcnl3wAd4hqRw9i8j1zsW1qt0rmr5JaVKuRcD16HmhAV9KF6Yxi3bpKC5RfeGlJ
/s/TwGb8AHhnShaF8EGDPhzPakuiISvJ83eM9cKtMHcaTubnWgXE0taZJbcRwUAb
6OlNnf2xWbRmNkn8u2nbWN5D0bSgsHJ31LmnmS5ISGKJUGBR9cHG6InW0MB7Eu4Q
9XyosPPXUQqZg7mBybMSjP+Pkb6WiYEzPyfGZv1vIvZbzFV3rUtFBk2D/od82I96
t6Y0Z2ot9MkieO2vAkSJEspOPiqpK34cBYfTALyrE87BDh9xTGGC2tk23kkkgRUH
ctY1lt+z7oGD1R1/cyhDmRqeC/72UYIcxEA/r9mWeKQzQOAs92gO4bjqyYt0xd8T
cBYdjWqp+5PmZrgV8GfxA5Q3GMB86tNEe9P9fczPuTklR1Ub0yR15Vy1CeToGYZj
mimj5Mjdeou2EGF9rUT9R0a6/EhotEfInHOdIKyb0cTTO9d+mFOlviLgvFo2Llme
Lj1OSnGETOLCKoUgJezND47IjqjPiNwB2xb0JSQdp6VsV6Xz19n4HAaIb0htvdNt
Z+5BgNJ162SLAbZ6pDC8JaGwB4GkBLJpRDtwWIU0C9rDcqZ/Qy7c+DL4h62EzQr1
D5jYu+pBIaB7aSL23EDVm2TE+d0TGtcWC7SAvaacznuYjohtKIgRUbDDoShdBxio
c/a6yjnHXr5Zjkqz+S7bk9nJx/WfZsufpg4I7RweGXxwp6LoSpVcIfJFI+2MNuQ9
ENfFgkI6JmrPE8kaC6t6o7wlhq+SDl+snkZXQ835h58007qfMT46cDvfTsy67dDj
m9zuaP74OS0HOx0EVu6oNlWgflQJxaGubGCjfgvDIdpCxLK1iovjGZWGA2ylifAK
EEEjATpM0nXUxPpYv1zzhUO7vTgawguGlNtUmex7We5Dkxh7MU//hebmKn9h+QdH
LxxSh7gyqrH7vCnwKcU9IjRdDdFNyCF6s5DX84EEV34AETa+osTDFyhz7TNH3rqU
Ptd/n65DW7jAN7QCY+MWJUhEs03pvXLxAgr1g9NDaDYArBhoMgV7xjf7E+tGxE7Q
qM1Brw1QAQyO8Er0zNgGv1FfbnUQRB+EYLqKH00qgV+DLuwG3AKNan93hl/nFEzh
Gofen+k1TqtPLwSQHt6vnSCK3IcYBoEFFD/loNUz5PFK9InGCxXrjcLUkcF+B+Mp
vwyjInCy0T7J4VT9ea3QfGGLYJGx1mX8vAqRHbqInL6V3z1pygjgqE3Dgadqqlyu
SyGJGz/n8+5QNiaHB8mJI1URLzwy4zpWQf0luTteq6fsyRt4AhwCp7abXvq4pQ84
SlAchBvPCcXgYbLQSv7ldbczB+tWeDDT4pm0E35W0DLHVAJd9ZgKLAgcpc25VPWX
+AIHB0bXL3zRLEHPmsQBxyZOc6sgLtCTNNxeZh7TXHJu+wmgJsaB2n/CeIhSENM9
Y2W7Xr2Jzmni/vFapl1Yt+W36puA1uj2Y/8Qq7Yd4GoaQ/5gEgsVIwUEuRm2hncT
hroGLRaIwJF8L2E3LY8i2Bjklnu4CNVEUeWz19dsOIKh7n2K244Y5s28TlGZV0/Z
REP1WN90Pf28jw1Xd9NPKsqYoAcOOwEooTA4BP/R16ajEMY1ku1xkLzJj5I2Ts5l
OiYik6EwIpaanLsT3Y0k3k+ZOwbUYWRy5floysY9Fk3Qm0amiVTBKkJRoZjrhlNo
8Die3MZkwnm+pVhR7jdnNv2+AHTBccdwIPm7bCUtMJ8VnE/9E0RJaI65QD8ZyXxb
iatRMx8OAp4/nr3tb1pElBwQnMmrJC2cW0BfFq3BM/GM3RWp/zjywgORfMnZHVHo
pasO7obU4zIMIwoujn/rEfDqHx95Y97GFtsqPhZVezcxSEigTKdvEKpirxTCbha/
OWp+ZbHmy/8uPDPFCDZOPtpY3QkL4jl1jKZ0A+B01S7/7cxMpT+1h3zshx0ejGXc
xML8xQ8RiihCA8fcjlz/ZQP8edzIGQPKGkdnh4CXzbLkCLXF0AenBZDR/7gO14DE
BLMiuKbYPvc7tsGya3LW/Uf1dXNJhoKPf4ON+9wxaj7Cr7z/oZsgJyXrZOPxyhFh
BU5lnUhCF5YJxVmnxnmGVsmUwtwbwY43/U0+i271Q+umXLrJFucYlnQ7rFU5yIsZ
O6Q+b89SGqiMWpzK4PdoZwk1agNoV1Xs6OyJksierfMcTfKEATkTDeVGzmMlD270
eGKOb8yqdC1kA60mtjjcW0qXebhkiBsdMrTaWCYosQTUfgemsNFAKr7bPySjb8Iz
1B4BwHS/pc/qbfzkL7tM4yMALSDCeWO8mJJcvici4SfpJppfuWuFnMXpg5Rf1Sgj
hnCM//rwlUbZdXIuapip0Z+BmZDkIvsIEJy2auPXzKBa3cvfXH8s95ttQnw49Gsv
doSYgb8Ue+J4fSgRfaB1hp/QPE+wbjQ903LmQ/Tsc+pVo5nTyH/mbuB4sNg2BABC
hQXLHdSiSpS6azsnmoqkdEZQw6/S5dg4l1JnkSrSZwIhQY85X4hRHopB0CRbHrfP
mM0qiDb1I6ZN71+eyNo1uA66dnwyCu+/bxgfZZzc3cmyrctTNPonb43rzUYViYpl
28n909qkEUUIpPoSE4Myb4IB6F73rx/gOtvJaCBB2YL8rrR7zhId8lXr2JqrzNDx
7ntl2HBsRAx4kfMe61QPzkRW8endvvZHoQjJiMSYaAu8CuVnwmrsNGNwagfrpFwg
laN1ztWmfDWq7ihEgCnczWrvS4uN230gW1qrfkQ/a31C8WiWmMv2IZ936aIXTowb
C90MoBaIiP1Q3HTVsy6j61I0amAf5QLKoruGqg7otZ2ysVRVPdtr1aL/TQxXUwlt
8LMqCrcUmwPRJfeJ1mX0AyqtmIIeB5gHeujEHB6X+uCKdFAsM3oLJpl6Gwc0plj7
+7s01ASzJPwkWNCFP4kE01NW8+QwoHizMwTeO6ONA256nl5jw2bo8TDbhqg5qyyb
DNBsp7rBZiv3ILuyCnosnvP1Ge7l0daIrKqcDNGTCZhDe8rxWfKmFg7I2LDCDNG5
Ag7j8Ou4bfvWSwimlm2gE043ivUxoyrkTqXdZCq1SGasERb7eHeQjrqU+OEVRX1g
5xELm7+Su8z0Pl6lj9ZKIDaQsLmmtyMdNo9ml6IR5xWz64r7zOeVvFzd8IjmQFaN
9b3aT2dP+9jk2FTgOitItnH32rfEoEqnRoxODlM0JH2dfFBbGH8ukjkRIuPMaX7J
j1Pw19qBitmIbpBfJBA7rR+gx1VtJJfKBrxkmAVRxGWJV03Lkn6ij0Yc6eP4rHPg
QjeOgLX1Z5B8iSpXDrHcAWjsdMAc0+Ya4Lm7FoW0I4OnQ9noAbQJtbBVD40ax8QM
uh7MdCzaOoGO/1qO5J5RYfY3Rew9dTPG7JwWS4ridXM7uYeF5ESQOOW2V+6tbQit
A17JMi8+X8Cqu19T9k31JLIRyUvaGtuZ9ScZCp+eQBkb3XjpJw9N5ywVlhxw39t1
wFxNAnsegyzXgldFcDY4N0ZLRVvbv5gkPs0Ey7r1hvp31VulvHeF6lsmmkACg8sM
SGqsHyFHun+S1p06uG3SkmUU/eT07tbUKp5vYh3j3hQ89orADrC/LAGT2Vb7j07H
MxWy/t/hCzFU1BSbvL6IUistKmIlZ7LrzzIu1JXwJgIiJ1CsZVoBcfVSNiYm+VJR
ZcUlHZHtCnjokqEQqBDTxV5ASYnj1MrL4eBwe2o1QaM41DHJhFN3dsSlAVdhgw/o
tmZUXKs3DUpYt5zezu/ypXyCPh78jPGTAWO9KX+lEn0kL/OQEw8DU+SlF8dOUtTu
4PQm3+gjdsnUiFcK7AtGMzysYj8LtjytkpfZApGuL03PRPlewmZxfejdPp+df1h/
4N7LyWzMIuzxmB1MBD0vVLjvM1rEHrq74RJYOypLqg5YfiQcFd9wCEgV8M8rjDzI
Uo+EPgcCCLyNY+ixKnyCPhPxytLoyzRLJ1XPiZiAM/0FCAmmjsXgN9snt0t+ctUv
I/kE8NxqqGivqBTJL4TsqM2JEob/orD4K50CFfrnaIOF/gSH1uDGSE/UjHbYIND2
YdDeroWpdld9jlnzP+T/t8LE+MfNpClJwB9dNKUWG59jtkoAqOW3nZufR0Wh3pRL
RV+1UHoTeEGquGEEPOIUCXNIR/VkhmXkb8ap6RhXvY02xjlZZvVYvacto54djpuo
ET05Y3evlXhDyLdLeWrUb49vpgkg5SUZhv51F1bAvr6fxDjRYlcTP8uQx8n9SOMb
bPfIlKytExRRL+nXIL0UwhhQ0b2Rm3+9xMg46es9RrvphXOr0z9XefD3u/xKqVr9
uh93qPYKf7q04bUvxw8YIuPdtVUKhgWXufailGEq2iKhou7KK4nMnhQqy/guyucq
x0L40S/SQRsdAhRxVNkEpaz0/EFM8PhGp7XjBj3QAZFSqHvIcuuXC9B6z3ERRqla
knktkkUHRKnDWVO5Mg27KY+l80lIXjRMcBH1HRjeATzNHHUNpHhy+hgquLWeBQT5
3S/qCQLgh25ZEcbQ15I3B3rQxeay4+PwZW758LDCDBGo1TwwSf1FILtZnDnNrcJb
9JG11Qhn0rDwrGcAS7RFqiNwfTWi6jUTsY+kTqMM4+yiS3E+MpddXHYFHzzKTn5G
xORLsE6p1dJJXocqyMqVVutxeZvEFFwxI+mmYBOhsXnxL0WzCBaDOZuwux4+C5uL
PskedhAo9Eeg6fzptcBSnWFIP7lGG9Zc+sIYv8z/J8GNEDQd71ViwbO6+CmvfmSa
L/zM2x0pgo4idLeNc2Qseg92Z1t1c0NyjYNI8WR7CVk8MkTNT4he7XInqOk7IfZt
NX5JwVR33gMVg2FLf3dsQZSke0hzG1clFPWRITda/GFVJUociJwzjN3Nw+Zo51qs
jBr4+bQjN4CqzbHQdc/2CtAo15wcL6ekOV4bE4Br2Z7DmX0238t4lIymT2i9F20G
BcFNn4i8xvjF0oeFhWEmYINbc+GBFkYltV2UtzKCIcSSSdJZ/he8+ht10FNWQG6f
7BIhxpLLrhT4AdVGJSSWBkN5vN9bzNGVtlYQzCwenrAUCNxLIZP0JG2OJEvaY/mk
WxR/o2HKc+GG2XB77YFl6egt6olahWKqSqDE8tv05ksZ1vrwQVP37Ip+DE7XTBt2
sAPQ4Keooe8jGTBzFwuZdkX7a/wFpKZyUFZlNBpUhTTLr2zXp9hYm4gB2oABYYTk
xb3ppMFUjnKalU4m5nXxSrhrXWpunjgzSQvIO+5PB1hk2Inpo+2u0Nmn0Sq2Dorl
dLGe7LNc28XNzF2/ZB6clbY1yo9eXprVx0Z1zVdLdPioVCIe4dXdHdgrwhh/JNLs
H0q43UPVx0tF8kV7e6fAkgKaxSaGMOGvuSe9R9710fYB7zWJGmsijozXp4Gw3KYO
cc+UAZFV9aICuny14SXciY5eWYdXU0Eiya3XLXHMwN97v0qSn34/P9TI4pnf09nU
/ZoI6sNxL5wnlwT0AafeNTPOusQSX1q5nGp4YAWXetAfR0/k3vQD7sY5xf30riqN
LuQAmeAGuidrcUs+elZPa1TsZuzqz0tB2nYZtwiIM94D3BsEoCT0Oh3/nYFoCJae
sgz3u8uQz7y9ztP+IVtpoEALaNoMyWkhr/DpDFC5mXkNXQZPcKcca4odWbNWFvEC
kNUs/pz9i6JNDfaVd9V65yCuYN+749pyAqYGcnVVo9wuacZD20Ys9dsrDx/xANuC
pRKnMWokf3ECNejual3SuFxQfQv8W5DXX31oKZt0OtQy3RCvxiDKCjDLVAJdAHb2
l+RCojCpXF/qofdOjjXPeYukyAlPlXCvXWD+BbfLnd36LW+dCzBvacKm4uULcXL6
0W4gejH9TmkfWdHKkPNVlFWIPRx4UAFFXCp/9pcTiuN91SnqgkxKSB3/h4WUW5tj
/X49HVev7woS3U7kKcFSyE6IZYSoRYn3d4CEpjjXwPKu5znq8KTxp+kiTqe+VhE1
o7DcZ+9MiV/Av8JqCeo6d7LbhzgREPEAGVNqJa+fwWAJZio7mOTwYpPb/hLxiB4h
34UC5Ou18Yt/Yb7ENP2KL7BtivsJHCfui3UadNxEkfz2TUNDyJXlCI9btzTguhzZ
MQxF7DoBjwujDv6kMvquL+ExMUledS0YPZEfRBkJurSQ6AdgOrYwXBdueOISK0ea
ooKZ/AqeHW/t98iZKDrXOnRprDf18qTx5odg88/ee3LfjfOYvbDKDuOrxJr5Fjk5
nuj74Nq0/o6qB6YIXHk3DolwkZc80Dt17H0alML/7VwXh6wWYz5/bx3iHUncvf+e
BDpKFZM2I7znRjG4q1ykd5QYHmOgrctIQV1BFdSRKHUzPtoPmSb0XMvvN4TeCi4P
EYNY/kggVbxmVeIxpgkMJ5cwVzYXTGxnzTsakpicaLR/JmnOn0EdL5/ddbqHf8EI
g80dpqLgtf6EWNRHARbZ1SRVdcdE+uaubXF4aAbMnZxeyB/usWNwelEfTKIVz2GF
wHQsl0aMxWNruRooj5Qq6G5Wq4V924MQZvizBZaF1SN51iHOMgfOs6hVKhMSc0DQ
3vAGUaVr1WRu0RvbBxgKKzvd4AK11pfehVHwflUQeOj+NiOnsgMUa+wpCjY+ILbI
iQJc0ZevdsDUwCMQyuaixRXsYvGO1QBGWOitOeVSaD1NXnBx58qtJGt7Og9LFCaA
jiypsmlRdkUOMIvQZce8It6s72NNQ8Uo2p1/lJgsv9+HV4Bt3fW1bsvaS7hhF28I
hUsAmFTcUpueD/iF9sg1vQJXtuuMSdfRrJaqmNUJVPNUDfqypWxXjwgs+1IntbkK
Mkd3c6abaVkONo9v4LNOS+y8mEPIyf+RFqq54CaGBbhGzX/Qd6pbBbMSnYiOQR6k
1Ou5snXjMgYHabbrSVHUeFL2kJGxEIG39cXSkriLU3MV3skdiw+2EgR7i2n8DHz+
1MhQ28bqcYCX1kr7EsC7fnjWKlXxOgrQy0t9iQsN7msNnjF7Mjb6Pa+m/W87wjlZ
coXYjdTtLO54G+S0KahmlQ4MsWI0R+3J5vvCkFAYXnU9MG027g2ZJUMoTWC+AOnQ
JIFq8tjMwWUrel+xxqGF0siy9HwEwZWeeMycL6xU+N8CH1TQTwvduNFATpVF8aTJ
MEVkhbPIB5qED+dcgM/iL+4GpeSEHy566KOeIMQPn11er6Ncu14idO+Dpj8ck5oe
GXkvtAWgRnS14zihI+k6Soz3W9waduQRS2ilecPwqhwz3/OMA9CUQ+QsD6pbHnQy
V9vZsfJyJlgQlbsZjzNCsImqvTaavbjyl7MbxJ6jjlOkXVCWdHjcHrVhOu1QT4v2
5WsgnHeQWEN1WbmDufd3Affau1Rbl5qPtpW1alcqutgVEk2h7LsrU2BEicuDWoBw
4qRTINjiLBS1V6sRH2amiay3bt47rhuE41m8pOTkEsqRAZHnFCOH4sHiR2Ph7V0B
qenNr7259eXGw3K50VDh+T+hJn6lw3ktPkHygvWuHYkTSIKXp0+qH0x5czI7BIMx
09ypSQtl6uaCXdrYUY5G5wI4F4I1tY/hu3MU+umSHpXp0p2QwUvS6bdGI2cdgGvQ
iT5iEr5jCR1b6IOck05Ke0RY0ekcfRrqgBBJtLTCWjbCC+9Ehanx8s4Dz/N8ALYp
IYug065P7ootBrzVOApiNi6uYCxKFPIkuMNKBsgdpJIUIGmR93DBJa4xgfnhn7nU
wsUs6vcCfyEuV5CM54aRIja+0D719xolwwPLzv5x5tv6z0O0dR63P1kg81GBPZiE
bl/sA/vYptarBIV6A0d49pdwK2CcpqJzrtW65w5HiOr+12r7xY9YjwrWWuxmjQy5
sl32TzNq02hfKjEazuoqLVF/k5O1+UC5KH4apPymwzLVXk7P6ZqqLq9p64taZsDH
pacBpH3HDMLuwets9lA6p+332vbjvgobedn1MOjVM7BQ9oN3W+SRdh1Gu83HFsTx
Wwl8k82F/mwze8UQ8j+8jE1rL0GWBFeNLZOLvS6ABfFYQXo/uGwDsw1lfm5FG8gW
4RjCu5myzWc7FMqeXSb3dldqrmrp5IWtVV32zHF1MsktOmPSigjpyBi335VceN2l
cGnQ7x371xaYCiWAL6zS5SzIIbMmYEZuAijMNQL/bOxjhHlUd9wVWXXKHbs68U2b
dZdDw9E6nwsL3NtsvmWfe9oeDD6e+DieCAMU5M/BJS2bUlozKD1t3Mz3fk7sRyOi
VSKLdEnwv99zwpGgFyzAhTSmLLIroWCC479DgK4y6WvNLlIhL6s9O3G9p8ySTugz
+FLRncSNPK2tUI1TyFKdDc2R4DN59ZUWZJvlAGVhW8jSiAWX+Lj+G9GIooMBJ6CG
9kFMa33nj7/PAWGWfWpeOA3ddsp8KZPI4uU66kal4a1CTWKbOxrSWKvEqyLusfZ6
FuBG4RaIH+KNBTLUwZXyJFbUU/Df9qm7f8JtIechDGcJy56UAb0EnxVZHT1D8HCw
t2yW+c0JTz+c7aTRxutAiMVujQoe05a921NzeJF1C63I8Ahl21Kl32AfKX3kn/xm
F6d4anqmmWMYm1A0uI8wm/8XcWl5wJPd+5UOVRRQs2t5Qr4pD97o3gL8ElrS80YN
P7UgMpzE9xtjcQj81O1SN+7z+u/1kQWuYHvhe42UVNXBzgElEDliQZbHoOUpVAsT
EFmMpFQwlE/4W0zV1CF//qC3kyQjMwHS/GQfL+qkdSg6LiliYYYskXW0dlX6Qt7v
aalnOUxUaYcshk0+GmdSBvxqq5rXy4UL0Bux1IQ0Q50exWzfjMNptNZb7iTCOGkw
D5ycr9BynCd2j4dZPREGEyRTuxzq7bmYyeyEFO6PlAQ2qsF8Mm0XcXc8r4VTmjNz
jyk5BidVNm7MYuk7L6n1Ig2kMs8VNeL7hoANj62uUFq4lcPtsnCDdC7DLcJwKBaz
fOZEcgbreC1i5szBlumJAYnNkUn7LqWBrcYXYu3h/kdYCus9oF8DnMIZHuT9PJN6
wBXkir+4xb84mlnIYQFrMHPL5hA4Qs0Npr8fmgzQxDPhZlfgDLPUUWee3PMuXud9
WnIc/5yPqg2ymudU2aET+8G53XAHEo5XYXklPgaTFvtYD1ewOE9YJQpDibEQJsFd
vGEL1HiKTdLmc+Tdy0Gs3Wl4btMEgBgG/o2LONWpWXSFVzHhjO2Syp0UiQaBL5lt
19W+9VlXFcZZzhtLzE3tJXhiSQ32R+ynabeC5L4HZwh6jPq1IDww3+PwxKGVRLo2
+fCSM49PrvC83J4RNxPjMXtJQ8DlIdodRsZc0+XirvrX15dGKKTFl721zs94eFJx
CyemwKqVBEhtgzm7CUWHe6lcORB8shwQbaMCc09BMkWbcyxVLJq+qYTwTxiiojZL
SFKpurM95Xd8Wmrib3jJTccZzv+uQQhosSCuxwytisWPrwZ+xBsJqCC7t3J06ECA
Q+qO8v8xFQKPAJ5ZhIhQWCUPaUIaZCYgLqgJ4LSQUEeKENqWRqm2eDKgY+GCWtH1
5CxtdSfaG2ickH11coxF2uxFZzeKBJNql9oK867f6B4sizcGR30+Cs2qUDRlW52L
qw+zVUoNe7NYhBys4MGdskh6vw8JTCTH8ddQtynkKOabDxy0vNx4AX1FBj0s7sHV
RqTHpKSGvnipGHO0pxttLfIPq0y6R29xTCZIdihHeWiTu5mBWDuyTeC3uD+fMa7H
PkRructVE84/pVjhRg11KvdILgdEHDl6KxfZAL3l/1GIzoxaggmd7BWOqnzoUct5
Wnu9odY6742YJa2tgcuZWEsSUGU9qEFmUkNpRRGOOW6dNiTg3nq7fSmbCCEjqGva
3WYKY2znnwp/2oXKSRM6umODUnqPv1eDGt5o3muE4kL0P691/n3HBq+uhjnT26iQ
rnzPWgJhX7kq1t/eas0gVyXbhtPcxSyVSPqvb0Xl8r/wlfmtRL5FWlSOhmOFxIAQ
rYFNAviGMiQ4Kz+a1oI9aqef96R1SN+C7e3ZjnzctlFWQEvjAgc0BO67Tb1k3Odb
w+85sErMR/rWVFM4b7l9Lc8K7zCOkKGwrZ03BvnQw8MYi0FDDNrsPy/JPMhGRbxh
G0lDUwK/IZxZRhxZcSbL8be0gicbo3NkyeFxdJi+HRSLY9iUBN4g+FNC8JUvL8Ms
DLMQHDRdKbVKOh4nySmbzgVVRIZmmk/8UCmoqQeFhxT4kiQEUYzmg3oXz8jT1TTp
4XzEYC7qrbGFNtqt5XP+T8F/JGIoKWoXzroPUQ5rCwb649XViM9SVpRw2damuG18
oAaI3Y9KrDHTvOKxaRaX1Use8Z9HVlswnmrj7iIGxbCQcmP9CRBZGcMbpKYWZJYa
/bxBRANan5SrjyfGo3QU6DKiA+YMelNpSiDqsYNqITCsFbbzU9qmgwvLsMbE9wzo
E9kDnDU7+aQnPizji218KLfjQ1zmS3Qs8rhihPuf6kWQc19uS0xq9PHSGQXLZ/9z
xsZs0sg8T3RH5+4Pv/DcI4smUwNpT67u9yir3vfmYZkhBAQaKYDNUmpkG9RtWOm0
TUG2uzyIFt8T+e57K/Gc1xyNUrXVImkrlJ8KIDWyL95xQ8Z3ACW7sszKDqsB1Xoj
UJDNd1ANlFBtwD3K9v3yXV0r5mOOPWQz6Q4TrpK8nfZY+Cc2qSnYweGKRbuCUETo
qnZfZzlevaYUalNm4j6619EfXC0UXAzwb2Xh+Cn2FJ1j2C7HxkfJjeWiZkC5iY8u
0KUIKjanK4dVaP6EQZnIi/7Lfn6HLhqtLHw+UvwTr8l1xPjly0KSBzwfxH4OlFEt
JjhiWlkUw9GhUMBgUX8f9a14eZaLBl529ZsoasqC4W2nl3z3taX54pnEF3Iwus0v
9X6ztR2HsKOtBG8AyR9L+L14truQiTKXFOP9cMMAK1D32MsueHTaYRHm46pDX9zd
BpYIJgJ9+VvUx00e3uJrM7Uqyo9xDrW5YdgNRjDYJB+DXwyweL2OmgQ3niX1Z1F5
uapwQ93OLIqlJbfiPWpa2piVkHl8MWBEA5o3SXr3Z6kDZ4x1eQCwqhoGS1KatQv7
cDDXLgzl6iTpjIKj3wmt8B+1s93U0z1J5V1EsuRs8n6t5gETw8G/6GiqJIHv+cAC
5zxpzJMVZ6YAw4UtyBPncZpOKzgz0cK2jtVnUFDFI/Zlvpf+9SaLmwhHqAaIve0E
/KERA/68ClwUFSH5bLOYg06TJaBz3KC+PVJ8Ysj6nlrCBQcsIgmS0DyAV5OJKvcr
qE9ZD3SUtGt0lY2Jj3bxBU0/qZ9JZ5sWkf1BtLW3zcKRx/XP34c+pNvXd+/AmH7U
ChQwCxQ/rETp9NN6HgnKLDFMmpE3yZdDJ9nUezmpc/IoyjV2OyLqwDKIEXnOlL1O
dBqMC8VuYNkNBxmtfivQ5qvwJS9rfV5VToOZm8UO+poI7JYT3VrfLMenHugde1Mx
8HcZP8qV+KhqdMphIyqnr+KLiSSSazv0/y5oE9CKWRzUGWl2hOmiZv1ElI0sjsEj
13adh9B+T+g507I2myHvTng2b1FFqTjPgxOxjllRz7St3pSRAJ1Llgj6jeovVZpM
TlYhnwWsejKQRlFpjH+F2Z93Q3KZCrwa6nnqTqXWQCdvoqHfcDRYIRzTWwtV/uJt
O9Ah8WxF2rofVY+dNZzTiiJiK4m27r/+RscNCnzPRwfGm6p07DuNS1lXN5htbdgl
Fnm0GLDgvNWO6t+RcXRvh4kA0HKsHF6U3wjrhFkIzcuUPsJla1zZ9ZDCdoC9WHsz
LBbU+4YpqGuMWHRlUdn1gnKWMZcPrL1C8WtTiJqneyx8AEey4+v/y1o6+hU229o1
nWtKQlyeRWyLwjaUSPWVdbk0HcQAL4lT8rLVwvTzsOXCXnvjwofsxZhCexgCR8ts
1YlEdwRgod/nsB/PPV1lTvmFP+8THbOnp59Ud/aaDPXkG7k56N28X2pBQFVbMaZU
XlOgYD54nvx1AQ95w6y+P9E43wkZJOgjz4DbdIpKexj4SyTmijJBtzROwvYHuQpk
tN5uF2zQNWRTlxsCdKYbt+YgpBPURCurjFW4uxNwUop1ZSYcqzvul4mkiqhNZI2I
UHr6KGcA/+W7zQJxZWQGOpUeQv3lOy7Ity6D/aLeqHEs6QXCdLsZjR0e3ATrZq/q
0fIULGhFH41ooEv57UlNQp32+n1rFLMpRksfJ38UHrjhCNEBycrUFl64FKra7tbl
MAOokyqV5w9NCxc+WWJb9nKoD1PlQuZCytY+2FuG/J1i6EWzCs2nIvvbGR2BZQ3Z
vfRIEC7jhVDfv5IOMXLo4nr85ZjTh11PREwPkJAfZxbFR1OuMrV1jvYCcguUYCZz
a2zKUIwbA7DCUlwhrPoQS+9zovZUdbKveNB80HpCc1jnk3qMf3C2km7IuJcLgdqy
TEF0Dr1UbM/HqSPtcOfSNmuCaVXzlAXJKWzkOuOUAPBlKpphz70/LogQsIXwau1f
j6TKtxjBRPAN7r1F2SPx406Cr+v8PStPwUMSTWfp3cn5VkjZAoEURMhqNwMH8d5t
ZpJdSnAIvzXAT2hDCpuCxVh+W1YkNrIbnBJDMvINe+jkhxjXp//ca0po6Sg4jC4N
/C68uws0NVXCfn7Eziqv0hRr90KAfM51Uu3od9Pg5v00RnX9WIIAhV79wVQx1nDR
PI+HDqLD6Q/FYfxIb2sPvWDHpvR/mi9bZ/u9nWDvE3Y0kF8ZQPQ475CBBJ8MKKYP
sRcIzO2b40aO1PQdz2YjUZUmjIr/86XBxCzxc2HG+kDrq8TnPdGyfX6+1N0but/v
pTHvU5sJkO+APPPzJhdoWSXy/B9V23rhfdpYULctogmWpuDC1FUp++6ueybcYwTu
R8w1fXPvrnX+ZpElwjWKECMFfxvUSSugTwbgsuy7+PppolXbsChxvKf8Mvy/3lGL
cUFtu9+Trcc/h7EhEMhwR3L7eaZJ/g3xuOTxDJ/6ijHjC9x6C2oUNZaFR2tJNcoE
Ewugvhxcp9eNuxY+BICnPOXQpNRBToVQ1Y2jGFLrU+ylj/HqNk0JbwrK5oZR6Plc
4ch5TX0zCdcIgd+PPlp0skQfSbbjqBKCid+LjtdA7k0Qn6kNqZlRZEuscpGMuRPk
nE72hxCVHVMHvLqHkQLLs/7n7anu8hUO/Yop1Vr1oEby/VP9efnhsKRbvhN5NkFb
XBdGr0Je06HNhtWBBz9ZL1+84B7n1e73xZXtkFwlxdiC5eQMlpwE9ZMIFzjMFVpp
YMbik9DBlK+tn//35E6id/SBJ6Y2kFLYdkWaHzT25ha7/v16YMEBR5y/ecst/DqO
xkbQsbbzgI1aKsAe6FuDkHLaiFMgueQEf/W5CVOd12PUOnSkeb3ubVLxWX5rooBx
x3+WhLCmtpArwj4dvkQ1N6p38f+W/nmRd0T8Jdc7EPvC20bsQeDnh/TqJV2V5p5E
mGOyDfFi486wSDlZVUOMfOX/CZC7fRjE2P977e2FiEeENWESEdWjXV2itsbVU1fG
AmaiMMxRI4Sj+R5Wo7z+b2JXdjiFyX5uzl8zDloVPzKBmJq5W7y+CBDcCf4drnzc
/AL2bPNS/vp1o0mxVPYzbx//ICGeYrpJGRg6NDVTjpcINZpzyfIFwU2tq9xS8wC3
gEW734lZRb20lAC5eFc7uIoNrlHTH9fygY/Pd7KXBYOnhsLfp6+bt0S9ZUHb0925
fu1FQr4+wWPgD2PXslG6Pk9eoh/RdHdOpepcHFWQFT+xECDAv0bFFK0fVrEr1tKJ
+jwkvTSSUTt5Sk4lU4EKV163J/8kjlb7wXYSB2DDDe2nO4OC8iz8cX3Mv/wrP9rA
n3DLRBxa4hCQ/z591XgTuqLpSy9JqTyw07Usfb/0kQCuXebJGLkUBfbQpw170dwP
twFCy0Uo2BMzClH6VXBAxfYXrV/MIiLDR6APmolKZG+oziMOD6Qeu1A9EFHiXCV0
RAlyvL5lk3kfFwgxiKm0ApM7nsRnRSqE5S3gkd61r1xyfdCmMg9SD1IeuxgryNSw
n8CE8hHAMhL+q/nx55nfMRI6FEghpqqiqrt0CVzyjDqK7shuZWqyKw6mi1GpyeIM
BbcQoXF+jCCKaiMI+UuFFYecOQ8srt7jNpvedsaoNYJjVaZ6GHoTFEd9gHd0hZSZ
NZ0s4TIG4xW/uQr0++8rF7ZI8dbVJ+PSPnkaIt6vB4bw2BJoNEsgcDEQOlPN+PRZ
x/vba+pDuFnyYDv4moZc3vQAT8eNQRAqBvyiQYI8HF8w1+Ky95HpvDH2tg1Ebprn
nlMq/28aBiCjXH44+gYWSi7/uhzjlRSOcX67ee1AY+bgk89hGNi0kn4ZDTI50vmW
w8EsJa0sDlaSPfmRm52mD4F9QGZ4kBUM1JIBxGOj4I8RoySC3RvNrwUT2pElN4G1
oXTP1P121bsJXB7CNORaBpSfJ1mk3U99mlkPALmfaUFEuS7Vz0Xvi/t//xAsTKe5
sRXo5I4gRmla+TEo5uP/n9bGwhfk7ACdstuPJEymWbqH7pt34IVlvJECUzknWSIi
PeMgrnOcECFwBNiIrUT4pfH22+P3tOHhSvuDMrLdp4H/u7N4w5v4jUHTX+wikOzL
vkT2WrFX9M0CcD9gIBjYfGcv7qxWZbzq0mmm+Iwx5SUqISbPdDZLfrpNW5e09Otk
tbf5QRSIAjZ4F4Cu8LUdKR2lbbt5akZZlQrUvEU2jFv3a2FEzDQBO0OCX/Egfr9G
DaplgOlg9Zf+j5f03Oy3s9U/A/9YsYVVYQHSF5NmO6PuSqCNkeDyn5qEThvwLirQ
jycnkHsTsK20mBEjrCDMR6BAowRMX0+Hrw7DbAWcJ03U6FdkcEGC3H0UwvOtweBd
91Ut+Ef+So5j/Cuea/c9nABDGFH4QDY34NCohGvSFCzYMYy2kLzlRsREgAu9vQPM
jUSJ8KxA7Ha/162Czkfm9ZN8efN4lNI8VXEakX/ZFZLTUWQQzZdlZEzeEK8rOn6W
yY1JHroOA7fF+HfrKMDGYenc0mBMJuby1oXuOlDwMpQxq/ZqaBrtXk6JY50xtDrQ
ug+31/CVaDuYShhnD6Z6nzoKcYU4S7wb95jjn3B+POBhxfvMdcwEBHNzKbkAFMcA
P/ysLExbsPi6qvT+4k/Wo1f9rBYEVrjKI12ZyAAd7yJAB+6u9V7R1awt7QjhHTXw
jXdbE9kJw0u8mkLTLIM0+pQN/ZOv63iuqvybNSWo8tAq0reh+0wPUDJZVIOyn6j5
lX0chDP4WWMAxi8orNLfyh/z3MGEE7giJuyLxz2AQvODXZLaoi4WXZADURDgm5HJ
yBZA55iPGiPQTSNGviPeNwOF5c977LvOSgaWqXvXbTwLRLX5mTxK+BGMS6DZ/XMD
uxzZ75ZvOR6mJiUktpb+DZs9OoaVUd6msGzJw1h1lNjc2m+nOmfuKBZXPESsrUQN
vKq3mrcPSBfIUivfsclUHSoe8KHFhPM+pXOeQvMj1NO0VllmYsLHCu7OXf1izEbQ
wc4OP8PC5gUftFZOHsc7Xg1JwuWlOr2W6i52XtzrnpPm/1cqyFh91ejSOSeSvLdh
MgXlTux0VIn8IFo8DtQbhX/FcrbIaDPaqZ4vKeFB9c9C2NcsZ58eKAhdasujE7Tk
VjtoR+qQS+VpAHo9oU2DzuN978jmAQMEGOesc7CZgE3EUPZCFbM2ig1stxAFu8Td
qHx3bQ/71amHlNOuhBrTkK+Bfc9q3IVOaxz7mHWG02ExBtZQTUEXl+vf3SajRooC
8cMwPGpTMU2w+vI9XtlIT+GflCfGy3WmFXJ9ffna82yAmizwl2VFcok+Gy8ubUJ5
Vvg5k1szQZNI/f7V65SkHGInMms0pK8XyWXdvWYLWAwu5WA0B4VDk+/NuPUjhnBv
OZSL7KFnfJ73PHZdKt09DVvc+YPSpZXErdMFnHDOkViFnCN5yQutpQOGrkKlEZos
WF5nFNQbebQ3T6wFaGcvyg4Q1kBsMji2DnNOzsZMdIyIRhlOl0U1+/yaaWQ+RJEm
M06laiBmXeZJzSMkk0dYv/b9t8YCiA8txgke1w/tyx5LunSkeGas5CM0Pr0Qlh7n
Ogd1yDeC65d/MNQ2tdtsM5r5KKGW+BzPN5JA0rwZPQfF35nB5vg+sRMEyP8Iu/uh
DaGiImaBikInmQNXvV7JFlAxB5sIvvF/fdv7joJmv5LlF53t+PWCGgE9Aww5FQwd
gXsFxjTAQS0tQCabt0OA1RMLKKJVKpWV7cTKift35pJLLiG9cpuJ2HQPO9efqATV
9HoV7i12a5GzJChQeta+vVl5ITDakAMYJZEsfqy3tiJntNJ0+N9K0RYSjBR5sp6t
Pqwr1I/7g33M/WBCDiZLAK8gy1B2xre7r+K2+fJOxwkg6yXvMGpU/D6/v85fKNKz
tPbMUW9XU8cAqraD3TulnIQDGCkyqr1l+k2nz9ofAxDtL0H0ub7Rf9HWJe1WstCu
pyam1Vi+/V4l9SO+yHLHUc7CBG5oaKPmWW6zCfhAWNLO8Aw+LlK+g8vkaHv5QgxB
L9Cz2rtU0le4ekfDZv36Va9TrFzt4u7dbsgCunfG7kI2KxqbX3DM09qXTireuZwq
U47AlSYhriUDQo8Xk/VTDs/aRjcKa4jzWZFClkmB1/uq5AHMXxQoNC+xxfuyH4zI
W2/mJ9Ta/LwbjkPC+247LYjR9PhVyEPrqp/0ohY0mV/tEh+wZPELVrBIv9+wJp7e
Noh6bv5wkozR7+aeI2SVPGwU+SuP1m8ot4KwbK6Rpn+DOL7DdDmwK/6mnrBDOtMh
KSv7zv7Zek/R2glpgV/VM8ilszxsHYXsElNvuvacMoZ44NSG6Bu7Z122QL1VIDVe
Ms+9GhtFqVEFayWqaYMfRCJaQH7J8l/vY9jLl77PsyeqmmUiJyeR8/fSaUhLRAfT
xxM2NXHSt4wAdoVlLOM7SruETrtULRwaj1rLzEhqm+VL44ez/AHjnTWlOXqYXqm0
54sS0DgyJlpf0F5Cci0MN9pnHHizCMwAHACUBBv3g1o1R36wKmIYceF4nG0KBUDg
R8LosELOI/zYeie5FWL6DGc5sVez0xkuy5huk5lCTQeHo4rF0OEzgtNibNr2bb8g
UrzST6I6mUHUDF9RmG725ZpBp2kSfq3P2eGlD/yOTB6UF6G0l9ok+4HgsiQ0U5CL
BV3EWXEhbrJ4v7yXvnqEjwHMRiYZaMBBHH13H4QTce2rHRlh0D6GI1Zz427lGgKd
FEDq37gRE0p7OO095hqH1zqjUBn5hT3OntdnGNBnuY9fITBjNWoXmHvxF5mLz9P1
iVKEI6K2Wn42N90B5Yr6AMfr/c2WgcpotY6PZS7r+q2VZupfbU0KEHw1UlVtjk6k
hh8W9g+hrN2ynt24Ka8CE6a4xPHll730/au2vMphIUvL5hxJPSia1dZ1ZMN5Ltp6
BovwS71BlMAUUacPzU+R/7oFhxNqynikI6d8JQuevOuIQ9+Qd6DOq8frtgxOYsKt
mAleZY9PlU8HqRGhTv4SsqY9n2Eo0u5QhEvaOWS70JgGiy/qXS2zGrszQ9P5Kx5g
NPV6LGWmOF6bCA34xTBYgslewMadwW7M32EEAkh6bN/8PF5s6gUREw/D+aqFoB78
HD8dMXdYJBjINHvyPOrdrhwm3i0wzxyGQoLwDo3VqbsEDF/WjCkubihlRIdOE5yX
e3T3WF1dnfmU34rXttvC+A6v6tfnF6HfqxP5r8Zd7o9DNgJEHJbdJS2I5btSzvfQ
ysfSEmKiBDGnuB1Q4LOgWXlOzzdJc48dYi9UlsYuvsAoOVJBtt3qTYLxkg1f2psK
J10uecEup4GVJpRjvB3EUPz0DH6/IV0HDoIcloKR3txS2Vdx0YlUPNzOMQaL6Zkb
UUQMXH98zBLRl3s78plMVpM5BbXhaaU8RRH/TJRdcdWITDNzNwKrzaqE3rIxsI5l
WT8U7dW4CADcRBMatDD31ty5W+2lWBDiilOkCKbRbAscl8IELPdtjjOs66MAXx9H
igNJJI2xcmywMOXPHCnJBBuZdqKM+3tlzX6vcfOR9SUOY2ODyew8gmxz4Axjp5V1
0YTGWxPLI07FJiail7l+actFlT9t64MIrv6abOHqKFTMdXi9y3RYaN5GlPri3tlX
EmxW2kTcP5lRcx+ztV122WyojA6ssI9knG+qkgg7sMdN7IIQe99txTHk7GkbDEEg
WdMITLkZEfh45Jkrzp9buI9jDHoeIDzzPjLoH9Z4k2YEli4g8Hvdhei4SBmhBVBa
aqm22nqsTSX9QQRKDCFldF73HNbIH8qwn1xdzEXfytCiiueJvC9ak2WtahhYLqN6
JfRwQkn+Dyd0zb1nFc+2p3DvuUATGSF7Gms+Qcb3BW2kn1kifjL8e8DkEyWezr8a
MocL7R5dXBj5qDvlpzf1qVCngL16/DQQOFfMc6LzAqmnUywUgxBslppplZ78TZx+
F1P3SsP/K02j8396Z123R8gw+pOsKFQpHaoG9+Y5Nxj3pbGmJqCGTLycnzyVeSRZ
Cy/gRPhQo3XauhQldtlpsfWoWl5GDfPNxCDp+BZhuFgFHcZuXDTHHz7cNteAMiAI
JXmWB+sHKXNFV9qeKZ3QeGRXjd3MXo/nFlmvQ8pcDEv/aczINVI7A5M0ndAfbg6e
xAUka/qv/QlCGtZo7tvFFuhh58AOxI/Z6kjYRniHYB2qRLpMmruq/zAo3Epa0Z99
efLo1KoWpbVR7jAvTy1KY9w0jTZuGvYbi5m6IF0l8NBUKmcE74UdP05neDC06yX+
qMinatsZKWrPNxaN/6pS+18CLfJLDaDdVo9yAamvE89U6L5c/NfjQnJuYvzahxNv
7YMFJ9hkb2AG5bKELly9LULMiCLDKJ47fTjqxBEMWuOjqky88iTGEwNExtd+ay4+
HgVCQZhOoqfW8ypeHYyQm/QOtX/xnWJY/630ttLN5IPM8zWk20JaHbPBNAILjDcr
zG9XXFLmlcJm5L/iiY4Gzi0YYGAjVfqyQEZJKLBJNsH+MqmefbSjTIEArZvcXYY+
BlPcY6PiUrxLaLR20Lu+vUnjZnjB+7VjC8dYXi41lvl43zD7fMLZQGFNCJnSY4aG
vuhDw2RsHkaqbJ2QEuet+fXAxZ3zK8qhaHH3SGK2UsPGA/eB+zLjzEl6Xr9oicxc
nngNByGN6WJS2fGYq7VicMn4+7aAiuBz8TeOnHVbUnAFO1uqOJl97daE/nHPZkfc
UHZStl3EXHD7RzrkWdhHfVcJTRtU1UbsSWZZRPSG59XHERFVe+bZOqfRbH+cp9Sf
2Inkcdx3qPHBicjSjoKf5xEzv686Yo2kHQOKQGqnAJKaNsOaHtbe8064QyJILib1
LWxLYiZn6RHMNUWmzb64PYJnFCahWYWMdcwf9RCfziUyXfZhfxhNhkXeaR1WPYPr
+4L7+KT/VbPn7GGDl61ICJX6MavHybOwWf7OM0JHQOQyzgFTA+O+VJRIakgP4BfB
WtAG5Y4VhJ4PVSPGNSA+cu1o/jPbIYisuAwlPQcP8RFfUt7c057JTkBEa5IJ3nBL
izRrenRPH3Dnh8URSh0HR6KpLu2B/og1ZqvjXtAnspDLZ8RLQ9Mrpqkw1n+9DMPZ
/WyudbqMGi6gEKYKrkOSommn5Q8GqYmlkafTrnb3NTC6P8AGUtEU65GtMWE/5sA9
B4Ake1HgjIbTo6vTKl+X7EYKwimt1pjx+diYuZXTNubJW0H3PAZLDPdCDZc/s9WV
Lv3n4gnq0Si/NTAD9585EJKX396viOpNT1CNmET3MCHUw1/a54Tlmy5OnfiTNwDt
FISwVGbSuOKEpuTP/9agmJCRxl03yMKHJyReHM9m5PNIkFa6iuBNVaRwLBzG+ZPE
ddRJs7rg096BgGbIeu/48q+j2TR5Zu54b7EBH/j6ziK8TjmiKgmqx7WIW4ePBubx
vLLnGKd7zagiyIAvpEijUirFBHsL4DGrxVRnKmWWeCNiI9Nr0d4ULjnSjxBZPo/A
9VyfuVxt06fonoTmxhqXZ3lko8TFYjNp8EyJgUZB5pkpz5oFSjmLWuWWvK+ayT8P
+VSe0essE4Tp57ovtLvpBqBqz5TXlghWb2NlCGx/4p/4Nk3980pdQh6RPecPrf1Y
yy4q9k0hdwNwd0iqtVh+oBEK1cxbT05gMhfR0iN8oZlxrAmmYYUBIpqkfd6cepDs
rMTxmlLUNd20mD/a4B3AsAGeEgyexyYSBS10BM97i6kzdHFml5gfbjAezelBjOKC
4cUFZ3DwUjTAyXPwz1Gw3OKRPAWvlLdG4WvTseDKpP5H+sgJjC//4pjkAvYRJRe5
8NzIEPxfploh1Y9IqRlObv4BB4FTZ4ZmIj+1b1k/9aUlXC+C2rA6Q3nW+sYRRuQC
3fYSlIWTRB7oeeasW4TAth/i57mVjqYmYduJIAvt6gDnahnGUwh+DliMXfY0Z/vi
1/Q0NOw7jVHguta0uxpjNb1tZnc/atDQX9mx7jcf3EcLi881I2hPMle8oh8fnu/7
m+yE+CkJhlH8OS+wYDVtCYfkhhxKCmTQpxUs5omXQ1zwjw0Z3ZsnQdodsSxdvXxY
pqhdJCaegJiCdIyW7IFCMocGIXFU6VTlve4j4x7dMQOedAUqSCrxVGHXNqQ4u9Wz
TevuftwI7Irca8b2Bz8YXCHqY7Hdho1U9MGEiMUQWN/Mo6caFZzySempr9ETFB8a
n4pLhPgM834KjuD6aVq07joXej6aNToLx0h9d0HBzOJ8OkioD14GqyVRclcXTtt8
55xYWOjBoYjkA5KWt3bb7z5xmNZLZKBx2tKUIlqh8ZtYAX95Ocex0ltu7gxErofb
mpm4H3cvXL/1pozTWb6CxXFmNTAYX4TKhGFunBgutRNr4QQDGZsm8Anv6V7MGWgT
AqjU5RLtBnpTSDCl7e/lSqwTeYo04G3LDqXuoAviJq7xU4vLIMsjh9/s0NKfj7Lk
PBFi3SE14FlRsoKZhQLLRMeM3D/QM97yAzgQ8x2axLxZxHmul/UAUrJZaFydfQPS
+M3Ut67qKid2No6sgR+zwiuSq9Ny2Clz+P0/hXJCOacrC3UekiCcQIq5zKLLjsN7
KmHOp4l6we+Fr0oA+CxmyiBvZRmlAsF3ecuTf1V9uh23sHzSzlF5Dxos2IRdhV+1
QUKhLUUBhRtXHIbEAc/6m4yEscAIohAWlS5GGBBewkuswgyDFiu2C+zJByYuCDbE
2yJYxqTy1xtFN8dUq5IXTQA1t9T+zaaWEprZ47Rrz2InDRj3F525HiFjqu+G/MVb
gEi7POUaGwbO4Q+JhfC4s0JTQbI0y80KwjZ2LwUZ4LyAA3orwyNwGqeliDKInjkn
QqOA8AblC9wrfQ1dZ6RT6qJwicqFAFEK3MSnI9l9yfie7jaNcYW7S8Q539kQNMaK
4MLDl1oYKgq0Ai4I0xfigdLe9Ykh+LPZ2I5YKvML3xVPgW4SqSq9xl2F1BLe0x6X
DK8EmX5Y/aOj87fWN8/9p8VW/T0Mo6udLeXDykFBVOT4LsTTj1pCjM2b08c9WG+I
gHQ0nR6jlZx8cLgOa5J+jvZZrvwtfwVPz9kxYlkkKUJgDBYs43g7EU/bYFxD1h1x
L0R0/LIM3E2RfYk88cDtnS06AaTQ61wJ3SjivT6UNetCbAuDjUEER6sC6g2qpYiw
GBqlutuHH5H9/mnEDmZQiuBsW/OV5cwEZQhUPU5h019ucl2+2m7SD69tuylEb+9K
TrWuNdn/rPgsh0Sf0UojcVofvjgRY8OaXBN1bzF2MagdGg9sYGPuyw+ezCzKfP2x
BUyp6FRkksTZJDcbJiwmceAUn9eWAqMGZPa711DX6OsoWKbfuazVxxBOlapwpAdU
bRhe3bfu6vedLM35i8AogWM1fkD/6M9oCcP7ePTXNcmlpL5KUD4DwI2iAeiYpTOe
ulxsvWbPIueqluBODmPvTHkXwiHKGfQLb1L08GaRYe1ExvtqXhr5lxuy9H6VRxhg
0u9qfl9+rI6qfQwRncMJ/AdmE34KiXaE2GincU4iEG97Nra7xftLTmakbvnYZ/Zi
BHy9FmuxSFO+k9DRzYxG2bgVVUFm4sMEZe9baUIsMLAHsVbKZ1xaLdYVF90oXTPf
ckuQZ3TY0IccxowWf7YlC3M3YpLL2mptrffRhPkkPWPbXydgf6JfPqVMsbO5pyyN
fXgvXM3oPg5Dfb9xk+lcA1JK8U98Q5rY0ILhNzU64Ex45v8XgQrjj2r3IAZEvFWf
As/KAPXhN1bXjPEx1Zh30KirCTtwleGDO2ZoH0i/lPWXaiwMZY2P2FpRrynQtkGl
Z4YJsr5f7z289Z/a9O614rZsae8OjihuO28F4VRqpRFI82HxYIvPVhV7Oq1vAYrl
qoZVtNsJHztBLkfhBAJSrQdZKxIEdGvTzQ61zeq2k87bNUI3OCq2t+TnRu9qy3c6
uYYzFIyCqXYguRNdHMrqxxsTCjoxFjbeaBCUFGuK/FFOs7tLrJdFf0aGTlMY6BDf
0/yC/wjEkDE79cWHuZ/nqJcP3CGFOQqhRgaJZUVXx8XbkTwFM0IoGzPRcy+c90EH
Gyd30VITUJRVDfJA7nfT9W+JC0QbyY3+SAFZYmjj4rGuoxiQIt5vEBGAfyukBXUL
9O4PNNVHp/3ClUD+PLZ3t9B4Lgfdw35ND0lDs7EgDHOAYkpYEPHs+TPLejag0e1u
GHcMiGVnNFmQU7tcoANnkP6sgJzxKzNcgmzPf1y0+1TnIlSo6vGv/N8DgjgDvaxs
Zu25m9FaFHIIIPlfMZZdeS2z0PHgSavq+QZ3FpDxl+4b5wI2ihYHN6fEj5n3OsAi
sDvCaioneKL752nQj4rHMpWBef/Lpds9JKn9PGfZc0EFWqnCbNlM2P5X3IKW4Cyz
SKbj1IJAb2O7RZU6egwK+LgALqNlk0vpwzU7KF8/0totyCraVQXZw4DbDlUzONUK
XzdiajL90eifogqWRCVGCiEbXyHhv52NLYZvYU4h/XmkXbodoxa7nEx7m+X0Egg7
XE0ga9WoOdcpBYEAAw1ayi1moUl7xFvczSV4QPEldTZ1g7QUlQTZbkZp0VVVtyaU
X4Lzjs+i75fFyLFgcP3X+Fs8LuEYuxjepQOm9iToRPSc7zvHAwUhbUGWOoeSFOCj
Yo3uzDl9gKh22QFu7Js9yjh0MEvFYVY+wGdQZvS2LNYJzsRpikSbxQruJj5kla0z
W2jMtKJPIRqnZMyMeJ6/C2t4O7i5CiCQG2wqokYhCx3Z+b931UFEnbKeLhDy9ErE
Fz9NA/sbCfcjQsfWpTdmE6JJxXdwk6OIW6D082kGVJkKp5uvLkGuSoXSRVxJcUz/
BxkCnVQxAdeM9lIOrM00DoLl6h50GZ+MmT5qbB6WtM4mjJdF/ZIDEUsAPDNxoyEF
+hhtMP9owpmXJ03B7SGqFCSMCd8reP8xagERcUfX12vToAVrwdeC1LUvlA6L5fA8
ZaxHYpWck7TO/2RzjsBESaZgNPNulcK6ae/9JuZTM8z7AUMTF+ZmY4Hfv2wrVJJC
21+cSi/HIvPe1C64pnwoMc7StNYbR51U6JCtCqW8vIv5vxbhUhEVPk0ns2UrN3BT
ZxkBCYg3qeP05f31tb2E2ItRzajVU/aLiZsX82sOMOYicFUg/IJOQjee57ejUCwI
Gej+IuQ8/fwe+7vKU34/ghbFnqMtqOzEnmFAHHwdSUSMSMJh03NP2+w42LrE5+ip
LTZA1cUN1cpfmZWn4DoghpbH9hIyCZBF0RUdTt39LOQ1tLLskPaNOyLUF3NUV5En
S+OZ+bKogbQyq7YzZC4Qs+d678BTJ2mqc9+vlFSKjHFw/d9OURgU/Grn9Wa1tOXM
d4sG1kfE53u5E7xo437YTzlmB1xZX94OgbB2F2J1974APCV2PgcRzGdTfxmUGLU2
FWyV+lHt89cDX6SvwpEGVPW8u52YGRI+ZoNG5ruQTxIM6uxXHiR8KW8pgULzVhjy
H+0e0wCtWQ7TDg40nHUj/bzNGqbNxQ127UrrWNjvV3FrcjrWPMthvMRGTS3J0ify
2qijCMJBw4hWyQxwUpgEBl9YEpfYSzQg+6NVzHNfsp5fJlMlh/91OAVTy094doKj
GcTs4OIHwj9FDOnquEJDIldfsxmTRE+sbDSLzGzIRmSEg0AKwgKrTROSD4SYKvLF
9TR/CY+A0acckSbYsuXxUkdhBwj2v/O9YpEV3eJd1pfklmxHYHgpw6QHFDJHGZRM
Tt6iqDGT9//couibY2+mufB7NDSWuC7MiimFFxlUDuuenDdp699nqUzU9ZdQreba
e0qXezfQ9b/lsveU6RgOsB+yoGRHoilY83WAUpHpODFB9mopJtGdCx4a5e3uEoE8
GfflC2fu4qguEikiV1PQtUgh47fBtpFcvS8+LZXrgirGbyFj3/f3pGHDFwdL+yBF
XjiPBFGlpr257MJR9kcbAFCYQ7WDVRqgIZ9qrTlR/2N5W7ZOPOlDt7Ve5JbLy91X
GpHjoy0sTgKnUH2JOfdu14FuJDSoA2Om+ccWWYFQmFUaa0R/qBEB8usHvSnQxKoq
jlANQQ/p6P/cReqyGeeRkxonXHx43CUllSOuvbXOXMR50hO7fqiU7iz1Spx3wrco
A+q6z/ew0avuXHtGh40hCTE/CuapsXot6evts5XD8lOHJYggESP+37hqKpNIW1Nh
TBtyR2pBsyr1TeDexXgOVFIOGiGPp1p+LmgVrLWueFPac19LNPnOUKn5X+SgbdrX
h4srBhibCWGWf6YUpV77pjjxVVMUxFU/y1DC7ZjGhlnZsF3VhIHr4ypkXEuWEhfr
zk7XOY4wJoekM4XB2jj91ADM3MMDUblpIRB3zjGQq5y6U1WsBlWoyiiNML5nczQU
FbFFvDQ3KiyAAw9p/2MtJL2I8FSz2xkGkWLbD38NatZnXf9Dh26hHKg5e7k/kxCa
Ujc3xBik0dXtxcP2akLDqKhd407NOPXvSHrGYfnRt24JvwbPtxSfFvy5ZDZ7JfA8
oDOabhO3gDcpB8gLmoQeQypkc89ehAL/hGuBfEDTN4QDnETBoeaHZlWeuBsPC/LN
M10Ekk2pTA7hQUicr+MDBEFw4NjwJtu93loRtzexNl9+GRqr4sqQFPMOJ9aHC/zp
zXDXaQADcsjNknZY1C0Bv8I+L1pOa81S9dfAJr+iZb0ptr1QVvw1mHxImfBy57Wv
RQ/ibq2tvsv90PjlzMG+NwE5Vq7tCuen+1H2wD36Ac8EUQ08npAOkH39IJ2HGH8G
7nUjAjgcqTHXnU7GsAQy/NeJWJDiNWpXixPLVgvnPVYT1/npUzJP6SHl26ZQWNBc
fWtoexeWlVYsWPgOKOIpccTQmxWoUvM0zT/NhEOtN8sMaY1u7aTPt9H1LEUt8P/6
9kmbl3gYZjTDpwOBWTQXZ6a9DQx/LfUyhgLwOekgGwYWcvLifLLF+X9yErfCeLbN
lvZrjUPSvZsnNGyvH745iJrdaQOHc/vUm43xQfGg8D6jfOMkbujymQLUZ/fpwdXG
krsqwnRlwdZsyYMkM5e1IHdyPbrsOwvfElUh+zGOPdgMZ9jrkFgCLbSA/gnTK93N
KoVkHKVO7HWgymg+njgfzBocifvUm11/bqJVVfCbP6OVqUAoaqf8AIS2xI0yp6YU
50KRpNqfjUAuOBxoLaVZqFwqyCvdfoDHG2RlBek8fB7H0SsUfRmqI+kn1kZrUGAf
/91rOlgdX1XxuWgcVdSCCg6G4Ly1McyblmMUX83EsyDpb/1fZx+d7PxexteIeFgU
hifg3/31cMKD67sxSYhITXQQgMJp3abWDBokg0wmtRcZfZ2F3MS4fOmZqSKi4PT5
0T75j5z0ondDclGOsti1FIdLNZLmcjBWh1vu5oPRzGCXC5aP7eEe72lFKQdvHoUN
pFTPExw29pk2wnJ1u/8AEeGZp2Dig0IDJbglDEOaOimHFZi7pdN8Ysm3/qwXbqDU
wOW7Oi6XpakfsEZ9SD0ckMBUm0PShQdt+TXPl3WBKdCaju2+VGHVZegIxag5qxa/
0SgYBS7ZN4MdBTk+HZQNKaZ7YZxFZs1fme9NsQrak9ut9mSivDDafq7WyyEllKrC
M5CoWY8mM5O1TrH4lrUK1GpD3DwyBN0LhX/vlH1HzX8rdjQNcygboTCV1YmNS4wr
+9Gf4hpmasCAcDyTxh6490u/Zj9sh32dlArFvgpQxMQSmS+MFDEUVnA0o8SlrkGF
LbINtDI5N2DxlKr3YDXCrjfH2NlBYbxrZ6ryMbe3HTnjk8Vym/8h4QFaSAODI8YX
l4SJiM0mnjvF7ry2pDFIjdxASQbF7j+Hr2CyItoIxu6vG06+afqfrGIuNj5yrCM/
6k1+gFm9vR8EKQsqpaO/lqI4IZhGT3rxbRFUw0O3tUpVbLd9J1A8Gz0dXQEigKGO
S5Unj3+Nem+ihpNVlicLg/T481q7CK6PrAB4HZI0rqcJcJR9Qwy+ZBPS2lC8T6aD
EvvbOJ6r7GM2BSjU0EwTDKqL1heE2IYrAwA0yo4iKa1ImlxOBll0MxzNqzWXJA9z
FkIlv0Mj4VV1ZeQnx1+3/vKez7afsra/jNdVu7gZGV8Jq6h02Gu/7/u8P9CnxR3H
0az7yvw6ov+KoebQmXTw7wU06rzg6epAX/92HoA8EWDmC1LezxdoYLGX3igkpz7d
qdnFS3wcy15U3wHyizqs/t3h/yAm6U39eVDQiEN8R+kVyEnYJU4N2W69VhznFzVO
Sj5gBNOBPqbGEzn82SE6zgr6pPcB2a58MDyjpNbEVPgk5vE/6B7ppw5dnGbMX4zF
V01PgmuMjwNBBWqENGf28jALT96m0RJw+j2v6X00H/STf72BSkVg0cAiK83gAKg0
kFHNzyZthrwDgwctiIHxabH4ALX9oBajmsnZReDHZyThyHH5ijoqD4hhK09we35N
NO+0rbWxO3kgt7EnbtfIEEKsePhryUt7BFKah4kcklJqfcP+QWCy+H/n0Z8AANKT
3du+t/qjwy+o+L3KZKW06K/vrwF98pgn8V6VIIPefFPCBLVsMaIRcEVkUb1dlAsR
7gJI/7zcCCSMTyt2NWOogiuIBJ1PXs/kENbv7xCPtX0bCgn0kTUh4jMVRjFyGr6a
5j2Wu7dYe0aT3/QATW3oZlLJ06KJMmk9pCyxDjZcyp15/tS0L0B+lpHu01pcUmMq
4GFp5rTIShasRXWLn7VpnkocMG1JWz5XCm+lCvuuNx+QGQ9gfE0M8D96YhHyRjUc
Y40K+9RUYL9lt3mugrn1FGjwuADHL/ibRKCmy+l/y8jgveOHhceqENkhMlik6ipW
jsHK8dWJnvm3FjjwIgm/Bxzbuh1wYl47ot6sj9B+W8J52N9PeDMEqnil2IQ+n4s6
8PuRl8ACiWPH/AN97DzX6CpLXIqjU30DTFB+jUl02btiepmhB+OWX3aJ397syEHm
E9uL1of40upca0r8SF75RJKnm0+Br1gLCpg4pdftF0Bq/khvLwsClCeXozdrVxmW
VjWthZAYTvUuNuY5K284clZMOpOhzxIDaMtv8ymYGWme5ZpsCsPUtFCUrdFxpa6Q
qOG/jmWzh9QvTPjeq/PacfVNuQ/WXDHNJvOdM90cV4xHLE4fB/yMZr0nOLNQHnh1
SQAx9+MiQoGoU+cXUR5jf8PmfV9Sy/+YnhWu/fMztSf6Ye14evyuqSm1wqTsY28N
QxTar32aV/Z5A41WQei9GDmfpgwCsIHc+xsDvdLxMVFtwr3Bo8c0/uZbgIYSa3Rp
s+AVQZtUm09obQ7sdYgJ2NDD61ZhRIuVjxJh/LQ+9oBj2FBGo6jBsoB5tZIX7xIW
Nu825/RyVIA7TYrl8XbgwjjmOntM3wOpPD0AGZYDlJ3b7V6tNdFy0gO1hfGJ7Kpw
hpg4z9JKLNsu5LvMt5GcAaFMS9KxwIpyY+rR0lQpqEBsf9lj1lKJV677GcZEaUKq
ognNqVM72eE2tckTJB+NpMhGJcKteDykz72WnnJL8cknPwsA51Epd+D7NEbvGWLT
sgfES7hWyRhMMKh8z3O1cBLCaTs0tIEncRPf4GsQlPossTkBg86tujVQjK2+1sOS
ZYNNkjoA++JqDDdK5lzKSw4WDuDlU8Ndm21SkUadZ2N8AzDMdEzj8kVwf7AsBnuG
BgNgnCFaUROq/jj+NRCKby/MMOHwZl8dlkgysy9K7aFg6zjivJgX/+JGG+Bdqn7f
3jX2ki0JkAbnFCpX1bc9v82PHKztnbMJZIxIaZ2qk1vqOsaosO8FyMuZ8cDs03CL
DkuBdIGzdodaW8MIALaQAauN+b21o3w+rN8IqIO+ZIdD7AWvdDFUwLL6osxGA8X0
MpgsjKIIfOga4ohJxnZ9Mn+VxrpqW6aLJDm1x5s+TqZPd1Kbwu1odCqr261U0kug
8RZg+HA9uAA6MKkJg4ynFi+JfBhJ+yGtB+zB3yETCbpuwN790a1oKzxj8OGAkN29
6DbFLaQq/hjdqlpOoj7I32VmafSfXLFKX/ZFkyEBv52hdDY5/Pwn5b7Lclk3CR94
l8M6Jxawl9WKXG2F5yR/cXJuCHZ0uuCZ6FNIeREsSmig6gf4v2mGEh+j4e+BZ5PD
OCrVdsuBxDkobOHAqwPq0xXP03qqOwyR9/lphFF75suvUhZOuJxEs9Aqc5Grje41
16ZGt1gt3sca8dFhkCE/G5Kk9GPT8IyTXaDAQCrFnL3lh6HBcpkb+8sc5sP2Z7ho
zWo8BWbMlU2KKEdrDp32ljgXqIHWfVxVTzgdPzNniU7bfm3/ITLjUPihUCofRQZ2
E2oT/LIDHkqgkaWTtFn1LdWa0jieoeeNqev7E6DUd0LGwtdFmRCH4jEISyC0Ko8T
h7hi5Yf6+Wo4woWmgr0kyLmLJnMHAYMYFu5WGEc1TBbLHsV9mhzTgajY2WVXN4pt
Px1qZIQ9enGxhkk+Nkz8FiyrHiewFF9Q0zySb4mse3LOC8+ozWNJ8yIMAVE34T3C
R3hj8oAbK1YM+VxRAJIID3IZEHF2ChLtXpMUZcaQmm0fI1mJGnYZBZgx4oAYXbZX
xk/oGzO/OtYX6fuQ8utHsVXJY9d7XYQShhb3IsmNALIjt9oXUqMuPAydCLBJiBDL
sbThj+zZiwmT+Ot3MMn6xO2pVHNVZFOxOD0k92OzVxrOPEQ2CV13peB1TUQJ46eV
5eOyUVoIWmxxMQflEg6ftuM/ouxwdnDSUl/FI+8ld00lfE9znGsmrFKbTEciW1lH
Zddl0B6Ml72CDWH9L1xr0mNY1WDqd1PvR1TY03i4J4prgWyzNPfrr9UmuLz02bbN
FmCBM1yQOl9WR4luIcIKs3kWOmUuFdhWfx2w/9LN6dIgulH4u0AB9ZW28Lww44kT
G5she8RbWh5iHgGn7JCZfqz6IeLdFhYVd5vPpRHlcm7vUo9xGd3/L4uJr2L08a6y
S5eNja7CwogUCeCFCPy5eCQHNCpjTfstAIynQPytA0DkzyXvGXSSLXGxmyUcGRic
/5SzMr7R0l9lHN5OTJZgni8W+3r5EbNqG5bmY99VMdtqiDuW+J6nluJAN7DqZoIW
3RfcO8pCQ46Wl/PiYnrFbBsV16vsiqPHsoYqvc6sYK9lM5elYh3XBNMvlKz8oyMe
eJ3olMvfe0yDY99qLPjmE+/ZV7fG5Tnw4L4rn+O0a+NYI2t9APU8ft+4R6FZAELK
vE8h0B9CiRx21j9Q1PM0N9jJuMHQslKy4ftTVe1ugqNpH413zL1ILM5tqM9lloku
D92EX+gHdxvL8WN9rQIPsq3kG3i6k3/aBXfKsR+iF6E3HaXPCPBlWxs+NhCkOjEG
Nvojvdj2jO0c4B+SZ2NSlkVRUFHJENsxbXvdToWPkra9876nUyh0oOjj/4b8mkQx
TlDLX9srbdPYezHPF6m6jjF7TUcUop703kTNVSNtvTK7pESSlMue2++gPMGBKK5N
z6V7/HqlThDzUqV8yQORP7sbcDPs1o1neOHE+iQ/Th5YB+Vqgd61sPCrMPJ1a5a2
pcWWWNsnd8T2k5QLOvdEXNBtRzPEDLNrG3in4YrUgiDFwCz8BIVhWirkRdn7nWfR
lYcl+5iMi+S6567fBb+biPVw5JBnTJ39MnYJw9+Hbgjv0RDpGGcT4hbLnRWN+CvN
P0nOP5IFWYPEKXfUUHt2tjEHUcSt6PiViYsGPq4n+negSWpAH7ermUE7m1u1aYKg
VFMsBMm5Gx7cNuOWRlrOIbwZrXnKen4vMY7sIuIS4knZCVrzcdY80xDPYeRbI2cK
gabWIVwv/C0BFmuXDL+b5KvZokfvIa8ASkIKw5378OOfxq260XpZVZMobRmwckaD
5P3AM1NrvIyPcktEzkfeipkaSh6zqgIBbWfOZMPwhbQBkDMZZT33beHiD5b1I7oq
Sav3c06cqAe+GXfqOqEc5KH2W54dFe6HFV+NDIqwA4ViE5yKnpntE0XPMq/SM5Oa
3DhONZ6BqCoEhxMgTwx+dkjntMKqOor2hNdXPcEck1HfBCcicuoDNj+PLUSUNT9V
3R6gKT64XdP2XwDGWdNznOIcIzNGuQwNN7PWDmP6AFiSmUGj2VZFMYF+s1h+4HtH
VbylU4w4sWGkE3SxUNcAhRMkjfp+XqE+2aRjSAlqe/LhcDQM18/aHvoXmaFfPBxN
lNIkaLdssRkzLmqTjpgqfEGX2eZd2MAWbDnXVgX+IQUq/OcrVWgDZ0dbMeYSJNar
x6wvjHPQK5DbAHmueRC8A1JmXTDEj7sga71SkxV5b18ASWVwKpa0Mge/r1FOFJjV
tlhmVl7/E6zsFKvWFKnLUtj6EzVFodQlgGOI6QtM6VyXRo9OL75hZYEJxRTngkwD
a/UNvpv7YnMyh82Z6m0BsPUoW00fNo2wqebs9Il8jBgcstqxhMCDfGE7OnNsdGLU
TgJ8g8Ci5higKtJfv1lrHsibvYlxOjMCm/qLKp7SMzOrM8G0SVLyYOEsfz+4xLZE
p1Vw1lSMzH2isghqW46Tgz8Cp+XVy/YpXVn01CG9h++QDSrPMZFCH/+IPgrzl235
LFlPb72WMaTY/VE0v6RjwP5s4e516Nh8wUjsjRMt+tADqXQUwhgBANChHG78uTlB
C4wKv8vZVr4v4cMsCUE17LOarHTDBxIigAluMO9VHm2f+cN06QmSOtCn/swTAq2Y
wbN1Jm0SLLlJFPNwGBhcCSpCsyrY8ZVJ26fu70/RCrWVgxtLVjjCPLcaRsy6we2s
oUD9RUTru9/faQGesUVICNNrrWe99HfNF6lxwRglJ78MnP6PYw/9U+MihamL1YjL
QoUDIXVoyiZuv49rF1FqM/73NsOelhujtiRaCl5b5C9El+siNFnZweWOe0671giR
GVbRdUhkrbGxVAwTOM+GGCLMPECXcBF+HZXWwRuFHGVMi4EpYn6XZzOhg1iaMQgD
D9jk0amYBQdaXUunx2liO9HcC6V4ZyEAHtpRivs13FR98PzFSnuDVT9uHnygOZuD
cbA+UQemIP/vr66WCmGeSTFKuQMo7u83YXPNdppmchi8ALdMhfp/zHT4fF8D4Fm5
F+sYWtzDxCfK5oml//MHe3bOomsE2brOU9vyTOwuoOXj90BVvQiqPt9WfUdjSDl4
pEwg9hCs1dfd6EZzUj2x3fTYFE28jp89ZFoB8/a1Q+piHu61wR7Isx8QdlOlnNfJ
GkEBVRnvb8oRjOg+Q/pE17USbyaWxzErPavjqxKf9tDaQSfvgFIumETIYYEWHJuO
SudUddtUlrTpK9NIhoPuQyzUBdWe4XKqmT6ypBIoG+Jtr0OQvutI2IhuAq8CtDQh
hjW2wTgPlS+dEVUXhgoIcmATKze35aE/+gIO1+8+tgwl2YS3OKuUZHEsUMox19Y3
BrdE0SURhFUKgxCDNiAV2sVtIPPVU5KfbLvHemx0Bto3dkHtJmMW49ePDET80w24
VquCeLPkT++StHgdM7O/xrluMFOLzVnfmLfmJ4rFAFoPPX/jgEgUt6f1SOn2lKSy
Jd9Tj5QGNmUvSzSgQqGdRe2bBlicW+kokW49t9HlWMz3IAQHKUpG9CYQ+xk2Eeo0
7hM1IXOx2e/+FE2rrMcGE2cwk9YHTwkyyPVxdpX6MOhVd0NlqdVqSQp2sQGf6ihl
24aQjr1fi3/rPunrCIDLLNKKcAyC8whrhPaSGbA44eKwxsl3LOSr1uZICTDOTnul
WUqQq+ubJbqJMccyomZF7i1SQnNTCxQ+bjCjMwMXLt0n0WeDZmcRIHGIE3wi0Rex
drfuZIdLoZUH9CmnbhAu/S+A6igVKLA1Y3MF9YifbRYKGNONFk6+naSRNxjuqKeJ
bIkP+t9LrlGtvoMrsiNJ2sM7eYWIBbdeVoEB5wsqzFUvk5BTVVUlgjyitpsYaNPB
QXVESSLfNmxHC/LWY6KrG7FCP9btnOAMsRX6b5VN7lvN4dr1fK8as3R9xCcTGbOx
Ox8WLXx/hURW0YSJHHoAxcy6OMe1FqDpk7gxnjiTy4zUjZJAHRQruj2FMa+8t3dc
F2tDp9IA2jrcJ+SfyFkZNnpmnl3hIDq/+iiArUP0k1Lct7Nc1lGuX8jd6StltiNn
t/jYmaaEByag8E5J1JAJJiRneInlqy2N0W/OsknR1AGUNWZ5abnWvNlilpnS7DvN
YxQWe8xPzDeM+2Bgttq2v6as2XPkOSWrH9pxNS7v6SsakHOcQgY8/eeS0SAJ3o7Y
8vEBIcjI1UV07FoAWJpe89aQ0xebyfz099x55qMeueHyMAJxtzVjEezj43Hcig4F
78Afs7NDtlyCm/N4FWcXg1LE6gzrLN42EfeG7UZNm+AiK14ZlYkrVjswvpfG2b/I
pAFT2u4ej87Ba69TkWlAnjN52dwaCHRcUn93f3QIDWyX3s+7EFaJsucPjQY9jNac
cess21LyGKdW8zj5IKZ9419dwnaq0cop+72Ilzo4/vU4MrA3pdlJ12DntomvCg6B
fkTaV4QY70R+qEG1ny7H5Xl4kVBO6ZGVCPvA5byr7l2TZGyNp12vMDPzJvzR3Fgi
d2MJn7LlIkT4J9FslGFRsOymTLTtkb6uq78xnwQtKaoK2mb++y9+82ZUQdwukRt4
Tse6p0j1YF5sixed7b0eD7ErBWwXOrW7ksYzA63ICi9dhmv0vg3dzQOsNtp+DvBz
DUz85pIa7AWBbLb61YaFrdQuWiFtbWWFlxj7G+x4/AbrqbaSOr19QYAmC7BAdsJc
2taGLFWrS6jqrwNFAIsEAJJRC6G+lhft+t7uxGPx1WbjkN2mWuCWzhRWs0uDcbqj
lDVMg3xe/9bXb3ohZmsAvHvWFYhP/dq5yQUxuae1WuINEbwc1vVwHnDcD7D4BC7B
n+9+NQTSLmWoh00XEZi3hOoPdScYTdj17vI9ESEXzm2Xh5Gt6KcVf8EyjUUTRjgf
R5Hn/siyZ4wJiZk5yi1V/+96ImSgE9ArX1YegLl3MS66NpiFmP472Ta2Cd2eHLFE
Y2hCaHigCAK00FJr/4xsS7jSidSmH45XQSEtzVe/CGSD9YrcbxvZw3qvgzPoYa/e
i+OE24xDy1X0xJJzJZ64mCVEzmCGX1EIlYemymNrpbNvw33M+qyOIiHzhHxNfHyb
Tzjq0IJFdTMvM3mpnfSptClqQ8S29jwxSZ9IDgKjPBpO97b6xLRvnILlJu3Gl0YO
7zwcF1uyr5QyX2aI3WHybcKqaCbhfjQwWYGst5S1j4nj92TN+e+tDKCPeCfDRdGb
591rn19zqBx97pEh2q6pIKQTB7t5/AAxDE4w7ukGebh14R+VHKBCE5TEAy/GGKHV
cIiLgjDANtBsggef/ibFMUBUOylR3X4DAHxa9Vxt9Js/K1zTHHPLVxiONTowR14d
t/P5kWEVE0D9vMyHlUEwmdtQVqUvn7yQmA0tHRIsq4XnHGzLPvmPANt9q4/0QZvK
08rN6ThYzw9ej2CV6uo4/qwBuOy3KZxxYeaT2JoKYpVcmfgv+0jFi5PPOWUnFDa+
Os6erGqMB+76X9QR2wYaO01OanIUs2rjcsNV5lpbxVpY3u90tCQKBJf8yPNt4aDD
61Iz9A8rse/SU5iBH2EfU74gry2bTeaj6rGjuupxdcPCAxpg4n13Fb0OlfviIvao
DoCaD1C3xq6Ngp34JD4Y2Y/h0kiVygjvOWJ0IRcnLw2IR7NzP4qperp5jH+o6StA
gQ48LFQkoawa98ERSMyGSPQl/1eqyntqGaf/8XPtz4WDFEkAZeSEFkO7IWHIIQrT
W7qNgyRoKPEXZo60JKX5cUo/mCtMhU3WegNbMktgjzY/N6rhyW1csAeClv8kKYN6
w2xI+UyiF9vCQL3ohpaRRynRwaPKE4MSU3pwOpTKlnLGqaXFcmtMGWaRvj94l9QM
DxwM5cmcnXzQnLdf0dtJa1StyU+EqY2zB+0jK76na0a6mFJPcmaz51fZWP2nmtnB
ABfnSTapkKJi/2ttY+H0VbK2xByIR17wsm98a+ReciiWHuKSKFpQxrlxBxRaptqX
CS3C2jRWSsKjQ1CA6XBG+c6fiedYzKz0n4wWiuvcEG+IKgQHk+thNC2hx+UaZyJv
ZXRlzj1yAMMpsRJe2R17dO2kRL4oPmHCpZYqyNMeABHqS/6VWzYrq0mG3tZj9lTr
ZNO6vjBAPpIPxPaBVmZsomvkImxDJ8DMoNy8Y5jWI/6jwUavx7NrBp22Xx0FVCd9
0x//1xzgQKQk0Y+A9D3b+iXgi6F05c/dF35ZLYKEFriDgBgDCnFiPNTyJigq/aCD
YrpPpb1fOz3mE0xUadIzibf+EuO5DVIUo4p9YnhsHVY8OZQiAmh3asMoAUzfaE04
OcxXGSrnWbXzYPHuPGVS6ooosNjdACdsUOhFw5Z4x0YJJhUj+ja8/JCJ7NDZI/7M
2B0AJqGItKtJpc4hT0oajR3z+Xx5bq9xc1JedqOFROx2qrEM8+9oLY1hm9xqS2tP
6DLFnlw//Qunu9TpECAyAAo0ZXoo6C5xkQkI2swMZ5JaZveMwR1BGADCYvkIZDL2
LOAHNl4EMth4kF2z9XHgNaGJeUFquadds0RylVYcHhhfSbxYfKk8hfG9mKsjZmZt
ZyhcnXmy00d+7kKo/XHD4AHlvwgK1LhA58pWV7VLfOp7bOaQC49l3emkZ2YvUzFp
uvbzsavlJzGgot1Xd736o47dkB8Q22A7f5cP7oloF8e9NSjriLrlB/R5Z/j/UCcs
iAZ6tr3m1v4MAuHgbx21pg8BG27aZ7jaGdBo3tgZDoZ5AKM1aJKDK534Yb4ouj7d
c0DZ3RO46qKymXP8Xe7OcY+PlDFEhFW/hseLPx/WKPQOV6oJUiff/HHcRt97jNQ8
QJzU90Nq4yDZruMDQRfrY5vGQ+fnfOKye8qmGdoiRahKEvU4NYpiDZ8ojpBJCUXl
0ZlW5l9gbrSsMo6qd6QiHildLPZ+t6XUDJWgQUFu4O3aB+JZWfk6NI/SQl2uGGrU
EkK4Yyg9NA9uT3TJ2AV5Si/smQLSAMtgMkE0QTAe3tnmcP/E+z5Vy5ACjp7rK8bm
5q+A8+thLmk72B8M3IT4AW1d8zQJ0M+saCBs4xqSCi9Dgac1dU/LckuvMfmSQOYX
8y0dbIr3OVUyMZ6RVzCsNPHH7XEEjmfTbX0CRQY+sODiWdAX/W8ioS1qelGHD8Ox
ZbYBR9VGVoTxjSpm5Iddyb72Vfww74HiArKtOc+c3lM+B1DTw5wBRXRjr67Otote
aTlN05NgPhRTdNUUIMIJVvSYfF9hdNAKgGbDUHb9fG3TZdsdLCtpOZbccKOI7n93
83oxvmE7vtotqTsb+RWW9X5uDKBqZ8+RlgxGPNnyaQ+avK26f6O7xDyHiEN+44r+
28CbEyGEObqDVlVc4qykmK7VoWBj00koItgJg6hEKWQfbOoOWxAFcuSCZcK/w7pl
KII6zZQlIgwdLDGAu4/e3JphZEr4lP46UrmVasoDD7jKMilDLP83fyzyLWd2FPTg
/ioNEGkn8U4jzF2qjt8EJo15i6W0NBEanX5jLFYt8XS5Q22uV0xPyXu8618IxyX3
zaH9tjLk2wLHduPJ3wyjj7n7iHv+JTqOBulj7sHUfPZQ5qNIMClvh8mHqbboU/+s
uuMKcdb5eOERjVYS/W4HKwDcwTCjtQYuwQVmY6DmMso8+waY2bHSiyPTeriUWBIc
wEq/VcP8f2lqFDq9InqP6nJ8vb1czWH8pTbrIoQfHdYvgteFvEY64fTkQv+AYjC3
GHTL2H11MgeO6vINyUhTVM7SlkUyTdPxqsGgUuQIE9p2Xk1MBdwX29SwqaLGtDV6
nOil1HhpkgRohrDKoMmleuhS8Vdf2HJv7YKTd3Z8Y91MPZ9noD0tlsnY/ar8Ol9/
jwRd/jgBTSF72c2YGOrhzZACWmH0vg0BJQAdVqJcUv9hV1ZL26Xgar32u6vWINIj
I21IIWaKL0F2ZIh8jyy+xdiq9hvOJR8Y+thXtcq2j7u694SzT+1hKm0+UjdEyzjD
6mxgFk+rb9pHn1Vpa76uQd8eEqHimSylUucGM/4YXEzzgWJYBIeojLAUs87q31N7
LXDiV8uxQngZt/9FLRBKZuHEv3IY+SRmaTp3E5HmewVpQ55WaKEql3yIqKHCVtTj
2XxbD9zm2rQUWdgEeqeQKWpOKAK9oiNC9mDz5qYnZ0QApH5gIw/V86QinF+WBNWL
sZTvw79Qv4VO2fyhv2gar8z2+5ib71rnZFEJxEekRNaPkFWVetTXgCq41kQjrf/v
6UFdQ5vOcqRZEXWeLNfOB06ZSrhVzz1Stxr4qJcLtbSUtYPu9rHjSIu+i/GIN3ko
ryCaRui+qo6wVnjHazySgwWNvqD8Via5ISeF2PjhJqeOLo6MS0ipfk/XBCpaRWtU
hvx15c9FhFt7BKcmJ7IM4mhYgjVe8D+BEP5eDynWNiugIq5eL/PoOtA8dhcxvla/
gBauCidka136ZTXF+0pNu2BG71Zesv3e5jlHRkWfbqGXhk3oWmrMbSaKcj+Oc8vW
Uo8hwWOJElte6rwh2Lv6+qOgDQ5Xgf5bjfPUTvxmQsIzHxKx73UOk9PLb+yVvA9y
1+96/YG1r7SZNorcudQ13YcrgvgD2J+FPaUd4ARhXQJxznCIumKrPBdOG5pq6gUb
QcwE38RM/cb3EB1veOh00YhFNRt9ICUfJkRirXPTJHaA5yjBUloHMQFYyCv1CDP0
KQ7QuN4pIfyu0txlWQx8uV4WPwfGcoIffYpcYzxxEmYaNDyOLosABhYawGCfB4ah
ZLh0YSgT858X1yOv7Ey6b5hVT/35yZCCUo739WZN39Wz5c7Ove5Hj9v7+qyWVxFb
mYfb7Tk+JGVDBxkVbmy+pSlBXwA/15TXI6HeVpGk/WywiTm4iE7GsA8F857a6jPp
Mm/NsIn88Rjpr6MLyaf9en9mCrMAtjDCCSFJdQhWoZpnLtDC9Kx4j2VYhVmiA4g0
w6tNQYWRerzwlktQ1JdMV2+1FMEg0fOEs/YyjvnAY+PK1zWoL6Kyq6G9CdXZr+gX
wXw0pjo27Jnh5YQL5RHjjL8BjwuMbrQB0mh0c2y5LFHjSxe5W2PRJditYjnfaBk8
SYTaP0wGsjelrAfmOvxv70XTxvREdxalT5i97l1Lr3eMYy0a9zGAbW1EdqtbmheT
Peyi+S4gKLhta1fpTM7cTcl1s/PEbTL3nuIU51VelgnapEkPjpxkeYhYsb+FHbLo
LW2TDMFIKK7aa27ZaNhzQtOtsVubgmipxes8SBMynW126dPcm2TQpV5cIdpgIITt
FRiwzQEORBiixd1gYQQ04CsYV3aNJ3hz8M1na1oHVpIQeZvmRyrhNByoGz+TxgBa
oUxQY9Mp0WREYonEW1RtCDZlbh6RjTzU5ij1a8eDTmEEtlzcsfLTYotFs+0AOrQJ
hP1VrO2ubq0e4KvVh252Tq4/6sR9DMg+q6+Q9FqrEW66L5rJq+gqj+MWQFTw0Wh1
nM6kdc2rugFUKAuJdMo+Fk/kIOzzG01boY6l63bkouYiOCeGxtLAG64vDxTYqNeD
j+n20J3BLeXsIgRoqewZcaLQVYzNUzzrediN57AHZIpPoBlIkz+wWDLY9YbGKWpA
SvtSTwi9n5t7PjSWMd378u+JbRJMvb8B0qx4jVpFO5ONLfOG+dWRFrYqbNdMnu1C
pvGQdt/SwZP9kPXnT36Wq/JPgvfSs4HM2N+I11e3K+UA+UtMqvF4PGk1vt12o5O0
jLI44zteSrhhVvKwpaMSzWwhB2MrpcJht1Qc2ZA8KjdZ8FBn34pELYguxnkIJOMP
Y43yU8RwI9OTkgUGUWEwol6yP7fxUrTKNWsShhrEdgIqtermdnWa6Z3W5CG/DeiK
+lwCWccOlKal2KYWoGVyKP9ddkIcatvdb4su5BVMxN/TnqWZApYvnVfdWhWx6XiP
Lue+EmAakPBiM9EzU+T8vNTIhjpsT4zXDnUpMXUYXUQk+d3LuEYfcZr/WLzdvh0n
mXtGBYJwM5UPiX8Z0PnHaohb2Kb2B1AY2BZVzwvXXUadClq7ZfB8i9Y1paCXNJqf
9xZ5YsaqBtvNW0VyLVnGclIesl2d341ggBHpZb3tSFxbHFbgb/+NAG6W6vdyM2gt
kfcnxvpYrS1aoDs/HSufyj7cFUnMuZS3QH4cgUG/KHxqerSLbcCcIZtEJqe6+C/E
7U/qDJIoJuQ1sWYZaPduzJO4ZlhCvM0bA4hszBGMloVHCFNZx319sArKNS6O31g2
7r7Hz64ZX3evgct3/CbvUD8/ZV1Ek9Y0su3+W6cUzLmdVPIC3QrYyz5Xb/dJ5mS0
btzaJUtZGPRNvW4XiME/AH7TOGpHhIa1MbLIF4PHJsCjjyKvZOQR+hWEsZa+STJ6
D35RBzT1xt9/b1v0JavXQotidNZHpRkPrdrr5X8rKBhrnwBtnUjzoR6IT8/hSjnT
lYukYNsPRE1sanpT1mrU9OtOBlsjF47qFf22hug5acXnTVfJQqvUTom99XbpuqD3
rfRD1ZQDFU8tvCOrc/b6lxEiD071gDG4pbeX0EhHMAbCWR/qBJIenglDSwek7xAd
Ab5jA32e8LYn619+5Xwn9HFbWyVQXc78q5z7o7DoWvGwU9QkZIKE46iviGvVO8vK
QUNX5B/Dw1+9wnyR/nDGxTDXSfDSfgGdJuklWhsNvI//BAONTXulYv8RfIEVW1KF
XMFgJ0r7z9f0R1ePZSXyby9EcUs3/6ni+8U1ExwyN9kZaFgIRlVDmA3qw2J95geQ
m0lrwWP0fWrLXTpCNpafJHlCyyGkBYdjFP8tSBzbtHSCQVnHDYMkl7Pk5e81sKnY
towCKN+FA6FQTsCQAcnMQhI5Kjz3h23IBg47LJQl00k6wIISwJ6YHXPI739slB+m
+ZV2450Io8bk0kBCYLTZXwRf6s13t0mxRtSH0f9JgGGIImHWUg3gC7hc6nXWj/2J
80PZ2mYmZmC0vjh638xC1dRXOcSfs7WRvyPeCND0okW6K1TK2e8X+zwIB4eJy/pd
A4VzZ7ZWu97aUsxOLBVSdlA7vNObilrUa+HDrlHPc0f2wkqnsaEpFFl5A+L8ioI6
uJNoi2iZkonbpVRhZi0xgorhV+8KnEGLFwNeQEwpGxMiym/EbfLzW7rluK8vjgig
h1BvwseortdSxD29CFSkezNp+RZG3XMvv+0w+nLVAR045hEK953hFNNXlxEPi2Vd
TapNEHIRPRck6HNdVLlaYvPfZrYnX78uP54S0gpdKSq4YAsgQhak1EN2Uz7For5p
UzAW6ZQ1/BEBJNTG+g2Qqm1zv7UCfco1Ke6pvduCwcbFUWeJhlcUmW1tAs3hf5mG
eJ333nINHBYBhoXW5aQCuVpZbw2s96D3GrcrVWhVm5rgNQWowj5lCKAksH1R2Ddz
pwMp/n+4j1TDVEJegTrnm7bkBBMrFo2OcO9xpt3Tij4f5oIt2bbgSCOFY0blAgCa
ChFSjZCgftZuWAKp+TspUupBkNpRk0cbsjBppcD47XrUI9az5Ka71C38mVpjdsca
I+/36P16rsG7WuldzzMW+syV+gv7bi+jp8aGIYpb8KFVMqdMXSfamqnz/5PQbDwR
8n2tvz+/bYH2Ls7O1xib53RkefGCTNi+PnZgdrO0vBEzoZJKeCdsm8znCHFjnuqQ
goxEC3EouIAEbIsfFIXMyUgIrNCDVkk9yQIHnHDyFFlJTDmKANwPIHrDN0kHKV5/
uPZMldjZ1rU8yBkS84fwyNKeAR0qTAtlj3u6FfbaaeVJuupbqBZuASI+NXLnGIXO
GVX/ktVT0q6k9pmT+W9D1rOryQ8YVZoU1cZhOHYVYpGapHYDlvgfy7nEY4/Fe9+z
YF325v7T5/qlkMoZm2govUlgZH7gG1BclDWCUwHpr67iXJDQ02Klc4tXmPhkdWih
WRtvlBOHi5frGbTtK20axuy2DOtemd7QVXv4s/y3Aed0Xym+jBVFYdRcWemqN620
rFN7EfbO0XHwuW45d7dXKNYONrW55BWkvHKmb2qVsBv59KJ8MTn41/RC65QwjQWg
RWo5LMeKtf4gtAfsf3Sq6TG1/6Tkf1Oa44onF8Ku9MPV8iiquDzkqIoppJaZ3Q4O
IYOQ63ZTB7a89IOa/a4swbB3/EOOhMeCKXl2rH9/T+E6eSw8H7jerrhbvjtW/LWC
/bql/OlPc+ePCoGjSAVL6QO00PC2uWRQKNUVtMieR/8XNZ1lur2cupZPE9RlbdNw
dBvamkX0hs1jlAa3LQkU24JZBwI3CZ3avV/9ZvhILu1y602m0lqGU1z9ZTNyBYI5
4DVAYkmmVpduz1UbJT78sUf9WewKtr7ZDcWz+jSao5IOnBEhcCKfkP4lEZFE4tfu
6woz18Q/khjeYaWGWJJDI7+cAQYJmbjMOnl31xen94JSycnBB4dEcvoNDiSqsktp
d2tkNFdYsieIioaSc/d+nIP423SSAJ/pnFGsC0AFUVb3fL5/udFyZlyJ9P47heOF
LR/dRWOCeCaUcQ8y2ceQ3hB2Kv5xKwUpijsBFUU6oTNgEj513u/SNiZsctRmIPRA
BRSSTqxMYIJdfhiP+q1mTy51U881M6Wcro2oUwORi1+1df2d4Y0iKVDvAqcEWXi3
KDPmymZlvURsWrEFhs1zUGVwnw08+foLtBrKGcwDU1qZCZXnVe3ZnxG5TELSbTh7
v0El9L2D7U5EM71YMKX90Jhu7eHDe0GR8k6XJXvyoz/yor3DrIfWvjKShRi25wwD
OTjXY99tH5+eNWA/vugvAXugHBj6aeV4Fs8lBXnKZfV0/zX+NHxL/t/c0FhErB6L
nbrXUjPufab3N4C82GJ8+6Lavtr/zInB6hG1GRgs0dNYWWwkRXAzEwbPV5grTo2s
NbCJVaf5/s8gHfej3LeGTGL4dpWYCAnNEFpFeu8eLTBgC14IEizJwpszaHGMl6Oo
rSFqOO0Loi3T+jwg61o2CZwDnsQ60vZzvmemNJO6mfBC3w3a5aGw5aHRGaCPcI1k
sSLsIKLwKZfkpXi/+KJveLhJD88s3q86LRgVjZJR1Lqn4WJAtjNI4H+JePOiwMf+
ddxIVosX+Ded0uOsOaBOd0XumfZ/ATA8p33W1PNOq4c8hztmfG65c2+mWl8KwoFZ
CjbkNoBtb9fIdPTUC3FRFibwLLgTFFpJNnW47G0mnCMQrP6goapChc65QpnOYO1P
FZPear09by2d3tQzmfHO7/l6UXY2c1ScPcYMREAerzS1Jdh8G5OB6aI4+ZkYEC9x
94JRd+2ae+98HGfCH+hyoR2FfnYqt2LCvP7QppxOHbsuzPKbIOj9G8uyu0JQOtS3
GEYtelOHeGYgXhG1+fv56qtBLKmyWHzxWkjnqMpK/GmboR2DjFqPbZP9Mg2n+8n8
gwO9JlnBSHT5EofupBCtTtp2LOjXhHW5+iWxuB8NtLI0JhYUCq+4SLMwv7Zf82Bw
5C0U70NyPLaxuCxEOZba5yWWYaDRZfKjC5gzTv4dPg/IZ9BWjYSKdi3W1xU9ZThb
xmYG1XHczJjZ+Y1xYv2+X0TYz+4BqOH5I2/Gnn21vUhE2vGVOYa7EGcAP87hws4k
cP1LLjYaV3RvRf24W93+Vtx1k1MIsgRbY/LW0h/uBzYjr4nH9N/UnjK5eCpCd9Hj
Jt8reqLfQi3ITISHzGZNCf7HjEy1NYBREr2owfmxMxCpAqOa9q7CKw7bSQpV9Oyr
KHTbncEWCzUQ0zd4Lav4fipCnjlElWi/GVIzE8vbbldCAM5nynNgGWWwyU9HTcuC
OcM6OwOW8jSXpi6puIMMB8YT97ThZAZ3uabd6I1HrC5JD3zHJNBKjDruvVeb8P68
g0IIFY4wOhYeMsncFZUJyJ7dD9TNe1qg6z4mkkZRBe+1Bc9G3rIVrCQXI3VbzhDS
0WwH6wGiYsW6LSvI46uWAzxd4kjMzFtEc6oKMbapJZEwwYxjGedNhFIpNXiaG96O
qUatyNTJ7NBXGJcsUuqsHe4VaXcQAWNJSan0hMbu5Ygjv5yIHlKGSPwhI80zcvVO
jCHScFgizVmGPSXsjQ19qa29dyqC1JUi4d090a5PVNgL7DFZ82pWWnbGdExCNTSg
qLw7WDbQgLHjG6pV6ttv0IRboYducnCpvtItKQfgWMvNVKQG982YdKL0HAmBX7mn
qpIJflulyKF0An/yHrSiMNhlYdypgNYf5fNWJqcpO7i1aMsAcAIs970c4uRFy2AR
E70GVu3WqDHByoEqUhyqpNcG13kF+ih26p5PVOQjY2VdB+w2QGPX+LDdJ1w/FHik
tT71/5pq4ayCBFMJ3OQbr+3CUFBUesf78+yWTAJyt+qAQx0uYDvVc+SBRfXcBB3y
rfjxaLBIhifTJnE+yaWkAzdvtT6ZX7wZQt6EXFeBsiCQfdsAE+icxH2Z7bsBllG2
AveiesrFEmA49ZW5TFsdknJ0v4iXibpkpBySwKNtOzRNTagCYDHavsZI5lyztLJb
PuyF1PQqL83s/BknKvFTMrKe6JISoElNQx6BmCRZI9e7NLpDxUabO+EJK2t15ZP9
cjNpko2Tic0Fk6lGKRYJV/Wt8y/hLKppvVZfVfUj+73cjTgFv4A0/pjd/oiOgvEF
TRITXc0n0y1g0O3ePLnC0ys6tF/iIO3rJbbsTJKUiiYoBdHB0S3KcfBAUn0Wt9oH
g8wAyvAk0xQjZ5brDExLsuqA1mx355JOpzSP9JRudLYZYCRX2CqmbkTNCbzPHNDk
0ttIhkoBZMZAVGBuoxBwf0nzFgM92tYaJyfbuNABbYfExs/fH9JcDv8JPkIoimuG
Ge7srIeD3oAJWQTbGYVokbH8OGERmKuTV0yMTIyvOxd2EQRztYd+eBFoUx4/pP5i
GQ2DqGqxw6p7nFpvuIro3X/OssGMmS4tgs8uymo4J6nCaz9Xg90YMxxVwnB9Y4dV
rrbIh0MmxgDJ8pP6Vfu8ANGraTPwaDVApN0ueJQrGW5tNBKVqB1l1Z3+8w2/z0uH
wpPu2saV0GH0CwFrqcD/v8pZ5fSLbXwDcGNenML68RSyXfUULWOC4jKWdFeg0obl
8WhJT/r1YbY2QxCgKM9I/m/GJtGKkon4gKTaaIqc2qE9XainOfOe9ONQ2czbtSLq
fs26BJMPtnjt1rFLa7Qwj17nRpyBX+7kTL1Tw6PxWdz8zBTCOwP9stAega9Qf8Wa
wYofpKhUWExzM910gCKQfJfjMDwrSxrR4fDFElVh+07DUWEw85acflnnNGn/PUZw
Vsvhz7mJytpjEznRCjoNv8j9qCpzztzh9XxbZX9LCGCzozKIrgA2IewaiHolb7Hl
0oP1K0PatwVMx9tJPPbGlTtkOMRA0QfhT3B3RGe4pHPBNjbAsJoPYUnMHTUbeLLx
vMMWGmTuJLo1HDgRf3lZu40fWW+dCeT7LaBIhl8mXAp0iTqgUjTyvaPJdXX+g9zV
LUP48b/GHVcrhMLBolVRSjiYkGNHauaN4r0NIPV/yI0xafOs0IR8o7pnN1BXt8If
kV9FCuVdgJZa9jWk1gE0YXvYfOaQa7PFP/eOhSZT9fehkcikDcQpv+I2wZV5GHK1
JuwnZz809iWsoH5SGv+uX6JlbmRZ8qCO7w33V+vMVjSWLP3XaeE9vpMscXFmifxA
OLvWXFFkV7cdFg9FV4f5DDIpplNFg0tG705/nYw0hlzIayNNEJVoN5F23e4qdqDu
alS2saQc9qLGbqqctwKx/6Glq2bHx53KoDHRi7SMKoAV8my9JLw/L3Uzw77krTT6
0/YKqm7fENrdgsZPcH+/uaZQdNWHRyaIbLitsxeooGHEA0tstXC/m+UXLnvVp9Gn
dPXr7Sxi03D8O7fyCR1UUISzBwLFLR0TsE2CZLDnzxdPIyDzGRBJTuSK9k/uMyl4
Db2rQ9EqQCDAoxe2ySauxQOrJTyts+qvuKeOLDHeLzB4jTFKqxS/7dujOuitdivo
S4PnGbXwiroA+aMRXf2GbpEuKVQ3miwETMU1Gco4h3sVbMkcO/yENQzBq+LOaGeg
Wn4sKT+lmfcU5CEwqPYyW56fanmU5ZZhRqMrVJMLOc23pF6KISzxC1GN5GfZLX3u
WoUP6iPuPQmz6x1eCdAs6XuET/fMwOBlza++/MH8iZMZlRtfqARZCu7zp/ce+TjU
2eSKUrzLHgDGfQ5mtnKYysnNNsOjJq5jTymDzr3uxqPM/L8SFi47RDyWbtxE4jh4
KfIEzb+5swLY9/5gCNKjjRxVbZv6H+Fe8YI/UU4aiEoJn8UDVYVuqS0P48RIJdZx
+g3Tp3KjGTvSKH1P2TETmLQsCIKh4JU2p7IQbHWzcFvNF3k7YnL2nfe+oRfgPbg0
ktc1SwLiQe+9nnpY48I2puqh0KvrV3U3FI2KiVrO00mkMGU5pxf4ShPn6wMeT+Us
FQUlSRef56f+6Y82uNvFxp1CeEtF+EAyYfdItPks2C/LIteUMNiHoh1rzzAiAQEX
PiHrl88ZndNpYtgXiTcESC0DOVsZWv3kYk4Q5S1BE3scE5ICShvdtbfQZFtILecw
f54qs8sj98kKktRXvIdeDuPXATSyze+okP2luIkbhT27wkvj3XVf1AlnE8FYKFN7
ZYXYhkAuKmblTyVFipVVRoMKaz2QON80ujsa7sSckDoa6VIWJ5oJUV2/71MsFAau
ruN2IlQvxMYdwIMViNmUviheSc8ogHbpjBTs5MegpKSa+UlHfCQoQt2i65EIAo3E
h0lVYoNERjyDaoQehed0jAUvjZipWyLBRz4p+WzkCDRSQTCfHTFEUEvjpoJoO8cj
g3twzKWMDHdSEhMT0CZkwPNtS5GZ4697gpETEL7sMQGlJOzcGuykMIrfZ9/vxV2Z
sN+Y8ebdvdrRh2TIlxVx5UwuUWmhcMXoXmRdfmtu/Cf00zrWzGYqFWdBl8Aln2EV
ra8nDdJ/js7PNv29jmyiawRccAbZo5BmvY1JNsoo+YBIXkKoCY8plDpLPtVmze7M
fRYqRXX8ThWD1ynUUBGTT+/rvUNzooujOW30tx/4/bTuT0JPfmsF6mn7OEmklsAu
4QDy7nRNvaTrYMvckmZxs8EZqOvZ0u6YX2vo4IqyTGC8r0YCRppJPBUA2TQIXQar
9j0M4+CFzVADCVHUeaJ0rruG53lxsEVqxRpRm2MsVIZVCGItA4xa0DWpYPAfcrfl
8MIdXA1PqEMsbWxEv9gwubrSxxOrz1Rzf+oK7+zv5OA81afXWspeh9/Kc4LZqsji
YTRV+EER0avK9r4qyxiA9OnAVBB5SF8wWfPGAzA6vpk56sLqaGOOLmx6bfZmlhzV
kK8iBB3xCThFyfDoyyR80SooK1PrzMKu6ihizFdwJgHMyGoPmkdOSBf0fPf1veE/
cq5vgJEXLBNBfkL1yzWIAwG5vmHnvP3iyKYSnafDdSt1ZnFOq5ryaI0RL2pIzPy/
AdVJ6F7FYGOlzfimtisKvRxcmeV6rWgEWCPmjbDFvagEKaAGHx6z0h1odiKaPr7P
j5g6qZw4152W5CYu0TO9VeQeTomu8oLBDlakPzeXmYALA8BPheZACAq5CxrvXTWf
udXpPhFNigkr8emxRWWsFAHS6AFRlgjgQn8Ug1vMBHbIwPJmvqjo6hTvO1Qy6095
zWep4o7dbzz9Yk1IfiSYhftV1sQSxjGfoQC/7MFpHa9Sd+pK4Zz4fFi8L9l4jPUK
8SGrknt6UZqGfkteXqXFTcgwu/bi8CK3sVDz+OqDoRzPUWgcDTeifT7uQzyWzv6R
CRFZysppRW6+SjEHdpM3JCqfxDw71qVq+CEfitVZ3MK1hxE0ctQHLgRKdno6q0sN
mY3BAzmQnevHzkhhY3WRauLbklvYfcKs2ewxE892mu5YZmBAM3sFHIGLV2hRmASL
94QUZG/3wha8HDI6e4ODCgSD1adw/nBoEb4XaEGASdYbZkfTN/DOhm0hLjKyG1gc
RCo2awSuYNdUAhpTJHSl2u4aMs2RvVjwotmwI7ceYtoFevYyEivXlDeJ+ClAG1Vf
6P8ojUDNlZMvksTbF7LugQi4KVgVkQfT9ACxYRkIpb7QU+sAKqJgYEEJ+Kp3ei8F
VqCAbh4i3SPNLmCjZ92Vl9UgkewDHM/4VxoETMMikdaxruvbEdwQGZb2DkpNRF6G
gpkHGmUqEppYJJ68GxgMOoIGPxKl9/0dN1dTfNklZn3z5iovWjpaoUmppL5oIKgP
czNTiRCw74M8KQbWNjRYIGH5sy2EjjUHN2GSBgBHsldxvTSLIc+oUIBSn8v27pHE
jrbUKezke5n6z8M36I0gi86sEEFsGjNoGAi/NSAvw6AP0RqjyIRe7l/dajj+vjOJ
vAE2TN/uVZxVp4B2vQsop5vvrSbI3eWjrbUyowlzkRSylF9gQAKE+1UH6h5Ha+tc
vRYstzYax8GPhh/gddQM1jlQByZogwBpK2EjadXprO54vh8Po0l+nP/zf5xnH0XW
M0M032uDRqew8azNMACEJWcNqDKCUoto1nMwDH5UyUNQnFCQoLT7XW7lLzeWZ2xR
XkkrMd6JCj0BZ/recFIrA4ytCkQ7nFDkL6P4l5iU6pHJjcF8dsCLOqZk6fBPQE17
imUQQVKU6sqSTYwh76rXTWH5AuOLFb59gCnl+UhIFGp/b+le7gIvvRsqR64E4I7h
G09n6Hs0DlncEkvjpNt7f2VguNteUAJ1gjxwpAIbYoXr15gj4AuGVXDPKN+0QiQc
Y3/yjx8va6W9UAAdeYXUtFIQKBACyZ0OVt53OVh9oyyFkfQKxzDwsiZNWTCQ+6J4
uCM4Q/wka5sGIiRJSF81Gs/O8xKy272/BaPtVMdl/gFotK8cLtzqmbjoVFzQrtHm
RCtqijBq1rZr5Gs/Vq8LGpkbNrMbyYZKTqkGZG+k2AklnoxeAzW45Awy4yXsBaHL
mLSe1hM19AllaAwvR7E3dPCFpxzw6ihkzxJ7flYR0u3OMGgTJWCP/S3UtqbeUQOY
3cJ4oGEygHZ21uwUb38dz/5OnUaLOAcXeXXIZ/3hmBTs6ZMns8hoRizlfPwnDRso
O4S37pSqFocDmKi8AcNY9+CuSx1T6JzNlaY866kfguNB+m22BC17H6JOhbAfBK9B
hnP1yF0eaKELPprMkcPYz+6vxPT4pMLzPBcAnuwPmpbCsg+VNOWjYure/eCR+EFJ
VgyNo902A7KUh/nhSkg5nJiyIylkjQd2X/cK5MkPTNvOznSFgKC8oz5Waw2t/9+m
c+BmX0hhyOhjp8fsAp8TX/ALBRBAb+/b+rhfV6ajqhxX9XcBxCdlZ8qxplknCMhf
SlwvG8yQd3jM10O8DgGQKAI8FkOHZFRZg72A74Ei3+ioDu1T43gBiccxH+OEkiZm
z745aPyXJHCMmE+rsIoxd42fISOyEHqEmZV3QJJq/iYnK/nwWK/3VShVLm7oW4gX
LOAhce9dlpQ+fbO/dJODbCLKl8CvEFWxSv+9zdE94vDMN3Iep3I5+qropecEQxZd
51SdzuRNzEQgbeXPwuKzMMsRFvixDL8/t/Ac24wXvtPibD8ju12HFh/RVamr+PZB
L03BDgyhdS/v4x0bhAwTm814udlINY1Pvwl/n2Nt1eLCQ9EUqoARIhu0oKGYo3tH
1zunsfETj/UVLNF11tQjpfa7ECx7AU7crx6P1L215PVFYvFBj+K8kOg16LCPA5zw
Nv31WQdgAFFPZQU+xlJ0VnJq4J7Ik9Fy/i05tGD18lbjqh2x0jj0ETZV4+X1lDDn
lOc30+Wgu6SkaexPuwjgVykL9YpQGIOomQ2BfrQRynWWYSBAoEwva91xhN8rLrOh
hhnpbqzhZ7TB+E8hG1gjWFWnVKw4uGfP+s0szdjBo2rIrERVsWwoni7T6rj1G92g
vAA3QiTtXYczZbTZNjquYLU3ZqG1kmDqdWLvUsVcCblXL6YgQ8Zr4q7ecc3IL7Lw
DhPbvhP5J+0uj32GmBWLWorIsvWR4LYEdAYg2uYIheqWSAlZXfsvB+4H29rGMYtG
XJJs4Ltv8lkYHxLqgPV6X+mMFehM2Y8V0wrQBpypg1RdTTRWpRtMPyvd9IalB2pg
A5vPW8w1cWWbJh4EpnFAbVeVGbtpGBam17WW47xJx12vF/ZnSNCfpzGfsPDajUu2
wcVxwoYoZAmAW1oU+grILBVNlXwrmmLXv+BzXfGSnvGPkCzHzOKBAMjJG1VVWttH
lxk5F+mnv6DKpOf1FnbMRzTTQnayJxkOFAJAlsNmGkolUC8MrmJfmUOoZHKzcChQ
+uY0DeM5EsdR6GhcqoRQmrmDsM18kPZBPOaxrYXabFomIAq3R3rsipU0mMBTTajI
J1fxIAigtjUaEXlGXp2YEDFf8oXf5FNmQkJ7fBS+CfsNj9tP02SWbCs7yzwH3XF0
4FTCKOejaz2W41OkBdSugVqTaIAZfGOvIvrdUNN4ThTeUK42PCvZns8K+3o2cJNg
T65MrlAdFhWhwSL8IoK2VVokT2tOnUZen00l08a6Pfa7HDj17HEsFr8/K5xBX8xQ
3ow1Fnr9uKmcJyjl/JsCMkILEE2i1liW2aEfAGEJDXFTTBzrFO0guxU5mJ/FaUHO
Iy17bM9sv+Dzhh07qvKAoEP2O3tslk7Eo78cM6yTZXgp/RQppfhzSW5DHovoBOoC
Oi+4vtJ2+oVUDsdqGiUDuh1HwSGZ0uZmWoWKzno6ulT/LFjJZPR6jHkQMIt72ytX
hQAPexzXWUXJqe38dUVJiTCqEXk8iCs2Fa+VGPVVgzIcNC9vP7VowvasKtY4dIPu
2AUjyUF2aaAEfcotD6DH+PfXYou00FqdZN0L0NJ9uch0VTWSX1VVYUm//AZja26+
TZK/+Zrq50FLkD4m6KS2Wjmj57KIfOBkOufxcwhlzTPkfOsEqvpS9v1yIy/27JTo
RMkk8ZBHUR+tA7vwOFUw4vx+ll4EaXo0teQBhxpPkarFrjZLM2zakrv/fNuz/4Xy
HsajEvfwbzkVdILXMg7FFBWp4Gb6QzMyAtxSxmKsXFyYll8haGSvn23+EVGLztFc
Ml+jHkTPzlPl8Rzw1703r2f2RgEG/BjhNFljldkhTz6PHJQVJzh1Zys4bIFNZToD
nhL+HAPf+bl/RCf0YpYyfmSC/YPtSOQujkQPkZzvyb7NKowAm+Ptq9psK/+rW52o
Z+tEkE73pa1OjVUnuFqZms0kKoKPwf01SB0sI98cccSFZ+LFNdpw3ikxL7H3z7WM
kPDnjoQZmi4vi3ZyILoITgRWmZYGmM5BIjcv9ni59+fpnUz/caPzyDUX6gXWh0MK
Odq7QFTgELVg0iJlqmIFOXtiXf+wgLS+BFSthLEoB0e/wPBUpdveR6ruzNY3cAHq
2UTjJ3kuvfUEpmT9dJJqcmmXkyuNndFPv6VrsOYD27iplOpFptJCf2lmGYD6vrp4
3In7srNCEsLr4w1Vvpd4AiGz8GIMVdUSaXBUqDnxi2sDW1bPze4sptTgEauKiA5G
CIlZnOA0MSQQYNRRYaNyD6U5AhTRXXE1/OnRn1vFJAXCtILEWNEVvgzyGsXIxkc+
BXLWwGK475ObuX1U1H1zBPcUxbYjfB8ByUrhroAa3ENUeFvO1D1EUjKSkFuQnioz
9S2GchEzeuUocgtmHKrUhP+l/xvJ9tv35mrfREozukPQRyV1NQrdNvZeVMDIzC7c
3gJGZV+jmJSOVi1NL173UQSPsXCgUjJJ0TIYNzSSQofuANGxNV/nKinfDNQO1r69
/aEbU44jasPxRJn1oIB74+EkTUsJsnxtC8dyrCBd+j10cJtXLvSKPUKRX5YhtInl
eGSvDwv79vOENaBZfPShQrOrYnKbzBFxlnpTvKDidjibOexKiAyddDwP5WQBQx4U
97Ss/S17ZmhE/U4qB96xSrS6m7eWO5EhZzBPc+URrr5QVWQ6DNrbi6DlE8VylmdF
s/iOYMbbaIBkprLJsxYl4e58ywzwp8Es437kF+s1U7IAxYk3cATyJlsdd4N2iMQh
2esABQjQ3Jw82ZkEt+p+hxbaUvxc3TZmQLhD98ZZHqn1V/t6btn6krtUxW/DqsIR
kH3vCXTdnikwR2MTRdEKYcFSrsFNZhrQW+/WmAMVc8YupIEiQmVsp9tRlG8n2wrl
+9/8U1AyqF6bQNmQR8hIGBRCma2ijfTIiSBrUwfjVwbS6e5ctU2d3JkZ+NFsjFMx
qy9ILbBPzTY4XzzdqicVcQoeVXhnI34kKMnoxv4IP+gWhKSQHTjW5EwYH45MdLGV
/Tg1WhtDo1qEKYkESslW+xzUbhkxoy509yZ9v+P0xnNbcLPWrcTlKrdj1CKVdsod
x3GUKM1P6kNyafq541sX/h8ZVT3dnxkfH97Vi0b5nfbd3vx4nmOjV5RPYjWfASkR
zIKzvCRd5CdyYUfpXnmKS3gp3VpiRooctGEHQJk0xe3IGawlldN9nIGvY4ITid4l
H6MzgYEIbjNC+FIIV+YDaPjML6J6n3g0JKI3LYh266BSvoADRV21bcPeEB3dbNbC
QPKGl67v2uPFSZi4BYjYcQ0FW8xsn2xE7ixIhJ1Sx2Hzjcv3JO4/V9jduH+U5qIv
QbFU5qnb5uzEz0XQEESb8FVNU8Cozhk6vLeeqU4ailn5d0RlSYXDPUA1xfvvi/Qu
KuMI6GuammLBCEKe8DLPTz2kKDNe5+Cx74ea83uqevzoxMhHoBae7C1aKmVczSCO
eQzXhXTn6orwFUyXNfKLlaZm83q24tEaMSo0hC07SQeC6LjPIauqwcx5IAMSYD/c
dumk3+o4rLZABoulHrXF8ty1/r0WbOCyvUQ0o6b3NyXFn8vyWWssb0F0pTkOucC9
FQ1AkzGVg0neg4eAxGRaqNaQR9E9LNzs1R7GV1O/9A0w5JKz/NVZX3+cSqhW1aDp
8tQcWDqiCEYRpdC1pgWI4ekpLA13ZNjsarUEpxpdutp7ehAPTFMtLuYCiWgY9Fka
dohjfxVz50gJRPLybBYtorfOZXGjdHMLkDr7XyBuED763+D0MPwio2vQCRfVwwRK
rgyd2a5CpzQwMmC4It838iX22qpzzoZr3wmqTJtkwS/jMsdpsvwtQycRJvIdqGTf
vsy44ItOmSzlsWHfgPRUia4xHprk0bdXTPYB60LTbASnr9/8v18Hbelo9QKSeIJk
WmAYOZqqXZAPEzWLLiJftuXgt4nRJvTceuZ+x7cvoAxhAt9a4OnPHrO8n36Tb1GK
SLcRa4KrNJBRN/1S6ttetG2d+QeO5Giy8b0aER5Zat92Q2dxrfOHhEyuSJet2oK0
IkoVvVD0SPdvE1d8xICeNnIqi8XGFFTe8U853eO/p/NObwzQ4ccsA3vtJMOzCTEw
Cdj3WoaG74b+zy+U7d0s+HIGCHzJUYFYauAXeZxF+AmSGz/ebU5KMzuCuWYb7mOW
8n5s+aWN1ikhI1NifSW9ozWaqZgEIwhKrKQVEnFDP0NnMYPV8SW/8I3pdlvt1n3x
uuae+Ff23w7vUGGnsEc5K8e3E3LTgjwh+vJmRP+b5G3rlP7Nwtm0/tpoGOBSlsYt
IQqKKe6FcHu00YhGSLdocY99IOHXoMpY/8ED8HSPNRzZmKUMG+vgeHTYcSt+3t1K
jpj+5S7mQvFxWINGAqwHWndk7xkcFApnfmweJ6VSIs7rXiq4L1Z8jTa9fddIRx/9
VlcNPR48hsR873GywnEDLkRGcgbtDDF7HH2QuGh5G3w/CzOpjXe+O/4q4FUjSvTj
k8ACNanJ2H/hgOt5tDDCYF3eksqRUM8uGwGYDkhzq5ZfmxKaNxLW2WeaSOZL2Toj
QqVQm2FzapxWDpQTVlZBn6X5ggKoQRutbdthfcy53vXa+MfI9dhpPeXrDL+gbpsX
/nSEbcdchRIGUZ0YY4RurdTurinmUngEz4DlHvHEkM9iZQvt15DAYPyu32Uh/xLz
IshKBhE9+nHvVO1vbJUbz9JZzwTMonXzBmKfJ6qUhfsHyBSqtwP1If1k4p2EC2ME
63WY80cOt5cDCbks0hdOWcdtj0ZVmp8Cdv/Wpg2FqaKN+tVpwnXbJRtu4iSE3iQe
7qyIJ2pq1IjeAGZRneDWsQWmuBCERT2yfHIDffK98WpB/n7Le1q97PaDZVo5HLP5
ubLDsAtsIpthjNzPp5CTYer6kLj8Wkox/Fy5KuV/Ib1uGGzIfdwmgzRwYCWOXIVN
w4NqGuSgOmOVIuMzCx5FKIZ98XfppW8BgnmQpMZGSTAqXIIagiBXSoSRbjmHDAF5
b4MwUJKnZc3hAbFJXcGfMGL6lsvylGxGxeziFmCPyLSuNxwPNKpuCud9QD3mB+vF
UhOxnTVyrxufE5T0ZHvHKRt6ml6Z8oJ5jC2oDRIbr3jcDwX9vwGCxjJc4dWgpc3l
BVlibr7QVJBXyuSPe1Wj5RMwXmqkQgk4ARi49f109sN+uFPVaDqkwsyZxjevUG8O
+uNTtMcVvQaO2LBwT1+nx79njNnI7DRn3nIC2L+ICMTWeFxWQanzvLbTFY8UEdny
rmFOhbVHzSsTmRclx0LnXT2OBCWFgl5+u0RslYiEsmJuNtuFHRyyS79tubC2kN0b
RBshiVcXBDcBjlP9WXl7W7YGl8QZtByM9ZPI2mr3tvxugSpqnFALubniDZFLAhxH
EQVSfAaNcUXOTeqeEB4ZlAtJfD6/ikaZVqpqoyjFv3kmUQlY1W2zWQXfsTATiHSC
2Gf7hZ1IH/W5PXDRuFjwL8J3KhWnFI3b3JFSrYWZBlTowWPL+CYqzTML0i0+DURC
o12qhrO0u/Ji8Ys3YmLiB/98uVymGRIA7gpQ9rSyw6JKtGoep6eAdRokAo5wj/ey
Q29vNx7VgPIPkb0Pvgi856IEHKaOz09mQpxP7YFHjKkuAbk6127VkwW/eu0jBgdC
M0991g9gXkFayjG0GGIobnQ/z40/UQogYGqHIdjbq7bgWQ2SLqEUTb18Ny/i5MrE
cYQ6gOtAOW7H37CywYREHLS+dq+da8hQcmHlrSdabX5LowoxHmW5ktM6Hw6RYhsi
OAW4wmnGEQGFdTgcc6D/eKlL/vlrDUG5AWM8VMu3GNBt9oXao1wnneF9+eHeI5pI
6PYedIhV9guj8zjvJBZL9P+ijBb17AHpsRSpE4PKMmAgQjgrPDIZ9Cf8DpL4J87H
cp3riT8uKDICJ5bWiUtHJ93c9/GqJ6kB0MB9DVSWo7JO0ka2VnAUSn46ACdOb0eU
21xIKlKf2tAtbzFEPGZevCCcbuEvus6cR0NNtBQV9gv9rcgdhlBuhxCLcaAZjwgt
SXDLj1xmJ6q1n2W7AO7mH6t18iGQLTSxk+qQS3gFXsyr0d+KqOrUiJE0LCFv9wAB
r2aBtJFjW1JkBb3c+pCDyhR4Sug4GxxjiDZH00tRlo8w+ZKlIUJc/rGt6MVrGKJs
J7ZAa6/lPJoYcrFpfYnX3i7Qdfp5elgzO+APcPu7epMMqMdI4w0lOOQkRiyzRqcZ
HMZLHhK5l3d1AZNLlwZ4WPMGbfpnga81gKyDqRrCIjK+5rvmcR8nlGzW4/btq2Nn
8ShFwtP+i2SOtuAtSLHK/BlhFvsfuHNxsA2QM7uzPxQ2N6fu0U3SgkbMHAB3611W
xf57lZ7rUvyN6TbJffIm/oDFPMC3WAX2buRGNu0u8FjZGPLvmIwxn0+W9dxrzcS2
nJc48EuNZk2KTwwe7mZidwwHlsxCsmd4jOMfomytillGydndRUQOvMFoh/6VZ/wS
aB1J6azjFmCIfzTMeg36mQ8SNQAOeMj25F+FwnlAjEsOMWQLaZjBiDQkQNIVxCih
pT4bgXOcQWArAgU1i/sQwLkn2P7OjBxVnv+pYrLc/aJYPdJicQeRCmgsxuLnjxwv
GZFYul+s/HPSlrqhtZRYBhURgHXuOodCWu4SkQKQ9PWJ25YbNW9g2rBRVk/2cM45
GWp+80sMhqzf9Omx1ul/qQaTyUmW8iypVEV1ipkPhW/4MK3zc8W8vOZUUQEYl2uj
ILx2vbggjikf+UbeoxIrP/DTQ/q+zXivnVQD8O1cQV5ii7V0sVTIOuxqp0aiB1Gn
Mhq2vjIKOPY6WMXs8tZJ91/6tHsxLI6TKd7GBDuaCIjtaHL9ggwegSeWiCIvvLAi
kJdQal3tas4K4/6tPimDY19m80fMlQm0nC09D8HKOeFjd+VlO8/mAnnzuukeOUBT
UWU2R871y+3RgynYj3w3EvFpffcBmyoOqFM4N4vgBgOgO7+k3AGEvFETcrjFcPBc
cEwDKQl0TxIy1gDhLhKoqD/pl5JzLQqEJgxtdhRN+Y6/3BvgcmsAJOvfJPd7Dr2k
3iMazPE5vGy0T/DMkx7DPl/F8Vj+Si2qGcoA294STu7a402csAmuIBoxUGg6JnSy
Eila1lij0PK14bKmdCicPSdivpNB4eNu/eLLJqPW58UZ852UWjsbzmzh1tImywMf
ONtjqzkWDvUzV+baEJTE0IXgTIIurqDc5UpSRpPyQmmB9LaL1A0r0nOMw5CQAZu7
JixYBUUlGANMywk6OnckfbnefBH3usB1sfnOnARMa2xKSnKRmLQODJcABLOHqX9f
52j1DD+guoeY/gfbnEVquld9+JffbasT8HAYucuUoHToAUz3VKv65uSAvM/im295
QEHYHsvDmbRp43wR2Kz8pgr8mhx2qkkE563+9sGEJTDc6Lf/JjTZzs0nLSBEgrAv
8yOehmqSalBcGMgFoejhfDfBR9ePFDlNDQsEM/Y81IR/Ou8o+NLF1hQnLIiVAB0n
XGjwIZk3HUqPz3EUoisTquTUnK1qanB9INEnYWPS+trwsm12SZFxc01gufl43SY4
UdMO4qRT7aGaWeddgOnQya1OW3wh2vTSOg/rY4RftCzFO06QY1TWN/oChIGv0K5J
fF+faUstzyL3n0/J1FFl4dkvBjL3nF5XH+vyPnED4zf1czFRZRtazvg29mi2oB/7
EkSxORElxkScTjeXGgo5L4KP6+LCnkluSDeGzQ9LyYrSm3tpq7ISe99dtGRlCY8D
vf17lRgmKkMN/ZVk3gCzw+DLuV1kzBbnFB/1y0KvDhBxQDQ5I4lpXKkQPlseUz/B
9JkNb65zk5oKerEzMoREeZTRRZ4K21X+9M2/ejXqC+QsJGQ0/jtusbczRvf8s0wV
xTSUkxVURDbPQ3KJFV909CpoK79b+2Sm1dOor1/v1At3GGlKNQZx4xE9pte7Kawk
N4931q9ANhMc3WrVAVmT1+k2tsfZX8RhA5x5Jh5rFmzwh/S6sKVWFH0q3NISyfpT
Ks/1Qh/Y25cVwFE1AWVjtQF3p+igZEYQVQqYEmh08LDNN7iizSG+PJiqCQjsvN3W
FQ7eVe5uFm4fE9B6gSlzLP/qSLj0GEWGR+SZHewraAdSgpdd9UEpuku8/ZciisL4
ZNzEwKXRr8lyCzqmfB1ZYKZYGDlsRfmKc4bIDMdBolI3ycUNTqpZare9BGsyeDBl
vDTPHoWd0g67HQHjOMSFcpn7T4BUxsbHXt5DqmZDSNrgKL7UiJyv9bk86Ojzo7JR
f/PxXguMnwwiDF7HapKEEGynqNndqSFJ/QP84vNLWGveuXmbl+NfYITlE6Umb3+R
vg0dd7WFD5ypAZpCfWDLynriDD7+xTCCHNAJlllGyX8t9204QRP1vL2hMc6Ai7Wb
LrHgtwfDKpsW1Am5EkCDoVXD8ZqwYVJrifur/fJGeVNLkUJdgdwjWvZsOEHXwVsd
Snoz1O2vGJ9I7I1a8r4WVCqRpOBDkO2uqAL3RF+o2H1LrK3JcU7soM60GvIi9AlW
0sZ4d+YzAoAJH4kgFM1mRxoKHMUcV4VhcwqhZkNgwS+4SgvPNm7SuLoQGuSW7mPZ
KQDS5R9hIbSga04UCmImpIHkNuOaFzVU15m1pxX+lNQAFFFmhKLfWDxH8nUXI1gn
unPeE2fazkRHdozOdjYGmIisU+pbtYr2cOem1kCB4/pUmlV2NjKr2DaKWPQOhNhP
0JzsTTA1GD09xzVK2su81mJZ4n9hy3QCfdr8UJw0IZh8OOJO8riDEpYv9cXEVFKZ
RTICC6lUio/7MLiVTCY+LOUyiVjAEzrnCV77eCmudcIGQlx9mz9uwlJ63KY4/KPz
okSgEThl0a5ZDvOtL3L7YWUpdlxX62Wlv8Xp8y1IRdEVdUIrbFSkHthQA1rAgxRG
a3xI2kx19gABMSBcSKIDPNNTpj2lyuVKnS+ZVIW8awjdIt3t/Cz0H3ERNKNbYrPW
AytaQTo6e96ei+ZpIebyZdD9x+IyZ5O6XwFaNO8jXPyNley3J6UhssALX7CfMZli
3WscArJVHi3p5O0AOy9Rgt8TEWS9IuTxBTmAYEGG/4fMEuVz58iGdlZFrYsK6Z53
o4Ziulg88jcL2/dz5HdhsRQwD0DHbYEZnGN2RhiaSjFw+ziwzXTlRfRuWjtqMmrx
Od+qgqJnESxdzVtoNXld591+O3RruwW2c8Zfb+Rf4lVphw6+9PbGraGbhR32aAFf
vsh44UBH9/rPnIZEsu7k+t2vVYUInBV1kuyvOHt8gDMi+GSmuycbEZJfLW4BWYlK
efDyWyme4LNj5OMVap6ecwgRkxZEqeQbaDtixC3rLtDKiQqZtfIWvj3qBxCAys1S
zclkp2b6OlraYTWmu9w5ymLmlnZg8gtsf7hhMwpEOxxv6uXHOHp3HFLZ0kPn1Tp0
mrf11OOmXxjm6l2KP0RW5dmqbh1ZpBVxdE/SkYQQA5l/BUklW38jxEEZNopkDbu8
39sgofio4U6fYX9pmsXSljTja+C5D2vGNcinfkWNLbODajhSivpcX1wRcs9bze/D
TV+r7RVjvE1g22lCp2haDiRlO2eQfCCl0N4/PyKXo3Hy+Ydr6GqSwj9Sb08wvTN+
Uuhi4X/4Kb+v+6+9BzMs01MobBveVwzOaRjqXwjJKXWMTD50zV4MQ0T8V2Vf2rPf
HPfNJaJUIEgSWw/N6pQNUD4j2ZMQJ2lrCdHXnwTWf5BPnbGQWk0GzwI1ORpn1H4e
m/z3caIScffPi8K7HzKmsHuOd2x7TKbUZxMfPCY4P9X3mLGIMo6n5yxKn8SXw187
rjmfEuxyOYZVPsbqq2MuABbKTwvS6WmI/qETKqwdjD0PbDFqJ5jAQvx5Tu7DYc+n
ZQf2Kyi85TzX4qi9S7DvQYWQUaHNOAOpHUu2DSAVwsvcnQwfbmKvHoLhmvLajUMn
72Uw81WljLKCv26nfgJHyA6TgfTi9YqalOZKykZHElNKZd3GPugYMxFCG9wVjhry
yL0Zm8QwTB29Bzk+/d8xSe+A0Q1ju1m+rqbM9zZTtJ837/tNUFdbEWI3heJ35wew
4TSl+5DlMcST7atOKdXa9mhNVqRJq1sJfgCZ4/uZZ4b1OtHFRcSDme4P0b0tTnjE
LzqSBIpOxQT3ldoGtU27oJWqewzB+pZ/7Ygwiny+d42WfrrRYKTrhcRltOSDkF8i
ANjWJwnyydom+zxPLAn7dgIZMFUiVz2ItQ/Q5WQrY5TEo+ZTtmJep5PUn2xLfGZ6
4Z0gQXCeIll6LVcFt6wbtFXbn2fu2zFRsI29oP8C8gZZlwWCSavB+EJKZ/vzKbqy
Graa4es8+DA2ytmBzpDHmtmYwRLYUT4jbTNXOBkNskb55w2ZidENnQcXha+AtWq3
Bpid7Ic8nfVI9k3eClihxM3UatobjBEhqN7VruJrFOGEhcwlbE2c0oTWfpTAJxrX
mYiN/kkIH0LxvqBhuxhrhh5yeQ0lKT2e1IpzPFa0xqZUQd1mXk1T/YyUi5O6pzdT
1FyGoF68ToMEFYfDcukdOj2c/lRi23epnMvkOvrnZSUvYEvoWLd192Y2qHkXHb7Y
xiNnU41YqfKlUD0v66/iO6dNmg+moHuy+alGwfYqRITlE7RkOplilYJbVX2md5aR
R/epuYacvRcyP5mL2iDG37XpNEg8wpED+skqY2qhcslUxwAQ9Hz8b8IIOH3YA+p5
fbgzZC5q4vdl1PFd8NcLamCTOnMufV8Wrn5vYArJJ4hrmEsU4Y6sf71Zzc9Cu0RK
6g8WbI0M2kqgdZilNMkx3OMPYCjqi+nM6/DxXNEb3+GRxNKKP/QfT+TPUGu1iNMg
OsUI9+vy2UzBgypAQiguH9KKcS+//Dcsn6uf4OAFGzlRnKp8sCiDW2I9jvO61Bxd
WpdZb96lt0Y6q14Tq6sGfRQqnga4L0nLGrGvSxG63MmDggc0oAmCGysIaF2xnn7S
DbsGtF4rmC4DhLhiYZ/wRXsIhICbIc9u+/Pu7hj0gtp7D3FaS/hg8FNSg1z4/SJZ
81UvQylZ3BdOZTrbFAWnPRm7W3x/fvPdu6jnP0A3a7AM7ag+fvbWLa0n83VMfKnC
yX4R8thpBqyi2rctk2DmVUFNdkaN9+zTRcPPVmDQ84gaCLrRkXAsS66WPb/Ok7fl
lo26KK2tsT1YPzJTufF++UpSC9LkE7BGTPC5XQKukHJTrOPn4vvuTWyzPjqhZ+dz
5eoeJHItc+3DpuBqv6b3zU1zccwbVJ7EndqehW8F4TiXERYlT/y2GZrwym78LpzM
hryE1/5WdaXAGFEJyUR7pMaPSXJ4wqVzVNsZ5hShAxAsyC6oeU6EeQaXEdcV+DFy
JgtqHNW3F3IzuIUJYfmZh63a9Afde9a01dqNkTOLJmvwAtAcmaKeWqlYPL8TTe/0
GqhC7jhgVwCZPNKerl4oS4x1+JnL94ycQMxij8/VtjdpEy3gqp1Q1wYp4xwT3oKo
X0FLeAdSGE1aElfwoeVVwgDPF7vRSHRYgNeGBSWJxObFZrrQzC6+rVwHBq6j7v/g
LWCLRyNVAekqK+upeggssTrSxKw7TdOEmTNWA76GIzfA8/7xeOknINwU9wdXXLLA
JEwNbdKZP4m33U5d/H0X+aWgSTm0lFg0muL0tKVobRs2vbLy/vHm+XP5i+vKI3HR
qPn0HNuLbs/dPkmBCL3MOSanP8ki3ZKlnctFxZ2ke862ZqJeOEsSP57Rz5+FrsoT
8cr+Gm+qoTJErfhGr98DRFVoodhOMtO0PRN8Mhfm7ygYuTLLTQagJKcKu+QKUyBB
OaA050gf1qV32JNO4/LJztbCLV3iaex/EEwmsDZAOYqtQ1+7oDkVd5CiihB6gJ0N
QCO+awduOBCtlR2g/5jPzPK8CcHWeqUmtAt8b5FTaMJWQxC0PSjS6C43xHlrw/Jf
Vf3b3zTzqHgPhsSDxPisb8SQqwVF+9Lxk3vAD4xZxkZALrjq8Hs8eSssg3L+jkMf
h8Ghn6oxbUYNBe0TxmOSj3fBo2EzvU29huk3rjbzoB3b9F+QVNmYhv7pvTcX2BUU
o9dc+aBGlJyv98reEdRDGlcE/kTipBoQqv1HiZ9XZpWLIhvs8McUoW7OqBfweyfo
zLkZKUFH8ieemuCZ1mh1IVn8gl8/tZm/b2JTPqY7w60gpe59bOy00S/zoaBU/MGJ
oIE3MYIr6ZdqK7C/WwhCZXsMJzJikKi3mARW3aoUBEt3DaSRFh0yPMgg2plEvaEP
q0znQ67Y7L7h4f/B0FIpsXC1UkK0I1+Xan2jQ7tZKGZ0mSU+pY5m4Ex/vcf94Nz/
psAictxRa87HIynWrdFPY3xknBe0Ej8r59BbiB3HMWoXcfytvBv7vtIxwckQcGO0
lp2C0fT9wqlOujOrivsp6Ak+Tsc7SRS2tpvsDfrqYA0piOoMvTdhkLb1uQdYsMRI
yiCoe/uqTlcI1ygnN8qcHl+Ji3Ofmil4VHLCZRngRohNykXotD3t4D9wbVaT/mSm
zLGoCiXBEMH4H0EgSR5dtv5z8Zmftd0mIXcVwUK8d1rdu1ScDNp59tTbdlyj5s5i
DjAuGEYXonYbR9AIO4nFL2ydZ6Xg75Y0nfU8m0GtYJEGSZ7KmbrcV+6ljKXjpYP5
8BzptEPVUcH0eDZwXBLVfroQeReh8MkoNCGvTlGFCb7WALFmhitDTAD8Cw0rX1nV
KoOlFZzz6JsGCtI6P0MJHCXjQIqWmIu14cMUWRnYXD7i5yf+J87UpCnkPuPqLNtN
V2RLBJElNukP5NMQSWb7J4pVwwfFMhYR51ayA4bOSuJWjhUIuE6OcR1GNtna/6UN
f93l202yaompJ3SYNPkUkoRToZ7nnM0yHvO0lAKckbqJ7C2a+0ifo8V++VvZBPOD
pDXdDV+/mQoMVpjHfDFwv1h4q4jesw+ztd/AvyQGOBfgY7qg6Kyf/pvZMTI8XCZv
PukS7XY44PR6kw6OuyypCBiHBSqzte3YRhzGOSRVXotf0P/MyDJmOPUWiVicxcoh
NFZlH7jNlF6jY4m6qwSfDrItGHklaRASRA0J5z2Dssln6NJ/nrna1NTBtZQ/tVb8
1pVT42Bfk9pLZTpUtWN0FU5t6NhCHIRHEqLxR6GiaId5GLwDVEFKI6bM1qdAvg8W
wIckSOh6DDTXhzKxZjqH9u675gjeetBQDZSgwg2rRwhugRcQGT3MbyJFZaEYLlBQ
uAw7yt20M7EZumMrz/zRjtbz1bUgK6D0yWnjaH7lCPiMiydN2YImeWueDeje2wG0
7SWNZtanZlizQW/uzx9PV0cP3EHdEz/5OsYdL0XI+qQXP0BS81ZwfbhVbD4OUzr1
F7MFfD3PFAYUhqYaYgF06QMB/f3FvGLGaokCDtWzUcfoQQq4nI+Bbmk2LkEhsMGP
8+Zoc6UIsYyh3VPLevWLfJwUJfuv7BAXeP5XvHdpht+n64oao9aldyTRBf/9hV3v
9rIgxNAOK9XtHAlJBap+WGVbiJcJU6gC0vdQyXNQSW/5zewtrD8//0k5RHLM+fyE
tuuPwRbOhsGT7V7BWHmLiKqWDTIYkpdUtpXvIWFIyiRzM22DejKBEtHvnW/kQwAM
9z0V7/bSQnJUkW7WBtWguA67E/mHqVZ364WmUQcQWdcAAhEaoVvmViJQoBaVfmx9
/NvQcTEuxRq64EuBeLq8coX/xe40eByEXHEsD/z6BAJLkt7DGtBJvsodq98nPehh
geEl7L2b4ySQQNkvG/ZvVXythwIqPr0s1vr3tP6A3+ahpI2wOJrZquFgj1ed8y+b
kKsklQzqZwvIiN5vnlYnxPiMZc6yvocjp5Q7BI30zYoMRLJ7eqP0YK7j4jl5KdBq
3SO9oS+Dzd5e6MjQMW4Bz0GO4u/phAgViJMIjmuzsjS+MPfpA96UezytAjGDuwUu
k3TED/L6WXgTv7huZBGZWsdhdwb2/hmQ1kVNCtWTuYvnylo0bXrjB3KipZcTBstQ
3akRyAFTb4FN/SugkV98WWmX/AtrhA8SGz3uMgwTgua4GHY3vI8ZKxUnK30aFxxN
jjTcJYgLS2hhwaAs0A1+rj9ETjX2K5hI1VmDygqOIhaNnFZxnpFW3dgDzVeQqxAr
zJQoWBmZWHnu6iqQgpcrbLBF0OkYZ+ffNjanTLcCPnLEZEsv9SPF1l2cYm5HgrFm
xtsJ7jev5yjHC3Z5JCj8dIsofNVR600jjpgYbGJW16m12LEn+Rt8QJShQolw6zb4
2JiI/3Kivt0EshHUmpWsSyhp9v1SJhizPix9Qx2LBlqt9O3wzb+gMdA+7NkVxMVc
VEkdcDbGDtV/GNyManUW4UZU+PKb9R3O1o8mr4Paq8yOpbnJP9HSvDf6Gn3vMqWa
yrjuBVL1f4zAxorHQuhK05dFw4Ajf38qpYzsEOBCf8NYeqQ3mM8VccMF/BWC57Ym
eV1qad0oGgFgBY7tYaGc+9vcTIxoZC8OdWV8Q4pUxw2QyBww9vMmOI1NojFmm8P/
FPnmOTkWNDhsny9mDrmkN3UMab4jeh62eh9RoGStRIGL0Sm1vsaPUy/U0Pn2/43E
eRV+axrfmPxtUhBStxhWDfJdMl87zLHWezEkbBpAUkiz+x61nzOJPXaTKnDSeHQl
8/S2z5sd9iyU1flA/U81MHdcvcyE9jR76DabUDDbvHqo/DJ0Ry7GCr8bHx/VWP8/
RspHVKHqGqoNlggk+UE9TgEbaWu3Uqmu1l48d8y1J68vLOcnA8bHK5HJv9q/YCU2
la24LWZUWQzYIgLTu0RTejTITsDGzSRs4Wm+ZX7donLwmGZUn1WOEVTsvYBXS+4P
6dy6v4NN5fXsw0q1fy7yR8dOHWjHUqdx/f7gZgVbCASMXOS94SF6ap5JqCAKroYt
I1nr4+gwkkhrzEYUAfy3Jz0ltKKz5Q1ZUqsl9peMfxhSgnFQhKbo49A/BTbXMwD0
D4TzO8AZ73qaMimiuFIsZrbPn87ttvGrLNrGti/wUiDOtcji5L0Z+aQzMJ5Zctg8
Mlzy2UNbXciGW1zkm025U7AuYX2KOUbkDtU4C+x0RkMbHb17b9KoTVpbF7ZDkXRD
iI0R9BLhIjyGBSEvpP2BLjawK++dYBX1kknJGjYTjTs8AEPLhP8q+VZRbiWL/O6j
BqIpJ+rbenf1YKs0wZXAkRn00v20pqU1AuohUqRq2mtOpvnxJYGlgVRMXKSGUsCV
mKFH75WXndoBFK3nitOnGS6exR1c4730ODpYm6QDS0PdoPaOKylu/yVWgYQCcK26
NnJ7lXg0m+7lXaSXEoiyGy/7abdXFEVhzFRvmoGhwfbx0uxunHCNbFBRSx62K6Yd
AQIl9JWpYRg2H3pz0k5dYjxGVUk5ExqH9GGQive3greCEpPklqFJSAl9F7O0bNI5
2DdrxONcOMAxbvmJAPA6qpnfaQYyZTqteEAOzV4XSVnXjXcclp5RipRqtv+LMn0L
nCu3WH+pumTDNmaW2rHnEOtiajjnTY+jgXtNHbhxJiQ8AbhqNeQxete74Mrco9I9
QiKVnkLZU7XnPgwgBFOCL8Bcw8qK0pNu4nq/CCfYa7XRvn5gSlJ8BB/Ff95rjm11
dx7BYgL2H1FvYNJoCHPn40v9tzb3bPMc9WY2tqCVEEsd6ROe/P0Z5cb/InMjeUh3
4y0tag8u7Nw/oPODmlhYU9ufATjG3IizoYK24D+kC87Hh0KvUoMl7NnmwSrwVZUd
wt0YRBtH0yITpNFBpP1i/tLiMGh6WdURj1j+o+G/1Fgz+bKf68MWrjqi4ti7Doth
QaVOOOYGRQfe9AXvZeyTBBmGGiPXPC5mDPTPGkLLENDcfKfjXrIPMJ5E/ZJrTOQs
elHdsT7UqBD0tnKsNb1GglpGXhNCKpzcBE6I/939K9WadUepzJn/568owHpfevpi
c13SVJaZKwmKUgJdG6uUTUd1nYz951WYB6PExjxdv3LRYye2O9FjILP4//MV7FJi
faJI37b1MwvOdT9QX/42VKpRQb2GVDLVM8VBc6o9s8Uwk0WfWn4x1QWsY86o5KZ9
gp5Vq0xZUQ8K4BmxSVCYpuY3J2g8fJaXLuwj6+RZG9eJuXxVRzBtqtbaRTOs2BDW
HxfQtKTZKuCduUggeOjSotC0u+rOLaDtGNHTdiSOzl1mvaqaU8UbmJgnLnRdMcmL
eSkH4Nq8+Y83EvltL/1O+FfUJ4Q/TFOK4eNdijPqobptdJdZMlr33hoXxpB6sqUa
oLdrvyhSIko1x3rYhX9mdcucCU64ja/RGEuUUG/99yjjk2zT9fCA3fuA/UcZ1Oi6
T1RNLMDIdqzGHPfoyHoEswI3tOPD3v/HX/EFp1eYWX+B2YAWKXOipdXttQTfGUmy
7UcklKfdvNSKSVXs6D/3riBUk9bY4Oi0Kx3ZUQpwxHgfs3PkR89hGFcDwiz1N19Y
QPQKAVITXxJLyoEUyHGT2vhFZuIViVYH0RWuUrLHevXXTq6CATMv6GnaaTLTBhCV
K7mUFLDEq27orZIEcNzaTTP6jEnkjdANkhKS3fN+NCWf0sj0WVdLbTS5bDry91+H
kEB9yv2K9VbiVo9eYRjhRac5HOMqsB+n3U6cfFTcP+XOF94xrILzDTriGIh5eRcP
QRleq2dGAFsqsQYdcNIsNivRAgr2Vc/slqUFOSjDWZ84WOsef9Q3vf8TkWBEbafA
KjFYufXseY4rqKqx60gK2gKCR27beCCHyLrRIIcTInddR4YkZms5C9/AktKBBlR2
7l8zWyhiBWR+D/5hyO0QrAvXaQioaySEK0zc3RtKPWzNcCSwk+7J7gK9+xWILOOZ
6RhpYgenIVOvQZfiYZ3CjtdJS3BpZBxBEjXWaVVU3OJR0LKB8t559YpHe2Jhtr3O
jxXc4Sm6ujUKtnby0oNXhVqjD8d/ljcJSvLDiCpxEZY2GQU2OShF+cg8p6dQ3lg8
CoQBYGu4/+wh0mDvKdW1d0C6nmSSQgfrGfA0LcD9IIMAtxHV4eoexzfxa4T/8t9+
zszvMsLIw5weMpD0QyMI/A9DMTPxBhJzht1EkuzOIMZQrQtTnffnX2ia7mWgCiPq
wQlmqZTCIz/riF72UHZ/ueOHSga+TBxcvAKx3mOwTJVZExrHw+aUGiIWVPiIgn40
Q6rpyspf3iAa1OU0Hb4LqNo0nDlPbKDTunSE+6givtxy8b0s0F7ja6htMFyjqIQZ
cHGkcyXviWlMi8yF2fLo1qstLKGGRCdYmuk963y2Oel2F9Vi6FxdQFLa35ZYsui1
opCuSQ9iWns+dNWh5GfsOv33nLa4IOeAXfPw9r7p9GhoQ0kZdJeYvRWgzYViT4Cv
2+UIdir5RAXiV3P1jY0HOgtJjk+r3BW7fapPDxmU7XiUjPLbnTrpryqXfq39HLfA
7h+eh8yn1T53N6oJ+xqPThmmNg6Pmcg6albBLTUgeQhue9PmW2jq3enFF+WBTCFQ
eDUah2p8BmGG2gk8oIfzieN1TfCIHMtkGmLvRg1NN+WKc6LBuaJsvhW4bFoWZ+LE
JbFUJCIUOk2p6qVxTBinjaRjPF5f3T6nYmDFVFTbgpve36c1pwdN3pl147Gh4jeT
B2j1OijProeDw/JNMyvAN/Im0ZywydTyUqokMs+HrLj/WNpAiDZZz7+1QGDRCUZ+
GeEX7Brb870iNXYtYM8OpbSyd9sfW3QznaYdakBrYHcPSb/wwr9iBRWdtXmWHdPQ
XUuTlu0DDJjUjifyvlrU/gl0UOyXXbrOmnP3BA77y2ljUSGRFVW6uj+prIG2y9dT
gCr5kIQv8DXTnNQB7FCEP5+a2T+pbhMX2uaaDoGp59VI+U1VGdfraKpKEJs9RWiR
zbmbmiiIXIuyLdfXWgstYCq5MEzIGKe8VBF59z0G7il7nwZY0M1XU/Pvm5h5s36d
1cEKTIGaDEkqfHLKdxAHkByWH9oZ26BHzM101TJ8mzbIEzTVhhVujO2xjS40WAxL
jXKestyn5eYcUhUXkcJUyiC6QD//cAI0gi9gLxr6UDv7wZoUfNhdHytCWbFswi1q
PLnniSMfjR5NiB2cASosaqIiKMRmqRDIxEzdTv4cdSWL7ZQm2QiSR/Zb/6PNPqCS
KrT8F5O2G9+NBPtBjOr/X23/cDzEN15K5sk1/RKJDx0ckzrwyU7zEL8C0ZC+TDvh
NdMgqhLzOPhvMBeFri31McqB4Sa7mT4zBPjjfCVe0eRfGE+H+PcFVTCqDLplnavX
26To6Bky+mW3IrsXVRLPlqol6FnM3TvLvpP1NziW82uLX/eVW1kv3rcHbK3yqPXx
HCgNpJxQk0lIDgfJHBx3lTERzaOWdoTlsPb+H9GhK0hZoRW14a8g/L6djWXuYIof
+3n1pj0YnnGwnxjvx4L567pgQsoBFQ3rGmRiVF8H4mIFEAVkP8F3KUnJaifEGFUZ
h7L5lMBVkeqKguZnhF3wWMMc2hq0Zs0VTu0IdUtR8zbJ/ArbOHELi/uDWd65rwR+
9PGeSCKSEWspSLPTcpttvgKZpvr8Be71iPNtym2lFWQFHiCZTuU/Jqkp5B4rjCMK
61ZzB1o1X2Dd/+CM2czKzj3i/oBSfxzIQZ1ciRpsjD70iuB9+vF9OuhHoQgCy1Kv
/UAn1mAHiZ1lvQXXy9fc4kRb8VpNyQT1nJAB5U7zjxByQQT5EgPHCs5FEU+8C48/
Ew7LF5OWwpJ4+p8bHdHxEl4ylwS/NGEI7si7UD3njZBI1iWIkNLkzqD4gHJcf9ZT
TRL6tublSFcTJw/NQ3UFRBJWT0Wf49XJM/6CgnGsA7ASCeyWV2G5wNaNwqkSN0ow
eJZKpjiPoXjpd/LwY+CtPBIIVe5AbTuNZAIe/59U1o6V0DhhQANd7l4uHrAYfNut
EVRZ4lQXHOFw8x2IE390FbQaAGEMvWpeAGW5LiwG9ARPcwI5L+wK2HoPxS9aPNW6
ifkO0XXLCCOPW9/1RI6uX2sTk6K4Fj00SDSENO6TYCXLDhSiSRENqlP4e4AgmDKH
15umTD82yFWl2TWWkPwlirMwVbaFq9KCmajIURJ44pta2K0K7ugAK+zMN7aea3uX
yqkOs6sRHN6mZDCicG+ELgW/yCotJB+/n0+8hAnzXyyAOPAk++Y8lXEt5ei9+/H7
LeIMmalXnXUb5RHhBl/QRAeFnrSWUZ63qiVTv2Pfx7fZJS6tNlQ3lH7RuTY9a/fa
LK9Zlm5lYY2lNkQMLbTJp2e0swBf6V9Lmav85V+ee12Lw+uy1KtYcuVwLY+mHIJi
rh3K8gLfHMe6GbXQWBfA19v3oGUSPOqCSU2uv+jFVwOMbQyaQ/2MunFQXhThet8T
uGtX1l+B3TzzHJiNvqFTVf+FxnDG5iqfkGrkpH0ngSDCcfIBRBTmBMmBjGye0IyU
l0G4Qe2QxE7LTpj4b6Izk5Ve5Vz6kflhN3IjF201OQpQDhs6RVDp4u3Q+rjIi8nS
lEPSIhrWuhtyElky0VZRXsnXwlAEA3TAY5ygTjigmHSDrxFndTS7ibxFQCCatMdd
AhyeUOamAMIJYbExXwZxiIuyBssgnoSkwfOkiosg1GswTm6wxMgIc2NFjdKlFvZ0
wfE2VaZaiwmT5XCF1261D0WFnEA4lGSD1VNAT+uPiXXm6Hd+KM9g9Uin3BJqPRFX
r+Pjim3rgikjpC0UiJihtJcg9EOS469AIDzNbRaddeBjkisHuiq0+NIOxMFOMiWZ
i5X0n7P7JwJg9Ng7gv3ETQkN2dnQOEwlW1NwqNZ4J4Wss4yRuAd06zpxe8rKVS1w
77udBKeW4gM2hL5Q7p5IAqbkjaayqSJUWBEAIWy04jGEJrJv3yX0ud7/Kemyf11P
jmwI2K4VvHfZqgFxqvCuAqZjEtPdYb0nE/+a9Gk2URptDNC725PMW7S6PkazgfYE
tXlR77YrZ5xnkuyd4kZJboqdssPC2BsKIVzQMUhV/Gq9Lp1KydDh7PBPuK42/2uC
+UBKL+4xmFpA9UPlmpYRsR3XJwaNfgRFIyKpbVXi+yn+M9F94+ObsRoV3bhywqnS
QpTDmamRe5X1jffnwRoTJYkIA/XmLq9Y7zXeJm89aJPXfI8Bd0rQa7pVBP735C41
PTHVXrUXASxo6atxU58OsXxI+nQp0JxnOLcCa9eIOHhk4JsWhliw9F1yY4JOYvme
jZlG0fcea+00abxEWF9pZX+B5vh4p47AYDA0nZiwiEcqCyC24y79jlXx6aGz09E4
P26oex2K85c7dPn7REA6+NViVkh6smDupPDL3cZMBcC9C8289Qp8X6v7mtnpsA3N
yX35o5HI/fu1/sbWSpoCdteyUHd+J3JOHmBYDWWR/aKdLpzzZSTfBVsQUdBFcqFC
3jAhE+wFrzXaCXjZ3F6VTDqDLsMVoaImMfwIGnJji2oIBtNx4mgyEVnp0gaP9Xvt
iCfHXy6Hx9j/zs/QcmaC3gjJ+8tS1Fznge6Y5Wbxa2VAgV/+rO1CkU5IDwfj9m2D
MPKyVzhz2nHmi7roJt4U6X/XlTCsfijyfzJlaDU6pEOzo/D8rNv4aG9lDb3DacAA
C7R6R8FrSZQ0G+G0ut4pXJNkgtl2YA2y0DgCjc+4zMlHjx6GWYDNS32hBB2DQZKK
TllCueZMisHm2Op9TmwDiQZ2qDfsek0TE2WDe+A8/iRBhX30BLt2aDDpM8yhlRj2
c8hbhM+F3k+bjWDfNQ816wH7JLiD6lL4zhX6SenGan9OGj7Yao5UHhEDmVHiZx/o
J/BAuVAbYHPcXIrCxdKoNKoItzwjuUGi13HywbmijsO3wApaPYnnIglgTEIv6FP2
DrobwglIaTtejoCfyVI5MHWJ8eVbeG1L51TGcSlv0syHvxbdGnXdxY08XDgty80K
cLLPLhkgLjaCtHS7qIhMPoTWefMI4V3hyFne1lAD3VSuE5pxzgg/IHjYZDO5xmch
u6M/6UjoX/qxHXD2VlAehcO84ge4YumEIPjNMDCCOFSuwdxlTvfKUqdwgUhyYJad
GM+Vj8DjSPHC6N03bUuUD+sR7i+y/4VQGsCtIE1ds1NWyf6845Dtn8gaFpMI1TYV
eESJa1aD+EIzRhHUrSWftMtQVoB44y7RmlOaiMfcwUxoGk1FYsLsX28zkflm++ST
+rsGDGXfu1z0epfIaqCVL8jou9i/v9CdWpcEoPdTZ4Z1+V6xBlR2gF2Kq9ebEo8U
8G9GRnzh0n7yoeFNkuMIwrYgzdBLYLhxoqrYq9TAyeBWUltbRpBJmzbJoHaiQYoP
tCyIKNKOr/mQuaWQadZ+S+UWl3NqbNkodPhEZRDdbxRI7tTJ7+hKdaRxfZscshrs
lWBM3/9B5qggmiufZm2qsBg83jyMUHYnPP8IOfxDDjNVBwF6XUMAbS+tDAwZkTVq
64XJoT1MeFp/83QhLW/LHZ8ORe4ZqoRSpqGREJmG6soA84z2s82uqAN4xa5qbgyF
hUdjEWlO7UotujyGyXMiEqKWEkDiV4qN7HVr7coPQf+y5IrH8D9kheBJCvprMYUR
4n46IR/9704OlYIZdOjGutWTgfsc+7tA4ujppDfPeMrlu4P2IkEOobK1AxYw5pWo
7RVzVIrFFSJbKkQ21nqADdYjhLEqb6M1jEZZUxt6RHj/iTs+9FiMERzSOo7ocsLz
SyoFFh28BQV6fxujoOS8FoFnyD644Dw2mXcuJxdf4erUTQxgs8qTrjSUce4o/Lym
xTzUzlREcrzNbdJyL9NIEfaZUZVAoLCaqnGyoUsr24ZbM4/ficuuVSxKQq6qg8iO
tKNuDtuwTQigKoDPV+KfCiYhW3c8jSJpheAT2/6YQCsjwNRYToS4C/U4RSNGQtkL
WoQ3FWLSHZTGHRFaDBGG1a2Q1AKFv8/zzH9hM2HVnJtAjHu/6Mb1HP1w8aMK7kzI
hQZUfTYMCCmcDHE6Li55+phqP3WUL0WyKBHkKZO7hiC6lIktN48hU7yGLaKMtt9H
f3rISNemkH5gVeGMvMBboWgnRZWkEi/0mlC79AiSnXBiBpfwoLJryKPAzb7XI9p9
YMvYugI04jui0jBgXKud/SVt/5r9itJXnaQYPTne/OnKZrTb6YneawtjRSiYVmEo
YRyBt0jvl/Y5wiuFhRRCzkvE0xEeYj3xtEql3Ysdr8ce2lu5LWSxIIDc1YKy/lc4
f5TpRvehn7rlvHhrxlqCFCjQh9zaBLLGZ5S7omvfpDuQEgi9xakwvWpxZT+gy1VX
PnLZtHiA0qeqit4b0+VSf9vIDuDrPhpKT8YNmJ3tbQN01DyKj/XjElfzmV0FIyvQ
+EquC00TTnfRHTn1Xfs7GRPf7FYe4jZfPoX5ndML1uRuiZHFncQOcUKyAb4ygZ9m
z8zv337qeEDHuJNXYiof/sHQNijf0OGm0qK60v+QkZTnqcnw+QisfS+ehI48LJq7
8YRNxDhap3Z4yCfKNaDr1WYYmq0gvKWSyJxOm4iCl7hTzkEe8yU5VuKAYasVQxk9
ZgOhsj2/rL0NHPjY7oKDhutolqomyeGUQ+diI4gqXWjP0LA56Txc+HM7kBnz/UKR
D2Vdzum7e5CQHtUYGd4dMINgcSB+oMrNYmy0lyg7Tc85+xhKYQmPM9ktEEOirjXX
vqP5GuxKUM5WI8Zhbvftu4gtJhQqEl/r82SakNR24lLgxZEl1dKfRaE7KX1Khiqw
9bkR844sTDSUdSp7kLbnYIXSa7szayyU48juiMtsvAOkZk5J0lSAYJxPW6kse5Kh
NgKrNtQmPgva+4ohN/68LSBbKhjbfd4860iCre0fyAPnN5syEU1ciBhCBYaAGrx2
t/NlIErXpdZqhGAD+237rg+6gNRhFbpOKqS6g2bZshIuOPGy65ijiAK+3mYkGWJW
KphoXx4+Jv5wS1a/nUVZDqxF0GEb8T6HBG0WGvzZbe12F/pH+Nc5Gq3TyHdW3swy
9HbrzRcUNn2CyNSnEZHj6Q8HvHU8QcyxTV6Do8K2Z03NFn+U1D6WyX7C5nxtzXp7
32lDW50xl8CYt++GKK+4/yIhwzzKQFPAavL9ghPBVpcGClU+PxHXn6qj1ORc1Der
CCitJSgyxxFKXKhN185VLqEvSZ7xmW/Lk+LPuAKRZEAxld+vKSkIs8aU2D3AnCVn
PMt48RYJI+nKvVEPCSn3wjeanXGaBPfL8HVVvUA5ovd/BP9Wzi+aTIhMQcsMdYpT
qwyNmlYdAMeMcfIi1AuMsZprJe4gaOD+7rcRgKZ58SN8WrNfVzqOt6+bjUpDu9Hl
51rUGFaehouWxIbqXZ1KBDBvTiS/sw7TwFhDr6YjaLxnf+0j5PXb17/tTI0l5Iwq
35eyWDN8EKk+hoUyA2LM/JWYaENaZS2YIstNKYcz5PpCL5VwOn1GjmD0DFPm6wMn
vwakK8ERERPZPuQ4AT2lNlodMczPyUTX2mKeRYp/j3gIh8RztG7fuhdPZNsQEteu
91b45Qjv0cpgTBxLV9M+J5HnfXuR/vUh3vuz1JD/oKbuiU2lqMGWkNGm74R5OKIJ
4HPbO2eVlAYxs1/Z8VTVW4CYrw6ZPGkNdz7kQhWTKz4vkkVdKf/SrddZy1fNHAmK
caZDj8hcprXuJWRCNGLTPEGK32JCLMSvqPFHMMvaJtywBmO6knWhG4xFn/wV6JE6
5v6iVmxAVIpGY6og1wzNMmIcxmcS35E9yCZWL0iAmaEbmdkWzsxJlZoo/Q2NQDyV
Rbb4pjAKoVEjq0qwxSaFzgwsYEdt9LSjJvNNLCMN7A/naUhaaiqwQPt5WgYRLVvs
udg0vm/A8IpfLxRUFwfX29sUS0IG5a/1v3869piTmWFIMIbn/NPTkzve7Bbk+xRQ
oHYSVYMoLUyUSpbwHLj5mnju5U9DTWlNmRtJybTyXfkm65W26RdZdPPcF3en5QXl
r65wnQANnOF/+3ghgyRzxDcZaAz3mA1HV1aOyz696a0h0r1nl1Wc49QvSQ5qOGdl
O3Mx2ejKOnJo2GaRkxDWoq/trGtF8GWeQ2MY8PolkzSwx1CWmcXNlxbDdaxW/jK5
/N+Zu/ewa0noSlLzRwpXgdnNjvZhYrZuk80fQpLoS5bea4BXeL9WRwWqmVIbGZVM
nzmO4FgcnRYa7Nuv0qypOKIWXoGKHFzVWLhbzpDFUOJu3oRc9IA2qxuDk24TUDQr
2Ar0ZibOlIuZaDcRBPOa1TviPFdNk7vHz79hGpR1LeysfL+Sn5cr7vaAXKcgb2re
VBAOSnU5sk0XgCirItsujwn33YFJKctHLxQruIna2aMjRQB2gczbmCxxNmpjZWk3
+V9oGoClCs/ovrk9xApuJDJ9V+YFHMyTvNcCqKsd4GYWBoViJSxVcL7pYmrVaaRy
OJpcIgMe+6kLY/UM17LVTWxv3T+XUohrzcbzA75rv0pKiU6PSYbnuf0/A6BKmmYH
DHJ6GnGTuHMTj+Fvaspmuz2/NNp+Wx43k9sqFfcKgJN3C9/7YCzTkuJ/nHRaaU4C
o84zn/EzlL2xeX20Xub3vWyQ67WLVTgSmBpWiQAfitU2CBt19i9VADHKY6MMVWz0
id5V0WV5s7RIyiwvPb3QyvP4BlkEgIh0Zlg4W8pG2JW73FLOicHsf8ApDBmGk+c5
wbN8ntr4GV6XPyK5th+TMTEEELeMEK1i/1mvZpuHImqgM0L8WAWkxi25NeiXRJDA
gE7ifB5OFL4MCk/K4yya4GccRI8hNFA6WqX1skpzMSHTbeAYxpOW5GkgUkkIs8MU
6fuEJ08bbronyysedZQyKw99nksepUXkgyKVUDRLz86zbFbttha8preo85L0PYtg
Rs9upQlFckPlJvMKTM5AaD8OhcHbd4vjN4kI0+oPuqQ4Q0XUu8hAEWeFzfZAqtV4
DvfPyCWDAhYWtxf30Qpy8IxFbJNaxpUSOmzCjabswJomZ81bg7CeyEntCkSODb7n
5JcpM2NsVY2DvU5G9kRGpOZoZc1CIZlb64wfnkoiGvf+7ANG3tuElNulGCKpOSpu
+BVCMg6t/TEnqbWDwep+LaX7xu2e2SIeRHpvxjtr8/cOYwyjnZzCPv7Jdm8E5rql
/6FIW9c194B8sLkNh5x60gYQFNr0nNkebOpwe5n/oAPI5n+EfWqnfFM/fVBPq/vB
vh7tYm62A4uj7VOEG+HEalULKETB+GlrQpCvjgnScfbXdChxo0BwzcWjJykXsILG
+AiHTc+CF5h8aEDybZTKxuvXmwJrQ/oxx/eHUIMs7/UlAvXZlVagt22s1cxuIvWU
1JZ8Kav4viOZ5rkYgJjV44pH71PGvpqeRJbb+5v4l40wroAMIbLV1PrnTb+bvUVa
XZwBWapwB6lzhghZ3vzsK89VcmoEDw9e8PDmPymu2kM2zfcDRnKJlHRgMBcXcfBj
h79NFT33ApIw1ofIZXzzAblwbwfNnGVGs0+W8ZIMRe7YP7qoBEfz4HudVu1bL5pF
4kpoDukbaJf3B70Jou2B/CjLw5tDhkejPLitf/HPjQlIlc+KpZQwyZRjxn2JhtPg
w/xhOeZCcfyFmf3Miz9iFioIXdFhH3lpdRmt0eHXTmOhGkQHlTXJxnMf08QGa8+7
bLPP27ZyM8uWlc6BFq0GmUMzptLfQbbSd8YQKHO6vScyRNOR2JbKV0qs/zBvKTQX
/T0/EWpMkW1gp94sAV3QqQwkQpbKEdyHq2v5mNifF0pBEKN0yGwvXxxD+wYZk3QG
2pQAcNfOyt4tJuGvFDM29NT+99JixfuLneX1HhmrrV0aXa9gpst05wvmN0088nya
ZWEjJOoEP+f14lfpNbm+OnBkTqd1eLnHZvvdpV7/5dsKrF67467V7ZKT9cgFYeby
QdPK+m1q/nONsFT51lYC3Fv/rmCufZRCNUEzqSuHnsvdQYWkfT8VZbFNckFsNEmF
wf1n9onHyvKoTvicJtw25iXSpEfAhj8E45l7zivivOqyLbfdpifQrHOTSmb0zNH/
/5Jnfn55v/h5HjAOdANYse7N1jbwLApFxm6OUn5L9+LcXyBlaMkeCjUyEdLqzC77
NjyEKUpCSZq/+CTyvJOUHe8cDF2GAEMjZhOHZ2a0VS9v3x1aZ75+qPQo5Rpb6MqH
AdI9/zVUKlZmLm7E4gHC3RBu/4IQMVsqaDg76ONtJTZCkp9T+o3DVRyozyZpI+Bc
2+pGwLRB4/e0YYk2qiTOl8Dg5Yj76+ggtFytQJAj6BbFzn8F2O7mcNB9p/SKNrWg
eOzJaFKxdPEYmII6Ea01sUUtxK+RRLtoKyGmX9Rhdr9YKuOPzIbG6GdACrqbI5JJ
Rf5RQ5ohHoaRD2kF/vHCse7RgKxoBfMV0E6a3Q8jAspDvXw3MZqZk/eWjwsXN9NC
3Da9+mDJWr6DzGCpMBJlUG5pqieqPzFMrw94O/Fv12PRwiHsOVZGibYDiBSIN/cc
EUJSkkQQ0rWGQ0afJnx5VBYZ4pvsWa7C/BGiZaP0hQoZ2JP2MV+1ci1X4Debx/sJ
MCDzgc+MqP3qNrRLR9x9aHoqepxidbrzczxjBOW0qStM4n4yh1inpwG/Mtuo2oa1
K3gjNGcoz3LA9G9p6jPbGCXfhXp+zA8/uwFdFcAgXuYJaVma8o4pUV8f9OJvBByb
oMMv0VUZtmLuuHJejtPaEe3njB/REwKOnUtMXjwwSuhrUSl4UwTzQtqTyXQh8kzk
zuiawWpd+MQX4rpkqHz400Q46ttE4jdfyseGXDgu9n09cKJ5hdtFpfTX/QuKu5vJ
D+5lcW7ROC3v7Ms2mghvdJy9AZXtz8wK3C0gvIw68EjMMqkRpV1trVy7fCpDCYSk
/qG54NTMoAysQszEXuq+kZOuCGGnaGzYairwGwfVYmn9wKac3VIVPKJFu7qqoyng
QtbuNJeoyeVKD9uGLQNf6d38SUIMFths0Rbigf2/sMjMVNZQmudp5Svvn/yp5L/k
Y0dF7MpgW/akAdSy7Uvx8wKumCHhGPnqXk4P8yNq9N+/E7M3Uz+ps/ksECpC0Yyc
6Wg0FGhAH0tXSKiTnN3hW97CcqEZ9dkwn/deuvsz2P9ubFbTlTWdvJwOH9hTiUAK
imNFc1GSaT6tf2M/LFgMR8wzVWH3Wv19RsW4aov4MwAop22luWl6fDlbPBjUICK4
gQa2TN/gpkGkXwUjHXGV46dA6qL8ZiPDOirQus/0A20Z3s0i6XzdFV6TMrh6ELF2
Wi2ezff6xS5InA/y73fEfctMN4zW+5nohQ9FPlDmjbtICqhq7IrSvRXOgKPleE90
+OyCmSg0+b4UiWGE5aU1Km5qnmskyRrBpbBbnnrORUrJhnR4VUajFjMHpQz9s3uo
PqRpQsd+mT7Kfq9VIJ6YJlvI9koqDTWOwUaYf3sltim1MmxC8UPFtUArxwL+aHD8
zdvrhrwfr7sVNdFsPnza+x4h8naNJYVFGQ/DUeq9YbUNnUyhDrSdRa2ZSi3KWRWg
Kxs34I/L9wQF3je9NyKZEdpxdeLKwUkwFbRCaQr22O9Tsdwk/8fnKXlYILdc5bRK
gd7QpT/Zke9y1RdUxpa0zQzJFbaGSie22TovxWSy5otqgreMTU6vW5ggmzJ+G3Zs
eBxM11sNhs+pcaUH4n6Ven7r9BZIdx+k2CS3uLJMN3bpqOUq/ik0joQrYVM9Nv+J
PqoPv11MSwb6jWOUy1E1V8W113/IRT4RnGneGlv8mdmnKrO1XdcwSWxFhUldRkcG
dlbED3r6T/cvBar4tRs96tRg2YxrfxyH6PwmVBj/8kkQOa4G6Etd+zQ+yKJ+UFNz
Hmb+NRAxZ9tieSR48vKEq1sBXyqn7FTrkoWAQ8u3iZHdsSAoRoZr2L1fjtpHaPgf
sXhExL5e7h2QoTsvxrqe1y7pKsYuYnpWqA2L2gMu63V7w+dcCdav4604hj49KbdL
uHA+ln3DW+L48cnQN0Eq8aUjFUHwWyhQmO81Ws/goMMrfdwYbPq0ZhlQhWUAir6b
LReaAsCPBIbE6SiR0CmcgFP4c6GSt6gGnDnY4jXdvA2g9Ias+PiqgFyQ+RRlKrZ3
AllRj1QoIoYkyc21GC79FLaX0nv0rJstz30QVs4y4QBAWNb8I98GZGMWCrYLOUhf
aI6WIttDVLHPWS4izbQ7T1LXp1OxMpY8o1p/mDYB1YdL81XmTDi+qGwz0rPw6wB+
baMDlfrSUsD27kmCydGcszeeRImVgrll+jWPIf5JNX1OJo36nIaMcniQYMvqSWSG
prt2QPd0DDq5VQVoXLv55I2K4rm689100lkc71Sj2CaWmEHC+k9lrWAZA5g0ymjg
JO254idjtTVQcxgU+024pnlaHhFQFCN8MpFGlFO+u1PXPpO9fRko4gFtBD7Fqq+S
2wFuQgZnq+upUP+LqWfKjVQR++bptd2iGXIddryqs4C4UiLZqkhWVApEG3fzYbRj
sSFHxuS4twmHYoMfNb7FtaDyZHhRH5emOEBwf9bWMomIRkVfJ7bcqyee5+1TBhI2
PFb1e+7ixIxtCUK1d1LlBIGwDFVkLvfrwpJOrg/z8nj2lzpA+MaATvtW7BCx1hfV
zW8SzsXfoSwX3ZqY6FFUrlF3sr+XClPLR4FHeMOrzqjJwimZ0RdRcaa3HWwp1k0b
vysyazq9Rn33ptoxSycJMu92OSMS/FLryw9UMMIxF8apxFM6vLswCLONw6x+GPU2
zPQ1EoyG4avZu0xDNl9tZ/7kow3wkOVAn2w5VQ14Eo+YtJ/hQkzOYtxTKU1h3CFn
P1uCHvE8PRDHV3eJjfV3xSXdOQpv4pPzJ97yBcNGmAARFf3roA/wPybTZTt2mAsK
fKPzETxJz05y6RIM2FHdOgyFP1lWHDzba9UO6uW9sBEJz5uSjwYdAy3q6s8PWINM
JY1xSe9N8U3iZNSqXPpQzzEYQjW6SJhGzvYmo1Wj6TRrsxEwk/KAifoYH1dCZVXW
mASMqy8TExw6RjzlqFDPr/kOliRmiSOpK7uEHJhW5Gm6uYoeXDCIeSqXy0m9dp1G
MaqQbLtyVBZLWSlMz7ct3Chgmryeh59FhbpJEZZxOjiqVP2RDjs+ztzrRExYnHGY
rAVj/WgC/Q4HbebMV1nu7jLM9VvzKoHxbznyj2JdAWZDxdr2BVqRbu2ykwnqm/RQ
Ww+1mWtCVDy58vYr3jjdvoj0yqk63PnBmKT2huNCgHa9Gr6R9pUB9BQjh4o7+nby
TEatS2JtXCdPSkD/J27t5ynnVJlDlK820qfESSQwk5zsKRuH7w4dlDpc7YwjPQ/z
4Mft07SHBsclsyRJGH3u1ZUh/3neNaEhYQoe5Ay1sg4eXqWSlUzjfz8yzWKfko0g
ZO4Jm/330mnczghxb4hQYwXST/KlrYx4xMkssTWHekXOj31Lc2qyUcgMxNTzwVxI
Xnys4o7j8k1SYgrkniwzVzVDNkNjQfsDgZKsKi4jm+4GWc9pDqr/pJgWf8MvNGAa
f6dlJCztJjHzxOr3qlvMnxPInoVAUuElSQJ6D3LRklPQoqT7a1XBqq9ga463o9n4
5nBmrcdc/0aSP1PH0tT4D4zA5hcGhzW3IdV0bpMwSvPeMXr+vz+W5Rf8dW5RiTAh
MyinyilHyf1uUh5t3Ff/WZq4sUFEgQxjMl7Y2LVatj2foZrT1T1Ha+t9skyHiV8h
NbdeVEuVSTRF9KBrhuPmbTmoeFDO8ZQMXiWYjStKVnFYdunrDRgNe8W4TLwn2utA
U/qCeXq4gHCufnPmkd+OpSkoe7JGnpfUyNTNNnwW3+Y6uDfpep3e07r35g6wwgJK
bZCt/rt4sxCltNS2qyiWVufnC8BMBhEMEnoW7YPMmGCjAZ+D5aPilGGe/eAoHq/z
7Thf7ObDyw/EtWPcnoiItgfkX5jG/XGVvwbW+pJ07KZazj8SwDpMeHs+SHiJPlc8
jGq4BR/bLO0krnV/9clr560+Zj4BnwtYVJMXUY+eJTeI190/EqmnXPCWTWM/Mqvx
HZ8YeEBlHc6u+HyfBGp0jDVgEr6QkounZbmQ0Cnci65JlLdSsvJjDGDPs/NiqIUL
YDcm7t2w4fR5by/uU1neTBS+59EeIo0vdDw3b3bhkOtLm12byfLvZptLJWN/6wR9
j5zmTS07reG8ym6lQY4lVPQQhJbruDdb3P0Mj8RvGL2Ku4ZNNF680/FjpCwUdOzS
QFdnSjcXm5QIliJmLEUayue9xTqJo8WEr7Jc9aQWXheYY3sDWadJN67i1aWItPsN
CGALZssWtZFNEWrbnBghVw06OljLq1BFiqVzHBu1ihSZOa1Y1W1NrKFS9twGXMpW
oc9wZlzcdGvb2UBxV+g9/i75yn+gcyZjhNJId8ZZ17m5mTLEivyS939D6DrhWA3b
IMdXfg+ic/+7gn4G2IXvSqSlSTu0ns3DKjeCw8TRxMpBXipzXZQZz3QBbaP5FMQ5
X3M2nCWoDr8l9z9XEb626UlYC7ZrvMOyWxjwkT3sJDry0RSOWf9sCeXEkTZiLVz0
/cCGQoiA71nRtDIAdUY0LYSm7A33jL1jTbO5g8x7cU0ku/zS0DnjN9dFVvMSz8Yy
fh9NJ1zLhlBr24HbdYlVbEnCjdNi4Q1O3hp3D9kZuwhXKqgbUiKmpuaf9VhhoZH7
rrIWXeCbuCwb++bD/vasV5DYqhwgvYpwTR8xcphouxfulCArg6g7yjKSAxz7SVRj
FPt5Z3F69f3XkbWyN+fKOGnv8oTKNikCvb2WgZoYedmZEkaCwblBx4lnJ2ua0Gvt
VafO9Eb/hipZ65A+pFkoMHZUjHWX+tWA7fctqCH4ADyKHgrnOio6445zF4wBaOEN
E7pHLOjnzORdkqI4uC8Sz4eOPm8cj7H0b6FoNSR0Y+eDOjGROHPxk7C+kf9zp69G
gwJdNWwZ94MnowwRbkiN/fY66XGo++RSI98Cx+/MA/GRuu6dXb62x5GBlaFMyEEG
Q/PBDdubpbOlokTG+20BdinxgPc3Tcu7ouq1kC9XRmX8HjXOM46imNWY0ApKXYv+
UpIJjYqWD8XrScjvBsRglxEfzfFJgPtr4iz+b2t+NE8wf0ZZbTSdawjnbjr/o9TA
Z0xKe2j1/cHwn4PGIAOX64uJib0/MOZRuQXA+OByb7G6Oo0je/9c9A+goBsXvM6o
7B2bJMlj1PhxRxOjp0qYq8jHI+RnFLG9HCymUrT2oEG22uVY25ZpuOpAJjbAMGFE
Lsv/Msgh7zCuNwI0jv0zjFXb8xFdGRPEJjKgjqp2JGB9QHP7rHr70nwqtRDtl9A6
c9sECEZ4RYEigle6X5LJKmsAodkCdZBVF3VJvWC/5HgGfZvGclYxLwsemIsvp9TV
1yp/k/49XzsMTT/Cc5H+ooHzLnesoOZwVs8i4zKfAQCCrfQjgx0tgOTHBDBOjo3k
V/ciWep7Q+d7auWXlFxqM6RhyoGGYiMxV0sz8nlVWB3zuqUOtELwjW7BvRAJYX6O
XqtztzARGtCrp0I44u/pXr39TlPmKPc8oSEkQXj/U3JcoohNijyMDB8OXNpRJkxR
my5Bdj7NhcFLRaGF79MXOhfUzMdhiLPLIPW9eX42RwkJZBlLu+18BT3PBdaRebmK
3XubJgW+i4kz0t16Ohb5a13/+YSkVtc089AqVY42ACr92hur5Xfs261+byn2C5B8
pXnhjNUlb3zLcvxHSty792n5Yxwt+NyZWqDWcDmmn7znaiEwUiNX29MXHWMXTxII
36HzOt99sGOPEQiBow+tNxqiDgNHaQzBHOrMfxxurP9PcxwWSjRMi0a5v/VIsvP9
aalvUK3hEQNeNf1j0b8MP82PLgLIDgrxDVM2Druaz7ALMXdUHxcWCGQoB2jWas9l
EGJGcxWSMsSNItAMGf21Q3np0KVmMps5K2JuuodoWg7g3u7klk9/3OY4XCLjle1p
zJj41nWJ5ZMDXuANDBkQMOnX7zJzSPG5dXgJW8O0FoTRK6DNVI/uQYkQL+PMhmlY
L5yLR8X3SoNuNjHYYv3b0lb5UcFMwmxqMaIVPGUbL64INRipQvbYzqWV31x0PEHj
nrtPNFiDZTPLAqhQg+0GtBX7W7c/iGs+X4+yVRMhRa63LKonDNqDI4p9ElJ7ZVFt
MF2O2101uARHq98et809AoYbMeIXSvp25rTyLIRDu8cZcJIBqeSzkEh9iQB5JinE
pYqS0K7MDuo2N5X/ZcL+J+nIldxvKFiDvynJqKQFNJare7EwneRhIrJXuberznIX
kYzT1XG90xY9Vrs433KsbUJFTJAiVZ8XjdxngeBeDXwwTiYrKz8FN6u76m2tbSMk
aRIqMzmS/Ii8AwZmwePKXKOjHALHCcvD524uVVp5rObRhK+y0DjGXa2VEGRNmh7x
jyEXSr5hNgZ803TqrS9gWOzKBdoitF862qOLix53mDKr2Lum7aOqDxW7aK4pgj8n
qdo/35ySiiQ7RJWvIu5YVsOPomb/13LKq1npPQ0KBa6CgUsqhNE988MwPHaQWaec
qCcwnblGzMFysVzt7QfU1jxPfEMoDgeEKFQPyalC5KjuWzyLIKGmExtvKVWE1uEM
Y7dluoNAOf79HYXb4gUAzwUhMWn1KB3sLNu1rSrSMQYQK13TKMRhsLzqWoPci7jI
ZEYxRsobub5HFPd7cAmzLTgSc9rKpcKyd5UosphfgSb8+ruKKgK8LBmwJg6LsxIU
7obCvZoL0aNukTWUEE1r9WLaEp0mRNYiYhM6olzOHSJwLZ8rADbRMUDwLMRRIRUP
McPJC30BSnkDARDOK8UZgLJgsnsYz5G2XtfLWDz7LlrpKEFbtYtB0LeETfhWP1nG
rv8TmadcincCgcVVEB+bKXpvA/RQXRcDPJocOGsqyvaR3EbwBRJvTotL8EGBlkUw
qEuYP1BZ6Mg0RNKDJu6cyqwH0zhXmE0RMz3882ANY7eSWQ9hM8H0vl1Fuz/MrtFX
qyXQBetnHGQFIKaue0fyKW+5gBfp1De7YzWBXub1TOZMVXgF2f4k9ZOQgF8sYnUR
SDkIfpcCpfsmDFJTjZ0hT5pOlkyTZt+JtDC+8D84B6+j0GV/glYOdm3jo1EGuMos
K5MtI5DboToHbR4Xjxl+nVULyY86sD+1kKa/eTbFEljpPpIA0t/oZAu0fQCFgPPc
3imG2NsAJGGE8Tonyoej+0gihBMnVkJsPpSPXdHpJWRUktV7AaxeJoenh+MGdxQL
6oX4rU/m/K2T4fwNWOxQ9ZncWgIFuaULHHsiaRjKTYAFL4p7jVkgJ6hwng0MBHaz
cU+FMNrMAVIn37FzMxteDtBwWPscIgzteZBtQWR6/+T+G7BWGiu3hSUAmriDR0E0
moWJph/4SY0KletMg/8+7bUgm0B1MEtrfQ71qAkzYDNFDpyXDuDOYA6SHpiPzbhm
lZeasnAmc9BQFBdAspkeGa1+1bJjmZKEjiahNVx/QqYVN7x9mRq+0LF3yIuB+NGe
7Q2zQYRb84ANVO2AX7AZIugshCik+ZpsbsVQQzWpjUS/vXfJ6emGd9VpqTYofgQV
TtauOey8y3dBA54wDUNl8cv8u9GZ41A7nicxwwzSAK+PreFKv9GC0pljuCIyB9IW
yf8OuaDkzi53JhaPBHhO4QvfHNq7LYr/VXrl6qIIRDTqco5qywoGq7BagIdC0ZoT
4le3qX9eIxdJF77F59ufoXxOubzoMaqbFXoUBlGiNGZ9tiLKPQvcy+68bNXLwXvb
IneqzNTX8RvZlCzYjTiB7EBip1f4bmmnfKDsRxdG7xYXi86ewFSfI8G6BkL9vwW6
8m4hR11yVUad5Qij8Eiuqu5qqxWMuby+3EXEP3+S1LWGRDLUstVRHKGtUOImkmQq
3i7hc1Wqe2LCCni+S5y3pvQrOeRrfqsWWWInwveSrk7dVGPYM9PbSLjZZEXoj+jc
7h42wShOndob1S8/bHvKou2v9IEMs9PhPn8W9D4oPyl3kB9nqiRj2scKsSPLwcur
5PilEZAAao5ymoAbBJuWf+8Xyp1x3A5yqzGY9kIE18FRn+NB0KWxoLbySf9gZWjt
2sWedIcutlWlAsHGjxplyIv2ftIJkMM5Lnpeyn/We+fYWp//NZsEKuRYwN4f+xjN
3eH4LfigqRDocTu5BH07thGz3qvMyRm0qMhKASwviyg9wIF/XloOMtakNODdoLJe
8jzxcTvRv9guLKFHVKGic3gGBy38iWL6CEZ1b3hQe8kcjeDyxZc+OqGN8nQ7aT5d
vAsDDeSmMqscf21LQRoNBd9aAdouVXYbx+B2+RQhIO1psCnI9mMOSciKdFP3CMlm
WXhBWDNeW/Kev3m+ySrxqRPcQ4CrztUaNlLtLSzmn9eZln0pm+xYyYhdDssUINyJ
XS226Vy+LghheaBcdJ5HZHYQSIeCOGzXcUyniJloczNUNgnchHzlpA9jHBy3BbgG
IbIg5GgBncvvmGATJUetFJD0XR7ACKD9C3C7EUIgMuBA/DVLFn/e2dkPZXRdbL3G
eA9NGraDbw4AlrieUsa6Oi7aH39Zx6zASFuDC8VNAZ1PMVEydKieT0pyRLxUo2ca
75zHFrNsnXU7c6vytdjf51xPOD724HM9woKR/VrZmdt0iqTo1Mlek15Txy/aSHpd
qMLhxfeLJbmYgSGs7AB0w8m+dwHzMvblUMYwNtTDuctz05FAuaH5qtmwy5RDbp90
sQ/zIxK7ScFJhfJvLgjM6gFbQf4UCu1ssHZs6YYmvULD8stoOxsID1xXm6G5/6Iy
se4RvucWhxuTBBpgBV5E46CwKkQI5V0yTdQ9As5iKqoPQ5ZvRsBugaD0Rki9B9xB
HGgCypcEbL13ZUoJBIpCmnD/oBd5Art8NWnPLK+P3fUYp0bmzlvYwrA/Cv1+spI7
L/o38abXw5pwetdMoyA/oVyf0mXVpmEzvhuoPYtZeloVwZDHi5MwhvH+BJL0QSiw
tSw4qB50/ktZ0Kqb7B0fF7LUmmW+89lWBAJp6EkGrs3x88/mZO1mXojSD35l4NYY
HpE3rq+12HyHThMXqSG99Hs+LH6P21waymtKLIeHtlypMS3u5hZUfe74LC9iYcCN
SIWdiqqlXYZpkWMon4uW6DfkTTF1eG7DGsyeu0MU2qasKNJtu1MC+5d8cyM7khsw
SfpxmSp/T37UQKWAYko6HE+gdgMCVMVH4rrz8rCkxDi+qQX2cj5+DB92w2wdNWEz
CY53lztUZO2CGiKoFxbr+oNksJeAvQJVaC2M5tf0pET8ZKME4Q/yknSS1fPpKraJ
9EqNUQGVbbVf5BAu4vzo/u6z0OOFunHyNRrJ7DtwR03Q+6NsZglKrAfnf2f4mr2p
xl1wH9dXMGw37d2legZWDsG5KDB08LMZ6mbvVc1GbV3vC3dGGRoYOfHQZk7ecy+u
yR8Q3ePlWdCBk8ExJfDXW9pvmLS7+ujASN/5OBsxqRtZ3UcPtnCEPjYyeUUgYj3a
1AqjxrOVQOV84KIvf+MFmn/wfmymcxGn9MfA2br4B0iLqiTg0Xnib/zqk3yBQUmy
DqeEXttjHaCIpUSALjMl8WPXtkJQvC4vfHaKf+IIVW6CVxRmgOIdDMB5WIXVNfEA
JjuMBpgU8H8Vi00fbjroGMYxLuQqvpkUCpYDKsn72bVY2DkrWOfgwQ1DqPw9Ivb6
3H9uvwUb+X1JlnoXbPNUw912uVNW5jWCNCtXdmWQRrpWKvJumnFN5E+if+P0/Szi
pIzCVqRfZg4aessrNIzz+y8TxLUIODA2muaaTxMSbNtsUMVrY2GJTp4Atc+HYYtb
Pv9eBRyvuWMJKC9arzibIsfW/TS5y5q71oylb/zSypv2rfbdY4jhJCTRJbQDRWJ4
XxOU/82u+eGl/e5HLHckm6QyJM4nmS9WnAsHODWvuuLk5lH2NFC9UwdWwMXtfYsk
rV3FQMCCgzWum1qOtkut9KoXRXi5r5K17qRdI+hqmrY4iKrQxH3MY/v7yJuk2kSV
9nYisFAslgAUVtidGkkchKlBVLnl457u9W8sHe/qFqNraenqDx482qIK8RcrY31F
h4wYeSNGnrPf5rhaXkiundy0r9ps5Q1jT/xYi0l1lrf8ND4En1FoPtwutrm3dJo7
6szyF954B9Uwf4r3PYoVSZri/zBIEy+iOfmb5u+GXkSiboaNiTgASQIq1Tmdib7h
t6M9idnZxhSSIO5AixayoI8IM/+IBYC0T5vbreGFUJGTTKB7fpfrwlMPvQOLbpbt
+x7EVXqvdr8nEobt32gZRWFs/uCoGdYbRMwj1fxVr++57EzkhDq4iXIeMwAN3bIX
VDefaX9QWnkhWDVxM2kJWk6GfSccY4yw2XKqDNkbeeGxCb/RjeP70TUiXZGlA0Ed
ZNtooupWQ+zz9sA88hKK9a+waQ0PMDVKfGhPRo+d1LoPibWzQ16EFx5G/YwrEZ1V
HZywtYZc7gKzuHrunwJi0BEGnWJKiSgH1gpzNxvOrRpeHqyfPnVTIW/Bo0P3ArQn
W5Irrk8uUDAM+J32L4rQ+t4UnSJrsMUh+Z8u/4M1SHHHkADHhm+W6274ssMhAFmL
O+YGkQMNErLZqKh0GQibTDfvlSCUQOURrYpse5xUeBgQwV0ahZcLyA03KGAMX7JG
Dn5IrvhVtmssSJL0P/W3zRjxZjjWAzK1ykrZXY7WHy4ubrvo3jVrlQ1legOFbJGv
wvbEiGD0U4ZkN7O40mX8mCs+RSojRz1ElCWwao+dg8fDjwjNSdmSboN6l8EvP2mD
9GjPPAb+0i24TzJbFcOS+dCJjjD7y2t5/OhoAVQQ/JhjIhth/Cv0z64YFsaL39gl
O/mBaQ6yFqJbIm4CO86sODU5EfXsfIGzRDR1Oss7yOt/lcsbNgDIz3+D3TYpwe0p
2WJoPDu1gBY7T3s/gOxIwPRjfZ6bqk8tzPZIJ9ZGRYXl8mnLrczWaJUYbQ5r/RRh
dYCIPIhcNajqXErMDj8j31BggZMLiP87cA73BFldRcNS0vBPTvN7W0duYmF6M1rZ
ZTcqAGQ6CZ7s1g4W7KsRlJJBsVj9GT7N519NV5y7Gy+cy4+OCiETrixeVhrguxJP
IfPDlHAv9mvNRbDXFwk3yozKLoK29Mb4sz1oKVtJ5WJwG+hJS4iHFOvaANTU01Wc
jSPcKMln/noGvUD+YnQU90XYjZoArqe0ni7Q1ClUjvqWIKG3B98ufe/N8YOw13oX
zpKNXFxU4Zf/mVlCPJsCUDy/8p32BQX9RH1BW232KvCjC2YmFsU/KZeBcgKT2qet
kCqJpaJ35whrarfkLCx2HkltdiybTg8YkR4F4v2YauzjpIdaWiCVR9GVuT8zXniU
yjwoTokM5v/rJDTWVWWsTG2U4F49S7hbNOlpsaYnKf3HkYF2bRI38sBI6tHym0ke
YkmzGsTeHkLyS3li7EizC1y7RMeFoVi4LFTkXBUOGgkzjuPVXmaNHl2ED83vHnPD
czU37GMCurvg72PCyiTL+3zIok3olzPJsImmaDIin/8pVVRVS0cOks/O4uVPiG3H
1AJXRSbP1KQFZLikjr1wJKMVEVmKog9YweaBPhdG9R96g5IRy7gfE+mMwalscp15
CZXlRK0F40uE4wVnL2edbldn+XW1OleeD3Ckne11LrTjS35KL05Vl3z5/EdCENTD
xYedxmBNHwrkcJQocUv/hDRt1sDWoZF0qFA4a+GaOreDQ6EO+TG7oPM5121qKd1u
Vcf3ySDvvdNUBvhmKBd+qKq0eQPiWDVvr5uHRWQ7/mehNSyMapztNdyDz0zOMaT/
ogQPvJ1xelAazDT4RhcdOEZSUNa8DxcvOwdhUdXKfs8RzKU4nlfXHD4yumhYzMeS
IaZrFkF0mF6dqrbMhVZCra2dPDZtXalziEvFEN0vVx7V0fVtiyCRDHQJlhWQJqZU
HKvN4X/p/DqmyYk2aPH6qysGr+aCADLYWTFhMpvsmUW0iHF5WHCM9Ol0d8/QSWaW
fV5bvb759rwUF4NQ8kf6XDz2ttMkalR5Gpw0Ao8mS0A4L0TbpBf/ZTBD/vnNQygS
PknXoSbSGfzEybe8Ci8Z39AAlZL/mmZV3EiiXiZJ42QpxYkUDg5MCMvllGUvOPWs
oW7IxsV9c0zZ94egbGBRyvKtpXV90Z9UEgLcI8WtpP9Q3D4Y4uWBCTe+PcIiVkN0
uIi5U/D3CLrB9hY62VkCmfTzjbyuSIrmyVs/psF5rKPk0VLy0mX6hiGH08uNrQN4
A5Zl76tlEqZOIC4+BheKsGLiKYnYByTzJsymq6JN52SPN+d3UurX1yAj9XkGPWYu
NBcYwZph+1T8s33OYLoQxPlgoJh4LbLjD7HDYde93nSBKVYphWkG2iuc9UBnDgaz
2mME3QWdxfCZnyjD2BxpGReXWCm+aGpP0ymq1pzZE1O3ar9CmyehQl4zvzLYz+/p
MDPh6/xCpvsS4Ux8GZnHnw2Ph6qwgw6CBmaQ3f061NgXrPWy3Zf7ae0V+Q0T8TN4
9tf49ryciOZfyrE6sd5mhgNU+VODsyDuIIeFePv/smJoKRV/ZQVssW2xmSO1QHCN
OnbbegbYM+fRAvJOvFUdqLt1pPxqdLf3hAAAaPw7a5uhLtsRzWTavhwr4DiyKN/A
4G+Db3DNCIqhaJUoeAFyRxC7r4iqpyLjNJhpBRXSg9pcOi3GksTbRd45LJp2Gbcs
MTl/SbTWJncRHpJ6JOme97eVR2bJyDq6ueal4+9nRbgLsTU3A6WeP/UZ+Gfj9rt4
ilfkjTp1o8OL8ifuztmiotDX3LgM5of85/lRg7bxHm3wUrpkun0coCllOX1Umomx
O+slyR8I36Kn3ysdznPlQqJS0YnbYFldgY0ptANW/LtXV4rWATsE/3wBS2zks1ci
o9f35qKSXAlUEkFW40wrdm/segToqCasdLLcqxmfgb4F+0hs6k6Oei/0TjtTjaGG
yUxdRtxI1/QZbTUQa9PE6LtXIsn2hLnvGdCOiOSG9Z1gbCG83vLIwbndD3aJJ1u8
pVU25TDCRncoE3nhLoQOZ5sp8+NxDij4KVof0KoUiknQVPTjEia0MwwllNF+5YES
97yeAgY8QhrIvSpY5aZ4MSoJth9h+dE4uNo+0bkbixAuU/5tTw5ZtWCrIL3m+Ae7
/mVOG4UAwW2gRy8in/8j3ScotlzewWGcngSQdpWqChELCTuVHUmi8Wd5xYvOqHNw
lqdEW6MlXVRTfj2LMxluqLM+C84ymu5YLPznjPgJ0Jt4PR2MDcyMcnzlwr71DJu6
AGmuq5xBWvjeCWgZCD8tuyy1wfAARxL0JQd5NoaGzOok/bpL6+21rVTWxjRO4+hC
ZDMismOcnBptZrANuTxilpID+Qk2Fk0bgHofSi/cqK4IneNpAcmvvD15wDnCAZ8l
dLDSDCrOmA4A9owkniYPtfTjk5Z16yQwKrQEDMQy2JMLV+IoCyLfMJbw6Hrz6UdA
YR4MXN2nxYdgu/Jsgvd04Co8mEVAimw2BvrB9vqrCyHjYHnZYTRV+E+Io0EX7KhK
1eGJovt+TzNUrOw3SGOq8c3jD0TvTSlF6PeTQO7x+uSWCDjyeb4tvOy7+TMf613v
s6XagBpL1SdPzmroU+S7sVD1+a5D9DkiH/M6brwrRbF1jk4BenUKC1asz2cExg9b
bKottamTDcE9C0BOoWI2hVjg2kLB0hEPXuXgLEs7tGMr9EcGYG7tIlQDxXInkAtF
8ebndTTGwhJTLn+tGhoZfd5t8v28dXtIngOxDELv9soGaa2Jmi9rH3TXQyi+fVkw
lIX5caOOHpJ5NZmRfo7b0At1keYTiiwXY832UHghky+ETpctNZ0GxUAmprn6lLpG
iM9TCNXHApMrga+mthtXZ1YWDnhcSDECe0JXTt9oK3Ea+iYagMour5VxUms7dEPS
RnLOLRt5e8oj+cLKIfa4i+/ElUP3PPuamX04ZDIsgo12OBnk5zLBk6gGTIwXTn7Z
veqTV7ymH+O9IANLeGEzdUfJGEi3CcKUjtdsw+sRuvWysixvixW/JEsUAVjvlOif
iqkwstg6kQY5bgJYrYc04hJxbsw1rdqR+Txi3WxV+o+3Zj85H3hfs88eHNqTmTD7
TghOw6lpfSfsKvz8AMjsjhr1ILwEcs/7IQxa4td95aewftSYypXvwNaKZIWo8t0J
2zF986Rs4/fEzvz0upwZsu+65SYeQzgUy/shDBIy/9vUtlHfAIdNd8MijQhJRn1v
eDvOeXbXO+i7wPu8K5Nm1uldutKySetiSEcBAnKP0uft8GoHaXUFAgRGAymPr8g8
gDNO/da3mvfgctDqdFmlhWPdMlkvVJdHEBNj5P40iixPpJq5Fq0DXKmd3Lyyg8Rq
J1PHtaTJ3ULXahOfUkHdiX3/nXe3V5Rfi9aPmXCfIDpX0v/BPNUxsEr27YRtJGQL
PWMfhwh3kzmxnPBA0wh1WEmX0G3pqToJNsTRSVbv/PWP8mxiFPlUoMAs8CPz8H3D
C9EOgBNaQa5EsurJ2LBR7y5XZ0tdmt+bAc7OtJO7UGMKXyzWhhZrayD02/9Nnio+
a89zZ/DYPQSdghQVAicvc2BCirTN32tqIFBFQCc6Z0rYAXv5kzOsLetxPg630uW2
S7ROk7Qj8dRHhB4FXfPXZi5lgxGDO0Qu4D7qZhRB1ieq1OYb8LjE27DFzPzBi/Ml
1WT1BP/whx6IV2XUHWeYiaW9rP3Fb4IxPi+pGdpQGYMPaCFDbZmgWzXgyu9yvJtz
Oa6cdPrBmc2PHoAd2ff8rHH5UOGHJsEOw1QAtBdKbxmwn2NIKsQDXbXKRHzghb+Z
jK6g3M3MDAGRksLzjLUW6qL9Nu6exlaVRSiyxn4l9OuTANCB1RXnz5GzvVfxq3bB
OsAlfV6cllm1PAkDkgW7s5vmzq7vf+wUpSpeF6RStQno4oNjh6r6HXOBpdlBZhnl
vB168lqBneguGS3YFL1N5NugqePcjGAwLtcpDxBJRv9Wg1X/Ig6LCIJAODD9fF/z
VvjkGbbwzh1LVaVg1lOfEulxdQKXieE2d0yOnzdoawNZ0BofUjY8C23DTuqMUr6G
bXwNy2PLE52HpXg4zVRM/LR54j+S3DM94i8OkyuCVmOEHtjrYs4dIrjUGNTlB0WO
VdpffYHgnYYahb2JQx/Typyrsbe3c/b2u3p+iDtrLtwALwApyEvtskOo5qFwZU9j
PQvlleRR/+2wgaKaM+1c1NmUF1rD15/zgvGFPlAaVYkP+APWdqvgxYTAo74PQcm5
guaRCcBmIodZ5rYxKvo704NJeGA0il0TBiXl0p5IOL+3H7iSYy4ZqrviBb5VGaow
iVY5EmA1+rBObSkpxsdwajJcslrBRTVOzLcW5WjHKwMEe8kpB4lWGG1kODjmgQIy
vYH0xcKFFexTYY82NYuyvj4xNBPKKjlOr5AcFEQ6miy9SEZn1pObLA6UllMnLJDp
XdOPt9kwZ/hhbvWyPQ/ji30UncwIpMAaO6xzlxXMlhGLqfExz7YdXeNtT0FzcW6B
7v9JOxem/eisY/uv/hEygaHi8JqPDcU5QOLG0qR1EzuemAtVjcLz+I837nGZgPqV
fMvhTe4Bret96VVyZUHXFK8MEAxvGgZuNaLSyegKqxSG7Lmm3ewQrZrkE3aiLgRR
Stq4CpSHJiHz7heJCcKgmUDMQX5SAsETtHvt790VZT4P7YVqfobJ4ZQJmgibYxcx
tMUkjwdN4o04OOUW6j9q6udy2P8rsxNodw337pZC22EayGDNbNdY/6+blQ+nu+2K
iEYO/qC3+Ty8tazf31UgW4RdW/5+2oZ0PzqCm0sAYYJNMLYm1vlf93H7kGgXpz9R
vZxmeERAQtjdBRvr5hkkxGD2gImv4RUvOUDT3eWeRU91Rf7UDKNbnStn8AYrglfc
suEGVzFf5Gwx7BW1PnWsjvEAxdw4aR9ffW1R9mA51tn8aXhs5qOVlAV45fy9ZOk9
BRj+0j62t9CPnzh6sjNBOBlzabFnlrfXzYntGfOnpGbupsSpH6hHfoM9wzJ46EbR
8pgBJyA94SIbYljZHZhxhXl7x+KXxOL+gjbQSjb7uhsAZ1eyQAdmYZOltGcTJGPa
gMMcGzY5PyZav0hfaHOAf5ZEE5qf029uVrckms1wzkvm0sEp+nJsW6lBODKt0OyK
t2Ezfjs7+kLxoc7F5vECFYMSXKGdRSO8rVvtPDkGJod0ABffbIsUczJ7Z1HeY0tX
5qBNEw4BOpooX5lwtD/2+CSEoYtHTqHh5J9IDi/vxO5bBYZippYLt8qCKYCpoGjk
glFRnB8uLCeNVjrhBi41kLCBey/FOuJ5tiFAJc43ooL9pgBzHaQYKJDwjqVNrSX7
TKsPfsMEFyc5F7NzUWFbIiYJLtBa8l3uZqIHp/ogJj5CJzzzQFUDKWT9rsMPTeMQ
L9XRNO5EfEvAY7xSJP5bbEEqcES9861fQKPmljEJ1SQlYQVZlJwuS3mAbyt1i3M8
XGNCgzKNAuBtR0qQV9rT3qfT0HdM2/72O1NC/MhibVP5V5zNH8tg+p07mfojhX/V
D5Vh0Mj5sjT09KebmIYztuhGNyNr4p92Z0qpdOAdjpm3XI6UnOU4IgawX2v7GeSG
iaJjLVVlVJVfQIKpLtQsU52OoTZsfoUjHyKqluG1rtqRPTWxG1Rs+8sRcl1QEAa3
x1hY85u1Vpdi9As3xMoJuJV6nd2iFc84uczC9Qfmk5+k+dPJIpOP1cu2S3SPXGjT
jxcmausfJNYwUp0kekQM+D9bn09gnwxm2ZxMOXquUOZ1JLGyThE6MfFwsgapVUCx
A8rF5D4A70w11uikwEeNy3cnjkJ6JCWa5VrMrfGVk7ewGl0mg0uDyHDdW0fDxmCV
M1iXxD75THmk2F/aLCHUYDnyNOZEHZtTByihpUFTctyswdW5HRa9k8RWVdenbB37
CM4X5sGVBOs6QYR0ipavfY0x5KWJqEw2aCXmtePFOgU+nJFulDKA0vbpSg29YwPg
mOkVVtnmWaBqrxbfaanXKKWEKZpmzNfvd/E6mtEjpo/GcYkU/gBmRu9RfXCInwJv
8KSo5HeAAqRf/vRx1sX5k22VjZJykSObeUfU8jXQqjZtwXKnBH1oCEToErpyLEk3
zKITctOhFaGomXjdYrVkz/s35Y+Qfhl2xBENT6k2x1UYPLBrLhvK6KAu50zJWkGj
k5Os54GhfH2GdKHVqFxTtQQj7nGECH/RufQOzNpgM7Kv9diC9+EfNpNIZD+6/K3r
eMN4cmiV8tyw/NRIe/V209r+BWpAc2xjXghikXtqad8OhZBLt5jU2jnqidzL9wNI
oRrei/7KqE+GaLzrnrNnqJZ9Yw5C/06gTeZygVTdvh3kIU2cUXXSbe9gqSxFpdGF
JDjrYjJLizZGaampGdp2hKrSlUt0a/iK0UpkCEvDpZ6bw4HfGVWU7O8rKPTRREhc
L4uPWgSJVxE+J0+EUF5fliE3fadv+jXwMH2nq/8ZP3sZk9Qs1NYaatxvdZ28F/U7
fnddEFb/FzdbdoKCOv/iiSxTTiOT8feNuVK1FPBHDgaq2XSb9oa+p415sPd7/13G
ONTsoUU0fNSouW1QnejmXE6WzYEeEP+AB8j/pCKBB6a0gf3w0ufMes5lG/4hYc2P
9vCGlciBUy3mLuS07iBF0gyOXVhxCX8szONanOyRQXjjD9HwlHmuerrxCn5hRDOB
ZlW7q5dVyxFMf+5Gh8zVCR3TVkevTAydwaJHxtZ4PQKiuW7ViS8cT88aQIqQJb9L
g6XArI3OVBs1fHqJMNbC7TxrcF8LvcRYfzvHasUgrWJkNcREhTzn6TSo7RUp186r
ALlTm4bGdFgGKRz3vC/LRT/gLu9kNFKYhGf6xBhgQ7xq8vUsark+GCGcgVRzgAwE
y6O3CKoES+AQV+zSoGxoGaVXmh0s9F/s7eMUwh4XsIuHMX5IkfP1QtrmefvPpqr4
N+g2x2Ozymm1NF8fTJ5euF25OFBPYTjVUB3ubRY+EUiVw23hmnjrctBtyTP7BsUm
uGf9k0vCdk+B0CufTsLZpDwfhI9bu+qJYeSYGuYjftZEfAFQ5Ae5YOW7tXFcI1eh
1YEXEzYBTrhyWCYS5mNHwZWLcxDiUwU5lxReiQUGxFaO+ZLs7ly/wC09LvGGbeKL
ggUc6IKVSWBhKlKrhujySQpQthUlfIfbsqKCj1iOWdDzs6vq8eGnL5Q5xEZyBTpa
mdA6TziyM8Gg6l3cLc0ZtS0oT86TXAXcdgSWhba7s6ySJH9vc5H3cuHnY1R73pGi
ufziPM/A7+Gnv7dLvV2kR5Vn0AdElckQLNoMIsrXmZJy/on2x2bf0cA02k/8Aal9
MjU5E5nZO5jfPQlirGApG3M6OiPq3Ia7vlcXEMt7XVmjDqvywMcdDvbGa/xHRFmE
+C551AfwSzOlMIDL28U2vbwE3vuJiFg7x5/rxHCC+1le7cTkCD3GXItCj3cc0IdW
1thjw6oXiTkt8TVmU1Sn96Y76xmSJtplw9t1bs84s4s94NC3kTIS0djjQkd0ju22
gqUr3flPy3ohQY6/GO+nONFmy2QRZnqC5cnXYNKkTSkTfxIfToTL7gphDKTSUlGJ
ELE4pKQUuJOPeyucDFjEsR4c36SrliN9DTvzaWdIB2ftV4jHZk/kDSznK/XNYGGV
tjot8BkaJrFgo+0rXP7DS0TuHTJzTV+SqmJLjPZn4GwanFe8HsnCIMk13O2KRQtV
Zr5ATZLN1Km5/fPNgXzYEW5J/hHtwJV86UHhrhB7PhWU8AE38aSETYovgS8UKIFP
Iv7VEgKC5NXOkwASnm+O00MseBFglICD5QGNBxjU/d8Ul7qpMaLagEjMHUMYznIf
PEZXe12GeIBSpkYo+D96bA8EIGLhQY2OTA55xw/Dvh1e9ntNUR2EpSbdSTgjso1+
KX+UqH2WUqD8PrpYqi0wQ3j/cfZQ2ecM397Dw7J1HhpiYIUEQqIikjuxG5a72YoU
jwyal7LDlQXlcml3lfP+/nT+d2lfUNqIfG2TU0JKFC73JO49BJ3IR8IhP1Mi+UjH
G0p6YpWqEqBsx6/yIx+DbBG/YLy/Ni1t6DqvDfJQ23fhs8FyqRCE03MUIDeO7mNC
gCes7VvwDw9U6jVFT5aNBOsXbfcgQRKSr0lhRAPeHk9Kwv+th4lAoHcw42ty9UOX
uqV06j+vc5AVlz+P2fxw6DhGNMK56UP+CGLIiHrMV8+WvsfocCzr+u1Dx6MFCLyp
toLr/wmiHrNHYwiR+YAMs27NKuFqd5abKsH3XXuEWavhWv0ywbEB41wl9pVTMxWY
y7Z5Npx15r8iFqDRoiwP5NGpXD1ynZ/V89fqTv6HsqyXAWRqTs8GjiJ/+rDeXRrM
HMXTKvJZvuOgukDLjYijy6XKTaNH7dyRI2AnvxezmikjfVxLFqAgHF83ejJDz6By
O2D/Y8JwUdZgNsJGf1ipPySSdlJ+VwsoJjvbjrJzDG7XMwATv0w96XeMWM57tl/t
Os5CXgB++NPTAFWXfy4rER6/CIUUoRSBKw71McGRYJokzkEtA5U3BEUgTfAscITa
Yh4oioPqOo3bvctqiBrFuYOxHR4Y/l5tnLzYPPjShwtw3gXMlOUmW/9rQ9LRRafu
Bj/Bag02iUtDaNZ6ip3GgRNBDjbMLr2QSa4jBHKx0dy6SEEqvquB1J6I/uuYb4fe
WJvI7pvTZR9NpEty/IUIGzyxZ7lzm8pIIOyaPWO3Ogq2jMJ+jKDkij191K5tGnV4
gBcRNFxOYe1CkqSnYNMYAQwjt4lTn9/49SV3sbKLCYLq8J9CUbp3FLSeDUjRpT0S
LdPzB0r2QbrqosPoqegYgmp3lKZdP2PivelMRIJaApJ+GBPmmnIsIcQf/PLvxDdX
1Zf+CQgLXk9d7x2z11HyHbfbQjbqI+PiV2l+1N8Nz/zWrmMGyPniFeYSE0qp+Aak
TvoJZ4fkScHlIZ9Zv1ucb4t+ZjOKjMTmRcZQyJpnt0LBhi19fst3HNs542Q3Qgkt
8MpYwbuFmwiJvgs0uLkeH3smet652SctRzA+q4Iz3x+tcOhfqzbs4jOVGWUJjCBr
LdPOYF2mp1ufUi1gY7MVj9+TDMn4sokahhqmg/XUhwK3LR5ZiFa355jx+ZhrTuCW
vyn60VCv4/9nDBIImaYff/wHUofp8HLdB0m6yZxNjMEQIipv3X1k+Vu6XIzVaPMu
ADf1NLsmr7Mfx0gWQz1HlpGgOlUq7bZ8AB7qBl6lJHNZri4DzIxNPJyGn8RFk1cU
SMr57LPuzoP3RRphORyuttrSO4Aw1RDJ55D3TTTXRAVPHJDdrjBS4rIYrADeT43y
h9yJlmVRzikVxW3AZLiyQ0Q9396lHzepIu7kPL3XGKhvJ6qgk3csLUezyoPR0wAF
4v8SItwJrhZlMfE+9a2AdbsLQ7h/l1NIa8gwdNgY9q0aZx+K+7uPCTM7ikFzKK1e
pJ8tWIF8GtT6IWrOKqHLhZiBe6k5614LCw282k0/I59wWdE+0CcumCQFA9w68zO6
gMem9O+6HUw7ysZR+N70a4aAOVXh8sv8BCznhvEZZFTlNAua9SkRaa2+t822J826
fp5poM54BnbYiinr/zkYrVo5KbPh/GeBynq4Ao3UhmSbhd8Mf+bTmLT36wtm7KSb
tC/6O8qrWkgiUwv+euhtgc2ztCBH7RDTJLob82wf8Kxf/9HU4xTYdu0xlBQ/I35f
KFYhhk8OvG9AsRSJPYFWwyWxiicAf5ncuu5YU/9gUqh9jdCHpCxcv4/nS9vJvikC
vUMMA7wUH513NzjN5O7oH9+QnUMI6Em0OogxmdGQtHGYQ2036FQZqo62YpPmk93f
8nkq7HiTvDF37LHan7A6I2B+8mHD9IDU/LhQAlULbs50LUlYnB9RAsgLKdelJHuR
WyUpFGzKswFX3IiePbblEvhckkJjMkpyshtHzyF3i8fAby2Bkij3DH9NgbXIElr9
Izrjrze+35YXzKZZOadj55xkenx90XpgP9AWItAta7sz9Vc6sJl2hZkHr9BHvJkV
kJHyrNztuZB6jvCORgSLn6G58UnmFKWbdG3KveneBPXBhASZyNiXFBjare0puDnU
c5jlE2wlpfZQ8AqxbAyr4MJ1StpE1mu0LrFf4Xw4QnSCbbKMkfp3lztKu5hHPtXU
gVN5C2xRnjQFxD5anKPYeyWf4QquR4jZk1QJzvXa4qi6KwKOiqBIpBYbDSM2Svx5
pM5TlHQCDFJStttFouTE6PL0N/Dg2qwsGZxSY+hRXpxqBClOnFEkoF21BakvCKkk
3bDBDcetdDXIZqZBg8qSkeUM8dJn47WZt5H5mWxePZ7lnn95U2i8c+YSf1bXGnpW
9EY+XMmqCO5stviBshjH6tMWiB/R6GrejTTjjsCutW+FrrhxPWeRO9LFZyq4qLBE
HFXfsE8Qhn7/wLp89imtIPGwW3mykIE6FW7El5ZT0Yu7sh5fnHVzKcRvgWf5dJ6p
oPt7w86KLSXPIGfb8wyZo5yN34oSZhzWhqdmASPHwlT5/qk3NvSI02inDCwbw+Gy
yIE+agGGonqW8NvJeMih37aytB3qRc9Yd8e29KyqbG19iVzp2XVzsMdPvKhk7xZh
FhHMv3R2RtKc+/JCb/HFoWef650Ww+7mNIKFlo9nEUcFLkTbokAaOErA3cPUIAfz
0Qu34+VAS+ZDhQ40D91MGEqd+D+s7ZcrRVEsOLpOJBmHdINbLz3tAYSmFufkD+Nd
F8DJV5hQFtlBZV/sISw12rPuAZ+DkP/A3wVu/YpbXlNuX1dY8GwuK8y2r+ecE7B1
rnGBQJ11DfOSV494dCRAuZZya8iAWY67Z9+YhpWmsQSz5Ob+wXHA8A4hIQT+AURy
8GlvefI6dPJDJtqnTef6CE5d3KuNU1mStddzqcBcWmEHlWPUwJWep/2pFwuyL1o2
QixITDloKmu2KvxS4hA4Y1Qp64wvGPq8pM74b6KsIXDXwX3Tw4UgeICGYt5u44Jk
5/oXWY3ywWADqu/sq0LNtUHF2NMNcqUZn4icTX6/nvADfJ2NO6S8hODtVi0bHDqg
pnMr1THhlatVmuuPxuAaL396RWLzzT3wbE+t0E1zLIFwlQLO9vq/cNR99pPdfhgZ
FZWKciif1HfTdx2sTKVD2OWsfoTx6gAqUhGLrb/N9NvoWdisGY7pPF5CupENFxoO
PHgRdWrt/FCPLJRyEaIzuUIFBrwN25Pz86/l0jBBXU1UgTOyjgCAMSbzcEnUADOI
p7b2OZICwbi50F5x1dQeJ9qWRX3fIAowf5jodfmHaeAjIURXzMtjiyVMQr9wprjk
BYPfuCC+YhQj2EQhhwXLCl8virRzUlo4fTNkYOznyAgtMv9SdxNVwtF0lMZQVEkJ
0xEQcaoKe6Wm+QoWL6X09J66I/mbABiFuyGUZTZDysF8RQeFdtwnWIrQ3oBPDgZS
LGS6exxGgRcG7ec8ZoSkgplCDRaS/nPyzN7KECLw69Lgda/z/uNxDWMJesf1XFwE
oLOMzJAWX8r8BWD5Hh5NQH63VkI5f77rZ/snZuL7+JK5X4pdRr8PWu/96BoY2XFK
Tb2Q+2IHIa79p0DvFaiDOMi25zU5gjG54P/UIiVBzK3LmC83wctPy+XTUxx0ln3e
/mhI4BAUuoSgNkgWo9cscSnIXiT4b24Dr5X9rZWxZe/UScyB0zUlfiZKIVCyHF1r
3OGkAS7r8YeEFSJQSoQ0RVeMb8/2OeiWqpu22qeKeqEMF0QuFjFvfKbmnkJkEltX
40NF/AWMxLXvytm4w4LzPKLUbmMBTx+66fAp5F8pPl1Nx4kYpucs5qkYrCGvRtzm
giI9FP2joCVKDO/0q1GpZlF+afVMjLPQyHc9vTbAhTPce0aJZPjYC5RXV8CL+X1s
e3F++qW7yf84ykkd1duc1CiAhaVIyqIrD4ENUAQYd3Pwm+LmJaG0TU47hKaecfHf
KxaYKjjJItXuomg/1008riG0Uo+dSdecZE714piHtIeJKou6TmJKW4lQK4TqaiOF
FijSNo7s6RPwJivJj/tAoO1mvIZyRyAhSz2rSIeOx0JDwaBpaBVtCLXSAm239Lb4
qnEuaABaYlIDt6cDu4pfVmPETHNwyuF2sBLv7jdsG22AACDzZsJ4nFTVk0OO5H4I
1pzi1wWhIVaOAvKv8fGivbZ8oJHDwS5lxDCi85WDAZQTYjaxAcHqj4PGqQtIcw01
yTTQwgKgTbPg+w/P7YhUrNgRchLxz6STCPdKkauecfF5QUL5ZjB5+F/j61ACT8bE
LwcT08381vDbOLVFnOyxmMj+sJYW0OMYVkG8Us9it5i/guIAIqFtkyaSaDptqt1t
4nmRcPkvKu/O8dKQc68lHakyOFLZ0yhfF7tfqH86m6e8f5Wdn3ph6Yw9ZUoGfgWw
L+KetmsmaijU26cTQslT3lxK3oSMBNRNB7YpDBYZPi57GbOipfk3V9vxX9OJ7VE9
252LVHcMt22HKsHbVFK/EVJQETkhT5PxHa9R2zV/hpEPI50OiDzcAV9w+M0uM09N
PquiJlllPntMOf8BdjKuhfNnuiVaKrsL95vGFszzsPEwNXw6qSSm6GvcbkokUmFp
HuCzz5wCLSSJikHIt5QRwO2y6kn+tSXuZbzRN1KfAcLdc9EkV6feByac5sCvWhbv
j12QnUYc1d7ZP7sBb2yHD9dQ3c507GVNaPo79fZN7yYAkW1XWLmo8r68ZoWVW6QW
JXQtPj9GKwPpngvzFqa7mnzksZwCt05/qK958Vr/iKqHJASmTAoc2NzPD3myqykk
Byvz6Kgfw7xAT8PZhL593SbnKW3mJW1fCaISWWKga6prwpGCE+hUpfkImq6VkGxb
zAzyJsJZenfJU7oRrcA2FUM4ZxwaW0wJuj5W615ABJ+zeq47Kqf9VCj60SaJjddA
hwNKGAuD+B/j5nKvYSVS+zmQwujrTUVfHO0k7A/7uFAQYGgBv7swcdQJJ9ZJwDWi
7/6q9FItRsOxbjK1g1Rgi4OTkmLhQAQThqK6FSCrRFVxKxzjGwr7h+mT/F2yOtGc
YsLA1Ve7JiQoSwhCm1pwc5MQB8OuVe05j42P2D7i+E2YtVu4MYym+6s6FEbLM7gn
c1bCwhIufcUL0t351KNU21BU9BfPdBfv2HRQ8B8MPuYDkEWzkFoU1KFb/N0tqilq
PyA/Ch56WvScd9p4tNahBlqUTbLX6sdQCI1IQvL3SgBsG4i4VDm7V/zLstOTG0n+
od0VUUivZxdspxsG2lulC1aDxbrXSyWcT4BfEuIawpuAH9fhV3ryXZHWQZyDLrKd
vgoVz0XKq+R0eUTQT4EYmBnQrRHun5WCUxV3qSnL0CwdlMpk2T+QDmT58Y+q8uMS
iTSW/Yeo7M40d3oA5XWFKHxnruBcRKMPfYFcDezlN8GrbXNdodhrDiZtfXoGZJcw
1DoAhJ8fb6/xCPjBOCAqMgZqMizJdKz/ukMXGo4GimvO6h0527CaSy6N9k11JLoM
wrv4JA/cKhr9BATTU3IFmUlW8Ord48vH72S7R2ZxTvZFNAwFvQEPfciUWwFw5cwq
VZX0N1oNRCbPm51qo0vQdIC78aroW7WvXbg8xawsPFEnl+5vDM5D7Xit0MjmRbwk
0qa9hAXtYhFkh0h0x56jbunNWnt6X0KQ6bwcy1j/ZOOsTbiuTSoVc+/QU4VIicF5
yrYH2o6PWtOcaxl3SjyLsJt/ZqbOrY7c4dNnTevdM8UIH7XYvyPhrxehiYpzcRWP
4rZveYb9De2SCAbILpdqpidSGTK2+XhFdjdR87lnXK0A3RGeFS9cHwUQs4Iluqwk
qn9flIe43pGqfi4ZHaqHwQgqiae5NfZEh3kpW9EsTjfpj71B/Dm+UtwHO/0AA2ow
igqcUsd1pl6lRHQQgF4rXl5wHZUfBtvNwgK+8G1QaU1L4/T+MgkGJNOXIIpc4dxw
jTKYE00yV7gxMj21P/SMv6vi5AL1C048mH/W/xSIS4437D+ZOAlcop4ok6cmKoyy
1rIRS0d1lu76aTpkrirox9wxoMGGw99RrZFwcnSNWE+oQrZx0aNtXfMoaP1Lp82D
Hag8OSwtvmBPkv53df1pixK7g7Bmkj3rQQUTduQdYCmAYPGQEcU+GooUsFhAVhq2
lugvm32VgBYIfUoa3kNMD+J8Cv+T/QWyxE4rllXVfHyTlL5Iwl304Mus1xVONEs3
uAHVX/DZ3swwwMke0lkrBoaH/JnIYHbDpTygA7+yAeC+MHkWStHbSfR9wsnbqz6Q
eATWy7dyCg44N5olkOE3KLUL3t2gtIq9pIsA6U2S6x+oGa8hScWqrIK6Wa+0RrGM
AmVJHO6z4wIq8NZXN13NLOGL+ylNJRq4881D+Qcopve/SOvNyi9gK1V5E7fNXORG
/lR2g3oWIpjNlw35JGm+SwmmRjsTRMVu9m4kPu8lPya6NuweltJlpJV7Q3E4QJDh
h9oO1wNiX/a/DQ8sEX2st0WtGM6JFawIdprZxx2wwr140hKaosiZAZ1jGGrH3xU+
RH4Xvhu9aSqzVfQdctuBTjJUgRp9+DPabIXGFAoEUHl99ASK5HO9lj1/8ZxxtMOG
9SVUJ0Lfdm+S/LtOZ8/3pURUp/O0sh0vReMW+E5MXyEnpsrv5Lm41JlBSjeKMWmk
dXm6/tS+6sSE3iZsBlkDn/39p3HDFaMulia9O4wqzdX/LhLmTXsRiIwSEcKP8pzz
LNHIRnEjB4nhgwcFRxr/XUox5r0Il13bO+E17cu2J2k7Pblv0In8ndXmPYJqC4af
J6uD+iSaKnYDCenYO4SP4MR9xJBXsZYeScGpm8Jv/IYe2L8bSkZVKXE1YcIu69Ia
h+iYLDMp/cP/smTIKBqrJx3smFIcznphO8Z2WiNQl/PZsj2/FwHtNZM7TdJzHobf
eKewOW5WnJJlyZe5VB/VMTjmufQrEkpP/YWuPG0veK+C0/dWuX0+GbbGbxvHmbfk
7arMduH9omVDPznvxOhyBxikoE3/+l/NKRWtXwNdVIB+vlb0TozQ5V3H6JdprIRY
uG7GEOSL5PvxOAbZTgZHaAKk8WK+78X+XDhvQXL/m1GDOkLtgHzuQF3NsOUFJ2Xb
x6zr1JDvO+I/+M8EwxLfWp8URuV+aO0FgswMZ9oNpMN2RayBL7CWVOWFIzZDM2CH
ldgKU8lqjO2XmsDTppgkeDmwi0aT2Y4Mj/xTPis5PA/9Z3n2f9cIfKYWacquGXCc
vcJ2HTVtu7uN41yY0Sn/z1NsthrCmLr1uJx6QET22G5HBp22IFn4RMboxCzaSJKq
RPQlWZu7F1m7ESIqrp0vELevR5WoaSYg++gFb9sLIu9ystNvax90x9Z+Qdp/FNiZ
9XuoU+AfopK2VJxhbsiQlhyGjUK7/yzcnHFvZOS4Ig8R30LJU/1ljkh26avAUsaS
OBoeoTbjlfC8xZLoidFBnFV5JreNCvmIIHDbI1qH92Udf81oa36otlBOx1tbniDk
G/4A6q0eu5M3MFDDeR24Jv33K4LQ1zxy67WTQRgkzLo68EgiRaLN0WgN9gA/qRR9
2tpJWGqvdZj2iaQANXfG31Bx9pBYYk/2yO78EGbGMO+d+5IQHos6ehi5ylYBz8lG
543rulwwSj7giBPvyWbMUwLw6x53QSM9fDc4xpITWXkwNk3HNXVYv8WCSVLBR/ur
DY67soHKkLsSGBCALmNE7FMGGXyiqPqAGEm79gf4kViCYI+hi5uTaCJzH/xghu3u
pWZnSTJT/Ms6Gsbg47Qq9cIcfjyXi6cID3xIjUmHtdxkfaskkALfusiNHcoEjDSK
/2Joga3qS8UgkBxcCa8NLyGuDmaoo7x13d3NjpWHaFBRGtEO3AQHKYhR6AZ6XR8T
13k4vmNGeA6HZdE+UhG2HZFh3RGaj2I2CGjpMnbdeJoJSFqs/l9GaQ/sprcHe+9s
mnGZbwDN8zZnkvHDJVx+ejgTkzXdE4rvLUh5xZL5TOcaV7UiRhaGJ7hest63WsNX
5wX6j9MLEHGE7senxvqUrR+RszjuPO4TG5yf+p8urZUHA0BDN4m3y48DYDsPPBHd
S8+gIYsZhz3xbV6Sg8zzfAdSyxUK5hvbDwptH7+VYB7++SIWi51EShxW+QZRpH/y
rSaiULKv0iNYIaAsDzG5YUkIl+EUr1L+TxLV8GD9+ci26eBtJpVXpVNhuthi4JPu
z9XQprmQqY5yGpZ0+1uNTdCMljrnNIVNx9rwiqVcUzejMxrUDx5TheHznk2MSL4o
HsaAORwT9Gz4usnp7IHEIldrdeuNOEYJjyUVFkq3J/upWIXq5HaEDJdRo3MT2UJT
f4CPYPuvSHLrNefsEJNUjjMz1EVVF4WsOtnailM/Bwm8zQkWp9YgZDfgft9Kp1Uz
zXFsbNZ/Id2CCuqC8BRcL48uGqa8eHbhOVZ3KV5ax6WooOv5FcPoAMcj3YRHdHFK
n9eGxgPR4QVaYXgHipaMaYNk2B20vFJMEzSm7V+6N2tscCkuP9GUCAB6bRreFMXS
QPzBl8uy01KEqunuB9mAX1Z75FgUE75FcXGhAx3yhs0ele0BqFmeJiFES3q842F/
TIJLjTam14uYryaPv32vv0Is2q1JVky/RV62p4UHkT4Ku9WPiZoIjQQ05ZbHvW4P
jlVkkOObpvIoLB6+gOmHjWt/K2GUoRbn70ZLopYc9PVTAvM4iENTyfSDIRc1g7Yt
cQhf+r2D9fD6DHMI2ju0v0gWMdamslZMZvZBpr5EmFcnQi6I/0P4aZtyUA918Ovc
kSk4SbdGKx9BVWjh7HpXmA01oJPzZ14wlqcyc2uK1Lqik2jlEO/VH5y2nOm9DR3F
m1wgK/ikYEMuR3JqaYj+xka+y29dNMB4UCQ0cPe03of1c+Vhw4bpnclRJyeUJFl/
RIWIVtq0zZ849HIYq1VYUPpecE+kwIrP09xyiO+U8h8e/3A0U1G4At+CBPmbyn0y
G7OvyqduwcUIT7y5dkxrdSgJpa75MlDUqji5L6ek56y7LvMWrrJb13rm9Ux1QPS6
2YOWxrtxUCXIulEkqRYX+qL1Y6KfZDb1BYhoTm7VxlLh4jjRAWTQ85cjdUJtM0Ly
rCCbOFuIPRE4iOrZsl45AvjvWP8/VxMc3bJTiYaitIzBAU3yr1glNeVEYJyYvauC
Odo8M+LtydgLs4Mr6CK9iIfGRUbLrjLBT3gvbDWNUgtlE3NEK8y0KB1BStRh9G+7
beRkopvCZfwvcLDmlukAUX4LAr/Uy9/n17y6b3Y/0FE+D0XjRDevtASr1AGQ1eqi
jkcjO1cg9qXFk7CJezpHsD9Nka8yKAKxDgn/5uWRNCnDhMJBa3PGFAiQhdBBchF2
wLvOUVy9E3a9v0WqXOxVpv2RrVsuWLCBUfYpT99RKNQOrpVp+ro5TOxm32L4evqT
LmzydZtpEgSe4ZC/TRyhmTv84X9Ukri61CcaAckt8pLW6Hotl5GD2JXhPeFM97VE
Jr/zqJvxRAgBc+UoTmYulXwlNOIdkQD2HAvAqVn6Qby7GQ1CpXH4CF1FcBIbSSak
UmrN84kEcnCF9xNqb/aazNmxGbb1vVSDFjZlpLdWgdXNN2n5FVBVXe9VfVeLC2+/
TlyD+e+ea1f7b9kirlY6s7JCli/2/ydqBwAl5AfkzrPMHm6K0TwAG3UOI7Q3ucsr
fotJRkngqHXdHFMeTLRDFOvg979653eZySNnG+VXRN4QyElaIqKHvKIslctNmlLK
Ve6dCKMXDvei4rdY27x5SIadl3ry6lDc9pKfAt5YnNpvx4l9BXKMayYY5udm5mx1
uDUu342diXNGxG4mBk2CGbMVazfXMFDhMvOSu7lbSjP3wXAAkiqLL0T6XfVw7cK8
fxgKYfgO+cs6F/56jmuOWgX+QUuwsUbU4miBmcqb7NAPjG0zuCzNX8xo0k8FxZ55
iwjCVuq/osx+qbtYLab5QbMgN8qgckMkDN/fAOPs7VzzflBly8aRgHATB5MJ2Lyw
Pd9OWUEvuqSf1gmMxb7ZQcecYo1w/fS8r28PN9S7YsHXsxeV9418/XJbhORsH1TN
vWNojYdFAm4Lp3uvUfSTqneDtdF0k683UGzmN34JpvsJUh6I0jMaWfgvpe5/RcZ2
qC/v/mDAW/8HovsgD6mYFdY6JtQK61VIHqmu5SmJ4TrRcp5zLehhxcfeBAcH6Eoz
UgPvsOdDNG5L5Ou49/w0JY2J2T48D3wNgLZ8AWzKyV1RH/SU1EfXGsHOq+9UUJRY
e2DDIjIZJu+rB7jaVXdCFuHviSjy1ZDrV8h3PGlT0Dr+hsJWfDw/vRWAtUCiNf5Q
xzT9QgcEz0jvJmV0YUliyEKATeXrMr2i0dAteqeq9wDaz/P9XDj4N3dQwsvfizbS
YQiDMZtVUm3mjTxpPl687IyYmuD/useeix5GKRbkZFfvOTBwBreRmDDC2c//wb4L
8ZySqgdhXMcwQiI4nEUtgpr7M44/WkSc+Ccr1/VKUIBUVMdVaxix8z8i/BnZ5ZxW
H0n49Hc/zHOanFAYd+d9RQ3s/OzJRKmAT2JMLnqV835X8X3tCeJn4gm/xz2YxLUF
MAhZkGiO8DT/VU9OboeMpNEyYHQGL8h4TyE3x9QvZCv/gpYAoik6Ua85DSsfnD20
4dvcxdLXskoo9n3+ngbSjsRHTteOiXFGUSKfo7mK9b+OLHo+bVrN/89DX16ex/SU
uZoGGhA7g+pX2Yz81zcSoHlpdeFBju63pq4Dp0Hu3pPbVlZVU6PLie1IMBSpDwP9
GByUk9Z3KcTrQK8iQfg5vc+qwrbGvFlcW0GfRlV+aOUCVVOt4AvLcy3G6n/70YU4
Zs/o25OxJaXlau7yemrQoNV2bJ89TEokstMirmpsggihWJMAvWM9M+u6rdliz8Bp
2j/Hi9Hsy8bNwQ12uJOySFHIDLluwA/87bVQPyDXy/ZTsoUtP4qwCCxs8ctQ1nSH
m2+NwSsC+1KRJ9ZS5O5FR2EWYBwmBq7NYocPBrVJMSX6KQ4lIL/x5kTdkweWGvbi
8Q/tMMRaXEqBMjdUVOIb1toFcNytwH3HlX0VB6lJLl9N2UfWkqJ3cIOVhbUEPZ9o
IL2JHMayCqQhLNkdq7RFWbcm4gTxS1QgGRM3rNRwAuC37xuW/z9f8zPS928Gmlyr
UyJKl317XeJM9WlB/GtzSOmliyzMrqlNwELjsBPbDXKMzY7ZYdEKDJQLCuHGrc+v
aEeA9SbtyRbrkfHVGa637nF+FYs6lcHviSXMcndEQFq4Li0mYhOFhRWiFEd5gyAH
28Seii9jy+r0mom+j6O/SndUp0vZY+67+T9MGecSHceqNhXy8zZj/hS4y5vZPB37
GULTpaOCnsQNeqMjmur4fg7fW2Bq0iPrWZ9Fy3wu0QxzsXwAXVYpCodwf04PqQmP
dZDj3z63DqjT9a7/bKD8NmViTt2Tl0InOVe+v80SZ6Ajv/NujO2AMOowBD0sBYD7
uNKzHPqwrlkeP18uv9pScYy7hjmOK+ic28ulBTcuerXjMuYISIfdDKV5UxNfvK7E
WCXY4kBXV6NBiXnwq1Cwn6KZ1nP0/Qu46ZlWTp6J4qzQtrTMrmx32qmBS2CZOSRJ
P1GKCtkGO1FI969COzWz9/O1psfqJ5mGNmaQ9TbOtTJ2nqgMignbQfyClSEpRJNe
vgEb4djbfzMQJzIvHe8xfHHPVeLUWkLywsaF9vtmpuggg1aWpiYmKHCTN2IWNxZR
wsF1MQJ1gvGJKqWUYkITvFiSOdaZ1PdF+eGf6wtwemYzvcyDM4bWmuxnkaI2kedf
0ynNngoQuu6BfyvWWysvRrCmSb5txBghgAftu+Ytay1igT2K2lSbC3mM6RkHaj7n
VhwH5DjTAgj6r4TdpXTBhZZibFMPcrgrWICv7PvF8Jl1y14Y9ieNP02yzSolmhue
8kkE+MQIV71YkJIpi7CAz/RqgUi2JXN+Yx75dRJCAMMUI/2reE+m5KFDOR4NkmFh
qWKU8PDt+n7pLzGt7o2TDAl2CT02WmrzBSJUo9yXh0VO8h8aGKz84YYp0uPekrvB
KOMzLL6A8OaNXlcnofBrD+LnztJ58Z8V3or0ZghZCjG0uYt+wSRt1GcGM9uUJPWl
YXGoOnOz2aUHMdqBV8Jeu8PYjHxOfXFd0WhG/A5htQfgGwRTFpA7ParbYh07nOOq
cvRDMXUHiOTNa3+DP87UHIYvqfeqF4lJwlmGcttZBM4bbSBINF+rhrh7jITiqznI
LXmdSlMt3HOt/UsDrzAt3bcm8hSS1Ug61UWJjVit6MWJaryj4pDZVbYa8xSXQiHm
IVOSx1nagKPah9y5PAfk2ZIKgQjU+Yf2IsgvpnST+xCRRxOJ9NgKLSZVivpBEJe2
0G0oeqkSWJ7PUfU7zoQ9zMn/kchZAfJO6nzt87iDepZOns5r8peWQ4Z5GDNA8qG7
T/6GPvtSkYod4fh3I7NImRZEKi2hyZ+gcbVNtfZm/4qOO86CArTONWXVRIHLwyOR
1WOrE0w63Dpp1fybkHs69+iqEGGTK6bTKoTTIct1Z73VTOHHByhhOaBdnfWk9FPC
VFb7d/VuFXpAW1uMyAX24/jBcjy4VJjj7e4LK/Voq7mamCmSvltNEmWag+2YkCIP
t2+e+q1xRrmq/wQvC+AcYs8Xw/ChXn01GULQWvUpMhXo+3gttiZhoaKdWEVkj1w/
RFhaMtd3SmkxwedE86khOv0HCVe5pwWH8elgWHDJrM+6HZoMmDphJ0O0P7+6rFEf
TWGTREEmPl2GvckqR1xaTb5YhSRC0KOj4HNRYtp20HEAASOP8e8I1PI2Y+N4gUGr
S1EX2XbYdSmNEtGaD5ShmBHVmGTtvf14nz1oZgaT5PWOphhb/IJWaPVK3W1/Ginx
n96vWYG72w1mFXwgLRC9Z1rHWq8v09ye9xgnaLUZnEcOAOAEOrKhU+Biqeg29VTn
1eOf87s0bCQSbez0VU7mU39wFH2Cv+FUtONg1vJx1JDOHL8A7FmFSFNgWYLyIfu5
pwgRC3t6qywmjCupcrQbxQil2fwWDCdboN2F1ltpOoQIoETOlxV016yoE9n3iTGj
DsTVKri7SMIMQWbr1bDQIP1HtExYSZx9waXCyQMcPY/PSXHOYevjk+uxSI/qqfhL
M+6z2nkMSVnmGQ81vM/cileNW1Rc4ytXw0ewKmWu0NbzBXorPytWmKGBio5NKMNI
KI+zM917syvSFpBlrG7x5uy/+9pET1AHTMarRkbp16Ko0Hcjj5ZvcrTP2Vt/dbWB
F8NENBJ6Q9MC4DK9/kAbGqmJvUBCIyU1gy5mXOb48Qida2I3LXobOygaS6hi2u1u
Kve66fDspBvOsjTSYuQBNR8/nNySTNBo+9mZUI4Y7xDp9LjxSvJYja2/rRLRy1P8
l1aROtNOfaflb6lPiAqcjyteYMZbUr3i9FboxEUMtICR8Qr0sH9lbHabtWKtqTiY
IVOs8/3ztP61D8+W7mdUBwgJdS37sMsPuH1wEmTSiCLduLG7hwXix1vVVpugZDA6
F/Q666RrnbScAgm3Wcfwcsy4lodNGVK49Z3giHuv7l6wVveOaDbrY5b5gKZPmbtB
0/hEoaq8JTpChiQQsF25yjFJod9FVXoTIBgiGmyDo4a63Nxj0vJXu/5KhaX3uPuf
7W6RFhPEBRPFbwdA3q4kccUtUKpM4m6XbkA0ZKLaBS/qIb/BvzzwfyZizbdXZQwj
tI+MHuibMknVnfinrfhyCOBVyAXgUoLSQWRawvLd4uepWFcO+R9wnMFH90JPaRjb
hmRGl2BqOG8E0V5IRhqbE3do1D8faSSFRiy5E0suVHoZLyr7D/+9T8RSB/CYb5gB
O6qoGPHu2PHozFqK5xOsDpQMyxLHBxdiD/6ZokFJ+xr4RaFDgZBTEqJyxgH9te8M
tM97SMv93n2wRtW3lIDOT7TbfZzJCQUnkZc4DD00WTxmJAJ6xU6st7/+9i21Be3H
7+xJKaE/PwcDqMLl3Lus3/KdjPOPX6dZ7Qwpq/Vt6AHI6mZ7vlfWfc1Js7wPei/J
hSz4snrLTjEnKcJFrYPboemHLrKxYgS/X2lXr6r/ATLF/9goZFCfMeWAwlSWsatH
gpEkenqpo1u+s6tfkz0dCaGNQIPrtXx6t6Hxxb8Rk8ahR4T6pHWc5GbfDmIge8ys
HSyT2tfzeUYke1IQBsrthCT4k8gQNmiIaa1mCIdeDNmrzEjF9Vkf/l8M5pHbAl/K
OIut3hj/ar+M28jXF2y5AV+hDOIbRG4CKGcHsc3zi+GQNkSYu772NQUjiekq/l5d
1B06vzzHh2Hmdrt6ilUpwQ6hciktY0KEWilLrP4ffvI1SZuu6MDYDcXMX1hUSe4o
QOzXy4NaeJXpQI9f601CnFQQSq0TP5/R5QCJLwuFRzBG6UQ9T0fZduNFS6T2JzHH
A4lWzGCGy0ZFdHJTqVW1gsr5KUygzYGULGxZpwAh4k/biCpH4V7gcl88I3fducF+
wL9JbrdU8H0hXgFbUgL+1w0kt+OZFD6SlSn9s7vA2HvosbZ+cVxEP+CBDHrPhWP0
uWtUdJhgzcIS/7XUqC9SwtCD9fYgRXbWi+yNLtjliWDAhxAsrnLQQJF58gQ0OBtA
qDOnkAb/56lhCxyAWjrFYWPVkvB7G048XhL0ABAKlkngCNaUuAyzVY8j7hzmMHfA
VNCDCMnz3smfrDDPKxC2Q3qOwQcnBibSEHyLajJQQPOVhpwOUbFwHzUz9iC994US
j5K+skqXA6P8kBvxZjpn6wcPPyXE0klfCbDHIZWAvededK8RU1ObUHwQu41CVObE
mTN8QsVkZHZPf2HSHBISb7G4LbY6uvX+zSiavNdqzdsrraEiR0N2rrGmQjr0OVUg
splJGN4oZsAz2EHjoeQ+qn+WEckM9ShgW0KTHkphNU3IDFzAmNGrtt3DJ/b48dd8
mx/efHJBBuS94iJmxI458cl5rqBalvFrJthq6cXfWCwQQsENy33Nofiw0O3OUMi9
V/q6Il7hsjPEXKS1mcH7wjEJO/o9z2yWFLUyLMS+mPuSKilGtuIPSPvmcQsQrnRo
54d4wS9cOGS99ckEkPQX95hCrlj0ySf4SeEHxq4mgjiwGlrRvftc49IPaivEUuUN
9PqJupkOW2aOhSHSG/7SZDSKjIPf+imnbp9vZFsUK7j6zZUZWvgZGpW7R8aJcRLv
m5Uvvxi/PDRJ+XUjcP/IHQJJS4RlR0JRA1ivzMGYBHHeXElU/nq/qIrdLtUdfN9V
mM31LWv1KFtseYzM1hPKR0BVbr3fa+Emxqy3przIYhFdIblHky+oF8YVuiMDNOnd
8CTHNCg488TFesHGg71YpDbGwE3PV468CMs1OcCk4icNTKL7/UnPSPgjA4AAtc6O
H2pL1Mryvsb9nmBc/HUVLBNDYSJxBC9S2PYnb6QDvLlk3jBm9zwlsPMjfU9GbyW0
eMCL1HH7LREP2ql2/p3nDsNEzAxsM7ONKy+vNtyN/wfTLrnicxcnS7+nwyizjjl8
dNhCIENLBAfKNK8qCtpdyOQMs/PGov3F+aBFRffpiB3zAHjaSsBJ3u68MU23+bYB
mmgVAHqkBwgtjRYwQrNo9QW0qAe4GQTqvrwCBKIMaBI2iLi8qmyJ6kovnVENC7cd
EmFxmKtReFAZhLdSwW5pTKXiGGbBfDBQ1wJ2xxbErecc2RuX2zxFVw/mESqIdjM6
dM9z2l5E3z81IfHzYpRwOyHh8ZxtC5gVfXnMUBB7vXbMs0rWc2awOkLSSx8zdaN8
bFAtouY3glgEO63ElW2qyssELe5VzwJmX+qVqAdQyHHxofPhY5mL9vJKKSo4w4kK
x3yLLkF2YxusbPQQtI0g5WtlNouS45dAl0U3C91xxSq7pSFsk1hm3Ln1onprrT24
LxfUWxzmUvYEfFcmY2j4ITApUw8CsncF47dW/CDwrHKQY+unxVPWiX1r8Bg1mZRK
/IrhQTwOKaHtAVspfszGsyDXMAheoOFtIKnn1V6z99OIXLQ1imns99QVcTKHrlyU
J+V0i0WFMWAxjiHVPT+9kNNZiTtMWHsGC+if3gK+DnmyySJox1DKyUIaheMV9NvC
mxU1sdceXkbhPYjiYTj4msnonwxxTnKjb/I1M8xp2RUAYH4O+27aI1Rr6ARfw7/3
GfmycjsEe4qOPkoSMuQR+ReiBR3Ud41XmSGqSH+rqXfuhjWrrMxLR+WEan5sk5d0
EJloaxqKUNO0O4hAFpSIJCXday+G0BOxmSdzkXA0DOWxAroO7jskOxtchl1rdIDp
oBZfKKKV9EqicOKei4zd90jQaIdE6CqpApHbnD8JSnLa+C3m9JmG+o+zSzLSh196
8Z6RX3RLIH9sAFuu+jnPPto0FXHsXn6S+ygwAKoMPiu+UczxJXyiYTMNC0Uy+EAB
KKjGsVgxH0b0Y8TIYrZQ2Yt4PC584lVFcLj60XWzYlaB5ok+ID+r/hfF32KqP7WJ
HVcZP8egmLeNyJD1JUniOK2rulVoE03zUu7+KCrkyTGk+36Whn+LSM+E46X2WG3t
7gsrJVoZJo11/kCkPaksESf9RbVWnFUOdDK0Ckn4SUQW0ntEwaHGfywQUgM8ce+/
Rm3M/bRyKrdPTlqjUfKOMHN3lgeokYJw9zW2ocDVP8WctYVG7aF63HMQ/yTVHQKv
oobiiFx2Ls/2nT3TwGjKBPEZX5xsqhdSLMz9tr+AR6pZgBxjsiDz5K0cWuPUjwYX
nsGSdZAcbHbBGr/8y049Ue9gysFfGp1sd6+4bBo3DK8sYEM2q6yejVatYiBJulOX
NzC58fsvL3qU53b6WdrNikSCCQHSavUUVD5xfz/uKk7b0lvcIv5QtM0wlsKo94Jk
BoBz3EIjQY+0cc+TBM43cnoc6DSX9K9vvhxddfDrExXX/M3P2EOJGEs1rAx6i0K1
LVdk8hRKsd3WI8f3CeYUYxsA+ZZdkxUajoqfAdAHMg08URGKpG4O+XMWFM3GP2qp
WLxiwxgjT2nZtal/ttDZFffIPwvd41PWGR6fecs7yBN1FKWytG+y80SfdjPYsBmD
WCEvExpT1E9EzLBL9oEq+I43bo6DOWMSXuvGXILRhejfdUKSpTLqFcIuic4MuZf+
RJE7A8SxORACwNKLpxZFNXASXuEwocQJWzDmoYorQB7uCY+yPF5Duos+D/8BC8+g
pz3PuuhCvNkMZcYcsRjthUw64ZKLRq4chYb1MM/sqiSvIPjugMIwopLh39LBANfn
p2q+CcQnn0shlCwBeZvOeC9nd//AZo1OYvcOGGhtpEXZIPz2mZXn4PfQjxrvc0Kr
cfWAAm7RECgXoeCpT1HAjyQ7l8iyf45bR0FXIklR3smJnYLEeUyJkYwSp4U0j2SQ
ckva2993xGjKQqjW6DAKM/omPrDjTqIPjlTee3jfv9CmzXfLcWq2b2rPFwiW41rI
7vqy0LVKhkCeYeKqxCOp231uPKJmKJ0zwZFd3oSVJ/2+SoSelLLNXITtDtdONXxd
1ZJH3oWLBH5EObOJIuDfaEJY3W6MCuZTGflZUYThc/6vWDZE5nUdryOWizAnF/JH
pDIETb66ePlVjIL2tk/A9lUcsWf2CrJ2nHJW50lAum+iv2Hb3UnKAUTWx1IF1FYa
FebqKHKzrAD6bZZB6LH2wWfhBiixD0b8yhXX5akSjcMNAqk9SSe6mU8AkUGaX1S2
bZv5mF/XZcRN2Wqgiy0lX520g019YOq+a2TTpOtHki20PNujBrhwbFxOjnkVK0u9
XHsnJqQuqqN5V9Mxc9AA6BE0v9q8OIND1pdlGXZCpDP3h3HWvtgd3kZx7RfqivBS
Tk2HOYtoIItvFXlUpPwjADByp4zAyKkyL0pdo5RrC2YvANGPhN7EqZibgI9hjkvl
c07jXDeF0Nc7rWswNGEZc2SbQbRz/ZE8tE8D09AFWdx9I1RcQ8k2RowfSZTwOzMY
6KffpWvscDH0SU7R8Ahed8SNwZdrk5NBrmutP93qaDI1VFQOGp1yQ8YUVyyor83L
FPNBz5nMTE3+UIAd76MJJqz14JALgvQlWoNJqcC4LVbYmPbg1yjQ5H81vnG9UwC5
TaiAF1wGwSdzv3iIZRZ776nHHpAZU5KsyDypavBmiTY1R0kJYaw/WqHY4I8iJZTF
S1nKT3WIqTcsbqksfH6D1H9Z4MQv+6J+i4cNN3omJeKhCzSODZ45fNYoUOA9e69D
tucyU2I747TzFAnbHvKcJudkx3M1lVfe+WvPsC/hLDbHKRWuEpKM3fUjpSiDBwQi
7FdDxzht1kwtu9SBt7EGfsGxeJ8FIyhsOk0TMac1qINLyTO4UL2o0lVc8IcjS4my
ydlV42Xai4ygpPPJgMjw2sbuvYN9HRple8MqpqjmdBw1rbQ8SgbMNDVPkuhn3iY0
OInJdatgz8or5KE//W6lK49FPS/36zmil9cme75deSofi5WaL+fgYpVE6uP2vPBH
jfOH/nwz6YA2oaRRcBYRc9CukUyIDN3UK7FAsnHdciQ61prxyiNnDzyP6OWcBMUv
fcNCvw9UoDTXPUxHkCXvLlMc6uOFvHU74wp6eMQiev8mhzxJELlfjC2tzV8Aozuh
oCIhVQIlU34m8IYCseUjnYhc1EEYG9HoVXjgSYeazz4WOUG0om9wTgBiBeowPzrG
mAl0cp0iE5VvV3JQRQvNr+1IxM6z/v0NAh8XvCUSug0qTA/DPeRxLrt14iAnW5ZZ
yuQRP9SrPsEXACjprmdUFwYgPysFiAMGMSA1DY1MZS5EuLrzd4d9LyvdpoRXvVLO
ss0ApjCOCbO/O1qQsYf6iWivTraVesZth/SMAlgWblsjMtFirjJB37Gh/dn6qk5L
yKbq6Uz98kt7YDvYpCPFt0xsfc1GT7WK0wrK0nAxD02mTghLhfRx36UjQGWcIuVa
E2Yz5HpGIukb3xj4IuD44/t7PNmkA+0AI/JeGybp+l7zjIgtpEmvKd9zEQticqRx
HzlKNqiaqoOsZ2wRu3QR+QNYJsD9n5/qc55AXyliy7HnQkwGC4UvAGQ0n/Jj3qDt
sG0YRMl/ul2DEq62xZu3NSFnW8L7GqDkmtvEp/1h0wF6s0lXc2Z0q8xw6v6iygf/
weT8KaG0ajW72kpD4p98sI9bZg4OnG63KjH07+lKesmF6A9hOcbOosfgCH5WScI6
1d/skH013OH/BQ22GQTW0ub0Und5JPQWRRI3tmmCm/ko6oTuOFEvaS9Njxz5vbGt
KOQ1Ke8ZFSpvoqiG8WKcgz7DLQM4LzaSzCo8/zorf4mDu8Cvr8cKyn1HygZWlOkm
GpVYo4TEfot5ucSos6UarsQtxHcRH7B90zucBnKLtbmeCR40DqlHmpo+npb3xBqg
w0NyPeNx1c3BUgBy0Q9RhzF9iXLV+CO/KvuD92dTvy7HdJKYzdx3whIwNY0JOr2y
KbyshLkqt6d2DMSFJTUVEO2YtqKyCULjdGlek1wh9zotQyDYGPL19B5FBr5Q0IcR
wR/XM/2God7+Q+qQFIBCwhlXZdfh0TP6VsANnR8egeyXT7IatYYZLT41XLiMRFMb
aPZuB2MsMWtOzGsfNzW3Q/eMqRU9BS/iJP52uBnMtt79YMEpBGAj8WWoH2hxKH7L
Ce95aAAYzJZlV5UfwFUcy4QMKUcI54bp5vv6ypoyC2fYcO/6x4ZxlVYHFdLxAaf4
ucDbVVjEKZRf+kND4nPiIhY6YzpYkuLhGpoenZpjzXIbeFHk0cMOqFH7iWsYtD2h
7TLXzbqBKttQtAE1632JxEJrxNXTuDJnqJAI3PTBf31kIi8SN6XKV/5Jra/3o1US
XL2E+da9eHLZw1/OOX/Us6kpBaRAzHlB8FZ+rEP17JAZrpO8gGBhFA1S81K3v9Z9
TFlSsqzPHKNV2GHl8jcxdSqg1ZvZcBCSCvD4Kgc81/p2163x6sVSrvUGHeH+gjXZ
S9eJJTSzYd/jyUqGtY5qn1XM1Xfhg+tVxqFV92tIdCC0QohNSuTTMlF9tUV0lEwm
d2FIJ+tuTsVPLvYKPK2J3b1eI949sj3ZVHK++QHsmeep6O1PsSPYabLONd0opvTQ
N/1Yc2Oe179I8KJxzAEQbE5TW57290ah1gu8U8LAq2jwZiT6g+f5kj30GXJ86ICB
5/htGyX8x6JDiTnb06VFNJN557i33FrwQeiFyfDoleG/VRKbFCItKtEHWh1I2yt9
T1N6g77rBG79mwh4rt0haDFsGzyTiyMBR1XIH0omTvV+IQmqjS+/jLSFv6undazm
8uM6Vszldr4nzzTnhKRdsik3HrjhAd+Ht8iRkU9SB+1gXsTWd7yQtN8h9u2htqNQ
hee2L7Qv0DUS4eSKVr1ClBFIbqr15R/C73HiA/WHDWuSjti5r2ULZEe7GdFl5oNx
ZwgJfHK8hpORw5EGDXzUrnPDaw4X/tCRYXY98CbSh59H+7iiG0Lt6o2B9BVLo6Ox
osyq0VfBn554m1QkJPw9dM0U2AjtWc8CG2D1MeLTUGs2Y/rmi7f4ICxeDy0Tsqez
SRTKhn2nn/iT7+dlTDHRjuf+bUBry61ahhQgdCerISKyixfJd5In6TROKZoSqT55
128f4lYd31LWw0u2T9vuCDvE7gjEz7NXHULHmZaan2R2Aq6ejJFR1fSy68RSPQ0S
5H/tUqA4XQfbRTN8a7pNhEcGCvoQCfHwdtSMOOWxaA+WmqwDG5c58+6XsFjx7lFW
7TzQqzwgxoA3nJDcsrrPa70LCA6Xz1UPeQc6EuFGObRUzihmqwPNFEABPHh+oGCd
VRqojbiv6gJzZWGfzziWOkWJlNb+d5xEzCFSdorRwluYsT1pGJQ8EL9Nl+7vWwzK
uhyqgEmyfl22JZ7tHAzUPkBtdNfAhq4clQIIAr0EhWvK4XCRTY6Ee7HgJEH2aiR/
3bxtiz5euF08u0xh83wMBqarrI0ojKbGflf36tPy3bNR+2FNa5fbzh9oQ3Zg6LVk
9wuZyo5LGLHe4cCaYcPrXKVXwuoOJPG/C7byT7UlnKLoSjD3V5ACpeFKA+vBKdGw
51UjQzANyOu+Ghydwo+xh9hhaTYrtIq9mTN8QawK89KbdHjOw9j4X5W6Gc0g2L3x
irq1PQ5OJ5fvyWE/pv1MlTTUr5QqNfdaTa6GNUlJvUf5EOIFmfYklbBb8y8siAXf
4RBI7ix2z1hdw4F5hYN4jvjzaZ8urX8BWtjvoCGbWA0pqlqQuZuDgr5gGg0+jbKn
ZE3v0R4YTEYmjacuDKZ0iHZtwhdf+n11tYTXliXHdUwyMsulsF7jwiQOAimOrKkJ
xQmkt3NzEzsc7Ya8lVZ0WCaBdcQBSRFtpUmLT6X/Zf2ntdIbpadQauDkw90UUlFD
qAHcbWSPaE6kMyBNBZtGUtBE5+jsuEHs84vqprtgNN0DPVZWz7C6WsnLhleAJYnV
8RCnaojrmbYvXpFt36mBk97aIA9Nkv/lpzwAZDlIJr6Z7SanYdQi4xyVojOK0Dov
ag/bjRJTDyrJGcuduCYiFvxpgk9nZctM6cWp7LkB7VgtbAJ5Y2Mh/SME1ml8kaMC
W/lQruIJESdfc4fpYIGdkQFIjZkLsAqr53y1VFXegGh8kczou65D9i4PPu7bcejv
67ZS9ndREb5fGJ5l46p1A0J2glO4BW52ZS0ULQjMb0wUNDZwGL6dFseMoEJLwmIC
iUddG+gz+I+LD+zAWBvXppuxPTJdzuMs2c1SM4qTAGKRXMnApcng6UBaXNunSEGd
IAvjrRFFJIIqu5pIIFz/71kVw6VEZ+sk6ow0KhOZi7eSapmOPFoKDezv4vimQvtf
Qu1yErQz3+km/XrPdsVlyRFskGmot4sHhlatykni8V+zLtbp21/ZSrcHQhIM5HqY
vQ/4JmdwYXKgvLvfVWJULR+qreHqhCmhs7ZojUgxNlfqa3O9AtCYW1GfdZHDITum
o6a0sguT66VsIhBo8V2KxXhhRLTDnpyy1Qfh7Cu0eV2WO7zLKLR2aV570jF9mkOC
Dllt0VEeSDe+0nKOlWPlghT7p/GjWU3M+8wV5VEuPBu0kZ/iv0NYO+vg0Ho5gj/R
/5JYbpTAQ2paAyJbKEOx8renOuf/kO05KAJO4TP2eCLsgSnn/x3WMybaR4axdG+L
QAuLjoB06USt9KD2ibIWfAAzoxNx0H7NZLWO2xfdMVnn/vTrW5A4Fs7KrJ1oN1E4
168i488rwu9G3O/ofnTsxQI7ipW2FCBGQmeHP5D4xgTDiyCBumvRRbmejIlXLdSB
tSjnDdP2MJgFZ+KTv24IxON9i/Bqf+22J7aY7IjraWoSfLa6LCDg/FqM9ZFdGtIZ
VTPWOrQjiEPky7ck8GBR86UPmqHKYyS1BDR7OHIWWz3MRmoE6ApmmL2uZlq2hPzS
1rSvhnGq6Chg05juVMYAoj9fsVPHgtTz7h39i+Gx0v/LxJLwlqB/sSSVq7nDzVrV
psOMrWXIZQb6qjmsljaItHrItJ4cTZMFaOUwRkCoNJ7uuX7C7kvhOlPvB2vUxBJH
inKJkaqao5ALsZd9wU9JphIgGBTmDiwdUqHAdIxSGJYxICf15xfunyD9jGIM7viH
TUDf1SS+qi5/0tYm8pGHg3OIiSNu6fz0Rhoumyc5hPe1UdzyHcJIlbZRB7dLOd25
qQ1xAzp6lzq6Q7yacOvIkSZcHKFuwh/SevNNhquXhN244KR0ba0Hu72TY6aETESz
00F8s5K8yJEDKteqmffZ+NrmkLR9EHnbXEn+4iHINYnk14gzVSFpySG7tuG5HVnk
OwGbk7lUnLZ5jR/9RVcMALA1yI89OM1EXqf9v6UDEtzTzPro2y12O4NM2fTlcb0A
z5k+QSzMBMfx1jM9XXcsXCV523tBVKzbQEAQE0OKnDa1rEnc2AViIkPjTE54Ozm8
zdH8VrpoJp/k/NXw38Io7piyzFnGFdzgTP8/MUc+WdVw+SoGSknC9QGQcAHorX5E
PJNXyKl2U58pc0Kg6Ftt5dPleU2Zo9/UJXvxus7NndGOjxLwoPAEo0qs4zKY1A4B
BejwLgHRPP3uIfGfubua53Rpa5vcPGjleEWpQl5HJ4+uC3WbC/9kkZStDKu+DFKW
v3bvfmZ7fHdMUQIwtzo+NEt923w98rQMpx+pvyYlaCNk7BIsoHKSJYbpv0BXBWQF
NerB02/ow/yZRNQNYhHP2XG6db5HJqsTXr/Pq86cooZ+yDhEvhExTuSUbPSLbJz4
xzW2zpkSyZNBh7V2IMuYJp08HqM/Fz7nHEge1ssGAaEME5gFXUy6nnJrYZ5ENNw2
38mZhJhFBahm59TyBA0SQwAzQe8gEk0WJIloFp+tHBmrHP5mpPk8KU9Li8VwlwDC
M0bAdh+k+tTAxvL7/TFE56L51pwEa6f/BpkzfC1ShnIUGpjuO5BK8pGFe+7+q/E/
P29jaL/zhWl9XmY8t30Ek5LYR5DfJaLyI2PXA8+1lDvuPcduFQ3acDVoP+s2YGvv
biLbk1nxVGpTRPntupuVZ5zk/TOClcUKW6qre81EkKm+5gSxkLxiRlr8c7PcQTPo
7D7Xs4vXEwqPrNJLGSCPeoQKdR4xwn0T5HGBCNbA95tRye4Xhg2qJXGqsOFqKCa/
MLr1IoPBh6kFD9FeX6sfjHf0AiANpSPA5c63LWvjXpLhr6CskNB9/LdvCvDUObbQ
l9xAsCdg16ajaNfVwkqlot6dObom9yWMsHqMf3vi4VqjAMP/JAHbO21MkO7H4QLq
X8P1/2z6nTuRiELICYnKFw+A5o0C3CG0yVyv6wWdzpgLUCu+J1ccK8geoipvypxD
DECpqMfb+o0P8RCD0lVA0OPm8LZNX2lo6n3d+nBTlNmqcTig5uwd+BN6kAXxWoXr
jeJsXQHlelmuOV90zVnnEEeTUBirWbWfvDyGDuojLMjQokRJ2wF/iUusV0cdm0qV
/uQDV0QilpYIzH7lH2S//os76oWRnZTcRSxuLXkCMOPKNfYlhQOKNVN8Y4rV4ued
FDdHHAEAXacqVAaaqZYuI9goWfKRBFaPJX7OlJ1No6YS4aBL9MOcanhi+Z5JX+Jz
9/GwrmpV/umUEKX3CD9sft8hxaLPDf3y6jKlnz82kZFidI37YX9w4VHP/5BnWtPd
paH6drrTe/AJZ3XbmyLQVHxrhvYlpyujXIg7kl8jD85lju440ywPllPbSO2Ozo7j
jOSgwQ721xcn465nV0AJgPA7c1nmTiI83WNJ/SQAlrth/Kt0p0mFRg0fNge4wCgi
p5CzaIN5CFE8qX872J6cpYLUG9GmoFa7TH+cDW/+uwavaHGjKIScjlVNR3EKLgK8
pOkDcxcCJSXntJ47nD87czdlVPc9e3npzhS8o7DgrqiU+Kb37Q0Jfxt4wnbgpzPm
K/3ctzwDple5VxlWJwPKrxVvlOEiIOv0KWNF5wbJWWjzU0U7geIQQr0DXblTc5Uw
djjWk70QjjIwKYHVEl7WBSGrzNPIbvSCOKqiD5l9hqAH39S9c2l7iZ/jr9JrL0gi
52Dzr5h3aYDOG98k84WUAh8mteaRfey5qdB/cH88pyRagnhHihNvVuuCwQ9IZf/V
pF/psT01/fdSn9Ey/crUa8zciMqgZ140Pv3W2V0eciCH1Irn3RmSp4b54m/Dbwzy
d1hnbLkX6LRHJ9H2TG91GCH9t9wpbJHXCcrNT7lu3fWIeO9f+6w27njBbDbz4PU1
ir0EDGOVgHBPemEdjPFzhrx79Ks5uBdSej0PXj2Vt1mG2K9zaxo54jklT5jJULPi
HC2r9mg8T2UwegTUumbmsaFrZRjV7lIMsK0Z/N0CprX5SS9pq3p1yfb1p+3nZvqV
W9HLP7LBS+wHwzeEqCdSrA9r1V+SUpEJk+ryOuJy5zXO1YDez/nd/FWV7+eCLIDb
Z+a82QDSPHbbZcP1g6tVNdlSqvwkSnwJ9ibc87g2/UkINaK/3a/xesmMSJ29mp39
F/pBsUVAf8/D4bjqA4oeYKY8B61+qk9jCA9vPOM0afb28MLJY/Xsf+2ujNOCO17X
qbR+8TgzbYZZ8fVV30j0/lKfQN+cwQwgYl2OzqAbt6U8N9z5/Pjp6QozYrVITWO/
K5WVskZiLdal7scXjWTzLtIHLSTN36UWKkKoKKCcgd83S1DKVm0vOtW/pvWaDXMs
r8Q2NpK7nk8qDk4ctFM6FcugpA0A+T1h1jaQfyR87qh9WndHrWFyLV9dL6odFDh3
wbm+91Q2N1adxeOmqPa5Cu2E2IxX5tPXPMPpWKUQck7KsTWzu066cid21AiRzCXb
bF6Io4BP7BsrwR3D/BMNMQKpDRSgNWvoJvmBtxVT/wsuRUD2h+RphTYzS+jXfEgC
dhUrTWYdsSi5SM0flC8e8vbR1s1TWMorpiiR3XkLWU7PqQcKHjwn0uujf9vl6GaZ
fnPMDy2UsokSqtdw9iSY0UTHbIk0lcu0hafveR7rluQh87sKzaZg07paE468RVbg
Iyl9wweobNDVR6H7dE+ZeVLK3DkvaeD5O+a+8nodrWX+2jqnJEtkKTx34alwmWUt
5dvswZns1TMOStaXP9JTnJfDIRoSj+OOckOZi2ts1LqM8qLombpEqtimxDTlpQbP
HUpxS2vV6TXpHtesJxhleAWvIt3Twp+575D3NI3eEKbkOLXT6/+4oip7BqQE9s4y
rJzMsRhf4Qy0Ga8TicMkDb/UZxiIIIGgI/QCaxrs+DX2HsgdMjKXZp0RQVAGBwb8
zQquhADTy0VLJpYTHB4XYTwp4QeVz1VLP9nbzEVDpr8tS1A/5KDBON6Kn34MToFM
qE66ikAX7BFjSf3aKHKX0qm1AWz8eL35Fij1H3nq2gY33FsdSirbovQZFjTiLwfQ
/sE+jcuj3T9aZQ590ku0ZbB77Xv2gotn6uFdAING477hCLfvaztHz4+A8PNvYhPg
/v4Kyq75G7MA9ZK/gOuUWZND/fx1LAvmqT4jX0qVrFsIzJrQt7nVc8LDqA+cdUqI
NMSIZpsXI9Q9Y5cIJeqeWXVJpDgMlqLYWY3IPntN+YJSm7lAYt5w3b268e8eZCYu
chW+Zhm8VrgbW0PgP/9j/kit6i892+eErpValNGcAmgd0iD5gO5uDdKW1mHO4PlO
4yMHQVnAUXww2xQziGeHvh9J4dSp97VNxQU9+CNjvLLep+9YXZtfN4PbWk1rzki+
M7omtgDx6DXUUuVTirpB+Sn6lfqdG81aSbxx3+vFNth1QJ19DyoShI15JZd28cgH
YZLRgeLSdqzeothg9I6AWO84vVEevKcNUIJrRGaeX2vJAqGc0Lmmb3HQBhVBJavQ
ZE6sibIJX1Y/h0wsVTc7r5tYbOKHb0mGviK9KmKt+YbXxeqH9Z6LsGkx6tCeVoFP
+vUcHpsjm54gLQxqcOKmJZ8SFWVlFXZFDut6wmOn8u6LYqjpKB4q9Ld7GD9FTsZj
kHPCqjQe9Gq1L4gMC22HJPBwHoWth2T/iZSD3/xjMfMidgKDM6afrBxrq9Djc0za
M4cJ8mVw8CqLJErdGYTVko11+c8xjOZlJIPv3Cd0hyVzPv/lidA9nEMQz7eZGRA6
JKT6iHKJfXD0sN15uC1xMpastFRmsIUuJA+6pZfjxRJqL/3GdwSbp/7Ygahesi3O
ARpZZiuzPpA0XcpJtfABKyk8myDaBJqrux5oJrgCZEf91NMhuIgvgvWcMc8UDBgI
UE3jjEdMc6S0QZ9DAoMLqnhCxQTGaEDrtzvWL1pISSK4s7F/ClIcKwFahqNVt5dH
xz74i+quXejZEWbeigOQaOmcTokH+bN10z5ErsGGgJLHD6qz9V9kynh2gCeLpXVV
AdH2UtDPUFmSXULwTo3NLvKORpoUBVAPKNs4a0MMO+lOthhHnPcewVu9C9KKAQaS
sbndZoxOhNqgFBttPbOxzIwo9bS0xUK/kEbp5ZrqJSkgHt1JUaNfkpQo/Qax7BXp
nA6Umjnf3BZZ6YTVvqIGiz5gvdAPDNBsmSs3B/c85WS0ysvY7y8m+jKoG+H0RLCk
ROGqj0TLiQs9oOlTemu3hbrMbfDoNWTRdxSjt7rkNssGvrTdSbQ0PAc+CDRstGxR
HLW7Yf2JgOf8+VkyICgPakwaSiMCZalfRnGCMp5u/n2+/DaEoz4DOc0y6wK7TYwW
TTBlCDNMmJXXSIpnakyTSe3yRW6ELTcD6n+1b9Cy5OWmqtZURIb8l2T/c6MwmA4S
3GrV++CjyrUfI8UWVvb1KGxuq24H4mVS4uSaStctRI3e+tehqpE/2jfGO/Iem97C
JZ2pGkW9XADJx7J0uw7QVi9jlUbYfHJeuB4IZbPdeSSsO3N8ldRUWmNIBXyLuhrV
P4EcJloMtTREvHbO2mOgOup0smZ3ExkK5zTFR3iVRyAIcq/0OJB/4mawz8FIVjIJ
6VXA3Vxf0HmUD2Jxfyws8xmeL1bwUBJwGqqR22LyrtiKBHbkyEwpEsicbrXfg+hg
cLuogNZXLnArW4PTh+5+hOFJrKPBO8Zw+uk5Dt0niH3R04QSRNBGot8ICa0LLNXb
2EmtCUeirYkkKC+bRSx5D0S9z4yt3ldSn+53DxiFBmG78RY9JvxDSRM4YQUDrzkx
aRTZfn8qae5ekyzSRk5FK4X4+zFNUv1T8IW8IGv8JCEYlhlqmm8yOGsnN2lU7wvI
y2fY8gJX/4q36Ybqd3I0oDNmiXDxoqLm69rhzp+TN5KLc4nYHw7bhtzR3pKrC67v
wNcSpmElRucGwRywppE3EvCvgAyMP+EL+5BOE6oyd24lxKrCY8tkEr0ZfQDT4TU7
4Nh9B6ULHv0Hi91fe4Du5O+Iw6FL15Zc7NqCy2+rlSakPo/S7HXLLNb/DVIdHp5A
6X3InCQz3slqrThn/Zrc/yC++1CteqsJcdBd7LLDtOFOh7lPPqf7ugoJm3h4DPjy
0FjXbTdFKnMUgEkAsgDnEVaZKMxSXiVKFklnhFfnVigXW4vY/GeQWT2YaQ+xBaZq
FTMpmsmkyMdaBrmDXWmgxFVHqwoA6t5yORdNG1zM4MtEZEYDMFjtq7IsRaLOAKMx
ihAljs+gTKrLpVvgg3w6YnWF/NxDGClN/qcAnBz/88IsPHJN29qZUrqhCLYggiOK
iPpBRGfHAJ7W6zwv1cyO6QwF9VpLGoMs8asf7v87a5ioMH2woaRddqagK5hBY958
XfwGC30zyqMY4XamExnTgEdI8qXI0EnZszRr/+cNCK7BnkzD9YtzcBk+sjWLJMje
7FPegbKjilnVsX9w6C8RYHTqyy4EZaey0NG6jtMJOeD/9lYwFVHSG2wdIQEgnM6T
VOUL5rihhmEt2MDiJ/iLtBr/gwYsIwEbupGk4XvsinBnI62SQ73Ztc51PNgp1J5F
NVI0Ikq1XAQLF2FLrx4tVzdY91gQQyPXk+YF1bipS+gohAxc53ym1YLY+hxR8a4H
/CM5LL9P24u3PaAdvq4C+HrQP5gxhqhKBD9G8sRysKB8rSqbl+egt2XVmyjK58dg
r1lj733UvS8h6iQx1ySwwxHKmf+dcSj6WQCq3fpAVqKWIRmCk+Vdhf0kwJ6ztre+
wTWAtZBzGYmvgThLQvUcGq3fhpwWv8u6PPXrNlhT4VeqQSkhnea/BNaPGXeKhPrL
dK6ZDtiSYrjEgbmt+KmvlS4eY6xL4DV+X2AQzlxYnp2qxuovzLPsvtfX0Fvih7DF
kd/+jqE68AMRuNJ4qQxtXvFzLIxIEw3cM0f1YPc4x+GcWGdrc7QVF4gBGq/rqt61
3T/v6D33aCOFSvPYPTGIVrHfBpsafHLGLh3v3n22M1Y6vY/phV/MG+7ipgT1aF3M
s4unycImJtUkROBkmX6nU4MvQj7n9UM9gyY0Snl8tjkgqZmJC86SMYQ5AaXVVoa6
LzuRy9+2vRj4xsiWoSFDMw6iVvYqXDXe63s1RodDgHuwAJTGFQ2blP1oI6ajZUxX
MAAnHV0ejDbtzofo5yjXcvWzkl55+BSKbGGlt68vcgm5X/3XK1YYqdfP2D+H3HmN
XAFXn+RUNDVyQE/X2XEywmoLwvaA04AeTa298sDmJuO/9vIOekKSErwmsZ6u+o/v
2F8jLEnsWY6AQogcsgFMok+1KjjshVRtCwXP8uwZ5LZ7Kdv3jkPgVxR7SKCOgbo7
DZi3+HPWrjJ69ljIKy/AKrXlG54gAvU+IRuOtE5L/LxASTPiuQtp0If8VmHRuTHX
L9zpFLSUVZdP5rjz1o4PQlPuugykDR1u9e1Y8PW7fVJKzxpisqfgSdTy0ClH2ZzR
7v8nvVj9p5JZ2lR7kNmUZO7Nw1BtSfJDmBiEt4kF84EmG3GaHsE2MTRjdcZ/Bmvd
xll/Ne7grJR8MDTsCI9lVVkNRywT3pxwFS+1FEzBv3GTFiEV4bEb+HqnVypu95ib
gNn1PAwovfTCna24TAtSP+vM3BYm5VXNelpjcBvz4efjPgsx4HVfA2JyTe9JB7Tj
L1KkU4Phdbf6gq1oBxJlOr770gn/nPrY/6gCD/pdupjx2fpB1zW/PXSswiRv71fc
vbtVv+scEs9GGns93aZoeRoEAqtR0tdGWdS2r3cmaJ0CY/I7RKq7JgVS7/dBGRp3
cq+vn11p1EPK1MuLPiUcu5OElIggZ3VBLTv41t//JGc78Vin3qqN7mJ72XK6/6CW
tkiNq2Dea78TW2+vanQREXy3bqz9fgCdhnWqDZKAcxECz78BSNChI4KBaML8Ng+e
1XyR6aCPn8jjrVmXq/I3LJf7IVOfJjIkUD1aXIC/F4NO9Gg615G174pnlRNJ7Bqk
C2+yla4V7wxg9RG5uM/pdAxcM2p8fYI+yIO/tunK95+VVEV76Zvgd29+hE5FH3u3
xebC9Z5/c1Jl3xhoLupSLPQgqkCxyw8sMFzscItzQIJJoC7/KCtV/n0vkMw4gqEo
heunarEeygBL/zLuQIShKusSS0xGJ7PFgTsPwmc4088RoOHfBG/e3HpDeKjCi1Qc
7kpHnKr1XCplRXA4O0c+hUDkyNqGQ3b5jFl48A630DospfxkaIBkMPQBm8hKNeME
QKWhIh6xBn2oYrDuWBlAFHdTKxbS8QaqWs+a/jSFO7l4/ZRYBNZJecK9WWa1kT9W
aMIckSBXnG6k05FhekU/Ycsb0xdqHzCuo5rVYPX2ymSEmtzgi6zNZ6j6h6ry7UEM
F/yf1gXhk/TnE/kC5upGHSRsffMeVFwn2UBgrT6UPg0iUjB6yso2z1YAdcH+R6U8
lid3DpskIsmjJsmK3GxaJB//4AcZjAbQZMFQ8wC3RQaAZ1UM1KxuVvAXptig0kU0
YCPI4x50zrqpy3h8YDkDnkh348D7nwHtFYu0npGkg8KlGiHVHMLR4PfsERHbSK+K
5Du7WlPsTT+MAvfV7E3zNR3OFdBBQld9sqoywmujPbzIn2Afye1A2VTxJQFFqp8H
zQnSPnUg1JPKDdRyHm6Ig73idCleIKFiZM8uW/zSFxdm5WDledh4ppuv98/R/aZP
QrrFiQAu724ErpUhV+xxbWtBY7UuWNDPLQ9zWBiZB6sw1hxRy66jw2h+M72laYx/
BQTPR6tL+FmaRFABCtUf2dVg9zXLBY/tEYg8BADz1DFTjwKMYgsKRCfnp8+uUmP0
2ZPfdetNMepj3oukkFbek19BrIjG3Wub0c91/GcfkNtaeRxRVwbhzYFEmhLbSP2W
2fiSlrz7s0AGwcNTHft2g9YRMggmRZcfIVjzRRNj+uWaV8n7vzrJcGbFLXiWwlNY
kdPyrvy2OEaTq+r1PKQNDEtC+6XBUKOsMKox/WkGrtr3fPEQBPLANjfu1r6dUFEa
/eyrEWQ82/CZb8JPfT59YKy+s+ABtjtSbDvdGjzNnSKavYdXEUtNV+04xBPkhX0i
xBWlUP5VAfaV9OOeYrT3LnY6UumQQ8aaQNY+9o2ygGZhT9PCE1xIbnpXWNXFqhOP
yzjYeN+oiGLcl1oqpb6/HWe39fS+T5LanLKsS9ao+7Qn1XG4KqWQGtwgXjsQ/7G1
uIyOSk/Nxe6Q8wazIsGzsquZfkHHVrQl0UAp795x1TjeQiLnv7T4h2jBzgDPxLtv
fZdxei9unAyKXkqwjxKRnXvZKt2QqBbqX4I/xTeJp8x5bSpi1TSDj82hD2H8NUf5
BgsmL95bKVey6svE33izsJbrtpCR+vt/2X2j/00lsbO6Gi6QkjOy3RA562mHSv/N
7s6Hs5XpGoG1TSW1M61+A7BWNFV9JYur8pekRSwCwiYOaHhK3bgW2f2kMEMlKtjl
3atZDUrjaVhMm2If7RCxFktvxLAWbXbkfARhn9ZIw/rC4vxODjFZD3XLXoOOFZkU
7Wd6d+e77XiHD+uKn9uuFW3fzcRMyeuZONgnP5vXPcqbtDesHhIvVBucReMomaok
XDyFDFsfJ66ZpOb7Xt4KK4P+ddO5qsAk0y/S3jRGdpRJMculKD1bULbQDkeBB3gf
5fOZYyD89AE403H1g6OBabTaKGkCtZ+7uHsTJEPmwskdBXUgublNQELlP9Q8I2oV
EYN8FZAWsLCDoKgDntJ2M1fglabkm7EsnjsrJ+akO88y1en/c10yvG/V0b1TI6QK
Xp336AxicN9hTh2gthAOgHAIFXUhGHiV4mF4c3bx1LmA5BPdc6ya4NgI+LQj7E9n
rMQvj3c9bKI+CN58yiPrXPN1DcNJvRJIUgE0x/Js8irv/53K+FHAPha1h+VkyU6Y
qNYTsSim/me0N1J7ja5qbZvVSaM+NQRBcHV7TbYYm4y2zg9mDJ0Rslm+Zc0lA+Hk
YnwrxIioUIxth2w96qhLog1s1Jo++TklMaf5jrNEXEH3tKevYuh5EiYfUBP1yf2X
SMpKDxYs31MJwJ8R/lJc8bac6ndoUIHFLHJm/R25mneIhuonsN7mnAfcTvT4W/cA
pJqZzmleHyUbFsZnCWT3Xmg9hRDsEjRDWVLfyGoaFyQrD0CYXr2mbBx+eLbim9hU
p0hBmEoOdAW8JGy8ZNU01L7R4uuBrPIjUe4KCDeVv6MiLe5p6RJInlg1Ebjzo+01
QyjzG6lXVj5xLO5ZzXvL0+JZjXEPZTSb+tdrhwXZYaLTN6uoqyikUauEg3PmzkE3
/vvouQgMUl2jqYofrZ7oBK9NWBGWCkkLmHcrG6JCCg/Y1NiNsrTYyBDK1cw0ktE2
AF4qrAzpcyZ4Li8ZN/Bci3xjhYdsVPDEH2PgQilYg/UM2lWyWT83inO4N1vCRh+7
0woxdp0cy1PcSS4vrbvYJ9HrI12zj/blxHiMjhyFqR11+Qat8X75avMtZLAduKVr
4RMvCPsiv6bzIlhXc2svBKB19a2faVdxHczIlmvU80pId6w5Ih3J9ZIFZh3VpEsf
0c+IDQVHnzAEfL6bycx8pz/AxnER2L28+wZ9UmSw7ceYZGlYSaY80utrSMxvYYx7
xPohXi1SGJFB3Tx9VJLsYg8bhUrffrQ/4WXdW+0eWPiLN9Gc+yl0oVfFGXK0/cqt
e/OD48+NI4vpmEnpEEli9PDkj6OnrmLYKyTcMudlPvqnOtI03hlIbw8EgUFu9sUZ
EshG/oyob7Aw1UbtGjs0RKQHwYBRwv+/VrlhN+e8tlXLRKDhDO3u77gQPPUKlUPD
NT0bZyaMXG0VVf4YwQO+AK28wuy45i0iTI0MEWt+PIjO35drA/Ll33jxYc5gZ143
gs92vZ53EZaZyo5ML2ST/yQmFKSn7ocx6OsY5oU1Q6TNMz9Uy/q383fjk+WSiGn1
vyCFMmdHAI5J7dGvlxB/hfW+vd4aUrYXlo4BdlFNfXoEpkVOkNtvvfyfRf4CxxPD
0hZNFsxmPySUsWWB1ezOxF4iVhb/xQrS30vE7VyzUnuqthmK8rFjqkueOdtlOuLV
HTqpKBbrhnGX3LHmnI0t+luF0hbieLbcsJfvAXTdow2NyNx0iUZcni3acBfAATAM
3z/gUqab9kBY2yLjfvQdWlEZz1AeHyBWCIFKw8BjXpB1pDYZJRvIY4CUyC7O7FKp
0o7DjGYezqNPQdsI/0VRhviRCsOFt8QFvTZHH8kL0QtxEA8I3T2Ox0E8QIhGygXA
/N9lq++Bjc62Grg2i54Lmm5h2gfPiL9hjNc4BkzARBV8UjxZO8Hu1lNRutOKOk2m
tV6DXLY3f/tEYf9iNSmG2gtn8rEfQ/CNaTIDQdOcOOp+u83GvhdIE59GjT5t1svi
7c6QLZ+8pJc7EUTv5118yeYMpIiJ50ba7pPTgv4CqXBrGzQ1MlgA6jIzZF/c9Uhm
vm6+UKZzBKIelgsI9L/jpqrutJ9F63tazAs+nQYHuIegoNsxO57O7CBKLB2k15G3
nwqUuEQrrtWFSrvPf5NokIQAp0cJef/O4pT1205LbEwde4rsBAV2OHpyabppcJfu
v5U7WCkm910JnDQ9TmthsrG70SFY0B5vWrwOrF6SdIsrF7ULhtLwVyzU3HZTuntK
I5i1SdtwCEWNx6A/7tlPRUwbU094g7QI9wjUrL1Fb/krTDB5dNPINDi6DmGmENXh
BLTgZ4FwBKx0Nwhczm/V5ZuiFgbYeKohcRjhwKwXHDxaR31AXm/SeJ434mxwFCyU
IbEXMpP1Zus8UWclPVlNz7t2WiwTh+QVQoTH7P3s3hb7TMeZQK3EUxdet12ePt9j
h+whUx7XN39NONBxfxjZaxcNHUhqiKpuxt2Ry3q7snzKz16DYygIJkuPCqL1mrVc
W9lfHqerz9BwxTh5SqDdpoq9ECr840nxsAKauPROEY1YMEGjOMzlPvMlo0V7I45t
70t3YQt+UT2E5J4LP/G19RM4SzV4yMheRSBUqbfI0hiCFvMxOxETdRIfscdwBtzr
T2IdSWloF2gCnlDBKknyMD7h6qX6uWvH/CvKfpK6g/3kOULyA0dt2JKU4ChO9nIh
4RKCR0hrIoiCT46zydblb8n9Qbea3Okrlh/0YO6xhCG/N8dc/j0NG5Qu+HBEYHTv
w6W/aAeaV5XmpafV+Wj6vkEf3ExcNx2CeAncFk16RClDL4UauWto11H36OhKM0EP
PrL3UvNp6JyfeYg+vbz44OxoAhh0tO0L76lXmD/kLTPwrk/E6YvenMM0WMkGhFoe
Ej+gjfD0vAZCkKH0CK1f5M1ytEXGiWT20WodnCxgL9u9QfmwqyAl+MzkHEE9ByLY
gdKKmva6HlmJkw95oa0NIw5l+9bOn338iXJVgqh9ab5PgX3IQQDtoYUfbjgZCjVJ
3DVC+YFsUX+rBTyBCuoa4tkEMzbVC8lY4LZRedkEGwbdo+JeQubaLPaBOusf3wnp
9/nf5xFZUPLT8bLXPxkFADLfbdYDImHS3kLmp04PI3BXXyEnB2j+PKw9GgRdHF5U
H0IZGkE5ixln3ybuWgMZEZ4qI+QdKtKyq26ZxH0j3a2HIPjUdidZhBqgXliqEdOg
ho1drUvW39pPKa7SH04oYXc8KxCVsAZzJDsd7m7ynW5KGBRs7Wqg56rbkqtoHz8T
XGM8NUGdmPuF7Lm4jdr+yygALqOP53u93yLohnV/Bcfrxm3uuqqKg3um/gTcBS1c
8ne/HTt8Qci5wJ9S7uxvAM7BcN27PeORuewa6VKdNEX+zLPRiX+s9DM9YQV4/Eel
auEOiiZnmzBiYmJghFtrp8yCtsqkG1zgyd6lx+7GNgMfw2FDtIF/csz9zH0LyStg
xQH64ptnILHTLz+Raem1F90z5YzWPw5ZNzkp9SPZDk7RJ5Bd8Txcf1fM5fxSsNie
tfQvtqNXkBZTJHZnIMaHXXwT0RdBqm+s/Xtqc17FvIuA8azWd+tTxBLmRg5WFtmA
8EsDTaeKaGOzWol2gRrkPElDBLDioRyeb6Cg2DJVsXrZg7A6i4t0cx2TFd78mZjd
3xrj8/QJWgTZOwkLH9ljxMqDMJwNRc01QuBkUt7Z56SMIa5UQg0AZUiAmW0lzeqP
MKPYmXkysn96B5v/+YdKTZ4UEFh7ihqq/VLzKbVXHI8ukqqs2yzIBoKJjRA7Ba+2
bCEHtUxAR1WarQww5TLrl90j8C8SqstTs1dXme1L9j0luNJwfLhPsaQMcYUhHRkX
ahaiD5wX7Au4SE4qVeNvxkMaWXu+TB2mdLaHttO+TSNqMCk75tBxVZMqRmRKzi3P
PqFntl9Y8DnrYFvzoJNBWmGWWMPkorxQvjiqPuwq97rKQFoFAu+KdU3mN7TvsWeU
/r/Y6rtvuHTZfjBj7x4jRh1RhZaxdj516RBSx5O50tE/dIje8GwbE8bQJeusNa5C
9IpI5teZ+jpV2PC3K/ER8eDseVg9NILmuDmWFXF5NEtLDkzS8cr2hHNMY/tenqMi
Ce0v4rmVf4Cw5II3EqSw9MdDd66MfsruK9rm2H5erFEuBNKUSilko3B2W40UsSOp
NQ9GPB0YLbuinvvRH3yPoa9fQIV9d0Jr2ZPZNtaeLFsNrEDWF7CTJpEaLesTezEz
HtMSMN06cH6QWFzWb1NMzimxFdxHjPw8X20BvjK3DbV8QNjpO98nfUlo4ubrIN2N
O9FP54hALj66Za0GIVvQ0LwWgCt8sDDMRfun0+2G4SZhJU/MODYtP+fQz218TI5H
Q6dzyLSI67PMejkJfL+Jr4IU2PsYr0AJwu0qEva9rW2BoSt1+diEQR06qSCTGxXl
vuT2qgREcwDtk76LAu8+UnuryIyIntNLMY/cM2HWDd5THe7D88ZV+ESDXCrDIPKP
2l74n/kBHvY1JHNEXGBWIL7pBd0sel6vCzomTnYlclxjCbnnbjsX6wvavcFsNfB8
IBVa9GshgT7pd4O30vabXpKbhwq2IlR+o1PlN8cgNk+tGBMZj+nwQ34+f9E3sWo3
/+C1MplV6qhQRUEK3MNUH7Jqdhf5xA1QktbA8dSodQtMnBZLTADcrdgz1OwUe0/+
xiHVolkNLURjFnI6638TzFMzbbRB3+dsyfI1FzKoAoI7lJIZdvWJpv+T2dJGoQh4
aUZM/fjlyN3YYbitscpQwLuTeL0l17wxkjYF4GwGym+v/kjEtZ1hGdr8b40fV+Yo
oRE0CaFtXR02PQqJMLFAuBAUdwCtGBU6dbguiCPFOSR0eXJiJanuv9NAljECrbcF
fAyaYpmOx94wJvXMommINfjNacSv1n5WvvCWev/NxsYb9ZVJKOpsZJ7PQ43i0xy0
2WZbxhQi3YxzEFkeLN3tCLH5Uo2kLStFq+/yeblg+Yr4yGBLicJTP/zq0I4CfQhM
SXTfwPwBlT7Gol30sS+Rn4qIZu9Cynt6QyfuWs2T9BrzKpKVdPr1KONEmvbYer9C
359i4lTc854RQb/luUMBoU9ZOTWtuI6f0TB4QyV2uhGBtW30QSLTSZR7QZXqh5IG
t3CTIW5r54ef9pu3M7JTPgpUHNPT0BqLK9UIQnOoL3QWyhYlnNpL4/zyQSIWV2p6
9djJhvZhKjW65Bph9yV+4et7+W5TDwN2rj8mq8OmmsbfHlQXM+GhFiYewV/b+xy/
eP0G++2Q0FGj6q4Q7tmF6xW0NtQIjD9tJvezdCWLMKXFyDhgECo4pkbd/m7LjGvs
ZNTgOFBEfxVSCOWyhP2gjjqVMni8nltH+vjOaA74US1AKPlQsai2k/RaZK+zqk8X
RZbdxuD/ZXEpuR7hyRZtIM+wct1+U5+0JwfyH/Ks+snrxnC7NGlal9hOyCl0Nbam
7TozL82/7rsrXmX6HFCHgxVrL+CLDbhOvLSXImvoVz4KiL/CNs2IM0DdSwaYqvIg
zhQXQMdT36AiWt5sbmLpQZuziz47B5j7KNAulyA382phwDSresex53AM4DKr3B+G
v3oHgQzmfeXrn0Lu74SWh1AMPG/me8aMNyMqXbQP44UYYZpsaL7Jf+hsoNfyuUog
Vpol+VBUCgZXrqM+n74zW6+ntqQ0Plqr3PA8QHyqb5ZCjYFUMUbf+7CL3ik3rRjv
gU774VjXzf1weklvpLChYoujhUIR7yUvPeXcMLz4yASicBrIAT3CqqNeoTV8QS+b
sU8yOEOlbhazLnFoGVqDdy8LwxGYVApxLCBlZC4ga8dO6YROkbemsCe6ofl5LfSb
soLgfUpmYDVzvFTQ2RHk2qd1Jb2/gGFdoOUyQxt/HODbGmC1iQK4l1NDgM/jkkJM
FDuauBYxYb5RVDaMGzsEl1ICOACY67eVxgnmd5gMhOycJxV1MWPm63/2DFKjVkF0
GHJqi7qm1epYe2TNj+sLDsSQzt3K62XTUAUfPSL28l5RiX5oQE2Fetw1pr0AETdk
G5+lXlp+fJH/CHRFtg9sSUoeF+C0EjSihDBoWm8ruYw0i6tcXPYIR0AGJwIpVmXS
cJ0XeUD7tojCp12uV7x99hGSVvEy/vpu/WXoFxUqnwT+vWpqXD6tqzSbspRNRv/p
wRLY9F6cd87Lbe4kmIE3/VImPsUJj7w2VbByv9f0uR9ugwE43q1xJ7VEs4ejrK1G
BqUARqNv5wsK7LeS0gZ99klzDcOTAViWKQxdVVjC7BbcW1QzAsKRO7oMFlInuDwD
SgpBksRXt9hV1pa1poqLKe3ZJmL3wDtc25BmTVdTOfI3J1xTWw3Cf6pV3faEX+I3
zpU0aYcxL0YwQ6J11zsINgPJ30JJJoFRe3TTbCVSPvIEMNh1xcjkbhn8GqSCrK4s
IJqcjzbISkEnoCa4tsrHq/WkXQ72QQ17vAxfQLJe93emqWuT2trpuhPO+AXGJh6R
5SWgTjgOCBtIJ9h4ZLekMOn4FJYtIcFhQeR3qK8L72L8FsHqSYxBwdWHF1gPe5aL
cukVrpUEagq1wKGkNEszH/8ICs2ONm+8Z1hsauI9dfk1uIb70uc7POVYrqbXPf3G
tMKynvVax5Rw9MZ998Zrl1wTCeBFzLVNngevleoQgLJyJnBtxaRe7ycL8mrL7O2m
oPh8bUH6n2GV6dwbZDmtW3l587MA4iYsmoO8OEJP9DoBcOvimot8lsFx6Wiq7suH
Smrg29boeavDizKLFSaG4COaK+VtOVSxvkVh36BWAUtBf2iZ6wTye91WhiVR7iJA
ZuKTJYvPIG/s7tSzB3sOm5YQY1UxVTgKR6t3nhYxohFiMmyZ6wwSQeytRPq7+t/1
eJRNdlqioeWImZG8ky/NgXFxASj6EKg+x+8C4C/AIdSDnpmUWQbwzOVq2XDsm8UM
R3oFnFE7OHFfAxx70apJSq+eJ0xHvaOCBYo78kczZe+riMV27z8Jo3jkvubse05U
F2ijTU+69WXCqSgn7Dj22rsJREzHuHS5YXZhdCTRlT/8YxLgTparmrBKuBGJU/tK
YrcMnEi6KE3aFtAkOjSFsn0RQKdeOPEDjg7SAPoBL4SH9m4GaXUI1FNedwKXTn43
pUdYYXfHumW5u/ODPLluRnRmGtte1pliQZSHtbfpmEFdpzEkKRZcRzrxJKhq0Srf
5MjIiD4WN2slf8eLV2ps8zykSAWT+w5fXBBWQ6haLUGleD0oZ3vIxmgJ721pMkZ1
CLQnkkQqG3vg8P3+8WpnLvSkG2F/R5gwDgPjyL2KaoTX9hbN8USi4emeTJ2wCgUw
FX3I5EC7SqaivmT6KqyCuCsKm9LmcW235Aj0bEC7ERgxc29Jc47BttD/Sdbzbxha
S2HJBvB7rLnVT/y4pjbb1u/3kNMg4jpNPtsioveiohwTc9Rq9MZUQZgTiNJ/kovy
AYkO2gp+KKr3Xkkfp/qtnXQfePMaqGrxvDV6eNmP1AUMcXSmjxXNwmkvYzboa7oy
xaknTMEjw60jpW8N7ntiHqvzWsfS7gqa7aDb7DELlJiqVjio6ciEATUL4sWRCQHy
x655zllUeE+JFHpxbfNBeiRzeIA31bl11oJrKVEbUWIzgw96Hal4IxshDrPOIjtn
UWPA1diS8/3at5wxW6XHmv2RDugK9a0AFK5YWeyOukcGoLgApvRdIPZNVWL8DBuz
K7fpInnO3D6mX7M96l3xU4uGHULhL0Xjfw9wR2E7CicrMm1DUz+cq89HYzmKcmaN
LbLhx9wfh8AtF2jW8yH+SUY+wpEAjl0aIKlv9uaPeAdqgySs/EXz8PLuYf+lWuns
VI8nWh8d04QG5gl0PlFJvFQx53FfGW0ANt+lm+kxubauOtdbArYSGxOODSofL9OA
nIo73eJaFBGFNRLdP2SHdtS90mFNlXkA+mYiGcdqW3eb2X90TpL1+PHPiaZtSpvt
SRtrE+pP0a5FNPzs7OVlsUsX/lE19EiplCUfDRMPgsoQdOsEOBvcc+eREGjPQFLY
tzakXfOTQ7b18x3qicsYPWn7LUpvI0/LQkR8Y5BhXd6ifdlFCZIGn7KyqR88kKL4
2mNo87uhvNMe/ltPOHYaNUcjU6xwzbBfmJ4PYwJ+MexXXjBUppAP79rRxsYV3koZ
JYSPQr94dENKU/KyE0H4GUv5HoVziSYLzRCKkTGy9fYJ+LS4Frq+zCQGCGYaZKJZ
C7chQBuEQX7x2iju3HtBh+4upChldl63HFHGCXIrVYaNIJjejMoLmid0NOKHoQk+
7gZs8AVgiwZoRVE3nE27emnecS5qWzMrG9utEoZvVDvL8X7aUv5tU/C70U9/Zx0e
YunT900NRUs8yfVAmnCPxFla/OCeZIAoOyFND154shlEpjRSxoPX11oL/orJFI8X
hYZlB1DCRipDPQwfLpvAzoWEsYE0RQC4eunqPt4E45Dlutb2G7x0p97UOUYWw9uw
YQvmZtMyi+UrBOr7vTTGwGQzajpORs8S3KZF89xdHBnEB2tv9vUp/VSotam4SCvw
0wKzXvFpYuohvRbjk9Jj4qCttHzvv6asGFY/4EahEy4yASG6KyePYP41NtJWMFIP
wQFfiNWfxyKalu+5/riNhRue7GFp3TWomPSFdww4x2mGPImt50E9IeKz4jL95z5L
ej0VkigRkE+0y6lX05hrIbA7M01QqSrzGNqmiTicG3MN6q2NQkc5r1b6CH9gSiPL
DSwfDKuuNSnp7LpAWyOwg31yBM5gSwNu7TaQbo6TUO/cjxPE/jaeYwP14BEtatgH
QUqlWUWGgMzO/fCa8as+b5TWkSAKntHYczKmQ5Sy9exfzgyMDP2yCpWiAMiuFuZ/
zv8ApZPZxzxBQqrlZs3DkRXJ+Yo+TBp46m+Dkq5PUTl4FlOoFgl/Ik8HGcDONzb8
wOczp2R4wLYDo8HludxisFG+A2VKLjzJRgiIQNplZ7//JY4bZfhwzS5EiisGIy1Q
3XwGBjRIYtlortsX7sOwNQ0T8QIx1raiSmVtge4p5NTu1omopmGwRqLON6syg/Mf
90X4HDgK3mm9r7AAS+pd3wJ1B3NcgBLrlATDT25Gk5bB34abUq1PKFsVcq7wRDoh
o/yizaRzEjAqMsd1WGUWiTnQJeq+d2o/g44HytRXgDLYyvUHMGDry9IUVA4PmLf4
knUk5Xe6vAvuxnMV8NPFOSktvCiS5cbyXK3K6305q8FMpImxQlWIs+2CC7RkwD6s
swZJgzT0Z3GMyEXa7KQXLQOmiGYjBqj3EYBpCuEQmqXq90O1QvRhCqNNIgEq8TT0
NmT9QoETNP1+P5jWY3TPWlqNUgDogjTJYKGIW2GCRligXy7nyBNLhf2Z11+1JdK7
z7v58NJLVCOuXbVsu0mmzFAE9danYN2t5nPPr15Ywvy4SXs836C6fGvBfeXU+nsy
tKVBLHOLj9rel4dpP7rCCc7UuAU9s88e4NfGU1DtIx6KXPRzUkYhCY50Dtarrulo
rbGDDhZ1shRUi4dlV+O0NmILTVwSEdm7RjDNz07grh9jIvbr88smrKCkJxGFYnn1
QPdEo18SvELJ0rdVF2XkLopmx7RnzLg8zC29HV44BourqtpFIhix82NL5203YQfa
KRTB6CKPSmqBIK+P6VfvJKuni8EApzOF4S+oaW7Nq7g+mRwbxI9b1+6QS1O5s4pl
b7sQvTvW8BnZ8H6JxhTaEcmG6srkjOfYXcwoeh/wJw+Amnbclb3vLev/SsXf0gcs
KbvTumT05DIk35YdtkcAubjz0Wtxfpmnvs/gcW9wuuDSXwXrk8PnC3EXVlZSBjJL
DN37RYGIXMv6iNkKMzCXuBi7OT2ut42tpIEKXaAZnhg7NTQczHeGZs6kDex2NjQh
/BaPBWubVkrwRFZ95kf+cO75HG7QeD8QsmcX1swtWqPXY2dmzNqFU8cUGBd7G/+i
fsGSyVJdlf7tpQ6VZHUVipUY1fg+vf/dI6VXgqeShLq0O+JHwf3nXWdNYWd2HQky
kiEoJbJcuwO1+C7zMPtFIR0dOdbDZXxlEYV3SEkmyBP7W8KzLg5rU68SdY2xMXBf
bAAPTLNGc61lGFK6pUpbottIixNys6KVoQTJJTSyyvQQE+aqbPA0rJNTG/XeJVSR
F6ThTfeNc6QzCQ/YrREbKuJpi18o5VJtxyoPblpY5ER6gk/4nwM6xSZUKcHpGU0F
Ub0Z4FdnZtYwn2PYA4wtW5JDlKc5CflAmDi1PWc9vjqqQ01J0efDA6Bb+K9T01vo
ClvPymv1f4WTvsyfDg9FK36hyySHdydoI8+RfzhZ7uN58wu9Xc8qGmH4CK1+cPE4
wBKzdOmVdreqppdqMvs2H/0DsdSwPs1T0CggPq4yIVRZ2W9qvAQH12XIH/GD1eXb
oxqm97y6UV/nT0tFGsipGaQnZfzAzRqvChFwuEt6SFyfI2IXygZScyfgrXaENh31
PEYZHnm3vNIYMKiJ7jQ0odWKuA9BcF9XzeKvaUGZEN5KrV/P0F5bIyGsqa3BpOHx
PFzve6EuxhI/BLWheg99SHefp+MsylbmmKkaC37Ke9I7qBluAgxdJjayamLy7vLo
7Xs/hPcyMLnxP+R98ga2c4bpxivliaWbcSCwovSPVDIeJVn6MH5zwBfzmEaAWy2M
Tgc6ICySEdKu2w5Gsj3F78JOhDTUIPzU1r9rjF0zh/RCbONgKo+Y/5z7lIFpUY+l
+T5Y3Ur3IC89ImZAgi3NwLWHeS730R514paNicB11jRdWGcjzTCRM4yt3yvT2lAc
8gSu3X9Edw+R7KlMIRzS8kdZQjv3Jvu6LGKkg0UqkKtJIJE6QXy9qmCvXgRm0mX9
Y3AYnQ5Ev+ejsxD1v6ngfPGuvN0cl35KAnqTqT9j/GS7wkcTSATmD4YkzJY+TJXX
Deucr/j8UWYFfZbvEZFpz42anNuwAGuW/oltA+jga8k//hjT/hoSjuBHtZATbKCA
4+3fPSbWAwTGWDuylUsiHXkyEYmI/oN9201HuzHrWzfjEtnbji4TjwN1B/giBPDD
KJsedLfFyvYwhvsdCDsR5rbGP/qslXZqm0vj0NORVf5YJkGQp7bnTlZDyeVf4ztZ
yzymILRcL8zHuab6mWEFeMRzLbvRdyw8jfbJdFYBUXWfdS0naSmyK7cQtzeZoZRm
Uqklt0nVuucVISO4J+keQHnGabFfL5WeLZHQFxK8Et3muFdJJHJlO3qcdOcLWYWP
52z93CCVoEYsZWpCDAE43XJYG+oYNHE2lOex9Eyam1Dd6eRbDyGH1/m0vQ/+Ky8c
/XhJNm7sYCblcN68oj+FAPKUUrhrhwzP6r4OOxm0yFh/AFYDmNYAwTdZLsnR/4ji
2fywqtUkkYyFm0OBR6lFr596q2rbW/maTtSkhfybU1AXNROIaqQpQdR0zn97o3oa
ylIUZn8a1zpsTV9Hj8y467hB6DlB9z1USGAuKMNSt9SD1qF4c7Xtjl172QKthii3
O/WbBCCiJSfH7HEA+kcsKCG8l/eB1dP0fIteybke7NYw3Sbwxl5tN7NaIPsJvTch
Dq63J2wND3kjO/UEg0eJW85PvSbvahmGLXdR9R8AosrE9RQGgyFqgYQhdYEKwwRK
htzujdpnHpKcS23ZAozGTk/ds+XhDmTRhTHl0ezNa1Q7doPsmcRvIFqLSvDnE03l
+bREYDHl5UThFfkHlDze1hO7od8un+swGUET9w3RHASAscfurYXUDd1678J0BpEs
u7h7e4eLp4U7Mox54v1N6sGsOrZLeThPtlpjVjW81j3clf3e0mz9StQHvHFPtIUj
k/ifSSO9KcAFYLNqlvLX9eZYga5YqWydYUFLTbLGGOd6IrKiPXmN0uAmscxIrqoh
Uuv9rzelBdal/omHae0/vARs1gCpvp4kw+GPEwqmPlUKl0L110WRnYZ9CuATWTr/
Ze/aWxZUwIUnwDvlgnvdne+dNteBKos+MiDhUK+83HOjbFPooT7qk8iJqVuk5u4c
/wK7vX4XGMQuspm9faul2WF4ItVpr5Iv8pJUBAC2IGzdsMah0vwlj+N5koQxBXAN
v4GFjHtpi0zAyFfEDxNYJhlTuo+ee8FVOjNpCHPiGALXh7QwiDBPpIPDSQMLApqr
MODekQBNsouUW+hY/CNYGzfhg5RrbcL//f0DmERCC094Kg0K0V7KrSL25zmy3M8Q
XZhvDY5rS/I4rE0BEFJDp0TwISuMNkwyEYcWxiw8G7DGp0fp7MEFNWujhC1ioiII
+gzMy1Qk0ISGUzBvB3lr8sExVi06gH9uImfThiZoS0DC0oBWMypQPWW2T9R11x6F
eeTGOkQF0LoRmNazwZ1088pzaqu7Lgp0/MuPju8Fc1TPbVELAamVluYLrf6qMCVA
musoKqFYBsaFFLwR6EJEeJzxNJAc8Mom9l0pceonXhNUXz9H41my5NY0kiWrddeR
E2xSMAhGzUIwvM6vMLNHcxC+CQ2Eg6gzydydeSOfbQ3HBU0991BfG4IChrY/WKQd
fqZKbFy8PVi3UYzaIZabjrqEMm2O6qpD31tj3lbBIhpuJzNCKs2W/NWk+cg/aSSB
sX0oaH5CReFU2wHbLx/yIwrcg/+XNVklzsy58Z7WBq0iKcaPVrFDhkqwMjAiKNfK
O9NbR4svcDQ/GkFzfwDjt3U/JZovRInnoBjfC8mfGIiEiqEatL9IvnvbDYfbWgAO
QskPldLx2m1sWLKBvj0M/ROuC68cWN82V6YiAnjis7yv1xMZ5OTtFAOmvfEAQTgL
SBtdoITTFsdEbw4VlYR/goMfoaixIzt5J5sXtBi26g6GRawq+zqk24PXjfg2NbUl
XrDNrih6bSxKKFvLXpI2YCzoGQ3rApM1f7/3c0XrV3XF3wVrfKTU7hIlu42z6K5Y
xemYIX1qIHn+z0t2lZlrVmiqezwyViimbm2wnvP3+olV6XiEiaI71AwM/ks5pg//
WcVLuG9ImJNYhtwRZhkWyWEGxUu7Z5IKzX0v+vwIb0fzCjRmVAAY01g+qXJhq3GS
bLahjXsWoXQvLDyjztLY1J8goiYzxI8q3g4bUaKBQ169zlSi2rxF5BQKGc5KdsB/
AECoFii9U7OUjq62TsejiTTRLi9uEFaZ4G7iNFcwU1FnhhtXTrSev5ZAzj79Z7Xl
HyTf6286e0ScWbnDb547e8/re2YpP9SVay/3g8CqgGtAn8Z40UIKn4NrkC5RXp/b
amEP7XcDyDVKmdpnsd5MnCH/aD9O2lmGJcnxE6vhuJTTFX35d4MxTEb0lAEDx5WI
LQkoMhkJj5VrZSxihRQsUWHs2WgUb/zlnDW1plIAPl+uSCgXtfi1v4XdSnd6fy99
jWa8FnBJYU9ZL9H4j5rjMwRDM7DR1pKzhqYt250XBeLEUYY9rVluCCvQaZ5cbQvK
rz3GJERjcsMoLXpRwUAOMx9tbomTCaxxvMPVESDrMA4EkIrDAWvaux5DIB0O6hXe
NV8ebj8OnktBIWWCab1LjkQy4zAROL3MEacaYfmcEw31Z4r24ZEJDA1H51z7W4xS
w+lTb+8p8szWNS83zSInSK7U+S0Eh2ufGy0V+wtYd5hbfUCj1IAN10/EdBbCCV1h
UUz8NKcvyDBxkoypwAGBw0zXzwCXPOW9lBgir4g+AHBTkyNQdR8aXrTtKvfMvVHN
NIg4Z2t5wLc8BcR6dy7Psw72T8BMUzzcy3JXtOIoGA7W2GofV2uVHg2BBKwR4i1E
3Ny0hi/mJpgyte0JTbfCosCCqUPWf3rN0c6Q4Nk1G8PwtFR3on35h3nQPJtDtM9p
Bc6GRt5y+e19/LjaxxpPaySpKSjahoV3oFjOcnrjU0DL04EjFRKoSgdrnUfDhC5g
0RJZf+BtUJJjnw2ZPqx6XDmGx14D9xLP7CrdEgAnmpNaGSf4UN3CwnEeJnLZJSM2
RBenax3AQi1Ql/QoubSC9XOmXKfPoKOvoBeSRVzFuZzfSnZix+IlSx5J0VPU2iDC
bpgSLTBRzJm/chKUwq5aEJUG0xsopXp0441IHdR4/nBtCcdF4tc+XmFEX6+peeis
8YhPOo5uwurk0sm1H1RJBrVpoiWsR6w8NIJdwnjFCwaKqO1Xr+doeosqv3bFsRNE
l69i4HTCiFluFzzjEBObEXJb6bm2mEY75Sam0NZ+5LzRvdMxkw0uiUv6LeIV1ZPn
z4SxY3tdSDfgR2kHGPt3rRv0nBsdZlDHjfDbc17aphjYSc/6W0IwOIbUTWGKSrh4
wRo4ftDOHH8iJow3C1Gsbs4YlCLUv674nhHJPtdvN2FFFeQiKYzd/2R2pcSlg0Mj
piqe+LmpXd9yHQbG4nzvV4cEHdkq4n1tdP4J2NGAYf/2Aqokgvne75NeuQSU4HIb
Yl0OjyjNi+1lPmQB25eGrwmnKf+lWxdGsx92/5o2js5/Ysi/T2l0HApHJCZpMcms
7CuSejiXjxATD/1DIpBoodnpx8CCOTGOyXTmBo2lPccshpbAxS9wtNsk/o1u+2JT
8Xmmm/vqVG6rpxi2KMivwp4jo1MWF6/IOkd7cmStTl7z/iZy5QRUSuEPv5abqxs5
yAD+jLoIx3ttH3Ov/vEdFU99IoqBHSx1h+KIKLL4MZzFFB3Jenl1YwS49Qt0JIFY
d9Z9Z+I/W+m1RxaZOATt/Bf2+EGXgCRQhjtA5EREL2g3UR4AQ5sKReEIzaNKySXx
UgNcnNMp4VO0XqmqzBvQ6WNpFWy64s0JM6SWHWgo7H5uFhXutOrd8TOE1X+MAJfq
JIa6IiPdp9LL+aCpgh6N14u9CzepNzXutId99+639FZgBbeDUA3WrjjSlni7GRpM
94aUSOKnep94Igt9nrFdEJJ5v77NZPyMxZzK3sT46NRQF+i5xhpIETo7BDqLY+ax
AJ8F0jmAlGSidNCrB+iuaCW2XsSNZ3qPJuF6wTrtt2bhp5scSoyR6UmJoG5bSopv
WrUUVikcsGX1dY2wzH5OhRt8pNf7EloN3d/ZIiWpFVuj9HAleZ+AnTVjO0dPAdD5
JZHTW638ZBDk9pOjeyvB8jKQfUoVioacWoszSwyXN8FdxcDN/GTS+kO6cv8+f7lu
v1DhZ5XaTSgBsbsG2a0/vQLdUsOzqmnggQUL76vGI/UaPKe/6SKVSGyQT7ISeJTz
Nr0jpSIh7vjSdAql726gCeJUzxdHa6ZXqfPjxxKTZhuAwN1wkaezqVo1mekjoQTk
wUzZp9QuuyBCEi6EUOufyb02m7GZj1uZTT+tQrXponFpgUsP4yPY4RdDjzt0jyGo
eSEfjQqKoPesGY28UPZJzGtWtoz+6esF+RitQ5Ysehh5sWTNq0efzAstP1In5+e1
nq2VcyJeeqM9UnK1trAnGngKtwyUs+JtyvXE4pDIM1jobcsoD8CfzsCXcZULhvj1
TmzrkjIk0Zpx8c1go97oVLoj+mkPqU4/Bt5XFUWXf4Oz+dfE8hnRqCFx6JPO+oUp
mh/m5pTG39X7ni2e5BbSU/8fQ23FXsaQ2Ks6CO9wbvNx6zHzSGptQ2VZhuZpzWMi
IFMEV+Tkf0EAqG+j9QKtePAjs+dALZzcMXGM3wgqrdhnDjC9tUwt7UcCeoE3JelS
NJFj/tx+hbaAqoco8sFeTfgcuC8jtO0QcQ8rRXZF3S5MHaKWE11TUn/V6BGytauc
y6rR3r8YynbEFbREXZAuTO8EmrMFpyOStm3vYL3MYiLzvmGHscy6Q3fPHeIt3JpP
KgTG9926SAuetz3f52TOfoCne2dKMnSq+vjqfXNVUPY3QyOSgQX0d0zsdr7cJ21h
PrnFnx1/WTES+QQ5DPbn/vi0PV18pLQMAcq53aoAcF1uTCQvvZtkoX5KyEyLFhgq
z+B+cfWv5aN/p2m+6P2kT3sfA8/PcHhPsWlAXyjyC44/+gTppmeCboH2+JLQ4MzB
bZxQM9t8kJa5EmxHGlquxG4MT3EJ9Rrl0WZ9O2rgNs8Z8a89GO1+G21Dz4sHLbI+
OjcbW2hAzY99Wo3sCG/lWkw1DLr0uWiSHp6TiGls9FODt1GUlMFMN9d2zW9aICGJ
9nHddZ71zRQmDvA6MNcZfxTGIavp51matcbAf+2Q8Utbt9wGbIfRXN+2HpdK/rQ9
+4XGEcIfAqteT22tKCznFH4A0Odxmkc3Lu897Ho7g1roee1D+ycK4G5eZBt1aEwZ
NKQ5ld2aXLZq25inyG+ljez2oOYXYIQa8ajH7kUtxGxsZLGd61OUOyKe5O2rxvfw
3kIyyx96OquaFnCXfEEA0ObzLM3xf6HHrH3dYF4yJKjF7zlFh/YTrc0gZL229eLi
bhsTn6YH88GRz/gDNJxjrmqYg/7NWAuy+cJ9AZBCrDhzZCRP25MwOjys+W4gdkuR
N3E/FY9/nnvfgOWfX19s/6eaTjCc++rDeOkOU2SDnQ3cGe0P6/CJzq4lqxsa5X22
yJ5gco+C7ubKLxQ4mQPpuCo7A5p9Cyt6b0HrqpPMF1qUpNQ+vXQSWsZjzcOAhrol
LxvkEzxt2GrxWowuYjNMttUZA6TRo16PYnFiOHuS8V8cqGD1bITkiFDnka4FIvyC
JOW9CMipl5nJgts5h2ydC0lygl5M8kMI27+bPYZC5IX0f2I4Hd1LB83+IwimJxFo
53P9aAPtAoqM4Uxgzi4p6Tyf0VTXtgjfsnhiFbTeFth+NR7spPWBxAVJKVP+ZD2o
VCmMGkH8VYTRM4ySU000otpzvgyLy0Fi1++iS3Jg83G24xwUWYI9G4Bcmq74dX7I
2qRjdSTLiNGUwaGQrD4Vp2KiYO5B5K9W3vH8+Vr9rL5xZl21CSqG7/o3kXNEH+Ub
CWmJ+FIOpUzwenFYEs8eXkMelJ1VF5AQ2iDyFLGhUJv2+tDRjfxnRYfg1I2AajVy
uO/Wvrz7e9zU5HieTsgah9szUpcjhVS9SvXCg4Cjc1VBjo2lcxSRpv+6txQCMOqQ
+NI5vMBV3jBM034MyCcAlHZISX2/UdGNvNVSM2CN2G15OV+LGxCxClqOtHxO1+9F
a3/E3hSoJfzYDdo+Q1F1I1/AWFpNcjjpO3mFsZcDzEaqhIs/kVSaezjQ5T1bT8aI
UVlDENSV7GCpPksWL6fvlWg1psx6wrjbrIUBSHJF9f0F0ZtW2h54q9/V9LX4eO1f
WbQ62ZOAheQjAFrktmBGQaCu4X1yOH/74Sb6TyLMwWEE6bPAon1iTxj4IjuGlVT3
WabH1HZ5D+z843G9T7UGvxtYKvRJ6RDulvCGOHsquQGPo3JtXMk2ZPOva/40zqWR
w7KHfREaE4abF0ccSfUXh/C/gadbCz3oWPnDA+dP9dfxkWEUnbL7iNd4AFgiez71
93yWzVyUTJmmcRHqLkSTigC80uUwUm9N7lPgs2aPQuJcZ6T55XSJ8jRlP3wzGTwo
uPp9I2B9TUEuALnynpV5SqXQecZ6+pW5hXATLR0+NwckNVC6VPe1pS29D0pboo5z
m2T55XjarhTaKko0MbkSvOTD4+3w7S5bgSTPbHKHUm+CJPzcPZOWL7u8zO2fKWCg
jZxv5OfEKQrHEYgoQFpqI5Xcy+02tTxpIVz5vvMz2vtYxsnXqq5SGydvDDevEctn
8OiIHR8sDqbH6BTit/yiMCokrW8Vd1YYCWuTbYBJTQajb17suVkOvk9Bc7UGQBDN
sYTFtEvq5xMbz5TFBQFXD28S9SPUPXLBXPB9EGbihklOE4p6Llq+cNx2fYcHCWju
9d+3irNJhDLpya7nB85Lxgvb8p4v4e/hWZK7PGOHTf+XrEfZPgr2ZIaBFVAZe5FS
8WefcjkdloBrDLJ49WVeghZJ/DyI6TGd3qCdZdp/KdHLtCNbcnb7JHGciDMGph0e
RjfQBaJi301LnPuwaNFl/sWqQrH6fwfaoaOoNIXN7ffKiBMYFQ0qjd3f+m57CP1W
rKpS6UFtb4I3ExkxJ59Q8O4IcN9Kh5eTpZfGAUG+jOi0ANPXIj8PfZp9jUVC2grC
XCkG6zqgpzaFPkDK/7OZRstHO7zOrRaLt9Lp0PI1LOydwEzJSXeoTfmKLMQZ/VYd
bpHUsKxc2+rj/D/5ec1ejmdIzm5xuzjtPNJl8pHbUrtGNl76uNnE/ZXXq8vinwKn
zVmtzW965zrp5Ca/GotAflKJ8Z3rruv0qKfpUlsEPSuuIn8mdVRzIFe9BFYWNFJf
GBy2gJq1Tq32wCRQKZlsbCGeD31kElmrxf+yLj1b+Zs6RI4nPH3LTDSSGQK4akkG
ZunJXcSpOc19Xd6Dv9G0Y2JgAyJ8YpSttf1CnUGWrn2BP3U2s5uH0YIhAFLN5fJU
kpaNm8dVCvBQj5E1sYvBZXHA4G6Y4sRytoI47b5ObthwBIqWvdBClg/A/sXybV8g
Pda1YlFQSD0kiY7YUA7/H/TseWGkXX/ySNAhMX9dRiMxiYqxLbMJQgN3Mo8WrWYb
DwFFIkBpf0Zv8ldMujiZCiIiFCCAU6vHBPo7DkGCLK2HBTFWn2utZp+zsO2ZeyPN
2WdHUawGFQDVJQUCQf442AM9E4FAP5Sh/ToiCfZbk2/vNwXPb4vzCryWAO/aB9Il
ZhHSG+ondumwDuLL5iHDERbCvQb2X6GyxCL8TqfBWJK6vLTnZh749SRUR+D7iR4H
+cBs7GC7ioxxSkTUesGVelyDMoKE2MK27oM9M4VPRwPDiIiLuNpB+oEyYcB9S0ln
xo8+vthHa1DP5ePtI1bprvBuUrw9icVdeqs1rp0MBfEXDEmLHr6jNuo1aGGfJzLv
F61lK2JbByvhGo6YLhIUk7fqZIAHj9m+J9bGnKeilQy3dAHhKh3Qu057Ecw5DXtf
2/HRApYEBK6tv+0shOzJD1OFzekUBzPfcj0tOgJTAEGGe/PpD5d6jz9iZ6cAA1WB
Ve3ffS/nE/6TITgnwSAY/4WdGRGcdL0vUf1zpmss04bg2nza9PQiRkaWFI8qtwDs
Gbl5/uipZ9kg45ZLQJfrzP+0CSxWN82m9+SR1ytgAKSn2nQzF5B0SsEY7Q728kb+
WJUaPFeIsFu+gXGN4rbK6xKpuFqVLIiTKXBqmTHK9sbX7TltI9zxnBTXLW/jMOWf
EhsWA89jixgY4HwW9byIAlzDYeO+LUwrRTq8weYhOVczNJGwV5XKfstwJUw6w9Fk
fIuToQbc3zo1eKdMgZwSyYgiGD8DYr9mtQyTRVefKrR+49cKqCz4bnPFw5qIBu0B
i2MRo7LZpnkhGou9EOa3FoRlHF1PL9507ppVrJB0LkLwh8TsXpsnrg/0IPuNp3R6
BTicDhhpjvapaIXb9SS8H6ZLGhL33/JbS0yu81wJQxinJY2+ei9L3oH3gCNnyDxA
a7umxPYNwIOXn7ONkunpyv/+A99HztnligAizobTq7Klbi6mqpdr8O1MA/FZrfJd
l3sJemjhiGM34UorQ4NZ33Hv9kVP5ORw2itWKsNIsi0wFkKXti/caONsddVcy8pW
ytqs3UPM/yaI0g97dCCqRDAYW7aK493xkjHsLTVuaz1JeWqrgSbRGHds7LOHEEYa
bgR4/po235k+yOJUNvx5ImyZfvGr7HZ5B5bfZL3cva0BPYOB1bxTuJGI5p9M/T9C
cG/MuzFahUkCom5QVfA+RN2s2jzVZzS1lhKkO2HHkP6DkCDVJ9pKKN6qYEf80/Ce
Sk6j7WkHknj0n8GIVl11byIyvt9t57K11tw/QFfxW3cqyF/6LuV4sug9xzxf2sXV
5K0e0XNqFe6sLU28WyUC8rKo/ZdiEzM1qPV/LGOJ+tIOSQ3rvOW9ry1i/cqqY3eD
6DOnfLaouN4ZtZfmcMwQbH9/37lf84/NEMUe44HohgFwXn3xK3B9xLoiLJdiUV59
++OzgUNZgEu/bpJXEhOBf3cLHoaGuLkpiB/xbDih7ThPG/dYutJh3IfitghSZAzW
ewVknuWqvNU4o/m9XUVc0OcQJD44BqbMT3Ll0n5OpxnF789eoolX4M+nkegk0nDh
RwHi7zwEWdyISsoiRDi3soJfwjPKcbPKL3G63XDUwFBzW1a21oWxZcmPGHEz3ZAH
+6vK2vPzLUIUVfRdbPQeae4KnXcTIi61sX0W1wyDP0/mKjgBhNBv8uil6EqI+Wrn
vDwwbRLYVcriZRJT9o1vv1mAv577CG8XkFGs01LPYmCZAxlW0CqlmOcprd4Pf4c9
pnmze03Rx3hUpt9iSUjlsnOu4zw9UmaH7yQUOl/uBZWRNG5abpaX5PKS3m3EaKCW
wtnyQCkM6LwZDDbQ3bQfuxQSOPukKkDQrRSeRP0SIfeVErc0RJn2GeabS00HPJIe
OgDLi20Z0liRDQxTW+Mpty/I7XiV6fWTSxdltvf66e7z4PjrhXBeRerIhfiN7VmS
jUFEcUBT62kOjuclwLF1uIaG3gtSBiqzTcIpxn5P72wyaO2+yDSHdpHrfeda6WMh
yXs+r4Xd+ROAOsYraHA0hSWBAIuZw5aOh/WTpveJSLIphPVQJMw1ip7ao6ajIcNv
TmBNo/NrdfBrMMLwVYzluk64OxYBlVgEcgL1qTrMOj8DVdA4HkbJArPt3O6fURD5
k5J1InbgGzlk13/KcbqVqE8Q1ySNSAGm6oA3KLUDnAUNcYvxEA2TztgxgoOq/Fta
KXQys2QRtz3pCWcLoMRb6Xok7G2yVIAr0lJrVQEp/Qiu9OXRcn5JZNoTYNCwyvZH
uSrBwN7tivwgnwam0EPIKOFreFAnu9cP9HWxAQHHIV3hA9YrSKDjRDlTXvyhO8pR
RxIFLKPAM2+rRzIRDTrt4WUttCuSbPcvHyQXsXNF6k5cutdYKm9NFPfyt7JOOaxZ
ByPisWi3tTL7mVQGz7dp+x3wmbl37MGeTZnEU4RNAr5xgu2FD2BnLMj0ZlDjuEW4
BUE2gzdG6LGI78642JcqbF0UdSaAPhUM/kHWyxvlkum5cv4l7OnUcCU1LBu5IIa+
v2OWBjPMD8BWpvqHd86jrRjhxVVuDhvmPDSRlAAFj8RWKgOrJI37ReaXpzNnRMSA
YfHgVeqQXh1irvRmzcUCdXZSYTMlsq27ZFP8KqoH+rWqlWIUtt8r3NtMhvnfZu/L
oHOp8K72o13j6r+ohwPKDzdAYqbqKADaNkL1bJzUfToyY7X3kHoSJIs48HU0OY5I
40ltdwJcRyIjzzu+eIjuA+BNBIeq4jeJwYkOtEv75FBW5yhOvI4IXn0qJ4AX56Zr
j51Xqpcc3X4pIk64YL5S/keNKAdjSYjR/uB0X3kHtEiheSPMOPiizca9DWTs/+7H
LqwQkwzzr3Cr2citfwhBtZWlix0OJgXS0al+IhFaESWfUb/p2o6tvUE/HSD4qe6P
MVkdZ/q9M7cTrrVJF2lmbc7wltj3Atmj9GIYApbUMcYz2FJ7dCGWYpca7h8c7y66
OPUpvxc6XVdw/Vx71eGeM6Uh8zO0pztPZkzCmT/l6zIMPOEtWvG8EFEzTuq6NqFb
v+cPcl834d2jZKOqeOrv+d0rAI3N0DdRo0C3Myqqrr56LKAXpbq3L2Ffn6JCxbRY
39+5Sm/OPVb3ngdqFaRZhg+qUukk0NbmlYDKelIG+F1iTdvFE8JJVsmrD5YMQyyn
3CDFbAq8/gQNJWEITomkJXyDT6V4GkK2djxMPL1ZUSJPWJmDt/UUpVcjGmdPdS4g
KRNXpyePtH611AngFWOTeksjrKCABaw09XnQKPrvgqojQOvzn19+iAgts09sjEgT
jWw3Qea+tZbjsxeB1nXXNU4EiyuyjZQmH68k9Hzr5aSBf4RfA94ky8SJT2rQhBMq
3gbT1Wwpwy7I4FSs5gKlwZsk3GeMoBqNKKEVzOeWjyfyoJzo2qpin3zYhC2YzJ9A
+ohMUiAegb7ElnohbbITRtd1Uuk+FnG+6nuYMt2IePwbNn2X3n/EdkTPYhQ9XcWT
pR63hafODi2Jv/vtLUGpWLxTBjxQflTpylF5ot0Ecd5BG53vHuEW8TZnFdghSYne
V4PNAGgqybQMU/Nvy2zkASoGoRoO8jBLj49AU5DVBa/G0lGw/GDdr5i7ScXp7EoV
NBbnrvmK9fhlGvbYJ0Lx5QV6xh7TlbDF4C9pOLbQZz7H/7Ghmd4T2rD+e0iw+OVR
udXuIg7M+wI2RuoqUUkrxID7XMuwKnAw3KwdNQB7Dlyp/X7vnWoD4CJZFKSU8ZqG
e/u2k26UZC00uOE0+D2ahZafqJRLmptx83rN74KSuRFToMgWlIxxtGjgQrD9xRjO
ofqxT8hlDvMeQ0s26ZDEyj0rFQzsqfNT+/F1hTGtNsNTY4thynkTufjJLL6A+qm4
msegRNTaaOHS5J4gv63Ii4Z1igjzb67lVBHKWkBd53oUOQrKe6lMChxIKQ9loKXx
VARAOkHLfoWRqy8seU3TH6t4/dLnBJbOx+In6M0LA/3F7wylZGj5hBA37ZQIesKe
OuRrmYf+Tv+wnhmS565qARttCqTeA1qVK6vSOn9sodPiH9hFjNFP37L7mPz5hdDu
C/OPc9RWWZJDLwN/C3JewVrG4Ll7OS0i+t+3CB9yQUclJttbHguhbdPbDXnn2cjn
0Z+vG9frCQ4amg4XBxWp95gXMg69VGZ5bw/OzeBmJLS+Mxk/I3nlOVFLUgJCio0I
u0vnbGeTQFZY+cokIJ4e72boCWGALheqSD2OqQR1SgSNsPQFEzw5jfKKDKpAdeBh
lpnlE0Sgg6YU0QE5NEjDQ2gWOXU5M1J3Rz2LhR2Nfcy+OMpmWyPYdk0ndyfnbHUU
BwFTUGPh4QOEpqFJlRVihW4OxQDEuSPCtWB9EoTJJ26JZs4F0QE1N0jvbjIjz1w8
pRJ4jr6RxouRzkbN2g6J2fCzm57FR2FTyOjt+a1PMkAO4s9R/T5KnTP4Hfioazi1
d1XAcqYgwHoWTn4lQYU8r359hvt+8y231VZaV6G5RTsobEdsQeZ5z9y9qJ8uT/vH
JgjXsO/hvyrDK0CkJiEwk47mH94DBe4Hv4SaK+oCTQv9KaBa+0LsmTjctVANfu6Z
UkkzyyfeKge+eGkBiANSYieSyTOnPoUjjH19ZNVnrrzZBQT4KbESqnqGZPNFdYZx
KOj8IYTAaD7qDKsWLWjQ3RtaHa+2GObspL1R+FmwiYWznX6dNBAwy+6KgpF3gt/e
3ta4EnboeRFVEWSb38mhJ0CQsmaFF4aDAduTeGaftqMuqC/wICsUe/BrS7d1HSBA
36ws5JvRwIk3SvdKqIxgYm7Zr1sh7BrNMhaCdI8fKXcCNtAY0LtdtgTUEMz0C6qv
uD1Lv/Eth4Yx+ck3Uz3kRHkYFS0jX/IMwRVoydEICHlasolmD+4XNzHWRTXnPpyR
aj4x6cB5uP5XKUhpOUPf6Fy5HBZWgKZr5cnfr0O1yCHRXZRQjhYvh2ZSpcq3VzfB
fnxsDzDUrGQjrHZpZ+5/hlsK+LJqQED8i8vkJYYdUIvKFK+L5uHN4lQOwzvVto4i
4utyAtVu7qOrmyKulfm8Z91IOHSpx9tX8mK0uYN/a5l1Q7GtgbzsSiDUZPYqSqk+
8uCqDiZtJMJnvngaqM2CFen+XoAkJoGuG5bStQZ59NpWvawOCcCek/vt38dnFHza
lTZtPxU3aqj23YLtmLhtGdVT7Y/JsVvvjdHY5eeZ7ZCgOy83nzHZYYdHbDF2r3AY
9M8fjaHjEzx+IQboEomMSPJHv32cP7v/d4Jm+VbJJs8PKC9tP9W/QjEHICNBTxzZ
N2RjrPaj37XYosHWQCVUfXuloKIfIvoI6wurYPgbsqWq/3dAmYgw0y6d7Y/eLH4d
Tf2RdX2E1OwowWIXjT/uPxJi8IeTx9IYuTseAwCYWrvZlsfTFdFaXxtgfM+NPtmB
Qlb/SxKnHorYMIQxzI//r/RtdbXQCKmXRbSAtqXKMxEMiaTOTP7jZqNqlO4M0MHE
OuToIjYQbJQzJ4iqIUo+paXt8GNxPx2WLS89xirSVJ4rKkHWFDMF9bD7HvTJOoKN
hXQT0orFojYKPqrKoPysyWDYLRNVpK0euzQOwIGZUBOB4ta0K6or1DTtBOJ40PqM
CXnD6qcvuXwngfWXmkdRgu7LaLVqXtHMO7ihWcMRDc9m9JVc+Au/TrqBbEX4+Jsj
QO/pDvwXYNh5ARGP6shF4czMA5yuunXhypuSJzmVh0mqBivGIcj7fiA73B4Czl2p
gG/XbWwXi5H647uZAl53w2d/4SI2JZbi/aNhWRYNfpk2W+R70ZOV7pJt6oimQFrT
Q8Ru++jg1Hc/ikFvBjPuqVUvsVdBjXwJf6mmaqnRNJVmRJCOuOsG6UQ4IAqadv2z
cbBkHiVx+ChKq/2+P/YBcunuVixBKzXB+SWIv8s4t2voqkQGM1CkDeF/JjJfBvXF
FiQviXwEBGprm2P5k0l6wyQcCGKyYlP7VB1sQHbd7zpOIM/nqydLM1o8f0KmtiHo
jBSUs+HAsO5z+Iqz1z1lFIhH6lO0ynmloJTjW9dynoMBg2awO1L9VE0bjN6taTVQ
1xl12xKHFfULMnNx9HK0EY+rC9LEUkKXNcc62C6XoJCUFPtY7mOb0OAuKY0uIp8c
AM9dIdJOETNg8sIwW1ac+dGQzqeQNxNhUD2nXb2Ddz/Vj5RNEo0JrJnblRWDXI6w
q2LiEldLZ8eXV+NKC6LgdaNmoZiK9lRSgqSNXplzIDcf91S9+lB5qsOJ5M+IB26e
PomdanI4+NFHcvb7rJw2OdpBkmBIfi9e7z95oMefPLv8LVak/gMrR/fYT7RiHpzj
skyFAN1yNNccly/4xgSYkk10ptgK1Ljp3iyjYaW0oRQJyY/DQeOK48c/EdVogtyL
kWPjAJdoD5oR2Hrv9jR8V7hTXCdTNs2gywpv2v3IVjCWqAxZO2vVAMfhb8JE/S/U
UmjzssozJwM/Rl3XSCc4INnKBMXu9Ucdk97FPetNZ1wCox1zcI8pybbxwptS7LNX
P02n7kAYNmJH7r9v0un7cFzwdCDWCHGo+xwat7vwxV7jm7cD1M2mHNDiJPXDPLQS
i+7jblJc1sP/ijm/aiytQOA64aI5prtFINFzXMLFiWaBkPf/SmNThxgKp+O/rH1h
gMLO405sMs7/jlGob5y0zYPZsyiVv5H1k4d/z1fiZm/6jUl9Fq2VwLUTfRfZQXKx
UgA/Y+Ue9dQnOr/SBaXjZW+hZ8jm2X+tkZiHCOi2fJI2+0YyapIuC0/DtJ+0+vLX
xMiVrM/9WhZo3yoJMwguUUEiOM6M3oMSLXWPygSdePYWJNRXPkiZTy6D4I4vHON4
z1V4nrWO1doxaU8JhuezoJSAC26b3kg+dtPF0S3dn7Bs3QqZkdoK56lI6aSKPwtB
5wBlb2uDr1TWMjmcoRkxT/2UX33iEGicd839ZXTszKH8pNAXmTM6GpUKhQ+pDsrT
4Z1V9VzQ4sBRsuqyjCYmGQCeYQNGVH93B5ZrSp8G+THjUFpj0Zy8YbDlFJg8u+XD
69qFt4hmEmA2s/N5MWKZg1qlxDVQ2xHh6WN9aO/QdKFoOHZoyBLzpe99LeR11g4U
3SiBQmA2qYqpTJ+cooKLIXCE9jSA/c3n0hE9Qo24q117LzTrLfregCp+z/tLKoCC
aQlNoJvQR0TlwmvdsydCbiUhhKoQgtCbM6+1Zssq/MCt7QtgrzvwRTc+BnzbYCWn
yrhYFi/qAkHAhKPWdhm7BIVeJsD4lnJdDVABUVoAtemjkIunj4mwQxiS4meHAh2l
u4HorutT0vFlyiaF6KmrdUMqiGZ8Zfu7zF7BhpoGrP6IXKIpxyytSia7238QyGxO
d6UpaV1h9BUJdh3gTlVOUy9dq1rMgVeoEPssn4rgPdRh4LXGn03mA28uKQDLa08s
2OxATOtmdiDNEo3E9lorKFqWYSLt++NImXfbrvysW2Vq7xsKcAPJcL/+FwL46i+C
+2Er2RmWlge6s5YDFe4wjapDXASV8SoPHQ1wJJneUPL0j9j8+VU/VZ08L2VkSI0y
bgIVGQKlc3I2GcQWrkF1fd4d2OkWF+axhA7Egvbi+2qONYY93cPlTZp2JEc3Syd1
JjdXwGEZsnOxkdVcyH0geIytB/l0zndDHnAUKVu5HCUCVfkuYHHt9wUOs47jG+cP
/LqZFpec1xeSqauU1IW+RjVI6BP4GztBK3b2M+KSDV2fd+oJ7KqmstZlZdNExsoh
prlOhWMkSvoyMKcUz14zMh2v9Gj4T9HUXt2IRdqk733xqR7RTkenihSe3pL1dLQ7
iiT2MjW86YZRh01er+hiT4GvGf52mirhQmt790vsiHFqA6SgEo1Dq8ZYPTIT//SD
eQqiJAYwlK2bXagFpxfAQ10GnziuufmJu1ob5c98E2/Rq7SqT6f8Z+RLLzR+QD4K
3XKvyvU8xg/7JeVXD9qRbrIvFJVWuzMn54NySTi2HonS+bTfMl5jSTvmpiwCejqX
UukjPxpm76mgigVxOjjZqBt371eXSD33S+XodoMXq2E0245v8rWdyCpJWl43IfvS
74m8dsaqM1J/S0QTXjwVmaVuie7LrJbLNIKDDnxTUzrJnyXVRD1NwAA79cQzTFsT
dxQmnPVae6SvQ399SSqmWI7fEMVQ8fxrNCxvQGSFWaMZebKMQf64xrrkjDVBDJx3
FQVTTKKopuz74CycTcm6s11eqd7MUsjEQ6T+kuHcMdim4w444FTf+yJ1zrQgkZgx
gvfptKczWVDBPvg7Ta7dPP2yBhj+t1j4urPkoMr2g9E+du88KtzpCPNZ5fHRHhea
Ht3PxI/KCEl2BMsKTC2KA3bXPYHfmPUOS15T4zwn4n9DKgincPTnmyyfGPBPOgNE
aexsCUPohx+yC2rno7qR55IDjFbd/qRt+FTnZpH0qhUCaPvbl/IMadFH5g4Xz9lb
OQDCT02krOfh7d5nuASomPor6duJWL3D1o6M8UGAQAi39TCkvsq+cuhdkFxbo4t+
pmm7DlbD0bKRTlI+7CQSygzouKtqVkU63lup9GMsXV/a1N0n8/TOhilX63mlzzZJ
wIxfArE0BTaPMXKaR7aWOahXIjsvcaJhQeyRhSDYnZT+GbDGSUg46+ZaR3gAzkY0
4fYAus+MRgThrhRgOVSCUUDDfDMTdpvSoDpZ3DI3OG0Fs+OGreYaGz0HacjnCKHc
fyGVQcjGGL1bjoFo3lTrFL+QLoj0GgDQ3HK8YjUSOX3DTn44sZKYQOP9Eh49sabw
5T2uMP1gNgunsjD2+kZy7cRazPXZBoh/Pezd/f04ygcqnfpAKqewa97mC0zyDXbD
QB9+b/PYa6h1ERhXz3FmUAaWAOKaogPAQpLIHqE9QZ2TlXq/kEFC2P/tO3C0Uu61
WDuBDAGAYmRuNbJKZmevFTU1b5CwQc7ca2Y9azlJIhNT63SdQiYv/sVwCLfJ9qfP
edVUct+9eYV1Q6104epwSBtXrK3CpB6WfvNCvfYa8Dc+S5dKqlfTxoHQWrGiIphV
JEkITjmyGoBw7PQwx1iFvx+xbfsr3MuFY7ZrD2VxSD3Fr87OAD+UfTXZmC0p6i3i
h4jx3+QMcrLKKrXMyFCd2jHavFsefQaJ4Rdy3XnU09kvJFEowz8NTiH51atlg6wC
aa5plJYaM1qpS0pjZzUaC4qGBexdOAu9qSFK0CLE3SIwjhmg5vj/DB6rzHc7f0TQ
to4iCwf4O/VAVWhaeZEl6SrlU781tdAiTRiBv+Y6Xi8Aj9Zat5Uvr7lIwHfNJLZH
s4ECR1nxdIA3k0idroOaiY+ZroysbSoP57+FP2QTVDxG3z6K1JRG75G2nCICHz5L
EgpHsKeYCX3BJ+UEsHubgRlK2ma72YLwSd/FCkemQm+xv67151fmKrLTblguLfyo
iN4ecvsb8e2nW8hc2EE9wyCGsYxRsX58Kc9O/qEMFeqsNh/oe8H4z+wf3gdJCzDa
XuyaiE7HvzQn9YeLeH3q9NriC51eQZu9oYaGkqJMRkIKgIz6ukQnV/McHFDjBX+S
Y3Ol6EtwSx8OZt1BD3dyGzFntxslfZ/FFXc9oRR+jm7Cxxy7hTdenZpULW6WD2Gp
tGYp6T9Y7b1/9acca795ZrIQ6BTxuJYQpU03otMqqBOMo8Tuu0+HIhfi3pClIDX1
vt+p1Bv2ugiznzlM3TKtzfs8anLZCrW5AN5OIyuFtmC4XJfu6GNUfU70Rmok6tvV
FpM3Dcn3GPFwj8KnmeSF24DbetJIp3jsaUoIqPTsM9PfnX60JCAW19jV9uVvVoV0
Lr8fCky2T41dewPKZ4vtM7TRYZrTB09KotQ8KkiEFBn0PpWiBU1NbX7JRRBrnPyz
IAsHVCcOsIZO9EjSS33q8/cv/4D5dw/iZkVUJVsTrNagFgOpLhDapZhbQHBmgO49
P1iOyo+vyXbRmvqRS44cIAIat5dgwfmLiFWbzf8UKHcrc8+0KRtg+DSFW83iqQCf
dwbnqsPfqZ/4+vSU+Awqn6mVIBTH5JZWCic9Q4tTVBY1Ow8All4DxHVSk3cHqNLf
FcBs679sRVjWMECsjHpnj3D5PsXkBxsq5sbHDpAcGOfTCDSSbma0e3ui7R0FMHV8
8q4AVTFthJv6G7h8CrD2u7f6jhPf3eH43BpWYcvWx7AqVenzy5iJ3voxM4OjNezX
xrzSagcCIkmblAPxKQc+HYZS5QGujh4zgQ6CeuuH1Fq0O2gTX/pWRwVJIL90lXoN
Mi3d7ONhHFPs1/yspZptOnbwmKJKficUpx7qCSPxJKCsa11+vjWHTlrVmqjPBIHG
OfOK1ac/GLW3HD6dGZCII2t4cjKqMSGx0crB16VsgmhRj/lZ63L4jVNGDi7S33XR
t6IlWPCjKvS9Z3L2XHJEvgxaEhb5gxprNSU68Tb6oSoZlAP3i8r743NBvvugncGU
A3zHzQCzyI4pZzND96ZCl3Jy42uBqmcrqB/H2TPd+K9g0okr6yJ7Nmrv0hxYn4eh
0iF7WXRPx6p8214lAptG+zEXku9Pa4bwnPgCyzDbE0Jbrt8q8Y9TDMgZd9lMuYMN
km4xS4/to2JCp4F5meC+Y2pCw16G3+Wv6kPASeAz7VXtiYaWQyBwRT6bvlwvzWMo
rfWofd5oZvGfV3PeqO3ud4GocUFr3fuZiFxjt0/qgsci1hId4MR68WyFTvsWufFv
z67ktOXuSu/4wxiSxUPNXba0u9nC0w3NHxgIJH/NxSEjbX0SIYfwahntNaBjyozM
fCX1cJ2hbQ3BYrKLk/kbN+PNBJYcT3VA6jA/2b2wZgopmmkEqY4PyTfLpomW7WQH
xsYGbEPE2h/kz0CxRh00taKYPGnLoz918DP/z50jVc/rt6Ssg2Oqhko+p9QEbQWt
gBqFOIYM2AF41ltJkT0zqbU8N2RAs7Je/HBlCqlfB3a7vhmqq0ir9rnc8DtxW4Iy
bW2/SNYYuonm+f3ESihBr2QxoIbFWtEyvBXFH59vwgPzn5HvdrCooIpyEPhqvNQP
PhwPdlA8zF/ewRquZK74RdIy3V1PNrx+uDe59n75uDFlu5KgJV/RQviKAejcy/mR
QzH3xs/fSF0oulX5p8VflpR5wQdk7pE2LtCRI2W/8IwpuwxL5AMwAelLHPYi5Miw
r59i2nujC/tVEdfjAngd9o3wWJ/TDyWdEDmypCyvW4N0J7xQw9bBXieA7sBlcIxu
XD+EJ6t3r+U9z9roPEiousukImkSg1BSnb8faiB2+8lr03GeAxct0YqaS8/+K9+9
R75KKKUhIFirkEreXiYP48zRcfO8/WkR6eU/06a2OkQYjhJIfXtAflKChkfA9e1O
xxFylibAFmGTr2sIfxgJhGRGsxm5jYEbvIuJpqv9jH3B3/XXhwymObRb98NzBBNg
3JDDeuGW3Pq5oeg13ls2auRV5c/WobGrJylNAnscgbvnB5PRwx7/aASYJHYSsdE/
qoAPtlsvhuU9ky7niK+FdzVwLVBeCxvB2kg7ibKwpTvEoBz/EugzVFFUv0wkyEab
El8VKBUlMe3do2V6NaubY9gswgJPBe6iX/cNGEOpuOwtI4C36Vxrw80da2oe1/yI
3589PloOcZjwLGbZ321dnWP5u0JeVkY+98d8mN5U5TfVANq73uttMDfb7Qpwaaju
8mri5kuDbvrKYNP3uolnDrRGdVWu5APNE78KOars/LyOEgU5MN4FhojgFWJ/FrNH
ohGnA1gEicR8eOUY7ndaPkLBAkz9ODOP/OzrnNEd2wx3ylQU2OgDK49yIwZOcZ/c
18Gk9h4Sgk44NGHwdpxjGXZIFPicWDiwbYB+XbQithiFywetKNcmDdQ08orSBYcz
yYhSst+h3BLpaMfI8YljMairxPkfYYXrZSdoqZ+C5X7AtrmuT7mBW/e62CsCd/Xq
Y3KMPKvaTE0Gg0bMbSItxYk4xt8atLc7YxBwurka8aO8RNKSU490c42k3GThAfDB
sRZav5FzOfwGFxPS/HjAuPD5l6MBP7QGt9GHLsFEcPf946YZp2TYycu9lo+q3zQJ
D3/xv1chScUpAyVNzIuf/NK5h6Th3OTLYpJ53MQuR243mIySZSZnXB6myjeqgvkJ
yUZ1wxb/L8Wzca2JDF9s4+Lf403tnRVCJ6Qvb5M4nOf5/dXGNzOdq/F9csTb2MmC
GIhqNHgOKUood84xgq5WDH2+/dD9kCbK5o9izQkQDFFKdWPHS8FasBA4ekPBoNjp
U+PeF+XK6wYZoHPqS46V24oqapjATvHIaSOAgRvCBa/M+c2bVrGkqDcvwItsM2km
/L3A5yTsTIqkHLpXDb1jmE6wKAoU09NPoUOBaAUoVHNvqLC4MIX1PbHbhyElJbhi
aAJfMHMS79L3vEqzoYB6nFQpvL/fG1Gr3UPJiO4A25UPgbZsL3STGyBGi24SrQIQ
JarByLoxnOU08lSq2i60lVRhzlV0VuAiU9JG75tWY2gNJ/hrFa45dquKSYD3VlQU
OZuEGVIPzLW0gxpIf8w5tL3g2Ow26aMuycGuEl8+gL2kSYH/IFx7rdqfuTVcIyyp
jA2BhmR7HvsbyFRW7bb2yPV6OxdukNVOxo7SOV1usaSQxQ8dmgmkpkC+0einmytd
ct/49Iib99PQMw0BEm/oYWscAC7OtkR9Bj5N0o+xeYKNRvaQ1NvGu4lL0wMMlegW
mOPYci/lH73FLVpe3notcJfJL0uKpIzgFuXVCmyMNtIMgFzUhPw5L0pUPcojaWl0
WzGUcq9500EtTWM0pWRdbgiyT1mEGIJg/alxFIXQL6stIpRlV5V3BQTAgeiO9E6q
IsFS5jCxqs4QTrXq1N0Go6hS/p0Y9xIUGDwylsMrXqQ05Yx1a5yPGxxIloNMDg18
VL2o7mRsDsSo0bCt+RZdd8oU9sCLhIA6aQS4gsHk8IVjS2N+NjlGdTvoTa9LuWKd
iW5gh1PTT7vPdkyuW6goCl2VbBpbc1KOSteXTKPgTQnFS724RCPnDrhXwHNUKgCr
Ndm8mlGjtVk+RsryCfJMSpv4jhGRhXH9/2w9OfVe2VT0Unxgf6wwgmTtUFiPJY1Y
F4APtqwKJFwUtbYyNDLxKlxy1Tow5rWXzR2gcm/KL4p5itgvZJtibIJGk9WntcXP
11LBseI0F71+5nFtG49c5bjnRZL7vP6XhweWSWwFZveECPMB6gnvA579io/k1joG
3vHjoO652PhKRl/XIaMJYdiiN7mO9280SFXpgnDy5+NAo7N2vDAutIz1+dE9mTxb
uLuEsw+yphSnQLS4HfWoUU7hN3UrOaxqwKZe41iSbp5MBzKzIebrCmeldsm7b4Q2
93V/EGMfpv6zRx0bxsZw8/jDKUT2g2VjSgq+uepQ5E5PCdpBbbGlo2mgN0hTzfJ8
jDI9xoCbk9uawdKlGy1Fj9YbvhcmtGUZ+wSAGF1KHK22osnAUXRnKR4XawHQRN9H
KepXq9eCTIY9ANzPBRbJHfWK82NqGV5m57sCQHPGv36YYra6gWpGwJcc2aiJhe9h
8CsBvoIsl8QkcoUgyJLjT6AudK/0cZFVs6TpxUKSjbftpIGg5MrxpAeWej82MFa1
tNCsT42vDzIvte14iEJ5Bl9gUdZaB8kOf4PJFroIlS9FW6s9Nuqm6qg8fPKOa2J9
T0kCKVbGvgoKg8r6Qa2ZN75wAOtpSinzVjPSc0RMzeQLA/2aUwpr3HKDZDEpww54
kbZdaM4NOzNpw+EniM2qDFtEcAiNN9e/WNjar6HbD4juqEuwbtGLOXXpdm1Uf1SQ
62SYkEtkz6GqgS5qYLqwBjonSixugTQPQLUz+sPSr3QRwu9iAJf40iwhFdpb/x6e
YxNGPZx1ywn70ngnhBHPmrqQN+DPb+pR/MPNz1dfFtVFqwilD7j4pm/kroczZ4At
qPD+/4sUtWOjDxekKr7hlhGioeSCCrtmGaXU16GsM0HcEZJ1LMueD1UqNprjQ5zi
83IaVNgldjL/1Z9q7xnzKmWDXM53f2fhcpJ/EJdOICwbrMJDUCj84Sad8sVNlPkM
e/PhZMyPwYma5JnI2wS7aLzJuDBvEFtz1SaRP8neCp+VLivzPKpircAqEjgT6PpZ
pzetiQVj6wgH33oVeDc8zZW5FuWiJb6MkNzeb+x7WUJaZxFFy9PQ5685YGt/LKtb
L6qDOwc0hza1FoFAhABhvJqnnEkg6v5CWoLQ2BEE+S9tBih9v72o0wIS8ay6tOl4
c9rEZ8o4uEArvW0S9+aFBPTCAV1Y7zAGZVaOXoCzrcZPM89hcK6dDEzm1FOCy40l
KZP0pt4UyHjSUAAiRAXjJJQiQS7W1yCcPlB0CRpIMZ0JFvY5/hD9XlvXn0Cf8nkC
6dMWk9Zt3XRDNlEbr5OKWSV8IxlU9FRlhaQCXkTvrq8NWuwxG4SiRXqE94Pe/GEN
ckg6aytKVFRiMiNLmfo3CjHaGpqRxUm7yPzirBU4XLp3WODZVm7/JX4hTNgcqFEQ
atEzwnW1oMx9B2S+3i/+l+aFaWREtjctXOZPEf8hWRJ2TvxYTJaROq9hrfILKk/A
NLjbQyXwcMMSeIsYFVsxNfHJMXqzOeplrf/yQDQHMNBkOlxVr4k+VGYaKWMviJi6
udlMynTqSV4vk/8CiphoeCbexJHpNUaoU/0pxk8+O7S878tSSOr2/WI5ly5nDtYd
oBnhC8x78vgzhJZzreRjAYt6HQNpMipzjmfKXf8vjuUhq77froWMS5AW4S0vvgSq
nSoqXwfJ++Qihs886rM/MT00ENH6mGcsaILFFCkMun/vhJZ0JyTzdxpcncG7smBV
fbNIcLPAsfZ3r1x5lPVaHDIKh/nemjejfu/QSgEocQD9y0qdZdqYSAFYBriQSowG
B9Z4krhSDvwRqem7WalCi3+B1ccP8UCshg2VCUy2m8WkOyjrn0R7OQP42FpGhM+g
DDG3j47J4g7IEaqdPZaRXWN87ZGGaCc2i9BEGypcNf44SpMGW++U/m5l+Zdt7TYg
sGaIIslV7wnWs4D6j77qzj+BuPzhr5nrUlMdI3hkqVLf0DSTjGKWiVdwaCqrtoYq
mlJeVStFRk8kTqs8sh2g5gSud7WCazhfaVVJLdmzZ+zHxX0yxDTuo06jCFgRTIDk
hgEuw6sXBzVfnBkPd+lZdaOkuEiNMihMKYjvNX4Zg5t7/gxTrzBnLPvivdTZ9fHg
8AeFSz5KyqVT69NTUmnnMuUluZTRNT8DyR+FvZoYbve4Iv+RfpWhUNK0TVQsuN9o
0DoaUXVagaqztXCu21SY5eZnSXIBV/bhGICxzvsquV7XBHqoafok2DgDFbObGIs2
tDYUcLkBFpov+1YDJ8xu6fFbGrinbf/wNpJnLEJSNisycDJzEiREyDChG6uCnJPE
usbls7LcON1AdSfMyj4wN9nJxtfKTmcFMaw3ObVzXETcYp4bSiCPXRhu+kdhC2NU
F84afDq3QHztUedzmOPMhuQnd0scRPj5V9ud6VZO08bPoKqca03cmmOmt8FMG1UM
alpHwJIXtZmGOzgXSDBux2hwfOo2dyRnhe2G5YOB4stNq9GNtEoyKUdnPyKbHklg
hNVP1JsT9X+qJ9T6I5OIeUdcdd+rmJKHAUTXuIqkNLniRs2l94jYOEnzem/v7cMm
tiJBgmB9XWlbYcspu9HvQfViK/ecY1EOIdkBK3tGsvKmby0+C5wnJtajnNgfeZW2
OkY6kncBEjUlEXKS/GV+LG6g8h53BFDH1BYAvJE13EnvBPK5SFSW6C3W41yroTwv
bkwpr52P43OBpR1vUeXmwPioju/27qMXKM2Ovl/KcjO3odNS33zssERvkC6w7c0z
IgQfHyc3NfgCDcf1vSeDBlY5W80Tpr+ZZ1SC3dRLcmfoeUJ6oxnaSycGS2gaOGJG
iCDIe4hkMM/xCVbX6+nZoeEVdzHrfplJaHyynI5rMkZu/Dz8+maLY6SYORauIrBa
KRTTHNGRWCiGOmnJtBFnQhRcICOK+NLCPo1+ujhqXK4QKPhHkmgvXGCld5eWmhef
ebX7c5BjQf6Z5o+LxRz1poSV9kBftH1fCpb8QTKXR1zeTAA9V4Cr47v3Zg9pqTx8
qZFBKcbHJs1hLT+lxK9jFLAPsni4ZVoOV6jRtUcLmGOZQckWfaasLS3u3pNicx3Z
G2GxU2o+6BiX4qeBifwXfzF25H/eXldb/gY2F2ebnfBYu8aYKkNhLSdSXi4jLdpf
+osXZv7gCLkmWrmfu6bs1BwihfSUMf8YiQkYwerPwRwKcWeBtXgnZSc6otc7laqD
6riDc8jRXVPRrfZaSWjDwa3U5I1WL00KlA0E/8OaJMzISIxrxbLc0tqni0yh/IU+
kswUPMCiMCdtOzhyeZrWKW6WxJ/kdr0oBtN8CkH5QbIFa2hz6wsGzmoo5XJCwdtE
NcvbRtAY18sylIXW10nCdew1DPAExhHUTNIkSGmcokUUw4vtnOdfT7rRFmeqyu+h
bZw9hkT8bGRB0yDdGv47s75ahSK+NvWxpE21ZCfN+Ge4bFtsNtgTm/ZL9KLoh/R/
DQxtsElKqAY+B+c0yX4EwfwFtf9JtYngGRqwj3WfU5cRFTp6iZyPPSLRWMamAizU
4nhhfJ7EFAuuDIIeEl1Z858BCnjapVoCfkqn9qyg5mfnJQ0Y/LzJ/WCI+ovRLLtI
Z4meDlqny7Gwc05KFOuCNCT6in2wRM5b+gB4OUcIbmJoTpiAk5ssRmNvTJG5D6Bf
VCNcBQ09Bx57B7qQU2KgW4FV8Ja0SBcAkqpxuO/AUmQMEKzMSSkm+BM51ABSP7LV
eaSjE2UDxP6aK67TWfCXvM2k8JErrJ+zPdzF5XqlR0zv0nFyFJjgm/npI2f++XZH
jjEabZbcVjR002l0z1g5GjkPC0uxjteOI7vLhVN1JizFj6fdrv02NoJZZf6Oi3sC
oi5k/tCmxROUHyvf9FWo3HJOBe4JHvX8DFqGvbzfpfqRpW/s0looo0kFTi2+ubLZ
sJW0FFKtxWXOtLnDxFx9EYLQbnheRMHPq2O/Hw5PvHWWyiPh7m8hbe8FDg9HEOKg
LEikBlA+opxVVZZdKj45KtFBa4YbBV90mueqSnRw3XgiBg8oW8hDpF+USOHJXUHQ
oh2xWdRqcDEMMy6+XKa4UZqFI+qiV+rCM63FAiedpg8rbErbAUnjjvLGzDfBdIPF
xtBtwMOKm4NCFxzXP5wSNd6feSfOVCC3Uu6wye6/bXSX/Zh8Bbi953zHzs2quDuT
dSilfk3c5b01VX3rxZcUNQquitCOsSycIDIXl0BR5UPRYPyt7Fav8X21ib8C2SNn
QGlu4uAdeIw6bfJZb1sRSqb182DFPH0YLFErT4NfBHjo3wGTUlsoXLF6xnMkR+/i
aGm1HxLP8de5WB7UpSpuVsE0p50qwM0PP06Nyby0nIy/hTt8hcGkCVtaL5X3ZN/Q
ob2oC/F1onIKhpcqf0NFlVfiYjStI+qw1vqLK1kwYLbkG+L9yTxMnfbU3M61TlS3
XfHVu5pdIAGMhZo/mrMlxsrLFrE+JQahtIc7/6o+lCngCkECUFpK7hUqr0sWbG5w
J202Utr4wIiCJRhBqZ7s451wFPKrM3z6AIsdCSPp0lXrm3Z1ejhc+4OXE7KrL9S2
e6mvQ2njZ4ZevlSbjuwuLei3IYwoT4v2kdPB82WlOjYYipzjRiF3qT4FeTMmj6uQ
X3TZ/mTgmIl20hL7DzQZGJri6RIYNuRNq+TjUtaK+BDYb4Gr8+kbzqF1kslMbViU
D21XQ10CRFFINhcxinjpgHdYhhtZaPavBz7UQIQzMz5cayAcmzOquOYJf+CvepNU
uU0mvXOeHeyzrdBKXhYB/uE1ukDMzjENIs3Hk3X18I358JcV4WAn9x2rdPEmK51Q
hP6Pny/9YqAu4HYzozz1Bcz0XxkkaWz0UFKxusNWL/SdG5wHdoa9MGK8fLS2ynCN
Z5Xv4AhLogSXVvcRYDwJz6/cDApviXGybC11I3OVzDCZIh8MzAQh9TSWyCiMHC+d
lRblvpt1adYjq39frXTPjfEHmM2sB7zuDbQhq1DSBmwg4n0EiwrVKMkfOhR3i5XU
Dzdd+buvXzcJFQt88VNZUfpogd6LMSJxbHBsO7wkRIEebPtpy3SkV/GRScwjhzqb
63dUU3tdtb4QrdOnvQEmXZgpil8Yl4LuXbn3HyLrDkVZDNIbc/g+BWVCcdJYnbLj
RObJg1Gf/H6Xs/F2CdMVSfwIR4PQYi8wINbPcpDaiqI4bmpPktbXhV2gM6LsTnxN
1+2vb0Gq5UDmlHUSVcTMf5heYzsypydrLIDnN5CqKd/+t3pu0KZc81nIiMsu3d3z
f7cM1Rriv0JJgU3ANyOLcYsbAWm8wx7fMAuo/78uVzRfkVC6b7D8HW2tA1qs2gGn
0OESwrd4TCHsbdt3AB0H9usWZWm7/G+NLU8Ge6FBVoWouMS4AnjHAnms/wxWGv4a
2XS289ISR2iHlvVD92qDJQVDexnwy/LXroHhTKbwfCzx5G2xdBYXc6y0W8DEiXVd
JBi0ukUCYMYNA5LK/cjtOqefJgHFpGpYrNDuUQH1w3+O+zfhHT6tPdkVHy5Q7tlg
0DtrS4rZXsSgEVZdC90Bzil9HYyjT/VfL5D7LwlvWKSi7oKqkIhG8MrF0iMoEdGY
aS+MTSB0toETx21EkuD+ngSZZf6RiqXSJLzksKUFdtDfcrgKTWij/apJEjUOFgFc
v0LjYhFy3o82Z3AZ8pvcc2Z4ZlE325Zt4Igol4dqKIgfMzpZtS51hikFzR0WPNcZ
xi0HtRdGAefLoPJJ2h6OJPLctOTKIGl2WT8J2uBqM7eLRVSOAIrrsc6KDM32ZS0D
w62kGH7sn9K1/BQ+R0EZhWnrRzh9JSVj4S6hnl3hXfPcEmLGEPdWbmc96L6y9xkU
/zp4QpGrtk6rzTBjW+Dedqk3ETdnQ9Vsub3tm4W3CIYmcu8wfApI/ED58amnkjCO
2E9Ihwl1YfzFY8ynt85J01QumzB5Bm/S72Y7fFfWThqsgwU/XT++Sn9eg8Y/58Ys
9Jlqq/pMLpHzYwI1rX9HOhgIeOxO8sj+5Bfyp+3g2u89EWyCL2l3ZT0NNjSLlQMj
sUQeCLsjkGyzup25HUsV2P/Zs09My1MFW6mDeqYei2zOZbQIXqQlBxX1b6SSwfXs
MIDVg/J/dqpK9SZSXcJh+fiP1FiG5vH0h+O/a/KBY0FSUQ2H5CUtN/wnYrD9uF3z
93eJPyQ2Yt3cGqnzFKXuJmVFWVHyiUmerAAnAEQ0/Mec8QDrNCCUdye2P2HS0TwG
r3gPGseDi7j8r71evxHKczHvLTfzAAnKA65L/U0uEooA80YEEpYf/XWNllXXd9pS
OS7neSDkuDcMHybltJH3llFuu5VJBWQ3vBYAmLH7AYo8zkCZxdT1j5b1nZDMInfE
QwX6jsyB+Cxhzhvm1g62VvuQC3U+fZvzkNubEWiu7rtk6E4DvirUORURKZgkppa+
kClH0JieN/wWbpDtbkVkApnAKNjP95Y/4BB4MGp7ssUCO2o2g56umo0xXmF+rCRI
Bei8wbt+InahcJtcRFpdS4FKmxv6fonUvyibiYyqKREzRxLF/DmW+YsM5mI76Q7L
7DK0pNEbKxwK4jv4/eUsWl4Gbt5g00IAWqVK7sCBq2WumZJ6+3ZRxRzkwJV2aYLG
1H0aPMI+oK43DmJRS04ZHyyVjqTPDxKaHBwVEP4HRhr7LpoykWe5Woy8O5Jz5d0U
GVHafqbzAo4CAkYSwuAjdUVF+6c+WTnQiXAus3cRt4eq0X0g9//M7kTJmbWz1Z2m
o4uR+A7sKmGiXMi7pOYH1+c8Ru58P66PFQHFIzK/rf+C9XpU9t8pgZgefHWvtmW4
SIN7XryFFPl6CKrIHnCUT3kttB0xM5sHbscXpgZ78UIhIhWw0y4/Hfgln3srGqn/
kwXCE91bt+H7CjF5KoQBpFhyEReMkV0qcM86CiRQEt0D5BrTDHpQt0DfcFy8AGXe
rtriDgHqdUHFWFlMzUT6FLGO8HT7p66WMyiRBMpXMyrohDvWBk41cGBguH57Ts7s
HRkzje3THDDQpZLio7ZVxTkMjOpjdimKVoBmaXZWjJD5SImwPxY0VxtYhpMKYVZY
8zYjdzGivMo483mFVxobd9yO7lglhZeRCxAtBZmJo6mVmYOSz2znynyzT42HyRdj
1OEwPgCSsYe1A0Pb+4kjr1k6gbfC7cipgVh7IUpKqAF101lhOzA5Sl1Cim/3XJI1
37Plv7wAyAX7uV8He3Pl8M25E5QsouPEKJQVT3dtviMxF2GYlbDsrNnjDxqPuJaF
p8qO+0XNbzhR/D3OMVcFcnQsI4CcI7AKrzmGqEM6NqhoWJYgwatuL+XkER66GgAO
iQmRfJyLtbBWIH7JmC/FeSEGh4W9hPKYNl2oIKnxZJFrGcxSowXCxEKmZUyc06uj
MMdLdKPeTBLniKdaVZQXtaAEbLisB02yLMsXP8QtL44zapcL65Hl9Lyca6f0TmTn
iDwwd5hYyNV/yngqi2fRo0LRfYj4o7KDmyYrC2kt70MStzGo/59Lpqs+5LRixL5X
v41gzsf5iWZtj+AnnqeybIHjNzDB9Gbnim0bYFOeKJ7Z/1Ag1u2NaY/dVftvqxD6
ObvwO89IyjFxJ1V/Idqsf6EcFAjPrvR83EoX9SiGOpAh2OUqYNuIuNKS1FxCCclv
M0gs0RKK6jtqVd4hUg9xcmlPofQgnc2N6SbXTdm4ETVfgVDVJiQfw4ylHI5hSgL/
U0n9kjrzM1sXFlgWXyI9kcUGcUz4sGhTcUrcWI2y3KoXM3BHpT5fqj7+J1m83uMv
uxhX8Wq1Ck2uGEX5rTrQ5TepMtCytPDGf2WzZynhIGqyHVykv8oePy8PMlXtt8Nf
xea3xJOpgUELOhupAdfcrlAtuPLFRrGgS7oW38apmG8Y6qyyyFsOOgw7ZiIOQ2R6
YuWayKT44mbc11zSkKLQi1DVU+3Xg93sgZGkhTqoWWrFmJyryblBfHB6BGkZzvZW
2GuVFA+LfYxUzmxLKB4u9j1qvDC6CGBYwG0jjmlyU6dsO9SgaEzKTrxXCXsATxak
L+Ujxd5ss4GRd0HlEuMxSVgTv3+pUZq1Yqhq0wybJl8twnaH0Sm4juyMa6MEn3AO
9VcB2SEkyRNWSE61egqeqrVKtVIDFsWU9FEPY6BpeYYrjuYR9B5Vkl1KzX+CZkx6
Xk/RaXQ9z47IdzsAFIeAs3BVIwamZbp/FobLYurXIZ9h2gjS6Z7f47DuyySTxGH8
PdaPxYJtl9yG5ilpPHy+TjCXL5L/4kC9rP9AD+7ff0iqp6iusfPmmDa7rRNTQREB
fQSwLi91GjhAO8oWNXeKbu033gKFMJl87h/44eiUFHzcHlXQSTDe58NPgMrFsYKM
IHtW0F/uakNZEpXmHMWTTrxJKPigl0YlUBp2tCe9nMKscgbzueVbb4bvWhtf8sH6
KEpH5VFm21/BcpCxU0XtzAPWzePVnt0biUsLGfxT2U/nIkh3SZ8sgXieSkIR1xBu
tmSGx2XaF4e0IihDUlYD7tG+JAfngKo2VkSKRfnn6fwpY2gu72NslWn0b28uaiwR
+kherU2DToxB+HHUA7AFXe4GiSbIMMNvjC7nHPySzwzh2FfLFEabn/UM95joF3fR
rAo6vFjj7nkTzS1zCgGURoyiJcvZW9ZwLaONwi+0Gj6TxWNbWSC+ZIQ4G6pYyyXg
0n79pjz3b96V47aU4mvMwf2G9AAln64KGu3/VjA65f/RD3iyj2MmaKwuEsDu627X
mMOG/pgnPw9lHNds0owYG1fv7cLCcqAaVDNGZrKbIdHBZQJIf6Q/QM7ckdj1cGNz
IPdtfiN3vLjTHKOExbT8YghoLynXKeliv3WKi26053NcuMOQbZvrx4aAJvG7xXh3
Qp2tx29mNCYueDn79xP2EQJK1r4RV4tSwkcO8lUA015AnkMcYiaG/+aWN2+JOJul
BpJdRWaiFpC/Qd6hnnC8bYQnewvSCF65E0XiW1b6JGzIKVoTTOeGEtwA3em2K4Dm
pepH+bTkfs21xhMoQ4kB8QBDfTuqRJsBbdRRNd8rct3Jfru2EuzEbuSUzCkx69IF
74ScFt8QzMMqqLkIhRqEfW5lGTSEoxExy8WBZEz6DlTZmotE7f6ATJnxMyUTYgH6
tKOF29BQHSOsue1iTM/h5kuHksKkHzVv+VtDDwHq+aeLLdXDqaeQU0oZrjtpmy6V
y7QX53KhIHvZWSd/R7eo3e1hVIDZ1jFVs5IfdFXV40DowngQ4e4zg31o3swjkHyf
BbWUROlFlUsOs9DdmC9o/2L9c6cb9rSpQgLeUgzz2iw6/jyqXC3QtfNer+H2Ms0X
uchyFqM/w1ZhYYtxXjIeYYMGLmHivXDL5g70PHUNiuc++U1W8ghW/5P/H23KOYoK
aXvgk+l0zTVnBtkyOQTjdj1WfFDMeLTtOM9Vrby/TEGBSyZPirrdHeFizvNMz1Wu
6revpbS66e5qZFKKO48/RoqC8BPiuscdwqTSj58Cei2XhiXPkoYlUhoLL6OA448F
BoIPjcsKpXldBDcRcx1Sb4PPnrEI7pDHIAHDJjx45V4gAdpMH5fqQgRJHLFrDo3W
oMEGTB7m5WEa6/yvcfoBeAe89QMTFNOqS/2/yBRnIBuGpsds50O2I+iuh6NQnsnX
yVqfRkG/qM9c0RcbN2lrKnjmNSDvhfmC2jmhsfAxLckJKx1bBUTm6dKMNdkbP27W
09ilNUlJAVb6DnGTO2Q1z5ZxcPpA7uw/vrNyDuxIv53oquXEdNGjCL9sSyfyunam
7+EHk6Z8yHw1NmF4FyqR03FiI3u9+RNtY0wpGoRGkfeUNkO21P6NU9CZFLrCGT6V
HYxzcQpwlGz+CQOZ1M5wotwvwMmEb9yZf1JtGAaLZgKRrzanPeRuSbFxioofsV8Q
csO7aGrpMy2XI09I66gV9MatzhnZ81Rc79zpLJJyh6/lBGQmufDs+M5Cbv+i/Oj5
cdviz7O7do/M9j+GHQOohsvtWiOxzLSzRGISVNPIW9yX5AMEsnXlIfhXI15JuWkI
cVpweWUSRCc8AdAKQiXZBhthwZH0vyTSFyj4BZ1+prZB1Pw3Wjuq+WdbqA/9YazU
BxKw9khcDepk43CH86utfoKWh/GHvxe+2AsmfqUZawPDeSF95RPjqfa14+LoPDAF
8DzexVqgvBfNGgn0K2FExLWKrK1OmfWORyVQMSPzLQPuO9+9ZHV3PZX7xuAdR4CO
3p6JVWlyqm+4/2ra8IXq4quxf1ssAkKFNa28MeZQzyGBFRr34STJkODP4SGL30RZ
060nksWn9k1c6d6p5ZikSfT+rHeSEPjvo+iRUTOHITdGtNLRcZsAbkv2u1zpt46Y
7JaGfy4ouO2myKuo7bXjX0XMKdNJsmsfRy5YlNztH6Ph+HexO4oBmTTFqeaVRWdp
jflZLbav+TNn/ikeBnve2sEtWVppIHZKS9tGMpaWGfrn/kRRpkTGh2pUbaYIAKvE
dpqhjE7mIAlPTUu7opojUYgu6VIexEFkJMtH37Xv1BVK3ruLwiBgca0syibF1x9h
d07NMWNElY9N4JlvzDj1rrte0p0Gqw012vonYtRlJgHcUMYNi14Lu/vCtUwauKLm
jBazcX51ZNwBhUXhFIUCSQDIJCZcP1hFvhALHpxYhBofjfPh4GvsrHfTBQOv0veZ
Y4w1PUDVeovOUNJcGjT45kfIO9ojeK4ROSkI7ckqeO0in/NYLzgjJKAd/N3BelmF
nzpwJjJsuT5YYlec3bFPMu1/QaEhiz5OCb+lkcqJAIXn+yHo3WnjgumbdrNeieJ6
Lbh29FL5j0+ykbYdEwpxlZW4ysyuwDdjfwRGaC6uWqe7RWDLRaDE+EESEaiPZT9J
onZZkYE07qxCQ/aKCw6X8Eu4EwGUq/lHxhO4BMdyQjbz+cDpdHnWYM0DuSD60NPN
vu4kvy2C21H0BUaJuUHU/TpFLejhsWvs/T5lyQ7J9OPwWiJQ1yeqrzcOJi4n+jSJ
id7a20Y9r2e9lcYYICctRAMv+NWYdC+TsUUN1+5AtbFnhAW9SltPaSHl3HZc2TJ+
ow5Fv8GskguBbVG0JDxPVWEtkwXSHKwbuD4b9enc0f9mSCK1NFR/3tj999J+JBPn
AzM8PZfgh97W5jD6nOTe5ZVm9mSf6cQ9Ujh4W9FK3e4/b9jnNTvb1FZL+AFVkLjq
AOrgaOKWTNDQH+m6qT9blTMYgicxtkpcxPOGiGH5EsP35jXVkscPFP6NcUpSU7yx
QvRwnJPtDcyHd7G0wJgbHOnJcZ+4SgLevuR5Gpygg0J4piZsHG8ucrh96mqa0xB+
7MzPHMw79s9rV9OIz7/eSceGiMe0qZKHxopz3+cWhHV0vyY78ckahu4GazFsqdTL
aglI1SBeuCSaoTSKvDn5tazUAH0b0aWzAWYFO4sUmrAZple+sp0VtI7y6nHgal1Q
9UBgWtai3uTir9Xqan/7hHXQyrFvdiOTAk92DB1lGLAkBNsnoLelo2CksUAIhrJI
W1hUAzWgpGmN129XjEf6rslNjaCMVKqgCm4qfXMd/FKqRvf3Vu+ixYkN5kWcPLWi
I0ZY/jwEZsA1yJnUSY9Su5rZaXl1xrBC/UqBy2XA81bRph9jXp4boh1ytAXdFM+n
lF0kBLxrlo4d2/JQ4RtkDKIX/gXDQSOWSLYXdpvtrO1ciEwnF8olaWbRQ32SaIju
8CCzqLhqdVkqjMvxNiv7Ds7edjYRmy10e/PzG8zg7nHsxUnoGVgJR1gfflGUnpTp
8pdKSsl7gNZH+ZjC0y6/kPjCgUWG9esfmpBBvJnexclMYLHCSGMFI5RetvSnQn5I
360ABmzKcQpJklw/O6dt/7LGsxaMa7f2g45ujZSsVnUo08vpnkUx3vvQSLkr81Hx
EZhrH9Z6hMnMw0Sh/gkjYDJGpnPQQPKjXTsDNyVJb6FYhWvRspNDG1kgAA1vUwo+
GUdSwbWD8LK1Pw2FfYNO1sQU7bRDI4B4kiuIe5FNUA3YEKaZWh7AwUb8V9vhhrqe
Ja9uP96h+BcfQO0HxHZCJCPAUin/YHAeLqMcJoJ/V3ZPbmGfIy9WlcTuayHoo8Gb
oIEmZyxGvv5gwjfMEJn1rtAs3c4e6vMVGv4vCSHCRy/lh3OpuvulmMaJJ3pXrPRd
rS6Xx3WWbhsOX0nVwM5sIQgB2SJnK3bOaaTKQE+NQmAlmBZScky1sIw5EGR4DV3A
XC+4IhCyxr0bsYtB86SrGaAMj+TkQQhwDNcX2F+pDmsi4CmmFv1JGEnttS0//GHW
+gHF+Zrtpkm2rIaSZpt1My7Ra/7V5LGPw/v0VTAg8TpidIQMJFbkyVxWKOvpT6D1
UeG/ESLJxeqilGs+bzdpNhrNdQkeX2FmN41PC9v/TxEJxK55T9AWNq9Q7xkJHXCt
8BllfX7qsGNyvEER27Q/0mwruAonDhn4y9jkU0fVnnxs6djJCqNKEecUIRyHAqOI
nNTATm/rAj3kN8n0l/xzxAlXb/b24+9uFqPvuzJcJzuCX09Rm4b1DsJ+I2KBH0bJ
SHAsMHTHIEBHXDmO1X8uOelhfcGW7uTVTDSO+skbLmpJc5OpoOqZJeaMSr++9kfN
oYQZBo8ZxiNbXNmvaU87RjtxFXuBsG/GvfOK/CYZIIUpIr5+aw0H9RNWVQAzDx+M
8Y48//wz7or/1V5mRj0mwJIuz+7Wv90287OCgO2DKX6X79C83eFonbQVCHwya41G
8MUASLV1MClE1o719cCdWeZv1Gr2payFLzcMHDdVunxdQ+Cv5GZ0DpR2Y0BeBA2l
XhABG6PoM6l6mII13jWTe0wT0+pG7JXMCE+2jCKqnEyxOoAdClXxMleTGvz8XMwt
VTohKMeZwRc52VHyU8zXVJtH28y2OdueIPcKvIipZpk5fp/aoiT6Eq53syD9W6ft
pJ91BVwpWq97woDQiGFE+hGfAj35B04im5Jkjjo7aIeUjZTmrylaOc6LSnb72ddo
4CzQugVaZzE3qrrKKL9FocRdRZae3gnsjH5ndNGcxugAVPOmXu6U2c4QZpy6rxgb
B3W30yx7/EK5XVihLl/FXR65gbfiuEhvkUxc59+OdnGgIpwfBEe0EEAhaKI0jFdp
9Ps3XcyQeZgiDnR/J4qoRNZ2VO++y6D48r8lQi0gx6HEwGjPLmy1IMerC2ct0Tk1
LjSwBQ1jfaMYeXZsF5TyUQYTs1en+9XD779t1CE0LQsuHYVXbYF9H8790JB+SH60
TK43pFMr5OqwDlebhwfk67rcfkN7zAZDY9PVWClsIEBK6y/QWpjlP0vlr90GwNA5
/qge3MmTmnPHULOeLZJhHWDJdT9q4LkJKtUgDAFj4L8JRdffdOrnPXff2E8X7Sb2
R/R/GwBJdODxG0dUz9pRj4CLsXpIQ4uMCdUuNtzlqHVhkdUi7hmkOusLldqreM/H
TSF9hGK/t1nmDlUsdDZ9BrQJWipFerecZj6ZLL676xZnIqvcWAh0a2pQTqm8gp7o
aHwbkcj1JCL+DWCVwhFN4ZMZdA02fraqbeBEiMW14J+EWILSQVyK1ehiBPyNx9MB
9lnWDtBmN8RXu4dtmyCDAztqbDP+rrdu6k9rCWlryf9wZwxz3tub2p4vz8naAzAY
ObFWRTC7kJRMtjG6Li1UAtipmNH3Wt+lwIRikSBtp5Huj7/37vVwQ44gARxQkyPH
GH02CwavTL/qMpHTK0sMyXAsW7cMLd8oqR3QN9rKhgFC/RN07CNGo/nwWhqeV1tj
y5KDp846DrRETLLQAp0t2BRk7Az9b2rXfa+p6Eogk1bgb3QBoJTAH8c7cdVcDj9O
+LiCOEjdH90AxsjlDN/a6oqJLN5yN+cKHQpolXFkcSKZ+ulK9CCs3uuoI57qwNFf
x7D39l+HBcxWIbn8HfVaEizZ4feXOWqojr4Opkw6t6CwIqPioU3bOJfRPBVIR46d
jmAT/X4sk1db8WaLekeRLb9O9ePuzY8jquDVq3aQLAYfbgCWzDUnUDbiKW/swxfZ
JNE+Y8KQRJh8i0fJUw/IOXcOPoxRAcKjMWrbMvTXg4picv33y6cgljgBBiOaFEoh
IvkFBgMcoKp/ebmu6FudF7tyrCvE206lVr8mCLXIGAhNmqGEExLsr3LNfMj6e/U0
+IvXN2ncnWapJbzeEUW1phXKoZ9qDbv9PkRDRezEV+EB/lTJnXqcK4o2atV1TPzm
DFIrgIeX4PIzSRHrxlTSZgWn9/WqxmlHbtITMUijMB8kGRjGqJECMeXwH/8a9Z70
yILm04xTHzsUl6K3+47CivvHEqW3hYZilTXGPKy7RFIrOnE2jmMx+iOHcus5GPeI
vpM3UA2zk8H4T+boyiS18dXbt2TX904fgN393E223UTpEla7UGU+UGbO10CgGI9h
fHQw3yp86zIskkwQh22awzjT6gr0l+ab5k0ZpSLDq61Br/iZbQLOxppa5p8Up/yo
H1J/Ia8lhKNY4ovQDVCYyfeW6Z6K6qXJVGlqIHHbF6dy1gNnbC7NsAPIfsTmCQub
9J0xuUHXv9Afl/b5S9rdf5wXexlrFzZBovpaQoK3RfUhx19Vi87oAqY0SW4w/yLG
duTJmEXFNaQeSn8s+yg84ArI0P7N8bEW4txHHuLhqhKL/4a/hY5ZTW0MLNpv20yL
LkXGANWEWC1ZDRu1PntLpXiJa+mlpgxZXX4rier4FauTNzLn30OxN7Z9qZ/RN4UU
MWejFScL5RS3TjQ6rvjBYaGxY2Ls/8XG7tH84xfz0aGE84v+/Yk8kiXvBvsfKzix
NBzIHz0LX9D9eANBzfCwzj25dgV9kSQIy3pHx8g3nAj8ZD61vpok+8RTlMobDKco
fz+tIRwSp+HhpQVCQx7qGmOdGZUObHPHtYX79FYEH7j4wkBcEiGwboB3iDTjrEae
wENslMs2mFiyZSV9+pdYDPQCDn/75T3KIR9ArnN8Po4gL2zbPB0G+GYdcyuUKymI
VOC/0Bwi8T3lbHvj0d+9zkQcWDvcN3Szo5ZyDu7Z6JiO6oTf9ITh52GHTI+j2L4x
hbuQvjOGjmvV60S/VXmfJy9P97RRzMSg1GtJzudVkfdGqMGtR5hcZXap9dd4hhYc
F4nSsSWCXPUIflN/dbWk2yTRrMZ2/D4/QS1gJoEhmG7jKwAQSZYeGkOBWDA+TdNA
j/PmkbFemfoZ5gOZkWVghkmXCk6Ntk6BIww9TPWoMRDMtoQGbbfToAoCon/Xwhz5
mN1anSWWr5ev/BypbyHGE04pgWeJ+UisISN0s3xkp0fcvOGYSLqyzXx7MQwVHn8S
RGpNJHwyimgX9zOYyc7rkBu7Jq6USiWJ/CDp7GcVprdCYCS22MQjC3Uaq5iBXgO0
lcOs4urxeErt07/pH01NhQotlqP+VlmB0WHrhKtMnraaATUbtVoE1NRoXsO4Cotr
uGLFkU52VgdM4CWZCleFGo2eEpvAKjx9t/n9SncYKrZsdHOAQLXuXUV+OQT2iUAo
62YtXNOTPAc+gKLtwT0MRHIIkup2sNeBQnm73c1SvN8OKm7/I3dQ5qVCxJZn2Vrm
iUInObveCJUbYqPMynFQKJvqrAY8mXsKUaWRxFEH2Kecx0DJwMpDtyodrumDIX/m
2hdYbyt+eEOiYJcM6D+HgLbOHLr8knL/4hS5ObewxNg87hDYwo5yUkbyOyOx+BXk
Xah8PVBIn/4FwS3tkOHXacJgXBIVGoylOXcC+tcOu3ek/eex9Kg+xmAkQNuPEZl4
dfYIkyG7S8QqYNQpjG6S6XJuOvrD8s8xeHcmjb8w8QksiEbUMmVLmxcu1X/wwq00
+hCiEU4VtJCM6ZddcPi7TLoBgEqluVOHcrfatx6VNd8abLUuGV7ss0DJ8nEz61MW
zJVxI8lTnHjFVTzpEv7fqMo8rBqYRfPczOKl9f6DdIesmlWi/S80kt6GaDI/+jx5
Lahd1S/0WPgApmDG6fWQTJZj//CxF08pZms3JdcYEHAPi8wDsAPE+PlKPv5/+wgD
Yv/kA1Lxfiz7Txfzvav52Pm6i8vmXm7GS5odvaFaOpfVwxOCSG0jAgGPvqeQ9I4W
5/EneNcY55wIwxbMFD7s7EI7i5MzNdj+NomWsO+Au34zTqx0DBjalrO/ea4zpNU6
dnOvwfiW7uHhUMFr9Mjy8yQ2LjdP0WJEKgU8/BVMZ1bamJxeOMl0jocPuX+RSxEm
T/jGsER/lgxpEFtYFmsF13ji9+ZgNB1P9x8f1eyIiYg5HJiD+bzwY9J41aeTP72L
yBwC5X8X5cB54+BXuxDO0RRnBMj/wcXjHhm0kL//ruzw8QJ30UF4XUylT6CbJMby
69eMhXWf5FMfVgvJsg7rNxayyT942JUcK6hAtWEAntRk1/STmkeugeCjleFj2Dt2
qNWvN5Rg8lPh3uHQ07iQVjTVxa20GEclagbOkzudkcL/oLtp+3BXEMCf5QjKvO7R
K7q+3EBJpWY67fKLhx0Yfj65CqsYMLMI8HbKHgEAf8EO9zAkzpj4GcR8HHow8TMi
3h2SE88cJXinGs7quUq2NmGAYCBvb/qHC6hpEKd9wyDWmNp20y6LwH7tzLygooV7
xlvYL7HBT9Kvhay+2azJp+PhVIYdhBfprQeog3xO3FxAXrG3DiCk8GFTChHsoVD3
/y8xVt63DFhrCPytt24Chk48oCZchy3XBLO9di4wHyTph/WDAwtV6TGrSalqiBcA
NjzWpXS8455WRXj5Pik/fpiaSTk+0QFqjG9B3Fxry8LUgHHZbTftV3KkUCCUl3VN
WSeSyYE1jNdx3ICIaHGzUOD5bTGarzNOhAIrO5RchFzswogu8mNgr0mXKW2lHSKp
UfMM5VeDo6MdYcalERyKUTsur4AZcKhqxsvqf/EJ7Dv8cHR017vSuwBARZ8okCEg
KNZB63A1UZGWlq+xVP6MF3X6RnrwGoqEpxy8KpK07js88t8u0JxcI8v/tCHiplaw
Jp/7w9J1U7A6k9AEh1EFeT5F1Q8IUdrPdmjOnc0iPPXJxgfCM5feZVBzj3ChLlAN
QKDFKgPh6XPq5LJxUq+tSY6BFqQkjJgCBfptrSl0kIiT/Ng9rEpcmnsNqmIO0sAK
7lSjQCmX8ymeZt5vvQskKRpiorcSfvaaQdcQ7DUL8APPuixYjmq2ecMl/+a8WRXC
8UDlmo1BHFD/FBfywn7Al2ZmYKy+C6e08bRIkSNTfGzOkHUwv3GUK6F0TDTAdhT3
pAhltjWrtkraL4xDzwKuhohHi+w2q7+bXy0byz1JdvFmmKHKff8u4VyZyT+5GHRm
d/zqguy7KAgRNANz4YQfn5loAE1KEi9+UFBzZcEOIkr7RY/bviD2xg3FBrndJwn6
5znId8aYgF9519rq8SZIdP07pZ3HEX7aktRsfijdprBjMO98Ak5GAx5SORiAQXpi
XXfNwWDgqvw7M2vGbZnZZbhFCIY7c3OI9DmNmKLWgfDd6CFQr6Zo7YyiaIORagbc
KCEKVEkbDXq+hxYGNe+7FudVPNSuljvhk1NYBKsKlpAr1rR74WWppSdlZxBiM3Mj
4SjDSOBIkHxOaKvjbKgRhov29tPPUlXHwmcLzIkL7Tdex4Azlo+BOecpt9zsuAHc
/01vlehbf9fgNmfwCVxaccX/8RBSNKgeBcRnYDeaGNboYce2qUVyGAUyjeATUNsn
ZRq00NRNqr3HECSFYLw46jzkG1ljKm191eYzrtWD/5hkycbXUfmj4EzLB9lmQ7Fe
h5Qqgdnm5XXY9v88N1dP9Ycm8OGTzu3QLodiGez6G4A/nheXKvMkVykdMkkePWDX
0OLKDu0Kw5HN/XHY1CY4f8/8k+QIeZcUsoD5LeyvsGH9VgJL/fd9A33p2Jw0vTy3
vJBCHS9eAgP01EYWBJjDWugdmj5WuxirR2i7PVVcpqC57cewITcju0PdiXyqlLV/
SGOAncPlu4Bnr6WuvhdIUTElkEUCDaTJljPj1W3qBS+nCegWm+Np2R9AAFfYYAs3
0ZL8mwfTDJgj3j1cSqaxK60XegQAp/znk/ykcPK+pzgikwfeLvtkvLQ/cQBc1V5f
zj3Lge5FG6Jc2t5QPVi7cmadl9NtJ6iwuNGjwZdKxaWa2WXnGjb8GGPp9VYeZ8Iv
KdiRQyvijoIjfb2Tz/U3MiroKjWPwb4/uJTFF+ohw5XJwDygPawXjt1scSPE0AFV
QqXx4ATnsU/dwaB76bHmR270A7NT2ldDMsYj10SOZt2JkFm1Flljx/b1PmyGVnDt
Z6zU5uYneWIoyIamjlks+5hoAwkoE7Y1FKe1GGQR0cbF0AbTMnsF1+C/5PLTwH9r
0N6Z9TIuDIAMHa8+ljurWF1s8ZBHQZLMmaQs3lOsbAAIEajVzdeUHFYH/KBXlvRu
rZyzX4a0WzER4Xs8vrIHhd4asMB0W1MbclAc46qt4jyUlFMZv2LfargZYYVx7CBY
MD4ccmJzPJj1xl5prXZUSF55SCFAePvXCbO4TDUcbHlVeWIYDJhu4IX4gneYkEoS
39mOAvhruYM9dSrN3iHTnagwwNcOWYxZr1h1pBx1BwWkFBiaiR03ErtGSuM8b46x
gVYn7m1L9K1mSsdCrAEQnhjXFPJYkl5e8Oj8Yul5p5SaaQVaOpJ3qEO6F/KrdMSc
oZ0TjZ9vAZE8WhhO8dg+VAI0cRY1p9sPcCVU4zToRqSpMxrlzs/hjDAMaY3ctm3n
MezrQZZEgxCqF+CzLmZ1l9mwZ0JPqWzZStCiN/DQRRQ+J+NYN0WzL/OcTMzhDGGk
XIN0X1H9RRhj91fn6+tYLES+pdmvaOSp6ErMKoe6TsrB0EPcuMzHa2azXq9tKVLF
cbFKnar8hLPhvMvzBS9dIuIOoAlDORxtS63x0NBwGCJARUPQS3vC5Idl6dVuGgXH
OEg146DZF1BBtUj9UW+FbVlfSZCNYeYvygsAGUzIpGUeJPA1FB70nJWFQTXyMFTD
7OmpKLGiVaxLPdk2WqGoYMUCvULXcsft/6bif2oqumE0MJqbYzzcom4zf0gFbvyi
5A3Lk99IyOBJWf1LFaYJSl/pIzflQ99d41hpJWAzMUA72AE1WwvR6d8s8or/EMIo
GJGkApP16K7D7Th86xjCA/nYohVowyQd1IukkdIamozmqm66OqBQ96/IgQOmysup
QD3VcZeBnpA20IBMvrhX7Gi5B/mA1/u9CsDKd09AMOk+y2ezcgZtHJ42WPluJRrO
z3gAOowuuVPYztc4zJDoYsqXEJqrJyOft1zuzHRBh9QIwCCx2bTeDMD34YleGoK7
S81iarlxc1CgibgVWhPYcQeNSYYifVyJTZzOLx1+i8m3DNRXzTKinl5Sf9fODWbX
hoqdIwD867PLH3yS6wG1E7WswGVpKo9FOp4qMq7sQdywCgq/zmKpcnKLuEs2R5pW
p4AGkLcBE/ECJC9Uym8hg4l8YnzAWjkjHFKoJbrVF4U8JCUFWM4oSgo9xhBORx2C
PANhhcvSSC7but23t+YwqiRLIpxYOb4nQxOZW2yG3auO20mgkIE04MaMOoSU/Rbj
mBiXkBAebqFPUffW6D578PzsP5Jj/vRhmtDMI7IGbK8t8UaiN5frNy8mFKW9Wg2R
Ht6sFcnR+UrMKj+yeBidUX6pg15TDe9eZatewRy2f0/mbfcES0X+HVEWIq92zdAt
yfWs9Ef46yNJuXsBtK0caPiswAa+NDRBQxnG/thhaBa8lVRx3qMy/MV2uHnY7HS/
EGV2y1kgBrphKWjykvdm3wZF62FUlObbKKI1Ubu1akdM6tJMY9Q1QXF6jI5L0FzS
zZR0o/hntH5mRg/N1tyolre0drRr1qVhCfh0YHuHtsHlMHWGk98BVQ3ItNfiouBR
iHZe1CnBdjDAHa8TPi68NfvQ5qSnz85+wu1TXZ0P8eaQpG4U7KZrQCH1n2avjZeG
h0AbB0yhlylEKWXxcsynxU45tNe4USj8jkaBJLag1pNFDxOtLdUGlmYwkHSoy9mT
1KQ48IySJph/FEkYocoIhYWWd1tFOw2VZMbwgoeE3iV5RwDDGrxJV6lolo5KQ4Tb
+h8wzxrY7BLnFU8WlcySr4zk445Pg4MQpUbN6O7y1WG1o/NfqhCusMfAmvNbZHOe
kOQNW+SunJGziEk/D873l8iZU80j4RuwE9ifWSCarE4EeO4kg7BNNJG1f1Z1PUgo
2b2xBy0RU6UQ5e/4gX1ZumPjyU1+P17bi3uY64zuda12MjdXY5iYmtQCU9GpGT8P
EdE6HKsH6U73duozgKP0OoeuOmOVuZFRrnQbvVoDfOcEpaLNeK+xjHMIM4koKFLD
1HSSnr91leF17iKDgNGL0vpwh1iXiJQM3CPpz/qDfarB2fxI98b1kA8OYk/FRjIX
O80YtIPmtrl+D8yDwrPiTX1jU6y2reFkrp/RB8d32PIoGE4hwoMYYXql3cxfPbbb
KaXYlZ2vooKnq+9835+3Z7//LJhtuLMggJn2FpUnAu7UEYEiQ641zj92WrV8SID8
DV91rxLYn9kFcuIh/9f8YaqvnTRa1ULMID/p1V/eW4/XqLrQSQbF1uQBpoBCev+h
Ufl0UHRO9inx0NQUkcHW9DLdx1Mte0z6hVSIJEX+mIHd+BaU0vMkYgnaiMa5kugd
M70CDpCpSaUXMoPTPqlgGaFK9DaPLOV//ZLp8j/MJF/FA3lnPjz1C3YNn8FqhXQh
DNSl3eoCPq2sG6fk7yQJVUazAELA61YjY8nh4S5CyXzZDDTJE9xDYG7AZ8dEIie9
vhmilZYSWKzrYFpVFDmZkJVNZcUR1LNDWkbv1gKqXVtIHB6UhUI9yRVtSXnhHdV+
XmwTCmkTtF3hqn9zZli8SMHXc7geHacZtc1ZLjJGwR70rC4U/oVyokrVeyXukv72
9E6w03Es2wNa+6y5IE9YxKgKQVrWyvc7hzhkLhhCSeEHJcjKh4NjcpvcA8uTbm1e
Dxs0oz2nA/d6e3PBxexfjAApOXfV5C+2cWjcgjtqf1IOIesXtRufg3FUw9IKe7gZ
PMA59zk15Q5UfMT6B3OShjvaD/0+5R1QKUJAm1b3MSp30z9OFCUNXl1yJt8r7R3Q
l3CiASGKq6l32GeiGhhyi3Veb1Ssm32ysKizSrx8SdoZx7o9X+XoMXnRbTo2gjwD
1wzkdvNJVt6fMFKLIVEdrk8GIZUiVV6wYyeTfjm6uzOxFuhaFqo8lD3FvGADlA6Y
PPvo5Ea6ObU4TbVvIotFimfuQCkbQZdGlB97yKc99V1Pyd4AUaus107+KGmxg31d
mJuxFedu9pgTdIAkMNhbMIkG57i+33IuhLTc+dkYrm7jWpfeugUmG7g8dM8P01qj
+YFl4G7nnJkP25/NyzJbW7S4D0Y8OcLnEDB1bIsKbQ1FZ9mog7Z3TgxPA8CPpV3K
Ywv/QBhPGpFmNLtiES4dK80hWjIiNvoCTMHyugQsQfRaGThukozVdRT8p2AJnccf
RrQzbeWNU4WZQwXQ/yeG/5john/nENsF6dF6Yd32WXoBdq+ic4aIm/clpNHKWiiX
1x1AdOnsisn+qXJi5SqU/BmtdFnN/wALCyDazIHL++f5Hs2yDMkWhTj3zUqwSR0+
UACajnfW7S5VFJ8T0ok4HGx4WzEuJPbPeytVkaONhp+p5XBmI5R55IWcL4iMIgG0
MavAdtCTkRrhoNgS/Kw8gi8SSuwAh1C8Xzz5vjW0BqTTnDJTOEXgnU9aNz6eP3cK
jjaddkS15R6LWIHCEBuQ4M6tGo/514m3YjoErBavGVFtQo6mMQpgF8gi2JWfhxRw
O89b4uc1ZYoQbObsP3o9eC60zs0rqfXfZ4jnnDgyMa45d9lh4Vphrx1fPv76Msvz
B7hzje2E24XcijIXSUfGhPmeDcAoNDl3lGDz+00R6GQltEzbdKmVfeNnZD0xecFZ
rmUkz0NeRmUIrTjf1D5+tHENkxfnPgdSY+O90fYdmgsVCRzksi/AftQgXiweIxVH
D8QxU8a5RwePu0JxNFmJiq5Q88cTC/7/k5mFTTL9LZB7+qkItgj6jNMxcdYDRt0W
MU44zp2es3nBX9UT7yYkHGJrjL76JARW0l/gAwk93tcawpulR/BxVIvtd/HiW551
qUZ4V2vi7YbtIMSpI/jufODbMIzu+Mjsu3YtVPrl+SlF45LmsoquvEWsNQNybWfV
ujQ5D00maSVjbGh8HqDqAX1MC/0pKa7qzu0roolDETeGBOyvFs9C/JmnOBcV5aA2
Bol5y6Krb1o2KhP6hKqN6ROuPa2Xa3cD1wW/hDZ1IMCc7yR3y5IFj3Xjy3QpmLrt
o4WA06v5CVxEA0kWE3PNaERaK5itt8bQT/KfBfOMq7dftj+fH25FbPkisTXtVHq7
brDoQT0hzPSIOP7GZTiqNSZnFrOZ4EHGgPD3LOJpZwWbOyVX2aS9dqKTeFJp3YFE
vtkTraJA/c162xSyWs7UpWb6NJMXZgBfFDEzQJT+zn7EGHoummpIuomOGXCPxkrR
6VoeRCSBF7xS3/1wPia96GE5wiFuisG1lt0t3M877sJTqLzbF6tWdpze+4K6zDit
viis8JEcOES121RvYz+NGAesUoOZeb103ZpiqV1qawrpJwzGSwHr76ydHgAF51Ac
ikUMSmI0habsgm2aihkmUNiynSRpB7oG054+EpJ+Q9uv2u64pvX1isFZGxegM9YJ
7jiD7tQKtty8SshqIqmWoXh3StnC0zINTqcgiXTRF+raQP+QxGyQsGgxJ29208ja
zwna7J2RLKlVIywmLvFF7qqlAY5ue0UJETwOCZApobPLNHJVoXIEFaMP/ausdoFA
SdHw7D8/8JAaHNA9qGq/xqXeReovqWJxHYoc3rpUg7LQzOXxiUWoySPt2ekbUUel
SExhhtxZoHdwMKUYDY/Api4MrPviobmE1fofOH2k+RYeLfbrzeCcZqQFUnkQxgY/
5GWHqWAzjjcG/MXIpZmABcSvwFCbKypcSLs2ZeSZTVyX/rFjR6DHH13AqAaNQC7B
HSc+M+g95lVmb/Xwd40WlBKH0Na+RkWJvZgaX/y2n9Lpmxa4Fy7rvQOJS5exRnlu
aTF78B9R5APfsLKU6HTGIvhm1RQ8lK/yOz61kreJo5nkcFVCHPdZUmWC6IOwtLRA
pNiNOJeqrJ2xKVMkblrPwG+nFeILWUELVDrimpGkZgXUHHPtQWMvOMBKe6axcx/g
WwHsN1rbQ9OZNILdeYsGxMqLciTSrNln8osPhON53LpamL5dvaYdGEhLJjxnAo7U
pK7sHvTwwgtcT1/MEqlDnWlnKSOYrxZVpg20QY/k1yt1eKRzgKZBy5g5rhfqPWWb
2yWeyk9hXdjIH2c/OXQPnSSjhQg+21jhJUMb1LrsV7s0hkNAanCSGYPWXYvugDJc
KJ5Ux1tFXLhZdHG7AWZ8HSu6QArnJn8TBKMDlgVMxkt1erEATCA3zvb0iwizK6Ah
MWAFslXfc4kPes4hCcN/AodX3xsYdhLVKzajwx/OqL4lRzWAEj5SKi0FAOc8/SBb
muVToijB8Ozg5gN2JhVliACZ/p4dWHqK3DvFM5e3b70OdcXkmQkC79Zf6VzXqmoL
iLvpzhXoUaVFJ26jOlPRGbvpYwPkzLDEoYMR2Auj4kFgVchr6sDPbH9hy0/JiiQb
FgnDeMEcX0Ng4ILHaiWIgN5W4QIweSgqtX0fmlDgYLzVPu9UOr3ocZaweT1S4ISa
c186WUbFMFVykZpLVis5KTbzBkJGBoix2tnEme2QG95hXuzZlHmoTYJAgSR1xN3K
UYH63Jll7TJQQyzg6iPDVLVkqdes+CduyOHfYxx4v1kC3mGis1WhFutaieHpFqY+
H4pfn6QrLi68TlLqwHPDnn6I0/XNSuspHR4+EZ6cyorv54UXjzbmdRUhGXOfLw4z
Q+CY5zZrFY4/ne9LiL1+ZLKlS891ovF6cTd2dzn8d7XYK865/Z7O0HFPAcv2ltl4
nPxgSe5A9NdYW+pbDjLY9S8QfNIok40YE0tIQrXufYEKd0DsEuFmLJOeuQUIexNs
F+dZkm2RdBJey/hk7P/LaL588f9EAMhV+NbI580Eu8xBri8LPHC5W93pRL1AFXuy
sJY45qysxU6m7d3muz8sMTILAJr3I/N7XS4EpnUt/Flnyo8vKchIjORBoMrjh6O5
S7Ot5xt7blm8RLSEh+Aw0DV1UBni3x8lmHq84EbAcpRsYWa0yGSBxYG4P2ngw0kP
JBHLQ1DPoWn0dd8sn70sbmU8n7/0WQay1BOhf2bUe2YeA0MIiJhBy6ElXSNYtK1u
K4kMkc+3VUUdBMsBXGYYcyr8yaoe5DKiEbacfkVf2224jPgRqDn/xihFJ4YGDk2x
SU9xDRosKYnL+rlesp23bV4JSi+9UQBL86SggbOuImhvyKTQkgcZx31dPoY4dlCc
eRdbvUJJFYcz9Ru+wMfxXtdKy2f+SWmbx4nPzSUyEUI5KIVIsEs79wtyl0KmLuQ1
GJ69w28Pmf2yfR5kJm6Ajk4oq4n1mfS8FvyFudyrcJbaZ/7UsW+/rgc8k9USBZhx
nm0ghcmgLJ9gFFJ1qA0UsQZyAEa6QF+EnQIL4kjWe+G5Pv/Kmh6IXrcst1z1j/HF
PGlrQ0qa4f0o8PrZD299Lw7gZ9pPpFyQDWOGsXfYGPu+Ldob78bQoAnsQtN2S8qy
9+29I9yHJlQ4PyAuxl7XxJBMW5a0gR4Z+FyFh9HMFvyt2QWoLfrk33klT0uYTEc3
7QhPn6V0KaOYuDedxnqaf2SrOPHDAMnmfjgkiiDv98rdtcZG0HsEZ3SbdX9+XZme
hGt9Sb5ZfwWmSXLJhOWPo+b3P/9hX1j6UhKxhn4qriVbkq02Tv+CklquWdo9UD/r
K5167uIm34C7nRR8svaxuKAu6OoZbhQYJLGnIuHI0m68a9LVKshCO9EriE2wOBGT
j+0O8IbY/Jynu5T64e0q2/Hj5aYcrK5aHMluOqEHNbir2NXwjiNwfVHLjsacrJbn
gFgJbcfJwHZmzAxJO/lbNdJyOz3sZsvabwfmUsnX2gMsWMdeWdgOxQXnT5Vpq5m/
bQ/2iID824KP+3D6yYiDgS/1CPJWM5BhE1OBgHp9e6r1A8l7zTjlRHVDPF1/ZwfV
iCsHlpxHQvzZaSW7jtKBfOyjAiDCm6FRTvVxukH13RudSeNL8vyGzloIX+AkVEDG
8u+f2NngmdzB/LQZIDFq2pHNUMQOQqko6KASUemXChClicKNKaK/tll2DAbMwq39
lSi2ATJfJkTmRUYntnNh9/wRn8nOUDajaFY7ROXlWYppBlp0Jd4tnCt6sJobXvuZ
Otxqd+KJvhHxsYYwML/74m60bBEZWCTrVeEdcVcfQRGkPhHVtFKJs05mUL2FmONd
YI/uMFa4hwCMEULkem2oqADuQ09q+1fqWokGx17Dc5XGNBi+9GCDepcwQDrv+WK0
H30HoBALvQIRTn/IhvyqCYUThwXHrW8Y9cYMZ+bsHwvB54+OavSQEN2jP5HDz6EK
KBNcIGoUMV1MKewfuJqXHp8Q8ViaNigE1ESz6Pu7n33EoOHGmjQhklAmBs4hvYcb
lLNC99LkMQYZIIp04/W4B4zeA7v7nJlsI1nXE299eF2B++M264ttf3vkLlcwLSPH
KUZ4ulp1zhXeOI8nPttUo5abw2zPHJEA4DvvBXa0R7uFWK8xvuxzFOAOO3AW83br
Gy0Whq0t0PX49nPheHrJyWIMSPJivIKnc2iqTYD0iesbJb3IPyN/sQGM4OiLArA5
ZViQYWdT+Wt9jW77oXDpHfbi/hDu45jwsYVKzyTT++iW4lD3J4EojaOxmFzVvkQY
t7sykE2OjrCt/RNX3aRS9KnZjzPGZ7vz2wkU00z0l094Ow6RoBjZ6jGyWwcsf8YF
IgXa7SWlA79doIt3kdKc5QV+OMXWrgxZA4xsgiN40nxVpJSbVG1zd2Tcit+QLWwL
A8/ak9g3fHUx79hxaLcxtCPd9NHMu6pkn3h/nyyTp2ttgO69Zc5Cnulaq3bEQ/Ap
tSA0qXzKFeNpiyv0tvdzqVIQRgOQqJ1L/JyPVTUqV24vxzXaF602iKdZ0w25U5Bw
BJykOVMFgZxeGiamOUDjP6TqHQ9JB9rpjPQaRL379nIIP0qxjCJlqwPFm6AHhA/X
gLLMyjb4TkEIrjDdjCc7WAVKeuq9FoGqP2/CWLfrb1KZWB1DQ7qqj6dxx9AldDCP
6mr+6hLbHveK4lXmARCHStrlOl/0KjRfQ5kKYLWcpSioG42kH6IXxmmFBiHwwaox
5YesY9G88dEeSIqXf5PkAjKVroWu5yJlZmDGJ0J3UZac2yXAerD8TFwV0qzfKA6g
gauZZ+vk+h61EPRMQjah0Fg11aRgYqzSvkhBxN6KQIaw6YQFKwm9h5WlV2eRUejO
zE5Hl2B6iYpfK3EeN5eiYT5V4N0nEE/0xc3bPRNhi3J9HxofpoAcqz4Kt9njsDpn
QjEwQvgdYnNX4g6Ih84n8rhb/UqOx7ttuXgmYu6mSo9LEi0bZcgO8wudkNRaYFpl
7SEJxfgtEEstqZDETs4ztjUKFPiMpDlEW9D3PQ6v6IG+MxYtw9J9ijHfJv0FcTfN
iv5xCII+NjVhm5gj5atSLp383Ja7bDBOy1lFZ9//IQLgkhDZaTjx9PC1ZyHLFGhf
9hu/itKyvsLi/PCBK9DJXnE8U2E8T0hOSyk4JXaDUwoc4fHgiCODkSk3YICEt/Pj
feX6GqReCVyNZ924e4icq9B6uSKZzM0Aahm9Xo2B1+BROxOeHNqhYN8FenbpmWFf
2pW57OrurOumlggMnKvnC0J8TSVl8eN7ZYrMzvyzsM5hdoyeh7Suf84qethkCvWZ
1sUYEr6SITYFfwt/+LNbHQFdAFra16Dx/aSXunPddZGUOym70Bh4wjvc657w1fQ6
CoO+hm+rrfktK6vxoMHH/FN8Kd3X+At0J2wUczY4AEfPHXjOVYLhemBKBNSoMytp
m5qmp8z+o3qo56KDF/Td7pN7lR6RJEnc4/qUsfO41FPASY52BDcu5meG1NwiG2Ek
StjTV3PzxgrWuUfvysiSAOwJEK/P+dSTG8cAD4pTxuqZiNeShglWfnqZ3ErqOibx
uDZCAMP9SLwc7yYzxvqUG9Z7FN4WuE5umMVxT+NTBg5h3Q0k/KSJaa4ejN21oaCt
l/XFPfIQHDpuGZQPAPbv1uWl7tm9/6a84IZoV5gC5boSxZBBRigEAAK6bxHHxhk4
BgS2RMt/J+MP8XGurJ7hqqs5RLOTj1JNKwTnQxacSH3QtK3o1kfzkpxtGL573cnW
Yx/8nmXdZrJfn+IimtfM+kRA8ZUMynG5EYKKRi3gFEnV14x5VLpnyPP+WASoVf3g
p0VU9fg8qvZ8Zil8nJLW3BNie9gdCfUGlG2sFtJuUbn4NsRwif+JLbutP5FZXN4z
ISIfF+iJJb4/lCnuW0E99ntzZemE5+ZmDLazkCIhEhJoWZ1L3FC34YEeQyedqLMw
Ofc6LMhJDR/D8Sg+m0BThPlP8JLb/Ia2Z9zwC7DNDDivA88bxh7o4VDnADeUBxi/
1D9HF0JY2eaNitaLyeFQTy4z/y8+dI8mR3mQP51Q74QgYjoM0M30Vva0DUcUDGR/
cPaDN++l4h+oWBmi6Q4+mzHjORIORuD4RGDfDR1Tshsa3dBmD0Ish/ucbS3tXGlL
Un3X9XVdZL2McP6MgJj6299StMo3939IxnQnxa1xHx+jxZcYyXFq8i8wmAOwilTN
dVg+Cuk3346UZUG0lYBRlcKS7GEKRJGxNKxzMsVhPE1DeHrnrLxtb38DuOFHxiDR
5jeZhWYiCQ+cHrRfXygHy+iDNXv+m9n69M9m0olekIS5c1/jaa3nsbdWNUKEqC0s
QkvA5vE4cInGR2w2gvOHhgODth3FVN9ycBvja59/Y3ntww++JB/SAZa/iv5R+R5p
pxejyeTZ5q2qz9Gl3fBsi7b07ZnRlAUukjvrZnwfsmbrpdqVeubwZtx7TN819Bp0
oh9e+9xOegIZTiAHUgRu0cQ1StknJq3+hx1fsDanrVW7SLqJqsNHEM7hoSxJTbPt
7MeEKZlX+T+Q15L77iKPWVIv3mxxlT7QmxPlhQ4FCG8A53EMKn0KRzIhcMbPwUJ5
4qqfdif4w++P3r1cedAV/x1/yNRjcLrqYNRQHg5Y8I75A2B15MkaV7GiAimc6PVq
GCdGaDPCB+NNFSlYkv1U44frXxmnVwRvqzsgo+PmZPMXjuKE3EO1712jswGoGGtr
jeIH1Aobq+JrzDIZyHNK8l1klsDTq/qCqRD4HO3SqFCt7QCr+ylh+XxD28NyajmA
ypYf5Cqh4PXLuPchm866hMuETpoXoEugY/M+ihUs3VQs8Ae1Ba4ysWRd6SwTRK99
WKBwWFe4mok9VRaJdDdIStlaOcVy+Xa/CDfu/T8iwptXVAcKd7ocF7E4+cQatMVu
GX7R6OH2d7pyw338j5F5upVbqXJGYkss/RA2ZchIFqQ6FCYkOusZnlgL50tLEvzL
JIXmOcDA3M+sKvH7LbrKmc23XFE7PyaCKEfnLQg+6qm83bt55KebE2xSw8Y1FKxw
WlJal8qte17sw8zG0HACADxeHSllssUf5wyyfgU0OXYFE6USlDW29QFUeeWPEE2c
Ap1Xp0Sn1mEgK34eIOPvaw59ldZCGh4FvArucBFwCtyQtbun1K2kFEdht6bp7q2b
vcKGPx/FtC3yS4mMzF86VWX8rGL34iGqhi2eM6svCi+NPC5cRE2q7p0/CPHi1c1e
eEi6s3ZHIC78i/ckxtOUML7XVNPSWG2oxcL/AeCYPToYXipBWsVqMpIFZS7/kT63
4jf3xgT18CMHcldiHhY73eSjWU+A+lDm5URixgc5kA9hKMHZUsL6yidzF0TWsZFh
e238n7J01tBRWe18wscqxez9A3DFcO3W3b2sVrF4fcEAzo08awxnE5u2ooZvJrgr
chML8/wJQp1RPu31Mx9cVeaPD0zbx4WdOrF4AmoHP3aZkaXwT1luNMy/LxAoosKw
CkvwDit8XUXaFaN6X5ppywyrADhSP1x75IJgfeuc7C3fiJ4s9SwC5dWJF7mbIucY
CWyMuEAZ2ReFQGWG5PzGSfL56WhXYjgX42nuXT+B3l3mjxPgQwgADU4GZD35Ogl5
6fh6VGXTp7SjNfTNUBW+RySMPf3siCq58q+pvqfpCdwY3RiEAF4ZXfsBOM5I5jaV
ep8QEEH7WPgIDM9gCXK8GrBRZ2VQVcGW7AlSqvhn8XOuhzwaQAmplKRZ5+ehpSwg
bEJNYolUsOn7DOVrESIg/cfGD/+Mh1J8jeU6ONhx2JPYTNYz/HJvCRJ07i54dLps
V3LjN5l1W1d1zl/Q5sGxv0nO36pgmGAb9guzW0qDm2cWaFLnICopp0l4zKADYPBz
3Ih57m4LwA/q6eUR+OP5uQYOjM574ex8+DbXxkA855/5lQnt9wzt0sZMfsjjBJ9S
hiDsHQqw4vNfEl9EGb2MO3Gf+zQlAu8QMDz2hcPH348xCkdF6b5yD9puWdgttTgW
ItH4RFTAgu4qQQvAp+p1rMRrmFqmKj+1Pi366PCGf15WkqFqNlENboykCZ5cTNkr
zp9pjgOrmQ8K4oNshE9o+crCKcjBVs15ZvIA5k7OkzaC6F2hr6CqFjro8D3jkfbo
mpTeJz3Eibs6yXMBGV9Yna5LaDbw2TpgIvJkYZdmP2c8EnCFO6i4VnQfKfkK+In2
FUSL7mOjHm95hmSOoyQo+rWd8D88MAv57tpwr7WaDoYjl38B5CMTJMMkgVk5DWP3
4m+GaifWd+fMJ0dMe0mU5YH6liKA71w9aD/4Ms30OBzJMIp/vn9xO9s7qcO248AN
rsP/90lc3IFyxxT+a0b/zh5dpoToxenJxqaMrHbzguv3TygWLYZ+6SQclfzNzJHT
0KjvT4Td7j4/GOJ8WDSKmBNDHFeiIYh3p0CYg+3V2DvjhhLJAY79nDbCLijDNuHF
qZpfQGz/Im7AUUfwpgafKlvUdUgyb9se/6bP7PVSJ4J76+4cVoD/ieo/FHQQeSPk
9Ko2ffSWCstjom6lAqCi1BnUAB5d/DEutmFqU82QUkkZlvqULvESnRyRrI1HNb/9
+L0mNxrKv8N8vO6tkDL3Bd5l7ns0bEgQJgnKTEHY5T8lSGSUkrUUjHDZl4Mq5JO7
xXZRmwKfLZKSVcPrwWxfrCfnY+Xd/UgphQB3/CCDMc/IGLJXJilQ0q6LBrbiJvpx
zCExqF79UfDegbkyFzFXRrpyBaOvE0djoSfFHgPB6GjGTjPjfVI19qYCFgQiKF32
uUyfUnRFLp6Evl1CVHQnYPmBhWx+KUM37mluz8gsBlnQR6ZZmsxFnTyrIiWTU5c8
koyApuPeXsYz7qR5rV0qLYhHbLeeh4GoRqC78PGI1BSCyprbdB24BZAYTtrO0zY5
C+/dBB1L6Mh1CXwk8RNj7PJ1/NnAXpEUlJLXJyKBf/oxaI/nrAUlTVfBKxEGbtLK
ZYpt8gCNvI7vaQMuiz5brKNUU0uM5ZXehyxKGqKrx5LSAlQxb7Ir+m83VhAoeCG5
+YGLaJMvmZEV4vCUdUN1ziSbhzwV+OBMn4Rz4xMFVbw3+4yCqEiX13EbAwd3sRQf
ByOt5LmYYhKvutNT9PzzN0nthaRgpefZFYZhrV6FMQc8jKdmRwfSpPgvSCOeKF8/
l2jB2wXDwFPfS2LifoUkZmxM5ouU9ecscbrPI10nKNBXtlno9t2cmF/Xjx+ZIgbF
EPSN+tYeDn/w285DgvVYKcFkvLur9xjByeiIGD2oCQjUfrLk9isqKi5iVySKKBkj
47MmdJsct6MvrYNMa+Gk3kTdGV4OnlZtN9LOh1mnHDgE5IkcKPfZYib0M5YzJUaw
oCCHXiY43JcCKvCD2UNHr4swC/UxFs0W78dkllsRl91rhPJNDtRNdH5PpuVSnxUg
DfNwqM0C87eo024LK8sYK7/eiuqt2adZSyADkCtVTcQ/aC+B+i4Tm+R6iEozRRM3
hqyW8rFtqhQCSd62C9pj8Ru3umbrYASLqOTB3bUJbke8YUrKwXN1i4jqv1oYFh1L
2h/czOAjeTRlLxwe4H9xEu/qsfpsSJPa4jE+9Cu2Yv5rYy2P2oQY85thqmmPELT1
TjxTYZbKVVx8/pwKyJCIi+H0hM4Wr0hhE+wao+2hZXIdhUHt2s4FZlq+3S5u2fSh
eZ6W4Pbt0Dt/u4+1YPqqiaiP3OtLtx5kfJJzwHrhgmF2eF6MpeJNdKOWy2zFgDre
0Fw9ZbPme8oMyBoavBjE5lLZIcdDjm0Ygc38yN1oqE33GgwEuVK8zgmRWNykGsBj
rRbzjs2W3+GVsMNsLOian64VP6V+qNZFkEWLNeV3NeWwkzLCzcDxgzXhhNuwW8xd
30d/LYCQpze321axJ0mu2UIHWjAkCys/0zbPauhXybyaxGrmcN8ETNJSnIuPEC9t
812sP20P5q++7ofCSrmCKhQfq+3b7xpc6HBGciWtFGgs+h5qGiV3K8pPHZapSv5C
JRkbpB4yL+65kPEAfaDuE+qlWggZo+fKlibgbpCnkj1Jjz6pdll1kJ8iUULcB6Fu
Fh0LlIT5xUePEo+T+HvAXP1RecellsIXr7ZhRJSYHNrdHU2awVbmDEC6Wnj3UpJN
XcFFM91JYlFOX9e/5HxLDE+g3Lbz0oHsBHIGtAx+m5n6NrAHCAGMYFDvCc6bgnuB
qojrc02bVAeoh7E0nIgAAsZLxKo62cZwOPxipYXB2pCXbtZCukhIsW3rYxcCHYfG
jAKHn0mct6qluqJBpa6vcKjMfR8YfZGpD2vi/qRaz2acGoj3c/pehzXZ09Vxz06R
FffZoKGXA2o0o0EOla85z92WdbIfTKuGZwfW04BpCYJeIyJU/Yejc+spp2kSwjwX
wfu7tHz1MhL7VM40Au5Dr01ImjtWRrEpUdylI0058JMvcJLq+uz2YAfbMEgq8ijg
S3L9pTVdc8o9HKimBppuMKKvzArZBnejCKmxhtH/0GALf9sJjWKxNZXxoxqsRui2
S0hfzxjJBLHv3S7NByV3GgxAjFX8d0FovifvTmO4eNbcSAvwCW/mlgN0/CFKhzvT
u39UZslltCL4jWz03fnpMFE5ukZFHjL8llbmSQ/OpzgbPaSszfGIdiPn4kbYxkuu
AwTVwsyuIcKKBfYUP71bSp2ypfzwVNSe7fSQY5riBYTamm8jq7yaCOM4eMis8WZU
ddH6nU5egnJbTCQ/DFTo+LShAV55AtG1nVkhSxtaKundCViITvz7Hn+aZSYsqXRI
mErRZ/bwxa81UEgSEpLk200oyv5fZf1GVX/Oopt7Z0z4LO4yPrYStsdH2P7s6AXx
tv6F0maQItzI6CrhH0WjI5uP93B+xd5FiRX+lCk5p4hA7UIZQFsbouf5YCTaggYR
dpWAXyqys+CdqFIYMPy1ITLFLlwLaPs47oiQQkZ+ca5BCN5unUQ+MdUv2gmyp2DL
gRzle8/wiJsuBfSeebpYQBlGEAxiA56YGj4V0qJ3+EH5BTslbeIrATAP7YnIFz48
+vDM+Rt3Uy51KThFGrt5v4oH1BbuCAn5j7ZjHHyfffi6G+a4XPZxjDpvQ8Mf1qlt
CittMU0mxbOxV/1Tw9y7tK86ergZMl30oM7opdnjdxc0TFWd/4u36YUzBApGFRTz
tHr7vBO6NE/U8boHMh2lfqbe+lMZt78uG5gezxGabnZ+MLnyoeMAiFQ1ulx0kEDI
aWw345aiotu2AgiL2XfqVy7iXWIr8lgYORlUaDLyp33yrtiNR86dObYfv6vxUE7e
j1nG/hfZX2GzOQtORQdABvF2nIN+unhrgVEUeqAfKcPVym5CDGm1ien4iOtiorxZ
fiCS4Vb9ZKq+H0MJBatKh7EiypC4C9ILfSYI5AnaxdAzQG/y4R5VmOIAoSfIIb1i
esfYXvEKnru83wOQ7wRnDK2/ToR3eKW6I3KWqdoHcFuWw4IE4fBqgkMtZNY+1qVk
YcPhklzP4iRnbM2m3dCnKXJweBQOkO6ITt/MgU8L/LraVD6IwM2tholFNNrbGvZ4
cfyULzwZh8Nw4b6nneNx3Rjsf0vQK0V4iC48ilgr1q3/fGIQrFMQqe36vrj8p8mb
TdixefDtTCOpTB2RXaJixVxIdM+cy/eazEiQZ+XKuzi1NYH8HYNF7U1ncRgQdSni
9ZAwnYp+f9aPjO3fbqtNodjXLHMxOsvDxfLljb+V3QXktoR8UKNNkBUQ5x8qbjlg
uAnc+Y+CI0SokmFH2d8ez+Lt4WH0bKbCO+z0TYIxYAHd7m57u7qpTqnursOzHp6p
AJhGNccTFOs1+NAXRSvddDSOiDMDN2LECqhinfdxid3jCMbSh2rh0XL1J4XMYtRG
nLrNJmnVvgeT8F7zeY/FaAbBD4pOcpKekOU2MReLHDrR5ckdm10RmaMatXPUpW1l
K7Js3BVy/GNFjtUvlZlhBUaxpNZbrwyZv5sCp8wT2eJ0xItbGTTcoHSpHVzsIbDo
TtsK9+LmuwDXpdyEiRRsnKoS6Qy9Hs7gi+ocm4CNkomMEf74LzM1rB0ntfdvbJaL
xTK/fuliv29qPfFxm9O1d6sAfv5YOrEAqyJWbzy2HSOQrfMZv8y14aVefo+TV0jZ
VJQnMs0cyu3nguAgCvu51MBxmlTCyYu2UncKY8xhE6z3RAuTObzF6kjGg7YHnQgw
VNcQ/uv5S9fVRhxTsjm+9KNHlAnr0sIybL45AkucD4EauRN63rZBwlUHYpFhrrsM
EGnrKUDUmU0Fwm+aos37JlfhFjSKk7DpilKtoS+fvKVj1/mSSMRO2n53G8vunvaB
oJYnV8rVYMNjf4zmYktLk9rf95ZblpqRTcXYHh5E4Xnz/Lw4aPNICuOZYNFaK9TJ
jbpFFUqa6438I+9RPAVSaJlsKS/nQJdzt2Hv4HqcV2ScEd5lqfL0ZVkQUD6DnRoX
SRxkdxK4YuTnEon4twv+D/yLTadVjRlB8z91vRrG2Xr/3zm59//IZ/N/Cqy4Yx1X
La1V1nYBGQDX2wl9/J2DOQwNozeTBtckNvlg6PcI6Cdh8YdFEjuVpAmo9hY8MnMs
5aaalrrYoNlJsskNNtQtZmABj37/bsMDqnWuABD+ODGaeVso5hbRj3njdMMl3+Ds
WcSCOLGyCMgh2c0hheT+Uh6epCLO4YMrKyyYWoJ/6rQ5Zr72B9dXGbZMQeJ+M0aK
VQcbE47qZzIZfZl8s2JViYG1tGn+I5H9vp3YAYMa9xLTlELydSuShmFONorfrPYN
bBfRlNHgTi4YmXZGfgMfrO4CPKL0sQW9l13lNxO1tNReiYIKF/p+njA1ju4NthdY
g4zhyzsuGOcNZppUT60rBX+j00kDmIe0ATuRA/bs1r2EuQFExlwZUZPwW/dcCIKZ
4j8oV4mgAmNEK1UE+GDXuUthFkdlHhWHD0do1toLoGsYaccDVqMvaTeEgyUOQSRA
2TTH9myUZCKdJhkkNiW+4vVerWS/F6Lx0VG4fyfSTr5v3kcY2zX5DwZ2hlBVcaNs
kzAwa1gUJLfNKZsphwRbV/NvOWPz1PHQh46A3xpVOUAd9iWjs3zBzoFdQtw4vLzf
8nJcjujNlR7a4V5C8vAbzDNQiAxVVQvBwZMx7Qy4W+9ur1ipVNJhQ13vXvrPOSIR
mmJ0W9uGhCNoEGgIUWVLJwI77CDJFFj+JHp7Nn4/TilF18EWrqXAPe6TM3g8lDLQ
6vKrfvmQo1VRkILUs/bRJ3ZLl2hNJLipnQjRliPkKCYIJNdmY3gC8DRoGC7SG8uH
FsTd/HAyVd21FPqYIxvzVICD4AeJh/jnjvMYDE2kbeUUwFqfN2xS8OB+e5ZhMbpy
bvF6iYktWaomCSnAHqoIpxqYiU1dCxPC2SiNUtizetsXyF5BwOY0iBE4uT+wgbcF
qCScy8lcEdYkeqVKTRxGQM/5ttLMRKACogzdVSdgTRksumC3kMarloqxbhv1upOq
oUkhupntSiei0LjiiP0QZFS2rI4P6pIl99A53Z38roQV/O6IaoGY1m2M/sBVLn/P
aulGTezWbZbcXPMS7ahDb4lgXB11OcoNvO6yJayl5fvsZSqWh8/alBE6GqbuPHCt
Xl0I6JWgkaaS/oIat6PtXkvH90XDZgs+Cpt6pfu0FqCmF3lLfhZNN5Lhwd9oxEch
G305ZCqrEtGfNpehPkbidDebK0BqKhMptKK4AJkJzuf2B5Fca/NJasZFW6VJmLAQ
SQY5zwGPRhTcMl9qKC4KX25msXMMRfVHqCGImwWZ61ZyLiHLguBGDNkQw8P/9zvo
qAg/9u5F6lWSKBkAYbuUohjGs0yBdcdttBZVVEx801tKQE75o72FkXpHzbKLj6bt
zv7TcGZKKZOkSmogQJHH2CRYuxJmj6/66MwQLQxMGw8s/449Ycno9oGQoPye57Ad
t030NyHDA0XfgNlif1c0cwbgNVWz2WZ9ShfRk7KQhMqUa3+7FgGRyqbX4/wQsDmP
jqXCyhdyYieeYmGdHzKEmbTnjq5DVqsJVbxpVDekkpTsOoeWNBfIUUX5aLnfc67N
gkwmSs6qxp7YGNe8K8VCptv06yhxue7z0jznWrY3uFgKmdChNZlhRZouT1irjPHx
BTvItFNKJaKtXPc5x4Lmw3paew3KQptV4WboksFSeZteERXMhY0U6UNUj0HrBCeQ
N5gfrGeUVGZdjRKeDc1IjvHw9tYSdQDuT8rJrPWRr+gVUQTa9DVn8QO98pEHQ4oO
zkKtf3H9u497XTK9quY58BdLZLS00jmMe9gDRRcGsQ1Rdgt7541xNNbdDeMoHwL9
UgxHQlMeAoUEvUwOLiRFzwh2OpuiDdGgkPj7aqGqH/9axmzo0Kme/ligRbSsxTS2
tNEAyrjElb1UPR7nIZJFTXN7RNGni1Roo9u8M65evnIum8K7XGVVolLfK+ipglHg
81bbO5qFE5KtlaNtGJJSaCLJoC8Y+iOyteTqFB44BVXzmBMr5oNOOiatc9+5NPUO
E+3qMXrfVUjN6Z7IrJDBAMZaYaPa7BODogmFk/TEfbZZ+LzLstCepv7bq7wRRHZ6
s3HZq2ufYbtQegjC59QxAJdHwKcIwNnHoOhbNYKRZ9iLGc19EznC8r6dldwwGeS/
fjMjOxFZLU5HK1mRUgv8A5ZXjhrfeFg+oAkitgwUNxe4OmFXRER3DE7nQCBRPqxR
cNCAvlQDoi+ICeeVHCiAYxGpKC1/g0hqFb5ELtVof/F6sPy5jTiA7MZ8qwYJMknH
PWzzJQBK5MF2Srebpoz3VY4nbHiz9ORBkDv3mY0g7dzPGNVkmu9dJ1V/vySazd6W
0mj/ijQO0Gr/+Urk8rWxpuPif27uX97f3mUBOM+PRkXyDOpI/3+b5muin0dwySva
83STn7AluwIvLzgSeCpjZJqSgYrnC76FUAqov5/DeVMpHUYzIiQ2EvEwXYNTze4S
x5oz80sjDxQefbaKuS0vWD871yhsskATT6A7D5VsS3OucqkzYpUlYPVDSoOQBdkP
4EGXy3Dhge7i7GZaKvwOyLJMZSo07hiuzA0QUHZsd69nMalfnSs+gotvqT1hvWP8
bgrh8Eu7c3Zzct3evIYDepaj31B2zbBkQOYvJTBNFu9CyonuTs5ImK63q4IbXMOk
KZ2Y6h2EjV5yrWZ//HpW9zO00uEvDa+QL41iuPuJWUaf+U8v7AaJShxjVfXtKwTo
snpyaYkZ1sxS+1HCxm7Gs8smX3fp8kQc7A9+BIb/Y4Q/yYWjberCQdyGFtDxANaC
GFanF42F9jUNsvYrH19dDRtGGNddh4lmWSO6x7Fkne4hAIUlMkL0OmRuKXJoQiZf
DmggdtDXLWRoe1Fl8TTexYm6/0lick/VZmrnzu7FozXAPUeJDajejz9Ohb1YD5h9
83Z7K3jPvmIbD8IiYsmcaRuFXqqfJCiM6pPttRRMSgvo6fibMli+8nd3r/8J9ePC
5rePo/tqJ952EePFFqtmzBog/UYBNn25b5PU6dKLtb1s549IHy2K7UtZt/um0kW6
l9n0Td8OPfSrNvbXU8Uymj+EvFBWnwpz2Gn7sXoZVEYqfEKGEwRKzqSaGSg9kY9B
DDyUMvTEXLQ1639sLX/XK3b8JSAEKfpLWRGNld1GeaS5ziGW/WfjIoOYlWPjt50E
rdEyI7OqZKXBwZ1yO0CbosUPTu3y2scbIahaNKX/7iMOYaz9X2FhfONkHqiqXx1p
EoKlMR/ip94UhkuMpPB+3QVzOiFFRnXGry6Wa8cOQX6QQXOfoi77xNIoLrBbluy8
vPDEKYaHErJ/IkJ23oYb4sjElXfyhWX9uJC9FNeZW0zct3srCUt69a8r+Nkkqj4w
FaZcxJGA6oDplAXS7wwE55NVV/3ngM5cvVRnFCdbihrwajRLGxUwF8XzI+sBo35+
b86FwTnNe+7NtDllmFpwX+kN5FRkQw7tu5ugdeYCLaHHjoa5BDTeq0huOWusp0+b
aV3qxVa2ErCBhMrTBsKCfye05a7tGo0NG4Sg7d/tFoPWdqHih8RUh5DlbCqQeaTx
4HxlnJd2dbcJA6sNCr5oLPMKjXqlLt33BnOiXqC+OfsXDgTo9RmNx+CFbirPZq9g
9cDHxmn7uiDpHNgBvJsxNMK7N5guZSTLKsMGONC59n0HPSGeE5JREijrTWUqBtLw
UkNJDPNBWZO1Yew7spStUYArKRB/I5D8pmWDUrKJr6VSrde/mJ+rQi7cxjtbPPS4
5nqTHuHOk65rZumuL/KUT7geP4cXLg/fWaLTFHqyNN0sA8X50ZCbkQxWiDjnZ6VA
VEn1ty09cguNTu7rVSCxYTqkRi4avw8LeFzC9JVtDMyz0FDq8WLraBz5JSe2m8wf
JzgnWTfdA+VXS6PDqKUjok3aRp8gtrOE5/QwLOI6kkgr3htK3w8IvGpyNJGxzjbd
fo2OX+ZmBImpmfqcGFs8Ruy+FqpKn5eyvf4/tML4pr19IvokdbpYFho6jO3hGRWy
A4TskTKOn6JvCA1jW/Fspm2S0hjSEzR+DLmJPLbOs1VURH761fr0hi/tlMavWW0o
HCUCWc39YODiPGk18KAd2EflG5ummOR9V0kLkEnFv4JouEKwB35zleLHWSn+B/xu
6k9jc4CVpk4wmJdsy2TNrjURU0dv/x1euWhIT00shn8Ye3scbwIfuoNC0nwAOb4E
Xd2RgpSXG6AVMLU2Q12/vo/DjVFCpQtWJQmHw+QeLBQgOi92eDYquE8wgKKoYGPL
J5ZbUqmwkl+dVvLkrydJgQYHdRDZRzY4l27u+X+RHAfe21G+9IzAV387vSjLkuAO
t9H+JX5Rk56zZRtyOZ/UBAvLtsdJRdIlm5PRYRmH3NXYhYCMy41caaaJQcpz32d+
V3nRBEyazXA/dR5vCnAFdDsQTuEEiOvXQEFXsq0gHmuKQRLWVFiUy4lzKmuBmnAL
Poh2MGpg9OwL6GHP7x1J1zS9F2P9p+z/iacsF4vnfHOoWQxdVRGOol8rpRvlMhF8
8cQAh861Y01sKN8oZTDfnb0twj1Q9ISl01z9I5y/32EEUoiS91PFr3vNbomBxtRg
OcUUp+RAsYsQrZYTknZhlIiRdhSJmLkn7/xnMTxR+F+EA4r6hpV7OcWGiXp77cwX
+5y3Bq3N0lmfQ+SRadGngvm8ysCstvy7YITirce5SHT09eW1bBmFIHmwp1XRHtIp
E4h2tasAwadnV4fE69ieeNGM7I9IxSp1d4i+S91S0Sns5Zty05C3uvss1ahR1Rjp
KI7ZJZjESIzS7y7s8Rwl4QufXifLodb/OZCo/6skfL2dloeT91qc6T+P2k+hF4UZ
qwNq8LBlYcTdu5tsrdKdEY/IKz7bAG+kJw0Nu5YfZxJkkQMk5+7d5FWP70+2ZkTW
0qatMlYmvSJ99qHmGpwydPPJHmnPZdgOy3Tk+7I90Wvc3YsUnRe9RtQ+7WfKZ5Vi
eeoPF7twedJh15yN5Rb7kXaof7iQhVcXDofOmqjGQl5K3TP1z4bUUcWg50AlJEyy
EPop2eaPVUM1xRY71TZwQ6vo24qugAC+O/MzZ0bHlia6BCOElXZgmHgTw8pLBy5g
suxXKNAC3FPbNa26GpCgrof5oH3ogrpF9ZjIfE3jJfRz/3NAkyLso+kpAXmfuTOy
hfaM2/lt20Th6YJ6ugrFimuaHnPPx2a1BFfVQqJnAJ3nFRPOEnl/BVdort5SiT/Z
Vd2OHiwTJoOe39wuhYQWIE8y0chq4Lv/kp91o2+B2cCLQ+tAqOsLM382J/lOYMZN
L9mkOMT+/H7zwABh3PRVYqvABZded7QF8MgJXyVZR/+U2q+u/DbR2u4G7n1ywo6a
Vj7Uy5PfajOcpMHFCiWCyGA+uDtiFDBLTyuY2wTgHi2vxyDWIzlAEwK6Eswljev7
d6pFJrw3qrwiRwUIWwYuCG2KrleEPTR+F4hF0ZsWvyvhrIF2bjkv70tnl/a+dfL0
dlR1NdUGDcKfQ9khT3p3Hv94paqCLzGGBxr4VX/iwtwoPyqCwvb8x/taAkc5ixDx
tkaK1th80l9yfg5ey6Yx9+MdkPW5mXGYP/eL0dgwClLEMxPYsl6/jdBEXAa9xvDi
NDTUk3xmw6VsyFrefcFytlTO8x9weVcmuTDX+fUBjuqXC8NaDzkFJ1q9gye/dFCY
8q11f14xDGxdWxJIms5LTm+658R10lcJmPGTkEbaAs5hXrH/YYQ453aThZ2WbB3X
UjYstwjBuC4Q8NZ6TgwSZawY1jZfjxvOZF78TMkWxzslLunD6WNcIYs/IkXaX3EY
WFOKGxhTXu6+dMserR2f142SNYmckaqmfO0rS/WW6228AQLHZI84MOVRQupuS6XP
OeH3M72yZFRZQAT3whvOvA0yyfogu2CJ0OAcG7kUosbaIwWRFQG2IvMkGxNrkZKw
qQon9Wr3jn+cFsZ9ThJw2Gu6Q0shfSO314pwHMdJUA/I+pQLdWtwx4KT8V7zkbXl
c7EmAlevM5CGGdz21Kz3etWmNrjiLEI2rrKxM2tUy/l9rFkpSzx52Jmt4NrmRKZf
n57UQcXHGOA6i+d0TZ6dmm6cyHs1QvlPyeR3rUXSv8OFXIM3RJk+bfhQY57VM1oB
uGW+VfAZbVoxaXQ/zCSi3lvGg3pAl8K3mmmpNyk9XK1pw13AB7vBCBpwltj45iJN
Vc09ZSI2BtgAb/Z7WFLxmpiFRbaMEotoABfhMI16OYO33o+npObkzyzaXufk0Cxe
DkpxJQaEN5OeTcichiygUBgi2QMe5nhkm0pHmH59Qn/51kWXxYl4EB+YZoeGM3m4
gqZE2fYGroyGfWelR7A02EnNtQFhDVHVOWlGFZkSx/35bb2qVCoWA6UCZ0iwq8Ig
kWybTJI33vfrwUJ4RGTzVoro9mSrLUdM7eKv/7DuorNVXWjlJdZtEN+zKrNq4beR
qaxw4v+scYH0CG9mjqdGKmQQG+rBtaeaj8jaOBant1LEaAVP9PQWbIBt8ReHjOYA
aan2agokGDlsYEgX6YxuuSzvlbXMuDIYKEdSM/CrvjguIHbcepR1CY5kAB9H5MFm
MxAEllSctFhxoHAd/pmDTgPXvFS4nyuX3zsiGrTClsdugThzypBmejyu04WSjmit
bhEW1/eTq/V0jyhYts68mOJZR4jKEwBTjhNT59emIIjHTQazAE1VCI2DVoRX8hd7
DuKm4dUAlReFaaYsOCi56ZWhjPJQw/4XgYs0JpISnY6arS+A+hx1q/jF7iJd5G5s
Ik1c5u1e7PEMy246vuuKoPVwRblEj/6pqrgwd9UR/Slc/TeXEGtIql+NWYbUHbti
KiWZ2KwXh6Fp7HOZmRSAb8Z7bL0ZJjqMi/2SoWgUFE5PZqn/MYG3ECWmQZ32T7Da
TMCxyxgq58mE9XbPXOiJG+ozHhviyOKxeqNf+N/1wCkNCin5uHrkWggOuDARQYxc
LuhGGpUcUUwp+lGIsDg7Hn8pcKa75u2DOz1XkIxB8bC/GQYu8N+c9t4TiAN6PsaW
+VocuwY1Wfra8FQUMtomP+vsm3oG2WISMqzP4TcbiqPlmrFpEvpmWnqEsv4AGcjX
skPyXlklLZ02L5VN7vB8q7SCT0VI4RL28Mqi9YXwOL40v+sNiA0g958YdG0/Mwke
qWsYrAoWacKbX/sYROzXve0t8QIjm1U+WfO5WuEo4uLQYmzPu7zacubfBMwkwW4S
7//8eX1cZ2vfq/99jx5LnDDnXTr5jGpAL5dq7INpfOoSk4ZtEaIHf4s05TTrspo3
pDabugfNj8nmEeBKI8DkyXSE7lkeFSJr4+kOAc08QRUfXxN4uYfSrURq7Yq/lL6H
RR+RB3Hc60apRsgAhK9UXzpr+I+mgLf/WdgJj5/JVkx4nal2LICL9pb3dEL0BjSh
bhbeQXbFAG9Id0L7YzXRc+x1vz85Yv7nk0dcR5F1ZTIWzA5zNPNaA1M/7r3pagbu
XrwxnxXL2RVqpW4zKDOxN6qfc6kc26NERhH0u7ehWmELThKX4N9h9joZb8QwqNnt
38WgFCyXQ+u1jydwuWNHHXKqJ6FGIINRP9R6zRF/gHjcdxbjnVHNHOBmro9ZJmBB
hwOH9sbU5zWslsFCy8nm/FnIghxCSnET2dhhsk6p0/S7BzU4uplQ38HRe7qoTB7H
Yydt0wUp+tiYQOmkPnSFnlesiEM+VH+gp5YvDSsio7u7HPaoW9yEM/NyWweAYz9d
SDYdTvyHgOothmyy34AfR4FqHgg2CxwmTUNWleJOzziVNC+5i7grWn4abExqjF56
OD+Gu2ZzJvEq6wBJ/bzgarsjkzUC4IZpvbBkNtK4nW6aJ6ebPcNbVgmdMmH4cAob
AGdBDTFT6Mn+CnzJpWBDflIkclqiGupkSJIipjrAWF1wU7vBH4GcXI6u0MGKozRW
SvfFrdvjud5IE+lFbgO7xwIWzVT2Zs0JMBKDiqmpKnLEKyrTV14mvwRrF7o1XOA6
W0ULAgSgiaREAsv//A6a4RIayDg5Qg9ynhfbDyNp52OPtBBOd1+jYR1qWGs4z3+6
rfEYsEt1rxFr38JQOil3BwGPliv2sxpVPoWE5ifEU79dvv8uR4wL9L/fKErzTd3S
Il88OXmUKl9uDf4ZjbV8sjI04xOEX1pgVSAKzX4eVtBgBnNGEtXUmTvrpuDdAcO4
FZI937oKA1ANfz40rEDQRlvXB61AHjDRQYFneRrfJqh5C+t8B7e0vb211t998i7a
BBNWJSQeI5BHCG5PZx6aG1ewT2aosUUBsDCIjDOIeijufhdyAEl9jY9NCCRLCp+F
t2jb3/V5vVzTbZ179gpsExbyE1ny0AOjX4nc0iiUhaORoKivKf7PoM2PM0HOYfGw
0sHk+VRy8ohvWL/ZDetJG2R9BmGyxgsv5jR77T1qP2OiurVkcB7iQ9pcTN/DyNZV
K5wrsLfRDAhi6fgwTaV/fbJqDkxGI/C/ZvC3a3TUyVXLtfnoeIIk6OxbF+X+zKyX
tNAsMCam2aWKoNL7U0BVvkazsTaL1B4q4EzLtBX4IYEMdEs8EDvo1tmWbUqM6o0G
ZMWKz57FVy5UGG5xA/UGylv5G4+MvJD++xa7LmhPWF8hhbRpN7dmj8QzPRvcODm5
dBIXc49RKzEFrr5WgV31ND50sYAgvHo7+bz8ls7FKP+TqetW9TL+OxDcuauVQXgC
T4AtTfgXGMkTpSaeN1lGGlnqdBXEIl2P5l0K/giJPWdlx4eSke1Hm1KNHRCXU1x5
ieBWHBtRZI2I37HccZF4XBtD/XS7dWWkzQWNk1k7S+KbWGMEgotUCe05v5YuzwRU
qnP4hBpcwmCyYYyXLv9zsQQa96TFTYI6Jk/Y+XbBEVUMfF8Wc3B34NWMicK+1MSP
Ek/lMondkxjlbRxUHxfIdtZfOn5tzIsqaQnikFDnxy+Q975wibW3Hhc8UPaymOCk
kq9lUKwOF7pq+Gst1PO4D203CkUXHz6rNfbzHA3iW0ph0zFgMGqR8Vp6b41Y9nO/
HInqUctg6ov1SlpoXhq6QGxbJ4JhpgLO8uCejOyxX+9d0/OqPDKZ9I7fKSdeUuwg
7Dftt3NSYNI/MjN3bld+qDs7cVHO6/ngXzaHMvmypsEl64YbRoHZgtdGD6L5N/lZ
ZrsBUlF+ify20Q4wg7+iKcdlcXhFYQwu6OrLu5RWyMKO6Y3K0yeK7dE5wR4RT4Xs
MvHOT3rsLcGVc8IkesLU/meuplRK6P8MRkIYefSudsv2CAyybnp962dMHe9870DF
F35N6uthcTzTDuXKpa13I/dudajLvFvJIWIXEtd+xlnTWqRcaWGYMX0NTj5BJSLb
rrsNsmOT7zC32ir/h8Yb0IRUATbEwua6j+Z+btPYxl1+YM8grjC/gc/2tyTSkO9U
XwAOHNBwtiDLnEcT3gxSpDrfkx/cO1nCIuqB5B1kKbHXKuj+3pFE7LhgY/j1TEkK
wRwp1gJZfDKJfh+ufEfQaItUmQL8gV3Y5piRCXBMQU8eF4HddF27iZv9DpvPH4N5
nG2FNU8S52GYe6PqmMT3YOoLUMXGVWhn7Lo9LJqpErhYu4LeN+2Ik/+kQTkz0Mgj
xJqC0Cg0pfRivXtQC7nu5np6MSJxcnmjAlN2hyo4olsYtihT9YIgOT2ZTrLiwHuZ
Q6DkXyZBNfK8GAlNv/Smt0ICPnqPyxdz6t4JYqtINScvErlaNo+nefdPKzjU3egt
bdzAU10tL0/owy1F0KjgA/5HN0RiTEXktdVkHOoQrQg9v+wo5Me559spVFl6BpDI
/rkKrI10jZMOQeqrGl2EorWvm4UHhktJCNpsVuKEsLb1wfiPcOpyHIKicElYC+Ix
9LvwV6HMV3kdVjSkd7PAvFgo1fzHq+fGRZl70L8S+fFqmPTEzCD50XKorzb3xtNL
Z80AY6qL25/6pyzwHV7CFhzGPUkct2DnYqCFNUUinvDztI8krpArVS6XtmSHQOBe
3ph2uHdK1I40841T2G5CShjplesnnMJGUBPcSsG98O4qfJoNs5zuC0qzRFVBLiP/
EnzWG2szN03ew+Q1XDaWinXpJdJP9qP2jZSrrCeBngwbg14lp2XrJSP3xXX+zhbE
jaiu3nkABd/6ypNwy4XMw+9R54gh8VENbpQAeQf7zQAESksAU/Unn/6PC8Girk1C
e/oXIHucAeJo/em9QhuvlfSRe2C2p1QAMiRkABylkn5jvuJV5Wlmqvuj+DGzpBhy
nf2yXCJwqtQNCOz6HEgS1LIcFZHdZ50uLyheRNVa85+VE8Lq4rflF+tburniqOee
xsiGrwUoYF0vC1Ga1ZkL/oc9iech6P60BdIt4d+ss67MHoGLXPmDy/xIgSGykYP7
6mP9RaLkWb16jKGXSb1iA6fyWPYiQ/M123w8UqnpjXVjrUaULPu1IJenTVtMVLoq
+tkWYqynJwruw5a8XdOfAFPd4pUK8WEkYaUXAt3UWg3cf1VN7E35uIPT7m2dJOHJ
WfxR9U7vdjKVUgaKLvl1qApEAYxHoxXKqnrt6w6pZ82NRa45rz44i6Bu1+i+BYMY
me0LsNFB+Zi8rv1lICOKVoqgc8BUxBi0wKTM8t9EIHnoaA+lSeG4hpuFrQAtSzcO
DXg2mIGS0pOv/SXv3NYbffvD8oEHzw+AubTWVMRLhXgd7qgDMF+6YWPjTlKu0fcD
hMqAs7ayfmpnKZFmCpQWGAiilMffKYK2INZ7fZoUHj6gAhZS9rbIr6balDHzyz2C
hy6cq8vzzLGDbFFStEHzAXPqROGnyqkyg6IrsqzvS3Nro+EU61b6ilkf4HsBuETQ
SByXcvsiymwfY12SwLxhCoDD0xmLu9ERvG8gIo6SCS0RTFKgI740hF8THf/5WAVv
IJiF/olXRs3OXp2m1s1zxbcS7eAG4ysi46oTsk8GIz/lXtv/9BEirS8A8hfE4++U
DmkfeNZJwDSAeJPxSXFu1fmf3vFdWyeHl8hFc5Bu8uvyIuT0IDYhKkDtQ7LtqzeX
XsOpaa3l46eGYuVRNkRYeiFqcWkaHQrlIJympewYBHs0F/UwBEy8EKvmCeKalOIw
PAOeT8vw3rJ7+qjw1TRHf34tvAN2JDZYhz2wwbIhqIviPBdlw3ljn0kRidE7yt8p
Cpzh3cAHdpMBHAmOyF9grfsBcnN4KjosIsVgv1hbMFdOJea1Iia+/cdZ32sanx0o
a7vsdFeyz49K3gdd1MJuuN1UjMHcPVeki6N7EuC919Aiu/+KzWVwggyW5UM9GDiQ
XUIxzfxjO/LpOgtpcWpQvpAfJiomQrG+3DgHtbIOLNLv6CdvJtvd9rEEt760/lGn
7Nl6k/swg5Pv21g3WEtq+VuZIGviPTEmdGyeDomXuqaZF72l95Xdq/id699Yyv7X
qgt3AVv4pw/XrjHYgYy4Y45gEizJ74IDwBj+0wBBaCvRXx78ro3JSCLH4ZRhRx8m
IQIpXjETpIiVWwiqCjXIoC+I6zBgtZPD59SmRLTL3hmN6ZQWPiAGrY4N4XlrEpmI
TK1inVCsFJNN9tGWwjl4L6iDAutFcE6n10WyEeeGJESLfZADlGN/fHH1WLp77YRp
MDBSrXkis95VX6PKMtxiCyLoIxXz4z7eajIeKpPMPpYR0J4oJg2cV5Tfk809t5z6
P9pzKq8R95QVuORlf0UPZCqBQfpAkRHuW76W9AY/8nMz8kBJ5sqiwEgePsm/4EHz
HzKDuKAFobruvP77S/lmbWJqnj5FikzGYEMNHr4eHW4u6EypWsvBHlXLo7+BoKzv
mqkAEUaix/q9Xyu3YNwSSKx3qgyX5od0ju9KaXd2e8Ctc7HPpR6Fmjm4wVGtmDiU
RkcTHRbdhWm7EB0GVHatA3Sy9fFL+YG+aant8kdjR5V5Iqh8k0cshwVxU7GqFXUV
QrrBU8OsBFAl7LM/0qJYSLGKGNIcBw9wnZTwfldWrpI1laZuqYNaYIC6cLTeCKVD
Z1Gf5PFVH45MzzFup0LeaAtJmd8T9935ZP8aOktr09Qzc3k3kaTVKB/WGKxg8IX2
XAxN84RUBPkNIp7utRIp5X+rMHYhiF/rM+bObqH909pW8ZRHAVLz55nc1tib2Lgv
FONlxBxrdPVfkH7jBFo5Qalt4432EZC5wLvbXShIh8e6STe5PwwflKIk4OcPgtH3
8GEBKGbxSS+GuUE32AwVn4GN1SmNaRwGpHVJkm/IGGpMoe2nousjAkqXzNFr9RK9
5FpaCuTtCXJfbkxw5P/je6J2M/SMw2vGa2UAO8zr4Y0Vaj+l5vifNOh+SuU5r76Q
Qa4crKqPnmZq4ajetJX3bk4tsY+gaZblDNHw4Lmyap6wWXXIQEVa7W4L2tqb5az+
Ho9r/0+1Rmk9LFrEzIM+efvDcYix9pE2RtPmcIEEkDKmCGgZXgRoDP6xm62HhC6M
xOGa37o57eY4E4UbfHFGGJQsMM2tUPeMO256Rb0LPx8tcVno8J/fcgAq1pNC7Rq5
S9HlGd2nJ2qL3UCdZrPqKugHD2yDws3iFGxVM3BAo4mtYAin2Ff3M/L0wPNsHyed
GRuH+oaAtgFLY/iHDm9PgjENeGRZaTfHqTYCpTeU2a91L2yqVnJ+ttEVWPipfrSi
LRV2YQr4zV5qOHpLNrk9sHIVVrKG012Dah2DVovBeL6ZtmqBASaByQyU5gFMxOAM
DP0FSoau9XzFDX4pziifeRBcds+QMZjkP3aJ2S5Trx9KDw3nRJeQc+Gx9Lw7EMn+
JporI8Pv/DgOhFs+4NsLh5m5ylx6WICt6+5GDQL9DteZZCgE1/a9t+O5U0x3Bmkh
3wgjwXFihDJTGa1B03k7zJ9yVXesJa+8Lqdkf4aFXclDVH+2/zuQI5hfD6+3UPRf
yFAVIOcwKlM9rbdaEZXQSvXTAEJI9+lmZOkFsi06GEhghDjyAX/0hrL3C0A7jxia
3xzbodknFOjKQUrwZ1lQUQwPMMfPiVAZNg4z3FioGkU2nrneQ326p/VIGAR9g6+a
F8FDWt/0gsWzzQU+28OxphMjlmUSkjGzu5Fp6zmpr8Tyx54SOaLkpJC7mkRbFTY3
H0DE86kjcndKTWbr22b7+KVc4CIdK9pq7ewTH6vW2C2IYuBxpvo8uhZSLR6XfOFx
DZeoLiaZoOy4hjaLeL1ly6oxCWAaI6BzbaOArivIva0J+ida0TfEfCMK2CLxq015
oc7g93WoiY1dia9srB1Y4Z4MHnwja70uAbYycjEbBfqD+6aVuxZXjuU7s+VEGZ+X
H73Yo9MAyzVfLPmMCaxFQNjVneJc/x8SZJFrN9Qw/su1u5gXUTOvoFIHq6fVjusR
UOTKknyQ7mv4XXSa3nAlBcLcyZMfR4FtyceLXKDKrdKdIwQMGJz3QwuUqg0hWLeH
yxxovM117bAqiMYUP2zpIs/SRagzYyKht/RClaQ+yYyyO76QGBFzeG21SwhTUefw
e5eqjXb9db92sRJAqbKIuD70n2jg5j9AOoKmbgDRZKlaXmbE7smgN8G3uyxakcy8
Mk33P27sAMxK6GKk48PuDCBb9XGQB7FL+NK36S+G/9+1t/+esVFuSTnPj34Yttm3
U71GjAZY+wo0TBILZWwQ4ad1V3aGtvpTquh5L0dWkUvV4qCLxyrLzw75MTcUcHzl
sU6F4OuoO71wWgU4KDgB5xJ4sJvtYTP58HwKkslH9g5fV/SNqUV5PvezJyQbGm4v
pZnJHFvltbuX2sFz9VByXsADNCL46zM8plsRkz7RFI6PQWWOtCRShpc17C8Daad2
glrHLXwu6240CYGDN5XpRcOWh4SKE2VhxaT3eHFLSs98hQG0L72FDu2aCOmn1nX1
SimoRuTXbjOZ2C8SR0dLMoCluq0onRi8qmRdw3jaaSSms2648KGxKfvNBnX6yMR4
3b/sK0Slvm3PLt2gD79R0F7No54gS/ocJ0wd/u358LyvfTnrG8NA6WsOJlDLzS22
xYgKN4VsGlUnwCnw6J9LabPB96OE5ocDhZfl+IRXNrtOWs8UTiTs3kWit7tc+XSL
vfS7X/ClEMWLPOzufDV3Wnu96OTy1JfR+eHQeKz0DFm2wrK0ZRkihn0uegB4OEEr
cA/ZUEd7epsVZvx1ZEfk4uFatvUd7dL4KZDJZScT8yvNmW0tihabCpu6eDR/MlZp
YXSBa1iSxqjufcO59lVj9tbTNhJKFTwaUXNTRdz7hxrI198VPntfIfmqtYz4vagI
6/gYvZXvw3RoHvbCYb0N+/jBQeL89fmB9oh5Mz/rOI05kgTVEmeM6KqfMqrSErE1
ygNHw4zvuA/78QoyKSy1nK2WNaR3f45tM43Sxo9X3HP8GX1DT+XvYjvQ0w5M5Rmo
0FGIq3X/Jncbx7t9bd5kbAEqYkgcM5ARnzYbA58VmERHdv6Ym3F/9FLKvri9gVvz
6ALdPCzLgOz3YFIr2qSaSE3Byes+wwfhkielAqQKyUuSuyVSwCMzJmf0QOvS9gLS
gWMHR/Eccnz2+Trz/xCgl/UDCzQ/GtPj7SxDI95/d4CrKXLGYWEx+ohISQlOYG4y
jKoCkG3FcZoV8Z5uHy3LhNCmTFpnGxYuLXj+R8xRTcTHaTpmtNnOTroRqaYz1iT+
uvhmPcSmve2z0JbUcfeD3XJNEL4PN45qk4VKjSyCN2saH8xLNG+zPKZxKAzD7t/u
bxrLYPS4tPtqBsGkGyHneOBxk5fJD26RBII8qn8OXU8jt2V4eo2+lFHqD8f8GBS1
mWXpTY/YWN+CQhDXVL2veFFD+Ly/i1v0KKw83UPIeHmb6H9LFPKt5NN8tWqzXMjY
3ENOIYX43fZ5pS1wm09/1ZojVhbZZB/5wUfTrMp9W5zROiwyTuvnwmLsUpVAp6C3
bFkSIhfasWfHXITrC/Q53c8DGg79fGAHzeYjHJBXFkhekFjX4q3TjY2Aui7KetV9
0ET+oTZogxxND3s/ZPP4Vo5xQ4jlNJrf9Fh4AunSASq9Gi01oe+aojLl8jy0j4PL
0cSJBJsUtPhYwKoo0JRzsjdJk5ed6K9f7LmC7D9HRpKZVXVnXi7z3jHbMv466PNy
AOavBw2sxNSNE0DkbrxXjYZyFJJmAV/VIOflrhTsxMN7wGQiBwUEJI88SbOQlIHs
bo/Cb2NpkFAvWMMUX3GJ9bApn/yeY54+N/h4ly4wZ2VuKUhRmzISftzwtX2C4ieG
/vyxkiDAha7F47Ve7nYo/GVNZalUsQF8JHXYpKUNnm246BTn1Y3rgsKKk5ZJbJ53
iFTwZGGtG1FpmbefXXIBh5Ao+9ZbRt6F73CvX2CuzwULKq5j5tciIxcexJalMLO6
0Ev3MoRSUrnVUqCZp3RgU6PDVGGZhy9OimQJMRZkI0XvedfYiI6ZQvYCKgVcs8oA
ORQuWzyxihCimwbwAwsgg5+Yj+5vZJepiP48o/c8OwSIn7OY6WKHhWzv83Bf/ovC
5QgfwYJ2i4OS5Xo4LKP/T0usy6ARul9klMQcjDoZidSqPtl0W8coGOmdMxPtEzTi
meN+f0cRSCG/oKyP8mEYxoA/ldI2SMbynhahKhxhNPp4TB3qlhypH8MbWvrgIejS
sX8SoGxlZEl7xyW2sXdJSB8E7aBTFsU2IIbPMiFJP9EBAZLoUSRKgWoLHBE1qT8i
s+QeVtH433lzlvGrrmt8SE9OtK8trMRYws+tH9WhQXrlTxh9mSA12do6MmeQxRSf
GmRib6Bdpjdxcbnqwx328XdNji3h0NNONldZ1WvTJaN/xEQame/7CWrsL1XbN/pX
6wH/lGbl8d7XUHGRbKEItsOAi3RqEy5gIB3zUpajtydKDmm3APkx47P4UE9mm/9V
xG5SE3nCwD7mYFHxKk8NS1KU75aXG/+heMWsjIF05X9HxlZAJmH4TcTj5xg+CUI+
5m60bRKZ2szBNZXTVWL9NKv+0FhZ9No+D6I7UfWQS/Vgq1O4BoPCXXRXrli6A+Jg
IUip7zDjsHE4RG27D6OFx3+Bs03mF9+eAjMw+dTdQj5GI0nZoUbBxyqQOMVlqdy1
L5XUk9PZOUCtYNEl3Hk0B5/AHXohQC0wj+NKpUCqc4yoDkAzSiQo56JAR4pEf9fi
DTKDCXcMmED4TAtsr1cOwL+KUju3gg9DX6d8wxLWgWuaqLb1TNfYP1M4Pas5HDSv
zXuH4wk6UzK1aHjdgwksQXmyoZSV2CPBTY5LYO8yed3loppMxM3AyGmLQgMLWE6G
gQDRiO5Nm19hbyzz2n9cKm00Jc0T07eoS1xLj4Hf5iVCGHQXlGnTXZYdI7WoicUL
HPYCdOne+dl/IeFgdP6dO3gouXVvSlOqn9cwoZ66yES6qCnj9f/N1Vl5XzlfRNVp
BLes/iG/gVF18QhWFNSC4TrSF8VnUWgqbCF73JJHpzk7ayYlCTL14n4E1VM3yvFY
omoo5ShcEc7mzeDboKcLBcFUo/SWdVRwhSbfn/RxfSEwVmo+5vWCBO+5LGUexhRE
A+dcPTlmMPuv1HjLlkPHfUWc9jd/mbyBxEZ+VDBkmNXjN7uWMo7NAxguQsjTBump
PITVgLu0reoTJA0FqABjj2DGVDMy519JzuFJXVH7TLrUGd+nhiZCpHzi2nwpze1X
WBBUlTTtHne/YO6vbSJ9aRdYCW4gFs91Qod6d2qlurWsm7GgjoA0+hNJBLSP7c2t
bFasoVZgA1XYxUdceEviD42/zY9Ri1TL412aHEFK1oP9wj77IG78UZjAIUIFZN3K
bdKwMFvr7pf7IljinHJ9K8bsvv+2M6xnvkKI0L2GsdZabKf8HITlczRn2eryaOgj
RrUrfEfgTCOe6fu6Irnb1P+Gil7TnVPCCO+QelOt+V6m55olhQmezdWK0ao526EE
dHSmEM6GcoY+9V7ylLF+olJNwMKt+nb04qWDRsPziKKorfVi11JPhhHkdyFv4gGA
r5ai5SU6N7LqTLhndq56mXjmoFtpbz//hfVBkSrw3uVNOS4Jl6CLhQ23lE6jjK2n
WXo/HsIvT5sJqyK1kA6BQIgTGtUyHgDZCxgT+2cSEO9VO3mmdBGG/9rUdbrGyURB
WldTHENJDeYIH4ewjmtjHYlZ3iBocAcZh6bocbRc72Zf3+mOxArlbxRiGgj9oDpE
fgeEI74SJhEhJMgYblldFpJyJfamsolQIMHBzaEHfZFZh732c/+0xgVPmMnHx09O
TT7/Jk9I7YwAFAnp0MnN8e5YfZM0HTj6x//wD9YnZnQ1IV8vOUyw2HW3UzsMO5Do
lSz6LdyrGgx1p0ft/0p6cihWV8ZrpSGBZ1vj1BRMdHFCM11dfrY7wuycIaYRnedy
W9/cd62OPX0Rvn5ZvauQxS0C12QRLMF/jPTp33TvbprI27N8KwJrvknV4LfM+cc9
qCjSbtzhIx/neVxpOvbdXiwhFpElDyWjDJ2JtqVlz458qQ99B+tDRJhdhzeCVvrY
nfhOf2jL9wxkGBcdjHNBTCMOZeAZMv6sn+GvXPoaPz+30y3gsim7vQIpyu7jlZmb
pT/G20C8NWVgsBSdZtFfLfW6Ns2qY1qadpmny8RdKjyzgSMGntmW7BAJtHhntcBs
NZtzBEpHS+sU++Li1hYNVigSnIq12/LWgTJZaI8Z/nXNNm4u68e7tT50CrU1KJZt
LrZjkVG7PGWneyAeSj1SXtVMTxcP4LXdDStItCwt2WWQgLchYHuiL/5PJpylMcmy
Db4NkzjoISt44TMPxLxYBphG7NHde4A9/L3xlM5w+jvq06EXOtKIQ12j+EQlNIqW
gNit1DlX87Km8V1bpPmI9udrvmSF56Uuk+YHm1GT6jTVbzmcx9pfMhrepD11uUQ4
0bd/xc3vkWE1W8gtSwAV0c6bl+Go8gACyO4kelhW4KdBL4qDdjqPZ/RKRpGtGOT/
NqMrziExVpMVUMRFbk9gOMimuDPdLrxXRG3927FVAZOu6+pZn8cXe+dncBZzS//D
eP8t6hMS5fkFh8f3X2yRpTQ8blBWBbDiPevEjF6+S4QF56esCMlcPG/061u8U6/p
gekQhiJGIl35Y2kQqPJUyuMK6SXEL29yryMj81w8pfQSEwVzFLUSZQQ8kpZGl6St
DTioRn3IXuGOvd1IX+pIRjJXd8OfcVDKqOmQoM7qpJvpr6cq8nQb68nsbqJ7EcoR
mXwCu6mxLerEvNXWPm9HW7RDDW1D7S3xRTTIme48z9g6KtfdSQqb5MO0DSghEhrS
w17QWZ5L9IEABaJjL9jrxeqmjpXZapynBagIVIEv3OyV+fUs+6BNeTKEnP3itMJm
OyRZD7KPNW6R0AAr8K4LQOE22Urxc+h56vr15pwrsYwGkqkfOMqilj594K2V5e4r
o32mJldzgP/jknMTNLn9gZda6eKzTYfmNcmgzFd639V38APXDVfs6QlbwQYq9Pf/
4ACROvlIJvK/0PCVzBESo4PsGMOHes/Wo4AdoL16Uy99BmbNUOxTUUi6V70aBxeu
cFQjtsEazpmtxPD4mAJLqq7nQlagcvRDn3r4G/l53w+f4XCq9xJC8PhmhMr9JlbV
J5wlT/dqTdT3UexSjOlh1Vphqc3ujvKCv/+SOBFjSj50BsXJYsZY+IFmsFYXNPqz
H0XnGAUc6iewtsL1z1H4Xfu/BqNtb8sWtMHUsDbCyGIvS8jtoyzXxs3XPJlGI06r
D7d/5ZvoF6SyA5ykEL+LpUUF8/9KIzEgXzcFt2YsAaTWYJfZJ0p44cImCW0aDww3
bU5yzJOE0A4P8nfX1jWBr5xnP4b8+ZMH2rMpwo4mz2lCuUQDZeyk8edkc1UV5Fyn
ibzEvYMRPbVtO8Vd8uhjZ1yM+T1URRnNiwsEzGOIhmVSr0qCj7IOS4R9rG72dqwk
GKJGP432HKCT6IQOq/yHxlXO+lmRwUaEI7OPz5tza1d5ckuIMvuGjIdoJWJe2fhz
KqSz6OQfR50LYEOBUZwzvblqvww3DwM+19/ZDV11PcnekzzlPXUzrGHZwwAOGlg7
Lw9cnW6leg+XpsMhqEOBGSWg0rZ6wS8AW4Rfu/Z+70aBkVjV5rZPdeh3OKruSJWY
S7vo3nyelfQnsMTDCUxfz34EXNrv6I8QPEg4Hgq/Xs1IUNdQyv8DP2koEElIjDmu
ARROp3MjkOyjvlg562DX+pV9mHUPX/dwqnNfM6uShYXSieVpSSEWWiLzxZ4esDEp
gN3J7WphfqDahMairq04lrFQcG57edHyC3NTjF+NYLI5h2T0tmvG3bgyaJHTeRxS
CI8NpElMQBLHqfufs9jZcYvjFNbhgp3oyU+qQjrqChU9/GyEaimZF5FAomK8lLUE
lcqh72ZRYZmjW9VpX5jZG2rB8WCUsRInOPXfRaXV812GyMbc5MIMBUuLS7PVxoUg
k5/skPgbekVChzI9UjPhjAwRa4dm+7PGUfso2JVYpduUYrSyKDsxstHSrm8UTf2m
edCT8eT22IEi7JucBqbHppDjiVt+OQc9a35t1ZQd7VlOzgEcOamiJTpZZ1lDUo5C
DYzgKkEevpyo9ioG6NXeWtE9ZX/N7wLccb+XNdo1pfCXX3f9WvIsJdQnqiX6a1B8
oLsjh+F9BBRiFJqfudRr38ESJIP1fS9ImLkZxg/aj8mB9j66+8omEhPCMPHAK6DL
wi2lWntH8azUbHZfo9OXZtdErw0PCQ1OS1XB8257g0NqQOsZu++K8EpwL7UJhKwK
/s/KSJMYmyUBUNdF5xv3Wemmc0c36j85CCte7D8tTAf3w1PawOCCwAWvbYVsTGdi
Vioy/7SEff+lMmw9OKYUmnWYImzTNvxAfDSuctYYTp8hyLb9G+H4F+VLSZplJuhq
79quP/lzJUpuO8XOrDbboVMPojajPoc6B4qWhjiMpOFZ0V0n7Gn1q/4Iu1o+vZ4b
YkYAyE3rgYJdlz5aDIevzAanGSeQDEBly0rsEXmn7+3BIGw2QQuonMaN8TQ6DZlH
vkJEt/BPlDirmgp0RPUPyoBgPtKJ1HNYlclPOqvv7hS+lMJjcxn6TBFaTiNzbRiR
xuzhAWT2Q9U1tHJj/uuX7JKow9qvL5Ot3noj5AzYzr8nXrV0li1mfu4ANxjkQt8A
CcoASZvvyHfqdJa70y1KDd1ue7boECA1TE/BGNIRW1cc0D7UktXPLDKk1a7tApMq
9HvnU13NY8QGAlYOz5zg4G55goIPrJGT/6V/lbFeiBCa4oOUf88GfwoJNAf4hgwM
BcoSS5xsAQcgjTP5UVB3AJ3a+uj/1u+ZxpLiuXMHdk1JTM4LVPGVHBLeHKGfA4+n
B2tfnBLOZ1PA8iAexeizryvQIL7EmMJqsYAB7bvo+/mgWgZiUQhyH5Cb232Rgi2D
pBLTh1GMX+tiirgLt0P93JqoKkIdiZTO4HdL0N+7rFRy03pN3zwVXEcTKgjSm4D+
QrMSHyE7pCPPBBOK0TpVTjZz/e8blz6ekauvIUOX3XzhhN9+Jn+OynZpqLIuArYy
0WRpZz9rADLDyuUjpZJjMKb2QtTcGMWuRL0QkxRAyknlaJQwFOQ/OtMcHS/7EvOp
8/rkZuvlc9WBhzmugChjEyNpx3Xx4ysjYAWZvqENHlpg+Ixw/pEwuDm2CRsvJqZE
VnRHQlHKRj05KDREaaDLWWb/l8Of5O+Xj5OCmp6FxWeGTywboYisz7tZjoid9v9G
CTgy7ihf/NIEulhK1YIIk4DlkCkZy5SHgodX0LjmNRhlaTkngMwN13QgD+td2b4c
6drsVddf1CEq8hsEd96iZ2ABkhHMxtLbtRflBv2zD4lLa7BFwkvmJUTXwRksVUvU
iKwDzwoAf53M7F4BHNMtaho3DfqWpJn8Y3Dxb115xI05i+DXqiKM48F91k+6zQJD
vhgQ7rWwYMP7Visxlv9HoKHbaH9D3e4ufJ717SbtgY4LzaaYddvQuCaB7Q2bOsan
HpGPJXiPLg4xjjoVZRaw/IEAmYFAbm27qQni/vpDFgsPiVGNSfQXzy3O4HklYFC1
FxZmx1MOiQ0GxnLSqT0PvuFIejFejcuRzpAlNAoNeJ8GHf9Wg73kOs36c8hAwYOi
0W7HD3Jqlt4D8gGmVOP58EdOROeksffqC/vYBJ08hfm1oEhJSETYHpyxZX4c+xBS
SJXSmcEpjC8riTdJnn8/U5IotPQdne0jIzE5VWQWqE5STDKytrUny4ip06P913li
p1pZ+vAXmb9v7oFKHMd31NLNNT0rSlnCgNGNi6FIpN622mrfVsnGJzCzttRLvMm0
aizmqNvkK95QEqr9fHY3ipu1/9oFHBYh+iczd9LHns4PxYTEolz36SLlRPS8pUKr
XWfxnLjexf0VGL9dkofsrvKShHk8DdCrLU8lPzIOWBIQYA4Z/c5akJF/BcWkdBnj
DSMtGM3u9UpWI7zmF8MK3FIF0DXmUFLc73MlSMzdySlUIuEsXJvMCXOdyMUFBqsP
DuLTrAguda1TaeXygYpDqAXCrst+n2JRfXK6V0mMSliCkxQ3PS69kuZm7eKI0pez
h/mZEnPr5Rvra/Q34H4RWZ7ipkJziaQJaan4RBrFkHIKWkXb74KQtpNqngD5NNt+
BjLwepqtMxjP/Rj9BL3SpgUC7+yX1mfrmXzOdwAP5+WLWZejIwdC+pwBgwT9YyR6
ykI7DhSBUKj1gTAY7c1uGzHC0ALky5J92Iu8D2ZKkrTa+v67u1DSgwDIMmbPuwcc
yuNccF+Ob9cm934KooF55c3GNDotJAa+g/7pN5OMPvnY0sU3JHtHkbBSBKeGXcLd
heIojRiGI5DtvtKdfnKCwWVSV9tCmUZuPpDu3ALcwDzjpCFjg7/RqFiQcdKPcsjm
zxkigq8SPNyu0fFKE+T2Tk25geyjMXqlwSPIu04fbetQDZEPlaEidRvYN4o+R6fI
UBj5PCu5HzzJrCCvnug+y1oqQzJnR+BnuWem4oKiSndxwSAshQpgFmTpRDztbir/
LOLrpI2fyUA4hWdN5afizbBOn99dF00hI1NHumU7TNL300xsk6w3shuYaO1nwvJ8
0lqMAb35oL+nriwYVLO29qA5fUvksJLJvNSedwbvR+PMYvLEgV1aZkPTx1iZBU8Y
EldEOURT7sukqtuHVughSHn3h2/B2pxk3yUBjndze/l4FUT/r/F1ukB/zDYo6g/9
XcVgZ2p5thvuqzABDeO5ZNQEwgYP+FnP/ixBv6xkHvkBtBbw1M56pSN0c+FcE7Lh
yCNAILxuff3HLVP7/5jux6GzAYNmF+xke2PGpCpVMujSlQoyU5IBhWLdTdowWDGF
8cNnnI68lT1kUFE5eKvHcqBENRXPhzbm8La5LPYsAId+ECHfLqo7Ti0ZHEv8wROi
O9dMLlg8S8N1SG82W2qfIdENABpIVLgX6HebfwevWCbQ2g8lZQrKvhGyN5Y+X+vP
pyBCmJgpv/A9JhWky0vY2lHv7neh/rkb7BZVp5bh6tB8FFhWqugcLc2J7mGXqEPK
2VZIYK+ZDsLEEbf1gbdoLPTv2zcO+TioQuSd249jTfAZShf+WtluBdWWp0J22ldc
iwnZYECPIgQC4jP0rO9L6M7fNZVAFSb4W5ja0LFphwXO0ob2qT2hGNG8P7Vj4iV+
ZrwtR8JbZX4v2JpsJBUSMPEJ/hAdvqhjfsQSOlyjpX3Zbs/4MD5N4h143qU0VrbK
XXnmstt+g+wb7ikoC1QmDSSAabzGj7uncRgD+MrfOAtuUY+V9qpGLC6FLOA1tzaa
QJsI6lFvTrhtzRWK0Iw1gPgoLTp/nACp6ToSEjkRFnqbdeBLPL9Kax+jx+vcbuZY
5WfCxm/0SocKLn2XteGlNVbbj8Fx9YZtzTJ/zmns3xirZ+pD713bxRQK7BBlmBtx
DPfY06kO0EARpPQL+QFW5rxoEbWPHeRTcT3j+CIzNkZsrFmAuXHXzC9aNtfXo7ij
doF/bbHGVXV6sEArFPfjZChPdShKWNBB8v++JsoVp4TiSQQ9ybPFrYzAki9xOuBm
Hl8utxGivIjOOSYU1iorX4reSV311fneOLF6zL2zF1fT3i1cjFxkFRgGWW1Lpy+l
HEcj2D+8/ZpheJZFVupT5jO/8u6quvXp4LXaynSYxIDtIwEkDUGKoY8p9vstQ66f
A6/s6LQJLW3GUtSCDTrg62QAOULW1f5S0smNR46Y+mDhSEeA/lN5nE9637MGy71a
kow2/u9/yHb0dz1ogpm8lAYQBO9O5JB1CY6IctnObE9j0WSu6H8vQNG/cgngkc86
EjAh5MXPoaKFAdw2Fk6YB79yKv70NOindNyKiTQXc8yWdCY3prvpbFiLHklhEwXT
8spAT0DbAkSoIJx9bokkTqQKKHjnU4dp6r3e0+jfQpOL40SgpLb/xIU6RX8EX/Jj
mEPMRf9n8xVl3epJ7vpHZHWTJ376Ge4mNLZ81O0qce4Ctb1FixEfjOob4OuengPu
tfwVm+HOwjTnm5hXJUknegoSRagteN+aL0YYiLTpJ+BxIgFXFpU17uWV658nmDo9
5W/obVALrgPKPGtFyS+BPYav3lM+NgW9abOr3b2l30fe7ZjIKjfPROKSUvpk5kIX
Pfjc9trX21sB4akvHkA0BVk4WdWgTV7Eh/W/2MUd5aphqV0x9BsESSzUKqKf6nNt
vwmXYL8h7GUQpmvApSiMhXvaWDkjcxVhCC58WUFhCsUinamf1duQKRsFrLXoQXli
C1i+gHjbCn0EEahtsF3SsWhTh7qGLOwizlQ8koe/ru1+ts91PQ6boQ6YQFyPRW/G
zBjDb2xvpI36dXZDUCwokNRD1ijGjJ9AuP+SJk5jMC0V58Olwbf7xwWh2qG0ZuB1
DBCa2vGrjhug60RL64GbRibOTz7SyxoAHmsABdlt0fCuqoRs8dpHsvnKUQlDpPcN
+g/D1YCxzQVTheqTwzsbU0T/50LGL4UgrxAwyVil7Lpq4eUiomnqVDIVD9lUviYD
9jXrAW3AL6XxTreYvexuzyb5XHnCshf03bqj0uyTraLCVzgGEosKf9Xsdt6otUkp
pYmKS66Wc7rLQzJ4zfIZUp5xHFVUkaRYET1mF2RKQiv0LzDxA937Joj0+sztOaGW
pi1D6BFI4BfgFwnFhDdBk1+sGECnLt5Ln0t+KLy5n7d2Yqjp/lueHcfFWI2fL7z7
507mjW/9+8+VEZJd/9nI8c8ZXc2MJdzjFeSuU1ALf16jaNDmmLWEtda+1sKThaCC
WxGAAYxDqZydyWbCpmWpk1tzO6F3z002O74aDtDN//ptMUQXmP2j49d6LC+Qzadi
2y/flqpVyX4OSG8ccZ4EvIEpYv8nlmySUfF6s/k9GksUgdnP2GyzlaAPceGEBLGE
w7gz3iKqDFgoUet9x94/zdTq5mvK2SBF1+jMZ4fGfZOlelED62ad44mfCB9Zd93M
86pWPt6OZ3U+XoII8ZuuLaEa6u0AIOi0kSAZJJB9fQHekmj4/cbW+fBSWqU7Wxi6
RVPFViT2qF/v0K1uveznJcbHjTvSZ0oyR2zp4tUQS0P9OZQoNZNQo1S/f92qZ6Vn
jdKMhbTs3u6UpXR+EbqzeVGFiG+P15NlVdsjJCguU65OaU9MbK6Wxw3YZikcp1jG
X+pkj6TE+6ksNxSwKYTDGOqc4Lg6NDKrJmjmGpgrNB1qWu2r3SWocP3NaXnqeiCw
e6ciBPhtf82EmtwTjC1vH+LCzswJjMLCZahFKThT/R4VD/gCKo6CW0QfLzquIn7U
Ah1f1EUrlMNZxChm1Ra+RDkgK2xno9lnk+AxFZrpIIZWB5LLKozP/25FMIUF7t5h
loNIoXBPyV0F0En99LTNTDSxk6uey6SnMmn3Tly0S5MZC3ByS5V9gufbgSEeUSVy
h+75k52Pk2OTXh+axQl9u+GcktNBHdfiTG8uAKJtDrGgDqZ1AMIUPUVRruOgqVm7
HjwG9+LW2UgwsBqQkHFw1ScbzanZBGWd3wXVg+esTYBJT101a8R+okqfoRIMRNHn
gXw1xnXs5dwYfBO6J1jTaQclS5swucoDiWas6wtuWqbNz/XVkWxoVlQsrdHj0Gaw
FlJSkMHoMqfULnyJu4COTY/CsXD9SqdS1cybJOqX5lUhHkW+XPWORHvBsHapa3qs
lTYTS8pSSi/0MZumlaI9fzyxXQyxNXwugta4r7WZi6rORs4Ps1LcRQlqb44e/jPJ
amk9lfgOQYLDKmxCFAiFpxd+/LVFQ9oGxNsh+KPB0L/ubx9iWAXokKosTwpeLHuM
PGeyJlB+4RatPPL9tyhLE1tPtA93Ty54zdgCdHyhHIBCFeMjH5Waikd3qIHKrGOG
JJQO2T/U65jl07SFE2P4PGDGw/H4+0EluF6tzY2H094m+chpFd8AimiDPWOHdkWv
jccZG1CAEZV84t25Cb5zHRQhEaxOPTB1toqdivHvoQ6rsCNRc6VSnao47/OcGBX+
K6riK2qiESpLvVSj9XWPERLkU0ZiAB84gAnKiRQj8vEwu37nWKqExZPrwI9780PF
8mTHOMwGGa6Z8LC1HjD3LV/ZScctCVw8qeEnmc7zx+0EJC9vYIrq2/Cn5T7FuX0t
h0YqqVjGVdZrvxalgxN9AyxIUhsP1ZXzGjYFut37X1GqglQPyzApq2tR6JWG9SnU
afa/HL5+SPO5K4BACVcFBXcZqRZnQMrwqjAzx3XZ35ypiMlQ/fwFzg0GvB40MApU
3wV/jJHZaxGszF6MjfPxhBf6M9iRY69U8GHseC1Tg8VPtfVrnwaU/V21FwhpWl+B
Njsez9RSNxbl9tRq3ty6zmjyQlk41hwDREaWhK/culMceLiTT5QwXzhYCUrapic0
ncDaheI8nz4NyywjKYh8o2fBGIdEPS1KIDKO6K+iBxVEmQpLeZJt4AQ9MteiiAv5
hW9T+pAuZ7xfVkVRIPxMWNLP/qqxdMKqrLNlTsF8LmxyMFmRoL4r60UwGSrMmZ2o
KnZNxF6kxBpLjVvC4YoMM+zpCf99V6AQlW+uTfYoIRB2CTVPD9maTv6rWWXSVqsi
95dxUGF/bLNE/et2YBIq58cqqIb6izPVKFtq7RSkemqnAXMve24qRGBkV3+nIvj9
hvib6hOilkbp8wfzyNi0Ung9AlZ+9Gdh+OvhPTROfOY/bas6SV/6sMNCcI1P5ngV
gKBu1V1yycxKoWCNFaiiq6B7sFidYA4htua163jdlj7bNV5kmwM9t0yjeqSHnGU3
dOt/0D9vPsdbw5tL9GzO6Ajh/NONpckMLdqEvYTir9JVDJNhQCID/dHssb7hRtqN
XhzU0D4BmmHwA9M5TtlNe3rDvdax5lLCeoTjEyIJ2IiqsBwTvOrDTfbTgLwUnYBK
BMTqGemoGVL1hxElUEQGxsHyEZmwY7atbTbf9om++1WKMoCvjEv/Ls78UkZWNOQm
aaQoAqWeLXmI2DRtdiTGiDVxoFuUrDEAlJtI0mdxMuvDXwIkPYEcmEfNEkvfRy3Q
MhXLPzLWvwN6MpTgld1mY2vHDlneRBVk8BNXAeUItfuGzKopB12+0Upoh3splHDF
upwaH/U6sNTlBYAURtUUqBJ6pVkBb9TshA899yo26VG0iaPJDimaFLJAaUAf8M1y
X1uSokJmlbbnsdyHaovEXEOMdwGpJm0MH2ahSQ4kve4vRVBg+Q9lGD79X40YTH2H
ARxWaN0WZim2gBSgvGag8BBPLtPKz+FiNRo8HciajfRRTdO/MJr3egSaNHooS/gR
sf7/pKSDK1BlP9jsbpi9hI3WCoUM+bDVZFBpJUfTgDRFTO6a9xUOKmEUAywabTKU
zp0vuLisk8PPhZx6+SkyotNGBKzSGDslw5yLvjfUST9qXHSlIYOPbDV0w+Atlh5m
YQnTieQ7+rEtnKMZDzU+YjDs98yYyJEaYwSTXVnKFjbakS8XEf0mTZpex08dzzFj
XNemaIsIcTr5nMJXt8uy2Hrb8KQler6PqctEjEs9hIdtgAOidUs/ylNDqR8A9VLF
ptl+nZb0dn+0CLG63pJC2y2/0JU+s26fOt7RRCN8z5mC8rPxiwnBrVTTaTvJYj4x
LDZAECy1xr+n25ObsdSTUd+ofQ7kGSj/lIF5xedM8jGiT3OKXB5BUDUT/9aNTDfl
16yWADZltCw1z/WYoPjhtuAEOOWBuEuyj0JbMzz+Em5+ZBjn5RHssqZSstnpqs6t
lLKhoJQhPHeYZ0k5EmEXbKOon5rR+Wvst6wn++yxLxQlaXGgRZybyz7VQtRpskyO
nWQUsVc6lgCMoAUKGdTPmIdoBQD8R4mPaJGAhXDgEiXAEYX1TApstryHrGzwc2ma
jLQH3G9Pu15praivk7jrU4nWR4U29+oDho4lI29z2/ruQU0UoJ0JfduzDW8QgCyJ
Jn5bVFVlZZ9lPDTU+ob2BXMco48j3P5Fg+Qz6iMJ7YoiAOzgrgmtdabVT5Bd7X53
k+O20ZuNvMaShcMNF/XWs6cDTDfcLY5S7sdTh5h1GMDjV23O/sotJlkwSF6/jdVp
G2cq1hPFC9HXvAgSsU6KFpn7JQbOd2f5TbQ1e+bnHYHpusF+xDUAu4kGTEFmnO/F
4aUJpniITwvTaXMfJ7nsFEx6MsyzKnSRHXbGuXgiweyR2G/9hK/5VUCgsNEb5vWK
WleLbdxjGz5a20y2/4BIjqeW7KRWWf3FPf6N4KD49z04FvoBF+ns9sHGpIGlBaVU
vRckyScthmO67tAsTJUAHN1zkQIq414hBcSNYuSVcPNCXAKpH0NPv5CMwpdHGwXW
JUzsfFFXrcjoPKSRy7afQN7vK9IZwtJNTAOdlrADF8eXQ8u22u6ZajJBqz52ASdO
+SfcVcrENLcHMX6ZjZKjWlBQ98vwL3pggWOPXAp07yGisOnqztPqVgRvZ4MvLMiy
qXtp16+BqDlnSRcps8FUiSalO4IOZSiatNwecevo3Kb1zkuUA2eeacwgG0Zpa20+
2Gw+/92N442+i0sr0PfTkv6ykVQ8drm/5ujXg36X3+6R8LX6jBiTrSgnciSEG+sK
JOsWvTIo6vqgemzjraDjYjPUEUjA4/vTYPAhtjOIkjY4RXtcm96DJxupz3v+QIrJ
kIBTxcW8Z5Q4KYr9CBxvU1QgW1jphoFqHluUR9rQq//uzd8w8fT/jEXjE4MuJBEh
Ibn3wZS6ZhFFpvgtfazTJuhVErkjpBDrlKtJCHIQFYcbE+4l8DKsBrE7N76fpHdN
moXHxkHHWtPCv1vZTPDkovLH3Fp34sZ+QkVoCJ9FZwtnwv2pnO3yoIWd+aXYTl0d
y9q/FPX92OlUYLZ8ePZwDi8PT2OH2jO53FNQ/H0UIYQQE0qbG2bof9HCJ4z+D+/Q
iZdFxcQRuqjtOXSRyqgnxjuodg5wVfcQVjoxESz77I7+w7PqA8wLKO6gM33PlEcR
ge6jKUwRPq0+kxEw/a8vS9n7ZJi8jKjxCzoYYUaquoaWqkgFz0xYGuzNgr/dSptx
VdD9UP25fLIWoOzeH5YgOOALaTcDknprbbZOuC95unt7VtiotGoj0V+7VAtnfseh
coKpETYL/YY8Q4w3CXkoMztsksGL6vxPFsgx1gmdxtC3E1fbePQHprlUcFwDNMnG
KPaDTRZc1sd+zdoA1IfnNPDX4PBHgGxhO27zRtBbD0BdKDTTFwQoVzilwgnYS8dK
GF7eJunBwX215Lv0wKMKEyixEJEJawtb5YH3Sn1HmvYt76cCoO5K3sW3xNIpMc+T
EoYMAtE/uWDhQ2Lf2FQMIsAUgEwAIzriU6vbVqyVHX0lBvKFjOU4Z+4kiT5SxO09
GzNS0GzppGdl3NsW0PASE59EvX5JgDtWJFwg8C95PBFuWx9GDnUB12pH7/fRqn/Z
t2EWqb2xAaOxrl/4biTgs4ldXoilubbimcOy70P5T2dF1dEIIMAkxX28vCnwKLe7
CAio6b+h7rxgu8I/7Il1dVGGiR0+y/lv5KZCDmBEvJe8gOXf0RabXEhTNtr8fabl
I4bgblpBYC8iWRaLcfGFO3IjqSiGEBloKzVdFzhHHbdW/eXyRrCIVk8FfO2vb5jj
XEx4qyz4JeeJziO67X951OJU94A7Ed7xmNdVQbVx3hsPZzdGXR9qFW/j6jb3pi3Q
N42mUkviNB8+cb5ywkVBGnQ4F4kum/47uRW4JCdwZf/gS1ycJNNPRxeGYhxcFvOd
p8ggCSmW7Y2BJLrvDOD+dXu7Bt26pgPAtaccJGRnTO/ae2BiW0LAy5TyrbejK4C0
lRUtD4mP+P75e+tO6tvRv6LrUWOI8ii3HU3dxjhaxEZDVvPL1E7K6YB6+Ea9wied
vpIRQtNA/91qnv+8xpAecs2HvK5w0ci+BkMGGmsCmyfDHo3sFwMAOnYIJWFToV9u
rai7pKANRxKixU5rB3QQhLyd1lVaHivvB2wvhB11uaDBfex4eLt++Wp1P2lyYXFN
2DBihS9ImamfEcJwTbJnb5cbbvddWn9Zkb/K6lYbQEzHvrO9Q5HLZN5OWtGcbrHj
EKbgX3w9U+WGA6n++pYb4S6OBOMdmNs7RWH3UDchM85bmvRFHXw7GLd7JNpxxWgp
SwmNwR+Lz0uLug7iK+Sgsrw+24vXLYgzy7a1/yBRP4py3gMroEoL8qRcIB5LsUPH
G+qhjVLEe1Ht8+PV7RkwkIvKAWi1Hwq+3ajoBQtVFluUUE0Fb5WX88PPvR+p9tqh
RAu8YXTOtrF3Dnj1CtREye3E4ty1k7UAmo7QE3+wp50Q28P7g0o7WRbGaTTpyzps
cpABY1Eg6jsxfVWbfJhST4q6TgZMdHi2Q8OfUHU/0bbb5HecQH4iKN8Z/U77jMNN
0E43qFk5abec017iQuwgy541eKMOenIKcofn0gPWCPo0He4LMaNgOTv/eTOFjsZY
1guLsiKxptYTS1ARuk0m/ZQ8BQ/iPJSz6RlFzVRxp3tb/Yk7Ea2hJ8lJ/f6it6yg
mQMkp7GYAn2uLBmH76mDECrDMaR3FYDxn8TpUMjmsbuk4YGLmd42y7mkfwzVcUi5
taAFCMeCjJQ1Dhj4e/TH7mq9DJ5ued29ZVfqslGXIETjdNE+fjl8eiClt68HzfH1
HY8DkhptAGaDvllEEYpFHA/7wTLkXcmYQ+yo72adXQ9vQvHauAy6+2S7Q7RIbGyS
6ATmsmDMsBzMeWXii4MDiZEg1thypx0cSczcUg/mwd30wAMxiheDhIA0MQj06nbb
VNl2Gsq3j3YE7zukyvS4u10YyjqRfR7+Qix65lGY+mKUv7HfLvCB5c1ZLssyXRXF
CXbqR5MFPvDb/IkWUt2BbrDW8BcT1bhAeIx9bTTKXBW7l7f/ehyacHzlkpZaS8Mq
TpbhUanXiKXB0/T/+tFLIcXF4LXp7Fg9NgtsG5wf2nxYWMmgWo3CPeMEv1Pma1mj
enbW1QyIF8RNbj2b040DmZOzojpgdhBB6f2WxTpG+OHmErl8AvY7lK0OOPM4+NM0
OYtkzK5Q70qqCmLaPeT9iDf3C0+3WYH3tvcdQdBA7/A0mUQDnY7AgkJb9uVizFjW
PrrvJ8H6WnxqouvQM5stR5ADfziIWw0iwIebToCgaaDT7xF70r7q4tr3U6ooGbAH
F0IeqnqyTKPTuDvPZb7HoA25DPWbd/hA8e4A9JixlVmqDdGBM2BLQyCsiP2advaM
UzlobdB+HVQpzoPOm0OjwafkTM1qv/q1lxyqvNxy44ZO0lh94MS1PjFK8QG3a9Rz
4rA/Ksjqj/bjre27ZnPUBr+TFkK74phx8SK1HlOJAo1Br6K0J16Y5sV2zirFG3II
Cq6msQXagggWNHZlJpr81TrT2/uYS5sH9NBzJXMgRfgoCYtcveAg7inMq5fNy2L9
5FX7BvJDsS+SPwQbGfF7bx7oYlWZ4ZNKxzUwxvy08eMwGqR6WdAzGQDLsTfy5gIU
VPRHjeFlDuB17pb9wXCJqo7tyYkJ5A9AP20FR34XHoSwWzdD+H/NMeZyKUvOIwg+
Xktawgu7lRRHDma7FH1sFJoqrLoN0jiAt3q6BGeRlLZO1TuX4/RoJiHnEJXSxIvn
1173cU7uC9vO497qucYwjlkNs9Lzq3x+3sGmb7vEpa0/INorTiAZUpzmX/U+/LEj
zhd/gfLvtfF8TJbBbSqLj7VdMJAuNAhHrfVtwR1mRryCtAHV2C2Z+BJTa2rRFw8U
jMcN2eRhMjzyQZLAjMYPMzTUFncm3h+cNRSoFshUBah9X4kB8/uk/FZMwKzEi0+J
WN4jZaqXyxQAM2Vt194tYodHCtxBFv6//GL9YBcgLNlRk7mi/BIhsZp5JgcU1FHN
tLDX2nZN1SXfPfh6UXi4He8tnTwzkFUw+YyhvNT3VVJzcvJvZ8IEv9z9zPD3iMEs
IxAqjDruq1/q+CI1z+oPVoqIs8zaVIv8PCMXVSCfbWOROoW7yhGfNbmrFcJvlNJH
m4Gbaa1cMNN6b1fsx2ha80Mv/H6/53/QD6ogbLTd4Gltjz6bRufoXJvHE+ZWb4Zc
YyIzrPdVblVC0LCcwVgDxpVbBI5tmISgB3XcAL1g1JpUPhvpmbdymbZDwMki1CqT
6JpmeMjKqK07dTMEs/hYoqvTPrKGqHgCxJgDfLu0xJ2EpOSZN2vfjZ0M6Ma9OkEb
ahxRy8h/PBLEmjDdNSfwkiNvVfDwm6ERKIldKZ4rtEcXKmC8jhnHpfDI2jFcJ9wr
uKzhCkVX0MALCRekBFjBEqtE9LG7EQFqWMH7YX5MKX74tEjzfVtNfCkNMkZt3bv8
fH5YeOz4rO5joOuV7YcwloqJvtCxBD1RXmgcqR/y3uMFSnDrGdEOGESqAwbZsaAc
K9Tu/qxJxp551ueaAiDgfSHpisfn48rCs3K5hhcsTpZzm/mUt2iLpu5il3AL6Wvd
5GOoBCrl2SKV4+l6AwkZiW1wrCKd34G2Y6IpS+jiWN+MybIk8cEeiLkZuul0Oh8E
6JVeNv3q9ktgbsA/9RsFx8wgjhB7lhVhexqBefqyQ/nJi4bshouNFfml57QPKdq8
uOKeXjf5D3rdCdatrSFFgoxB4BhFKKiqT+SA8BEsmv6bwOp5/wjXAJw03vzAwabx
JbsHzUFbaOJ0kVryiTk3rt6Yg111WhL/35LUiKvjIXuC1IDnamtRq36dUWCHtTnC
vDeGOoiPm6at5JSMjzSrE84yTajRqCV/zewPrYpNEpM23TqsK88woTWIDuJF0DzD
xzabTsO2hqbDSX+IpcPm+KiJjU8W8kZp61jbtD4sCdTrJYf+A3jIBFn03PI3jl0n
6PfHYYguAmjxv9T1msNis4bJfRDWt9lTtdCnUcEoRAP2szWAAcVAwF0oR+DNdUSS
PpE9gHtN4deNsUGk9/TOHxSc2nwR0sln8NB/q+yUOomFH2feudxdokO36Pda2ZC4
hsDXgb/8ROvF1fvQMuWMdWF3T+NBvz6s4n4WqqHlPL1xp5OhWNT1ynOs5kBbgO4m
Vdel8esrZtJZyUDz9Uqis8hbg4bk++I1yUJo1PHFpB5ayCeWJxo79Q2KGeKbFOdb
g35ny7p1N6Dw20z6yyll5ZAhlYFqk/mm0WEpNWIat5CuyX0TycKBkDOMoJS6Ec/k
6TtdBBYQrBR8qtfybhfzFE+pTrK7hDvA3cy03XTdrg3oqDm+6VsfVCMDsr2FTgok
VxFSMDYvg1HDeco1vNFJOpQQiDZ6jN+vQNyT7q8x4xdMKOdxt2R1fTL0tPJqgvNP
zqrdYl7IGRxkNfATdeyy23RyJAgQI381/alAHOQMZ47C+s3FrKi89V1mSCzMUfFJ
bfqX2zMBrcguymjhk+pI7AmdD5EeK5JnHOvIFgm8XomJe9l4cHK70k1UEFu9f2mg
1ziJEZ+f3brV6Sm6ktkZUrHTKZM8qBuYXCT/Dfz6H7YuODf+QJk/ML9hNddFI12i
9tFMsOLcw3OwUOwz3T1GmR3D1f/NHvr9gN1B22X6Tck6cWioz1rrov2b/CqJqoGg
0sywL0nHipAgdvJDImRGuYD1f9dF7ng7C6DmUGWvgClEx60WhPL12CUhmy++l0Qb
aqOXYFJfaiBpoVKLSIeSRAqdlaaBmwhT1RBBx44NoZJ09tBgmpL0yGk9L043OTpl
LfMEtyqRbwepil2U3UpEM+o1wg1ZwRztdsDOulA3OuNEPA0hqhjwrAk0xIhKOM09
S2xZGFXwZXJyIFmKXcCimwy9MhbAaVspmuEDa9gh9wf03BZgXwUZRfTGNA9lgcDm
taxT0XJFXHUBGCi9XG3jqcK+f7NeXFfi9TahmoNLgcc+XpdYussn6RaXGYmlGcBi
KqHNMiJrkPS7///PHM9x5sUp3eAUaatclfkc64xJ8g9/jrXlOmuy+OTVhqB9Dzg3
EcB9wG/2pG2n5WImmn7e9VRzAJen6C6hVjEgVlVzF+g94tNfWmQKXciV8p/50qUi
9qX4ps55lkimDPVbR9M+WkAXDKLPLxk+YNjuv/4jfiKw55HmTZyKnvPOAxz3DN0S
xtZUHKP2dw3uhT4aGYCVzQJPyeeM+d0l1yTOj2uFR6sl2SjYP1oBKg2bG05mZsOI
TeM615a4zRfGO9bRhanrs+lJIKVlQUwhdWu5oo+dEBBTK0S5ywBiDCpDPFSDH8Nb
sS9wJiBmVLt/aIammmh8Z39RBJjeLAZZIZ2FJle2TK9GmBtJA1DitMLBQddQ1GXh
bM0NzZkd/5SD9bYNPlKmO6olSqUJCY8dYJU9t7DYnSD+NWCi7R0RGXj6OLPjVLG4
WV+2gnXAb6W/gooTTfZCKRixxvtbDnH5SJOvmjPSvgJlwZ2zWpYQtmJkYcRjB680
5T779jllyFflW2hi0J9uxfODAuj0+2oXg0KWduwv5M56XscUPCnlkdiezoZuI0T3
GrfP6e3J9S05vW+CnP448xmZd1Zc4I5xS9co7ibAaI9ZTHT7I7eIpcaEB3V0KhSY
ulGJvSrXi5EU37BMIclxmvdGx1bQQZWY0DNL7AZt67C0ACn/ZwwuisfiRoCkA3WC
s41ExuPNK7SFCN5mE1yZIGGwpTXcoA/v2UIdD6xGBfsEY9/wjoYhS6QU0rO7/RIi
Jpf/fpvcMV4FgDgV73W2butdkvaR0M+cd7206QmW44gFIio7oSx8cPZHlQY1glSb
hho4VOeAIx76fTFNqIGRtQOYImTITQ0ryVYUFCOUBd6CExwW0lh+DUhhfbqj6YfV
1M+mLKRDB7stMX7pnmJk2DV9PlvFA1g+v65ihZwnMHAs7tUFzpGEKSS7aOvjKYU6
J7Eursj+BDhqsPX2M6TMAMwGgSMyBw2GsWyNEp2Cb6r1m6n5JB6KeVVL/1QSxpko
HmZFJUeDXUx7TWFl5quj8XFqOuSfcaHyNUvVuO4Bzpd9Sbd2XAu7jhQpN+9hHnSZ
KFWbLBo4AK9FkpJ4v6HsZmUMDhvdR3JmWgMzZhIjNiFNNnuFUvRDqqdJ0vd9XOlL
vvpjoH/O5SSz3VWibQuTZWQW0LZY7PD1vJ5aWEd8nkkaCZ8YQQdnSN/pI9Jiv2KS
o0oKu19uftLiGFafmPUWWAzVcEpGUr6OC6CWVTSarCJgdp6CRtMGH+b2Vt/ndHe9
3Ayx965Y06qHxjBtF034j/QToudDqdhfqxDSGYEOrvJMk8HXQysRgOeHEOKzEqpl
J617NSY1gO8Xt8weaLB5lJlKwrfEbwL6LSnjYTr6F1vts3KNGS6f1h9aOo6hySSq
5nF4xhfY3+/Zmvfewsw8EURmp2C2ckuRsokH2U0NB1Jb1jUhtI/ofhIdH2F3eUH9
NZi9s+rAc9VtSU1NBxhXHCrwxPLJhYl8fR+6rF4WCyBaJszS3NZyWTXNst+2/JZO
Mt0q6f5J4TO/l3/LypWfxBl6TQJxG5lnkJ1lYkyupyIXrtsRG/e3seha5+8dxThh
RVywpqJuIb/+mE7g/TcM2HmSW2hvFvDed3Y+eQMtKZDc8e37SyEzNtYejz3LMl8m
hOpIFxSgfwhkMLEh/S1xvaNFV7jt9WgB/8YTn5LXjYwr6LqLPiSm8Z6te62xktxo
0byyNCuOQ/8RPZFf+4VDWS0N98rQa64rkGNQ30uKT5s7stWRX/+G0ZXpVf4HBjhx
Bp0ZPtuHt1NMvnXpwXJHRT6AZaAMKG3q/9/m3yGrMQu2jpo/unp/zemRILtqRLv3
UjIXBTZk87CYcfTOQxJrBcV7DhTrqghFIgBF+BrAFdGnv4s2NOesLNyaW0VTGiPz
AD6E0qHsWMdUHNU0nzgzvN4akhEs9RAZD71AdtNVVwHebKnQ86f/un9LEBzXnTVT
hSXw5hExgakH+IpgT6H6WMezGKVhuJiyQ7KwuaD28Keba2KqWVQUIUavS9MUYQHf
/GRdOiFH5+bV4yh7FtuM2l9kXw461/ABGDaMlrnoxIFQP1SPhA2KH15IxDayuUfV
3WOhrFetoCPm564iCcPZ4UuGvLKl8zjoRAh291WuJN5FbxGZ8zExiScSSqKoxc3D
fmy5TsPWKqWM3p61N7kkC06zN069GOMwuhWET/ARVHGatupBJC/MIObTBPn+46az
NP9VR8qdGp9F7OfkjvaVvqdUAWs/3MIIA0T2JSzbHF5N1PbF0vtOXYjT/4+lH7Kr
xFXI1O+cYYw5j5dovky+iyHzplq8X7MWTH3qvS5+6l3ksMVzxrww8mG0NNWdHWm9
eUgWjoH/dClnaNW9hOyHDcmqAcutiH5vNlwjkwXE+K8PcJIhxXbNoKBq2jR3R65N
faHVv8nC60R/YnraYBCwkvuFDMjQ2jL4A19uJwf0Z8rjM793kSd7W9KoePrLfJ3L
wb0YRB8aXnF/+LxJ4rqyI2Xn6JPUqRv+gvNSjc7Pb0tDkjXTs9GqEE4U4tqhHm4q
sU1ENZ/tV2mB7d0tbckjlDbFi+Y+xa+30Mdg4m21ifQ5MhxMncu+uCFy2UU1X8zb
6Pb25W4pKQrAkjxCTH55aNGFKy+8B5Sn1NDpG4maT8QHp9KnNjtGdkE0giW9W7dQ
cY/SeNWXfQtCJKCaQU2Vt5+q2fn3H95SS5F2AGHf2/7mpGou+QjZmeTZzFzXIwXH
CdWog8wgTc7Q2k3e7erXL2ctJOm3TUVFkK6ZVjqFc/rFCocXnP1QVPcldB4AuIjF
AbRvpOUglYHPFsu/SnpfqzlgJCeClhB0ATuXGYxaym0Fk3XZvSL1l42RJg+uovkB
M+flMHqFdFS/P5yLXlxtMuhAPKzCVUTYvx9Ml3m8mEgsylmGYV/pv/KStMQyxDFU
8VYyU9kqi18mLz6lkeIAIZZ49XqzTUOnC40pZ2kEJUnKQ85vsMLIr9DvpUpxSkes
mEQVFYH/ORYmKlvZq/8YFKxQZ89HdvQM8qFgamq11vNeWIhjEeVYzOOZFMDDF9HX
WNxfWh4zwTus+EhRPE8GRr8Lq6IdoKI8UP9dV5R3WYM5pZnIfvroVLI0E53gYg56
jaDcshlYq8rPIv4T8t7l+5iTb4p1YiosxIbnIZLx4cZgYgdJ89u9GFkpfXoTE6SN
Ty2nvIG/I24o1653h02O4zbbCspBSWbqe3MrUeTdsAvq75h0+Za9O6QMeTSAb6AR
AUxACEbliADVPgY50yqQL+40S0atr4buSIlVNUS+v5zi4YsEanG/0fq4C2y3QqfE
UaHDjKt+Phzokue5YBT8WuCzji0qbfjgrhBbn/nXxZ445QG/deqB/5H/5G61o/6/
PkWAc7xdn31nJcb/uPChLWxCRFhTTHyP34AccK0gmQnQYT/mV/myW6Tn7CyQgas9
+joQ8FMTvnFH4hE1fZ6m7pSQRLg5QtcoPNgs+HXFK1eYYRG+tvUlpx0HHq6wqP4S
dinEtkRRsIjKmzuEQBx4pXiTzlbBQ/+xXYDT5TnBKs1fSpRWg4wjtlm3R1dIaXfb
5oKUp1BpiZhlN9ZTWQve5sLA6i5AUV6kr2QZ+PiJrBKup4i6Fo5KveBajVNHovXE
dAPEWIA6HAGxyxFhNJ0q9Cw8Y7isG48M64BcMDrzsHxEq8CQmBYIdtq2UCxd46o8
saeqhlDPIofvXLpQ5xcwqaG0OMqjgwvprEtnwBJ6Da6I6ftpZJY0Bi+Y5/kbNU5b
1rfAiURnxP466YCX+GX4kxrekGN8CfI+opMYPbfryT2B0x6m9LzUvlTAPmveGEOE
Q0TL0Y+zvWg2gQY/66PxH+d5dlzecNHfebUaULj/2sc/gv9eLH36p52D+CxsYkXy
qNcuUpjL7aiQAMjQhIb/HmCnQGsypAU5SJ7T+E8lFCgKED3PDrj6MBIJMNGNtqM4
XLcEmgyhaEs2gpkVNDiL44QlfuhdszfXQev9spLjtOAff0PRut/wmTgcXV46daHS
m0NUSlLtit4t5QZDdAuqkhbS3RShL3i9q8Q83Si+V8ZtUaU9WafLekplAaoxOfNa
npIGdQm4NHzXdCL2RFXxemFbrZGZlwZuJiuNxwft1R6xWpTWBJ8uSqpwwzmOVBus
DP0zJmtVk0bOZ0cHA55GASry2k9WVlIFfAWUWtJtXfimOkAJZ/8TMEoCkkUGZp4g
CuOBEmf8BJnUOj6i7CB0Gjsje0y6OR9q4pK7WX5HS/hb4jYVSLJVazfgzqYYHwpv
xhN2sVtS4rrkBzLwpYhVg1UYAGR7txopybGFbEtKDI+6P/JWLV4X4IwBr13IqDrD
6Wmtd2HL5hT71jHOlJiizVUs+uwPYMeMByyE3aFq2i9yTvlA2uW1bK92Pdfbj6P8
r82Vn2kWEk3bWkeLUMTa+oYen40DT2inEJAUAfiJUFShcYOrvPQ2PPIEmSST5bbM
lAvLwAYWdo+rx6Ff5hQ81TNHOg6c+quOu/MOKntAGNmq21EqkwMZ4hGbWvo+VV8d
84wyQT1oiUZgkdLOLzTjqGL+e6NxfX/yFnuqwO+rKSKJzmhfxtUeJctZO65mXxQV
rWnISfeYpmm35oZHQ7x+dfwsEje6WKa3Nf2zPtF86Nl+ZCGSlpXL+DyQEWSPbZLn
0P/vNFZzaaRZa/kcFbu3QHcrzHd0kIRpoVQT9oOI9xRd6AMDOfGcD6luRi8Irnpq
RCikts13YdG19xA6ZgHFnrPyU1BC41Xs3OkEQxWxT75eYpHsZ6tpqJ/UPOInLOoh
r/J0ns/IOOwdsqslUbupsgkZDRrlKwx0lKNwhCif4oEVhJgYYyeWkThRvYNrxoqi
HWaJ2su1gXNOzMq+yh4qpfQFtxRwyxP5kU6yeKUre84vDwKivKH3DXG8ZgylLlIv
JtqncPfDGL2uqRgwAlgBH5M5z0H5YsrIxX0e6kaRuCEb1ChNQwLVPtHlFHTSOI5j
OKgVmhfifiBLN67HVVYf45nXKk/gPKIerIbO7GBYGPMKg6vrJPxxSisy+wEUw9zB
xEzcHvl5QOV6bxSbmFTn8DzRS2C02QK3XPujDHNFAtQXsdouLO6RhwM9vFDgCvQ4
i0Wad/EnDnT0osYO1oMaokET7JqnsHHgjZUYmFUO7gOoBdMos76KC0tUeVtVaZf3
OInW15sb8zG4u+OirLqljKNnrbMzhtKeFVRBehLdm+lQ4GwO/V171GTIHuLUNHmO
wFpaLfZpPooYg36q9rSVGQ8Qa9p6+GQGvs2RiZceywGqG/0KbWY7/6uisSRo11WN
V6blf+Xw6uRv0xD8s7Wzyg0P7pAJY616R7QLoGKhut4y+MRM24vUa2u35ehVutqd
Mqyn9kLdvsSMVjD3SOIx1KLaKSf1QFBrM6g4E8qBFOVTdBWF/Y6UrOWQq9Tn3N6N
08D6Mfa1msM9vX7Ky4rbX4s09jTdJif7aGpcokmw0rxS6+KEtNanQGnz06jNNVUd
FteDSM6N+1AbbvtMaWoFUAEBgOPSsDel2TnJVfyglcntsypPf9RqEhERGN5BkTI4
5p4tL6LkW12I3PpGwPwBRewg2OHoId8ArHLxqdwxVLP5l9ww6DyyQRKBeRBPXw5H
tls4tz62WfscDB3xfaIQ7iMgQ8cKkdsDkF+cKLxrYPPFGmm5MjhOYnZsvyhuzgZq
3KmXSouahAdGsSwq6yUm6pM8vX/vFO7JqwEXN6SZZVOWgETYWE1306a2d1jrw4Zy
U4l1yro5yrBR4oCF3RXnx94YnpfuEAKAsXN2tIJaoMy1my04y5jctL+yDX15Ovid
D8swCZ4hzMDtBNPvtYQQTpjT1hkiSpmdyiYyH/kDbDAjJGKHUmi1VKZIEHPbVszl
KsZScPoQTmxQELlV1GyINFzoaSm7Ac47PH1Ixq0dKLIEW3zMqsInN6tK+0Xk2Inh
LD3RcMbXvhSZJ4boLSRPSnrQUX9Nmwzy52qdO3/Wavw+cXr8eXaRWgDn6cV6s4HI
OMoUUjQ7DmFcJcdJmJp1jNASzJ3a266aTxSeRSUW06p3z/FV+MujAF+xwFSllSqi
qZ+O7RelykeBNxs65xv0JMxIgCzZX5rwpk4PgFkApnHvynBkbWYIJwodtem+gs6j
VeOmHfpzpkB/urwSYm1TJJp/n4GY+cASn9LA2j2jNVbBR+gop9H1cWDwdsG3pINM
s1fqaBNkptTUMQ0EJ7kU3zuRR6wlWUl4GmzH7Xtj66yok/Z88B8kus+2uS6c6+un
YcZyPgafkHxNKfzZgO5JJMZS4/XoUBTLqgEvL9CIWZBDDm/F4M3KfTKxVNQKhnTH
BdW9XwkVjyyoDiRSHJ16mkFbuaIHUSdzdSdfll7kkThj1zDj0YV961ETeRqJUQUL
7ivCe+H8ecPuXp+yXFirKsDtnSEmO0N7Cz5DNKlaDp/mhGMckg8BFdeUeh2bv0cy
gPiri2vpFNdDsKlTuWLaCqLA+SfNitJyn37Jzp1BojiAT8gshZD0HkGyP8B7Ihrv
FmtwBOzqF4caBOO3xly7zuH1QMgiPQMw09+j22BRjVBRLRNsGnBYAZm1Rf86Yroz
AF1UDeoCyWpReMmR6GwiUq8/mGPKxpxqSv9PtbV6c58AZP5f269fZRM4MXNZ1mzT
0ZoS7worOo7rNSidXDQs0Ts/fj6ai/tSwlcwIDX706ysPC5WMG/86YUkTd7c8Dw9
Wa4MkGXCIchqM8ZPNuaFtmiRCXv+jLeiLd7vt/CreGxF3qPhs83yRDOGH1/TLKyD
7/baS6MxJUfhSBr9UQHNpivz0vOhsYdTi1eEfCO6RuPH41k0X4/7uCDiE6aEBm+v
nVHVy7uFFFcwyL7RoHDmqZSx/vPnwJew81uFn4wETqnqASjiUKqj+45QJoyhXhPs
GCWgI2z36v04yU5cCx8mmEPPK0ai4ghyiCkLK+sTVZVwpltce4NEet8M2X6O/0No
KKSkud9+kvcufqr0OUM2dzRX5cpWBStGfD8CY1pyoYzyy49qvcWTB/wjJD6+y57j
y4lKbmj9f/3JZMHQWr4tz1ostvGqmkYOV8Ae+iEPPPeW/6/h4ZtQd/eU3F4itLSw
P6edhYkxMbswPyGBVqEkV+vGfs2YIbJhSNrAH6wW/W9grsV6SpnuAPv9nL5oxHZR
t4xFBb2FFZ2pXETECEoyfj9D5rzUdvTxfl0XDJWN7zFiwJTeqMOx/i6sfsMSOcSq
EMulOrprs6noXN3m6I+ME/+H+gcTSLST8M/DmwLhRHuI7tPCUtYvaBEeTJvNiO9k
gtWxAwsDsxkvno83yJESsqvJGw2wWoWrFxuiv2Se0P+b1UbGhFfz8DE73Xc/Gdyl
8+ZlASaUNwqO+ENqISC+alYqGn5utm13TFZaeD5+mSuJjdeVFDjDlyBcpFuoKdgn
iyHisW8Dqk8lg5JZMFTuitXEGl3eV/SREPYDcllT+0eOm7pyug0lpzM8oNTVFDfs
Bkfm33NDoMs2Xzu27H5h7AF3l6i+4iyK0W+XS7etY3S/XekJTzavB9tKKludV8cK
aFZPkijPi2Vg1YwQjE0XMXvQYooS/xN6pRE09DAW+pWAGNu8/q508u+fXGPunP1M
lCgEYSQThLyXUGSo5CChzWtOB0Wp3VcveaoXy89u6PU2WhgtTrdB1Zfkw5NyfcL2
xKNeywV2E4ctl3LzBJ/3MOcnNE0r8DjGjb6l+T3q95GIvRW6C55LFVCdpT3H47In
QQrlb79F7t7IwEmBs1+dIpxjPlKSDQfkaW1idrWJSDZthhIy8DZ6sOwaqj4YHo82
axE2qJzKOm1BH38Avu1Nov2xXaUbLbxEUvDOtRLiS386Li2eDLMdcAMO5SwpDKWD
PmXaQxZ2oqorlEy212oaXX3Qi6b9aHodH4H7Ja6mWsOOlJqSk2yvkRIH9wy/ss+G
7osmEyuHL4atuEQy9mZJE263hQvoEOOXzeyprOkbJT+fnptIipnQF0FJRo2O/UVL
YPFYezr4aEDxG9SRV/FO1FrIzrAgD4BX+UjeJfvUBaMl6c4dGQleF3++FPxvma/w
//oXQjQiYlcv6UTKWksgQAW2f5dDjEI2aCI2dcF31B7FthU/nYd/LJrrzTCiwKgj
FZrGzCNd3uZxff/fJm5UhEIXOlbBrdkIYoqPRfOeaLBLNzBcXewBo9OSix8LOPIw
M5JTQX6kCID2tOsTaPa+5h5VrT5MLJHTvxvAu0ozTMUEnYFnJ7i61BhG+3lrjVc9
bFUR9zrXwSjLyrLs9qey3ZJZDbtudC3CIWkjcBYRp3HmN8RqyIm93Y7TF1s72BPi
Zl19pfm604nSiGrum2+UYaPGYTIhBUzC2ClI2YnaRyxpmY8krNsbyEQWBZjSYN7O
Fx2IEgZgJGwcEo4N2Jq+cXLC6p/hPiJBAGI/ZtvkYZi3jLCZsenJCKNfxE1EiAZq
yPkawoe7VPSfEnV9OEZJl9CoTyvupvu5P17zzDtWpoQE2GnnoZzkC5cc8R2ZDCTC
yXOc40Jmud0GrE+Z+GYHRkKXjJetrUA91FBuwMJ97H5EYQ0hPn1IZ+wIswleIL/G
ZvPyysITDVN7N/rDHUlwZI1WUEvSjVyPWWfXFr1cRuB8Us4PLhwXIDCIADTtwSdA
dBlCruHk0aGW4QPV2iCOv7zsdzR+GzInMXt2DxH1xsC+SqS4wIGKWL2a1Fh669pe
OnVzdSoPIAo9d1ol3MfQPCl1xYjgfq/b76qttKvcoXSpc1uHPKIWyNggt9efe5JG
/qJBRzIuLApD1Wj37YlMZNJ5P6ZEU9wtW1rtA41jQY8gIXWQ1PyfNLhrxs3d2aST
BYJH10H3W14r04LyqMcbGyfg2f5epVsmho2UgBtGz4tyWumIlwBt/EYgjtKxAKwv
XLecWicMz67vPiMWuEnOkLdA5IURnL24/aeEuBg+0FZPVMwkUsINxb7OziwkLW55
VL07Us9dmP8zGyq6HQDBtoVrgQyWcwTbPPdI69qEGojhSlCx5p+ANnTL9R8Ne/LV
Yo4IgWmtH0DI/wSutVfEWdxdWZxMqKmR8HBfGug2BsbQFBmKMcxQ+vf39xiw8vKO
8jNxaW8vadF2PBbdj+FpXN9ZwBaxpaHPH0caZKRyY/ekb1A2A1LBGBLM/E0jglXq
Y+cy4M0YEahzewS8z8s3N4YUvys/5SIrqpLbVunlRQAcAbldNdM3EweHcZIXwes+
ZhDrlZ4xpgtiOpLOSoE37hL6ue3ZWTcy23Cqrfu9jdba/8qUya8cwUNjDdWlIr3j
AaIRWxGx769ahTrzAL5RPzQGHI48TUs5MMIshipru10rDg7sGkltm3HxSDglupHD
Hzw5GvM+G2DrU/wioD58kwN8Hmsf+JnsKjGrkRhyuZJ5TLb8uRqFUhZREYL9ogV+
SNdjUgPnCH1I+/X5RjU69DINGd0Dwu/gaqMTej2E2EVuCoqoqc8aaOx/cFyJ3piS
pbnoAEQhXU0kGrY4gSDGpW8zmiXZT9xzMFtfgBH1nm8WV0HrctYyQ+lKijFTkjUW
rj2VrcU9oFbRMoXKRjvUb9S8xj9jp9CFLiRtRJBzQNJ+qEgcJSXS9daOVSbbe5xT
LAXn+MnZ060M8CI4Q5u6my+sufxO7qkfQOMHpzy91ZW++Q4P/qoqhvK0sCr97BSi
SF6NgCGUyWP9s9t3CbfdXsuX/vyExA3ZouhA3KKOgrXR4/iSlg+z99+gY9J+Z3Na
CBKwaA3U/91ved2j/q9DzBY4YbuW0XdhxlNPzpA6ilKCRY5Egc2FjkBPgsGhw4Lf
N+cRWLPeJpkhMg9pOPoftyoTdAITwWXBJkFpUBZJ3BYcm6Vt4+gbeCDPmvkZRmOp
ceRky6nN9cP2YIVtqLl7xNsITBIKDofqnzdiWTjZydrSDTR3VAdYGeG2Qs+ql5jU
CTtv5Nczf42Z3OgN3F1jMmkowVEJnJ/JEz/TF6jD5cZNJOQBtfwT24zJ4Z2yDJZH
fkkdyq2Sm8tlLe0w9j/3Fr8D6ZtTySqI6F/kPw6Lu6K6IZsXZvmMsBdkZMZsOvNB
QBhGv9QxSVJ+2zn8sm2AHuhu/IYC2IYKRHxKY3HsomGMYxYoplvny9sGO/TTsQNr
VvFQRYpbaxRCUPiz3KPWQO1wzuVTNzqPSUEB1+SEujLH/51LbGj442GQZBMq8Tni
z1XITW4Qq/gOI7SW8QSzfrVwfS94eAc3VyylIy1RhfQaMphYuLVleii07KlgIMzJ
5JfHQglata3A2Y9hw8qytb3ezt2OEP69sTSKyalXFU0NDguxSqXxvMW4kZF58CoO
6/dDNhINOKF1ZdJ0cXRUEK3fgRLRlXpbb5pQQrEh9RJM3CshhukLd210058NIHpM
0VlBz1JgENMinBQD6xXpHtgaaZvJxzwvajdo8Eq4Udl6KsW/ZCxWnZ6JO0h3m/ct
JycuY1mmXaA4aD7YioC4Qr4MnQYKUSFn3MHQNTSsFWOvF0HKDC7DxVNqvr7Z+Tio
3YCHk3JbHDERwuq8LE5xsaHyH8IG7su0LTHAuO9dr081iCm/Pe5Oe4CYxhvLtOFj
onIHxzYXZxaLeIgUtB1jK9dV2FKFNeO84+mkIcOaY4NsdGLzp15KL7UkGyj80ZXg
cvaBL0Nv3btqifYWP1kPbHhdbtquBIe+QxOm7ZhSKdMqAKAByuTIGWLFLpAKYSGG
klbcX9WOspQC9BG400IhaK8nvl1JIFtroVm0dFzcgWos6KVLyCglv5M/8L6G2DUi
JFxpeE+6HOS+Xck0JqMTB+H2ivDGYzMHF5Mp4c1+zOx/sRsYFsrhpkyzUmhxLI4d
UcUEMJ+4GUdqZOpXD4foaeKMFF9fgwd/aNGZE5bcu8rhWmfhL9bwQA1/pnaOjD7v
504dCADwQ0rKyPpkXyC5WEaNz4wQyz537tjiB8uATNsAXGwgRc9ecLXECc4l+EiN
TCixv/A1aReCXqfeM0bPDTDMuRH7hEQwKKLXWHGGC9DhQ91vXTkgZhwDSTDYIHtk
xObrT21+pCc/z+MDG/g870EI912puIl42QuYVyfquSh6Z/6JX4ZRubaDdnaoYWEn
wCKYkKE+nNAoP1BbZn/zIz2g9ekgY+zXpDANE++z6HrVp5PexqEw10mx9q6FwO/Q
iRzMOADI0FgQTCOGNgb8w5OCHmveVihD8R5bHelSvUlvf/GzGxXQpOCIBmoDZSKG
5gJy2YEilga3drn8zOtiBgClqoPAPRlZJFi+MdsYZXAlat+m84yGxnZIxCz3K9Gu
J16iJeAHa3BcDWpKo33ifQf1murJE9L5VdCi1DgAGLTpUSy8yf6O4Gh/PPCqruYz
LFl92oGWVV6nj2F/cQ3hguAcxNDSnsa5yaokKZk828WgAd0+XVC0p77vMzBufPjf
ur842CBfjmTvJRV+Ob2jpDHf45FtDakM9l/BTruE8yyrO4BXNS/wnkiGdn0rQekR
/UVjzlK+iFWfT8UqHOW/ClInXoMohDObcAAA5Z0uRLz76ki6VkOTrDiHOPAxxaiJ
c2W0q6+dXRYSvs9kg5mTfeSqwN1VowvUxkYRXkoFb4yZkgSw0p97AeN6Va5dFO5Q
bCfqEUXp7zOXYEVnMEKEv9MAAJuUJJwxDlNhQh0nXkb+uXbT6+2au5bmVIFjpotk
PAN+lcYXbkObDCyH8+7Czao+Q0mTHrdFkS4xrcQQntO6S/q4FWdHhyJbbMeVYQcO
PLhGWyN8gVKX9n93jgflLjTN9MKhU8mV7PlVTWZ1WXCP+QKcz60XtCSAt4pfj6/A
AADlOxx4SE4rvTDkbP1KtWeG2Zrs9eOB8uJ0vOWufvRTIwAKNeRG1F0DHGaVqqWm
aVSyS9g43MF+dFsOL4KoXluurT7IItXjXBZSDj8zVil94apej2+gZvLiva9wz1b/
Ya7vKXafbI76HXA1svZtC6JzXKDuDX9GwYwH95bzAJntYCc75B3uwgzJhJTh6rtG
2PVV4jkQ4Zk3kP7fZw5QIgThAYpj3STOkMzzNY/qCmpjAUvbNZpESZwXUct58APn
EiBhRQ7feUUwzE40X29wT2HAM/1xWKMXMrTRAeYGjX4BpaK4byXi9EJRASn4ufV2
VjvEthwAZqrbnbXn7Zgnop8S8BB1WPiNscGUZNCTgm5nvtJsrbhawKT+w3GKXrnR
HZRdUhvukLdGTtz6aPPNDNsQ8GTyW7ws36WY8+m+gYHOMONR3yMSWhnIcKAWg4Bc
pXlxBm7QRBv/sYGbhJWwdig594agcnrHBnpay+O/0yXExd5GhnsKjeuIhdOUvwWq
km43X+bNV+V+QI4r7lDI5WYteicBc9xBl7lTg6gZJ48FGr4K5fNYK9UC/Oqn9qBB
/N/ATJKLvX9iWqoFmujbriICnSYntWngYFQS2twNyE27c9JYlxivlrz2c4MaePRt
3T4y5HNQG8UPEugOkXBxEHxhGL+GRCIfztrT2tHSY38/3MCOVAtYSV7VKk7sHMzw
oJTg8WeFQ+czkDHCnb9KPHAKYlyaaYOuzuaHAMBzcB0wZP8lA8XNv/xYjI5ahq4I
iYucdoL+W+Ejx4TGCHr6U5jbYsxI5ns8O/tYrwS5gHuCPk0+gUcMzxZR+C2Le8zp
NTPPtlIiuSr1tONxQp3aFSEC+uvWrAyADnUfnRauWf8Xf7tghM9f/EsCRmNaFGMZ
JNwT8+znEErTaWzz1OQzpM/B8oKS5ycQwV8AdGtZad3Z8blHL9pDVyH8KWKuzoBc
WlIzHmz+XzxtOMM/isB2HvbMUIlVhWUGGDANH1bXD97iHZcfjGLnoXIMxyC70Elz
cVVaAL6syYuhBonIgV9GYZFtPu959MsOFHs+g5HSeYa9hXpohtIkIbVS7VqIGsYS
PSGUJDo7L0qacqWM6fl6ExhVLNH6uIk/iHO6+9xPv3zihFzA22rvdkJhHG2wK3rV
JAN027tdp4uB3wkwpdusAbPMCLGW9avKqQWNvSDemWmq/t1J1SGJFdx8ktDWSMyy
yorSSaRsXhlZuJT4VENypeqoWpEvi6V+mMm6CJ7e7CvD+ltEgvEMnJtD67YmndDP
1zuM1crmdulwTy9G9MsUmQmZ/FfFlx/MARmOrEpiKs8tITaazNF8f9Pc4hGskPM5
drPbVWenB4ZQzxvC3QOf9ycGtMd9TqAp8pogwsnzyrMmSOjjxI1eD0YGSWdm2iwS
Zm+uFF1Vo/LdyvoJMXNPGFkmTJq/kjC4ZaMokN5RI4vho+BvsyVTygsvlMxhQO4+
6Y1+ExWvBDVi+6/Me1N0PTnlToVGWSy3/VGRa0OTw8/OJ8V4is2s8xKuWUQx/vVe
D0gEB7Sfh8jAFp4nuqKgArMZ7T2nbhuAJ77fB6ihpgdl19FA6k2G+4pC7nL0A5Bz
CdFhbeL2fEjFJ/Tf/fkJ1JkKHlbs7vJm41qIKk0/yQvUgINdUoSi9UE+jXmv+4pv
2CuVZo8RoHsHzoOV6e27HW7ZffQzm4lOPmSB5/7A27lKNIKr8CJrLhBIaiXcWURk
4ytDOJaq0UQNIiRt2neIt0+A0YKma3mYr9pbcecmKnP4miH/l2wkAVjqG3TtFMsn
k/iMc6+h2SdganxW+QhLgpePtTm/w/vytqhCmnsYaaxyF5joxqLIzJfgB5CftuoA
3R7MM7/BM3sfdqlqzdgJ7B6/1Q/ISNaLJAGTYMAunU1ZCUurqP6ifIX0XQVu8bxa
bws3FWUKrFngxu3uSiTtU3sq1+3gyrg+wf+4vXDLivpY8dx6MIQ50UbJHvgWN+Dh
TAMmNHjAchY3hzK3XK4vpC90MLvr0OpX0GAmBZc2vZU5gI7YXwcRP9ManVuDgh8c
WOVch3ZZ49V++JkP0jTXKMvaiiMXDUxZzwpeU4cSkx+7CWTBXFhD23yfw4jUSJzo
AOHxEFCaTJFBxPXNa5leoS6n1sgrJm1zxNC2vVoYnRC8+/fPmhoVWiEH/FCqrNmb
FIjZMoHAt4x4UcXLRfZtUB7Y3NAWixIAK6EJGQY/I2VSZIzsxaj5DR2YwZRj8gUG
S3wy5wXvEWiV16kyirSmo3F/n2AYdT7He7XsgydHpdf3a+iCEAMmxOF/NzBayZtW
Arm2e7Y775Gieq/4rop7Ox231y9PsslCePTWKAGkkttJtZ010X4Nw2G9JWH5KrFs
AxxcxgMDgKkl0PoWFigeb6b4TneG0XiLwEqLsUXaBxqhh8LYMKHLvl02sq5fE2Yc
2O6gctBF1BXZzEp4O3kwE0brop+xvD4/YYylcbQpqNLHibgC8tJjCaZ8UBcWo77E
tm0n53lXUnGS7pyE5+XOjnm/wTRj5gbs/qvclrOyglsgC1mTVT19HGhPiN0iOYlv
t3CC59C02PkOavtXAtpQciRN2yh0fmxLnBSOPslKqRwIrt6/B75Zfb5s8aRR3gfj
UEgiSYTPjV4omn8MfJAuhnfARVkZV486kYtZb7e1iYNKHY9TtG2zII30YZIByMuV
Fvxz4FBUFNmy6PzcCfNyNa47jPsvmid6miw4qfyx+VSSpl3lm4/k7FA1NnYen+Zk
RRdBEfcKC4Vu4HXVNI5o+Q2PhgnXsbAHI4Qj19gFtfXCTM4y1DPlFlCXqdE6P11B
wAR0TTSMdlHxormoV0xq+1F8GgtrOVeOd82Y7TcWMPZ9n416XsCqzIQdBfzagtk3
k1kVmDprMuHdC8B0UHcvVB9stiQc1ob2RwPSs0S17rMweHhk0oII2nR2kNTI34Zq
AEXiYvIHS7bubagcpVVi83y0kr1p9J6P9EYEJ3QaYo7cUgNHgxRo5ByMXwt6xQAv
ti/3KV5xvRr2g2RA4nUDyM0xVicLNGEdIy1RdOe2QpykU8o2weXApa3oB1UlTScz
TnpeKQ3wDW86W0hfziddSDaBAIbmZHPE4LzNAkiAyVZ9hTT7viEal1WIs4NJ1Mk3
/rgW/wRGowowt3BRGe/Ffz/p0AY1b9RqyjBGVJzmmlG/jhhbCnodDic9oauuh0Eo
AlAycRNH7nEO75C8Ke7vP4Mmigr/kpOw+5Tzslnm+sbH6BdVK1+pOpKd1u4+eJ3x
kvechMD9kL/duq1RdH1i19xPxw58B6hNviQ6NuZOSpeLqRNDaeIFEPG7B+tH9WW/
LLHR+jcrmEImYhGktaxIzJlgPDCVgAveZCnYHYLgHUno8X6cM2bDKDhLmnq2eb4Y
I35AcVKYJSoma010vqWgmGLwi5wtthjVLiDBb3jO2Z4EEywsS6AgBUcjlNQ+CWcJ
jnQnErlZXJCk/8ltuT8qvxtOBCmRWaSJtTAMKLLw2FztIyluN9+b6KMufD6dLzdZ
y5ENiG8oBCsOsVvP2CIupAX2HNIQs332FxZI1xhgf87eN3+2VuX8JBa24bWL6Skh
RuCDGjGCfgwlWAJaFitCOK7fog69Y1RQ3YvHjuns5wJA8r7cWJd3w5UDO4T3WzH6
s/Tywab96z3GpgScFkvhW1EkEJKtOW8azDBFOFKq/mAm0isr/jBHC27RnOzfi80C
LkIgbgPNNf7D2iOvjBcJjY8eQvVN2keybpbmApGtohsDRuvCqQZ/gaNlVvxXNKfg
Wr1Yv0e076FT1AZYUKx4W3Bywp/cc9NeIgylmCsCtXLsGitYQmghoyL3WY1fGNn2
W4khAWcf3lcZhaTPNMpkWv/UBicrZCygpGLy5uP8NIUwHAVZy/TJinvWjLLMv4fF
jxgMP7FvUCCpJp4ApLPzY0LAuReiWQZ8NM+aJ7zD7xmiHhtSf9Qbgc5Q3ir157Jz
t0Ek9rAjvuKJGo3kHMOM9fkSW2dIKdi4Y3JAQLz7mdCM1WjoBv+9OWaX6N9JGUkp
3gBz3ktzeB+pu9+i0/fSEeUSixQD5pJ/dijzINUoPJPAtbESMeWTU14sR9mGQSdx
CANH2XBmtY7/+qIUA+4MonggJiCt1wrJlbG4asNcf6tU0j91rscj5GJ/9MyRiUkX
WE6gFtkx4jyjb5t8uYi4FHulCfTYkeuLr9ctEux1ouUMJ8n8l+g30cxUToGe1k4j
nanJauDRQshSRVxgRM/6UUvzTaOR39r/Q/m9IIamNxH1CNETwX1xXwHwt75ffII9
0nPjyffzt45CRLQcHgXmakJX9s3cMB45LgGD8nrF/On6UtKJ608A7Qm43IcB1TcJ
r19HQjvsqVSQ1NY+B0Ng8Zjl7EBZ5BXfn5njI9TQ8zMXhSCP5uGguVeT/MRx/XQD
A5wAMA6x7Vw50lK3CTlIwRHPXgYACtJNYsq+53/yoB/Q0a6SKQAXlANbNxqWlopY
R9W8J1RWokbVYn3jsHYao8SljTiY+i1/Hoie26O5bnO3ELjHMGbwD+bYVX/fJ5Gn
dsetbw/wy1Wd5ZS6l7z2k+m5nVvyE4vUMqLP7jcGKpXpVIzN0cooC26a1TYTZQMY
hA/XCa0ayb+lJHumCmqqZkTxpbz6LThjdWKF4Br83g9aE0joG6eYVP1BkSgwezzP
LqQEwqsKRjnhGDQjiFiWaV+rvnI6ya+lxxJG3iwEKL8cVzmtJPx0DhdcN8ddtCag
BAI4IdcCYrzgjmih6nlKY6yrc4HbwXfPLIrSZngn7xhb1BUtrbEjC73iqZU4CvqV
gIPJiceywCHATAzgtEpmxbBvQNvs9H2qKBWQ7RBSnX8I5FTnEYkav/IXS60JwSrE
PH7um1EC5uZCoiP2hAcyZrWCWYZJW5X+w6Fw7KZDtO4z9aIPzBCJ4IDwriQYHwGX
Viho+B42+I2U5vgmehaGCr2c3AlPXcI7ek/yOUYcQLCzIorn9sGCUMUFiDp3LQwn
Oqh3Eo54WvfHj4Inc0VGjMbtpau7AYnJCV5lRmRnCegpTGneUbuG208JIPXZ/oZY
2lLuumgWTv3TB+UMvEZBZAn+Ufxyf+lSf8M1uR+H/SRZmHALFZ8Qf92lmEIwPuNK
3lRSonZsI0dc0S/+v9pW6lNbtymjZgm00nZw6O5vSaq11UH0q8GT0UfRxq8MPepH
myl/0GLQgWbzs6n8y5FtC7xb8QATrKbAXccjdEb37QMbQ6/+cH/JOdeRNPCJjpLi
Jprq+BJe0pMLX42itd02eGn9kWp3fOjg5SfFeuHNvYl7otXXKZ+mkzjKKZhbjQr+
tw1Qm7+kAsQ8eRxmq9yeM7BCcoNin0RLghiQbeHY0Igd14gg4nwdYsuabGTsVvqt
NOeWhkWXWmitrm3lbC0VthkudGBn8FGiokDRL/0luUnax9Kuu0rvhc3mm2d8w6Cj
JVBsOskAt/1NsvQBLaIbNLHDdu8tReBZgIG74xVrA3CDvC3bvR2JwCTZx91fRoum
uy0vW7BdXx3dFlYnVDRa84H/5Zt2NAWA16+nGNJDFaFOiv32fGTZTrHIREdP++NZ
zoAsAva+DlJz9JI15jBpzcVEYtNCnsBvxZhfYblF735u/uSoEu1X22nhYMreky3Q
FPBHfFx+usl3x8O1SAP65hmx1+V+xqu+MVwLdFn4X8jPSO7/dW37onXX7WB5FHyF
Qw6ykm5c++36MV+0NkkE40FfEWSPCFkRhQOEI+P2W+I0oe9WwRUcb/ETaEPenROP
DMTrhSH6Z+9WuUbfrSRcbZjAABYqIkfEtWk9+EmPbjBoG2bTLE2JQpxNdvkKQKDv
dKL589H8MMFh5j8h3TUhAXJOcn8RzhVEQxO3oOWMqahJU/0mRBqHJrUod7D9dH0d
coaZdygG89YNq41S1CgMJAm0k41YUhfo17fnfsNX/eftDQnVQ1Yvuqi4+6IKtil/
h9BNvXlot9tKyEZqO1614FkarVak3jjUFd3kbLtuvIeags4uMLVmXCy2WSHcf0HN
nVayBoumt1L29ed80DrHx26zMZbmBD554roGiPbByPcw6DTArZSgpO9FDmGAi2Wc
YpzkjwHW2ie0iDVcYdEzEYEuRB6tCTQiPIrFZeYnmQLA/pX2fAy6uWP0SLyNoqpA
geXiXk4TPJQZFKkC6AtEXR9q6xQq/NoB+OiL/uU5+reytSok+2/HNCwmB8CSkF0s
vQ+Zj9UbNawbuLN2Z2q8vGXJBjy1+Rpy+9MsLN9hd4xs5xXjLhDqm5N2SRO/YwtQ
vWwMF8FOqhKPHkISo8liW/8e28b/aM0YOtjAu0/m5N7+wsvN9mifI7ZQVCTwKZO7
FKBhvEoz0Y8VnM4xJUIVKhxwrKSRe6peQvJ/8/Wa+6TSF+fnoa7kep/7IvYd8CS1
PoB12F79jef6lpNNcCmuyXA+86I+p7LHEu4BGcu7r6zzg6jMIYfQAx+vqgDQm7Gv
Ng0Q6o2qI7X9iZnEY6+m2WHuvVaRiuV1AyxFZEghKug8+Q35LV9LQbDRDAZUYuD1
PhPDd9xLpYsJQwwFZsT7ufxqKZ25mfxdoQlcUfLfhzc2HkthdDGdQXyUg2iyrJ2W
ArXO4PRGBgQvyXAP8W7BESlnvW8kPQn2chpucJktWs3vLR8OAM1fWiuHwXamDuYE
mA96w1awuRsyIW1inwBKdvTr3T2bUlPQgteuNuN4TX3RDZPzfPFSiGay4+01hq26
h8ZaA9twPlLkMn9YJOlJeD6uunuyDDXVaw+6Q9s6s8nJAxSV2LFdfI5fvYa7H0m6
qxWR+s7V+pzs+79B4koyHN080gO4lj25dR/uo7f/fTti5tNw7+LCKBOScAEMsKij
EIS9fv4k5Jp4577KSbDk4CW6nqNrKpEWCWe5tMhkI/zY/JETvG1O8RoEor9Y1HjO
8ikdjraMajKnAmK9+ZEJw6kbhHO+GsgDY8SowhJZVyf0Zd6aQAaqEWZvrANieix6
3faQPyRpHuRw4WPdxG/yF8zznyb6ZTcbKIjwGFU41IOUGMGdK6qupgSLEetrzEH4
H/E+vl7anCJvuwR/NLyjlniOvfiLdgPZ3D+NNDVJkkWYIuNwL5EhOLeq0rn9HN78
2wXVNArRd7numLsfyWrYmGbpIWYUE7KQURvyGe5gX2lsFaB5KcMbMsr3o0nYG8IY
8i2ZxTb34XaZIP+xRPqjJ/wsq31H7des+f3N6/9awjy4ON2iZ+qUx9gZUd+gyvvH
9HLAsOGKMFdrE3g8QZE6/elXBRyUO45wcOCPDfBYI3UbAvLT30YTNm3Oc8UQ3Myr
irUeIafiGw+IY+q4xzZIPSSGPL1HKoRo8RVWcVCZz3iz/9o5BIx+JuGpyPzSNWPC
yYesmRu7K7HIQ9cEHpyB7SKxTVZ7mwVqKjb+OQ5NEntplSRJ0BV5iq9YDtdyGXOv
OSNolfCyD+viTEz99DxKT9WgA93cY8s0hQiN/aHAnBG8PD8HvTAtX0z0T5G/ibzd
Lx9Iblea+qV6dDESS14fMuLEjYumi/zfU8ikz/KY7tbZjdlEDlw15ZIeg+t9K9dO
30+v+2icc8TY1A5E3EUQoQAo9EltBr+MZxweU+5dcFb3NMZtIVa+vzWgwoiS+3si
nRJtCZ+4+3kuOAOM4wDImQuavr//9eiNUlr7lW3pi4ukfDnnMW831T1qIgpwaP6H
Ov2w0CyW5PYyc9XF+RcQ0mhmGL+JCDYG8SFGat/C2FASbiMfM+0f3AhFL5Ujxx50
mJmg4vTfJXIW7aTpEgui0s553YOTOyozkVPWnGbPQmRbM7gCGdengrFS90xv4TRq
zgrnucys4n88dTFMRiPDx8rZS/uKJb/w6Sv/Q2CJEjIwm4SsYEfhvT7nXLqtI8QG
z7QeTrL4iyw33SOtE6G2ABZbgvd5Sec6vUVAoPfa5LMCzjbLI/nevtofh5554Z+k
DHuYfHrVZRHA0OdNz78hPa7sZz3Yvv7rmAVb9V/wGl4Dy74QUn7HPSPDpyZHussb
5f6cDRJ1At0WTa9ChBFvZUz3uy0TEVzZUNyn/BuLrw1lYJLVeLNzHOykkKuZGQaF
5DoEEsA3jRHkTJ4CaBWMisLV8rhcM1oENFq9SlU620p4CMcj93bsljB4xeA80B4o
kXSP80JugT9jP6SdRKeW7AvOs1C4dOuyq2uVkPiJttU/8WkDQctbM/oKv+xTujE4
6/3P6rTuW8AyDr26TLoU2pKgtdLVJS14ClRRjJPDT2re5pL1TvvqhbhqWFi3//g7
Uf9ctotw6UpdQSHoe2VYDy9j1mB0bBPGlB9VSn0d5mhV6Cm3+aRqfH8IUegJ+VoH
fy94UOVtIgpztlVgzxzzw6cDY819627V59e/70Za3WYi8KE8SHEApdCpx27MjKmo
Ns5lcVhmhYp5jAyHmL1+KD3x0N2SArCHYcgoxYyvpmgX7Piw94PXlAxWUB/69Cve
EaGwX8JyFOLWYykN3YIPhUdIgRUDlvjYD1uXUfTqwr2AApUPRAjuYQSisqx47XSp
3OhXANO3AUd7UAHWZhcHAh/ra6g9q46bCZDkrB4ARFKfn7s1CIzXESrQA9MhFe7W
eXXj7Rfg7gbDa11QIDPsLCOuSf29o+nSl6N7u7Dv4jzKWgxcrCu+30kZNNEZbi2r
cQrKEuzPlPbCS0hJ0pAcUKGu4SmPjXjlq2S48mWYeA4GkLpKHunwx8ThdYsMtq4U
fNU1WU2oOXeNhHrP9Xwwhdw8qWLopDrOVF7ShU4695i/eTJk4FvL9uzXfEjv7bS7
TOoOTidndYyFyFYWU8GS60P4O2OtPBGu8X0JkMEGht2h95ffif1ibGvxoOmSVL7D
FUgBbL22JRalY4MMxXsXytFdoUIg0WsLgFoTy8PuKGrFMOOpXNqZT2QZfaehBT+O
ATB9JrpKclu5ulFqpz86Mkz6WfW0cYeUhNy9PX4lUQXj1E8qFoX++n8+3CX5W/fM
w/8YSeUxvj3PGQo123XRyZfBKy0Vp4J9ED53GkAVnl8M7mYuAk1/nXGEG6IXzlFH
O0GNeWUPpEl0DdpKQMLeJwRheT6FNR0F7QaJkBF9yVldoy3ocjcu3TDHhzn2ZkbU
eNcAxDI2E5AHMXryjh2zdt7Yy2cJmZlxh0cJmvJ2FFT+2djb3lJsZN45u2C+ZNmp
vsf31Gg9sQq+z1qrHyDMk01fcEGeY0jvv4c0Br57BHEa8QXDQfN+P9i+lrsDsN2a
DM0KHdy2kVNkDWj6DH76fqosg7pWL1x4KOA2ypbyhuBrh0KJQBl+7nO7O0tILQwA
89r2hE1LdpMoEQMITVWkTdrAGoU+fIWevsNBfnI4SdJwFg5hbZEW2GM3d7VfIWE8
R2eLa3QLvDPmiSVc++22jHZXHUaz6yB1GdlimDdqGDMWeARofQ6DIDGjnLWS0j6n
2QUDlcx+H+z1E/TE+YkspQqPpWssRE8LDoaG3olLaqOuHRIVzzPP/WogXdOfZo/P
b6vxZDlPc6GpFw1koXNyWqPup7nw76NDm4SRULrgQZTF/IDNv8ShbYq7QN/41VXt
qaGAwka8kqprmzBbi80Rgmk01HPd0ncRfialtOlvUfhL3Qkbft7XDlBsDsA/q59p
U8skH7rOLCLnRm4h1OWgRsYXszaMy0qsCAsYhZ1izglGBoXjfn8t/iw6mQYSJO4O
Wk83rHzgnTMhzyJFkx4/y908FCiC4aat3M6mOc8sN4sQ3/nngsZ6wtIv6e0KRz7F
0Hmzjb96CK47dN/9D3rLkhHqYr7f/IVNmIxk55syj9Hibpi1FA32akut83bz2Bnt
0GR7sXvqxxM0FKxCh4yEvm0xJBPn0xAVWVevOrvpZRXmkFHN5yCJn2+fEISwgfAr
aGDhMAsJ7TepGaYnEheX1PboYEKmCPJgI4U0CF4Uo6Fb6zt482jbbRWasHop5Q5l
5cySQJ1ruUPUdSeczIRc3ZyBbc1jcKAG0y7EMGubo9YVZpgLjVDuJ+mlSfoGnkWx
IoaZrmd2t2U/4lQPZ1IdODcQnVo3OghjiC/EbPYLPJ4AZKVJxQz1nZQnqR/dZwdq
M8Y5geEA5uthZ5odjN5QPM7Zhs5kcvX9Slct7bm0ftys9Pmaix43C+9ftlDfU+Tu
d/OdLO3AVoUNvZYjjxukH4DMwfHxXLq/ekzIoeM69LwJ5unDmT2nSXrRRXIDLJaK
MaofaB43gkr4YGn2vN18MGRoiUoaSWt+m1wlMfoQ/XYL0IRJxvU1tTbGxrR2LrBZ
6n3WdHv+hsXMWY4DgaJS9GWko1fAU1uEnATKeeBlDtkK+GqeA2eoJiKY8XU9nVbK
uzYEz80khhahfjRE+twQx/HOZDXyjPzIg+DJ3mDIDTQun4WV9bq1inl2Cm0LNk8N
yCacz2EPfyLfSj0uuhAPSIKpJv0JXLXiqzgpbg0bwXcoT888Qs0MV3H5RWVO6TEs
e3ZElXx8XLiTyAVlN73v+NchAbc1YBhpoOdS+BqYim0Fc2GaF/FPKdOfYBpNAFcg
gAlTK37dCzx/WnOwSv0hRCW7VxKL0dFQ+CGP7v1To3Rn438JnrXyypcyVDHGka/s
+ET1Pk8+WJP2EjnpqAK3Eocy9XoygDKJP3m86sK9sUWtTj/eg8jMLVw+OjsC8UV1
kvGILmhTVyCPwWetHkxSFt9pvQhwliiwvzSy/AK6A3HTuvsBekc4A7f/hFhoY5Fq
c6iwligYzr7WWon/ZOb6WWygnImD6JLat+RXGci5ofS4ixVjwLwt+yoBG6CAGaVx
LO6svlQF4ts3sEbxwht7kEn2ckbyGerucw07YHl460n1foIAreiZsC8MUJjq2nVu
NoFF4L3KFWUr2aOlXQMYrOknshbdVOYBKgHEm4dNcihM1ztj2PDisOiMyg2+7z90
c+dYrDmNCNHq6w6IJayVW9yuuOdUgjCvXJY9xeAVTuRNp2Y2CY4aesRBg/jO9313
2DThxhTjQ1t+mcdczO0hy9x+OHELTuQbCOyCrXX7WqsCIXnL2zqbGyIStdXtUTRO
lBVi/Jqo8i20AIdLWWKWYkB53kHc0CbyHu1k4VrItQs1zMYGladnJkvvE50uDjJ9
UwQRAQj/7bTVgIB0seqk6GeiBTt2gIRPAZgjHcVf9r/Xa+HQi2s6NoOqAzZLUijd
ibJ61HsVkIStBffSuGpg26G1EklVmtZk4ME8+9TR11KXHn5y78cqjGnydA7Lw1mB
DnSFD57meMYco3/00D7uAEMTfquC8JFbgjUaGf8edXjm+6RhJ0OEG8f8m1uaVMa4
MopZj0/Up4df2IUdpGh8u/n3B2wJD6rQelu3UagKBz13vx+qI1Es+mO9ZE6rq7yT
LhHgHEBObXDMVhgU+cOnuZlPafXzpvdlxblHTv9bbYX2JmivcaGisyzBDKrfS8gw
iDdMsbQk77Pyk7uTdFnMxent+yLPK6/97R/XgY5zul3hR6snN+qN30fxJ8/kqeN8
0aGMyRK2CUnKKIDRfNBgpbTFyQX9GM5meOOsMgyy0kfTB8JL17kEM9L2DTAGgkTX
gzjelGh2Hpg8dM/4jLC2oG/B5OBr/n/yb0ea9/xphllm/QB++lsE/1u0Cq8eGcJx
9ndNrw/UfXrughFYZKrmbpZ5/HeWKP7R2WJ97G0wUHnMcw/W22pje5iyKta0IGD7
FE5k1SJ9jminQK2I9wzwy/71kbmvH7nImVAX/pnDszVoQQp8WvOArdK8Q5nGS6Wv
RSLrgNMokIpZ6UkDdZkflIJqq7QLZb2myLl1qr/3taZEEctiBlypk1jFy3cy35ul
X7JKC5CQDuLpL3gZwWGLVQqTjVYmgLWyxRLbe6eYKtL9RWE9EAD7APvYOBi3oM9C
RLxzN89u28faJrnCYcjGKdQDmja3bwrtlpJxXUGZbaNNKWVNOwgp2snHEeo+uJ3+
+aeSr2HlkRlVCHajDGA8faE9cziYgKOW99CMUu6UmGH6iX0Yx37bBIY0AgXUWnC9
4BjbBHRKc2hYaCEgla+9StUXzfGr9Sm1wdLQO/mzOJf413TXmCWefrdyjtJiUNM3
5gKi9o6eOrIQlq+I75TwwqE4xlVSep62XaF1GfIh8oOZogO54NrgjH968ytgNvLq
TOP6etHqVrhtAv8ekZsgKKBnpeA1DqJDtizj/vmhwU6bG4m2UZhHdMDoruhvOd0F
4EOIv7MFlkAA6cP418SVoBxJq+XZuD+nDtmOesJE+BSuqdmJQ/g52F1B4mw3vFkq
ESlMSl96QCkNt9XeHwnESM/khwCxjcNs4aTGtYNYUkg9JaIqFK6IvIqb9tJ/AQeB
deElxukjNoeNeOvk1ee7b8DhgMiXujfN6x5cqXb0UPMdeSDLnjAm8JG760V5e0Mg
EDItHYyx5Y91dtOgCy+ZwQj81iPrVtjBSgPqmcRy8QchUNtEe0e3O1D87s5Zv/wU
WlQ1lg4lJ/ERsvRRQq0QZM5vP45pb3tyn/cBiXaVaH4WQW4005r8Db71JmYRgMOD
MWxyN06FIAoa5+ZE7MgSfT1RjqgpOfGCaeffCwGKCm8x+IsfuYiz3O2jOp9vX4OK
nZ4U6C5nc0XgiKgymrp5vwmR0+5N7acrXlRo1Ks2i6wDktE8MyKzNYjAck2vjBJ1
dcheu6asIHUvD47gbM+bJHnW2bwC2EjtGsc0uvqI5QX+0VBDbrjD6CwBHSzUOdsr
6eBgNPJcdlMfqzOXkpxL/r64ZmUcDg/8i+oRYHEgrcfaP54ZTeMj62AkPwlXk/2H
EhjqI8rQ0fyLE+HY5g3Pu7nPk8a/7m+26GCNX7usn6aHPKRyJKsc8eko/zSTS9PM
hhr6KxLvKmFev4ef1GGRrmr0a4xh2AFgJW+fcISPcfz6J1GrrBIVLS96wkZxBOTj
bvFudkDZk7g/ctZ4Em9qczIH4nqJ5DEyvJOIcMK6A+AlsxkVvrW4beCevC62qw5k
MPws+Iq3gki4B6MLUXm3VmiuyUdLeBY+E3EGmI0PFXfHDuIY6+6T2LJoobI4QwEi
DdmT7+CPwLr7/Jm1mUfflGGbTN90Ld0eY+ypL3dqwR0cPmLLIOiyV3E73HXVd/Nl
kRwESkVpIqpTODclL214aSFK80X+yKTTeOV3QBkQ5WG7XD4+M+j2r1Gv76UE26M8
SecXQsTZI804lDNClR+3rqOBwOJy3xUzaoflMfJ+HFQWG49X2B62gl2Xrn6XxBgR
e2JOol29j3lRkYWbeDLDe3KuWSY5aetgf/SXrYVArCPZYSqaaVSk1zZCxPwjM2p9
MugvZmFMtoLdpJYFBQLD4YtB2BKq4Y4Gl4FUdrqO7q4nZqTYvG+ae/fapYdm0nY1
lSOD0+tp9DrJyUSGq42lOv1FQVdbai9o878YWqsd6wOkzIwINCIEoCo+GVLjkTbs
xOl5w33byyDE6cl10xbUwSXS25Cytb5ZkX7gqQUJoJwHie6vm8t1M1K5u6nPdpew
KVAWAb7B2Jmghq0mxU4lt27rYYHIQUZYElkdzr50vKdyROceEzViK6r7yduvQpqS
T4VP/S8Ma7wY1z3sP+GQ3Ilog4DrJwCsC2HCfflwSqmivMfu0EWIBTkz+c7WDuXx
0gZCL0+G4hLDVYx8lkDjvzTnVwR8ngITdB9k7upOJdrPz7V9IhnK3CwI3D1TIqGu
EfKOqzEMW1HLgaA6jYaR7FbWMTx4vLfgm9+n9PIboyR3usRVlXc7LtlJDEZIdQcA
OxfQ0VXwlUOgDJ1BKKuoxBgMHTw91ay0omGOkWB+AZ77lOAnEc0SpvSiOw1VSmc8
PhLxdL0YPSoO1btx+TTqol6NYNqWxUBFvxZrls+XjorR9rBLLiNXdY30pU0hbcYE
h0JdOR9XlSCz3CbEbqDDu0Xa1QJC865qexUXdx33IZ/4qjGeQeGzFnHYYmZLWPJJ
7pF7mMzOd0Y8LHEQ0z5efsoH7loGU0ZKSiwQiXPXk29ZRTaEsmKJ4qankQVhxG8X
SUPzldCWf+yOk9+mDublNZ6/deggo0FLQ8AaF/6w14nWzcJWT64566nG4kErenMg
Dhes705GKDg9b+ZWB1UGVbte0JvD/gHSn9p09N+YPFHoH5+4MznIRTE7rwGqUpna
ECnByv17R9rZ/QVkDDgMfCgCPp/G/PB5MzYpaA5yJOVhBqqM4FLF0kD+nTZfuzJ0
olQ844zH0yOW8u1k2bK143CFas51Zva+Y9NJcFNSHP5xnhu8QLj3shkioKIbDjZY
7krQxAp9U5ClmexGVYC8lYLFDR3Id93rJRODcVVAW0/zTtW9448+krzux1qAy58n
HyGLnxNYixGmaVNh6KGX+HXQA5BapSf9To10U+wlbaF5kZqb0lU6YapVBJPVZCCH
L2Vfq0hOtf6iEl8K3D/LWi0qFmBc4oHz/LNyn5CkAcIyojSIGrCV45WcW3ZnI0TF
fQ3CiS8ItJZZedLWroy57b3uK1YHPfdEdh1O87mepN6vnJ5Qp2MkHmPvl87QthrA
biaji/WddK4l2mibjVnxZ+gyEurzOgkGr1De8lUJaOV6MlUUpfNYGN3sQFTS4xTd
CGWrta5lqkjeiYPJNaDLhk2AgAZoJW2ZP6yBP+fRpZUBllejy9jX580ZoRucY7Pj
3NC5CmPpCj+Pzdco0hMYsAJ2DYN23r2MpHr40+7S++RvaftrmbH1jXu7VCeB6A64
NI9Hd0TRB1FqxlJLu4DJMz9R8A1slsy8j1Li1glnXaFWXBtj1b5ENptyNyvZZvj5
t/JOQeIMSOFYGVlC7W+DVyV9Ak5ErE0DxnOjzzCMw9T0I4M7L9iIwC+K04N3ivAM
447lVtEDOpIKRnuUxlwE0oDHdMr1i3hUXgoY1ZKC7GrZqEOCND+QLRyeKg98j/zo
a72cg2J5pwSdqR4oh1vLeyjrHCvYH8naEbcOzsiL7GvDPd5nKq/ahtXHV6b2URNq
THPWrsSUj4SVWqTwpXJSItOUxv7FXIE0SZxVv3gZ+rY2YHIy8fgxi/els4wsKQxm
YH1dsHpzIZBnpaO50QKYn1mA5nbnXwgk7QwdBnRJECE1gZQG44OkM/7pYT82EiuT
Ivrdd0xR+lMuc//yKtBePuEiuRVE62MPpn9LOuUzZo0yL4sfwK8dXYO+vemJ9/cR
rEDrKfnCus0b7duIfWESWgZu+iXd0RS/sGMPxRw1cYfkMSAzuU7j9R4JBqlcOcGp
WRM4+yy4BdyB39i+7JLwq3Dz+wJ1cOLJmUowgHURmeFZxJvapyXHJQj+GHjnhfow
ENFCdn+7OpZIgtQcTJl9vKlGEWP69OdCEz0px7EEg1rCLUmepg4nJev3vy42Umfb
C0ILAptSZYyliPSApIDdS8PDEiAiEujbXEApeZIjsCh90BFBzbOzxEbSI9rRB/QN
tIxpdyaqcH4gzj42HOSWlJ0o4Ov8JwCG0DsDZu35OHpZYAtC7Gpyy54jwdRuLK/E
55qZVVGxeAgJqKj65PvjT6aImwe5hjSVNBqUM2Hs+GHv5aXS+YtcwCuxwmBecr78
GxRPJHR97J+CrL+MuEbCS0fJRPd3BQL0PLsdzMvDh1QGTUDj/bpzvMwW6HcaeLkW
Bv7BjDKZLDAn5SsawkbNN9NuvXhbnpa9D+szaA99Mq7rEnH8Qbb72iEMG3uJMcgi
6DzCZt+DhigidlwvdZ+CALPbo0G/vPjLJ9mef3pNpN4QWPeyP4NNImTppsuS/3dP
iKCKF+6AuZODlytoMBh9w2q3mvK3EuyGXZunP8hfmVCSh9Kfm08RZnYThrc2HrkI
I3yy3wYlBimOv+UdNM058ovU1a9FqgWPc20zBQTpv7vlJlmRLP5s7XE8HlarVfgM
qy7VfyoICg6Xb5kyTDc5WCqRhs3me+sVxVVMXY/4+8Y5LKZSHqum4DUHhcoghfzO
9lIpPBfrJDjrWXeUPFQrlgn0BBMdBlDPaM7ANb0F+w6GQ5WJTLxfDLzaxfZ+CpDx
PYcjaNlUtSOnk+UuW5tUqmz6ikCeTA8T9SUdULlsam1uTx9SEfpQT/86uUaMREsg
QF7w4B6BeEra8Zg/n+z6h27MNmOYwr9kS8+rl+lhlz/qS6phpWrxchm8gzutt/4L
fYOY40RzGc59Bx8Dp1Daoi2I87XJptAruQ9IToT9GUBfgkSub/5JCq/5s4mcUlrk
8X4c8vM51Kvd3vLw/IMt2/RcO20+d8tH1+VgpA4otcUUe+qziutt3bN0FUQfVi1l
l90vLTNdJdEhKUEhLRpUq6oSgWUaiSLD5rXAUlm2qh7LXTDpF8n9R/SAiylKaYvG
2lRSYUIppcn9+A2YOsUL+KWL2XYeoSc2gMc0a4TaGV3ulq0f6xJc5qxUUFV68D6v
BLZrx5ogM8wcOikJybAN6+YsyDahcmeVyj+bzehPSOzMKwIi5DhTx4Iul4clTKaS
ckDruBueyZQls8Svbn036tPa4GT2Z2fRxNS3E0iql0B62GW3+B7xpwvv/xfERrUJ
BzVcb6r90Ms4ltfmz7MhswuVbnWd6lHjKZEkIriENHXT54wVsbRDNIo6XUH/FZNF
+Wq+Pgrir+7lGvlEDaxRpWet9D6UgHW1P3625auIP8UAdcXEdGNTNZCFp/J3xlz9
N7dCEkUT8lhRfX32YY1k0G1lkV3GTy2MR4HEmWUtdslUTcakcZTUMPPW/gwVKjxH
dBSFc92EZrYi6NoOeJDx+Eml4ShV3OmaRKP6JVj5BOrMY066nzaIS9EspFbwBJhM
jKx3iU7VuWWUF9WOI+aMjwEPLaLwq8CmUgrfBvoJoTvTqXhROxUphyR42JUA8H1R
raEXGT26MCa5EiR0x+aD2AJoXR7hdMcjU77CQacGJqBFY8Xz7km/0Cigw1fVIM2o
MuP8KnLajNPr3veKqA30mVYK0FXUtf4woCtntIj03PWSTC+7rBBGGaJWXzudPoID
3cpDt7ubSqjDAjltjy6Xm1VISB4h/8vlGDJ0NxOMY25alsQGEInekByKKyKYvo1J
jt57IprPoeLHFHgHJenRFVklQh5CHlnmdQypgdf1hng96lW6I+cEWg6R5mmA7czK
OSDTVPNHezKAGsyfA1txjrNPaPtjlieHwvA/AcsxEBy4v21eorwsVCi0PEwWZ+Z2
ckuTn7pWN8lwc6v2vpsolfP3xfcEe6LRGA9VLEorxdYcDWesooyRhm4AxW5SGrsl
sgjj7pZBgoUEeMqTBwshhkRfrbW/zdcj9RBk/Z5bu03G0uTc/+5ldHAvHPupUcDM
/o1gCQoB+UQbneoavH/sgcDZfb4L03FwUqpse0b9D2DcJLejwiB/wBm1ctqP+6lx
jHu1YreaKvt3ZRhBNdM3Gt3ED8UW7R/nwx2ViHvudmZz1/u4WIkzhDDAMsRRLzQb
svypbKwsOS8g6HZ0Yr5Vo8FJ+YVDCVxazz1Ld0uy0I67fFple//kQoFJewr+nsOE
RvYMTs2qiBwmV4nb7BCY7S9TFb02cJ66RBhgBTcvcsfYjigcHAFM6XjwlBN9+m5n
mJRxh9tdi2nTp9nTSoWbH2xeCLr67Z+xgyKBqe06h8+1eqKqfKm8Zaij+WqtlZnW
cq4Sow8T6PGeD0TQQXBWAn3/ScKdUP1UB8qkJTE7RCL2RMn3OrYr/sXHN+9ZlK4W
QS6SQfv0lDHuENcy1DfVX/2ATJ1b+rNZj/Qn7scbyiokW7Kxz+JKBptB4BpyhruW
d9XB5Bsp8XPa1Ok9u/sRg9OBkDs8H5OGmod4hKCGMJeM4evP/khrd9R2kt3ymb8O
t4dWsrxdGBCsEx2DYoZMniNaqIXXfSRbW4bIlT8rJ4vQreI+1NOpPwZrDzuGhJwW
afvcFZHpcyCWGCle+Vcojtaz78Ok4h9SaHhHjCplNcGG873HYIuPdlUZdAKZ6JED
bzAXgm1rPwBquLWXNyAat4Dl3GDYtXkW4KFbWHzLCrW4c5bhhgfFHemiIyvaDl6o
i+hvi6Ndk7x5dcWD+SumixN+9FzWwOZJgjUZa099tZgXpy0dm04iJhMrw+ZxFmlw
NcSL3C0t2NbOAxbM6DJnVl4yxRbZnhXWvaSHXxb5q9wHIf1guYFY32I+5gxG5koi
vtmqmTC0qnjuzfIoHW75m15RkT8CNcSMCqjjOMlI1DSyfZNi+wgCe3RiXxVV5+sV
dbTrJRluULYQfVmdmjrSsC2w1CxUZalD1MsgRYIpD+NnC5jhLum/hb1AiiQ5coft
PNsvE6Aa0p0F2rro6SmGuNJQJo4NxxqhDV+bCg8sCQTNARXgUSk05uQVWINfeMEd
1EM4aUXUkb/+8h/eULbOw7+IJl5SmvdUlxMGD5Y/0zrZOJg5R+qCplcJcuzKZIKS
c1M0KiDtgRmyJYp51khCETAAjH+qZWbHYPzdNX2RirD63NON1AxsIvpwz5pTRU1t
f0PSc+oe2XxoCJIe1m4NfZN6yJZys7r8yCBd0+YgL0n1mKJVgdNBOrgGe7jYTIF0
2hkigY+HlCrrzQaRJ/Wb+PW8I+xABOpRa6ADwPVLBfth1/skfp55FarGdArWfZGV
VqlrXaI7t+uyWm/TqRDS4IB94j+JC1Z487IYTtJZXzLtw9+RxnjwPXn1ot2Xotsy
nW98tfucDSFFgcexURUIVA1y6Bpj0w83v1VHAh1Q+h7RsEVns/GfbK3SBFdOM1v3
ssQEtMLL+36NSbJh31QrvU73O9XhABnbd/zE8kl1gK8lHxkA/kT5xUcGb+W6UgEU
lTSzHddmAOMy4vXh7FVBkU/D0+/ci36kNcSce37g+Du9ZzAJuTePBRDlZ5oS8eaW
uR3p1VFHoEFZruyo22zB5c5EJF4WTXrqLHEkABtKpTeO46oqRfGoj6rG7dZ1QR8L
zZ8gXD1h444N3KAs0t1CUzoQcm6uqCbqAV5KlVv1n9a53x0r3swNDOuxappbV12D
HdVvMbCZEo8cSwSf7cJUKm2Io7+VY5FqK/LiZUB66voLxgI7SPwxEUvL0qaYazSQ
MvoeAuAEmsY+6W/ywo82lzFhMRLIHxc/ssjXYoSpvwSjhApJUouK1KFpPzACXXpp
eMsEdVPI8yLCiLUEft3gQSQ7Y0l/WCeLiZU1WogAYeDL1BWN6GNMCKvq4+AVsMFj
f6I4BZfgdM5mFOmI/4PUsrms0BhcSPf2xL1wDfoyyDhanqEbwm2wfMjlADjYBBdw
OTfOjG0MwrcQniGm63L0XAQ6t3b715xVNlkMz9DSbJ+vXwG9p/Xv9GPqio7yB+pP
5i3l+3mpCM/9etb6YhwxLi/nmXwA7Qx/rHjhA7MLQBBCf5YQqaQOxiOmrhZEMMRE
H1WElhiVVa6Yp/IDtkwdRFUQlMjAnDpjQCVXiZhp7NnFMdAFwkSTDaiGCmUN9e2E
3/J1NYV6KD7nwmnBY9N8fQdPTWkp/YodXGb1CkyZF9nod2S2BTuByHrA8sP7MHAl
ayr4BBLHt04RroQ3BAoavDE7wYmVGnCyweqw2bUm7q7j+47qKNMSMHFyczQcWogS
xi6DUElFYfPIw1ozzAfahaHdnuhXEx4pJw2H5C9dZwRkPmMlhlH7I3CyPxQrOwKM
HaTXoINehFW/Y8DHOw6yQsnL4ycYQQR+9tgGSRVNhZ458mpXevie6dYkxxcztPk1
RPIAyXIEkXnVF9rTl6/ZE4G61sMKPJsLKIaWyFPtNsyftLCKe/N3eBzrBwbDibAB
4QS/EzBLFH7Ua8YIwFhJApi7GpOyl9Yw602grPvv5pn6lMC7oE5pI5vGz9eHKbd/
OVapUsyYOHCe3AHyPQnTi9Jcb3QIj55dn1xQ8HK61Ph6bBHxHKQWttDMUAtzk5lh
y5JO8+CEhDrEtirwUtHgXoXURWisjVTdpwYx9wyreheRVrgPHlAu0Ilj5A/UHqTu
d1x8A+2NNLL/CzyY1nulE6v3ug3cwQrdU8depSYISRaGasOe6x2iWHbQdh8a3JWC
tWn+XBJCziBtb/Q4BTmgNKOAzA062RD76dOBiTPzeeo/Y0U8kWunoIvLsrO53OmY
Cub5wvT7YnyFUF0Sd4hWF8Cbac/jZybkhNhn3YJD8lvicj3dk86s4jY7baQ+SFjA
TrsaXvnYO8eSQejb/DcHIJE/t9kkEFzqAJktLP6z2l6pC/vAzSIqyE2YmcZ1LV1P
WARSe4EgFijubN58FrmKULc6gNhTg+8SnVm6akz4RzCrxfZJQLhDw/+6hIgYRrWX
c9ookRmZ/bsJdOhf/DeVBbF844urw1iZd/fblMnQ6QgpYjMuRLszDJL/CArtRjJE
Sllz74My+J8O/yUaJUkU1dx1UzmZTiOlN0qTwo0B5IOR3++WFl2sx7Q2HFoctgXi
pmkUHmhhyV0rFNBL+/qm8RiaqcqDf9Ey4y36mNSjbYSMUyEp5UQLvMbKrgIdjYIH
w8BDDUZfCTju8paxrKfOKuNG9tuLMWdD8KEYmw3KNIVPwntOpouOsypeV18iLMj/
M0MX7G/ddEejyqMJcOS2zbP9X8ZDt1SuFgaR9OLFbsoKhXvd7nZ0eYo+BpMKnNSv
g+sjK/i87F74ayu6h9zeXQjbSQcxiHRgDOC9Dbvc4L2kop1MPMPI59DTOSmwwGKh
owWkqLXZdOJyK1wdTvjAiTprb9FswsanzfgM9KAUQGTWuH5M5sTlqz51QXQt9OM5
Km89iqb6frwgw4H/YwHidg+xNa/auEQjEzS5SQC2s/XyCIgezahIIx4JHQB/BsMO
Yhjouf8Vx3z1bZWuJ79qHs1oux5bMRrzpAcNCEpqQPv2Wg6rXy/g7UIrLOABTazr
qembXsfoPXs/uG33gHLUAoFGWl8NaXk3hcfi5Dz9GPWUAHJS0PxWZZCZx7o6PxZf
RRb5eP/mvfBC3mx3LpQtwxvSkOCSyH7+iEIdsU4bcNfcHzlu8CxCam6srvA/jRey
+S9BQ9vh42V1tzGnUMLmZONx4oQB6CX32vEILuMZ3HCMTP1pZ9FVCkoQ0XvgZvjk
2ElvpUqT4QONrgerk2qq7IInUaVlDYAyhQkg9Tk3Z29CRWsdHFFHC4cIlUwP+VPd
IKBPqm9PM6jnjjaf4/dWBvIiZCPi0rJn+oFQYDyDOh+3ns3CAvj2NOB9Y12bVTuP
Llp2WNW0inkB3UjRgkaubXeD74D7WiUypvRVoaX+0Zy0nWDaEmK9SiVJla5mdWKp
cJL227llMWrLciVvwvfykveevjKECwvH/TBzartaBkH7FzqatHSffgTxD7AmhY94
oRVp7j7iDzh5s85L20tepszqSjMuKYx1X359d9rQCRxmiCPfW/lLxUx4cgi55L+M
ynDsWXo8YH4ilXIeQFBrgF6jf0C1dMudzCjweBAVd4PI15bcOzxWz0PuW1hvK+2U
Rz0psTZf95RPvm5Ay+Up0XDi8ZFwx/T0VXm6bFhlS+igartStjQaQyPQZ30qJ6U7
D5YA8bfqbu8y8JykiwObIgPuSLgN63YHPAF3XXTD+R0xZvShNRLU750paa5D5g0Q
maR9mZjD59BZIf275g+8QMExL/ThE3m+eXwkk9HpBth/XKBrwvZhdUAoXv2ixOfl
wJmsG272eAiganSiYYPwhw4wSUkIeFhh7yhBOMUbOuCYegeBTu28yqyd2509WalH
irzPWWoKqMqkLUhdI8vZOJEHTG4A5i6MuZmR6dun06ePa32Ej1tq2k5wUQPynqM1
4sZ1fNe+Ke2oQGm7LRhfOTlscegtEKN3ON1w6cZgXB8aDGD2R6/z8E0e44/tHcyv
aMMBuIFuYhpSU5pa8pdpW+0IrANMD5Zb3kPvww61G1DQ2ENnMTgz5eUuwyscPSy3
mNSmt/+0IZCY6UgTcaMoMtCbbRMnwGstQYZGoVV0ccOgGDWRSMLiZH26GSkw3GzX
YmAkk5enAAw+hzmAkIYnvTLoeJznN2ecToOfGQWO/YubBZl50AtnavYhUKNVuog+
qlN8sFvTch43I9kBSx+0yBG55OM5McP5nNl0Epu2wjhCjDoHpheJ0lUvMvNgGDYD
5U37yQN3xsm0zPnh9ZghXs5EfJ5zZHtvPr1nZ2RTbJEGNxXUHa+XzlWtdK4fN9VY
gC1ekRZkJcfyOpqfQolQ9OYDjOJ8p8OcyMHhz29AeMut8f2wq1TkbDj+B2tnKifw
QGss6uC6Oo0WPHt4Rs/wvsMtUXm2exOznyKPFqG+4hFGyFYofFoEXH5IE9SgpcSw
06ZDIFOLb4xBySBaETXBrMyXQRutIkFl4n330hqy/ggHZgqaYtqD9XaS+X38VQvW
7c2CHWbL6ZdFLAP37yN31/muy5v8PKc8SMoaZsnoEEQBKK/CfntpGQAkfsb9gxt1
+u8jbgowrn7qslJB1H6Ktdr9QYuPG0faKm1xnomYUdyBvV3DgfPdHLgv8mwjKkmM
aA0BTHdMtDxYSxLGMUmU8jFpgBm5gobuznRoh36+s5IFtHFaHXOpxllBfFHx8LLy
53+FlkBrVzrGD7cBYNdRfnsE0DJ4Fz+iSm9NjnxwIQw0Uh4g79RpcvaC56Big3Mq
dy5QdIbZCqSzynLlcRCrG9eapv/sj8qZ32M6hicTH3unYgb34e16yYe6dz0aEKKY
qJ7AMohd/t+ma1o9sB3oaNWO/lqljpheF4zMWe4dSxSf+U/rTwcnie2YYhKR61yF
zuWDkH07Zzm8ddIK2RozEsR9lUsghm5wJ4FoH8BAlJbGtcGddU3mYHCmAbaxvaDI
4O7DhMtgBAZLm6hM9zOnUE2/ffq42ZASiRsGIldumYrG47kaH7RtETFBaSToy7WQ
cSY4XHzQPOK7E02O7Jqzhxl4Broo2z7fAGNDzxzhci+fzBXi5VCReKFh+DceyxoJ
cK1KuyELVhOFelGwohdxeLwLOSdxcEIB66O3eYM7ZU0cYIf4lhFREui2KKbzTuSp
SqJeahSe9Tpw4JwSsWZ8KIMJx3afbvmsulCAAqZoUS9hKn1iujwBSLMHrIILrSKM
ZkDLUXOGDLib0Vr6r4sGA6auPkx7yr9WEoL9tm3hHlB9XEvrJt0sTv3M0szwr2xz
dYmdEssPjxpdHNKZVtkIT9dDMmb2SSp0Bl4xeEMQckB74TDYTKf7hDbiqtfyvzN1
G1le/sA3Qe2Q4RY8PK5cD1aUSBuQN2wClndAjorw8SCycekot1z000mK+3i3Ztdw
uhGZP38vZAir437jK8u6yCxorDHp0Gkwvt1oGOI+oIPue3IbV9ZU28RKmg35Cwg0
8RRfTZsGIMcn8KaSb1ujPGyff6mglp5hQsvLQoYfshTqGhKUDqsz8pQBvRMmJIC2
gZCW+FIaXSCroHTF3ikmNT9G/RK3yfpjPZ1xacSmyGAlRDb3mBEC0zTcALhZ+8bS
s7l9u3TD0XvFuLU/PPsIw9dy/wuK5AUvbFj1K2wksncxdVdXWq3SMF9MhRpOZTUq
KMBRXaF4NfMMQZ2m/+iuMWIEFUZCU2lHI9PK8MytuFPJyONLUNWY8yC6kn1lB3TV
UlTYwFvJYu5AxXyocfY1HorRy2uGnB6xRG5/4FthdRyDMi7nAV87BvKyzLbuVl7W
IA8aQLaeadfGYMtpuvUZ8TNPj6vJnoa92gt9yffXIrJ7ChOUpe8e0lJXRkhVzc2X
rA+sZOM6uSgSiSmZbOZVm4X/WqYuN9nlrZ288afTWQhGJPz3Ll0a40B9x5wXD0tl
eN0kkzipR9xKnsKZBVdN6+nzm8Pcn//jLmoclsIiM0Hzyo7w7u0JQd7D1SnAHRQ3
mWpiSmP9KfpEuLl6sW7nMkFOvPxoIbQ19RSxOjKvYlHPYfpapoH3Uh+cWLesRCQ/
RsXigqCKOwshyA++HqdG/bVohI1seojWm3QIhU9JRHQkI2ztDOHE/xwNmtrP+HCe
nhTz+GuITulIqi0zqIpRs3WwT/YHzE422Pl9lDXvEAwkghthqAya0FhKiqdrz5gD
ZMGUECidIN0m4+yZrbz70PwmOhuyPLyK67T3xinURnryQVJWyQ2mtRvMjoi8PKZE
fTvmvxp+Jkq+IB/lpDNb/XrQsr7zP1mH1InoqdSCqOuAfwe6V3oOZpihYrHHfx1q
Bgi7lj2lqXwAZeOq934gja+h4cjQt7xbky9xpYVbpPhtMD9291OAhLVgmn+2NzN0
BPTjS4qvLJu6LvMdi2rM5AuK+ex2r6IN6BlwzoCdedHPEIgeLPM3VZ7Jx40XI+K4
yFa2AyFSoIJFWwPyGWZaN0S1D3YWEKB4rd3oTUp0Pt9uyeN+eelDBktKGEwKjJk9
OwHUhJVQgaV+3IN38ELSGVBudQZm1dcZ9JFmvc4irHsKPJ985aK8F9EfadtBRYlx
TP26nMDK5Hnmqa4i9/ICDW33EzUQDCX9QTaIdexh3SQuocU9hAnXERciOnSEdQDp
4J8OrwrU02A7+C9ksz1unzRGVfk/5UmpmNVfxtEGxy4OELISbTYHQNKaUMP+AUoj
8NI76VcBkZLlcrLgqJC/SP5AchIlgsG/UH5F0J7g8TgY2JfwAdVNhzyVmyipVx3B
RByte98RfAQYQZ+yHebL8hElhX6NtG6Rh11iv2gLPI3INSZ/GvahlhD3O5CywZDx
aJuSJ8DgDG/Ykf0xQaz7Hb0C0ZZDYsi/fq2tnWjIOHvXnn1IAlYSqPYgOZDZUSI6
+lGNaiGiUDZjsZZb6YpM3o7ziCymqsSLvIurPjnPnbt9pCpxAxeBefa5NH1wbPNP
DmRXpXAnTVO0Ua4YeEW/jmSgJmottSLJj2JT8psWGIdlfSgNTMg4GTsCLNBOR18v
bWhKi4yfVyFxMd79BBv0iknT9mFjpH37UTQz/qIQJT6MQxSegvk1dnM1tzzcTSxs
GuiHHiak2dmn6m17jrPxqp8ARiiaFS0wMkDz+30nAxruwKlSJ8Wu40oj6hRMxUtL
LkuUXxlhlVsRxb1hokNMK/LxQo3iDoD6YwHg2B/1Pk6i37RZpteL1A5TmSAXFruf
anWszk/KrKekZtG9CH2gizZ435fk4cLDzhTSePzedYdi1zhereSR5fm9tb6LlxY6
Qdf7gu5I8ovSx68QIa/yGSLN537y8TSm02pV2zjuI5V22v5TwlUEjLF41tJ1tDNI
/+zqxDp1F4TN1NSSHNcBGV6I7iSjThSz4P94/G4LMSnAQfvtUyr7E+/1wYT9OSqB
FNcPs8VQM4WlHK8FpmIHMJi0jTkvjGKuw8MDXD1sGalBw11jswXMTVtUOsWUrgHq
3ydQSTA2ZlZ+GW+xQbRt+5kmCaObQTd26mjI5FNUxQO1Rfb8zRJCMlzsIMRqOWEB
yadF+lwGN0VvsgBFl1n5xx+64uTTfXmB6kVfsM38epo+y1766D02pLZz7tLeV6H5
Hv27EMGbx/C4z1Ho2QfTHC/1dkeAT5+lh9Sh0xhwuxtiV0M/ICJ+swIXgfIFx3fN
0KGCLp6wKXVIOBBGH0vRKxcMm3D5c+/a+fvEssK5tSLVKTkgmckkpB1pMgIESsiP
h36klneAt1nafz9LXSFlFtQuVaa4u+7QykT2EUQDDBUlXx10hT3XDbB+ekhtoH7u
P93v8Ql8yDxiPWUbXBQ3TizK8RwJJ10Ls6Zo3tifTU5L2YA/nme//ezLPIN1KSUL
meQdyBRCDCg+Uy4bqYfQquYDwHyxnsJz4GOrGmyIfOEBImkAkFZ4YB8SFzEZrHrj
qiMy9Yn1bgDCga4QPJZG3p9Pueze6i2KUOHjNRXpJoTJowTh4zAEv60kQ1HVbyT4
EQ8zTrjj08XprYqQx9spDCm0Xfj7WRGrM/mMt1P2JJZHNixqBPOQPO+Mil1oJ0Lk
XkmLmM4xIfwtHEWRR4Wqpwqknwn10zN5o4ayhdf84suopO1REL1tm6T9cE6Y3zTo
BUBMzISxC8jYhSxzglClsqOSqRkzvN4dafUm9+HZPjNgHnJYL+C0d1+gvD6a6Q3F
gR72rEWKZNIUpi/aB/MWHAZ6ENwp/2gGSRZJKYu6Bq+8M6A4MuneKWkvlQ0VsvOg
1N6IqS968TgYhZXSq05itJxjjb+vf6959WyfwYalsOQdfsKmcsfeRVCQ1uM7dj6b
G/mAXperWIe17Szit0mhC7o+BMWMSFXlYZ0trP+j/08bxo3LLj3rR95cyU6C1d70
2uhFMjUofRPXbcEUoFJetJcsrvkwNwzZdY+fZNE0/5uCNPSbTNz1Onq+6xQVkQgr
QXAYsRyVdoUGj0yLoQ3x8rcftl1s0ZaDJF0X20HvLeM3ekvwSO3tUhB5QG9N5xPX
X6+YUTT2i/6jhfxd3CWTyyN9njbp3E798kQX0FsRZuCXJ0acGC+xR6VHKISHguYW
ifvatKew0OsKPnFfQASJ9B1DuEXoPLTIZMr31ZJbc65je4AN+f6ggpcn3GJqyB97
mHS5/206iSppwM407l/nr0XQjIEODhf8wgNjrMOQKXhGDIPmELWzn7o7PtcfcwL/
crLx1sttQXPdZYpiMp726kNkM7i7dSarhl5hf9rryk5zQf6a3vhIjol3kU83huev
jr9+1XbUDIuMAY7gextIrmf+AUNcxQeCRqitqE1BqazBGWpR7vNxyOkL3IgiDFly
W19SRshD7iPkhnabxH+zYRoxQ6WF3QV0WyiHYKk0Z3MohGyBc65zFJ//2dWMxfmO
dEYM/LyULlUbRv+qwywvzYo5D9hcCTc/Mj2pcqjPLYWRuHGYPV7Llf5l4ja1gcKL
0zKnR6wLpq/5ktt6mDr8PEDwei+LlKphEXFlzWiNC+D5TspgtNpABfWxl2KQ5EnH
JC7BYBebwH/Yl/hHqYcg8pnljWYjvZyGeCeU64+wywgtsC2b5Jwu9KMwPaQZt4sw
X7hu3PPYNCs22MWGRXJDIgs9d8so/9NOi8XEs3xn7AMQNpjrX7xgcXr61+XOJeJ6
tMdtoKkj8QjLsc2v/AeGLGsRfyhCsJ2BG9wizgP/pYZiAyad6uLabltHCFWAVI8h
wL/1LwEyyUmuZ2QRrDiSTVacalkuT8wNpqo3LIOqmOoUN5oUK72REQbX28LpXgeH
zYkd/tGRChnpwYg2pafVdA1/ZYjXjMGN3h9pPk9u0IPcWnHayl71b+15JNqOQBPv
5utF2dpy6E56dJiHpjN2Vi3YrIfttq6Di5L/gyPEEzn5YlFp5NU1gn3gkAcmXzdK
FBimHYU1aPgls4FyBK9kvqFn9hsMxk2WTfNX/JNaVzmg6ULqWW4VilU0z9ZUIZft
6LztI+XE8eax6yYbRGMTBMChMBUcVVPH8UGH39dEcrKwV+ewjLRBQ904ZdLoJN9X
HIyoq6WZ7kLQPU3pX7KWhK++WJ1ZvDjULbqxnkOi0Up7DwpHpFsTbVXH7Uwj31MJ
oYRXzJ9wAJK+mZ3tieqHxNKztBYj1e6GBjjwzC8ly2H0QLGjzhgWwIakWsfbHKmr
di2LsdycM5JC6xkGEeMqk7AyNhV0ZXvVRlWGgG812HeDfql0916d4rvxqrhbxRC5
PUwxG0fqxH5vXEiKMWwd65NahxPejW742XUL93YGnteyyU+f+AS/N17S/KZjRZnE
jBcEtAbWxJkHviPENU1aRB45kFheh9IxjdiDE6fOxiTSsIsXlDCXWitaK0j2heql
WRJhCnBT3j0Y03FHV9IkB/oN9lghkdn6/unYpE33x/otPo3UMWgWcE/Nd47Cvqte
fb1faYNyrRYyahk94rzVAvKCe4tikzml8z+wr0ZzyDTB0g/5KH2omBrhTCpbyeWr
Y+ewYGgSJ2i1Wk8gDmTD4bKEL5TH7WvxFVbTZgT+c4aRDNKnZbRvQgNtN4FoLIW2
mJSRIo1KfYpB6rboorv27kmU+0VwgHMBepQjLJkRgk8OCDMogH1CBZHOOzebdIme
xbCaeLkZjggqCknVSuKDSezUDo+KADPwIi5a0GRv1bKP64a536GM+Nan53lKCCLu
yx9bFxV+YpU+YENoqkLjenaswWFiX25m6FgQ0XZxv53MzjazaAmbwe/fQhL2aVaw
BYnk7/r8M+jQ62cGNNZhh4kjgv+ZeS5IWfmDdapBiz6p7+hdUAnlHOVbSOPIHL9v
ZvXVKjmrjKgoVjKdvafatGDWu/8tFQOknncllvPU6+V8U92F3hNWDG5b6T6efZct
KjJSzfl234EVFCxtWq2jKUeDPD9BtTL5xvKb3z6q6ILRNlajf5INZARyKr0rq+mT
QjFMflXjtUPTaXmcgpaakRCibYRjvUpZosRyuPZgagiVeyWhHboRsGV+Cur+tpO5
LwdquSi9gKNoaxlznjtVG1lWvtkgtPYBJ4htwk30syJC1aW7fybSkFh6bouT1TAN
nEwWHpUPjDTjPmUqVI+v4H+cPfY6MRZnP5JdMyvk1Ows6c/l0WnT7IMnIgOWT6nc
ioPtUpnzG4zstH9Q4T2Nd3LqWHhQDWynehO91+1/AMh4OayI+d8xc4vMdyaf8keR
UOLCE9phC9nr74U7neiAPLBpQAC31qdwMSN1KLY0QcfhM2pH47cTHPY9GPBvWh6v
TJUL8gTDBwPKoGUXx465dGTqhnVr7w+ITL7sgbCAGx3Q20Wlym1QKMMZ1FQ2ifOq
33v0W58xc+6FDhoC+46jpdYh627vfMIb2IZwYH0rcFaFLfuxv8h/vy0RC8liIwPa
SH64l/oOnxuhl6MD2omtOfBhxIMzvYu/q8EFajOGqn8avgzys+crSpJKiM72S7CF
5AglVV/LbhKBy4ULXSLQjcRtroNn6QIZvyNAwxJkf8dwyi2AM9KOfMhhUfeLbv6h
YAL8IzjtO5W4Yc8zQGXg6bTuaOKu6Kp3lWWN1JdSuP2PoAQI+oNccwsla3tZCa1Y
fBcDjL51y9r8xjvQMkfMaYqBIisRIupmw5u2Tu1lDfuo4NTANt8YdP0BrCzI93gQ
FIx+avhXYd3/vG832UbbmLicBzvw4PmH7ODT9YWc1cLA3e4z9Eowa/CuHzoOp/i2
loSboF3m9qRrF3uGSu7RGYlC92ANbL3unUx/0D+DfTplS792f+wE6ojVyTVajcfl
mHkVstRLp0oKII7dMPYBJ+mtQeNakj5iu6CJLRjx1DDbkeNF9guBwHcUCSeulXjH
ZKu8wgnYjc8iWE1bRs0/D9yBiUiXZPPlEyiCGDQQorMiQvoyxMhS4pvn9LB2ItSu
qfvChqnwaIEhiM0oFMmvDsIxqaGoAM0VjBZDZe/zqH1WgZw5YUt7eTY7uvSO0gww
bQzFaOXU8qTCKTolXSDmtyr0cypOI2U74x9NA1oFHLaYnuB630DkEUJFuWb//X9x
Y7ziOXIQqZGAov8VcZDIb9R7EWc3LzdbxbL5rNWBpDM51BKeZi/j2V8VSi4FsSPa
NkZQY0CYgV8zhxN5+Wd2h/9TF2Om84QxCDcx0lN0ORB9Le/oiybOmKaDdXwcK+CN
HWRAsQtt2AzOiQM7lrdu1FojiKJviMjYk/98Jw1ecTtrVoHPdC+xwg1jo1XMq6eD
Q5Zf6/W6JE9/qoD7uweg5Uqw6VH+Xj9CR5VuEe76fxNY9pnA1z1o09FgMv1jiXJp
OYwwGFKFbZah4jMz3hDIOjQyGUWtKY4zDaMgPe7eQ6AcKaSSvWRwl4V8o5cF4OBo
C7/z9+8H7cSywVUy9/zGAXDFH6lrcAjuhiv1RoAtQB4Jh25fiGEZE9cRibYmTeN9
kEfdCPb6rDZbX2C6skBw52uwYjRmHNonwmyleHXkcVWih2XsrImSFonwGtRK84No
MI0Qg4gZBnHOJ5GO/c+9Z9uvrLIQcn1hNs1iR4GJ+LBXLyLE2C2nk9CJ+Kc8GzHm
hLW+2BNAZuziGlXtYCkpMhZr3V1sjiBTXt7o8SV2zAMRItzYZ8JDZufE+MNUbBKm
RAlCqafFYva2qTT2z7DS64gBJ+lsieG9RbEKR1nTrN4P73RSOVgQJ1srUquTyVB1
p1cbNtfbZ2bFYUyTXiYsRkTEgfBeLYtdUug1t2YxQND7YCoOJThQoG5YI5Mp1pkA
G/624z69FUV6vFNufkIEAkHhF88FFHZCeB5c1ImykIB2VyVY8ukKj++FYHHaHMTK
PZY+3aNswkvzucP35PsqFvDcmCLdcG51kpDaTNQGFamVYCG75xjroseIWx6ZMT86
cto9rt2qNfUhxjDPZbGUirVJJuZz9VDgWfMNgtojHaG/3+MnNFSQM9mTKKFPAV9k
7xMYPwVx8KP0g3QrOd9OmymiUyEDM3tvvbSOqdsvt1oUXEG1wk4wSp18ouT0d1P2
yL4Wj9wnthEMPD0H/whU3P/RuBdtNe/geS+daERK3xN5Ved0RF6TXe1sWijJ9Z9A
sBud1bUQ1FfyP/p5zlbiP/YRPY7Cl5rMi9wbc9I/4oqMWphT+G2QBrBTqNPe0eEB
CFDAGe8JeU7USCXruA2i+tW4EJ+Da+0RjpG7YZee1faXRvceBQ+WgeM5Wu0U789Q
CeVDXFqaQI6hbJ71Oh2MtVG+JEUlzESX/ynFLNRfKXDsXCIMFA4VqISvlS6kF4qv
q/bPpf8qiFGGXABl6AX+p5n6w8WSVCEkpyhBFQbKafnTFPT1vK3Ie83+4kUc8FO4
db6bdDxmnAGkJyvG3sc3/0zyWo8GuKBd1mINJ/Gnvw9eFa7aCtA3SuCCVLJ7TN/v
am9ioTunN1jPMQRyLUBgtlwqSEnKfoYDcrO3rukUXntGL4pWYOpZPMLlLfCOWTmR
FeV+IFRUdQ5lOxMaI6Kmph03bKhlbr0vU49cQCVW/HAJ8x7YWSSX0XrwzopHi1HL
3KqiUWQr5RM7x5A3QBRvjJmjS3sS/oIzmxSV6sKUrCFHT8oN3bHBxL+ZWoJFRqoL
6uETXDGTCMlkINSpMXgg0NMARfpeBNZ8TOT0Vr3j31Exqe4Ve3rPxdvd+THUtC5r
jrvL2UMbKC3BdQBeTQjnSTdNbKQr+fU45NOPmQGLfRVZYixic/58cUVA0NpcYfa/
QyXZLei7pz8ryEBIB/o3xqWv4cbIooPV2Ewvrnk1n1ND6pFdLCt5kvYWRC1qrbMm
22c+KNfNdEk5hwsel4iQ654vvtZVJ0cPANpKIR240d4msWmuGgx9bN/OGEm8mGO9
jVXJeAk4WkaMaUH1hUHvlwk0hkW7UgofQTn1CuysKw+eym3Ypkr6cQNxPBkRucPv
f6XQAbXGBYB+i8Zvyrr22D+AWkiApjNXmyZC8qURJ6jhMLjEqAQbxh3KIkg4IUfs
7DutbmRnuQVi+FVfJWKnjFEQQFrB0hWOyrUAi7yIfVvxnoMi4kQSJ5knFdo0wreD
xFj5K5UDX5ioxbOBaCLhj+mZYlNtxCwEqhWFwcxtbBDJqsSBPijND04vX4QEliJV
zo4QShg4xHfAVGFB0lu0aTJeIBmxWUlUrnQex6dn1YXbhfQP1plvYGIzIdmn7cPP
bn15a4jPA8a3nP8lpv/Rk6zdS2CrTvHnYAMBhwM89hc48pg4S1j1Ex+zwgczuYlP
IExEpLM7noFe5VE+9xvlTgngHKXgRL7YabG2oxVF1UTjNofAu9GCC2jLY6OE8Djb
eiBg3+rsM8x8GurIlWeRUZXpmq7/pjj9UkBY1xu672Ziy11mC+V3Q1T1tppyBuLg
Ea6XSWubU0a4J3uJxSENvgMbko0ymnAZb9frsw+VtiogLYXMyKsteAaKnSMNaZVn
VTvRY1YREyn3as4l49oDz4jWirqVKyzdgvyJVsJhHGMnUXbhru2zhRdwAJYr96L3
sZvRrRdyDrKTYsGdDD0XgfCuVmPk7QWL5P1+vgXI7sOLkBuqH4KJUPhwMBFqX/YK
RefJ9xMZJhCFzF+PIUL/AY8GYbnuefM1rdmFD/kkoqg7TeTAlKu6WLeO7OuKAQA7
pmyiqiH+834acri7rwFl82QVfxyMNakeCNJ8Vh4dsplbi7iBcpOBJFledu7kj61s
Fkk/9oiZnCXWxFrLoLuv8MjGcfuciOgJVWOQERGuAowVRXPmhQMEEkyOhiS5amMB
g81fHmJTVjSLNrqwn5h2nC3jHxNBcpj4ywvwd97zvoe/mkwspY2HX07TsrVwNk5t
S2y4pK+QPcMx7jBOjXOhLUgXiBb8woN2g4d8cO1ibwAE+ZKvgGu92c+0XUWi/6g3
Mu5Dd8TAjSCiA6hQAgaTAGHzYKG+pRIVo0NyMHsrtpViwxZJSIhlnR1yJFbmMXja
7t2+8cOXxKh1XrDgeNL7c7pM9YJte1WIsB+qPCWoJv8zFQA3mlKZscYKFj+URNRW
AFc+jooUAIdujO7qHDvnFFioyW6R7bKhMDvaFYvZM3xnD6aTCJGHPnEPflG4CjA3
nFdU0DGrIqtXXDvVCjj0AR74HzM0E3SjX6gDTVuBVdy8ncy/jyIWAeFdQ7o7LMnj
usL24lVEvkJXhUfLQE4HRQ2RedBzBQnrWnlnyo0R5BioFBXYIBCsq5mYbvApVG68
DX9J6OOYvnGhJ7l4sBnQ4DFKl+ZK5v8HSVzJqPG68EhuhxqQ4pol9gfTcycOWT3Q
121fzf11xhvjBuyBT4xCfg0pW4N4m1sQ6W0fh6pkg4vlOTB09fEs+wDm4yQUZiaL
3NJh1t8PPyIq2JOVS7rjYiv2pMEkzg8yzoTulZPGZcB8DxnzKe1XtReB+nuMLYnW
5ApE47AduuLTI468AV2f9VDkydm1Eb012YfGx5GqKq+SQhzVpPLj5Ra55f59P3ie
OYzxGOmiMkXnCCdSrY1HGTh3s8rb+OS92pDEv+DDusAx8zLm2ZcgdsZxugVWk9AR
QYCN/6fLcZQn07zPfpaqncUzy4PazwY65qvqNT80301H6tJ2HOmRZjRSp55Or9hu
ABl7rehwQO1CB/v0tRrpZUwixXg5Kl3IHg1A+CqWaItcwpLYY4AOTOYwUA5mqxCx
ejTjJzU1J2Hca8KJCdxTypA3MZor8UZVSwG5mIMerVZeCPqmv63cF17egszeGf9n
6Z7lWrMHJ6RUSNXXHCVIYy5Z+4neexqWf/0+PXV5O1+lA7YAcKs4DLfb74vvbs0j
Eumg0cIpZZEhQDzNYgQtp9VnefsLM9+r4g27ZKPO4Vv8+/iMh8E7aBAai92vMfED
rKMt1wL4y16Yd+cEYczRHMf44uVucbH8VLOdU6gAJz5V13hJE4HJct/2ACsAe5+K
ahFSo3utZshV9IKYD6F8GPEFSze8OBzOY66F87tqWTYviLNp1Ud3l9ETWD9RQbFL
QS4WgbWi36/zm2wb2uz1DPovuj7NDr9A88cTEaeXE3HRwdHqfE/PRGzfNxRXZN7X
d10b2lZiSvW3+YOZpo5VoVCPk3/cs8QmwNqV8SpqfiYWwIFpH/43SmNKqdek79GA
FF74rr4TR4TE+ZvZjnChIX4ZhtWKo8bUyJTOiZ+hllA4hurvQT9ET57su1WFaXRN
Zo303EhTNRSMo+GKpniUZrOmzGsl10aeO4uSBRhd7f9mWlgHA2Y8IAyqomRju/B2
m/Jk5UnEqWfStoiniltpHZY5Yp61dok18EUOAI1GHSEuXx/CBrP36zSriFd6r2Ps
JMhfrfZl5CggouUwkCbUjW/qG9gnS9aGnqd3I8jLlK8obYx8ar7MLOfsSCVb+br1
5rV5M0xWeKu0uiOIWEQjkPAEZGz0ZnbA4++2s2XqQ0Q1pe5d9lrD7yJOh4F1K+Ct
pyfciXX5LR+NWRKSRx3V02+r/x7nnBw0Qo/LbgE9vxpHNGZejYc9qqIr62JF1CPN
azre+NntEcQD3RLF0H8qIpklfS3IAy7omxJagXHq/hxQFLtFaTbgrl7hw/7knHZF
GRm3A7s0b2UKVoq62dRLlRzpaBO3TlsC9vWIUVq6TULC5yM3E4TOP84azz/dHuru
5ceNwQS6thQmuHIPqaZEmoGRg4CLO1mHhFTaVdBOGXyVKFOAoi7GH2KOOu07eK1E
lGnMCEeqnCM73JizFrJcI1UV6XtX/+wD8AfdUvggTS22MFIkh+cW7a8x2SzmAvDs
um/50d9DAIBpo0z2BXamHB2985VIMDxFXgFq05Mec7Havj7R7lOUeaISRDF1sZjA
nDKIslMpogmeitFVjTu0dKAMDMhVvT8b7kz+bkoY+80DaVK/7odewFfwEYH/dc6A
Fy/ps7t/YxvVfy4y6aEB/gYw/mL6P2WFWaJ+IlH25BMcYQJvenP2wKnV6pMn68v6
2ajT51fVYL+lIdXsENCjgsU2vLBuY5ctcryYfxiCt9K6oIPOsqeQi2a3N4O+02+w
B9ArfCbzu8WtzsbfkbydOi85grHrqaKUKPgnFvYBWPtjICdjCY14YfonhZ585f1A
NWk3uagSozEWoeaysC23dCePz6+28Ye5H2T4BDeXzmqQZpC0pHM/m40fgt1bHupl
e2abA/DkNo2stmEK+BIQfU+rzohI4mOWkWG/nDYW8m6dCOVqZWIoJIrDBTe6Tv3h
I7kdb34qsC+Hb+/UmSoQ6X/EWTjOOoqQL/VucOXc3e/NiL79/t1MMDMPj7YF2S/B
svriw2wE9azSf+0temsC82xDl6JwPb72HRce7js8OlHNEFSS+Zaom/QnNvflw2W4
cP85masT+JtNp43CEn0KGX+ZWHvV6g8l38SzF4EFfYEQoVRiFnbZm/qUk+iOWzBa
ndsbM9Y+JNFv/dxGtuG5r15VNlO8iTCWPDKl9N+NvLqx54n8nJkAc3kiLhbW/b/i
VBeZznCCsaBnzXN920diu2orY5f3R8ROrYIgUEjQtbn/9xzM9uRwZnmqkFAuLlNt
TGT5adhtLZjkmOzKGcZjI3J2WnOdVpyupBtMGF1kXi9IXACJevT3yWWwt8nvjVsk
G2874kw849Eg4T7w5CoHVwiI8RTqxCA9pVhi8q1EHNLYHZS7iR9RdfsEHJTF1jwY
ZLXW+220/Pny9qHRc+QMJ3+Xq8u685PKfDyF8cDHVgBedgc/Xha3M7Qh1uhfQ6DK
f0B9YvNWdIpEyq15UafCH6sdhkh/TBYOPBnUP9wdX9zkkNVYA20fw9gYMiOOQWQ9
d48lKx5pqAN0Up2TS9H4X10DeglSKSlqCjRUXkYbSpZI/+m3oWshjhOsXszjp8CF
8jrh3q2DsWQPoawsxfd6qHXQRMR1LkaMvgK715TxQ/czhWujlnVvXt94eMQiOZov
d8UCNASpwBUIJeK6wlrg5MywPg9APjpDmwhHGEGNZBpipk5dieIEEhzJbzfb2RtJ
cwmVGtk1Oi1dQA0offBMRGRWoP+Z/d+0PDhOXZvvtuEylowHhcEOE/3ZMe625SeC
zXHPcb49BcPWxztBss4wUCVkooqD+5WqZrp3g7ltus7Obps79MbWPR/RdZa5Cg48
yUovgGEtq70yk7r0iZj6v/dW/kgAnOzvDoLOt0fuUvheCmnT6h8oLYzGQ4yev133
yPzRV9QyP9dtmeIao02EvGXiEtQtYtP6lZpzWbAZsYS9ahzfAsJqq78mllh3MU5r
rNGjmBoH1xt85qRBwZXvhedSq3zQ3OjcPeDXDXU9WaYpPHqtEdlM3YXINTpEhyid
2wZlsKPj0VAVbXZxK/R/Oi7/yC1prNHAjtX2N9GDlA3HJQcvEPHkAI1Kop8O85hg
Pny/9Eh+HUPFpWFIi6fycMa5dbGZW4/Ya6XyZadEX37D7w3aRN0rYO/BC00HC+2c
0z5VQ4rgmiuBCJsSwWVMWlanSWmxR215u8r10/zCd+1F/bhlYWrZKxKU8zDkq3Bt
ZfuKCsN6WjlvZh8VWdPC0P7nhpRC1yrAUeKQbjqIm6Z+kTh4fXk3yLQ8Zd2/G82E
HRWsw3gkb12r+TPI5y6MGbR7on4ylnRq7RyUsaoeJXJaZ7YRkpVac2fAo574ykc0
kJkSJt+tqYZ/wYXoza2ZqwKEKNqjIhlhMBqfmatRWkcS5tEhZFW7IiIOaf7zL6Ed
nuHGrp9+tRokLtUGO5q6abvzx8QeekV+0Jydu1+UOOknj3clCxHxL2z3MLQLsIcM
CeoXRD8RvccBzjPs64lFFYUAv6cFT/mjFzC0nge69kpmGQEH8jd5Gb0Vpl7kCOdD
Pdndt0kgZzjh6mSxo8mGYzM5KyjHB9jaJklXjglsM1aAtOqAgvvkywoVHdErBikQ
j6YmvSoTdYtDJ1uVBfVbdSvC4l2iSliRrXw8tyc59a/+d7JR//MYloCUzP2deu0l
M4ArKNBXnFWJigRPJoMEbBmtDVpKSGbPoRYs60Q+AC0nsiVJRdPryqFRi5pkFaLC
K0X0TGqS7WgmiioiYswqqD3LNsEGFbacex/IKQ/iWwWVxw83pbcpjETSm7UnWmg7
wbI15pxgvoGd/AGk9VLgSYwJ7edeFUE2b/r9Jnt8Myvuj+Onkj+RXJW59IGX73jM
755B/gIg7bzAJDi/YwXzpY1TNziC+cw+9YfQlNTzbQGEr1ZHBNp0AS5qOT8fED1L
diIT5GfO0kKqHHoH1gMe+QWKo6i1ZgmfsN5QbdriM9gXIs/38VnCAXM/ISOZSyat
CFwSohUXVa0Mm69UltoKSd62WI8fTU/VTPtnrdEBx+YcgNw/CR6xT98/RXm2agGx
8jtGG4h8mLfmbAsjtlwgo8Qrtg6zU8lL1VNUxYWkIx++vxJlPu9H4l+dZQfoqZhj
v6NQ9P+WRejvI5OnR8OLPNYD0yb4Zay7L0eeMGz/0ks3lTT3fNIJmJVpzLtnSd4R
UucLeefu5XmV85In47tiM0VCYhzFB9jVtFfVE4Afr1FHjF/iDn0fCN0Ye3bTs0I5
LOqM+Cu+y41aGPGa7VgjZsCQ9fSma3NiX57Ng0G6vOpKaz7vkBVhMbimSQaiDa07
sSvz8IqvwTSrDo1UWhgXkGoz5RkmwGCYG29cy2GVpKofaXc6j15HTIHIgMOOTAXT
RVB5Og2uZFr6j92ui7arZe20CIU7WBiarjX5z9LiPx0lw9vQvgTevKPOuaSu4vcO
CPsUlXdYYodQTk2fQb6Zao8cbnVxJHJH1EE5mnKe+gTxgQSbRxEY4LfuPFSJvUru
aZh5HNIa4R+idftB4pDvGq84lInoU4S3uymLk7jdyHvrdUSxk10nOnvqncgeR3a9
5PSsRUdgLAt5LLzB74rgjQY4iuWX6OzYDUbxN+AAH/uKowyC+grSfVcW76v5aI0K
bjnxfhyVI552ST4PwAO5qzBFgZXRNILokGZ0saC4aCXWK+qDFR2se7fEAKNUa7q/
it0rCgGE2SX9QX26UNWUE/BLx4BUKd0IFIhr3GI3fKy40waRf3dWl62urLLKxWbN
wazDz30SKBsuBFWkeR5gSCsShyrq7rJfC1LqK+qh+mbP6JExFtz5myZF6Lu+lbpk
+DDh5gMvuzWn9R2WIafVH1eH17Oc8oJWZpOPKCwkybCobDDrXNUh2fx/0uFD2cLj
EEKkpyKWIBQYHiPUM8j221VdRdnH6/gG2F8DMLS9jHriX3/WERnRBR92VFJnIAxZ
LbRbGYRXipLNso1I67TJ+1U2OznL9cg598UeQWt0OY5g0OnEhuehsZC4Gvxnkdkv
eUDsDzML2cA2xzyXmZs6G3TrB6orn5BY5aiLZnWwLfm8WS40Y8xrPZGY3stpIqMC
w/nsmVPqtQVBScmPEZ/EuDH+AYg/4FEf3CjYRAUFnzMeGkpu8gwkO3ok/6jPs3Kt
+EtXNqt8hPm5mkxtDA8E97n5N0EB/NLJm6zsmUvxmTZhW1vOvN9ZQLO5N6rCirfW
IM1jpIaJakskbc+u0RZfEN/Pf5/eOrel5oReW/ULYBQQNF1+OPFS87IAOj5TiBiN
fDL0Ag13knP5PTkOT8VXhPTO50lg+FfeGwd6UNGDbJFSGf0Ouar1Oq+C867P8ZfB
jdujFxtt1uLySn13LPT4bUEEJA9jAwhoVejlAuesnrkvBJ+iBiaLxxvk3HXMM21W
N1riSZXhEjb11aeQA7uWLDm+fxmFrCXQgJ3VHfyoqq4smeNGRaAN0/HKIQSYF50B
KIrsNjZZztwww9rPRN6N+EFiCIOOURO2A1znQk9s3vAxiCj6+IJUoCIJxnyohqkh
C2MtKcRtSVVRX+vHGVV9OxgWqWG8MquzTUZR8Qd1wY/ekxHEBxrLEVco2TkGbfla
bHOjn0DBuZBKUexFcZLCcqH0Qlrv8GMfiK+x486HJqnBBOdUOFEtsZImLGITBAwN
h3fS4XDIPB5Q5I/+RusiCq/eIhn5MZJiBPYJFZw7fKiAC4ICtIVdtCvbjGDASVgG
Rd/weMJ9MxqJV+5/0ipLClWMl4ITNFfcGgnfHsXn7qD+PLTBBp822SlqLV+CSVg3
QxnMwcBuR2BmLosHcF5GrEPRfoeryk4fFFUwld+1EB7EGDVJKToYcY5oZbJC8L5V
9gGSwvFtXYXUiELP0Hw3wtFdlz82VmqdqZReSkleIRMxNx+9IB4vla9ftEHIjbOv
UA3V+i6IeCXl3M++akPZz1+rLMB+UpLj62K4WwDtInypUVWMfZh1jcV22G98yudr
JNP/QZWZmUchLZlo43Ay4rveo3SUsXril/PaahIG7g1kTlWCPVjWNSuCuqACv97i
c7UZJg2xKD/cxQs48Ux6ow6soCz/bcbQXhqeOPLadP+fRM/FZ2Kk3fyWkWz0x9g9
hv5zX0hjNqfpQfY47zen+1JmH4Mb4e/iVEwKlkKe0J6ei/mIEo4LBRcewrf/8s4p
NWy/s+wJHopAhQ3GJzKmLbVJUVArOIqXls3WXBRAgpc+XP0jitC4GKC3tqzeELfC
dqOJQrOMSCnVqJ3tQDHIKAjdB0QRl6R0FuWwCuwy/oYxAtHXiciulWBQcelonSyc
dcudFl86qt2g+MArkIRVKjGMA7poMh6puNHXPw+ilmaEBrwtFRy4OQEXGvwsNyty
/qkTppGdxGRXQqdeOB7M4ZMnvjMcDR6tTr2bDv3GBGHZv/W8ldNMxR3lOmNWUYmo
2eakkXL87/csymhY0LxdRm9CT/fCosf6ANioiEpJ2A0AsOsLz8rWRQNxku+ex3nS
mpKHs0w9sFem6vggXiz5WwZXZ7ve9W3VkxPW6UIk4DTWsXKrK643QisL25ELxAAP
Ag70DZZI55p5REVcVG8XWA7kSbEspNEfpYfyE7WlCS8YGpiAR4VNR/ADW00cgXtP
joA0eN/8r5eN8wbMrKoWpr/Bcg0tXXxNVvpCSjm8hom/9hQLtTEBIqBzTrO4kY9H
6BJy0bLuCY9wu5cFtu50DVH2TLLnzbSDrSnqsKPfG/gcHsrkrx7mrlB/MRWinXHv
WYmCMCCzF3fSnyRLZviCJSwzLeVs1dk7oLUYTLbU7lCaOM41mPdZlwA3dxJuqa3M
TIgy/OXVaDslC3WKeqb5Ky8B/y8Kk3hIREZvXGu3N/X6VGFvtHTtuduUXGvFY4UJ
IfCo4NnUH4iJ0m/LjXxeJF/D43ruAPKqQwOVh24tRDeIwwDEpqVW6kgFtJgNmY/G
9lbUSF/Kto7YEmsQb4m1DQN+COQy7qCLJxpvr/FQ+2D1Xl/oj6TO4GtH/7dW0HVn
6oGrKcSz8J7qkf4g602o14gyRA6Djd7JMYRkrlxA0VYbWF5sfQL92nVlHm5rAhIn
3VdzM84AXTEcR7D1a2bRcvSt/deQCKwllGUAygmIpxbKsVr/SO5Q11VZ2DkuLxFf
+DMiMNpFr9DkbASC377ubsRrkY2affpggpBVPqt/fg9RZPxj/y3WzxnxiGffMzNK
NmBabfqdoPlbTjlRaTWOfX5uLnhVCEOk5YkLB5gbgC5lBxdFgw1ZvbC1rA92iKzv
q6x2hSE5WvkMQaEACL0+7bWNStHKEH7ZuP06gxN+b5od5mkWK4WSPRbxlna9LXyz
zYi1LGInijQHZT/PABcWwlxZTwM5uoZgdgSQJwMCGKzUys+EgNU0zg/7sVGgBpw2
6eIq6cpCwdSHf2dN/9wH4OcQSAd7RGdG3Vd3C5+iG7j7P6Xn/lCIr4mPL6qDMFBA
GtlXrBsufAHARNpOLxmjBNhCaPif4NOz0vCryTty343vxW1yhuuhPiuhxkeIDKAN
Lu2OwB4GhutGDYYojkZUoKg3elWtm9hy67oSeqiWdzHrVKkUolvT+ShUQGYvaL7e
PeNEJ1yV5jc5wh7kNbG6UQvcapILMTQp357nN5cBXAtD5ZFU8hEimCW88alYdQsb
q0aHRK2tTJRwZdJEufgun4Io/lIoFjqawXFOPuPhB0Wbs2izsjB0K3bwWo3RaSih
6x6jH6zm1v1jP0db+bNq4xocTIxT2NqcufbsYzJpx4a+R2lURV+oBte3mQ7/Tlq4
kjesUCk+LaW6869rFVojDDemk8KBz7HFhaBcbeBpMwNd7cabRr4WhVYah29f0uQ3
riRqBwUrWObTUJjWgwrBnj8m+8HuKpFva4FMoOKo3aNp9w29zd+QY6U3regMBgi8
rkiHfZAhFB+c33HCVZoixwcMRNCuM16Buo1gYg6UEaSwea9NPO2TaGq1GLsW6OeO
L/hgn5uvsusOKvt6ZYPqGPuzjTpdn2VjvcN+pB1x7ZPGe4iLMTzLin36LIAzMUkU
NqwG5M1kvAscxwSgLdU3Sm/HkQAre5EiB81c7NiOFW10VpzhEgnCsA+NIOg05vuD
E9DzqhaTQY5H9fOJpFuMqQb3Va3nWEl/6PIY5qBRqugAFMf1aKzuKG4i7go+nYRo
JAkb38KvDEIGOfTaOr5m5fTFv2gOxBi8PYCzk9szVIaYsZ1ZrphuXIUEwHgPS4nd
D7AidDLE408kIVcmL9TjIHANzyGkj2uEHM8U9aB8frAaMKXabguTbe28xbb4Udt+
Vy/S4ApktPo8GCRIMNvRjacniP6kF9p/ErkOxU5KSaRliGy1W6ZBCD04MKMp5Cc0
04a91O5NYeWOlhxIPgYSHoFrwqP583BgD6y5OUosDMV5vB0FcWTD9kTV0z/SX4hf
GBDG470GOR2jFxrsNtszG7fAp5JsYgpfX6b5o9byOOrG9F50+y0cg8Ye+DdsSIA2
qqT3d68mWqTJ8PgXEhBiLh/K4cfxgjz+ch13854a/C5wY0RjnpWLySLiml+r+q1g
KR4mURAUhlgsBTaoYICfdvRDu3UrgoWS9lPvzcjFnKxhBHuY5KV6NQoSPJwULFQ2
E9ydq7P8BJcCvHXHKXXv3DzfelU0vcL3nC/X+FI5FIDyNe2RxcX/OOEiFxOmx2nO
2ClGSkbeW446aqc2ayB5JYw3YH4s5pIh5mgKJQlWLUt4RybN8Iqwal+ydXQQtbIw
qTbosckSYEKPCgr/DSJUuQx5af0eFawMvc0dFbo6+2cweVBe7itZz280rs7Dk4rz
J5CgyApoteZfGmwi9nRxXQcxtUU6CvRafkXQ4Wz/j9OY0cE4tvJOQBsfAE1lWjTX
3KwvAt2hQGPeiWv+TCSWVsnw1memEzaK0qEE09B/N4q9p3vaphiEVJzPUVnt3m+w
2ROeVIxM+gcqXR2YCGRun8OfyRPx+tJQlbhO8NpUaX4rypFGxOrjFy1R/ROz7pOi
/FAkLR3oo0MlSsjIQzbApNMqlcOrGZWbIQ6pBZE8Y1b79dO8Zpg7e6TfAHry/ZT6
sqj7g68DIRnORMJmWcPNlm4UiD346JH8hJKhcOpKoLeEDzdcwlNMMG39oZz1RT1C
8wxdkRtjSqCclFLzg1nvyzjazo9j4AmF6v1jyxfrWHVhllUpOUb78B9uoPAcgXVY
FhZfEiAhJe0REd7xDAjdbpTADQ8rr+CodryiwH00erUYJAb2txyxh21f68GyHWsQ
0oWzh4AqsgYjj+8XdqmcYU76/BV+JEiee5kdqUR/l1QBZM7W9NzmEn6ERK6/Rl8P
L+SAM7PuQFjE8thY+aU6SdYlpQmCevnduYTY6QlRvAN5Am+b+Uq0NHOsy9BL1o/7
YlWHqBXHBpWbMY0IESLLzHPKVx1ew2xGqnWfBWZhLqWQz9aXBepxblKneQyzCA6+
6PMnv6LYisZlVulD9/zoFU4Wq958EFPWgDJvFd1gTDHCyZ6k3T30Kjvq0Osam1IG
IGouwdkVwn05OIJ+i7l3e2PFR9BFlhyGMLWN97+HuAJ2zLUvgwsE2s6+TCqnIMeK
Y3ObEhR8D7P+ArPXKpDe7AbsoSxVco9lMam03yzZoyjOBpu4Fm9l2p7y3HSFxK5E
I+UIQOPn5CBA/5C90htm5/152WO7AULzJV1AFbQEJS/caLKGpfZL+je3qi4hTSbn
bQAnw9wFCLF2Wa4e7tRSc00SmuRhdvI0jepq8Es7C0QwtTBfqmYIBmyuuEKYNyKw
ZkKXQA55h6CJ/vRZtES+CB/NTBr3l+51+v3yQo/FY6VeaX2govqhf+CFgPIU1IOD
rozskUTB9MoJYOT4Q/4hKDNEraMJUqKQrc4OVandh1/uCWNgkVXqlmGb8WTW+luw
XuVpGTRY4UCNP7cIwjBoCeCeB8ovmG4QPqRuEvtNTxI6XifmZLEL4gKu9TKQMCht
/MPDlIj1BTh1S/v7LugDnU7cg15SmRuXK3Ppq5rVqOPbL6cnOIdwM6Yp1MISCoE/
ZG4DMRbZMcXgaVriBao6eSp3s1m6JPOfjyW5ayA0mseoOuKaHTEMsygKCAxGMPBN
9GK601JaYlTCLgSwdxzKVhXy2jTh88Hwsd9r9YASN154qrfEq+1xD9I/QaZ7OgUn
kbqDXui1I1U9Vs7KwZ2cwmGCLnNlteuI0dWRDKofatjNNMCxLTpVWEnQyYWcirbV
o0y4/I9M144N54L6TP2+NCr1ySS+EmIQWR0tfh7U680Y/6eRjIDob6rvW5PrT/qc
awWfwvTCPrjwKiI2xr7lcmHyyM9YTNObowlipCKqdcbB1sRT69OsPywl+RvCGvw3
BeX4H3jTjnnswgJ6aMD65ZC/ZW1CuZNPt0EeJrfDNt0xWGLLwf1QoThMYmyH13QC
lLOO4YyxG4rrH6ZeNyBxBHvvyIBnnd8fNgEhGkvo2Yzbs4klNokIoCaD6zhiMJ4I
ZyZV9EUWG9rAHf51uB0GEGD5GL4BdJ7jG3Nr4JaH+EyR91jOz9IN7xCUqRBgXa+k
rF96S3Jwt7/OYDgXz41MHKLxjt/FTwovUywqWaSIp6mRGEEHLryHX/6g69D3ARqC
NdPqwTSqmwVycmHI4WmnRUCJRmuTFz4IwyQldRtky8xZ0NIv3H42aownSNJYf814
uvtPNn57IEx3fY2EXsn82MdDeLqSE+9mc2MA31E9yq1voZznOfjy9NOqg0i0gG8M
6AIZ4+QUqUVFLabKv0IOrvEk6vmsj9FmzIqfGhuZhygbOGHUHAXFhRyWaK8JZdxY
qrhVjBQL/uA22pHxEb5M3jFyiK+uQ7AG6lbj7j7SBScHsCShTGjsbI2iyK+PF5gq
mUaulL1eqf6QHksOv4N2/bNdKp4jB7j8M6aRy9nNu8r9ZW8d7F2CPKg3fXJLQ8bq
UV9yflnaYL0h7++R9qehpDdEqd9EFbZj0cAcGuB5M6vwqcUEbFRi4Rk0gS3Chvjd
6oB9nqNk5Vyyvx3tQw341lJMgo971A1fnLLav84Xfgd/YL0l9V4D9rAYLcshsfe6
Er+mU8QRalmChuOV12AmW3aLW+HSIwRA6u89c1SJ1KRH9PbUrrqh/eigKbhtXtIi
YAsrQ6tXVo5u4wNzJu553i+/W8U8sPhNMauVg1PFXhaNPJXMkFpLrtRlROecyK/m
cYReq/nfPjiAK2pzh+Sz8tLcqZhMzO4NSO8iM7Gej9IBLuZqlNYYAW3CzPEmBgSD
xQG2KVWJfuBIZTdKPfjLSDBaM0ncaYIFYfl4PpIhIddzyrMqxAe51NmJvZTCmc5d
GP/24zaOEqcgyp1JGFgb7BgE0aaZpeVcaGjVf1RjYCDp1XKU0qocS0oXe4161UEs
1QOlfDwvaN8UPqZSF5WJqxrWvS6WPeiwqldrb9BWC6gAOkzmd1c3L+0DWGSkBrca
RqiW6OJN1kK63ACfKgOMcDQdgIfYaHL5kfpEYwMezmRQdpwKMQVCjOmSwRzl4dVX
BGhpIyhaUs1NgS41s3qBagcaF3NwtoC9vTuzUZVhixoJaAxIaqY49BSNVhkd1Y1O
J9AOSKmRvKrj8WKcoSVIX+uPttMeAF7eMiNnChw9os+QuwMZyXSMartdjpqI5ahx
AxVHTUQpHsAARMsft8dw4oezAcGbLxEs73GgBMjAuoJofGnuyjghHDUb1sHFa+Y6
NW67cbpPvX8w5j9k7QqJ3S2wRh5OnBfsvC1F52yMVXWnuEguDe6A/q5Pz0/+leQX
xEiJMFYy7Dhs7bE9w8eUXqxuVTNErl3+GOEoidbWyciNEC29xFYUTxLOnFPN9Zfu
YhIOKZtB9oKjDQdLoP7llQAgNcMN8z/0GMCDNYpvZik33GM0cqruxYevRfC8n2E5
uopa/40lddfqbNuTNrsch4fTsPQlFSBh7GUezdX3HVvH9JHtzP1nDuYsTvX1thu5
i9QotphaSVGSfmbvVmLG2RNUoHEOBSJeP9Tv0Xe2dyR7MKKj4sv5raH9pywawUnE
rsRpTyWdm+FBwuOHOnB0Pod1HT7RiIHhsNa7bIjsEhVb6mxg1kOU9obLGaSVqvW8
egVdRiEByI9imrSwWrk29RwC3PArvcjEbzKYE74AMB5yedg6c7DborADzdOMtb7+
p9jKAYRIxJDaGODiMgtNeLA/OlxIxYXFJrzF3Bxpc1LwqldeefvYsfqS8L9ZYWGV
cQJBshA6OLguYGfR73a0iq8KNN9cQzROMCD9XLK7Csed7z51tklOgiDybd1FjY9x
s4E8ZZPjqmMFNnPJ6R94HAYIz0upDwCVsuZw8Uv6xt0hE70JgL3zgt1v5Fs6PJBP
KAoIcnCtZvMAQ5QJXZVXLQaoAgWRc3OKhA8lCteFPMxMCz11bsXgOYs1jB+O4sUR
8DFN1N1OSA3kjkvX1iwUSOi1wwwFEjOmlPujW3qYurEOlDUtfUuQLzzojcSew/3a
FA///MDPjB8qZT6AmRAcIC3AI30h7gxgpUUCV2Gb/hu6BGf21+PN6CjHyQwQkRgK
wYiQSItL+rFJ67zTkWLs9v6DMIgLotu9eCiLRoEJJLnFdRWmA8aJJBbWNXDGoH1Z
7lgJS9KNNjqExaGcb+HkWuCfXsoeczuSdnhb8s2od8RZ5VeGXuuI944di5+nzpQj
sile6apq+gyIUAy8g+rVJKIl5bEnh2VZiJRPYEZutjDvPNaF+5IKt97wB1LNazl/
ibNP7lkbpPe24TvTm9NuOw3MgInVZPkVZ1XFcXYl/aD1kUwJDRsRt8SHhSbC/3S3
SWtt/4DKtUjK5IqOcOAKGqm3UwHXtZW4ZhjeBZgZPgZM9YEFSJLccJhYuYA5qP5f
mcp9hSP1viDW1ZfK41g7Kr5aSpusM2tVFaQZ1J5R36vwya660/n99sMCnT4zliAu
btN/eQBBOQkDRnbrfhpae38HVi9oLy/pIX5m5tW8UY6N0KRibhToNNYRkgPNM8/i
7nKUPZTbB3ZB33BWfzog8r2rHQt7bpci2YSmEneRp6Vt7RRGQFsPBH2r/0Dtc/ru
YoAZSaMlc9NolbbKoJk7/aZl1oceDLN1quoagXHL/Lxu9aS28kSUn5Oc/GI+xUnQ
SkzEM+KXVzCpLUYu0kxjilP70P891101PiWgBygPsRtX9k21TMmyNLlUYp1N66Hx
foHTdZp4kfaj4RsmOj7nOjpdE6Ejkfo/s+e77FPwJ79Er/d2iskZGlk+GK2hVpVd
7dnLKTFHMUN8U52bWnJntd5OXy4Imwfw0R6bfphiH6xU+htscK5BHGnRDbqcYZ1+
6P0HOodm6uzm0WQv9PvCtsU2z2/CuUR0kGyZx5zKfIMbU21zETARidbm8JKTkIzd
flSjEgDKe6k9xJi6mBSyHFyYWOc1tzsSFWdGG0/SEEGlI2ebq0wcttTSrxGnbirK
Rwv7Oq33U2+5U9asvqWmgrobt5vAH4OWCrJE6POSWOA3GkJIBteI/UujOHlLS+fw
lrQ9PYO9XqHHW48IiU7YbpLpNVWmuMcFOBnTuX8aVKCqvBo6i1H4WKXNqvr22u8J
MliLrNkiqYrva3bG8Dx+EhG8ZgUHFw7y4yq++tFw+wH6SgF585UKh4CrtTf1s7i8
lEBffzeZl4qcm3TT8s+hkSRyiWcIVhUF+aGVSH2Ctsm4Bs+CvH5CsT4zrbUg+AGh
mnCqk6JNXfHqEFEBE0Gus9YgFENoxDtFax+zGCVPOV2SLok+78Frgo8ngGkX9ccQ
ZP1bHgCZwPL0wpH2Amq1aDPSPmosDEjYqgHyUvogk06XOtV5H1PqngT3Idjr0l+P
NZ/UGaiIJ+os9HIrqpkBK5M5X4S5ex/wp9TUtKH3Q5stwpsoiPcIxBoUPmHqKHGz
iNdOQIdED3bY1iKTIGYNPkDUkt2H8k+ZOlGh6KjGSGxnkDFBd5rFv3uWPRpLsE/m
Xkt+jpygOrYJqv147xaIj9VqztWl8X5G2rRpVJ5K+sy2nEgSakHeV+cpDU9EtipH
cp7waOM883D/mI+Jc6ELNY/cD/b0GzOp8ycGZmvyVRlziFQYXCnRx1U/Xgz3NuWZ
MIs1Q5mx+0juThQ473mzSt7TT9Twz5NQpDVu6uupk1V9bvC0zTDEVLdG2/Htw3xh
WcZRcmIxKWmECR58+LLctzBFAeHyBojLVn1/4/mN0auqVXC+i+XkR3kj4YqOOHCc
Gyvf2KM/E7Ir5+aoWl6gg7ZSGkwFa01YWlejvV1zqYywWLk3ZKLssiFS6KbRmSQQ
E6vVIbzZ4Ll9ikyoV3qice74NBNr8dnIQZyu04sBaBbjwsLrDnItD1J+fh5oUbzX
AfTmqo1gDIxb/7wevBoGoKqqoUmgTUDwEAxr5uPwF3H5kX8EI4b0Guoy+F2V0A/Q
pA6sLysxMs7XDjOKMNbaxneZW+dQdjeHC0zmjjhXFKlzH2c96tut8+di1b3/HsfL
z9TTe7H/RSjGMrp0HnzBgVIYL25WkBFcIkkVWroieLMbyKOT5Qg+3GPybrQNvKOU
CGgZ7liSMP6pIajLJXvhOlco8hhgJshRoeeLSmlRcamXcekL14YfOwo4qgUCKk+O
TJfgswEss96nCVBqDyv+wvmWeBEbIaq7vTrXO68keU824K6hNiYqyLrVyMVNbl0x
4toJdqMKz6hurdHWKO+arAnQekCN8HVheicB5tR9qxFdVBb0rQKPQdIgsSBt8Xjv
UxxfuexR4TXHYLXQDONL+b7wSQWi7Q/AIWGGwn2pYHSIIeSpljlX2SUlxveHOeby
2B9YHHivLPGn7pv7GQHuL+6egwY/4ZbKksyuH/S0MIvR6YZDaRnKQUpxbv9nDLOu
7uaz7elgqF703nXAVczxvnHZmz/AyjStxxBDHVDxiPTXQCj62hbtbZRUa1CQde9U
p2nva2j90x623H9XFJTPtjZENLsqgWAhCqUABzXl8pVAZoQDflqdexoAMJX1PkZ0
p6T6vfhwzo4G/GAk+rgmF8eea4v1Mt/cOnup4beuBArATbtAgankE0/xK6raz1mO
MgOm2ImItU/q3aDYxJiG3V2Zl67CZbSS+NWWC9iTBv8AMA8L3t6ygydnC15aqr4p
xGYE2aPrzYoHwPcV+3FWDpD9UNmIjfYetsUsTepuRT0s2KAOQIyT7C4i7Z2GTLz8
rwfPsGlO4FNPKeK51EPrFZTnOaaoLreS22QruBv6REmDHFIzH0lacxXgmUZgYXnC
r9JpnU2Ns5zadUB72xzSAbGPdJQup6qoEL0yNeskbvNu7q5RC/UWZ4qD+IvxPmRs
L+HMX8CyQV/lPpYoEOmbdh8gV88hEFFGqobtGaZGkR9yd/XFa/27/siYpQvd0qa8
ZX8st3pI2ktIFjy8cs8NO9kL4ykkTrV3Iy6NauLn7LCfHgEbM/mZGI56T7gQX3Y2
ArFpBwXiM6jj1y1jNGNuJotJ5ekcVuRtoLxauwGhU1w3dRKgaDsaYtG4nHcaqhwo
fhFKF51Topp8hMmni98/LEmrI55uTcb/hxgwMTDKIMtGv2JZwLWgz6r//eXW6wwm
UuNcwaZVZgPrY/HGjoV3ywije+ZdObwho4tL+wXukvbPcXZPTRUEj5S5pVzw0Mv1
oWg6/C+s2K3pupimczLlqdfpWIX/LmhQhX89ttw4DmzmYH8krHittWfb4JYnC4Kf
D54v4WCWPLNKuEFIc33K7QPxP+A46Os/UlkzkJW34cMPzHcGs1WVQrxA9Q2v00XG
f/Ytv5q5s+KVD0Y/qfYzIuzU+3ptmkgAD2LkTC5NR+gYJB0cX5OHEznLkM43Ls4P
kSpFEYnLdaRWckiLIFFxpW72BinpOnAIXv1L+xDkTyh2UKWpEcqgV2WLILnP/X9S
XOoeBed5M3wTyvJYrhw6T2GZOz9vSA2z6u77vSnSnS+SUPetpJEbaUmWdvLbIaMx
nSBjaXDcpMB7w1F0oG1WRdZ/2JCpIo2gkOebjDO6quG+HCdOfyhhekN/bhJcNuqk
WN83KGK5jwigmY6Cc2EFPup50lbBRjnfk7IwGuzhjCHa5zMBgRWyCG34zRBw91PK
evmSWJy18veHxEYADOCtd5VO4t2scJphtYuS3pZm8TAdnSS6YMhQhDohW4wNkoF9
peabZYRmQcQl7Q1L6sQmgFjLtafuNiQmKG5vS84fsNoE1FqgNxEIlC58lI6Wixs8
o+HO9AAT/TL68kDbfGdXVJadYqQNZ0zUnVekKTL7eRJdDA0NaOoajcZ2Etti6hwm
Zq41l565l6iOPaKXJIxaj/DN26n68GWkN+0lqIkT2W6EFXmIQiVsCdiiZozW28Gx
vwY5vZd51aStc0oOaNXGdHuZ4mPCijX6X+hUbmD/WmIk+xUjpToFyaAw7S1m5Y85
TDHvifklmrBtZz5pjhh4AycE5ZKhNVB9/mr1kEY6KNY5BSRy2EL1ZQbEU9ImZUO8
CDhnJWU2R7uu7mHv9ne6UdPl1YJC6+rnCP9Ho+W9p+0rkcVyAsYA8VHWQ1HWOvJn
WuhMXQoKG5dC4Y1wbZwKavjnQNzv6G3w+MLEE3TlQhDOeZaG3Tbeppjlf09udbXk
1FUpnWzt6HQJUS6Q7MfZ26ygw8RetEvwzM2gznrMa5kS4jvnBoZwVavQxwd5oqvW
motr5w/XmoxlsFMFvdaHFcyfafd5FU1oR/UwaK7dnCTtjtjIsY3VBRmo4/HZcLML
oZbBkLQgVjleHDI+Gk6VjshgypodSuwGo9qAGHxIokOVbt6+NSAHHA6q9R+jckJb
losSAqRobIg2xeED8F8BAO9yKJPf8hw8eBCPexVDLzaATNgSAinJ3f/L/PctOeE2
6vnSYGnW8gt4kegwxGEgmAkyz3XZ2clwK0fceiLMs13gw5SRvK3VPy+Bqcb2y+A7
yZLMm83nEgED664Q3ygt9sAW03pN+3Q+gyMgDgUc11z84qc0SPnQJU1EC+J3eeWe
Coo4RjgDwztzs9pWJ9MZANUAjZZFLz8MLs1a4X4rYNkaP66AiT7q/FSK7idZL8Q1
8HStCiZSujqTOcxIWeO4+qMi3HElTxfz9QM8DgZtLuSAisUvNjoyvYssTPVwb+l4
MWqGnFayKt+i2HSZhyMf4Jg+DIbz/qor8rU/Jz9j9jHNVg0LVAElcQARFCApQvd/
Vmtzf/4B8jCorWX7xBda05bSVVA28pB4N7MqoZGt/6NgousGn9UQzbTQhS10Lbmv
iT2og/QnPL0NGPETY9tLuB9N9BOQa7mA+4oq3ZROYnDIuowjjoVKezMy10we7veJ
9xUAaknzdfvX4PuwxBdFqgJN+3v+WcpbEOgMdUGaGiU5vv8tbne/r0s1nMk5KKGy
h6Lg0E+PbjLhCPl5EzNljqJz5DOTVNy284CnglhpoC9wpjyv/8IiKcoFBwwuHSfF
L+jiFf65aDyWftGnyie6YIKY2eeKGdCuEs/CXX2OMRWGin2fCgb73YHNvKs93LoK
8TkPrxWrGQTT82Gq3mNpVk8tvJe0X/r/YWotxlBN8t7jxtxEJIJMnqY6+FDo0N9P
IWToJX2eQWazdguGKrQwFnCDtGk1nirCV1vg8r3XVDiVEkoJNHzW52Pq/Yfg8e86
HeO6oDlSlxmPkzdvKAorrFuUN38mrRjqpjjyDMklEPCawTZudPqNzk8o47VhWoSE
FsYmwvrDw3kZaWgf/A6kVuHK4h7lh25X+rFFdGid07i5AB2+DXgn8NmIytqvoiYO
396b8QVVn4Ej7DSdWffmczV3JGG587fKnpmt+nUGye6FpTASqKQAwzotavxGCZui
AUr0weBvxApp9Vow4TIC/5NqHSVandqznn9YrWMxzD8eAH7qwhCKUS5HIBKaGMCU
z4aNrLns6qH8xe9HsQrRc9YOT+EsXMvG3UrztGDuhWMpwQPbNtqo9Azg6awDANWo
MYTR0+BONdty3HWYqsXnSef3WfirCpfHPBB8MB9RPa0G0cW7l0ZN0VvptPJxcreZ
p8uEp1lhSeD7R25LVpi33UvgQfIIJbmK1wIPKdHIQXnfLBS6+Rz2p09aqpGxIyW+
OrBzpIGPl/1xWEbRaVReDAr1xS90UwMPLVZF3HtnMdLfQegir7j5ASlQHHxhplcK
Lx7VOikA9Njfz2lRppcXIAmrXoVR6Nht60u7dK7As74dxIgJwV2g7u+nDsa9B/gC
ikJOGHPk1ufoKihkmA78Nwa1EwpVnjRgUzK4/wsHccHFD2REUlTQRMANWhOHDZWX
wBte42tbPN/kVw1BD+ADiMmHf58kagrpbU0hAmDuI+ql1UArEUBigozst5SD0Afr
qaNaoNOuicd+98h7ZIoP6078Kh4OkHNRi/GmxkWNaYKnREsiHQa2SBAMFcyNUvxX
zDD1d3yrKnU3guN5i5GspLIPMlF6oysnCyk9t1ZKx3KGNWRbKL130jyP4J5wTAGx
/NP/G14AmC9HOB6UuyB0C6UkMp5l9wxlzWpsiHjkQkA1jv4I9jDac9VphHZnMARv
TuuIiaO5IJVdPaT8UH2e7OZMnxIXmawTSdbkJHOSETdwTpim/rzYpE0pywjqUaiX
dCNj4S4TO03/wWrt+oIRfW4OirlqrHtVQ8+FE3iNj+a95rIYf4Rybrn4zK6qdmwz
ga5l12Jyz0ioEf/IHmmNTFex4d94MGMuTnYuB1FYbiyky8MaMjbgTHTaqjyKk/Q4
y9iNOM4kdu0DtVul5ovNNClLVjglbGYBUWy+G8mN+nwOMNbP4uswI3jTdn8LsIlS
cLNLyaAxMVdWkGOZ7Qo94d2z+1HDZK97p2X21fcu01KuFfI3+O1Hg3qsT57CrGdj
hiItWNKAvCMGhtmtfRQmZ6nzpAFu5emy73wpMOzRN4UL+fMQcXAkHs78uX6AYfTl
NNL3tEl0cOgOS0gZ7EG8hqoeYmuwC/vHDz+7CqxYrAHxki0lQ/22dlF1sNt9xXED
xDwrwM/a83tEHbxXij3y4GRX0k3VONbeWbR5rB/K9vgSJSEDmWdmKVItpndzJ37Y
/LCV7YU33rtv39mG/kgLw7x6nWctr7s/NvMwQxgm0leAievaFbnUkGIfE33ghn/y
Pl/CJi+UfZNBM7Cgvb0xfRg+RsWTn1GaCswbzn8YkWTvRvYdRfHekVS5WnkbhBzL
b7FPjxDkn6d0WXRISkgNpFro1wk48T787pXYTjxXF2A4MLyOcwR2e37QAoFZA5rN
NlzwP05o+1eIWAxSMxIwAzGNrujmXvQO46jKYpTiHU9NGeiK/HlBG5r4K6rOawcl
/3E/e1SEJdM9E1HGjvuPoAjhlexTi5McawKXj9rE6vB4EUh5691FcHCOmVGMgEQ5
CChH5yR60/zRvYCWEyULxJlIcyxPvP9kBemR5DeqbLteSt0+ZB5egjGHYqliVd1I
MhWnpMgrUuEKx1FdgFrPJtR5AXkS7w2pZwwudXC+PxDv3vCJJ3DAl0bEiNRUd7b2
t/9/LivsymmOB0/erqLnTo4hS5GdbJYfx2o3YhNScaemSHeoF+ExAtzvvbvfNe5j
+3MgMKAhWV93qBAejjewERGoZh5uVIODSXnqSY4tSzfoM+eVYFZp3qztIPvTu6Ya
vLPPMCMzrAKAmUvPJPv5MzHg2vDOeZwSJY/IumVgBrD+Y/KNexQleqjPOBN60xsr
CbyL1R3y8PXSD2qJ0rokST2HPq/d0srVA102Rq+zffMGyWwkfLsUUpHzMcRVOsMc
6spXJxewBhIye6aekyWgES/9jo2F90Zuii688l2c55Vhz7+zqz72owD/S3++C9MI
O5xXlA9LgtYI/1s+/X3WDwFFv50DBIeaAUxxWnbLeCc8m7cyu/TQaduT+jcOySXk
x9ImMA9DHbxRLvq8O0S6tcR22gOtnorOyZP8Q/+kqlfmNqQ7hi3ZHYzkIwNIHGLm
h7lhrm/rSf+CjtxT7iL8W+mkqr9bTq5jQAeyMojpkx1IvuTBfJ8d/3/uEu/MOeBI
jvfZfKQIXdecaaT31YMJZ5qldQ42Mo4dlVeRFib9U6hdxcRaT2qV/Tib7oQpDEZ9
QrSdmF6SYhQpn38Pt2KmUWbtWnEadSlhlNT3we9Lo3oNhp8ng/lj1d5lJOpz3vVA
N0JK5kUQpZWEf1ueU9FsmMFw8GPZbUvGfUJ4+0tt7actcL103c4O4NUQHONqOESj
0FdXqqn631eUgiQJEgEqs4up6LmYJG/sr4hW4b/qBR9xlBWsG0mmto+sZWxBlfeW
3Oh57CicNjkqyb1a6IwC46KnGeInOFvbH6jLpvqzzqOVqUl490sWzG5bSh7m25Ta
JdMLXReXzr5MQrQLDrkzD8W+BIRzLcFk1LmlKw03+e9usDNxIJqGvtWGyv3Xzs7a
95tCWYKpORoFht4wFDcVBRzNTwHm5X9MnoqC8xsPVlZxkBO28wdr4s0JZIELi8RZ
iKM1bd4/Kv9h3h0siulgYTmShr5SnE7uKXTn5Lu3O6KJ58c9iTXDBLV9415LFBab
oWuwPenrxxZOELMevIbOIXMMpbOS0vtM+v8liz95P/p1rlCVI3viYmWc3kYuS3qH
s1vfwDzzSvfaEBXduwMB4VnhtAzQMYN5rc7oUO56NucvLvEv+8dZEYcweNmeHz3Y
G1FfQHJJVnTSRdle8wFb5tGVlSBXa6+TIlyjk89Y9ox2r3CkdSNXRhUxLtKGF9VD
ay6DlPV700fyBSx1QKSO+oVN74E28Q4oHMblKHCCM/58goXHhrBB9I6I6C+KK7p4
XSTU1GXOWwL1Ebxl5z65d2v0AX2Bf7Gho7vzGm9LGY+Ng5NgjVIMUpW2oXoU8Rc5
96HYMQCS7NUCfKQ1EbYaaCsNQdfYnqUU7bbEQX5KfuFC6mYTcrdeOkURV5gB+ysl
XSEYmNI4XJBh/dVrSt8536WzZSBs7XCFxSc+/ndYQ1waekpj1y1OBmBvBv9XIf/S
rweK4FCtQRGR3Hh2ydqOyinFc1MeI3I7zjv56I8lnatQ9QGG7UtXWYvanA9nNYC5
9DdIWjQ3UmQT26vaooOm81g1tl2pwv5Rq02HNUA7sHEFAcaXH1zsAk1xu6FpsgNd
9p9oQDrrf55cr1+NzXtyIxi92uVSgzpNcAqIxT19HhWFARzjp2Rkuipibef6EvZa
CY/Xzck+hZsoQVUr7FSsk3CUK0xBJfxn48p53sc82edgDk1+9yJGLE4Iwv3kbrX+
PiJEoxNtx8u/itfqhZxhQVgzM37A6Plts/REQLQcvCI+m1zyGgHf5V1brEDOmOIC
AeAIYOmenCs17j2GFTqBp3S+vOk9Y6+wgJDqk5etpYKZajmFY9r5XYoG+yGFCgzF
Z2I3So5W7CU/kflOor/Ra/0ybd4sYDBhido6obYoQimIi67sw82tVezHE6AJqMbj
eJtTy6Kmcf6BjyWh6jKk9tR3hyMloePA9L9WFkggEG+k4BKyDFBRXQCnYXXK0v7G
Oax1uw9mIR9U4eGvUSpt33Il2g9DR3grWHY8uvm2GQ2MgYWbIlRIqfzvoJVS5U5l
yEFgVV1NV9bSDSEyGTxY6R588AF/CeCMPtMA9FRNxLTs+I6WuS8vtAJ16PaIuNzs
qS7T+dnPdKOd46yC73j7smxHxwqtUUCnwKSSiG1wZYBZ8c3JA9/3tXqGGUAG0nAE
inIFMzp3bMTyTCtN4nb5JhDOHtDsUf+zETrFluJw36xTsZV32kSbQt3Nj0o72+FQ
8nb2IAlJcyuTIzFXEKWXLnAovLTigzkHQdwy4S/cBFvm1becq57GQqZgZaQsS8Fn
8IJqIMvtYzCR/iwLdXerfDswVaVHsxU/lOpSeT8xGN+FhydVl8R7LbNp7Db5d66m
gJis6k2QUp1d+psnt+NjBAwktGp0bP3aOqTNx5H+U2ReA9XLvjbCjPodLGVw05gM
iu8vixh3+DuNQdII9WVT3+BuIpTrUgPORUM+URUvr/E93utLq60G50Zn78CtzmOF
1lreSlGeKr8FIC7eAxqhIfJgCFdcon3xY3+WVQjJDRMGVONg9n9aZfZb2iODfj1b
vRV5fJcQ9wDfzOFzImJXt1AmcyGnfc0wnq4yhbnEvR3/QcbLMh7ad8fMSH47oe7N
1pXWIynZiHxR/frkFJbmd5uHPf1zFGihriSXsTIpfw1DsuVpaaP0UMvaEcF9C3X8
oLZDXzrcRRJIaRS4SSl6AIeubYK6yXh23DdszhvOy2sZsP1DXxL6SBetmpalb8v6
uFkzlMTQrv7ABQXOSkSC+znJsHsmwNFcR0czxufobCbVjyB/Ah+GGGsDMw9N1uHC
t9Q1RueO+v3bD3PdLK392PdjSYzky+yd/73aIM2zyE9ugUJy8KRrCGLPS8foSWKE
h1uiVcCX6GiQ3UPhehyEVXeiOYTfyjhmFs3KTtowH5RdM8HT/40uKIVOj/tDLX4k
MqM8uHy1cSDhmwjhevn50OD9XYm/2ZFXFqFxX+XGrFxB1DMhdjkjgEa6txLbkLTB
DJ5/EfpJ95TJG6WH8gbSFfyreOVnQ706rlH1rHh2Vr/MTjGNcocqTPKvkYpSci7f
6jpLGUnM3CGuG4bzGZ5BKKZ3cTKAD+W1id76gBA0lYMhIMSLEao+oNgDNI+L2stO
ABazds60DVjdfuR+HXLjne4Bq0205Jue6LAE0hhSi5BNtva8sYufXtohJe+Tk3Jj
KlYQTXHDZXPp3JLWunjUvjj000mxdfvylaVnNmKKVIq5JHPBamAe4YYxSQ367UND
eJaX5sAsNwx2j2xD6498zrk5AxqVOez89fgBL6BwexzCWrxFXNWx0gu31xJEqBSw
6uiLJz51SUNb1XFel+0Aj6jZALowcv3cHl15SHN9E4LGKlAUEaunmFt3FHGmvaNX
bQxyvfQ7URSW+Ya9312/aSZRQtSsoNNwhADh3UjObML/x7MZKNjT2oWbrk/Ghewm
+dB4eJ/brLh3EJaYNES6qahxhcR8wznktLOurA7XbCr29BneV3A0aept3Cp+Z0dG
wqZvqcXcl+61dtKjC1twvQ8wGSEiZD5VGFjZMF/oPC8J8msEyUkOamdCW+jRvh0d
8bFyK+6nRRM1Xo/4faNCWFi4yDDyZq8orTA9ah6xjDYiYfyaJVg17Ot4h7R4UMcN
Y3gMIlLip4ATCLRz4huikBlNevhZmxS8ouni++3xG/DHFzEhlkg2BhsddWvufNIG
6PkPNdy/eNLNReTlqCNGy6HG4eFANh5K5YfwTd+b3KA6JwphJ/PnaQoNIyjqjgDW
vcerMjZfuUmeOEiwfQomfpsj0Fx9HXl9JCtR4XJn1E4p48IjxqJU0ODwjLFp/MXY
sA/Z2U6W36r1MnjACQBxCQg+ysVBcNu/tsoHd9tqt1JINnJ8VcKlM5F0glVskIzA
IbPp49IkCu6v9qvcefyLVM9615fEiBp8t5GJlPjCJUcdsSrJ/Q6cndjNUv4qs2Jh
o0L8ZoCo3C9NPfxxaFvxhh/ahpY1P1vG7aqgaIUETkbjK9z/Xk6+nMNEm4OMM4tE
JE0jo5AMJjLyOXV1d4JHOSdnwWFW7aF7iKy3jXAaFng4NawpNQCBulbywE2/kcYt
lnbOyjxiHQhK2+bYuCxRtUTemVTwlOWciCedD9UaD7lIQaC4cB7n2dsEzUZnyvxX
lZDn4cDX5stC4pPg0UwgyJGBs8VIrVPPQqP6p2+BRAi4ByZL7qRhVyMvhjbffemB
zH+Oz/Wr//K/sLN8yChAODE3ZDUTxAfL67bd2I1VaK3tpzW/G07Z7TmxLEfBYbMK
v7yRTqlRV3XLl2wfuplOKvw355mS3Y6btOAN8BKS/X8glF4b2Ud7hOrQfsMyYMWP
i2gcbYunVy2CXRU0z9lhXdOPifqhzbjdCgLB+NEx2diuZ7cO/3lA1vQfZSooyihE
wwybhe1oOIs9G16WDtefGiIEfTynpGhyTSQEaRp+CvDgUMEz4YS+N9VArDXwKhbY
U7RrY/T2Z0oWTuaPIho/TxYchiRjVHkGUmyK+wMfrdFW1aEqIr/GI1BGYdE1i6Lx
cwypDKt1LOHt/Jik8iXha1+yW+hSkcsiX5BO5OIgL5ZgCxRzJVxMMXh4G4rgJXYp
g1xubFJKgx+T+ey5fwNGnt3IXXXgTcmpcJI/QR0MxHwcaFWJYpUc2Xi3zX2yM/i9
V85EXjZScWKQvfrQbRa1QmX9GfGXi5/FF6I9C3ljHTGV/8QngDaCknI+uJ4AwfT4
c7EmxCLg5NsuwVU67V9zYTCq1n4adbToQ9kR8vtriem9QcUB9+vcx0nD/Jo2SW9s
5i3fRWX7NVSgys4uEBAX3BZ1g74+hdftpCDZHnFuJINBhYmy4hFEXgBjmy7SvPqw
qWPDPUH2Vd/q5DnDb9K61R9rJttVJMnjOSp7dybXQ1/VnO1rTeuW1WJ3eS3eHAFT
mclQ6GLMt0cuRGQWZWlB2DsIaBbyJtCto1o73zS8++Qt33s+UVbfs7R8IMANhVKb
jNKu5U2vU6FmzlvWb7vggt4gusQPhj7YZS2emTLu8JOvPBRN5V2syrxhMrMcyLCL
AGL1vEEdlYh7MaQmI9DSr6t/opOXCMfWRoNG6Ho0Gbo8JhjboPqCfvW+GJfl6hjS
Ewu3Tfe+PjJhscHjSsa4bl+VAhnoDhhvj4PrXgGmkrnyNzyuQQoDn77UNJMDt9NX
yHO401PNARSHajM+9C6ZOfXIklBAkD2HBtQShtLYyC0vzcr+Xn4Q83AP7AaOroSs
9qLuPnwS4KOJcWZM937f94/lK3ROFWnWrRtT+lxAg0H7wd1KyDXpqO1aZrZwOASO
7Zka7TWkSCBDozqcX8S1YjFj9e5VwJdgzrcXZrTPxGYj8IBoVRmsokhUSIiBwrpe
nxOmLKQnNE6F1aJKmV5sJwlG7cdsIKnSH47lSgOLe9JX/aU0tGMw1/S9fCCxBqua
H9HDCIei+BOrQyxX6LT49hvWEcLDW9XLyNNzKWU2Wp5zpZUFGCKnzhOHLFmZpOEv
aAC+M46enOFwk9EHnPFrTb/aDiq/TSDILko9uhsjFfUYaW6zYMRSzfKFntwultug
mvg15hKkFkOIOHkgyrf/qqAXRb8npLBV8GYbOGK2ba57Ly0rXsLNIuckFrIvbQb9
+sUKd4Pt/74zTS1z9MIhVjLksFN6D/Q855IUCHGV3NmGOZDcIFJni27bmV0VCBZ0
8i3UKOIDCRLRqWljew9Rfu/MLCp2vSQppM8Bq7Wk9UcVwGb1zudt5smVzO9bapUu
ZngqG/0NCZ0eaPWLwHj1F+OXhflpiRCtlB/ZeD+CjZzolOnsS8mhNyvW0StDXL83
mRmfTa3E++RT0y+UBYqMbQ7yL7eC+0aaFjcQphGi5/zlr7iH9wXpOVGiyg8FJbZm
+/tApAy1bWXPTw4XtQeMsoKhNnzuqjCsc+FHFYvASDzXJmBrYjYYMVXI1Q2n8zBz
N3oQk7yzW3PYpaf40z2hDnSE1mAiY8Mp7l240ggR0rWVRFOtd+S3bU9LA51xwpNK
SOyM+HRvnAyCr/O7iujAoohd6LOAzejqktr8xBLOJ6UB22RMrucazCV8j3XagBsi
x+g6tFXavcVZ3jvnwN/5Yg3lCK0dwh4d7kRglNAynTOAh3qPaxtaMNX0ewMafGZV
iRHlFbSJgjIFxh/NxR6N9xPi86QX3LV0mbw25+l+9UZolqCjeTTZkaeIsG03y3hQ
jfKSw3RhX8MuSv9z7t0TqM/SMk2C1pq7mx1y0qoH+r1IZRTxbds+WvMoPT5n3pbo
qxYhC7CiaiFnaptl61LicasBazYR3vTSMeJLqdRbaLBY0xjzM/6H47qzYR4Ruahm
LI6wcaiDCia2ckx61kngH31akYWd+u/KKJgdrN0eMHxefki2yaFqJwJHew4N/3T3
PgcxG/g0jXurAr5wj9TlkhfV1E/PsmAwb8kWATb/BmayD1BCBAbktGj/FElppxo0
V5mNw7QPk/xJlsA5AiGaPghcsy2snnwQu8lKxT2tWoA00fxwKvVwL1xs9ENDRLmz
zyLIVF/2jDLMu68Gd++oDLlD6nr3ucePT1b8Ckzba/hpJEGoonK3weiM0ZsUkhWJ
o1qoY3eioxypeTARk96HU9uvHHPSLVtQQnehcu8rVs7ppHeEVX3WPrnjDwLlWRpX
uQcYQu31iGiZQYIN3UJ2txBxxpLkAi9xpJ+ZWW1sQhHCoOFMDMPK92naJILIKorp
va2o99O15auqzzNkROhYGjARUrKLwtjZUSmH3qCFAVrLmWDvhuLvX79MNOP+pg6u
FJ3M3D/Jdis8Qim3k5tBmzyExHb5sWTx28/V+80QyWBU3P4Ey6m2I5Lsztureqkp
T6ypyKc4HvoVUxRWDMgZ1Pqk+rVckXth2ekHnnJ2XuvIh5tbpSnNvC74VokKzg3j
ZDWXIxTeQkVNH8ia6frXuP9MeR1rVd4EOjM5v4u7qaG/bCCIY28/2BlymoSI97Xm
ZdrsjQmjBBNCjJCGu6nRuPoTGI7p8KnaGylBi3TljiegCr5P8bRjDzyuEd1DV1Qv
+NJD6e6fMdvYYtnuBGw8fFZjIthjyPOm8nI1ASGNwOp5HNgchyfTGuv4PsBNViqF
4JgUzg5V/ZRXKWPAGDzUwftRDpOz2w/QYyFEmvmM3qbGxQRVS8ogoKzzAjI5u+8K
H++4aEHxz5odpTbHQUyUHBqzk/7kyKlTmUkZlXrycdJ8UFD817DU/uiWugvw6gth
vNkDSyZXY+haOE8hFbrdjt5sPQJmj7sdtH7KgumlDAuV2d+ezDElbHv9vzZ0PBB5
suHZYFkOzivZnBcOXpez+7Va/FQoOCvN152qMnD89sqZnTY0yvdv1WbIqsJGfkwa
r2mJ0B0FvANa9zIZji7evG7BQMh0m1hKKvVDUcYoi0aYPVRFBEuslznxhk3utgZN
TLyw9SAQw/5KDmX52fJ+7Azb6jRifLf47nM/n8RIfesueTdXSyo5Lh3GT6FO5Qal
EXfa03eKtfk5PAmqaKJSEoJ1T780U1EG95e4zqJcTRQZSsZPAoJpQWz7aEFgK5ho
zSKTdwqd85Y3aE1WBDoaBxu3MZuMSQRLNxRGVgDqP/e115pIkXwf8VfnVbiKWK+Y
cVRATJJmrHGN+iJeKfkV8Ee0Ur6n61OpYEhBmF6qh94ipCuyFDeOs//fJSBk84JD
A+Kz41nsVXCWVg45xc2R4vwWR2at9gkNuT7Mdqp7hwVeDs0VBqsg61Nqo3hvW72C
RQGhADJYR4mcLVzvGdkfHIV/w6A3K8gO1o6bnzuSgv2kIhMO+UVdnWooaODl1Bl6
NWZqbnFERaOmDMEVCq+1/P9Sw9IOi1ZEiOI8B9K9jgPdPMvuOyhl2ECiR8bUrklz
U7Yygc5wKYekxfxOtd07B/yGbR7DdL4PAiDD7gUALwxR5+9B8jn5UR5NgsYkGcwg
zQksQPlJqwtZIkS4/aiC52oC5PpA6TGvG/g5mIAATnLx8VeUC9EtDGvwSa1AvRUq
hn8Lw7tTWJTwnDRsM6NXd6+TOvDbEgxUXKk92t8wY9FxfVmdK86IX3dPzCeczMHD
C7l2JyZlfePGkhy6kbA3RiJdwIAZ/lDWzzr47V5O7sDn8WVDgNdjpiD9twebpZfZ
ZZYUf4z7b1beoY2Pej8y4v05El0NyJ6FD7aW02iHDDZZ0cDhhiDrPN2ITDozvill
Fqj7Stwd7qBdmDaUvsthPM9P6rlvNa/EY6/fW4ic7+cOT+0u4l7kSqFyMgNoeVWO
fe0dgPkhivFCS9nvt2yYIq46eOJZW+lVcHN+hRt+gj85Je3kNWwekEdvqy4+Bptp
g4+GMOooF9Duxb1kBWeT7OnY0Dd6mYEoB3TMAerO3nmko+us8Purq90j1eEZ/mLK
0dOtWzicX/6eU03Du8oSIwFMu8N/dRiEo0dF4n7nkLj+oPrq6KY9cNQ9cMs8Ydyc
iRSXtfaqsszT/aN1D2uvnWr+zt/itzxMlU6nmf0jaePYf7Ql3ajUl4wo5U2GLFnE
suVNQvYYcw+3zzpXfNdxKesK9gSxEaT7BP+O1DoLnDc5Vz2889Qlmck9XHZUJOE5
wLIXXwLCid8SFPi3Sq3xshWydAFF2Xuo4l/o0d2JW6HEurrvxFccHP0SLJsXtCH4
HQT1DY1hPImhmucnuqxC2gpuRc7q5vyQKATRrpkT7nvl7mjyhpjZEkNiWXA4nTjk
MDpSFqlWdIMlMFXrA7nN96/ovFwpML2JxfDUNiWyrA37pGJwD3+WyXVdU9l1r7k0
/229eu0UcCPVM0n5U/IQlszxOt+wtgjC4BTxDCZXvnF2AulQ8iO7d5Stacb7gr0N
UclpMnR/H690iUEraRo6+g3anV15kfgzbqYejksfQGmnbnJD1ZWDxYWdXfqQew1o
6BRrt1qGnGcbyQExFS63J/iS62AB7rKUWihoNRf0Z5vdZoPDz1eM3/XFFKsH1AVX
G4z6tkigusdH0dr2dwcYLYsc6woYfahWp3Sh76V5GX1HyZw8n9Kmz/SqRaI/hPIT
uGa6Z+tEjADCASt7lL3qvB7ikfIGxyy+M2GQd7U/1tRGJNigzFgFGwunlZURoW7g
/eFFAHiToN3/8e4f8p+LA1hg7HN1QhjMo9qnIfOX8BXpKVpfl0Hvxj6jwqfaXSeo
+22iNUL5D8ekTkW6mYbFMTU4etwAfZwxLO5n3pamaBbVsNx+KCZ7tP2NzaBbQEvp
puAeSKp5SxwElR6b8aSfGyLmEmmIBxa1gjxzeBbcj2mJdSMpRq1bFgTFsF0w/Rob
zAix07J1Yx7h3guVwYg2JM2nDsBDPFfG0gLWmyBGbaMRPRB4xSO4BCoNqgFZi815
vPNH/we7JW7CZpOPk14HsvDZC6snAqHKCW8OBNqGeInsRmNnidB5zLu5Iwcx526V
fnPX/+oL2gbPrNiOvtaVxHBAZYk1CePRBVpzu9O/0r3dTmT5/DDIKCJHymc+5pw6
CRpMmw5JfopslSrWcHZ80yYGsimrEympTMDG69CXY5L7nQIE+LPg/E+1eRFcqZmk
xACeokw5Z8fPSHKE6Uw+KIcDua2FzgqlPmkaDzcoGMCF8zMJiY+m4sQ240jTx70a
tznDLvn0//YInYkvXLS8WI1jCNn0c3nxN1O+KQ/PiPDD6/KbFG4bH3LZuiyk93D3
Oq+4YLOitWbOlOUFyEpVyJG5x2CVgBU99h8anF06Lfb5S+9cgnuB1vmoddNIp+VW
uAstTIHdQwbtjhAwaMbPd7oUBSovvpdvNeNozeSx3n9CoeIN0VqZnTrsyeDtshnj
uAXpu2Rz9dsKHWPFvutVbDMDE51BLwbmaznzZGoCojVBXjx/Ust+3D6xgYyS0Xq0
c+SE6aysbge6o4oVCMwsdTy9XCFQms7O9YWm7seloONOUld++ckgealseS3CwIur
rkuYB2J4YrwBDsfSb41d33G4TqC6Ixyz1UyTsX21iNmJ9hkTas9jNznByIeZ9aWV
j8P63baQ+JaAnjxqDFvDFrGVjtu/O/lIV1I+iynmSlvJ06/rlheIl190k2yxTozW
mOCre2g/k8xMZzStESd0Sy75xJVNVlvBRhhHusN3DxuGmzaKsy5A6cSXxU4KV+VG
1ggfUmk6lDP6QwzdKcgO+5CxwjZVDxEvPXpbxz1xdG2acqZUPN0BoXZF5EV4IotQ
XUweMp0M3o6Ug57nTTnnQ4dIxe9w1XFAKyndzEr22qxWkGjdbBWaxLtSaLhlo+JC
3gwAjj9kQOvbQ/szn0rcVVRU9btoCKejVviZT9xmgpaNMfcRVvYhpqcQfw4brPNk
qUf2jidZDdCYgQjiiM5y6EB4//Jl5zvT0m3Q1VSMx6cbgBQ11gYnbhfLZCy3SggI
x6DO0HD4iEMSIboiGYp9NbvSrEXgvY3kDusOAv+ysGSsRjDzU0tHiRbOgTVfKYWf
L8AB9C9t/4n/2bKTL/2S1GVpsr4SEobYxTuanN8vNdfyaLRVOHFgwnZSTi+n5pHb
qOjF1DigaxfH8PdErSnfZFQcHjsLZVuRZRwlyDRa5xqTCrMxTFAZvSWqqdLB62nw
nVrkq4O6cOnDuZDUufCL4tRIOPCDElAJ7V0+sGKofxSzOBh/RdIZ87hpf9Mn08Ek
V2RCZINoKytCADSedfuXskBAKm4iAzn38rt0NsV/cZ0VNBJtsjzB/4hsTrKxB6XE
afxlgmZaDM/PpRWOIiEkpyrQFG9Erul/T9feqdwu7RGURnDhKQDb6sjj+WD725jO
rRexYhzoZALjH5t0vfwFKLhzi+m1x2qZTKwIqufURiv+P6wXrxvBgwFBX8pZQg19
NahsdCfX4IHIR7pa9mrEgnOz7txq6pJXUT7dlbKAuWu2xm5Qz5Nui/dqSWXaVJQG
sCFVwoCOgroBOnzXXvpl6iiJldoGHspAAHjqAo5a2sBoHeMB1BDG0gSA2ORypCg+
gOw9cvF0eXmJBDIl7bsK64FjWKbij6+3WCia+QD2yOKeDV5GR0Opwr85ZnUzpULh
+Pt0bs0eHJN+QYBGjpfU+37eqrFUNVcZIB9IxcAodfSQYcTkaD3pK4oXIvl8cqIw
GXVFr3vwMA65ANiwfLh3pQ7DNdkfbTX9Q27XqQ5A1m/iAiggSRnGsmQOgJdvzkak
k0JGYoluuc2nPD4roUAcVyTM8d35SWNgq7S1o+n0pgbzXoieCleF0dHuFm54JEze
ypWXM47w/2UKXF0Vy0u57EZpJCvIbNPK2/voBvRbsfOrKLghvpSCC3ei4Vii3G5f
iieE/MgqnU/BuNmpknyftdXhyo2bzgSrQrgnRuumDtXTl6lOKrLg2QfXmoIpjj3D
cVd6SzXRSsiJdsMsVb/ukdWp2H4JD3JGx+zBGnKBjGIxYXHi+r8zxljH7rvpC+nN
LbZy4a89yDkkyAqpLF5OOdSLb3K9+qXt+JVJdC/8P98qTIcxJIWvrbbHJO7o9euQ
h58TnSrXLPk04dbeJIcJhtak0xrKjnvFvK5JcLv1qkHjazwIoY434NlQbUx5sKWH
4PZJsS82sRd+u1EBqH4guFGTY8Wq46vb24BHczpggVMG0srfillDj6xJoxpjd/7u
0pSU85MrFLy/oMypHcHOM3fPzZ0W4OAqGYPLMQEwFpzAZkAppvwVvSdkdv5X9Aae
ppYZl6VtWMXHDqqamU/PX/KCtUQdORyPlWvA8KcG4eNLOnYiE+XOS8Hm/DJKQdos
1iW98U584WEXY0Gz8YF3O7Q9Q/Gdhsx9QBZ7QlSRiQNDtuMFL7HgMJODUrNcY9gM
HQ3UnGH0D3ZbfSyI5+Jh/PFiOVooxJIgsjj6KDQEumBnNlracSh+t9L2H2hOYXrZ
6d52oBzg/fzi7VkmdeJLdB5pMJMGUcOPWntbmtQTGcM9j2gibOuEJf9YiJO90RIk
TePs453KugYTeY3rUDd0pkZRiXyj5cxEMBB+qb57J+hF/KuEYGyJLAmtJJ3qRyVF
+gh3nq2SUdvprYbD5BhkDLzPrK8fPXlzjTWm+DGcSV7MXyRsaKVURMsoT5LLC7vu
iblHbCIkr+eSOx8AXen+zXZWEFNV70q06LGHE5qKmKGs4ykzoSlq/Sl1H/OLqY1L
p3O+goOynE5GKdyoMm8PIMRyvgmS1zwl2IySXuzoVwy1jabJzwjCGiwzHpiApUbr
/cTRB8ZdvgjJMIS44oQiz6OmKGrwvVmr/ZVgCW+i5keS20/Nxr8VgYPQaNze6lBv
i+BKoCzfGjyBz1ldTihXUNMszU6cZz5Y/mE8z5zIvKEunj+l+613+n0yqo5YmKXS
VZWnCZAjmFOmJSylY5FEYzvU0SHPStLWgbTfUJQbqhWRnY+YPXLmws6lXegdMcGZ
tp6kbMGb3BMxmrzU38Up8WrtiIqE5yq5/M0ywK7nJGeK+sKL9BwNVXUzW7GpKXDo
8Zbs10f/+mz7LTczzqSB7ed4rTwXGoFeU7ekcfNjFGSvYoQGz7Lgqyw9mOdzAN4R
k7yhWPFLUvSm+rnlvqP4RDrX98RrjNJU4aluRfQ2dWmRzgNfLk+3G7BNIxBTyQp+
VwFJk7OpPNoBHY/K91A6OUzptlMeYBe697mj4AZlwvwFIIY5FbPUeETBbmfT98ZO
3wwzGALQIgF77xpsM0kZqOS6J7MeD1a7hXt+sQ2ONNvI44AacUOBBuAC16dbe6QL
j4OW5LDyRRfXohALI5O9cAtpMC/YH6SJt1m1PItrE6i2llua5dr6eCZrc3xK+sKz
LSpmSgExjedAUFuUPHXA1yUFM7Cwa+zkrLKL22E2RlBOBNavnosQjGPuhrNYyWZC
V4K+zTIsSSk2k9xqZdWaikKNndCvQfCpdZ5tLZiUJCWKSq3zvRBcwNnHuaTMi9lz
1IWOJwNBXjnlxGExvQzHoNLHO7flbNzv77BXa83EMcRt57EQpG0OND6HvncJLzS3
Gp0fgfrRCQESYj8WRAAYf7MK3d+CZDzHdipn2iKSOF5kBLsKpAhvRkEx0s+96cns
ivCQyDDvDmo2Q2QBwi7glX96oOj61pursJw2UiacVwmbX/HU21zGhQIKqPIEvZUH
N2G+ngadpEJo9U6ra4AJEaRvxVJFSguz0s3FVI6XqI39dxiE9Qu5y++g6shV65ls
uLE8e8LsLoJEN7goeL6d+pSOpXxvTo6zyZIAAp2xuuhyMllG9fG64DUS7/HQWYzw
wAc1lTqJiLPs90a+KrqNDd4vGdEnu3eCOoNuCXkqwzUk8qYVCF36BekxWd3Y9qor
L14sH1Ijy1FVpRVVmi9igYbzzq7PlypQ8jA0YydwAop9nnjRjRcvvBYOrHO8JACG
hkIiC2H7YOi9X6Uj1g9WgIHA/jxD2whe8fJYqBmvTetYfJSeFLR5SALaZk+z294K
BQyp1CeV+O9xhAHWnrjyg7N7WNYVTGE2cmza7x8ZGxfc3jNuJv/E0W7Xaio9xVHn
Vu6lN7K1q5yGDTWtENMV9s6j6yOrWbmHMQ19H4ucJWohVHmlbeSoN2ueW+0Ay2oD
vMN2FV8L9EiiBGrfxS3G5YQwA2Q8QwPdtTZiuHiUup+ce9gAsE08aBCTNYP2XOX5
zgqmID4i4qpcpbNdWkThloY7zvscEBbzNIhwTa1zlwhxrAiGlXx+UnvRXhqNoxN3
Jccx4+jWiGAQDD+pto9z5HmA9eYTHboWKojQ/8MxU7lOcWCCYa0XA1AU30DPwRMz
SauATPbDFKTsHpQmV0O/Bqf1ez1UzH8AIK01R5yZ/b04TQ2Zom+x444kS6h/WzoU
I8gtj16KsVA/mNhjD6CT4Y3U6/nAwoNO+qeg7E2XnijCdLWQa+db5O3+fEhDDiU0
dZLkKVrioXLwYKQJU7N8th5fTSiTJrVLEojGqIPPzJCfJ2fR/WmHg33vI6kFZpq9
v+iR7iKRxNwV1xWgDOTq/ZqVPeDcMap5jYH+JepMBjqZRdawF+MtbKqmxRwJ8QNR
KJUxzCQJQOQ2iXP9sXVKR7AleIGpIsKJTiOC6+taAF8Mk9hNtJlPpypyWkORnyIS
SN9nXSG5t4yoS5vUDJdSrP4aiz3HYPXOejb0lVcOlcOPPLtMqszSRuZnqYPs0mzX
VR9+YLfoNk0zG5DJjMhx9H90NHJp60YLtpRzj3ijA63F8AsQnuCqbqtAqXEaKYIq
vVmxEQWycfQsoegFU970QmGVRI3/mB3ALGghzTpKWVIOIQsCsIV1uXCoo9QGWTdd
U/Z8q/cL0olRdipzB7eeMoThKKYvICRDUK3neogLbOxqm1zKpHLGUZQpURjRs8ED
E9ue9mPeuYOofzylPiDmkKKliNtoNQXy4h0xsqwxQG528a7Frp7LzcwBuqGHaNHd
9X8fWOIlE/J1Pf8YcrINVCREiztwXYJd3qfCY0P7rv8yx2WDbU6MSHDhhKG+XYZ7
QY603/O/gDkaCnXIwIbZpdsfBoY7VZvq8njt3OXg3HI6S3P+tDPIABMmFKbtYoiT
OAWakSWv7wQ2qrmA5Vroy7cZSbc7XJwvcRpW4OrX4IiU5+Eq4fzJjF/jnP5P43ti
0kEdJ/7CjWlnyB4zkqfv9RuK9RGiCg6kBRz/uYMzvv+z7zJ3rSsOEUu/mDNlkbAj
2yT9u0O5ZqzA2OLhR+JsmFi+rRlKwLg8dsrg4egmFTIk69GcFyUzg7V/r45GpzT0
lZXiBKS1ZVQLY/oobg2a3jvNdkLBN7ci9MDG7/K1SDCC5qcWTuMSn/mFbYwHjf4h
yP39dit+yh7SMKObA1OUFSMm2Yb2WMmuV8BBwvIGXu6xwIFewRwcMuC0RtUlXRPr
ychgCWyleU6dtMQVQgAbY6+f8TDYzOhQ8UuhltoOT2EhoBVL++XFtgki+YWtDtSQ
oLP8jMqJaObNC4RriEUcMq1yrUQTMYw2+WQcMSXlaAtKvZ26eyh1BPqDmJBE9OxW
lupSAvHxTG+nzPOk4rkHYVFwg4nsCKU2+9vXKxyDfKsJhKB3aUuVCpwM/oUWZ2n8
265Xjh1Z4ywnOD/0Q65Sf9KjbDeMjU4W0edDzselj+JkOIdMPKrd7JLP2PTQcq47
VZBSGnGeryFttH6wul9fMA6M6FsDlPsf0SjJ49/nhwT3jZy3VSJMJscuD5tpr04K
pxtHFqCona87eXTJD5AbenrcCMTc4ZG0OhzUcCSQClmkA/4mkUaVaQfwIU8E3yXp
Wz/w5LwjqsXYUGL9VoBA1jMEIiFqprR1fdl4nKN91YklRTwXotGyo0lB8qQzp1+r
K+8cJlOvKJwH7GY8kezsNPV+9jq4fyHil9Q8hPh3AzuGGuwjyXsnuK1AqC/WQrPk
HK3gxM07QYMcIiY/1K1fBXDBuHIXJ+WsBDHZ1iU8ZQAcsD9DHta+LGpi8q/rykh3
HMCEwtMUq2Z2JTJVh4TzLV7hKwtkvJv1ytgWc40kFltlvbh5SSKDsjZ0i1pZxpp8
e/otLrVb6ny56Uy/pC776nYYUomb8xsCSkw/PevHyFnyzQwgE5xAUCr1PKTcBYY/
Sqx2CTgZcVJDVQxA57WDJLaBEaeylciJWTVFq6zf96tRHqmYs2r8k3HA7icdKNdC
zc3JZ7ev27q2B1R8b0i/eEnoROppU0iNdGETrSJGyJSgyRlSP7/h2zkajLBRYb3v
Impez78v5EirSk2AemHhyqfHjKmbIrF3WCTRbUqDtpT0pD9tbbuOBJDXdxnHTddb
hJ3EIxchY4KY6UXaZIE3SKp+h8JmqYrEehCS/v2lel3Q45o1PpdPAk0z2hgWg1nb
4qYDZk826/USiNvjRbiZwgqGe62OI3Qv9Bu+1/ny0rvCMrdnUeAW2OZK5HUcv9qx
IVjdl4IcW17wu9U63ph82/srbtWtm76dPCizlh2az55lvKTlE2ZUUjh6AIyjvn6z
6Wr6hu/w4ZKgtSsJdqEKNftoYN8/YUzxu1tJvRCqKT+SOFZfC+ZAMitXhVDuxQhW
UEzmJQ+qQn6D6YwYSjnsAcy+isVsno0D+kpPT1ck4ahDFUKWUjdpSU4ityRFMsPp
2WRTvrK9Gzh4o+3MH9yNWfcVys2yt49bug0WkzHnfw59wA8R5ye7HpwP8vM6gxRQ
cRAyUa9H/b7RNwLvVS4hGob6XzGXvKBvUOVlrqajGytiJyk3evqmx2sHBnDcg7YX
AhzqLsvajhDC6YuyJz8mF1CczsPMimXugk4yvDqSh0C7CFP8+fpqYA5tiWLfHAHE
0nA23HCBLLin2AiKHL+/UdWix0CRSVJwYmnr18XJ71/92MEWgQaYGvgNcuvww1XC
j50KnlPYMznhwZzuUCrgKaoneEtrgbV+mw1IB8zt7sLB+MOINh9kpSQBcUbso4kj
la8sxvL8taH3Z3mVXlk5HjoUgj5kxD8BllHe5eRbk4f65RvgZ1ucAk3fKUca9Q5f
Nl14XtoDwM/lIVfo3oKxHRiVdg9CL73j5OzQw1zhdzvKIzOoObdTZvSbXW09YTC2
mKm+vx2i07MKYYf994yV4CzptRtze9UFuJGj9KKagJVBZ/tV5YzOoNzz64LpBbtG
LfdHBTDROR/8pw3hIa5zZ7OPcNg/9NX+ynHloKLR6okwcv1ccyMTwpzeYzOBV6G5
QAuPGS50X9QUZa1+NrPFg83kD62JU6F55LNRWauOiNXMB4T7e6nf+/WFzZYkOzQv
TZ7vL92Uw+ttjQhS/LhBdxK6YSxzRO40dezI2o8T3Ro6kyq+RDdRmssD3+q7bU8/
alCpgrB4OG6ITZbvS1dWHO40+Aiy0i3cVX7hsw60qJOyPhgKBbrpddyhLtM9LpJK
ZpcPQ5KK0QCcAFxdjHcP5hyfT9qHW93FkanwMTpVYzSlMeV32XMvaaQ/JvmTwmqC
eZ7KD5VxR15BkaZC/Y3xZjqavP2fmbDpSNAhxuHqzT+ucaskFS6NkyXI4/Ut3/oG
bXMDksXN7v6+WZwNb1+2l+xNQ2CvFo+c3TBGIeCOQnJPdN6BWTeH04tzn8zJfjhs
SdIjZoR3/6oIRFq/LElWLVuJ72526ODVzWgoI6qT0HwCcTRD9xdzdm/pJYRqGQbX
U8mr45dYIEoJKIIwFr/yMi3am/dEI15I2OlghOooXrtSJ0I/rpbmri3YL9+TpyQq
hpxkJi3+E6wY75VQpnF84TiV62Zz2kW1ucsOV3bsF9CFE8QwsG7mtntHNDXHIHPG
etF7aOxmHLfJz4TzKXl86d0pKUU0M1ABmjIncMwmxEDMthTT0D43zVeNFkQuPa7g
2K8LaIvZzuHPgBS/s2ayjdp2VOawUkmsVetoi/xxqMrDALWuGYTiaYss+n28mEKD
mmDMIn7jzUyU7tYqWcrzojUB0zhz+t52BKs4mkVH5DeBpaKmwG43d4ctW37OAbL7
OB/m+PwFck+h/hnTPhs6oNP3OhAhpkKYkoSWEBKVlM+D0k3gdOU/rAsy8e4R0YZn
kyU6M8S5q4Mk414qOSQZuJgdeFi87wQGYM9mFHPEKHV2zbekQVHop4ruoYsOOaB0
RZgFMi9rdHHsyuYAw0JvhAekQq3/CLRfSytO5wYenodk84NS+/L1ZWVDXuzMnR4f
MhFcTG79HwqHPMUOLcH6LyvBTnbjms2ics9xLOEzkZZEFHY2mWSYHK0rwraqnQlZ
fobEvmlzAWHBV85ySd5NOjIeT+cdVzhp/UukjkGUxzpf7r+sTIYqitca1iRPILUr
1d94+qOB72YWSFnNEes5sNyTQB6DHY5dvib4WaKrR2x2qNr8vyZXRoctST9p9uSY
GAk9wUTVgmI3bEhFeWio4RUsIUZ68QWfuLDGaYGxwjY420nHM4t9nwndo5x86tkg
wRyIFmAdLke4CbcrKzRF/Cyq4tnQBQk8fTXyuG4fjbZykGIOeHRoLuFx+gbTIEyz
0gaHJyqm2Xiy8LMjDN1RpBJjS2LK0CRgjz1L2yMCOZ/tV2s+kX01hZpV+JLzb0v1
maiKFFNxhcDrg8s3JxhuSL7KL0eZaMFQ/k/OO0dXXUg6+EXTX83afi9WiZEVy02Q
DmEDBVyf1Rk7sMjKarEawfUt50ufgCriUlnSRXxIQk5xu6A9UfgqfrRNvpXYvcQM
ebtzYFh0o3XmBiAGfg6El1SGrEdXqqRNgny7WqoNPYq5UZF49C0wUcs48FnSUofF
KiFvKnFNy/km3A7iGyVdaIAkuBiJV67mbd8KF0nqV2VZF0MENhGg7Mn5G9SgvLBk
hbsfXfAdg6YWYrk7gXf6QCV+NHoHDtZIj5Afj6gBVdffZLAfA+Xg/Bt+fWgDa9Su
8eSAtEF/KhRO8aVtwXGcVYcSoQjMvAJLk6p30q8FSvUiPCgrNI7FKyktyb/YIo/m
UB60tmhGzrbK4u+dGGXvpVeUVHiF9HCqPHrBG4EJXVQEnB9tuR9NYA1CsYreY9hP
yXWvFXGsc1ToX7RBcMSjKOSVYITFQaATuVbzwOoUysRrPiABxRZ4BiFOVsubyWTd
i5NLoG968YA36ej0f2YB1ibt/Na26I1XpJxCKOiye5Xib6/BfTMf4c+SFLRCsscd
VVqQly3oLRmjC4MKUNEa4Hok36x1Ua7lOU/U7LgKnU/VGU7OwecvhVrK6/P4FLo+
mBAEhATqNfuxXq7q+EEs9SMn5DaczeYXFADEmZVGwmDxcID9faLKwkTstbPT9Kzl
OQ1V9bBJYxFocF+64Z1uyNDev2S0gUu7KDYRl2zQ/SIWIBhAw4ytf3eqjczsjxrT
WEFBKky+6tnYrkp/5fseRHlCxqdet5PrU1vBHJ5DITTj/LO4WQcUjB/pYIDLtPsk
JeDgvommyDekgGpf6yX1IgOap3Hb2G+dPQiB5VJhGL7E8644/1U8uYVv0Vvht5tn
gfJ0MxS8mqpDoBqhBsF9mHhi3Ty+x6fwxl0hKjO1LJLxLB0CZQxJReoCajn7ka7c
KZc4SQHG8GP5P93Iu9yWm5Fgy/WgdmnHz50TunccV+9fvECLq92W+6F8lbdhRcgg
Zh5C4W7pzQoBIpuwRUKMZQ1tqQNEpPB7Jnvp+Hbs1LpNXC/VYPy6eOEMz6HAwJdX
xtGRwwNOPj8DEBxypzNJo7KrQxduHoXUs/DS8fKaEJCL28Uhz5LMCQ10T1H8KflU
t6TaimdZRXqcuv3PEMFo6c2Tlhff3PhWtonIaPWz9GY7VXAb8uSIHgix50ZfIXcB
IoxZdyItUFrjm/63TgXoDOiOaKfEdxLMZxS6PVlaFOCICH00j2qvujhZx/zFx2CK
wlOQXJEKW/7jkbllwd+O8a858UeDw9X30TCB+5PWvbobiR6KaYTG3gaI5nNKrAGP
Olb6jqfcXFoELLvLBYpuSmi+a4hsTWe/Zjv5qeVxLAUNYsWKb6QPrOdy8T7vkLbv
F1uiy5Kfs2hAcCRidLpeFWRWIoPtp3JRv5Etqw0Owzpu10ORHad5NGu5cy9ocUeT
GpL90TVvkH/uMTc0qyhUMEytpWcEUsBj+L/hT5uIbi6lNxo4wB02CVAri0K6nbHy
DW3YAOPsM/75jgx+81qqKKH4Kshc8FbNZ6p6MrOvGvsk39mm6myljwPHAPTbDNtl
rKAA7huVziB5vmrwcfrXrk7yYYgKFaSNu8lgshsVYySnyfEnClyNisXq+mobDxVs
hSRSRY8tGz7rY4jP79rEhZBU2bZ3DSlJdtSZ5BhE0rQGXosEFDZRvTKebrJiiHP0
Xjc8BY3YxRGXpzoWGtiXry4XgnIZh7UVc1MBHpEA8vxEQtcYihBWgpj3yFL9rnNW
OCoQ7DuqRQDiKv5K9ZTdE5pWwAKS5CxNI1UPArJy4FCr/gIAWJlVI2nH4qqMKacr
MfOtqyLbYdG5eVE/FvQ+xFfhlVX7axeUDCLJlRaOh7TY8ilo79wyNP3IvPpcJMcH
OOEnA0cIna0daKdtASfewlQU43c0EIBt8cxfmdnqTbsgznQxfNFG/ovA1lEwxJiy
hF0VbijH3CJp1uYzgwcAy0W/tLWFh4CPT+n7ltcv9KGXjjs36jqyFoQrt8GtBPvb
+9N2n5I+x16R/53QWIFPAVCBLRVs0XawBAgud8b5SNYo+FrLrir9/S0kGkL1V98g
RtbKBjXnq3Sx1NMUIJBWxm9kFoCQy5pAuO4pcJeXs0EPnNG5C9+yn9KDMeIzY+/D
vINIGq4WbHFs3IVm3w5Ok3iTDnHEU7d8cpytHRFZAXLU7q4av+IMOAZBbfDpDj+o
bx08RZ88mjWvPeON+uQaJAorHPr4XffRmys/fRlkphaQbBfQINhmFC1hjFuHOTis
skegBL4Pb3U4t0cH34B2Joe9IFz/prYxbT2Lg0BN04ZDoIkNpeyxa99RXkP/e+g2
+X+mNIIvnRNYiYHF62GkL2d3BnTUah8RPQtf96d5axu9fr8WevzbGe/oT8umMvOM
e7D6KdQQpMdcFJvfJtdsqY76avJCLUPnopdS+NObcWW0BOBbNdeLyy7HzFaFJpLy
X7xyBpaFiHYoIAkkSuu2lRfwabaSvkCg+Hq6wq1c79ixOHBHIg3GuyuRDhFj21Cy
rWwEEqfnbVDEZTRIlWyXKrq7k6NG3YkrQwrk3Mbi8lOm/4GW0mU6XwK+yHkkWt6v
P2gD5Rd+vT286zQKe3rUGJlkxd+Bm/SfUggl319Qn24kI1gTuasU1saScUOoCkKu
bNfi46mHzjPuGnNYoBlLodD/BsRDeZZdbFO4qJ2I2tNU1BfT/Ixvd4IIVUPQinqQ
WL9N0TFuyraUq6Tzjxp+j9AA9w/kBSyY+vGwhBjmotSV0Rt87JEVr0o6vHckpTAS
RTFIUjgojQTkbl8t+xuzm8EwN63iAZs39Ud+vgCGJXCGATvEqWUuTX8hDSySaxub
xdxy8jUtn/Yk13iIQos+iXTfgR2x9nkeW91uNiuJQBVNZysQt6IBFp6Gi2w0nMAC
Q2R4GJGnf10Cea2zoIsfmeSJ0To1+UqFdrD1gYRBUZnPpdAaZGo4nCXatagS7LdC
+JUwlfK7+MSKN9uPNDcyqxBSXwOZLLNdcVJu9uvGV36ULiaXZR6BJaPawhgoE1xo
doy6yu8Sk5xJbPxo3dvySmG9CWZPVPRDpjQcDdsv5oqJ7bgR2PN8edWZBlu/y+f/
AhghKCxBhdEVx6sAns2UXinFLJp4I8w/P5ec5yMrELoSL1qOle1kKyHviaVI+sgy
/485zOj+bH8/v+to8odqQjLJt4YwD/DfrsRJChF/vaqAUYksStd7qKpFV5SlilQc
nXxokSBXawGTGJ+dx4WJjZ0LkloVUV+6CxQqBUroBUQLIPkleLaCwZmAzNgSnUbU
LyoATVlGw0mi5ygOl6oCF3U6//Q0gZ1N250nCtJIRGIuTxWjenThvzbPIRHNJe9D
s7z4/J3t+o8NltaE1yZMvZugirACjsIPJllXWmZv2v7hrLhU/OruSr3hHFj0vsu8
w2K2k1jLbmce9d33MwokfOguGrbVdYaA/++ZG3qugHFoY1IBw6QpGJdxzN6vr17s
acgG4n6/+EudkmxFSuInY/cYzcX9PpLjUtBH2TWscpSNcdmFzFIK8QHUjIttyH6v
C59NVmWCVMKsxupmZAu0jBtfCd8rELcxD2HHHs7bplUKxFzolnXmHczF+WBv7kvs
JM4JWWfULhp822iy4mLcPootpJlT4u45xLPD8TtwyjOQvwF7PeziUEYCR0oHw8dJ
4KMUO8AntswkhH9PzBg1JYI0vNtIy4IT2Gn4cyNwK8gvSlv6esgMWQngBP9MtUIL
Adj7/2yjHpTxiU7O8DYJpCDNCktYzfY7hHrad7MXAbGJfbnR9Sgy37HvbX/yp6CC
2DhjQSUe1AjTUD4eJSYP4vQrjH1/IS7Rpv9m3dwMTtRPhsN3y+6iUz7RpN9YuWKs
6qdpQZsCFe9qQGqi5HgWHw77ZYwGw/0PpQLwcbogMnqj63BtLqyoQ3MM+g3nLcC+
GQiZzjlRJTiHbictpP8aWvjkWzHle/qRboRUybaNHc/IwAq5JW8wGag5JfsBi7MA
vbWrOb7Pr2SDhc+OGYsXjGFu8PatTlglxJ+jadhu/6UOjSDzDL9cHYN1mRPExogX
rYJUZMoUtOI8+PlAm5EhMs8mZZeojAo0Re0Et4jBQEx7bfqcjyzmk/jyWY0skScg
QgHuEDknjsag8Yt00oXuZxuqnxVHDjmRTxMUyQJkWcpn3O5Ya632SMlMzNJb7aJs
enpYRqCo4Z0FZBFPwdhbJ72PBvaO2OiCn/V+ex8Op8Oq50Jt0qkk5umCArxggFHP
tZ4BKYRjLWgzCypHLP95Cv6pfosUgEihSyelzpsHh/s7arpY/Tcqi+JvTCMOcMGd
iNVq0YuxbL6hvTciOI+LSVqoFCDaXN91eCuDWi30xI7U2jL+C6KhhyePhR6L2wB9
+uVkZxN/E2IB5ZArIzyjvVHwSyBOKHuRAqOTBGBIjMre4lTSe36uZKzAYYQxQtDy
wtuptD2LBbmuKzSDp+6nvwnl9/jOvIpyI8MoiTj1sL4i0vmeFbRHTGakJeu7af1r
o58ABm+YIXRA447vm+yHdFTU/RExU25pxzzUh3Utea0Zb859KOdgN1Z3JNnKKLXB
GozwvWvQ+tySd6rFT7/6rYaeRZUkWwDVAJdp3R3vf6yrh1poSAVWiLesubiXU6fy
fO0+Ht85KdWRTJ8LuFsruXW7rsBtU158RoAz4q5AwvPn8RHPbZv49autHH1G3idD
Foyo6lAhyGNV1ZT2gTJHfOxGaFdk1D5QxAsrOCacblhXcgaR8UPZvVH9K0Q2NRVn
XeZFoWMkre7uKLMQUNjng0QSflZr+oWN4BlSqapmDrKJbUKkbJtMEFmDA8xZeUxk
f4228B1XdI4/J1EhjX4vZhHUnB8xT1GPhZh5EDPcGiaW+LGvcTeFacTID1xEhr9s
BApgCSRI0qXTqRX+T5qXD7ney2vPlo2hSurF88Fw+gT+IXisW9Gj96C4mLgx0WzP
z/Pq0FcIx4G7hBs6bHzuZFnUCoe/wOqCSytYmc8Cc07RzBA25+rngaDdMUwIjEwM
AlcF5oohbaUDCIfBlYlnbrTX/HZDP8B+6Fo7sAV6gxLRJh2Z6E8prJqL09i7lb6l
gCooxI/fRTaySiPYbk6PuqMzZFIrIEIb8lamGOg2ABGXNWbTO5lB8GypY1mzkI/1
3SdVM842RO2jofsMfx/n4zYe27XkxJJSJJBUMKSmgb4Y//99b0FraQh7ShDgpDLF
zPGWaUFhTmpXUGbaZP9avvElgZYmeDY+AjdK3qItv/7n5xpoWe6UoNHzoydSHrp3
3iCn8TF4IMO3kZkjPLyLrwoeX1OiO2FAy8My7N/qu0hkXgOioajFeM1MBRt+P4ew
DKxLvdZFyq4g5sQ4ENXhPROBPliomKp19G8pekQQyLzNBI/Fv+BLkofNjw7uCr+E
M7lC+huSFVja4qmWfMLtxyOrz2AKVJVLWGrIPzCBRsUa1Hhue3X4Op1XyTXemy2k
M9yac+bTYKaQ9U7fccv5UBSmE54s/XvAJW8+uOowk1gg1YJiFPdknjSYbhc2TRm9
65cgoqJasXiSsD0Nn2L/4BbO7aUCEYl8CpI/2otHtlUFVkbcQ326Bz+R7X7NE6RT
nKGUPpCz32WXzLteHU749MVk10ulv7/wNPumb5VzYxFl8wZxdJlK1XCgBboRw1Fz
tzs5wMBwcwrPS/x03d9LMVdzzdbYz1ASfZrz7nVgMpaW1V8/4JDxZ9+r7vskGDvm
QgWkAr5akIMXN3OliYlL3yCf3iHhOjkE9cekVUY4C4U8iDH0rdCG/xoy2mBKg8ut
SsHRHQlK9sIVJwDghKdp0+ZPEEPsq8GMECQrW8DaDKjXQpWeLey4b7Jgyo8lhnOb
iAoRr9DzuOaPK4sf3NZcXT0cbCPiiRF4dx87kDhH/Epfua70RWgkcwN6R1HbDkva
mlfLAN3oPCfJXH9IT2ApBtcAyGZZ1NUas4z5mMAnUqYdJELPZrrZwa6v8+eczTWF
64MV/woaQTl3D2kRReRdwPjxu+ChbDlZ2IO2dsMmkQ1n/+MUv4GrZ8VHCV2T5SbW
uY5UTcoubOy5FjDKH6JHf60Zt/ME89uEJXBzb9smt2iYEbdCRanRQJi56vd381E4
ATQhguGcYAlpjg4J8IeSd2SN3uS7rnEe6gKP8yPsiVheyd3W0Z69zupFrJLJCgib
EFGnSECF3XIiWW16CUwiUve20NnSBZPGA0ZO9zPXzHXaYPwuQXOqQlBW4Zw99+sA
a+psyBQzIz5nh4+TKs1NQiUI1QiiI0GiUCGSBvlDNJiADg0fsO9Pu91z0+P2b4o/
nMtQNpBnp7Lc8xvNLZdMqfvlSNsq9pokt45ztvYIznSlgHtzYc06usok5LpI/LjZ
jSsvnRff3VmaZeeblQYo2S1VBt86gr35ykUVYeLKY+RDh0nOZbQuyvts38wu8D7q
WNd4h3pOuEKSaO4BIoQ626xtieSBiYH1JsB2UIJThFvtTHwKy8KcqY709G7S0o6m
ZjGhPoe9Ko9z+y1GT8WJ9qwEjwj8FmsdyX1rR/8SDwbNVWmQOuFEikUjN6Cvq2fe
+jjI+gaH9Sm4hhh7EyzfTz4TRdmb8zag+STFzLOn0XHPt58Tf32k6qEkT7nnWW3L
GsVhM+cjf2EKFvmFCZJIbmsgrQ/J5sjYrMKmRB0RimZqnvmSPZ6HK8CWCEmAm3vH
3sNZWyTO1aOk2y19E2VpGV1VHyzmkgqXJqf6dQ8x/WYD1aytLeUD9QCfNjKhCtry
+lwuoQvJrCzS/14ldgXMhsj8GZrODWK8i1+cIj+Ua8LlS8r6KwJq7ZlGP/mifWUM
hZgLHb9ea6ksheQzCicdqkpGRTn9zAFa7evffqMKbPBI3536ow/C96Chi60b/9EN
K2G/szci/McFWJgwV2eUr6HMlCqIi7I9IRYwn10giysbVZwVqNcER/TPWHx58D2B
60lRFP9F0zeoh+0iBWMU69x6A6Ueyvy1TMK1LsiHDF2/zeQcpgstSzK/D8RNiKSc
u+217S/RD4QZjGIEBHIy7kHRBaUOGjeBKNdwFuW/pedQsylOWyFmI/6Rzh1RX3iC
dFBuhPZcw+UTftycOxuCa8dx7SmCO0C4DEfaAKivWZEF7pshpOnW2N4vj6HOZ2/n
FewK8zGj5FjDWc9EHpQHo020r12wgNqiE5cvoI/dz0koCMz9Ie9xHTbVyOc8tkLb
rTl50RpamrhN/yVopnXHHv01IhP4LmxXHhGiz7xfTVp5YX5X6yITAEmZcbR+hCma
4lWDqOrEI4WMwdb8+NTBUHpILc/i0vhyB8uIVF+Ia6CYqSL2jXlZ5N8qqjIogXze
W5yDw7WMFqvT+mvfMAIknhU3ZrqtkIjMHzn7Wyw5N4y2Fa6LtswieTx8Eq41eyWb
X3fOl1JUR9+H0+AwUGlrb6UQbl8PsymOdSsykHGFNnthPlCOkGDW081yPg5ViyNo
TrGasVJxzQ+k9kkWf7Dso7qqY79DYH7mfW6uZVoesH9lT4dMWEwqxbfN/BxPGEln
Zqxm6X7LJMRdPo7KJ3boKxFuLP1wL64Wy283o3FsbLqXJWEdbv2+sll2gjPmm6t1
fOoZIFXX8eVl8G26Gbqa5GiyesDAaTpjtMrC5fvt37R9GZHB8BVsaBYd3go7E0qT
0rFFtWLi+EMKh8piO4Jw3kJoOvjXKlVFdeGzwTmV1cc+YMDUFJEZOMSZ7tcWI4WI
w8AH89wzfyAAE9rlj8WpXAn9SID2s+3MiV1N1weP9EIK8/kGO1E/zH9aV5vQk93K
eRknHpvXT6MD5snMr1UQfXyFnmY/pAPrSB0ddO3pFRUXnqZiS16Qnezawo1WoN1C
PJQkyJh2s2AvgG7rELF/BJSLFJgLRsYwux209eUGmtO3WJ150DWKA2mT9WUUrJmJ
5VIyFCmEUEXdZZcSwV0FeksWD5kWcs/FxfBTbHQb/0Y3foeFYswIAYigFle7+DK1
Selw5akycn+tFPkCo9gmNwAfW/NhCGvZ95qBeiMrBDP6btvOCkxxAq2AmlSGF7L3
eOi6XfxN4Gb/2XnZyshJonHbhITiRNVj48W/lAlJFQ9GXXSYIovicnLKjdnimhUL
C1KeyFpNkQAT22fDbIf/pEIxPonMoIxfuJPNAv/wStvmIeCJOVHKhK2OkWytbeVe
tfBRCDn1d+BLrwP4ivdWm3Hb4Gf37op2lWWR0rAqmrUxcZHpSDTYS6YHo6G6Hb5n
0A+S/vZVmrLuwttPMsGk3KkXAfUYwxEC4iwTS9w/v4cm9PmJMxnW8FanTVM7Q/ns
nCMX3AT+JyuuUbOmZkG7IlTKEV9HuvvouIu0FathGNf6aV2ezMspCDo+Yu/EI873
YurMe1+Z+CdGf17OrGelAJKNjQRT1Y4U2iLVYCEcQbf0xQOHYgAwXRyXADBy14ts
V1PqjooHN7T5huUEqWjFL0f3B4IdRIavdByBrmYVlBUyANFljyFvgcKU07IlWKUk
Vmf9UU9MMl/UZmmsAM9xGSRZ1TtwvDaFGJsODaO9d4RfwEkfsFGw4i2d8MWgbBEq
GUH1FMFOoH8kE3yt1eyueuOZXonh6yGUr5mHc4izVbuiSqcW3hxMIX4kpYFYcLyK
2EhFkBelwmsSiEIr1nlzDxIgd2yr/PqhVCoOUi47V9u1skXCkAjIr0pczxjWKr5t
fBkN3dQvQU44uuY3fkZkQqz0JeNZXN2F3ADA0h+D/ab+3auajPII5OzS4R2UVc7J
8QqkNgOBsOFyYbd9jFOzDMeeK/Gx2ySdP/pnuncIkoAKWgFHq7p03aRbKBf0R54y
11DjLiNOx6gef1/pww41EWvbLplvuNTlNq1uNWgPBqY0L9mwwPPhZ6hCP2EAJGGK
id9/v4PxcbBopExPhLiN/3lg4nJBcUfsinIdDHGgFGtrHxAnhEsIjBLY6eOf9BRt
9l2Bl1qQLVcfYuE1ikihTeNn9nbbEgOISbyKilgAKy1ZmziFnwXQjRl8FVFrVWAd
nIV2L+8AG5T12MhBTKQn/3reUXSxp4ar1iGOPE9ZFvtLGBkmdphdr2DJ4qkSvV8Y
tCpHs3ph7IVTHpLQzgz8UuKprsTO/jGkaKfSlyRtJm3tSXSV5qNpJvWOX8bsYpCc
q+MsmJl7TF6wcKTvo0xgNWrBqxRVPH1ygs+aGW2AqVc+Y54rO23E3oKArtcedjEf
Vy/OvTaNNxgnYLnKsUsana1ZRUm9VkIFnwlwgtlvywsanE0xGxe8SaZucE/DOgUD
EnbAYpF+tLwtXfp/ZpVnREBYpH+syTU636MUKay3ysxOykqgkUPUuLhO/Obeph3O
meXgm67pxgD3VST7c2twZYu/EhmyrfV5k9fQJt8BWwQAnekcREBgJ3kSWvbPvlnD
YpLWcgIWtuNWBhRW/lqZN2JERSDEN2VoSYl6Csl+1FZYa9pRkk8pxPQ61cjOW8DI
d7RqEjF5aAo0xZDDazkeFFhf7BM5jUA/QXuMcpKzRHv/GqjqKz8PxBehHm+ROT8o
jesAuBsrXO2Z4TMr4cc5WiYyCRjExCQyTAEvXRQr/sN1ksqxkpV+f0bHvY6iJ/Vv
++yReCS4MqrTJSA7/1ZXLAF4E9QE7uDPjJIjQphQi3PAMI9pRw22JjFQ3zyxxKVr
4wVD0Hp2D1gb6GIprxgrEWiLd6flZ+KV92z9lPAAlp1n5UZAxu1BZkypvVAV6i0e
+oFegbJtfRh8pWUUwUcM+MR4lzU3lwPZd50VLI6ElroGkhGUedEaV/k2lDjtxTj7
6D2ZEeOexLUBP2DYrrp6ZKlFViZ7iWAViNBjHhZceS0diFzEYBi1m3DvnuXPB+Oq
TCeypFanmF+qo+qPOkxJjPNlLeX4/Dng/IPJZc2xoeRzRNLvK/BaI5UX+vdnL9e9
YtPVYCmYJ/2yfqtzdxN3tuj+dXZ2yJsdHv2SxcsUisk7pv6s6vMuKDBLKlV7YSUr
HbwX4PEAcxkvrf3/zPXzPE51kYqQ8RXMqG32jaG8/Qf5IjAKJnEdRwGGOZmtJhGq
0x2XozQglNp5Ej9yq47ZYvFvwsv7fAq6qQgi4SW77wUPSRknbsa8ri2u6+qRpr6i
J5ooMVs8USJqoC1JtupdDVFQGZ+dpG2v7pgMT79si6aWCx0Gy1+DoPv9furMlbLo
bxL2/EafSHIE/lkCCr8pyMXV6MgfPx2yZ+VYYvG+OUD1hcANwE1iwCo+NVl0sh/q
ElI9Ocl3v9d1i8YISG62j6ZUUBS/ko8wqcZ7zyWU6Q006dBH9nGV4Mk5hLQxLNxI
lguPDp864W0w1GvyPgdz61KH60xLt/CcslaDpFTxkAy1zKX5RAu6GZaO0//D2owg
nHorPG2YKzLcZrkWKLzajUusmIn+eMDX5ezvhSm9mQzidAO0DLArnYMUMU7ZTt2T
jGP4dLty39Ups59L9wFjPklm+dlvbsrAgIzwah6jlAXBjEI/Gy2T+6POpwXLlJw6
d00rXwL7cUtP5TK0yTeKi5PzjEsKKrbpwv20YzJ78A35HUPlr/EBi4MT9UPyQp0t
jVEvli2sorI9tcN7SI+76umCN/f2yWimLe5dqtHQyJpOE2GsLJQwLmVjCYDuXRrm
BXEJvonKlJqMgPqr4aMCIQvQHlzv1Z9uVNOhfexyu0C6rRuxJnfadE5Vvp8aXh6B
Uit5UuLmZ5t30fe6rotSRijaXVvA4TfjI6zHOd3XYlx6d1I7gPGCDmi/tpVqPhfi
BPL13RRWeOTUNV1d6TUPQKvXewO1W2qInthC+3mwByUy2ggZ6+bi5GJMOj88uaUF
VMZzhLmBA/Ji1J2/E22iWt3rcPhP59txFnbPeTlla32F5MaaT88LzvOq+J1U1AbO
blEeD3Q2Gc6NSdJNCVNhgGYwjjaBdIQNIyHKjTjSRaX2mE6N98xgPrZG9Yl25GQ7
8splW2SXO5A2f7uotUekcmiR7LjxEy1XO+0jLCb8QYQaWLcNcmnlTcvgb1vBfkI4
4JXXxlnAY6apHBnR6Q3PoK2pfWgsLDUnKfO7tkuV2dDnT55SVqvneE0jZclGYr1u
/G3iZxiBhmCaMy2VtGnvIG5KxwkMmA6DWJQOY2+qXliGxKLFgRVcRv5NJDDJ4Pdd
/p+9l1hyGLZCuMdr5GwPjnmREXWy0qn6favKkHIMA07/kOGp8xknfsW7t9o/grqc
41S7Ho0mOIjcf8OXfmi+0BwHQ70VEjX/9oQmRziXvgNHaCNdWy8cQkPyAqzXPHw5
3pePuysC0TXA4UyB/9SJ7Cktqu+EdDYwsiGxyfw4A79mCGWT25rqfT9E13ZZFza5
7HQRVXQ8swMYl1mPEyIQmIpys9N3evCpv6Y1sxisPN5GR5w4JR5DCF18PN2mEB2t
vuJ+OKoVagWyPe9+YuKj+uiBEryhFu4yNOOiHl+ebknD/vHD/Mk20B7ikEI8rcVl
MVpB19Jvg8oat1qmmxK8qR2G89iE4dJU1EJ2OpK7GHKHR9YDi1Iz0d0mOOHWZyU6
Rq/rt0ben/l9sFENWE29sgUiIGXyNimO2zg1k56ucZh8oSCtfXgs4E3s9xUIh1Ms
XENlU/87FXeNTNO6NxIZExrKUNLZTWUEtdZUJPAy6ciE8MBgo9DlTP1XlTVGxFoT
S1aJQkLpvs0O1DBoMQwc+PjFksBFJhtgBv04b9j+5avoBtX+e00fgWvR3azUQQVF
FFytfTuadrG59HJv768sXe9GyvlXOGNDuEv1NGB+3M87iycXuJGs47pti4BDq2vG
VzJq27Ml5NBdeRpwfRe0PbpxRib9KYUqNKWn4+X/YDq66ILqRuyf3ncxgp/gMdou
Cif82uR+aIlKJ+VyQNvp9WGkYRvAGmTLue8nSjRWb/5j3tr8o48L1COfC3drq3CI
1OhLrfIH/xMLztviphnc3tZSXXffDYzV5ywYetDyKRHIuygwxR7Dx9O2AaUmTp8j
zifK8jz+rTqeP4QO9eWymemJgAlEIBrTqu/Lx/ySD009rUCV9gNBnehbikRymrsC
ZafDQ3SpP/oSqBpF7thARRv7b5u/pjExdDlrH57vzoInIe+x5OOL6lcW4EeOSuf5
9TDWuzO4bQt3WHJZSzaJS7T/o1W7j/lMifHFbjvvY4l5Kj2me9P6sWq6zU0kbNV3
sasi4uAmzOGbLTX4dMtzQS1A1hoGEg3urMbwe+/6bXHIKjsQQV+6C/ZVYNd2pFiA
DN1OcPUnC2HGhC4LTaR1h0XxtyD+M1/uwejykgkzmCPsD+gYITwO5iWouAsghYTj
PmoaiJgtGB+xlB9/AbUSgcSz2E82M+8JbYtuJ6rOX06edKlsuYX2PCdrowD+nQJv
gA9zjLuwXWKnWJ3eMW9x/i/6b9WYOADd3MoyKNNWD7WvW4E9Xd77uZ7wVMNMTeIT
QnXtmPgMYsC3AsOXBVuKot1fcCsMBYpAXa2PR21Vscnd3Hgkk7w1sxcCRHxde5n3
t5bP4/hco8hKHn5ejtoqZs02m/HCmjemOoexK1DnXBKm9Hcoes4wvvhAeSDqom5l
lrUl7wWo5xfsgviSrBvc60RfVDN2cYRd48eVe46L5uGVumECrWIYFX1ovKmm5+P+
I8Lpt4yVseIlH+mqB6fzt2GMObZbL3qzBuSYXEG3FTqbB+MWfbfzFaQpWAuiVltO
FpSD3TDGp3+w4uh8LZCC7t8Ur8GAH98QySS2FM57NYScW4NPmf+I3wJokgSYvj4K
2bimxAqZv1DyEh7BOHDUG9Sk9gyLBICKK8i540xvJ4Fl/XWTHAzT86vekJtmuOnt
i5PO3Z3y8NZzAE9386bSWfrxkD5G94HLRtODmKOHuODBnxLWxw6VsEGLVjIjYRbe
QCW6Sc3hpTIjtq3sYpRHHqNOYQf0FNkPYUKV/jPxxcwg7ZeHqhpBKat6nhqSOw2m
oicqIr6Vg8MVnCXazyl+Jr/Q+W4NpxS0rHil1FO3yS8OSzkkCkB9BKdavwEOzIEH
EaImq0mPP3u6Ln6j2ngXHYDQApqik3bdGTkIM6P8k1Hw+1t9i+woNt7KPS3OXMn8
mKj/MzlSW+q9B6VBSnuv3L5vyxnGAECGyt6FR0sUi4QWb23xpzmducC/x7k8kshq
+dwcJlJC/hxRyCMBNOYnTl4wv/Z7QgO4UgDwJpWcmGzINAKM5I/RWav6+gGgATNe
a9H4VgI10f6vAXjRi0RhxmG0vJ2Sub4Fhn5Q421lZIFz6sFlqrbJvY+4ItD/N2bU
qfrAWs4W3ITRkni/3m0vv9AuhrNCxyKT5onk0S7LQNgmNEgfBBcNSBNEelzNvpW1
KqFFV9DGlXGACTIH3TU/trTYlTtwB5B5SgEIpoVXxgcxuFRpECbOt96Jgw+NvRAj
mgOllrtU2lTR/g233Sfgz2MXkUzKXkrW87XgPSf9Kxe+deLaqTpubH5jvKbVHIOV
R7/fn59TpJH3eoDMGFbQLErg3non5Sx3Zo/CiG5zmwJmaVXzlHIIZTR9J1yJVEhh
8gR/OsTncoWt7Mdmhuh91CHiK/7mk9Z76G/MNcQrRy0JkcBxsNmioP3jHOPf1xDx
rXR32XNGuXStFeiIDSOjEM0yeyeaCP8h6vpLXlI9bVsdJTILgm7HPJbBtlyJX52d
B5fuQ9aqaT2oSZzuaxMm5SIjFwc7LD15tm38AHFj+JRjN8IFPPM+ecfE/x5kh71W
rY7BKOEqfrHo4+0/ldLPA6uHqQUHFxr45dQMpycMdSBj/tHbS3nMRiRJWEXaEFnb
9WLeZcn3H8xV/aFZL0L6qfbN2bMDQEpz+ppAgWnKEetgC5cu2O+sXrzUikgWwpLJ
uS9S8JUehc9PWNJzRiKqXLL6bz0Xl3R6bJHemGOrCxOuCTHT9oND+ovZ0URDMPzR
McjFNPXdR2EUWuON+Z/HnJ74qjXJRtETrfQZyV38SxfF1206gsC8oHa2y1BCUQRv
G6pDtEsgK5ANw3BWNhwjUX/i0GW3Fwbg2XT3fO/psSisyaDvhPxwRERYpW6bWF2z
8B/QArhgxzCls2rtdBbj5UgxtwvKieT2I2LBjGaBRwzfPNyaSkqGxD+HsBZeou7w
yAIBAZdxL9Au4OwO/U/2aUmcvUkOuVMCialNuO+aomn2pESYWQo3+F2gzi/CFdez
XznWsmuPRRhodXcaa2+nXfJQ4lMrMWq5vrW0hB/YRfxQ0F43bOOAJh2ejfbkOtdj
jVLP/PhovIoaBRZ84ebA6w50GkB7HA4C2KWxzDaRj+8ggZANv8Hgyy+u5kAKObDO
60K8uYo3YbwAhze+uzDx+PdlEibbx1Qm0kxCacr0m0QZi7aEkCNdsyx3lB+R2lyB
Z3L89IKw19v0CKB9xiCfcjThFETu5d+Wqolx667u+1RrdfVLTkbbOpt8B46xoQMQ
JfqCgkVDvZ6iCvGyI9YY+bmu+ueRrZ4+aHnKc5/kmIrToTHNDFL9tDs/JcTO05R+
zDQpqybOGsOqzLwAIDddW+U8sGby6wRIi3s2Sgov/qXZBJvUSxiUKYqOccD9gKLH
ljd0kEUGmmmoZpKDDskbvtTSk0L+nAfPHM4hC8hQzKrLYO0xAQq0GZIvl7p5Qi9z
bbWtBzHyGmF9SXn8E8QRFX3LLeGGREUUn5iT6V+j6eNWEXbdcQx4kRzLXSlmhVxE
qd+a5uLCG444k0gnzHX0slj2twCG7ydud+15ne4panzQh6nVzKmtxC/LfpOYb7+/
ijLO2tQplUkY2JGnOkl3VgRWuvMD4ljSzZ6n1mrTnHCpP6hILT/fd8oOHaMUav5q
CshakKyJkbjhjJ5K7gUUk9yLJzwPUwaqbHYafHLJfQlechiuPSZ4jhd+CayF6058
ArnYXzTL+7zzaKgtgOV5JV9kssK9B9oOuzlOVnV9A7MmSGhzti3uhUeVJZ0Ufc6j
2SrX/C6zur2FXQYwjrnF/X2rH7jLmXa6Z4ABhLLHKr9Ua8jvZN/a21V+fEs53nj8
zdRzi4vAlV7OeAwBSP0vlg4pVj1beAEfNchdo8tyaSqxRilUHsNDFEuh+T7VfsW0
35UTFTEDBX46AGyf/Q97NzkzJm/kTPhEBh+H8OGciUyd2cfCSXlIT8INpBITygVR
d8FVTOYGWgXBG3KIPB5rLrNsAkdUD+aQpPO99J4tgCjGxZkI3jTnFRobCxq53j78
nTfaL6wvw4nUsGOJa0mjGFs4sKrvubQlfsVBK8Gs73+YOVlg4yWBhhc0xSvsCNPr
VMhFVEHyC/n2TAe3bJQn05GegSjGAlld9JqKFSR+IqToFDKFybmLGrZFZ9bc4At0
j9ADQBZd3XjvQ+pGEAoA740BU0dlpP/8hA+W3v2nl5bVKD05VNy6BmVfOqvzHu2Z
G8NFgZJS4pIGtZJ2iFljFYV+x8s9IS0o3vie3hrGZzhCO4IpYTeiQ4V5t+gpUCBA
Tks+AHRiozG1eTbf5nIjHhPNjTXbLTgg6s6k5+3LEmpDnP++dFONF3Dro9hupjgr
jNgJlHfpXGCubiUfbpVao8B1LGPuC2fuEbk+xiwDbLzbHZjv7oPeUjaE6MxiA5mQ
YRbBrlcI+VqGw5I8PMFuM+GbU21wKHOrtBf9XmH5jl35mXDGovq58gn9s5xHYSIp
aOsJSnaXJug0988oY/IDughqCQk6fbBFp4snQUuTAth2EtDEpGKhgFqdYvQ4wrxZ
SQKx66d3YWD1BgF44Uk0LJgYwd7CqC+/bWPewVTuRxUUtOemNX1lTbbGOwEFm+uD
hy87Pi0cpbn6xBNhBmglA2RBpKlBMf7rWeun7niDWgZd8E93cR7qFeI2xeuD8XI8
0C+Xrpd1wR7PIEsOAcG7PF3Gcv+JfeKHSpG+QI2ksbcXcllWg+xHYEHw3c3GoFdU
o5olRJduToFTMaik9j9mCfhTC1VzpCcd/xDu0h4Md1EM7+6F3+UI0GNQwSAFer8B
zjdzfT1Wy/Mztn7qvR/4pRkYep2jiJPTcJEa93S+aU5au1FqKf0W32L3q7CMmCXY
asoKYAqOT625LjvQOpob3Pyp8fbEervzjaZI6GCV1NmcMR8OkxBssm/Wug8e248F
CFsqVMCX1h2WlnoFQGiajT6K7Xem03rqfn9SfksvSOyjv8DPCDQMV21Vuctq2kgP
v0wY6fPUGMGxTen+2mAU73M4NGHlSj0j/ziKUM1gDLRMhTK7n3fGYgHsIyvJStIw
xp0ZaYgVg7e2ILRHVNxedZmqRGv8zvWvMAivnmGh21RjWNbmYBwNRx7VTseF2knp
bUgw3JPgVXnTO4wic5OSN3KMcR6EQR7MOBSN1bEpgDJLbqKzRu//AT0zd10hVWAq
x9iVH86EDklgMd4bzLw0SIEp20+ujxR9nB86T3/+JBTWZEFg7Od6ijtNVFmjn+Vw
3wc+6LyCwjJvBHFAbJlxqGI5jVtN61eWS6tgplGqsMcjKrzGP4FcFoA1wkRFU5Vu
pvhItzXTnkLhoHG//UqyFJJ+2HT+yD/5jYTUaHwMKSLlBlcVzmAs+FUZJeU9kkWl
IoN0tlQSGEw0b51OvhKPyM4fDq4r/3inycSXACEmiFUhOw195Jfkz50Kw9Rhctpw
kxDPotJKDOc9ZoB/a6gmiNgVWJcdC8h8o9hSMB/3KIU+RujcXFkeEeYk9kl50q1U
o0WWsAF5cUPf2XgMTx8BG44fwQzD/+rxakswl5eINF++esaFeZ2Vow0VgOwyJdqc
NBtEXquk5DoW+sSaT715DXkNPuYmqRy7Up93ZgTXjGQYpp8nOLXuXTyy+hRlN40P
0/cI+/7/+MPA/llN3CFvSGNz9XS5O6FBnmO+2svkCmgjqcP/CFxOGSZ1D/vNm0Rs
SA29v7GUd311ZsWknAh6CsjJfWkDtupWI6voTr38Sz9rEuTeDf/ge9XJWs4TGoh5
9cfzzr2OV7/fHOXXAPbDlBwW+CWl4hMy1Y90hf4uRCCiYeyf2Y9k6NkVQMTqjpo8
Clm0F2sK/+wONV3bByRihfJmoiLxWjYsmsYFb9MpNCl6syS8xF7GohryDm21jXtu
VBKDKgcHfSKzMoT3sjYTqMcDT3Cy4XtT5rcf2PT9R0sJnQ0Y/G+uR41ioUcD/y4u
OR1bIIUZTKE0RB1YEkW5Sj28eBmGiWc2a2J1tHuK0vY3g+qfHXVVTJCDxBhUO11c
gm9b5aOEbmG2Az5XFyskxLhS9wdpg1hlZNpyaUxV+x7qInk5bl1QdgNbZY3mA7cA
O26NITKmUNVaY0oChi2EMjL9AwLeMXnvDgM8QJkzhnQ+5I4YFqHJFJLu9ajEE/KL
vou0/q3oTqsv0+R1uj1qfcmety2DbuMDiyTGi3ujC3K6mEOh82fFEzOxXWNs9eCa
0n5to7rNJoUz+g13PJyNvaH7uSFbvUraf5CUb5bxdJQzU80XcCohBwAhXqc+2Fxs
SoOzi/2098Km6Aci6SEeekCfER0dBDJmfhEdxvCMg8f8b7zdeYuRP30xcH3P+ZN7
GVDWOkHKOchkbUDDGVxXEP5/z9HkmovqTH5xSJoVRaNOWNXRCwpmeclwX68T649d
3W9J5e+KEv1vgFBw2Emb7kTbmoZjKr0U4QI+copcTA2qvit05B4zOIE4o8/g87Ty
HGxY5AL888jKbdtLSO43Rx0Z4U+1Tp8TeGTSsfk6cqMJ/2jjf0Q7KBen/XIQnK0g
L29dR9ZvxjX6auucq2BPuQ6JePVROhadVj6w0B0axPlaG3P1TfcUbYufwWP/jotE
eBIlrbL+42q8FeyVqyMEwpz5xn6xTLgsFryXaueIixNOJRJSSyxGXG+KdbClXRo5
zt5oFiI2ovNrtXJNT1YS4uls+OTZD6+QvzJV73xlR2qd/qnw5wqUDjUZTbk0xTux
z6NMP1aVaRNiF5e03R8kdEd8bYQQxPBRT7a7tNTuG5v1XUi0Mt3lU9BT276sz9Ml
/nH1vzeqFqadfJ2MgCLtyJv/Q3fiqv7fsFwlSz34QHtCZgvi7LyfCw4QsBlkbC5p
eBZTz+vTjORSowUTChgSiCVCMOFwgmuX2tbiIHILw8JKQQ8Tni6PTcSea0SStiAD
/gnTmwZ7pmPGzS9+eYoNbFhcTXh5D8N6duLLr9FMj7YBDkOKnrOAqz4K16i5+5CE
F7PWVlRBKeOSws4/SBRXSNov9VFL7a8nKZkmaDLGAvldbeonp6fUFZIXqezoSheW
6eeHgiabiE4CLR9urihOHhP/fZtm932sWxWP1Gt/JdZAb3SqxvDWJqw69rXu2/NY
V51SlBhXrGZapor9tGP21nCUuWDFEcZfkFABOL/D+7Av6rvL/FoNlnpMmVm5uKJU
NebI8Yon7UUAmbqs5cIPZPcCZ6Buy8JrqlUUuKF8cmxsEpit71ommSKQ+++D7Wcw
JuXrRzBZkaWPN9w5yfk8NG75RTcTRXUfx5iPN4OvxUFKNNJEMyT42sOKYpDZA3r1
DYMK/eRmMBACdRo1bP1Y397XQvF4tByLxH0Es3dazet1InolrGVLwT5oSrLR9CUr
oE6ZPkzctwGrKoYlnna74qYx9/vda/pQ9N4tGZ38Y0fnBOPC8fuMS06D8MIpbvOQ
iD9VRf5XEfO5lPBHtEmlfTWaqxkgKukqdm0YbcnJRWl90xzJlo6R60yy3huVE/AO
XEi9IPak+ei5FxGHqtEzNPRT2OGyqZrAk1FL1E4CNP5jZTF/zTywidHwTb7/X+kj
8AG8J6xCyJr5NRCbI8Xw0+6e0Gn09/v6cRWiMyS1iAleB5tTa0rIrEVsa2QLjF55
tbk6Xc71lHC6AXeJ/7y55uZhTSihiHRGrK/RP7RjfujtXL6DjrPN2CoWZGMNL8X5
fdbhELPCxCcX2ps3hM7TPgSmY8PL+ZLAP52VdhlTVr+aC0dEVglLYjQl1LNcyeFc
rjPDU4Pa78pFeFRuTPcsd9VPdgO7QdK8PEU3HuWUCr4m1d/ny3tLDuwXZywe1Xew
lnXPB6xGYlGOKIA56dy588HDuAOIjT5SXrWpi2Pr4v7KXrn2W8IpTIGikEInKs4p
Z6+VO/hrpTNNBnLjRxZBZZVIlDrfEdzg5ssArMXqmG3s0pBtvlfB7UkZheFC4gaM
AvDCVKMCKf7O3MyT88gfkCG/UqnFmPOwEg5x5ibsjpDdB8NVm/CsYgYvF1QoUce2
wyobyW0rS/A6V8UvOJCQZxe7+F/zGWngi0mudM3hNk8q89+DVk5PY791WsfJCaT6
4Z6XlTzNoozTK3yWOdpKEhizLGejEQr4JRoITEPGK+AIgMwcu5dfhVkgM0B7m+r2
jx/+UV4FxhwrSl16TQCtjXTZ+Dg4I3Vl8N0ZZ2qtA+4drv6MKUqJuEOtpoC5LNGv
kKH7KP1v4v6OXUPmO82Gli0nXuLV3DzjoiHNyEDdkz+R2gGq2EC0dqdkEz6zBQ3B
PFX+urWCDvMuzHdWHKiqd8XxOqPxktnl7a4uN4L6Dai5KhtaZmAMPJMQ7M/3yLy9
djNPhttmfSPrPIOBqQfgSiyBFo2nNZF3aw17Te1H+0VD65NfKN/2oTaOSgO4Q7Gh
8exPsK1au4pCw3iJMCtXR1xEkEHDKw0iEl6bIBx8IaxJbQONuv4VbhqUmdL5TZMl
gy2shpvfpvGQukmymMDCVHjiyUF+3ULaFjBAqNevRhUK5fZRdr8SRnuvo5CmhlOw
x3AbF8u16CQ+ubIG5HriEeBnPElSC7vciWbFPFPgl+JA4SmD6JYz3jRgIel3cung
1DEKldvwXWPtFJKWXRNqsqs7O9PFI0zyhd1ASmgxPMgjxBbxIyspJz+rg4c3YBv2
rpj8rZRrQuXBKRuamlxzhTUa/UZt/O8j5e8PK70fDoRMZugtrEEvZA+fVYJtlObC
ZmpgAyUf1RVLJa72ESaT3/K9wrKL+3xrXJ+LhfkPRplCS1YTNfi6K8Fp3o0fkj6A
n8QLv7MhC8BWYk8QtIXA8GGA6S6sDylWUUgdsMt09omO0mzqxlGHzvhu0lay+W+/
OcroaovxC0YoreCNHtXeoIKGWxruLFSonxTHn/jybICIEarFuQQL0gtmf9PiovIt
FYDjeRczoJauG7Wo/Dg9k11tk6fRhtEm/CuGnav3MILyBmyB/rS+6uwkxhYNjCLZ
s+ghI1LE8DVp9Dmaobl/Nh2wtzPT0FQUTx+8d1vtT1OQ2pArhMImJvhBRsY1f8r9
kxs+VkmQcdXetYsZNvIuVlkAYiQcNAlsO+Hd52xPDKvoQxQmSKfcNQu9t29L80wN
/fcWoS3I8oamRJZbm/lsR8byh/6d1lk4CgqqALKIR4Sw2CVjtAX/oG16Y8Sr7/nO
tunBknFojUzym8aUVKCAnuQIdVjL5nDLvnPZcHrF1jFG0Vxc+njUOmDLi7thEe6v
aa7fRtXvc7LcadJK8qHpDx2xnkghtjg0668L/3eSYZcNHy1yew+dOg3MNp/1u6Lo
fj1VTK2P4wamLxn5G0BzQ7LiUwTsVfIphJRUNL8rgGQzYwel+S/Ycs0dsiBBW6PW
vXdgVwIF9lRcbPJ4Svsbj3kg/fQWJBXs5BYzZFr5cSLP2NSfsu+LP+59O5Abxo1l
uJLk8K4AyIb3pZtxH7BDZpJz63ClmBzl0TgYWi64nmGjpqA/dyW8Ud9obCDRWWwY
hiPbdY6mhK/kaCrSUE0YUtnSfKQ4qXmbczgAlMrvhnyduVao6sMAxDB3GEMh4Vee
Z8RAXZSXK0SdfX3CQHLimG7anuY1AHgIrQxBtwGyu5Gl6SqJ2BGuWnWlYqYPmjyD
xvh8cqMFNuSozTbPooRQE4ShNRUoVzow8HfYEkwuuCJuAOALWQpba+YSZg6HaKGv
5Rj9imVJMMvDvEyIeGrKi2zsdmfbN3fcT7LdybXxG9RCgUD7j7ae5aUeHWyY78h1
XGCMgENFbTRe/xR5dI9hbTuUZaordwBzp7kCH5LPEEJMYZPnAsm9Ov9T+vN/NKAK
NqTnlQsciw7a8ws/7R9zNYEne7RKaKfZ3Ez2af4nVoaK/A2Gi7LV5qZ9yoyrckf/
X2jvs/M0J5xucpcP/NKIubPGQRSnHsccuwjlKb2jRLRDVajfQ8EKfUh0/vRWPgTH
IW9nqW8/PQrePSO0QMyoEl/FdcapB6C1VNumO6Z+ZfDPyNr2cDMevkwFcwtnraXS
TM1G3KuTejGxmAqoM+LwJ6sG8rAUlPj9CT83lEpq9GrimjADBJHfYoI3cd6S/MFJ
YavoDoItLuO25tQm84K1ZqRAQBieYlO9UT3ZskOPJYUlNsJWvT4u/6tzLWI1EOdg
hDAwbyakwDugPBNif1+NyZTdTsQ3fsZfqyoTLvJjCdvFHbWy/+JCDZpl/Mgj9fjM
jjvVa6Ue0LodKxiwzzFzXAYqjtcZra4+mVgPUDPIAvmXFFx/2+07ki73DpOhn/t4
K5aofrSWzXzAsGZMc8JVmpPTeIzP1O5zBjLUx8eQiswsb1hipggr8icFNRQaPWLR
YRl5psAz7l8+1w8BRUx2mUiQdTFDbM1pSP9LmxCY8DtS0q+e+qJ+mrM6y1d+3gND
/vn5CH6vfMIcrFe60e86C90I+DcLOLB7TX3LKRIHpqMEqrzMz0mqqEFWZHHIhLS0
9+Gylsj54z9txn6T01RUGUL0sOsBnXI2zpqK6w6TK++b6ECGxEwMtO+M6AUoptuu
DPW+kdzPIJWRoP9TftAUVTM/oGZ7lVQpnTgXWKqDcCcwSiWDvbGGbUoi+ckpuJQB
19/h+FTuxEBCwbHMtCplKl4I52R5dM0GgXFw8IXVv9yT1sbubzcvrB5+jromkMAt
bCYbFa82t1dgj3fTgVm98p8tfSDdorFc23JxR3t7X2HXWkZKwMcXfqjkIp6mKujC
9jMKcxbQ+IBMKDIDuFWfyPe1lHYBME/akNchdlY0fhA+/aEmliBjWqqgVUxk0JfA
b8UnEwuupIH3JlN+didSPrUmogEbxZCMH3SdLxupKEbeaPC4Z+TkL2yCmMMWCRnf
bEzIU0b2RCYRjhAjQXrO5shZBU+l9UtClEyG3ovtKs6UwUd7j9x8Ju3cVCN6I16e
BKkYPOnzmc3jPgPP0Y7v2PXm4jZF5QggtibwKdDtU0CdyI0NSSnIy2nFDvZ7VY9H
+pKpM8JyQ+/O7hoX/YMSrXFGgbFnAD7E/FLQ1I/dyp80RRXsPCdIuYWioFqpormi
7YW1fu5ACK+Z2jEdlgeBohDj3r6BZtXhr7cuLE70t6HKgO06NboASi5CZruicGLg
A8WXjaF59cTV1wBrpUnw6XGE+vtYtPoeJ95VSXxjJX5FRkA7WvAMrbeDna0diT/R
UT4IpWyCdRw1HZEn9Dh2DMoYHJZfQZE1xSbeK8lkTUax0aWBsu/VjEfrKveKmDh9
NANm1tY8U3iK619q7FUBVX0lW0j5wECS+CQOoMtPAIvHWPL92GTr163dTwlRl6p/
jF9K/STfSgdBQguvDBEwp7nWN4+moQuAZJRzcThTYzaAca0KYHmmuPQ7JR3Txz4j
QWi/QLzkr12AEhFKa4uqRdnKWrhge7zZAAf0VGvhUQ/bf7jiKEnrX1W8N9EgK9+y
fY4x547jb6peWtRG+Lvzyc23Qpo5g2BtNjJKMVWg8c+6ciWZFhd8D1LjEY+iEq3c
ecCDX2Pp863L6T+fNj/7b6xm+Qjn4YA+vxnXsQMLn9ktV19QRcF27X5wDwsmCXsl
wylPGJIceDX84mxrgyllhI97hNiH+cb2LFnEjI2VlQ6K34FizBfwHI/wfkPvh2wm
YMo0Kt+wWj9lHIMVmqCANQEEw/6PYKN+q5rLOf+pLh/Cm3BTMojC0/x/CeO0g4up
OzKXTh0n+zOFjkSmbTB9baxGOsjRgV1qcIswfqqUoVZ9jHMzyfE19c4Pk8SpNil/
6Zyi9xqvbE/7otc2fpVXMoRVhbmBBP8zrOsph3f8XmwaH2WTqs8J3CoQDNjsdPz/
9kDGWxXjsnViC+4sIhiCryPI+jU6IjodDlTIlIVoYg2Va/Q5d8l7Oe6GhVQcJb7e
Gb6yaNEIEShry1STEo3BIGeDRuHymWP29j4GPAZNEH4AN0/3uCmZKU0CGbsVQcfU
zOQtPWVl8dQiCB5eeS5DwIQBHHsjryTfhqFpC06qmV5ELLYB+WhPMRfGKTnKmymu
udxoQgKJ/jM7OZFT7ULPl8yj0SwupokVUdUpAXqpE90x0VI0rRtPivJtDjBb/YLd
5taFebDljDv5fb3NbSd5HupdmH8IZg6ITFyrUlEN9klkan6TPpNmzmuJQa48kNmW
eQzP9mreQZK0bMCh15tbLr08ARATkUTtUTNB/+anwIbzSw7gOTd1WTfa0bNhAxA8
bb++68uwURIWVXD6L8WSYqvTPrM4/YuZMYUXQOGlizaKd7GTP1LVztBbVmQWV/y4
NcRC51BkaV4MJ6Gbz24dCW2r4Ed2pSwWQo7AhYN9nQ0NV4m4GwoXHRUSN5IA4DJx
xmulrTyJlo3ZYquVyzgZ/x6JQfuJfwmUvxONDmjvqY4+2AP92FVFZpXEtGtwDz5W
6jFbVdgNfS292Dd67FtKWIotUJD9y3q8++1UF7TRGOsEhoKAi6qvBEzg5xkmzlsP
Qir/U7urrroGrheFH9pkbu1rOOTPLru24SYPZpS0rAfmebNd8d0lTM8fnjDirKvx
d6ExYdFRttdhrSPLpTXYxbNhBSfEI1t1XE9PmowrOWR4Huf+FOaQeEt85Tn0UCk2
HwxFb1Y/imZuOxD6sFk8EQkp07NqAeLDrlMfTbxT/m8VuBE3JITdfvojUbvRYwAX
2cnAWCm+ATsyfVd0k6LShg7P3r/NleO4oWaeiiVYoibR2n4sAmUnPhJPVhyYL/9P
Qawssx9QxFhtsjUickmnODK9499dVdnEvIou6NKi5gVHiWCLN7d5tlMwrSRUR9QG
vElg4XKQqJaocpUZ7u9giqCQ2b+IYbuqa77NHAaGTmeB46Dirm35O44x035umttZ
m4Kb67jcaZbnpDnSIhlpFqBUq9ah90NnSY0IMtIsc+2dSi7oALpmdN9utmVIEJYO
hQO8Ennk6HGogXTcim9oydCOhhussIAX8+XRJ6kvtck7fv7xairtZYG02zJZfIkc
Uoacz7DoURub3apt6pWrBYaUehEP4IpU8baOXuXxaee3XK0EHKi6GnjC3llI4MeE
PyvOrZeE5Jx0/tytxhIraG5iZFAelYvKZHxLC1X0RfuFyrzmUXutZ7KgXTh5LdAq
0WsVYbEWem9T9uOVh86UGc6FeNTnCvPiqXTrIDRsN3ms03muC516oCtwjdsz73tA
mNNoPCEQNOp/8xofuHuosOs/L9FoQtprHjp0HFrT7hEPSG4MF/fHVeD5FFS+6oNK
XZfZVVyZYPltAaTnS90k2yeUpcl/FZI86Aui7i8Zieq/XlouD5GLEfubwNCn3YYa
fO/L9L9AePOtMfZvinD5oQVHnUFZYzwGUUHWtahtCNbyWTFSc6Lx+4wysva33EeD
yFFPeYoVstEsoJycjt3eTw5mnXQgteoizsackSpSpoC2ebibiAuQ9IAtzrz10miq
x+DRBDmg40XpeFYcisTmTBe1yG+HMuyxNw6MqRwpid9h6mtBnwVuYUBnurxRn0jx
3i40j0rh8OjtD7+tGBkl7usFF1NixennLtsV/VFuJQSHE4N66cFKzFCtLrYg0GET
VHwqOOiBrGNlz/99gKb3n4Cs0M9fGVlCIAtGDEucWUjVKvAJEy2PixtUcaZFEQ5J
6iLP+fgh7Bild2h2U6wS7NhnAmzANmb+OD1J1KdPUxbc0Vk9aAq9rBFipfFK96rr
VS5LC/ofY+ZY42tL/KQhvUhaRQqgbdSK6Gpj37ZLy7NRWcTFh/g6du/Ski+5Mh2w
G9TRwk7CxL2urX9SndAJMPQVOw+x2Ex75jwy4ZzJnFqfY5nsGqfrlfy+QfRtink7
cBAj11ZE0CmEzQMcPbL+JfBaVG06vIP+1s9f20AwwYY0nnxpUy6OdgPzjlTCgtMT
juq6UzhxeGlTNNpWr01udXgI7oXc70QDcqmGWgDCBIGk6AB4C+TxKngx7/Vu77L2
jup/xeQ9diNBcAZ9Iu6WFEPTsp1WF0qHRwIKOcoJw6PYna2626itjEIcOBF9vxnt
uYYek2w2yw432LCbCUv3d/Ih6hZbtVogI67l0tQsK/6MMvJuuFPmt2SLL+aQF43T
7yNVYkXKA1/HYpxGcz8XHkCRB84q7c4sAqGgOfZLoK4UtXK0V1cUmR9ZlOwLdX0i
e+rVJbjPZYfThvRKTqyIzj2yzGyMyamdjxtQ9Gqedz9/1QWfatevfrjyTQ14Gmsb
Z1vRcqXuaOW1nN1Wsphm8qIZs4jUA9m6fB81nx7tLipdzSf2NOqtFnr/DujGyiY/
Z/+qjRriDfcIiUrXAia0HD28QBv3VfJUO8tNacAplHbiY7zt2WQzuKV93GSnuhXM
xD6GMY7ZAqz5JmYkNONAYFfMXFwnnCCesNATTm+IJMUWcIbhuZvQzoNaDH9JSx1W
6mYY9R/y1lphVTXb+c2ORPgy8WEGBfpCH9bLqSbfP0un2Wjge9zZ+FJzNbA/9HkN
UDXaCsIiclt/aA6TOqwsKseNKdqB/RAWi/L85mwTAMxIBZ/xt4AQcoueHXzLu/CD
6b7J0+E/rDGB0CCZ7mWVxz1LdLU+mW5MguDtEOOb+Flfz/hNenxJrlzuSU+qY5/I
P+4jJuYLuqaK/1SYo7XW1kroBG4wWC8oIjHZkasawgAwnh92Ys4zAvOHw7OESxTV
P3LycRHdDmMr1RGTaVl6BYOYboc84/YJm0qHPVhl1rb46qZ7UE9ZSAYCqXiibi9z
73uMWdt9VeeAZsXOxaHqL+Spfl7p2YoL4KnXMXiqBqnpw37GFE3UHXeqniPJw/xd
KUoRPcLQGYdC7yCkqDwWmdQg9bFmmyItkrbUO3stRPSIwkV2K8kF5kjREEs+GJAu
YUqV2+5H112poSg+IAPFDC07d6EA974Rm3EV4alo3Y82enorfnjTYeRAtcaoxY90
aFlbJ767Ni8qCgi/uWwRnzshHBf/bytWz48pYa79Bx1XiuyQpC5na+9NnlMJx/IP
PUpIO1YwGTF5nfBNmbP2iGBZoIYoK6Jlnyh28SIJvbp4NkyzKfNeko8T5kU0gsLx
7vce569wL/kqaf5ny+BU4wkX3z6tt+InC2eHwaiN4DwmIRV28ufsNJDa17MYeVdA
N7Z+w/YtRYWEvshzvmZpdYC7kpNYk5vldyLlr7FnCkav4mfTWb2uHvtPQjjyySFG
eQLgf13OoV1LYD6ckuqC9X/sUFT0jL+kp4IBoW8F+6EF8t2d4UqmZ5ffYrSQUUpF
Q+WHlgIfnkljXtg79qvz604wE5OQDrHisoiX2M91Y18JBGoX6bnklvfaceytnJsd
HfNi3HAD8GbdRMqIUXcbJW+qDr1IK1DwnaTYivkmVNb41GiUGey+Om3xkiUOOmKF
uYBfXIYM2C6/r1wV4Vhlyyw+s/6hVkXpeOWnd3P1Ltb+aiy0/mY5aTBW/MHhD6P9
6wkTUiGrPJD2dCi9f5iHIhb4jBeOs2VkJ7YJkyvBir0H3xBsmf6W8DYa7fnVGNG/
9IGoKp+A+3Ku7sHRMiWBO4SuJsNk09AwJVOXwvU0wetsRXT3b4Lvbtrn5CgDL5G2
ZaCWtPBS5mH5l2j5gvDSlg/HIYG9Vbfs6/7QGAXEEc+foj1274bVC2UMmGmA/8pN
Ov5UkLHKwyqYWMr2VTU+IdGY2IfTx2YH+NfbL1Cq8CjIGCESeLotWETfyUleTkIp
HRxD8eS4bRqwDeA4ht829ioI0+y1VXfSqseXfLMvv0wjPRSjrMz4j/09GmupI9T7
T7Kk3EFNDkhJx2pkift6BQeiwS/DCBR4ksPgjn7crwvOUimHMH5P8gzmdy2tKZsD
7p7MCMt1pXRW1pU3dtymD0Qexr/mz3YkAifN6ey1SbEsmein26oneic7sRgbYgMj
xL9x9JSquq0dAleAlS0ADQy6mqSHkZKYYQ3C9EB47UPHtuXF+CXuFQs+4bKcJYkT
3FzMDbZzN4FTm3YO8OfzNsElWarbEElT1wBnPLNAt6/7nq3JNGClk4+CYkClyrHx
VHMiW0c1fWOHDXgaoUUQgfeh2kO6VqCQ8FAeoGEaELNtNTmApUmdLQkC2E+SM3F6
Rga3f0WncRPl1sdSlqjzjq5ol+LhX1haM9pwl2Lv/XBn0VXo7lTRlFlBd+9fROXg
8FaHbj6UiSsyDZVxXt7cCAk5wekofM7A6srlU5z96OCx0O81bxp9xMcdSMZBBkKb
M8Y+dEIr87NvzKMrqQFJzvwY/yULWKDaShop/pliDpcFnp08KlKTSS0qKFP2CY2n
NnXEkAg/oIPQi9FlRYwJOHQUF1w5R3DMDO+vYor6u/Pa2Ysn1TMR70h9sgRGLny/
BCDcaG3tOyRecJvibzh/5Wn5dMl4JKukhkqddqbdd7+4DgiZGU5jKd7RmN8Fl9SN
D6xjupBc3ACjgMnGfCGQLHBioAueV+sAyPYG2ssiLhshbKfFV1RU8AeasfTS5yC4
hGIr3YcVtqdn+HdIxagG9qUN1e8/pt2FTPKDv5hdtjk/9DB2dV+UyzPzxG4YQlS8
pd+C6FVrqnchNwzzYB4anFm8BlqjykUr1HCvNini11wQ2Cl3lPEywV6Mc55LJ4Va
+bydchuP9FP9zReE5ZOs608tM6PAWcx7p8g/MXqmZgA8y6oioLtS15Wy1wjROZEL
Zg+aQmtu39UfMUZGZOnQRTdLNMWZWc7iKOyqfGaxFPnaHl1ABWiZb3y0CgTmL57B
FxF0Ouwo79wrYAE3kTduKXfYeN3fY/D2ZxyxUWxiwpUt1FJr8dFB0ihGQeR++uqZ
65W3t60R9WSLTkqG+VP0qCcb+sI0MhlOmSS58mSQOAG43krkN/FYkd4y76lLmu1r
hRkGMfphxu8XSJD9nKBCnz5RXNG7XXa28tEBavU3+f4eXaJcy86jOf+9acG/hhDe
UHatyJrsEuGS2Yu/ggbWKN51664gEyxndEJ4F/jwmpxkO+pxejM2BsaJdbE+hGuF
USWoIQfoSpff8R9HKsckdKwbD9SnhyzK/kiJP6VRBTvDzgCU3f+2t0zaehjn8QVK
9waIb+LRW1WKBTzDupck8NgBVX95810rpIh6TWT4eDZUtrm5n8/n1kPZA1uJ+i6p
jq9ePdHPuDQIhIdgSIZ5pna7iHUG9lPSiVa1A2EWYAd28JSc8GovFGhOazZ31Hrc
DvZcfFnXL2O+jLCAPrwhNhYcB9JyRyyQ+Yyp/P51/Zjo7jU2m/IP4zmNcQBa86v9
8d2yJzYfWWvNXapfELg/zBJhQv38dsfIEdHCxGcE2MZzGGNlZp/sfxc/ObjYwh/f
0JeS+18uD6N5buJmaycezzueAMJkqL1t4bING8lkHRV5ltlqju09MjtCir9YML5k
gGkr6aOX/gldZo+wpLRvbuYymd9J0f/koxZEueSs9M5OZb3lSdMvcmn2dZISqdds
jc+v4iYtu6kfO9KOQnLTkM7jsgmdrdc045vqjSJya7HNTLZQYEsyjx97uS5U3mKR
JGg7vzy/OIy37G+GisSurCDv+n0D2Y9VOqo39Qqzfxfp8gMk7/lawAr3bn/WaIcZ
QmdH/pd2FlA+bo2Eub02AhdEJXrtpGRiRw1za21UyIuxopg4s4uUR/Tp1yg77jdy
tJaYc5ana/w6e53cARbX+EKb8a2YBXrkE2nr5S9lUWqLkDx1d+qMN/mnU9ea/Z+o
dXwlNDk3fOYelk5rlaKSu6GvEPn+NO3v69Z+O5v9cK/R14v5VF/usqulDkwq92Mv
m0Y4w5T2TvD/dpaLg6BtTodNmfMz8z/iMTc68PZ8JUMQVE8FLSQD3+ch9RYB7IxY
p9bSNo4cBR96NPP5EAO4bhJINcr2leACP4y6Pp8yxviBVh7ANn9PoIHegC0OOnRH
mk8HcKZ0bbbYO9lG+67aDszMAdRTGVjLDgH5rfcwedrzfritGMdxsxF1YjG/YEgU
s3IewI0YTDwQZYQEBs/LYxgWWIqSUd1Kg8iBWfkB95fu+XglbcsrrQy5Iv9pRP73
QtkOjr0CfX1MyB/W442Mdho1p048tvGMBoZai6xvFRINRqSt5oOQ8IXxg91A/vxj
Jrbmt/WLFRakIhPHYfsW9p9qNHs/tv9Pv5xdVX4nubvNM8HZeIJ2h++k/j2LTrFt
aUFNrADF7gr7ABNgKqdsJ+f6z1H6D410MZ0g7NdjXOfoGX6D1GB03qAKukkyqIG8
T4ALFV9btONT2c/ymMXFQUMLHopEOTTHsFspryvkufnGpaNqmzyB2Yk3Vghvhwn6
ppdbTD8/oP/3JEoLj0TzLHBIonF5atNBMxazsDau+bT3pDcX515Z/zph9C2V4ChR
breFQcCPMNwDqeX2U/MI6Aq4wb4X65YrS4mydzwEg2S66t53q984eesbd6q6Dhe2
sirLSRPSDsSHttpD5+KL3J0Yiehm6gVQ9mzOWJICWofXyDbXXV8KVuWrr+x8DFks
l2GCi3WhN5AGkiHl9/JF6Fc9OGgEZ5EJJxu7rSEgYi8EyT6MMwazEPg9hCweN+sB
5Xu/Dj5+ypYxgExRKjBVisnk1IAT8NyLH1y3T0dqa4011lI9z6eh5L83Qqtpc3S1
zdP4nkjDdvWxsqJNdQ89fCUlNq2ZlMzQw+faf+s4JbUGI4sRY7SBKAyp/6No1Qfc
CB7VKkr499KfuSbrNd2pd5HM2hO4Ca2ZwOmF612Au8fj3B0ge1gFFkHF/8u2ukW9
otGF82M0PqYXZnSWoFeXPdVCcCFasLlVM4Z/WlGC/UkWQ0QJz7Ihw6y9yDc8f41p
zoqKgCPs2sc2YWAqPGkmr9U7iLjPbjvUd59wfMV5fQ5ve3CUCNXcLcuGOdiBEkvw
gjNr1KIR44Qouq9GRm75gA9I01aAeS81shoAZAqt38EtGFrnrnixMCPVrPpZu4Fz
Fivp89o+XNPZ+KpitZduuVSG4YUr/oJP+k1x9hpzpufun59/aflCiwQIc28Lwrzr
lOFiIAVfN4SwhQQe2KbzB4EnWmnfnDKnZEiVRL4X3vgg/ZCEV0NT8m/HGQLj6qhP
GZFPg5Js8KjncuD8nuNMnZWfvGGqVKKQ5js6i2ADk0dNi+ZJfApRJqGfkbmPiyor
+ntIJDlalX2GC4yhP2jCYSA9i3mhh5pYKHYDB816vlliTFaXIp0+1K8F5p228cQ5
M17Wd52piQBxJr/ArgcSeH6cfK1G/7nOIqeaF55MWs7CQlcKB2x2VTvnRkBURcsT
e0Y7wcF+yxFLGMoUWC67SEJ2xjTytbJ5GpwRcLUNjagt3fCztDHr661FB8Ab1s++
3xn0S00wa98eGRJJKDOjY/FYLqsoOEcBklqN3a7meWonSsYze65yK/3XflD3BXBA
9Km8GYxEcS9MKsko8PTzUGgYKMDQgUR6xy4m2xerYK8wnXWZ6106JjQpsroJdQGv
veJfpsPk5AIcHIm6Bd0lp//sx6cH3zf8QDEVVaAW2kRg97nTitgHWR/Qot6K2Sdu
LXOUZoF8QoSpJ8rMJ5tMZp65ANExZO4MAXLcQXUt/8WEMPCBcxNxIkpoh4AU6s/n
/0Zn2smGOvhTFMwV7jrJ73PeNjYGvuZwoNjOetbxoZV25qeFBRu4wXZFZWCw6/xb
smeL7Qgj4h+8E6YN38gBVbSmUCjjnyPh/2ynsMh/FyGQRsovpuiiNZUspUd86aHU
Q2BlGMNDP41WMBOZB8NwLHjtx4nJ5D0edpGumR47UM4OmVfaR7nZ1glJeSTXFjiV
1Wd17KkCN+WjjnbtmuVzyWpIka3XAYVYEAY2xAIg5Lw06ygGvVzHgC5FRE+rR+ld
uW6cJIj+J3Lezmrl87N11679afRSzRiyR/fn2B+J6HS6Y9UvuvMcbo4/zUSsHaKv
ZK8FNKXyjGPAZlSaqqnfHsM0sZ0iTT86r7J8rOsNBNzIHPato+d5Svu9u4cqLAYq
tbq4gxDIo0B4AlWZbg+d1FlsNVNA6nHnGPZqbPIjmzCw79DviUKvgkdDu0jzJU3f
hTnDq3HK61159+PTvBIOozkv19cAnKNqO4g/HYac/ejbZZi0XraNWYk7kb/mORnK
8lGGH+KlU6JeDvVMXPAoGuH5xeZCqPuGJ4yv+NFzotgApN5LpcgrqpGjcSJd9M8A
C3JLJ5y+ByoHb6ESmJzZlNheqoURNiXR7A6og30FjdLgQUrrYvtWMNCT2ztR7iTp
SDvzz9H1Zi7TgQf6KdgrpkxsABgIU4Hzhlvh4Dkov9p9Ohxg32CVGVWJIb6tyM68
cWZkMgckfj53lzaDYmwKfQ57pWguQKO3c0V9Y5y76qjZWWFto2oZq02MD3w0LuvV
PhQPY401o43OtMms53RNigbnnRoaDGa1dzoMkdcLMd9Cc9ggYRubtRyKokat/NSZ
pPHLlKhmjKDKodu0H8Ww9gjS5a+aUSNrVAD7Kp1o3B9wB23HGBcvHmhAkeIUhODx
4NatDsvtAxXfTM5tO6feBnRQZlICasgwZXKShUmB9ZqFxxYF3jb+W/jVRArAAg/V
2Nq/iS2/gzvFWz2/fBOe46h1nYOXRSRzxe7Y3C0J/7M79M1taVmzaJsNtjHl0L/D
6wBy/a37JwYs9S69U7JLxYyW7lwNCU1y3cFZ+3j3chlg4pBf+qQZ4U2bhk2gZVjK
Wq3CQY73pUccBUJEuxJAyvxR9RUKJZH21As/V7NM4esbz2ZeevOuOoDL16xv2qP/
UrzDLU4372m6SZZLnQARe5pE8tqcdTSiJtOH2976CFbHVd53ordBeje8hZd/cMcV
buSoYaFIzVS0C/i2wPzHM2+UC+GLpGSKRsxSWmgI1w73Qx0Ad4sPMfFkt8Et17lk
UPdB5gxU/15Q8ETsOQZaX0RbBSoPi6e72SPaRsYxse8dlTNs2lC8QLZ4PaeL8DFX
n1HWZCnu2YSy6q+2l8/37vkFL1y0LvofWdEwgb03hzcbjlaroBXmOdQfADSdWZ1p
+q2mgRnvnoNwJQKy8qnfY7g6bTnKU9KWf5iypSJPJvWpCCtnbXt7vOcYY0lx1let
6LponC87iVCcHLpFbSMf+CJKa8W7BCQqh2axr3RNXrKmKuO4oJNPb/GthOjIk6Em
pcSvzzy06KkwkoiqZUTumD4bBED/dkudFNRf5Z3Yn1bof4QWLMrmdzpQXsbg6s+v
rLIgBkkfhafJQID56T1rDevWy8LNtis+wSl9tTMUQYAOZg3Y2o/hmCwrf70yHLzB
h3siPsfjI6WKK6YJjLLvXTzBmyRzcD4MjP6dbW2CF4T/SX00FymEA1yHiRFwIxYb
MSpUPESd9MuVc5mqHaPIG+wBjpCr+uqkSLC7nnTig464xwreWoyv0e49FP94o5+F
R3+gCcIuYnfonXRCO3lN3a2A1Tn9gIA79lICme8uCGbmLpIl/PG0wXK/Yq5A4e9t
RkaBsTVLWsGbkBeDk6+0EPPpWVtdUBncXEr4R/CHU12WDMq4WDi/mHhEh2hQi0Om
8aLJNQUSRjRj0tD7tcTUSBHBF4111yc9lXnqx/HucWDYUnEXQVw9HmxhdWUYD2Z/
nlsHVlOqpyy3QyO3Cy+12GYYq+Lm9eVBAkRjUvVWQxc0tQwy0mHjj4yr9MZf0NwV
CPgHIGrJUg0ORstqSgCBfD5EugaIfInRC6T2Pyz7lIjxFCcdtf1zWhKyvFoIF4V8
Rm7HX6IAP5rfGK8vie66WDwx3cM1JhCfER7prGgbD/TVi3aJPdHIYrMMqG4BMkag
DEXZpHK1XxbJNHco8iH7IzU16+FRqhMK6k25SR3oMVjbhghmoiJUC4EQrnub6UKt
wsmOvmuQad44YPjt5NbiITOUwrMkKCDBZPAFLbD1BcAU9pWJXdbjdzPFx/aJnKBc
8O5czaNT61JS5ooCIvjgcrtpinNAHvdCIFCiwYAHAeDvh3IstmcJXnCYBYFWYOUh
Zuzu2UfvivTTsKO0endBzH45KSIl4j+9SP6leA1qac0wsl9X8bMjLL/2EdqnufVn
/pWuZWRpZoIlgL/jHYU4cTEj4B6yWtIL+Jxa/p14qlvhK8XZHOvuewvi5p5ppwY+
bdnY9sO97/Wvbe8HLrYGSe3nJUEI+KCs6UTMxjIvCCsjzbNXOuEr0viU+QpYBszY
FNl0LIrI3+O9if/9Voi/M+2aDK3QYKNqRNuUYDwIzPzzoo3jKh9oZvlcEOF0GvWB
Ja82A4CXMwE/+laNuZtBcZIfpbAaI+yh6OnkpJ0A5u96tzmtrWeePSZKvOUGUnDR
Jw5XbaKFjmnIMBgSCNewdcsKNlDTjFLuI8y1nOm0g803iFmtAGmi1g8j13+JwxGO
FGt4mGLI7tvzLhiHUMXe7kTa9NcbUa6H57o+Va1xFR9mQujOXXlnN6XwbyndoKHL
AvSmx1ehZnvY/9NOHFp9di6RlLP10loFCX2pUYB2pA+Vmj9LevLgzW4ZJxZQRERZ
+Q0I5u9YGuNWtYnzGG32j9QpA2CDPjdehgGY6mU/s5lU1VrmB8NH/NXV0IVK8jjw
h5bGYj3dNcOxt/BiLGFf7ioaLH8wOcHQ4W32Fc7WOgPpBTUVpBazs+DlMaOo8uSS
0Wk0JasMGy/nBl1gV3aAfd4iImsG4EMwBlNq1IdWwe1OzrxqajedNDtLJrNxSWtW
YdwZFLBatfXtmY/5Z1H562MAv7LR2vn123KExZgV3/ukWpge9jSEtFNndlLs7Zla
2IE9X2ETIZvuduQn74R9wMkvvJ5kQ06XgVXYIiN2yFTMYWb72Bmj6wqEXEk/0fbl
Nvu4dnAsSbi64N22KQ4pYRvurQUe/gM/lB4JYEURCNnI3aXsizuVoE03l9GUBbVg
BD7fSJy0OhQeINV1cTNwPIi5wU1OXkZFXNbxG9ZiJx363wzKjytupbKcefC2QOBr
j65g4zPevvvIfz+IIcnYPapeTYP3KctYJ3qinJl1IcVxh+BJSCoqvWlWKQOYaLPG
lzVp64bzY3XGkOXUHIme26cKyu+//+O1ORio+fZvqYEJXtqaJKZXnP6w96iDd6rn
lKnFPdU1pB+wKUzJ2uz4ot80zscfqyTrPOE0JnFcPi6OcfYmrLWRMOvIuLl6WQxE
v6QkD/kytm0+oecaGOsQSnHOaeZD0IhwRROSjw4B27CqTdVZmzPftzAO1CLn5yuY
kuPmecTBx+VYWztrYXsMsI7ZqtkvUYtYV8f88cf35Ym4Ang6O4TVG6ZumXo9hXxY
ZlpNLpvsDrqT9BMwM4ZVFbrz5XJedSp7S/KStJaLUMYdZ6a/Tp1kS62WEJLgK9Kp
0pG6rDO/arX/LJTc+nmey3GUh40fQxbBt2SF3kmAqMQA8eTTu+Bn9MDCdOIa5rRI
gzYkur+m5WyY4flI64YXN4APxOTRzSiEp4v2vRn3JwsxzpFayK0fL5weX6a/VoIw
O/r+1r+q5oye5R2lOhWwG8r54dsxM/nbb69MiTEBhn2LVd0v7YsSF9lMvGi/Xf+4
srjFd7GlRDNa2Qqca7lodWVov2VLvvlZ8JLygC5CHNCVLYZtYyQhDgReMsMQeNX2
Sb0vj1Xd6/2078sPmTZgcGXC1bcjDpXg92+9qs7667rLxh1d8U8nvOMisO0edOeD
DV6HwM0Zp+rdEHoxd+mnfjMcdLQiIE4NOToaCOnR5O7/22Rcid6wt+vX9pabTrVx
EsWlZOgO347OqclR+7D7ECKBlbW+V+OIQPh21Nly5K6uhWGErHhweIL9McJbuhqL
OyztWnNYtmNGicymlyCB1cZ0e8mjdlHACT6JGgh7C1c5sX7ikqRQ5A5dg047plTA
XViHspxIRD0nW1NDEx/mN6TqnMNvxvPKeERrlb2EAnCkDdVVuNxhd1XzkmuFpd40
3y2moU7W/E4n7t4vN6bJNvAEkqGnyQtTSvEGp/YWhk4CfM/ZuxTNwlwOWqGu60kG
Xd8Sa9zmpdI0whzXf+9nvAvuDglJCfd17iaHnPSwgZr0RHpqWBPz4jIetStdbMKW
gGuroVF6A+ZPU41Zibnaw8qDRBSYqufUGWfJNe3ruSFDHjIXEgEkiHtKMYHpWpbh
C/EKaMshuo0xBBYerzTyZRZGh0b2QCcw1MFJi3wBdz24g65nffBEVRty7utGtqrc
OLDT1z6Xm9+VRkOidTeCi/d8ZZCT70xwzkM0zWZi5ZAtm4c+FVw9c109M1S2jDgr
VoJElyUOvXuY5UbOZLDkBWfF8/Bf+hFm9eBaGVA5Rc7mvDy73UWxcEY2T8cM2l/W
oiKk8T1O/ACkZTp24UIHD7r0iZFLAGT1mcGAeRKBb8gTxwPhorEc0PnSp9Q7sBfN
P30i/hWA+yAA3A+03G0/vR4uvf778Ki00kBhOM1ph5qYVGNl2JitAPfoP21kvekg
nNNmhKd4LIrAC1b7lTiRM1wwAR2CDCk3+aHbfImfrJjzPz6jmnDoXqGHKkOU3yzV
uy2TxgCNkC90mA1mbsr74wMbQ3ftevi+SsP6vN3CLoXdiYdwp5eMGaqSm58N/qKa
TZw+G/8ZckKVqeEmmEZdQt8UmSDxBXKMj2Q/pJRTKEBqfeUefkL5mn9rKcG0Zn7E
SdgyS8q4u+53ep67qdukTSUmYqkxhO+Q4eTJVAZVJwFpe8u8CYFewPCHb+wVAM4X
1KP02Sv0OlU6lmgD5geTzN/HyzC1NkZTEAyCssbXEAeV4k6M3vZpHfSxQ+zPy+AV
HDKKSxHmYEl6w2qwhlQ5keVrKoekfBIG6mEMNzKl/7hrK9U3BxBkRkzSUvKndbum
g+K1cvQq4F69PH66+CFSPU6ngzYEpSVk1nNrCxdtQIcRXhh53LelFpSxR0btkU1L
hdoS47u6d7Rqk40LoJqfF1z8RTvJsX7x+SzcyjOCOiX5yhx21LBssqWC+tuf7oZH
mapFgPQOj4neL8YfBI7OV8UyxUU1yHV1Nu2nfK+/T0TcsUZZ27CBmgf2TfZRlIgo
krG8yuy434iwIc2/NWqSDkCruA6Ye1WY9XzZrFOHkeyg6WPX5bJcrAXvt0H2+iGO
mkgbYviRQQeqtKd8jFgZZMOWovBFGurJvNSrLPFdKnu4Vktc1D1NWMJ2LLFZ4D3B
T/122iU5ZiR4vrzz00UTnx6L8Pnd/AxNNkeBUgsBvLQSFlbnT2BVlIPh9ky6Ysk6
K22OnKAc+sVbHBHYa/w9V7zIJxzonopP8Z5REIcx3O93i6HET4Ltao9v5hNrPWKc
Q+5mmUrv8TT60Xoa1V1ZmRTySoHkodauyJZmFSiBBrKOlV3+gCahQVGdjDZU93ID
G3J+pqlhm6iyLWW44/YvMNnOSXEXwr2faRFEky1ishtadl6BKhI9/hcB0OJw06We
vIQlFtpaZFXcl+rJMEWsluUnbgnosYJZG/nHWh2aqFShjMxEiKKDjabhdy6DCBDN
dcqkSGjW2NXn3i8srVp6jRfDEpQNIyYFmmvw87KUmQI5b3Kup3o+Qr5EYcE+Pn4d
ZiNBjunkBijFYdVV+hLGz2wpwOARt5N2QaPvuaRRBqkAeX3umKi/XU4MCj684QA3
x3/3nw7e06wrAqd0yVI7tB2TQetfNr9DhJkRaPkzS9DYaNOgzcstmMwOleAwiKu7
r5Q9Z/vF8mnfpbq7ezyL1TvibfAM6/Nxr8DCBi/4t+8mIcMFKGBczQQZTvYcKK2x
7SUbOV2s1CCW0+d6T5LtolqfKhRSutNeH1PHazFClTYGBA2ihsaT1Z5oQXfBOisD
A+EhywSFKNJLwiMz0oGFf1Pt5GJEw2W4pzFeGObc4R48/14nwLEMf2I7v45w0uHP
au5bgv3msVugSBjXapX/4WRV483PBEDhh7UrMxI6eCML6L/RRuZCUiHPB0RvdcxG
B8rFVd+2YMz31uVy7HEGfSB9udoE662Xe6dCpaB/NWJa8I0F4ihMGX17jALQwAci
8fB18TO7itQ97ove75dDO6IdcMCUDqyPq6LrEmrsudSSfXxPoknxiG6BRIYMaj5T
A4Vqwtl0Ze5CPbdyGRf8RrlZUHx/w/yisqkFLehiH1C8e2myh884eTJ9Op3Dg87i
Zdae1W8NKCrKW2Zm/KPUh50HBr3BUU71r3Wjl3E8UejiQ9bUZLfluZxS64s154D3
K9hh7FO8Nux9m8vcsuH1k7/Nf6ii/WZzdr6IuDywHM5pOQxCeUN0kbLmFVnMsYeZ
LAKPoggCfO1t5y2xcRiPTjb4pmK0U5jdK9iNEvVbI7wQn3qNZeZ4YOopNYVrDEv2
yBBGx41kYWS0PB5RN0rApksLCGGXT0VkiPPWC6ZgdiZKsiO+kOqY1C4j9Lct8ntC
BzF2us3jgbkXrmAuMy0S38FQRDi3cPOS/9maSQJrQMUf5Y3kWMwg5p1anVAdxmML
kFe4xZn/VMadRG320UD2sT//UbRIh7tQOAJduo2ensTBwkZlKFgxKYlTYfqgqQ6F
aEzpkIi2IB4SSfdiFqIibxQMAJ6smTKFqim5BLCDDtuISrX1pcH0AhU+iv3SZGwr
6tbwS1EfDRUaTqmeNzS5XI23p/dIE5TZqJHLJ6UaaCMcoXm3xf15Epm1bF+8PL61
VitnP8oPv2qv71O1APeeNT5lJ04HjHrQSREw8xKTLrztCLnNy5m1RNLcL+VG4nWN
6LebjowFNJSYXAx8F9KpsIDGbTfUI/TOpPpzyV5sON0olF4gV5W78VNIZgRthvC1
345FBNfstxAaHIKfw9DWpvmGn6Ea1yaszvBZRh1317FOOSMHEodVLgDcYZVDs7e7
hL3HOGkui+0leSL5098068o8HtZ42xU6psIRzBzuIOIDMQz2O8SPEgu6kvk8Fvb1
tW4PeMyCjMDtNuxL+tz2DnRq8rGCl0pkEOACuj/lfaD9YdbpRnn023cF8WXqaB+f
wuhHp7cWvw2Indz7QnQWdMvQYBAdnMR1mkQDSRv+V2M/zSKuGz7Fu2VzmARnP1Ye
NQSufMkeuC06q3NQ1aiPgfU4AUH5+taXRntmA/okJzOP48m2a27qlb2dDZpHbsN+
7j8TxdBkf4Xzpk+QwMYAMr6DPTRJemIgHvtjytD5j0QVP5DgrhqBDCw925Utptpb
OHKA+FAINQ0EuMnfdDXig6QBjTgWlDW7ugsR71Ym8DL1/LhdBs8YNyREdzWROusy
YAy+r7KZrnj9sLBl8b/D6dyM3ewmCSmfRQ6eZwJqaCpsQzodl//F4PwRlHnXxAm0
ciwDklITGFaR959xgkL9cuUD7skom8AC2NNeiMQjZQXwdgLHYNadNjX5zLyeMpeh
GRTLgampBYQ1e5i3w17pfihqYM7/pVvKUXyEc4GPENVy11bt3WKAvxRwsAWJlkSk
NNleHsopbs3lhR3nj2B6R/RohD3XnNQPN0EbO9ux7gtYXg/7CsG75FnwJnO++csU
FaYQaYcGa78yEp8rpj+DnYAHsINCXM/3j/OEbnpRoYl5eQNau7QzjkbTetsnVRrf
nTPAEukixAPLsRDIWyRAR+UW6OSm4Sm2JRd7WxxCh/RCVvm4d97cL+qgcwlSAYh+
UTqcFX+kQJNs/gWHYD48q4eR5nRI3QMz+wwPC6Cp2HcvsohYFBFQVOhAOzCs8Bmt
HY50y75Q+BG89I7mdEd4l0m2uBH39mdd1rUxO6TCYrPXInHg8QMIJp0f5jB2Cj7G
Www+Ck4P7YJvpSTckUyit1zAypNKbH3urXlXVDWgMqxt70hRiHXlRfxDXybSAjRd
U9J3TWjTKgk0Z/G7fqbPJuVTvgGb5g/ThLCloD58132tRPmjFoqtN1X5UPpMCrOB
pkIr8Sqfy9+4lFyy6wKb8R2pCeKjjIuJwuN3upS8A4I4gRtmI9yL9eFiK1h2FZkC
VWLzKmMqqXZ5UFac5yDEsVS0s3nWIE7zO7IfNx8jRwipKHaoPvx7tGIVRhBXGpqB
gNADw4hT0rjjlCQz6ZlMttw3Mw7PanoJJ/6mYfdc+AfLODOlYEqQJKf9LBfTPQKS
zDMSmrJdzN1SVIfBraGHOHRQRxapi8LZy2bF0rBH5b3/sTghHLVpZW/NRFyGkkvV
EsS2w9Qumcsy6g5iOkfBpyBdKpHLMMamY3U6SXZy8BStT8ac8OcMYoZnXHZWETit
OOcsWISbdzPVBiUwDyNtcQAhMwC0oyjlugY+IxQA0J2iF+pty21zrosAv1Y0wcOA
gcjogpYsZtV/tVuoHZXQ6KIIZPWo0174lN1rubCMBHJvLiYjU+WUxzj/wda4vZNt
QzJGLA1MVrqCsK6mcAhjLNnYKd6S3FPz/n2x0WyVcvg4Jb7dS8FjxGPOcUuygtg0
JDdSbRozJhfn25Xt0qCbA8I3YE7yckol6YVNreRuQOOuWLeyIEBCP4sbkLJGibYE
xC6V2uJxnR8bxHMDTzGqjOdF/aMGCw/8/FSHOyywn7FLENMP5FJ8ti9Ab7bYJGih
VdIHBsyulYpd3L14mrDBaHWuRMPzPB3/OOP8lkn5YTphrN2trDMJjxT1iyZf9MK0
yTdkSrxFHiKu7sSiQdvR4whifi8fTMA5eCqDuLWm4ag5qSgeW77owzz8zshRBvEq
gXDU9DkWujTsebO5Kp8EyPoFvk72NWW5bKtnG2UQ8HSotn+wxXstpttQ/kY6krQ7
EiGisMsuPjcNaCvphIGKU7t01ZLdSDIby2RquKfiFRDdr3ZClZRvYTapt9qB9H8a
U2j7sPiIaY3bWkjjZIwVpbJOlsxejOXL0d41HO/Rdm9s4GK+T1P8SeI4Lyz4mwaB
6/5iMjhp19tAYVj8YitJPIA3vevWUxVGl1oBnmpsL1MalK2oMwRZCD4QxxwpW2eV
j+glWr5trzYNu1eg+hQ3qU8q2wBuaS1EdH2W6wWVX33ThEKaNumU485qys740530
naF140QD3zbQLovWgH6ZFck5+f9OYBWkwvuTt0IuZtodgDIvynVvhhOpbXZu2Leo
oc9+jiDg6Yw7C3xlD8U0L8FRgqpUrGSbvtgaU6Akyr05se8LOfX3xT2c345ehf/L
XHPSENivIOAMAwOK7q3IF5xAn5Hshfh8Z0YYSMq+0NnNv6AUrgmU6NsRSAStisnw
2ec2EkbOo4IarB0kCimW8UoROqmZRPYFxFPc8UBjMB0t8SYXQXdSOJzPnS8QsYR5
UcVhbJw4R8FP2VKWaWc1EsTjd+t/el1h0zgA7ujMhN4OPbl5qx+RL7sMyZvU9ID7
+3XasjMF9cLosQBkUaAQS3e9Kg9y39bhkRSFEFa7+eSuel73GniolRO0fx3MEvVZ
dSSVZt0b+JH29r0ImVQT80A81waGbd44QsxIWwExqNiaDFBzk3Wr4orttJe9e/id
UBGZzIxI6DDPge9mdDZdhjlXQ3YQUVxLcLH3vol+kO3Vz6OXJR5SyUzkJNBP3MFN
wQ/51MsOpZepZPV+UoSug71TuKT51t4q25OsCRHqRI2y/x/6HD2UlLYujSuPkdSD
dk+C+xnj8ygGt5k2BGIosFgO0sKgUKuwmJzili6RihXP4X983fbS8C2IlV9ctoWn
h4QSkkCOmxBhUHwaayPmPIjatynP0fwGN9Uc5mDgMBajHY00s5bzF8LsekayqoVT
z9wEhRpW2ogjGBWgu9p6ea2cTDvJgoTZn5flnvDR2UhBvKHmH18hgac9L3RlDp25
ZuDLxIKsqPUZ/zx9Qc3euaL8ocpM3EpXgsjgRP6Xeq/xk5OX8VFTEnUTHaOlxdA3
lXEjyh4Q6U+RegAZFvsRhj7mkEgOhWQTtDJTxSwvCkii7oYlkV+G9mL13UMJMLIv
wJT9qoc3a/3VSvjKKCnRObU8Y5Dx+GRO02eR6aV184D8EOFnYBa8eSH38pJ3Pnkz
pmgq6nt22ESYrNuiqrDIpN/CRL5qL3sPIE45U0BhX16Of045nHL44RbPAAT9P3C3
Emx4Xp60iB9OZFr2d1DCQLPJ9jXN9kB5MpWJgn43A+600NFF/s2pbPEVCYQyZ17W
lcsTvTwT01J7NYeEAFSjZiw3Ri95aGO4DH/1PEuHaFV+jV74jubYJvh4aiA5kJnY
3Dc6ivArvry+O1Q3eCS2WQlcONqSRzZMVx0vKjf2vgnr5lCuQx4JF2q/xCVuUKwW
fBWouqs0+gNCOyzxiPHZiG9sXh1klTPKFm3bmsBXQnGtswXb9Bca4+qYnChGriWl
2ajXUJHx3rRNFOJVhHWwZDbfWdeufz0k5ROZBh1S6I6gWWtke5GBqNmOma3oUQ97
bbG9mtJyasXrBErNCbEaRmwe0dxzxZ4TFr9GqcdgA66gst95ufD6sX+v4fZmY91c
3SN2becq8hUBVC5QvLzsgoojrt+xF5qi/JdkOAjmCsOQWMEtYyWlwIFvyYsJj+m4
Xa7lOtm6oS3XSRz/ZRDjtAaapjPOcZ/lLrKqAoX4+v0GbAmOgSnQTQ3qhaiUQYSL
GGV5WF413TsgrpPPW9KwV3ENuBrCMPpmEBpy8Z0O9f4BnaFFiWJSw1XoXIiELt1S
0GRVs3hlh1wL1jt9k4TZYoTKezFABeOEfWgu4+F1z+1EU4iUB5DeNVlVBmldyE/z
QO1lMcpgvaL6F43xPNl4MTz+GllbWC1zvpdxYRaa+hRHcbWwyWGEgh2BJXcEgUla
n5FGX22ky1GBaJa2TNQJIFAAedUIUtSnFuEeC294ksKRnA6NGx5VaGw02nkSpt6V
KQzdV04NaxGjYRIUks+Wu+pcjjXoqIP0t2JmFaVBaDVANsNs2a9ZB+VQ4ctI/CBV
CgYgf1wmsIYbQJo9upwrQhO6Jte2szi7mINyeYj6Y9BRZIeEZOA9iORlZSdR9zZt
OYACtLha4AvtJCI5RVIR0/DTQ4GLnLYfFWsD3qfMt+JptobU3HKgTebCPF1jl4+a
1ZfYgsi+ToiSTPxqgLBziNYERUnVLUhTa4oNh98IyR14ISC446E7rsTVaLHeToRk
a9vmV9C3jjACNFxvzMSDOiaWKxO6a3rCDUVVSQ3m1RlJA1XKOK/UczfRnWydjsw5
7iFl3jNfO9m75wgH9UV4F0amx/mD/slbShThn9TM0P/meHDjW5pQuCQq175YZU5X
2QEf2POH0bs3gx7zw+rgNqBMYt4+VsIFnGq9iAplRKfjqrPHOPIZrcMIi+/cwj1Y
8AfyewQxjKpAGVQhwVG10uuRbN+rgLCsW6qJ6rMybHqDZ9si+QivmrOuF2x2mxcK
IvHsIPd7WhWMrIleL6268YNx8f+R4dhUvL74rEygKvFYuETwZGQqe+ax37GgbsD9
180zrClvsmvYh7sx/w/fud4Bs4EKBkcS0Y6DVr68yBULSAi/B6fIUM11QkqstPd5
xxakwKDctrcb0r6WVpGp5JxqmD3XG8qJwxQnPOxby5BSUdL2JFH2eOOIJ1fOar8g
kk6qRHTZTxBotXlvyVuoXATg386naG0OxBBoJ45sqAfx3jrc9+vC28u+l3cEriSy
i0/HwM8bjULcpv13QAUGgQa+TSPBvbR+Ki2evMStrxEfZ3AWgrzznkeglSjJjMxn
uHJnz6O0vfEVzJ3ocSqfq2EEXCEbTMekzZIiw1FhDzpX+V/HhYthVGUz/HlGaeWp
ij51KRZ1q0UbyDSkY8LHXHFv0QSwuVbkpRGveHqEz2aivw+CMUJjpNIRgHLmPjrQ
dACH9jgXr3MNTKkPliPJNo1JYXHIUgaAffqWC2cL9fuqbZLa6mMdf/5IIPqhNDuc
rXxNXxiGxFlP6P1rDRp80oLztwZLEznkwwRaczc7fo+nRRktzYydnrN6N+gxE/V2
1Fw05uUmU9atQByWt+6o9VaXuo3l9UfxyJEc5bWSH2thAI3sjqaeeJFd/Ga8m1iw
czz5WHmP4tGxQ+3wC8V8xwNByzuLb24Iyr98pebySlwGtSwxtTGJYGYMs2Bp7zC4
JjSZeTg7RmzpwpWsJC0vK3JUyd4qFy3zSZOhxlIrafwLkvQPKpR5kIM9c6cCs9Nw
xZ9lbAliIPsBw1SPyRUNmYYVjQ0whh1W4iV1tNFnISsUq1AHWc+CJAL0wgczCGDi
lIuQSPmzNpsHHx0VRfoKMppwzsS2L4suLztWTYnd0fJjwnwL+6IUh7yPz3lmQt6E
DgL1+wNMCtInmYri9JHQeAwOgMHBFYpB46szHFZoZz+j6tmn9AehAtoP7CukFOSL
OzCeCTgzsRiat+8qEQuunBNB0yaq2d5gprI2APK5op2g9hEtAFcfkIGafnxiLtTt
t75zCGTfsO/+riPqC31czPwOe1+4wc3+ngP4TWXEKEVlsPQtJx4Ze0u7f80N+wIm
fZkJeyZL+bD0O8YPo9M/WB3Pid8H8mzGUlfzibLbsw4OVmkdtlf+7gpgARTUYiSc
C6z8yNk6vY7E4HvuGyG7lGS/zd6gD7s4/e1JtHJI5XZGlgoYTtuqKJ2Ru8l49/s8
HQBkIlntSqBSRTjaB9/1zqGEvNFuK3VG/OoLwXuv/+cmFplu3KcTFRkMMOwmdh91
tFPeevd8uVaXYvvaItfCGZMDCOe6Q0utoBC8qd0h4PdYmcV+ecUJDDt/CldsoCzy
RVVW/1YRCFkfNKHXftoXDDLG8FNff4jU7x+57mNN8mjfrfgfDSfvJ5Ma6tented2
cR49/5+raUZQFQv/kOQI3vENQhne9B/htmFAVdmp37UNGUNhXOG85bNaIykROZCq
dl3qHzWbjo6sg2yJ76DG7qSqAtPBdxEO7j6h5rhsmypGE6NxOdF8x3qaS46sSv4F
3Q9eGu7YKoS1AExlhat6vr/XaFloD9Oweydusqq3o5UdQtSvRObcaKvZKlSxq8I2
ozfuwjop+cQaoWB5vvJidorWYcCf06tSXVmpQe/KcCqQcKDtRVFQgpkrNOdPNS22
FeSYfsP1uRFrJgASRYH3N39ahW2F8U8BlXuoTe14UeqUKFgJwlMN5sxJ2m2Mf5IE
6qVlgYbOxCM5SCtNJ+mjMMo1AfKs0hzJQArsFMUC7lSRAoWpHjrNCJZf1U2I2W80
XrSUSwSIQ2+Ef2+rw6FBnlfdUaeelwFVbpeqEPtsOqwA8SYPImkWJlF+DpEPTs89
01UxDezGvwcNCPP6pyIzJ3YrRvbPEXnL5rp7pr1e08Y3TF98zu2IaDMKoVIbYKki
NF5Vqufbbp2pATT92aG51RidpjN8aMq15bnCmnH09OYRZORh9pgYHpD2sG7jKdsC
FXhUiZWatDR0Q2fuDXb4f6xE0F2TEhO5knq8SJHH55oIdYDpP+SyWLsnW55SRVdX
9bLyKt6JuZopCWsyaCr1ZA6n0yEwxV2LwsWySblSblbq/6JNx/vG3+xwssntaIrB
UgsLND6i1Ie7cqdO3xfzEIsGpg6U5lvhzf/3yZXWhVP26+P+/kZUwNfww7/f3KQ0
ybd7nU6KnY8/FZg8e1MgPPienZaSNAVSy7yJWTtBkheCXAmlE/mlzbwS99t3Zzyf
Zgt6KlRhehfoqkfu0KENea7jo77KzlwfdIKoRRAQC+56I+VoMubLCsJVJLmadqfn
ClJT2ZXDcNhD7/dCI/W/P/8p/NTZ/JRMaCZTbz7yF5ZAUtPUZXjNvaE2RVfXs6hR
2sZMNf/Rx66xycq1ObR+Sk6pLhk5qNsL35701ZuxjHqZ5lR7zmxtjxD/kkZij7JJ
diL08NxPCcO6vHe78NzoEHS4NUDZNxVpWOZCzqQ4ON2yEwSnw5jNe2k6kI4oZiCi
JGrSpKRD9yns0LzVMqT5qFuQeLx84QIuytp7QvEhySVHJUKCD1dzaIrWgDhGy2Ly
XYSDKE663S57wtia+TVLLZQbdaXXXGW9DiHmKSd5603Fbj7qOmcx1XlNt3cEsYef
sXunmFiK0FDxb48SPfBE55XvEeC0wG0cdTPBwIfIiqZIFVK1+u/svXDqpttXCc49
FHZW5kJvG7GfUSh4PKgCI1QUSXWLirP+e3Yr/5B69NUS/dhL3AiDYr/RmIAmPdPO
erDM6VLeABQA3c/JWZb6GwKr4X5oisWG3x9ggVZ1OCdF/ADy5DZJbDuh0qFC5WiJ
PskaHz8qci/ZdYhbaVx065Fbbm371YSeXkP3Ox7YSacWGbq/qviuwnxQ1oBYGRRl
KN6SQWfPRJhQzprKG2ObqKBVouqH/AyjCC4WxVkFtFrrmRWkGfkb0S4vqp2YSyKS
EjNtH6z/kyIHzb5q2vgVT49MmIOt8DBkkdjXmboUoOq2OZzgsuBhrGmalYCMDAW4
dURuGJ5TWTDXaaF+VcJqvnrDeXL5QwACboKrnL6rDS6VrmvNLOBpxq555nD9Lm1j
HGIZS25VDCWNkYYKOhMBLtZSt8KuXF9OLL/Zm+Iu5GO16mmWF59TNRgZcU63AuUI
Zlutv+A0k0RCPhX/7tBjB225nMO5k1I74rim6yZJqAy33Sh29fo9WHw9grvRVz47
pKCtwj/J620PDCo68B29g97EMA3RXc/12EVcpYZ84yUbcOpy0ZT6uCXti2tC6e+h
2/6eInLMGBzMJCpYBMSZ8ID2SZF4Rmz6EgxlzzKOA4OzmSDDSkVyvmbT00LkvN9z
iAc3z9tNh8kAl/uyKVQ+9P+RctRJyd5aIVIqNHB+lQ0W1bOgbfsjl5KXsngYpoR0
igyEscF2BVVSpU8CzspDUcvDduBaQ3V7ymmPlxw5eBuPHmF5LhM6EPuogIjlyBRW
B2msc1qkUBCCsdh5Wd45NtjuDB2zd7dVqwwA0eTN/BiZvTeN3hmuoVOn5OR9rlTV
bf4yxdMQLbaZSGVEUtrYKYuqXegwxjuC38P4daebJYJ2rybRsNrQVwkFUF4LlKv5
cGYoZT8Z2uOVEOIQ4ubU2oSX+R5p5nPplD/gUEGsP1njisYtUAByppP8HtikoCkU
drMGCk5sE6uEBXsagVyka7vLiHmNLrBcIiablaS06tUcPBqzkPP6WLHuUNjlzrDm
pF8+9B45oe66k/8fU5/PVNz0VHmdLamLZLLKmDEj840Hk2erpbueYT2pAmRSpsae
8PAiUPNgbkq4/4biCI+TCG2QV7PKoCpbYyf6c52c8YeSlgKV7xkQLCUCw1ixagye
xFhVbq8WaKQRFFpioBfIQ412K24hIXUYWDHZrOZ6YbU2+2sKXnDSLZVFSxGncHIA
xkIletBQKwXIGH2Pd0iThG+aM1HXWNMiRSmnVrg9TBtomvmJMfHcIv3Q74fYhzQI
S9D7scnPcfW5sLcWO6nYTJ0Y/bIBcLSFHijlyk6sdVDkd2aE05PI/YczpkwyXiHd
FvC+Z+4+lfZKLDV3AGGsDuW7gQcYX2RZr4V/3fyOEeCAlk8TMKp48EgyXqYx63J2
zNgLTvWaISnNd6NcSDMwt4ghPWPbJIZAd05Jl7OvjL8PZjG7wHVRZddM8iSoWiVC
JLKwwf+HOHRuyKZo461Ew4MlUUYvTFsHs7xVsi6bPu8NYEQv/68ZB7MVkC1xhJok
Ue5gpOeDceqityUDRV5lPzCnF8cVFq2QuYcJRF3gUvEdGDiQiomr+VWiFxJv0Tw5
9uy8V29rD4lp48M1375aEbiQnVkoBkSc2A2sWqBbvW4RHTBY7TitwTYdHGecH6Hj
8LnVgmtNvcSw/EbdlyJUwyhOouOtAvw31Q+ew4swN/oTV0EB+YPWzPdMFzvZi0aP
ITtmzUa+szROjKfZQg1LeudDeqN9jFTlZXxwfeBX2V2F0jXGcH8Ein9G4d2M0+F8
Rai9lqEmWrFgvVsdetZIwhnKvz3E8FgrPZKXY8g2USObKqh37Nrn1Gokm2mTTRf7
SjZnTtXS356w/tMjHC/ye9InGN8AgeO6U81XOOKBuHrFyAlJF4dPzR+jShZcpvR+
3MzzbyCxN24b6NpIM7Es0Rxw6Rxqn9asuGh2bGdnPfSBu3IsXEql2WON5Yon3fLj
sDOCvT8bnVhO/IzTEeY6Idzh4aZPCu/OCagwjYRCFDn80Fx8WfT164jfkH8+2w6K
ZunkAZyuekI1kJyiSMkDm1rcdWdTCrrKkLB28Aqh/d6uzpv2Dp2Cc3R2wada702l
Q0zFQ+jOtnDwXcvjAS6/rBLFsPU6mI+G/0OX1roo+VKSWth5pH9wAK/W/NSxtMm4
v8RX9qi/3Ykr10yfpCOe2LcaoG7QOrjUFfBNScqaN3OgyCJ5n5xro586fytvIEIl
ZplZBp54nhnRA3/ptD0Fg7WMkne5lWrtdChzzn/qJtB1ygULymgIZEhcKH2J9UuY
zSYO5KuKAtAjhiJXRzZ6A3cSi2/pvWfpzaE6LpqxJOSqFkNtm3Rrna0T2QcLMY99
CUHqsvWYv3rWgbM0OWGl++8GkdobU3ubXljMQJFriimUwy2GTimKk1LBcmlrgPNV
gYp4WVUAs/cJsH84rw2oFrRIWZW/yG/cPLX2SCI0htSzgsbBiTqxb7zmhyYTiWzb
QIckY7VbC9uL2YpMIm+AzTWbdnsNY5qeC54mk0UUQXfb3LBKVvbDkEUMvWsQYJr/
lEYbpjXSMykKpEjSYkTTxnvNfaw6bUlaE3w2FTypiT/HUOgJ7AepVKQqQitiK0Dd
70E0k8sP0ivHKqCfUwzKNRpMemCiElXrWZQtAWSiPjZEycu/dv04WOZ1sfAsUfgP
uPfred7gJV/zCMmWEJwIpvMoS36XXF0P1gE+7UvoeaxZS23kqjjBleIPMIv6BC6V
XEbPg9+M/6pZSryFAo52JrA4HN+HGSGG7Ud1gymFRGzygjQC/8kHjB2HTRpd9CUt
lxcmaFsyWPp4ckwou8HgTBSFKTXN4+6LxZTMCrZIhHU1REpBu/vTPMDUdn5zX7VG
/808STpXaUyBab8GK9UUL4zR/Qj339sToX3wu5rXlLkBj4Znt3v38s0tq/81RY8G
J8n7qSxp45u/T6gWM3NOBRrLo/dfLw4MXLm55H/iFNKRxznhjkRYmBdD2RO+98mo
XlnhDTsJ6TLzZpthozGkAYoS9zy709koY2RhGCedBbxT1o9gSf9tCfhzewa4mS25
lZd/xQfr9lGDb1QhuD7Psf/xpkuaDTSDMQS13lvnIYK9B/zhv2/JwQbhrF3VYO9b
L+zj3YqdrGmLZDTZbhVYorA4zI8vKpDO8R4CyYboV/aH/Sakgc0AffLSKl/xIL2t
O+pGg3JlOi+DU1oQqeNOqw+bPeI92ECaT6w7u43tOwbkzg2wyNAoBjTzTq/xJb0i
khpanSspDYMi2q4mqk232uMwKo+kQenz96MDxqVOCTHGIQIOFnrsOmqDKWJwDUWw
4iWK9qkzipvQdjIyq9Vezv2nAHsEs9w6Ypqt0aYwzJe15SM88wBJcSThO8pj/cj/
F1KXWrM47x+nKm572pY1C0dQJNCYze//JOefQwvP/C9KMZASObAq8KhZYkOgNkqR
XnHzvbGMqxuXAcMLL+cF9El3n9St3a9NlzYU9oBtZdmR6Gu+8Kdw7CTrM/uMYelK
Uq0rUDDk+7vd8IzuGfZGGR98d6eJIhTL6+8YR0EnakXZ6UvTpuQBVpt47HH6SE0w
3+BmXCqCIDUeMrRdRPc+l364PtxnZVtuPruPwDSGmCScSE8WQ7UgQLoIeEG1yRnv
oBLtHXD4LonpPatuSoUm5WIFIL8IBUZ9V5mTET+wRSTxFNGAlbWXz2B8o0LyxAWq
hyjYT97RhjbRuqmejjCXQo1YiEs/fDFDFOblCfP6JrlIryok7JVWi5Wbf2TZer92
s7ivcr4hNuM205/EUtSHlXshEoVSghyTYRrfQr3m6dN6vD7Avk0EmwkPb7SudKi4
2xph7yntX7JIZceOtWNRFOZoFIvEaPbu2kX3YqJB0L1ge64jRR4HmDdM/QC1Jq/f
2swn36qn+20qBWMjZc9I7f/r5MEvJb4SFkLF/niLcmd83IT0KT5ZyIpt+BJpKJAw
EUq9KwoadnLPZ9fvruwjNEeZYdY1C3HZIYaJ7QY/PKzEWo2jVZzAcIQ7bfyoeMEP
mFE/IjnIvUojawY/Y2OgT1pAQtaCZix6qA3feA5G+AG8od1G0Rhe88nNNhAOuU4Y
iCeX+RIvK4WLHLcU7Lu3fTBSRRWizYCcINxfq7fbuNahEMOGU4BGfkVZbMg3bjFy
27g24JsbBcKd3OceMm08aXGlbBWBJ/GpXTqbEhbTZTXoLZCfX04zisKKpWleGwPK
25Y+zogWdHWDMZVt0eez57+t+dsPiHD0fysKA0XlBSmVBOoMwuE6LVjuFZFE7nRr
CSAZ3izwPxOWdsDrC/z2x5S8LDx3exqbIyaiqKipRJneuodbaNSJTTsinQ5uFoJn
CtMD30Fe9/WIuiKhBopM65vbSEu8NYvCFAmYdwoGTI/MPqckTA4/yIsy/35Yx8yk
pWdYUGDGNofhQjTY5ie5rS9cWzClRwRf8CXqHlmFBQqZaonraOSVpZRgZcWQRnF8
drqrp7I4e2n5QaKx+1QH4BW3U+n2v92B4/Si1OI2bzL67nSWqWgh6BP9KCZ4dkE4
JgvFF+pH1C6JsNvLeJ8cF5zgwb2Fo/Z6Kw0xf2/2Kurcqu1zZvpvdbaGkR2JwyCy
JlDgplo5QjcXSGXyt6IxYjMqFiV+Z48MKs2woEG7nxFRuswsgRl4z6ZwtinKz/7S
tMA5Z12ArkLo0KydWM7d5YhUuYg0FjjiO4EYIF9tegMxkNG1881+cuL3ewCF6HIC
itFPs8HgZsnnX80w5uGViMFlBaIeqWlzuYxbm94QxnT5Q0LCTfORn0bvhi9+T2ff
NeXdCjnzPrIIwENJML2hE9FHfMcHJyMNBI3eyFeCCq9RrmkPUHWNVScCzMLVR3mi
KdT4GkMKQwrCb1SR5q6vaQ6ux8UwVEcIkqyUfKRI4f0u6YTPn0FnN8wcBk888GVe
cay/HGifu+EowUESRRcpTsGkWYTygfIFTCGfn0P2iZ3aLnr8B1kt7urBEol7Ri9l
CejtsAe0whSpQVBdTkPYeg7S6ps5EyqsrCPIwmceMlsnwzYQhbixNrTb6aFg/F6/
xUkFAd5zGbiVdKAM6xBjSb63HW7bWuj7zDNJgqjoiko/YqUynHJHG51hZVXmSvKh
siqPjw/Q4B5F0LagzIuCUGVX45nMslcHlh3YXziYb9z5x2XSIWH8pBwDqLgSXMzF
J7skK/XTD7QkL75zo+RWCpUdlZ8KtTc8WQGPvHRueSYWtdXUWwyCxkr7IulGEzqo
gkn8PLQ1mCXeiVAOyHlqJv0nBrGRhe9jViCvrh6dMd7SxyfsepzFNjTaTwimRwJl
TaVATLTcB5EKvC4DjZxFzo1mtVh91msbeA8EgJB4O5eC374taUma0y1tPWx7Mxkn
hsQAmkgx4AsD9EwVV6NTCerk/vMZg2G3/6Zepw6pPC3EVUbFrBYGfBEC/gCICuLm
aLwlVRZhepUwRLLJJzvPj28BlAZHND6N6d88ZtT6E5GB4sjyaS00jj0C7MflKxgu
qhvDKNCBJNCESOemclr6nP0FdmPqKH4kithrP2WAl4n2JT22lrraf8Wn7tJmKZ1I
zEPpoi2dz8JYcqcluym0BoMtROi2tRTwc4lSlON0J5wcGrh1HgSREMSOy9aIOyYt
pxDN7VsrGcrtbwOJYbiB8wNU3iaiTrdff53GmokNh3P+z0E3cYQGPONvbsUPky7O
NOMDs3BMfGPtffhGFKvTbNoLVa0A6R4AYfLp9duTG+XP5uz6SPxYJBR5pGjl8nrF
qXbEJzuT4QnHcymM18gSQKCxRVrmEhFZVZpekBkzFMutIWOW7GeFHgazsCzdj+vr
4VHevvQQBBq0YC0hHB4VdjxBFw23hVniqxMEHyLgBz1G2XDK0sxK1eJDNG5fEdrG
sB2MOEp4nFSfas+wIsBHfcGA5A2WFjS3zSH+HaK7Q+rIwQxD1qJzh/zeq0ludMCs
eifHco2S8S2l+OE0xQIJynAh1RixCDtd7hzmO31nGJ/DsJJu2feJjglGAofYWpi5
Jz0z4KQUFiBZMhsoml5O3DlDkR3L0TTWb6HU/ARSKqvnRqCkDmm9RtxOCQWaZ1Au
8GYSXv1SeqbtVV6vg4GwwYjCxKIq0SftWA6QQST8tdYJTVWf+R9oAReKHpNLfrD1
IPRaL716PUSjTHIYD5hwu2TTtspX8pCkisdlzOOF+Ak/yru4V3GYdQZxHwlJjn9y
C8LVaaK0VGU/owmaoqqJrw/tCXZEBxzMDwZ1u/oCOilofvD8y6UB8UBQLq0MjJGa
JpMwJGwku7EAfyWwKTapMZuNOkIntpXV2lOSuRjD6pfxz0zK1b/0pLOygCsFhVeQ
zpTjxbdqsgZOotRpWGNJkzyY+07s6nq4kfHNfvz8oer98Yz0NIFoL6YX21DrApjE
MHW7DX9tji3QvF7OQXX9aJ7anSnEFTarhO2VLN34j0RFl2wGk0Cj6RT/qRoq63tR
KStxcrdJJooU6Dbai372xpti8vx91duR2dPGy1HPEMJgijwseYBQ0plFq2b+RgoB
VRqvXxs0K0RKIYduT687SoItrM/67JlNAh9+e4fLGw3i5U2uxVktfDnqUM2NOwkD
ryJoo4Mog/32pwnhIbc3FYgRmkJLPFvs8NNtDV9zrYpChEv2XOAXnpG7FAY6MwBe
tioaP7w2Waw1h6Wt5mGFaYGulwXVcbNUggn9W5PTe3kvzJJktodquBReoHAhbfkt
6mZwnSzdlDruSV78yxZ8SbkP4/WAkKT93wXnxm92Z4bN12d8clU3HCsIFCKoDZmM
zqieLashorh+CwU+5E8tlMFPVVR1fGfb7mLbrXBASyXFGqg54p5lfMsrrFy9+BpE
lzP1r9YiT5cptNuEIrab2tLPWaeXWL1zd4q095GZwu5zFg5IJ2LUBGMwuWYSB2n4
c8ytZkiHcyGGOY6jsKlRaQuqkBerqHdDjVv0dEjrPwosblbwigJixeCmibRG0BHB
Bz2iSWuZlzwY9vUUn77Uc8rDEvgz3k/Yyqtb7m14mWtYEYz2lTAwG3V8W85uHPjX
F2RA9X7j4y0ssHVXydDfREXtxBaF0CZCu89B9jsPV01rDgZP+tqTRfmURzxLNeU/
gUvxqJTCmDZsYrcnZFhlDP4wtGvN+2GCc8DE5OPBSDevmRJh3flJT+ofJPY1rbQD
8dQTZ4FrH0zVtwF8A3zWBlXXIbWIobLcwZ46dZ7y+QKABANaGsG/8YSuRJ+OX+xW
3VCUAeQP4XU5LMRkDJWj+b7sC7jX9SyKqokNlIGwdDZe0C2GWv/3k3uMf/K7m8yj
Xe6rRrsw9aJcqzKtpEpAS5uavzhmkdBXt9lQYiP9zBgZBSxHyTC3O1D8p4P1+vuY
aSGPU/83/eS5vutUwQmrGKBosSU+6Y8NgmNLuXR2KORlgXYD8xG8PfhF/7n5xdGv
Y9YuDGI5yLDTOGX8HHF44CXJAmB2InG3c4dF0ZMKd3Q5qt5HcVd4orAj9N0hrlt/
CvXlUKZRnnvuLpfYaaDCu7Oh4n3O0zyL/LMh1TDHDJRX7OhMjQj5sszQzUM99YwZ
d99NkdkP65rVLqEDdCHW2EkFM8+AO//mYYv5d0BYxzWpfd3JKfEGfSaVevgwPYGp
CDSZ8Qsxp2BdLLYqeRWnWgnv2vza+UanGhyoEIElXfh47PYDN0ilVuVQgGQOLXQ2
VSLxb0HVKPITI7z/EI/DHIJjH0kk5ebZc9IuIC9DRQW0G5juIHYF8v9HorSgH7k7
yfU964EDcxpL93DaPgwzXw5vuXsJvSe5Vr7yrG67WpGfMSr3IJoU46XNakU6sYBS
nmg/Fl9YxXWYMG/+YJEGhFx66tu+Ktw8GbSMNczcVaBrPEiz4juAte76xfrV2nxW
8u93O3Zza9U9S3KReQs3c/X++N3fDDAoqPJYdOVCVASMNkdwqFjiTvWHvvzcBYPq
mi3mE0R5deXRYIWw8NSmx/wSTwOJSZay9JKQzG5OSfUpu7TOuWUFMJv/ESPTms16
ot5geakIm3v9igjY9kLLs6HXoxEFy2j1zBQfmL/o0Q4Lpp0q7VhTJNAEZXIqcAVx
p7bfmLYHEhI+zY4xaWyWz9Z0dat1kJmqH6iPe7vgzGYjDQ9Ibysv2+Ry8uaXLxw0
WRYXOSoUFAw65+vI2wWGI2oydDM7osw+5h1JrnlfwIsfgzz1yXygzGZsvxBYAJpu
bxvI0jC0dlIvdSKRqUSKYgdBP0F/auEIlAWXBGGjSjuxiloFg4b2pl1bidsMGq0H
FWMO9mo9h3QYhh7Yjz0kVbqIT0iyqg77tqgnpbCFy7MFLzp+KTOMpAS1r2/BzDlm
v/d1a4hti/8XushWnXucvfXgXuIqlyCC6VuCURDgAijC+1VNNZcwPk50nwcsgxhb
5AndKLnWTwutYE8qnAiBOGpy0Vwzf/z7C9666P+oy8R+OTko3XVB6IthClWTizgi
zpZEfsUE84qf5WDDMvmbMp+/7nKOR+b6UBtTAAy/WHJqc0ynk6N7hOYQ0atK6X6E
a9Fk4LtfAg/KjwoIYqKtkNRMHtaGHSCA5u3mXFI9hjRHege9nBEkezd5Ef1PqW70
UKL+ka83io1us9oxAKbovM+fJV1bAR413ywiHvfNef9sO9xSFar9A0Vf4T6G8WAc
9SXAgUWjRIjHppJ+D6Cz870KFnafQXzH7wwe4rsiDepuu25jB1hqjMMIfp5O8eWZ
l0NszPYS62tzxNERMJtzvqudy4MiEg9UKUxLi8a6TSn3eRBzJAZJu6bPFUFDc9u4
fKc0dAcMJKWOryzJusQ5ufozBKhcgECb9isxF2tQQhhqR0c/Ng9BsQnvosagmgb8
G5bQDdYJXaKuosaviyLMdkm7gEWPlK/hG3Cg1zB8tG0rLod5pMPmoKvE6jGD10ah
QnjkgKGInaHnWW32/VA9/RNvm1kH3bTN4xCbegij2UYLifHgnpJUT/VDL1krsUtl
2vEEdky8xuQp3rRnQtU0+RwIZuQruLkmiHgfhE5bIAs4p/vuHqrsbf6J7L0gSsl5
r9xBQqxhs87jU+LCAYYr2JjnhAsRP8IPygA9JrtrfZ8nNlRnj1pODP8uax1aTvbf
NLnG0sVjJ2fWjoCzn95kgPzIbxCS2+A/tbfquM9WkHqdaB7CP+n/KEeapXALAURT
oFVOC2NPpF3pgxDCPImVKk2JMGtYBUftRdcY2xGfPX0ImCfJLoLy0eyO/iqZjA4U
7DwMgz5XslRG+WSzAjNo/cRlO7xjCOeYVC+YO52aHgNDsY6TRvhV3TPoJELhYja9
DrCKXaWLAkDjcbHcBQanEUDlQ2DNHAlS017v9e1mKkui9H9DItRCueajRZ2ZwXCY
EldKyLBIlQxtrR8BYT/T2lVvX+90uy3fHPIj3wKYQZA4VT6bQguyKCwwPI/grnVO
tmX4hKohriBWi2x9gSCY3PPznuCvxmq8whQ34EZtzbe9kaSzUM7Vl7qR52Sfh1dX
MWXwLBuqaxQz4sBl8TJ4EfDf1DJfJJoouAsadQN4Ys+d8kHHUnNpO2suOjL4xVEL
X70yTYJcS37W/CX9zgrul7IL6psVHzBaIujDjAcly3rvz/2F2FzaH4rsuZCXFxFD
Das/wd9luuwb0qFvru4r/SZ3tV4CuQQxhLP9KC066BA4DTl5qWofvYINdoO6Yb2w
gvoaDyjx9zQsRK3ru/3Ytcex5jJKC9+AFRm5R0Vpw+vNUDXmer+e6IgZtScIYoyO
S6ZzGxet0rK0FUODCTq5OQwW0UdLkXjZ0JcKZzpBT+4v5WdSfGuKPRjKFItoufY1
OdjyHPUGaWY19mMI61JG3tk5Vm6HhcrLYULdZlgj/16eQ/lEd/KoZSBvQQIeI8iZ
BaT2wiI3uHVx83vy2D3Lh0K+tpAU71yc7JNLep5ZMP3/mKhXKEduvX8p8BPU4JLX
+SNXcqKNTir/z+glmt7qYGu5+CbtfImHQvP3ZU/QgIg6PTdtv1eiK3H+rOP44TpF
OddAbs2apCnO1Sann0q5tfFERQ3Pzru19kQ5Q1zk5dTcdmEI9a5sc0hVvFOoNhr3
gYnktrbV8BJAjGBKvj6Ui0p8SN9rF7Ylzu9PAk48TKnFxva5Vn1HjVm4gwqeqh4X
uVJIVjuQmArPOXrL1RHHc/v459lcV4vDHyWgLZBrb0Aq2vVLWo5ycf9pI/Kl5Psh
vQx4hcaNl5yrmig8/IUT+Abn/AiceNtrs6JLXN01YZNnS7XtMufo8YussRY5DAE7
YOCMCSYrCxCt+lrYX7FIq2fFGJUBOXTSfQUagOceyvcpxTo7WDKW72W/a369uGdp
b6IE5BNWKndH4rRa5s73P0++JyaGZhcuqCx8GhyPrX+Z9mWsAbei49PT2ScyR+Kw
rwlN5TRjUObdrFmfGGH7F2gNXlvejuh8TWAJK3H9Ogjg+htHuhPNk95UhM3TwolD
v4UWMWQca2vMpLHB7iW7Q+gpM1tyigEFsLWSfSfNPMPwmCXPxySemYGhCRlLZZot
AWlSBxH2AANOOl5r7asB1CdbucfvhkfkwvxWLg8QQwxNpbiIV8XSrwvnMObvFyfS
7APO/ElGhE7nk8VpZ8G6gOcZglR46A2ZWbZ/gmhKYrBeDUmEj9GFyHFDLqo2jCm4
fNrb6ggck95TZdd2q157Za8I9HR/U3wccE2TRXzvISo56wuUdl1F50zkRfk5iAW+
BIbr/F7+eTk2fIInHa6NbPKVYu70Ajrz0ETbYH5Ol5zrH0M4RPkyQOJYVyZsSrpz
0XZhkfay29NecFbLlBnSR+P34c7BCey3ax1Fi7lDt5Nw0yAMA1NqtXsnxUKzrkwR
NZxAzjdFdEYmvkeLlUScBG9RPWVoqeuf+moO3jxiKzlKiXiHO3GDvcvsmPV6q3o5
WzKxjGE56Nz5SFEf/mpSLs7xSaaQW2AJmBK3UbW3e7KqTylRXALyzQuGfDm0lodZ
dWZOE5I39DmnRcb45zHzSmydbCC7tf7bjjAptaGFK2MLz8UKqi7o6AvK50RyYOVP
h5eYDgl4o6qzUlXIDj2XehejJ2W3j/oajRMEzgxvdHX6E0azBiK5yxbyh8nwNs8n
9+uOANwRx1b+zPxbpx+iHObnbyPi60nzkprdR7Al5YP0P0EoKHnqH9salZdX7+sI
4ba/YlMrLxaWqBiOArctgmrxvBwHesbnMG8RLeliGF00wZNa/9gDYddhB8cNACo/
iluv0wH5pWsT7cV29sK9pVSyH9ZNnnUflyU0SOyVezbJQGddqAJ3ieE1H5Et/KZb
H0OQu52ApaA04CB8V5ffLFH8Qg6F6LdrevUH+4sEA1X2wnZnWNHnw3POnwA0bMtJ
0f9Pw6pPe403RSjjsSlo1pNxYkFiEvoG65RCglljG7cP3a397zT1mVE2V9CUWPAv
nCKuKZXu8NCE3fcQLF3zjOPhPLH9NGzGLbx/6b/70SFGD6S5FHeK+H7yBHd5Zlpi
870bloCfs3keRg2qmdQqUXdW3pWxS+C4uWxo/dWh4Hr50XgMpjkj7xLfisJjOoNy
uPS719O+UkPLTOsQRqYk2gbEmV6fzg72LdtkLDmoxHkiKmer/SL3h/ev8QK5Q2pq
sGBx9NEFostfMS3tYY1E62BNyHyrM5nYceGQNPzCm7pMphxTqTffDbNtNRL3TaHy
901pdLRoFKqa3A7jq0Ihwo+v0510u/oI7va6FPA1M+4FT85OKaRDpSKpaOr91t4Y
r/EFT6J1Y3S0xf98Br5TYnkv9YfgBOQVh6p2WQtH+DaLiaM4rz9zbGZ+WzZCPrdb
vDNvBvRAZqN2ohU55zsv9/qLMXJfX1BpGISsMpHULPtvpfkU8Rpi8ws5xK0rhE0j
+pf6h8XmZr8D8ZRPhepCxd0cRkXgascCg8zzHI9xdPKFAsvSU33iGWKq+EWJ8E7I
fYFj48UaYacyJAwTKpYfnwCsji7LA16gNdIaHPUfqypnwtfc2R3XPWsle0tshNh2
haw+gfrCOkYUhBz6hFQL8iEFXQURnk4opx8WTfsdCwGJAe9U5cUcMoK/uylWFjW0
il7ol3k/rw2jhd7nOkQcOyZjL6AAlV+5AnvuombFJEnQkZDzgnbdplYUllsZYtDT
nFC7j7DYlLzBRK/EBiR0FL8ePaVtHGF1yBhMLkf7Wy3+7kZlfspYi363EemCp0BX
BvufzufvRz0w72LNh5uQy3wuGZOntqgzdqZTgoNOZlO/koy/V6qe04hLyOJqloem
Ny71O1qH2TyxNWwHcaOCTUPeC6G3YX9lXQD6MeCwAYE3WdMqBMZvNMycHaOTerAo
vUsiOS3qofwsqW5HbQ1PJrLKnTVHaxHnvnSJmMOYGNck7dO4e2I1FglN4tjVZAHU
9f0nqSiZ0PTAqFcLApW/2ZQ6rMNN96cANhEWXImNRXbv6QzbRs+xgdFrsk6w8Jws
UNyZc0so6n/O9qaa/1lX+hlGHUcvSAISk6LSiKJ39TrF1WuY0cjeWLRvr7w8WN8k
HK+ufqImouZBQYjPKmpJH1TVGoXEJNQoOZde9jfVXheV0IrDu5zia1u07KBXAEHU
gdb2nKlyjk1ri5g6b0pw8JW1fmx4dE2QgGFFSyElvsfdXe4ZtQf5dwp28jxQ9d9H
Aa7etYaZP6ltekibMskUh1Ixj8trn2AX2jWZvDkJcyb90eXOiOdZ91Zpa4tu5V1b
ZXlyWhK2mhiB5D93qF6SDxEsyGxedmdc4sY+nUsgm10Ndwa60q8GYzhXW1eIH7Sq
zsQSlSOOA80lmee6EqTMW/WoCaiNxcUfsNL0s0+2+CTkWEx9dPkyVtgaq2HFPcCo
1lKsqxoY9m5L46imY0TLhYYUDzWtiN/mfhUPFpW5JTlUFLBKon+nMxQ0t9hqOAK8
sNtBdkatqICWnQbFghioU7AXbsHO6nhoRYpbCo98GotOPSngWTR6k/mVYpHqfJxn
Tb2gxCEjZqv1b8KK1UCHuo6Fsgl8n5LVV7/4rDjBAr92LjTtkhr+gmvuODBXr9LB
SW1C+BGUgtVFzEn8Q5Tijs4QeRbdG6+/MtwHy04cbdEo9iEr8fI+bfaIh2RoHi5/
zVfDPVPsg6we1St7ZJdIsy5vxzQ2dlq9fgwPeWF+A9WepYbbqIYgD9aFb+NQ1R/1
bgEKeLZ2gZTP7tAdiRXyzJJKxVsMtgYjIQ46+RrpujyKcZao9a8li50QfS7FECWH
e/IZASI6idNVXtQoD68eRL8UVMv8ksMjRpGMMSzq9r7NREMBO64aXqn3w3U9YSto
ckOk8OvX6WaErcXGNH0Nhfm7GuKz2qTO53k4cvn9tqxkQ5xy6kgnFnHRqioM+E0C
zsSUlzPGQsxLd0MK4QgLB97Ljk+9gspsg2JRwPCyFi6ydmcp/vRkOZMdDOCRj2Xs
DFJjVorVJOYq0sIdx5dMvoozo8IXcaitRH1FnICtHnU/4lC1VqvATvzn6m7CGX4R
rHEOQ5zFKJvDpWJnpwUifF0FC+jybk/3CTeR5En8nOBN+zcDiHiK6WYxLCREsDof
zaFU47lf1EupP3F/rkroavfw8ViX1V6ILOXgtfbvtpP+JwI9eH0+q8fiD+JqRUR6
csjLNh6robCnU20c+wREvzh4KEb/DQiw/E/BRbEz6PyAYiKkUjMTsDLgFoTovgo0
Sdx6B1VmZHIIP3M9ywj/m6pD5Rr2UUzgjrRkccDgKHJJ+RIzcct8B60hqfuqokpa
OJbRn9LEoSGQxYaMD5CjL5nDlyv9NkxCAAMGcMLknytwMP+1+pJl+y41JFaUL0NT
EwpbQiv+MW749zzZOyarA587I/GLUMxxMNenJFXElYYSLvAUjTEiiWFXdFyFzvZ+
l9QyCLNy5CZzS74G9q4LQQCBs0VH8trgnCnwJfodW4NUH9MOufy3UXswuK8sLo7o
V+T9bSUaFWIsYG1aiKpIbpgFUfHyKt7PhvWplGRUHB6H+MBLY7cLhjgq1uTtrb5Z
6aPd2DcD7BsWR+mS+dXxXgX3zX5Cvrc4FqZFb5juuRQWcA0bfcGNr1W9c+oMV5Xf
97KhSKj5eFlknWHZNbw2VOdZ6LaxM6VsykCc4nliijzl02NMj1vHPjRMc6eSOyhm
F2hvUjgj5QoKm3bmJcoGTajKidxWFEp+CcV+4gNJOLiEWuhIZXVboZoCRAn34JAy
maaPQ0b27P2xGKR0cEpVbTcGhN+ocXMMdh39UllvYXn+eJpW69nDsaRH9xgZZsyR
4R/a0xmPvOFV3oY+MpySxvi8iypsUc07fn7wVUk5PMpnDBZJ9SI5SyE+CMByif28
E1X4Dkh0SbhsTf2XAMhkgkrK7eYtg32Cekc6UA/dVS/IRykKH1kpgplSmtnLppfZ
2s0gtiU08dfIN2ffTl9fB/XIVIBSN899rnXZCLvjYXv31BeLd7i2E8wEwElPlsGW
IPLrYso0B8y8+C9xn+nZS7Hc8YVwCS4VAXJZIN9lRTg1+GKRXydDqoV3SCoxZFoV
I1tpc2VcgNPa4P5gQYNGlUnFj2GnN9lTnWDTqYnY9hmOZIs5QD3fAPvOv4sfMGbc
FlxOfbuPo5U1AIcdeFZnEND4yW7Zy5wNYs34qEcHQ/rtLf8F5J5FzCuLuIFdtmYl
AUE67V/uWhHTthetCySLjlsi2vEmsgyWCCAlQJPtP1JvHW9fmBqMY0vZX5uEu0gw
XOYeYKjyob3zU/sJqQHF7TRLctZFLX9neCHi31MFaFOgtoLXGukELPw5RL6xmgsn
DnGutZxdvSsUCbu4sEh2WUmYPxNhwk8YOncycJCME6OOoM713f8KGfGiBDjQULXU
RJazzqIwV7zF0aC0rghi67Rwik679/syreSI1KULYJIvWhBPpKGaKwPixJahNSl1
C6oLwHyrOOvvsJiU+dUvg0CmvJC5IYnu9zr69K97Yar7A6t/kyhmlSNmlkHSa4xA
6X+J7jxj0A544O4BA7L9Em17KqkR4TigVdcUjUyTwd8R4ZQQICy1o4IeW0C8DA9h
eaS1KRCeGMFvDEPpniqbmKuDflwu/WbJL3412z5x8lWx6wUFbwlFu76SDeY/ki/c
L6XTIqpTIYRoG3YkBStNF8G/a9tV7qLYHA3uAsgI6eCKnUKVEjdg21ySTtc8pje7
O+pcudDI0c44l5X7NBuGJlOhXgRm/HKvnaaWySmg7XcL2wbkY7FyV0ngQV+O8OIX
vVTxMVnmxKnSMFZl2V2C/4d+dDdK19yYpBe6xDjgB0VzfDSSBsiD43wS1aCir/ri
W8yisl0wGfKttYOgx8uuyRT+XNvAXWq42Fx+MHIYb6sEI2Gjz4aDyaj4VnSL2+Yr
TVT7nRoj/Zy9u64EIFXS7M0QaUKlZCcLQJ7S+y9U96+MrjLccJAVJGiFEt9a8ySi
EhVx1bnqkt9O2e+ehyghVxNNyi4gNYieYxmueV8w7Axe3LjUJnaYpB1C8iy/jKHx
DeBQjYIaX9KskGkvKBT99DRVSWq9i1FUmg8uy4ZBk9rLlJBfKf+PLFLwphobXUoq
ORolUCEU6ATEbtq1eROMVXfSVAhKjMWFKuL2DV8E283CafN+eiRMiz+YOBARqWnB
HbtpPih2dcc5TOPy+z1kxs1MtTwirBV4+bYv7HBaKjqwWHlMbERyFu7ozivrEYiz
fENu3IGwTXjWgE65RMU1SjPoHgAJoWpVSyGK+3Bt88cgdjimAc8Cd7eX1MZaOxxg
HCkLVpqok2luDrBd33g5qquS4x0VKGYVTCvKaJ1Sk9kh8gto1kwrl43XmifYCHRj
woYlKCyoC0ETsey1B9TOMLe4/emVsoUUcRgQ7zR1qxJN02PezvDyGiwMsIlscymd
pSwHk8Ah3ZORQqQ92fkUehTLI3SigIFK58iSqvnwuCH0GR6SqpbsZTG6uBkq3Ybj
KKuMwm+3MwD/AKefnPiJMv6EW2HpGGaEQJIOkrZuUvm8Qetc3h7MWaFaPTMhaXPF
4o6AGz+NrFQ5+5wqFxvsufhsIKz5/QVbOjFEIYafGYChmi4Lah7JDWzP3QQ2+nuP
KM+U6RSowxnMf9OTSx2JEIrEV+rTXKpE0Hg0wpgr6WA13NH8S/8F4iInk9wvC6Gd
xHO31nIWIIWuMk0wvZCNySN+9Eu7buN1Q1FXLx1y5GKGkvpI0Okrif6ewoKc0M/g
0rEpYtDeKIrHBdE2SclPPGMoPM83YZA+eGHky6sqqoMoZJa3KgEfh+TIiqSSlQrI
3dEPpr1Y1o4+zXKDIxS461BgqmRuOiIhVAgiGHe+PoTSnziZ4aBC+7Gr0F0WXpyo
TwoZf7THqnJ5NRFycAoCIkfvk5JTlZdXT6qI4JIgzA21IxtARDRYPUPc0PHMR103
iX0uBoZ84Qc8+VlP08hluFpnBZ2kAZ2uuEqijseZGP9u8o0aW0jlSJnNfQTyCdY3
PbZzts6ixE2FSYnjZjU3gJJ4aRpkw0malt1zSdPmgMKFUg1cUBG0m9aJNUWtrxq0
brRDL0x3fydN5HC9RY11KK5aYaM0WoX87FN4neiA9hrQXK8gSo1KURUyZjMAyPWd
t/AtnobVlpOstNbz0gxsft/9WEaRlUlXvuS7UtuMzdmYxtUEcWPDuGMVrM0uyu7a
dm7+yOm8rcenz/QOC7/jNPgNqRUskyJHhb/xjwGw5oxfYN20t1uzeYvs0GIpJ2/c
ELpdlYBKa+fwW8tp7MO+cNWcRkf2716t+lfeo6AJ2MJl5Fdzgo3RCEb8PdppHmH0
baL2RWWfuwjkZKvZvEOc8bHfr4knuQ38ymopElmI7Cqa02P7DU+gutzs9q3BmToq
uPJrTj57iSCPilUEQXRd2W55aw1TwRq1KhcfvAvqwiQ8Zv5QMzW0OtI2xjKX/cd9
4rDkcMY0/X6Ei+3m8zuHFm0AxODukuZ4OtZELxCdMNGWBxzDQEtxuFXvuCKbhIFC
LZGPijQoJgUcH6ZglaekGJnlikcP+8fchpMK4P5367SrmTQ9aKUFBzfN58zC/KE+
dqZyxSovd5PAvP0hWvvBiw6Dzct9kc6ai3XOBHMIN5Mmk1VuWdMh4hIxvIm8GK9C
7qZ/aHgDbs0zj4xjoS/9SPytq203PTQr+/woiVBBB1cM73HK3o3+sKeiwURMDULa
Jz+tEKn7Xszzps/GWnemFXSiCeQpLTVOPsudpMZOzOPjefrhf3+at9EpsK0nNGr2
IZPewABN/Wbo8U/340RU4MhAGYBPuCFyP5fjrVCJhV0Dyr1AHH1d/k9j8UVYT73j
yOppHWmzGyPOQCtZAA5CZZ9wY/ihNX/K2X8RYv2RIhahZBijGXcju7o+QhS5xXfo
fV2Wsivh/rdbmirhi6ovlCXKBxtlcs5EISpsLAVtJLiShNrMjMBEsGIPXajlwa5r
u4OXQoCSZv/D9IfNoQ8ZSJ3INiJw4iaB5RljP1ph1x8psWlPVTEr+rOZWOA/tw6P
7ukikFGbzz8P1abb812Nur3BXw+yegNbtEguYyxb8+tsHkIBJ04s2NpJ7IkCxA5j
wonPS6ErE/CQo4u1L2ruLBRktble5ZNy34KorRcp65PJPKFQtXrYIjaYjthZFrw3
AdGiNu+xtEReaPY68rx+4/UdBwScjhZLr6cknLUwgx6+6RLjDxOErP+ILPm6oyGa
RZ9ldgfqbpfN5fo2EJHj+8Ms2+dKFYR7JDNX3PEKyvjlABm011wz/f5rQU26hKmr
UX1mZiBYYsBhB8lLOPtoal68Awhvsic5x9G9CEP8LcD3QGwDUHKUE3rv9vrIKZdG
TOIMQKlJ3ks8bq5aJG6eOBnbk8qxoiMCY+Ekhlrb22sov/wY800uSe0NMhciKfnM
9EAeNzDi6n7etLbwtm4dnHCo9/vxrxXiMKEAjLfqz3BqyQz2/y/UgtHNTXNnA+54
e5PH0e9cNdbwb3DEnQypiCcr+ERYTckZESMw7y/Ir/03Fw8oYi2s7DgDcYPUNXJt
IEeMEmICRCJ//t5hH4npUn3Xu0ruPt7fi8+RrQcIffwXC48OZVbY2BaztV2cgBpY
gNbLGrIu0VvZtw37JPPo0RJwFDb+CizAB2+OcB2EdCWPIrwd8bLOf+7fZ0+4hNaV
JSGy76UoHA6zO2ToaPjKxPPKNtv1U9kN53Sszro9KY8DzmZMGnEs4rRuIvoe/uEO
+FzPDyhjEI3LKCjR/jOgU8XhcikXBndS9MtaNd86XaS9F0uT0vnfipL6VHOirA6S
IIXFWoqtVaB/qTEfemSa1xYMV4GCc3BqN8GBOI2df1e1jMWY817YmT7ab7Gge/Di
tUyfkH2smFG+hheAt0zE++/vihhANjG8ncjeKGP6FdyfHO83gbPW/9xCmDYUxySX
Frl9FffIJOGixUfCntElM3TYUTPGf35TqHugvuiFx5tpyHVMG2teAaY7MzHhLh5d
SfW3hxat1Xgrt6ZAJFKItZBCsIJ86WKRYno6FYyXQBVrPThNsEJ3DxMDeBh6GKRP
3rikfVjL0FLna2Yy004py+HebCAOQjrmvR6GCpdyBvj1RDr/9Cq+JZjB9mg9DRBd
oWWQyLt+KFWciv9ruW8uqWb9KeQcAxc0QJPwufoVUaRKPUf/VLbVCJGLakv/Q60p
Gtj+E4hpWnWdBXXhKJo5FnRV4Y15wMe9ohh13JVuaXdO5MOjzlMzJeREJFITLhHN
Ly/8We24No2taAXBtTtuqOmP8zq26qMDyIGHzNIEtbYFR65TLKy0DKkbTrKu0VDd
K3D9xo6oL71SsAoeCMvRnpEioHJ/GLwHrVhlWQSwJTIj9wZdAd2iNP4Ge0mwwTwe
oXTxshcC1dO7KqY1s9NNQat864usQTkzcU27L1NyfI96i0ddfHor9T1hz/U8KKC7
cTWuc4GZntUrwh+CTRamTBwevCKQhGgXZgc/UCDj71g7QHlflQSBXG1/V0lF/CcX
FjGQyhCljlJX0aN06pv8syveQ5YO6r9BVNhZBhGGCebOWwM6zMLF5pvk33VOocju
6AHUUFVw6YJluxMwbh5/OoYvGF4vUmitANTvR8JU/00+eNrM92onjjytBz9A/iMZ
R9oPFmbvyhP0X+PoVfv7cQ1qtyDgeA+uUBbehsfWgNcR7zWOyKQj/2Mi2uSg7AeP
H9JPE7hQiuBBB0aFRrEAHOAHknefiWdLo2Z8/36Zi/PkMWZb2t+uxA3TDOcmSCpm
VBxgkkrI3yW/0lRQnH5aS7TsPuaLLP49ZMlSB1LAOshYUDFF3moLeLxvl/5hiY6u
5TkXSJk1RBcvhUx4j3ERYEZTM7B0ecrJOSW0NijjE174KFKLeKT9MpZ/OD3NzxDa
KVlh7xuHsPWdqnsIoHNlCaxnfxrJEbyYK9RrdkkKXQrMWKUN1Y66BfPakpROPPLf
QvBHQWOJhTwo495nkf1nLugReTRn3tdpn+1t8j4Jg1svJcLOhvSmdQ0yrkkF4Z+5
NnMnSWJALMrV/AvYNcRm8n74lFWYVdmpZigyvOsjakZkGIO4zffop+IOMHCqUWvD
4iccOzZ4A9xC5v/bDn1BESUJnIQP5UuN/bVKhJuXUdBYv4g0ZuasGF/ECxQy4NkW
vh6eIJKhm4Z+sbsTsO3OKGgKorswqVJbM9Sy9sELp9cCsNpiPl0XUi6LJqi/O/VL
e21GjJ92pC7hMfP/qC1xybMnOx21SBlX3JjXXJKYGKtV3i2W4g9GuHmno+Czvwe6
l0VgvDA7oKxb8T8uEFIconp73Nz6YXI2DAYk39crGunVQOoEJq8xUgDwiDju0wqC
KpetkOdxu0dmm3eYF9K0dnkWYYPXprkjTYGr9cJuCanitKuwzJAPqtqupQsrzLKn
OOEyanaqgb3dqwBuqzuYO3QfwrXzh9TJvErjMLHX8Fq1joI4rxe16vuLvXRE3QjT
pQHMlvIzrVVkVRgMte/ksyVSQnpV/gFm4qprZTgWTJJJzM+L81vOcBAnz7gf/oOG
gXWsEnEal/0fpDSvQBQCvQwkXCug76VgnPfGWW9aklZGWwSPRMU9oc0iVVLcacyZ
CeVTD8rZC0POo2amaawAPZlqduujIjbzrZ0PqmScBHNhRXFlAPw8ecXSVwOL4sEf
c2YvabY8lHo4PjlWurcKAFn6CV1iPCEFyA4F0vYmnHNfqX+XfFXNi0p1dZ4Yw6KH
6p8CAqbfCp3zTtbomEh/dyUkjIObIQ5SgsrRNejEob5XbgiEwDDpRj3KJJvEq6DN
aJhsF4HPi5XcQftJrMmGUvkzInSJNjhs9f+EmwI6uwEuTu1K20mGxKezDESBo6HK
YyV+ubJ5UVYYhzyv3D8wAUbY8PSDw9fUlfXIF6UAv3jgprjkzwiym893FqBGagxo
zOYGl4umKM4Kq/+cYlPwxYS6JnvAQ04FBQrlh4rxFajbDxZHQMwSiKAxufQMbsht
qdaoYHxwpfg7tRNKTr5mxT0K1aFhzdbeQN7nUHEoWWzbr0Vb83btYVgwAT1irgEO
/eWiy+0ci8fWjFniwqj+3ZTm+PwClm+e4ZvzZyRsVSFYkZfPKgWY/KA0jWoqVErZ
3sLmoCTzYymEbWLPAJXTa0kWQRUJWTEoPjl98aeErBh631jArdai+9Ts8P7pbiG4
XjeSzcmqTNadHqOr7iz11MIOnVc476zofGWeb4uIJsZUHaFCzlLvVoaHhvBtzYib
OH+CBZnn4BHTY2ICMiDUC5/JHtyzYwz3A6o9jkepkD7dZbnNilckZZ39yj229fMJ
77e0zbcJnD0/56mxxd0jtzBB3+t0UHUayHuq5eZBoqvtMpiWgdzkrC12IyIDEofW
s7wR9ryJqFVepJ0sm0N3m6udV0y0gPYin+R4BcV2bh9RTbXHLioAKf5wEdbKnu52
+9koG5GfHXeP1jecIMC7FL+cE2C1ywXQdBNPlRvbME9uCYatbbAMQsqTtWcQP46L
emS7UCsyGYUc1SExL3RThfx3wKOaZgI8KELjmASNnFHiyI1nj0aJc4kHWShqSbT9
94/KWxb1L4M0KZ4BG9iY9U6/BPEvHRQV9OilM0hBPUpjIMpfVVBBiw2u7jFbKDCV
SjhOeV0kEcAGzHZu1FYZxzia2m3/GeB7drVk4F/tjfzwsbCPdNSP+hXa5WNVdd16
XvZS5HOM7GpRMI8bUoVUO4CIOOwJphgYpO/Wsb/HunXOt2TDIoSHLaxBBIWc2GuJ
9Qlz0uDaXDoJuLqhPjHGQ3JchnviSX3pDvkpaGqzPmlldP4H1HRSiZnvRaPxwnTH
529ZcQ+7i8QGdIoDZADgX5ZbrnelsZx05T6w1+IZYEfoe7pR/NljZ7cI9ql1tTpH
qTzsuTBhLKOj8Hl7ydNNK/B2DieMD8EHeyjczrWLt5dRWsAWjR8LCm2ZpQ39QYeJ
k5Mc+vfCbTb6p7L2U0zDdf4h842NwobFUe62Lu3PxiY/P6kWJ4VG215YDLDVcIzu
Ba6OMsVWnFPmpNL+2RplN8TSJYZoR9Fy5tDt4VaFtLZrbQrWwg4TW7bPNPWW3A+S
86QnTRZ16e91Lz/zZU85pWAJ8SMr0dXHDnn8HWdH98/ZYjZu8rxgaIA0nmY8PIPI
Al2XOjep4NTlU6HZ5wfseKpGog4NPitu+1lzIfn3jQypY6YF0f/THwNM3bQhNpPI
A3zlGUhfjUb21d1AieSWRLOIefjTUI7833vZ9G/3rPsBzkT3kOYe+MlJfi6J9SRn
5UCTKVfIF5f4qsR6Mn6cVjC6qydhHo9ljdPqHa7sTTqqedEG9GKVRmhhb3ORq7Va
v1OJYAAr8omp6GbhR2K+HqoiuAXiKwChNfYksKEAvGLoHFiRVrOLODvEAEqq3APM
kAmYKwMZHAoGo9h4Wi2uCI8Ly/v7gg8BB0MqlYFzEUWgY50Xgu13kS0x8LeBDdMQ
5uM7G3wV09Sw4RoTQoJt8umTnlIxFCSxzUHqy7uaQfHA+LDCsJnvHwCe2R83q2O0
E/Q40oDyR64W7haMHHPudCFaxL3OnafD2x7RL0QqPfcEIIWT6M+6VMESb5bz1uQq
0QiCgNt7+rnbiyIafj4QIM20wuMvyjbTSC+LL51KGTYbwxLR+/cLG9YM/f4gOsKU
El1uKKtK3FCXWpZ8elt/WZ1qAcoUmL2GaTds38nef7NsOT2rWQjzT+OvNsIZyv2N
6DT03qhePstY+6ZdBKKKEbMqWZHzUdXY+1qdMeUiIc+cDlYiUCbBbsLmid4wA8Ih
WHNgEAdhHlBB2/Gz8ljK0EfOd6M552Qgpa/F7hB4Wj1ADcXUwM0fti0xp+XlAknm
9GwyL5dqy9L9OadQmwyw4pJaN+PLl8nnYpda0mehT5IVfospbJf2yMCeFs22o/hY
tWM5dr9LJsiSOHV/lQqPp8UDueo/vvvqEjP/t6vvbr+xJKAQvRFWEr7zY5JFU7NQ
rGBkz2rFCCByIgCvK6oomb1qDKu0UOPJ/HjORvpsbZEh0WtgDVBSGLlZ5BqvemGo
IDfSHOlAM3exgdq0/2CiTqb+a72mG7cYDbmdB2eKFmAUfUnABVS49pZhP6wZdYC5
nnZ+CUxXPSw+wV37zfS99wN3zS26LbCuxCLqiKKVOeAS+Yfm/iBQjjGiWWHrOOfZ
XC1DvXZueZIAmbZHoKm+djtdIABxH1L7vprpZtbYAGJbSrh6lQEq5mmQQT7sbrPo
6Xm10lnRQamfCD0zA5/t+NUdtykiGkuETf5oKcix1HixmGc+ehAT7j+hcvJVnMiL
MJ82p4XnrlRvghRSTWpjTrHNHj2aoNu9BvNGzB24P52qR1BYWVJevwJsMGrJEmPv
+Yc3wqTN1UVl+nog+sis2vziPc0yvjhPHNmFUESYeqE1Q36TTrKuDOC+oy5pqFm0
3InR8f9jAElL54ZMgSGgg2Ap2ttptKcHnLwuww0eRxoPvvKAM5oOUoEWy5Qyfvnd
JPLictHqR8wUP9ESyC42zSFcKbBhudX8594poXgMvy+lzICKWNDIWcFIfZKAqIfz
HGw791jYiKwZAR4SOKYiQkVKlIOf5RGbvSwvnviSagJl3azyW9ZtQ6grA+owmzDc
KLDFqG5RA2HlrHkmLLRhg/rxRlaQNFm2YBwL+JWzvVryfvQK1sTQ6iX85jnpbFga
B7xzsEu1Zq7D8ipyeBKqCnZRWX2ursM4mjKoyXHBnPxVBaqhzVNSnF42CcXdkN/a
WKRy6q1x1IKmlw8vundlwT5MFQevc8ZqLVM6/Z3+bFsAKxgKuDZ3+oOH58OfCoUz
Cv9WK+WXdqo5TMAS4fwD4T4U3NGFJE5JjOMzKuQ5rMVr0fyR56r5LsD306Mtlgxb
ODWQFr9hvfwtqkKOz7NSp6u/78jyOegFUOMsisx7MKY9FAEVVOGZcu2s3zz60/yi
T4eFciDfEwFiLUx0AWVdKq+f+jT0e710cmM1M7tlHWvuJQNckFA4bn2GZhJvp/Ao
GRZUD/Q+hxbNlqIIO2klyKOJY97rl92zA/Z5ppES20M6Y1DtAktQvlfXYOMQWPpx
M58tCyua+3nO/FcQ5ZsnJywKSsSHLsUtkL9E2nhqvbYMxtt0NZ/mileJpyZLM95Q
vdIhZL+edzxFtH4yE5GoYMoOwLZjt7lqAwhl+dJ0Zy7x0tZKPSpqQrGtBXoZ/Cf/
E4FPiE9xG2Krm5hvd16H2DBHbvrzDcHx/R8DVzbgB2jOFYjHg6pAV03NlSJ6QKLn
tLeHIqX2IACriUi8tE3HSSi6XbZsihDPJZJ8xeoPM+otgtBFs9qBdh11gnzRjfVK
mB995D5JjSKwxqerouE1jlPPr7WLfn4O9gfOk4u+RVR8Hgl9igKrc0ROvQuikOmf
ONkjLNapXZ4pCxlQrHG+1cRseWSyR10ipnch+C7PHsps9pM7v2zoavUHIwUT3uKi
C9z6w2GJdVEBaeXXM5cnFnVYh5C291fVlQAZc/mp+8COwkWwDk5WSiFCAbQMv02J
KTNkCRZVaStsSTF8ruJfDII4zspM1nohbD0tj+HWZT2BAGuHdEyyVzwLqNeGlgPN
mcuCM7JgL3yP3Oj6BcfXw9fjFQvZIxrJtEpfoSMBvkCpijG6N3vFQa66XgEkmamS
1Rs8Y6HALfjmS4tICR/BBwjg13DLFXkcgOhWLSX14YIBYxUKuLbUV2R+zCVX/9J8
xhfBXjbEqnQ4ROVDNjmHwYSp41iA49znOQZ1G29W0wrb0ODRet3AppiRntTRrckH
anm15d7vKEBw5/fsIYOnt2FYpE2DKU64pdnBK+m1CpCgdab0abe2cmyuR04eldEL
L9oDm0tzYzfmI7WeCeb6LrEnEgr7hspNA4HJOMBpIUutBky37+SmklDsr+pZsQyu
EGnGvpQjvnJTPXNV6Cw77b24X7M/LWYOst94cn3QYz3xpzAWoqy/VYZvbPS2lYUL
yUBnd8LJoA4x/4dHn6hhR0fIXx+JT1NJSDuPFORXM1JYwRh5w3sVuxUIbg9oCM3D
7cxvA2Zprme6w75/A/Wdt9IX1jYMoWfNGkeMBNLshwal4LNNFLOTHNMYZrvqPyD5
Ufqy2Laml90XzhYH3tcZYgSzEmwgt3sGZg9Tvg5B1Tw9jZMdVyxPevctjtrUqotb
cOG4xHxVQwz7+UIU5BxtIQUrT2GWE0KlJQRfMVPpsWCbgiY+P8VAOVVYGplgcU0V
kLxEddtn2TfhLD1ffd+0CNJ113jDBrxb88LO8d2TR98l83UJdQqjbnV3flaLhp+K
I6InNZxYJ4Fwc1UZqbiAQwSLMmaXHI72qn+S2f6kUGRMpaTdd9YCsZiQTg9s1/Ln
KR5YHnm6qqL96iUxIkBQ6tBUJtqH8d5XHHCq9/lszbO2St5HNdFIch8JUoyg/7kT
TPnbxGdAmAnnscUSqY+y9mKL0smUb9hBgyocIuNXZ8kFYUzaP9FG5EbeVNC9RsV2
YQTVU8Oh6NsP/TuiKw9zaW6dZu2SR+mFjOPZsSDvJ+pYNjV1BrU42WNjVGVO4qXb
z2Xw7W0iIYMSckWuCDuWLUbOfR74zFRSl0Xys6nZn29y0wR0HMEERkjQ1s3UtuqN
20ZZxdlQtSexb13wo8ouH/c7J6H4xY++5C7WfzCIaHLq99USUIyKHvfbmWJPafao
atiAruZWgc+uly/JB1MSeVYl4G2szGxBM2M4AIk3bwHlV8bQLJiJPiR6JDieSLeD
WFYOOWob66GmPA6nulZXypLV796Uw0LuuOIIqcHkhwa9HpZOWxq6OhqZwgYE4bcw
y4X2lUFgnILA9YxzXuJRYj43TZ7mKf02QjfbMv1V9jSb9Yowo3AibNmRwbmw3QWq
8E3QqcjMkKB6gCiX5RRHbQK4SXNB2dMGquZveBCAKMzpe9FAaDXFPLoKkVpbleq9
oJ14euAZwcKJ3ncPp0Caa7wWqFEx5NYNlpJEudQGbU0mwu7WcL9T/rmuZmUxSb1b
KNSzfl3/pdupfL+vvKsdcOL1i8XwdIFjf/aPnkxljqOr9nt2GYJMGVInGGhNfNEM
6m8dShFh+yep2/7wb02mX08hEZsrf/5IsWDPy3a41WafH8kYwJonROrFMbLZ4o5V
0ky1MXjGgGrbqKydDiiHWHmMtTDaZfvmL9TJordMxsz6IaRJlbqhlvnUWvbTjblq
U2CeaXelAkNPrgJJYc9CeRPnD9H5Ft/GFx0y9tDbDFwkNI4At1NhkkEOZxRe7uj2
+t/UL2hQ3oNMoX5c2dopptM8ckEHDzJ0YiZ4m9UHevoTKjsuW7ijNxMrRVXXCi08
yBwqr5meSqvnsJzERluVrQJFShZ1HN428HRFvJG9YLVvs8s5MT1SSF3n2GoFOkhS
QD3OGaRhNVXADxmP6hXiaexop2lhWGUDrtLBSR7HgJVi457i1UtMgxKvfDMXBXHz
JjzUiaUNNFsNGLJBDUQLzHn4grVxdAalEez+sNamHrDoMcPxNi26ps6jgcyChokd
PbicLtd5B7h8xdxsXlkJ11V4YvPkyE12pYj4uF1nZbED8JfiFVmt5pJ+axw05nF2
MDyPkiwSXB+//khKMpMBO/CnXUBsxQ7relreZtl5lBXYGVYY+eQ1nFfii7Z/t3rb
PNsE6X1zGxq4gXaKin+gH2CMG4okknyDf4z6Aoq9arGTRwalSa7yNtpS5wD3DeIY
UwfoObFH1jaiL63EIq9ic1uz5N3VHd4K1c7sspfFlX9a+PFPbiplbhK1Ht3RUa8W
VN/apWZ0u1VuswlPqaGYCgOe1ITgtIGhLd7qL6uvKx2l0u1jqAxDeVncdYZXRCIN
Bu+vw0lSDg3Hgm7MUA1z+RLK+gfV16r9pmUFW4y65+MKXwZnaMkht8hAKZn3IEmj
gUPHt3VRMypWXbN+bqyT/mUhtD2vx0r8jkueeAAjD/L2MDiww490pWAHUcw3QYYY
7WYOgH+//asaj3Mlz0FiKjROwJzAgs4mXkySVZbeDUpDrMsF9qReSV3GF7YAFdWP
9R38S0msssYy9XoVuZP8bkk6c8Ue2wBFmfeChEeuLsJaBgbHWfHpHjpD2m2VVUJI
H+t1ePD4gwwzE5ZoZXYTLgTXQzPM3SFriouflTyM7UkgcZX1I8r11VYi50qaCIae
oBL5fDcEYl/Zhh0qa3n/tyhH79fIMJ3xyqPwRpnlICYkSBodp9SmYYASXu4l7K1j
1Lrkt1u0rayOlAKVRdQG72+lPoSrcMytd93Ja7Ku+pIkGnF6W34Gur59LoGZJfEM
FYPU21aK+qKznOC5XrZyyxmjkL0ZTx7BFntqWfiM1VBadxjxHqwl31Bc3AcRC+K0
isB0cGmU8HNmb6IXlOj9P2rLwDxe2zZgygnbgPLsOZyW9qMQy6vciolaE80KgMAv
LJPVVdMslhroiWoOqeJzyThfG84QEzMs5v970YyHVUFByl2poynfixBsTlKGF/Dv
JFaHQta5waYXCsn0E83F6zJ5CmgRdKgVz5YnhNfye6NTHeunVSF+sP5rZxRDpjqs
5ygczQqBgq/CczsOssnd2iJQxnzbs8Y60ooE1fmu6r8a2rplQsMoU1zlzHk+2Gia
d2dBiw1V/s/l06m7cI7kg9FdnMANRbRcWgCKT2RDwfUjliJodeEfPjc/pvDorK6Q
R+dVli7jB60nGkkGHkb0dAJzG9pkeUK0TMPFAiFeHTznk3tsht7s0Gvdc20mjzmV
ukQW5YJYN3928nwe7HX5JpQSoeWFId9Rq46wglhpf1HUdA8KznxjHbsJ7HCYNPKt
MQbFE6Ihq/Gi4RdGXOXj6g+xyok8nhNv1RXbElkSwlCDBZRSDVvCatLW6hbkV+3J
W835LCfMigtYHEvtEvKHWS8ExkCRDLQ526JcC+ueCBfpH2NoqIzU6tBxpLk4S97i
hoEl5cZ6YR4j0B2Ercmz7UXQgSHy1MTaPXxAjnRsWDWq6AMgIVyoBrv9KNpEBNAD
O89K//Q46fN2e66iDyKufDpARa9lBO+wGsa8XFmL5dnjl0i3bRRl6v6jDNKmCZym
gGb1hs0rv/JhhOnxxj6WzQaBOnQgpjsmMt3gI9BR7rTGT9p5WxoZMhmRlIInsuvo
zkLH8Ul7A9j8CgSXqYUe5fvsIkSZG7GXort+3i3+M52PejUPYE3da7HnNcqpQxXy
lXhA2Zi74qHh3YgFojkMG62UEsgjyk4uw8kCCGySPykl5W9r7j0xoOi9TzfrJbz3
X2k5sTbZMQGAAOv4fw3HCOHFBPUfFBGUOf4aQWS1zqalXCZHs/GlXaTb31gG2FAV
XHmit2hzodiqTnz3JQsZs3WAkI+ZL0YqPXstgkFvyoVqmJ5qYODcfLEwcYRls+q/
PJlVCooUSddWqNwPzyOt9DpEvSv4dXiDkzN+xHQNlaGpQxajr/7VR9IRTZYDspfC
Z7oGwJECKRuAi1M3kCC1+iqEkIKhL44LDsPg3kuRGP2nnPTa0dTJTCcwBZhtpmgE
/SD8JdA6m9G8lV9l+/5E3E9xNMJk7n5jHbJ64sfDaEDBU0S51EqesC3IfRxBo4FW
Nprr1XyJ8TLkpRX4CyC5bQkj2Pbd/7z+UY5IdyyJxQeqYI0eAfIEsOme8Yo6K5t1
mGk0yA3TQjiNT1KRNWREIDlD2sgAX/j8Rm0h9vGaXoeNsmNnCcibZc2eVLQk4R0H
u0hBFMNTwr2PIdjsU4v1OFuW2B72tbOMApPlxJWtBH1AqHS9LzOahAE8xChLVOvY
DbAu9X+zb0Jy0XBzhbUB58Xkrt/BFW8vKnOdTbPKupZNp01i7Mx48rC1yxNAHbca
g/ruprx2z3KzAAIEDCQX2WMknGVt5watTURXHEsCVRXWkvBYi79yEFPbZzNJOVR2
OjdR+rBUTnF8anugd3f++y5oUKhje65ivK1PGQM3jfNSd27FCphpz2hcst146QQr
P5p/rX22nHbvhSbOT8L+N4oB6/PdZwjS5kIcIfXMgUU6w8AoAlhL2kAH65tt0NjO
qvKACoOQRYzuTflXYundtb0SkqJaDRSfQrIMt69Xkmh1J2SFAeMoVBOYYEKpk3bd
h2OleqdRanlxmXlv4P+XH6Wd/flGNZ+4sWGedOMsChanHUrP4iTefB9qEZaE5fm0
wh5/FTE3XcIqFoGDvZ3QzISShxDK+tOS7R6luRxsRMGCCL2PniLX4ZVqvpFyYK4Z
BpUZcGEg9/o/SLZ6Z8rReD/pw08PXw53DlguSqnQJqFtz1U4bbR4MhyJ8u4f51/X
rQulTcLXqFhCbvnjVq7+rWrSMDh4ELcawm3lXLacT4YEeEWNJAlH4jwB2jOA/1yc
lttmbBhNOyeK0VfQEmRBD9rTMirWvVeQqv2QUv1jzGjpwwwH4JtmFm037aIGNn5R
xTBPGzQrGv0CqjhInLmm5qEjUTcJJI/vNNIXK/FxG9COg70gDAGprRyB6G8AxpSk
Q6n2XvzN73wiFQhDQdj/ehjurV5KgleR+WPENzdD94qUqpbLvmvApcOmi8cB8a41
PtadUS4kjBI5ZG8rsMQIZfM75nklNRzjXAcoz0a4oW0DEHCw5ohqKMcpyqnT9vmo
khH4wp3O83UdKXeewG8PyXHUQVnPGChzMvjrA9amThknskAb0tL0bhdcGUYPWRDP
hIkcxoGhCbiSrxennQ8gwddbZX1RRyj1WhDCrDSVvlEs7sDDUp3dIt9P953poVnq
bzOMy2CbtTMqOfuhckmSHIIcjCFcj7orYDKH7veO8hr3FFGdiL2Kv3SBfsmxyUoj
pnnxKfjcZU0ZAxV+3gi77hI2wnqOESzx5WQeofjUw4IEQYa/i8TmiXRofRvoTqCB
ce76asfPF6PGRDWvzgPRxGnwUf0pfIJP1xVs3NHBdwquuY2DG/BNDL5sOfkTSeVU
NlHuoi5Lq5pwy6wtcnhfpCEutvxqKI60slEAYiwi6BeiXO93O+mdVd9K5CfhT3ND
Eb7i2x9xshpPxSLDlQ/fmuzLIE28zDrqlvv4oUEVDRqCYw7TgHyN/yx35danf5Yr
uuTyighkVHD0tvouw6aTAHlLNilnmqRHmtFWDd+uf7RQHPCeK0IPxGqtZundo7fp
l5gtm6SIqajy1MSGB2LzfvPtdFaXJm+g9p/FYCxSKcWU7jft4fuvr+IOu9NOXhiv
tpVkfFPC2G1aerLemVdTp3B6vKIJt4pA3RedrYr/vaFVcXxajY5yvikRKqQ8MxEO
B0NGxmVRuQWTpmDpOxbuI81y2BjA4cMrLAorSH0StASydzYRIcy5+u+NVT/ophVt
KxIAvtpGLUq7BkMTRheZjAshBwYS9AaazOdpOsYWKOCsZp6D4ugr9V5Hf8hZCqCD
xJnXF87dCRgp6SDxxjlXHXIHGi/7Qafg2EK6fLA5m/ASwuFnnVA02oSmEIcoOQVp
38HoQN1aICFpeqfYtO35wxOx2r4mFottP6aIz4/YIjzRVHQOq8JKlYfWi9zbUEOT
cg8l4Pgf71bHAwExds+oZgIi+3FRU6v0nuw5LcalzKS9l3cxc5OvkyZAfWWUNv/g
0EoMiyhbSq5KeXuaH7KYoI/3I0tE1vTC9buEQWaaWcwWokeHag4W1178xPGJRbBU
9kWNhLrsjar40uRldKRIRBHAkHUbhpmWvHLdn3tosMiCndBaJKHCja5W5XRueU03
O/srpchJ82DAXZHZUayddlJ3NYUq6u0+clpeVhwdn4n+aZH1BfiOaBPf6UQ9HfyZ
Unj28PsiTlhmD/5Zb77MhL5FAQ+nTYnGr3gi9UBYYXPUWY58wyqS6XqIJCeT6yzc
cIqsrKJA//e33bNbDi7M2ezdcI+ibzDM8DbMNqvQhblO8OoPitGAmveEj7Z/LTNC
dQigrtw3IaegA0Yu+exP5/MiojP/0vQpgMyr1O9kyTTRsXTcc0ZoRGH9DPh36uNE
ss4lSxvw8cH6jOymm8EW2wR4AualCJYoc5IPumHW4J9bzO+KGGZhJEWJJUAj0KJA
kpx4+E06zP7/WO9oyZDJM3J+za9Sv+M/vEZ5pep+cfDM4vljQAM6krJNkiuSrxd9
TgPad44gJi/FGpSU9SiKY6ZxJ4qej21wmzDSi8HCzRGv//8bZ+0Zxa0du+jWeBSY
VjbHa/RJlR/Znjd/HhvG6HzuIgcDcTLxNXcz++2DPE774Y83RI+s2Wf5Cu2mEfLZ
ouxnUcLFOoRzFb48XTt+0BM7RZM2L2873rJZSjZIobYI/lQU6o+6/P/GoiCprY1b
POnXSZhWi/LP/67RCk+YrantsCX3GU2xeFaPRmvBm/NqqTcfkxuo/0htv2BAraUu
Vw2Oj+FYsCQfTmpX4d4CkH0OSewx0vvqQwpS8Yt3eIVQW9UJhgRKszftMDZ1w20z
asQO3sE0LW1R9HEYK1hXxTkctJVWZHCLdkwM5xcs0Zq4Mt7XZcApL2XJh8mHRzTL
W6lejJGZ9LjoS3NHtZN0uPxYH6WqSfheEEghRKZpDFC/xy+fJWY0oi4Iay+0atpR
5KCntIyz/7WzZ7AA1recZ+38FYzFvA8untcE/hBUm5p0sylGxvuKTp4FtSclfrhX
w46/VgtxOy0L7XN4u3QA0J8bq2NSi4oX7CFZqXLC+fqvGS0h/jvumb3AD8pKU6ob
yxirLAe018vbi2K1YqARMgyd+RqmNcn0SKofII7a3iHoSb4f+DX9E5sJeLBUJdmy
A+CeDX0WFxfOUuFHKcPqBoqUwsQglAdzVNc2B8j5JDjUWnanpoTuYsFfw38uWOAf
FXc38Z9pYcf/8zVJhLcX0vE77uQethXWeCRfPhkKr/iswaDlICduz9Bjmvx1/z42
KikOpcGzBR3EkAQLJX1K8PpBZILsnbBrCIvUri8oQd47yaL3AiazkwHBJiGZ4AHN
C9vky7IvBCmyROJEyLw7fABc7P8kYKPIkNzc48d+y2Iifwv8/NxlMxqN4lru3L9m
w+jZWVz3VpOS8Jw/eT/bohazty0vA8SrdQfYseLTrSyCVu4SBjStQ8grYlsJiawh
+ywjsJKAver899R2jY1p1WkNxQLK7BEuOp6cq+jqHZXNd936ToffPFHcUaoQd6rg
Faa53YfANsN3lg/r7/ypJuqCKFnP/BFfFqxvYZzBNSJfzLAanREUCyeGMUarDD2i
mrVqxEe/n6pTsU+WXEVTt5ulgiGce2nd61UlpOFFRSYkdc6wp/Np9CT7ZrDqCIv1
+0L1i491SZz2Ib/r0KqfthD6DWNTZLEYsTumJp4S+4QkBZPq34cRlBnWQEgIurab
TXSgkkrU+URd6xIceW9KLG7GGfHMUFqZfgxpVyHv/alRHOaEwNyNMT71YW/X5FAN
XdglqlJOnW7y6s/X30htp6aLphzia6pnBbxWXLc7ePCxZaVrAopAOa9OJSgeXGnr
oCGC7LUMIJKTgcSSLyR8cqwhc7E/8gnnZMyjv3l/CH6h0nR1FX1qA0iD7SOc3XSV
W6Yx8DZuIQDO7N3SXGa/IIp+7KFCU6yP/BREoA5JMgzingW3qScn3OmvorXRfiea
e6c/hwjrAg9mK83guA4KZNQxa/Zho58Rz7PvCSOOB45jaS5tMYOfKzK1pgeh75P7
5aqiR2IPv8umcd+6jOlFw7H2/oNQM43pHRxWGtaza/Y/B8Eqz4vFZgjEIZXcRODz
RwIba7/I2gIRPBYvy8u+v7NSMes1ijZL3YybWWA60RrENSeyPD67jAU6+zsTQ12z
hd7Ux2Q2XJMM+obeAoFux4Do5hWLeM1ZioxFFd1BtO+TdwmtzkWSEFnd+WfNHGKk
NMdBN5yQWulVjflD4Od/hQYrZwLAwioQXAXcyhBt7VPbClRTtcnTMgDvPTiKSk78
Reft3QGKfgK52z+DMH4D+35fIgyO6i1wphh076KHOIJyiwyP7G1/vK/rBZNBRS7V
7nfnWA2FDdWbsRI3Fb7oq5KXytxppihy0fsmQeDBjMUwJ/ck4fCfAUHJ83EKDa67
NRNFmLsAl8nlR/0n2lRJE4E9BmOmlPOL9gWGjM6VnJOopP29fP1++ApehOfsN1bq
dKonZpdQyKzATy6bNuGPvi5kXMPy6dgIiroDATg6APsXjFOFP8++oWjy7RCb0OOT
oaj+SO4b9DfJCssD2MQJa+M0sTy+J2C/8X+1pMxtWicavb770HKW/IAaRLnIghwl
JbJC0LdAvQII7wQFd6jyw3yJbw+Doufo98vebpZWBDETb1ZiWLx0V76goDDK2DRo
AhMW1f2Dxi5E1TpWEvPL5JLnOnWPl1j/4r/mjhGmcqUilVYghCofeVtdAu9/3W/+
m3DjK9TNPtNDChZpliuifAaYMto4f+E2s76N68th3aBoPWjWKUeFuq5vPF9WM6Yl
/Vw1dPLhD3bBQj86tSpQWxynPwuNuXdR4aJ1KPL/fS9V+xBsHPebQ16WpRtub8BX
aSLIqjikM/g1k+kutMOHSg+SXjAzrtjgkBwd+uV2WHOSWixcgatwp6EoZCy2wnPY
1H3N/3sngNHbhb9tsE6LCl9SXv6eURyamKche3hhEh5Fc2slZ0+uFzzXgjf1tEEL
wz3gqiabQSjRgqA9k8gnrJeVHxPUSt5ZRf+JYMjhsKV/OxQjS4CUDWTPPbTIlLy4
AMGQEuDtT0onf2Ci7RUY12TAmoo0294FPYBAsvxoJW8lxFAU4eSJ+4RYsCROL5Jf
dj/ekooqm99i79N9JyXuPB64FsEsPFm2MawVz+XuyxonamC99QkdeBquOlVHR44t
VYTZAhBFPXU8/oNwTUpYbbHr/1gjlPs4JXz4KcC/tiwzW0a3GodcLs4vdarN/wjg
Tlw8gNmt+QJjdSVf0xG72fZ/aNs2f44kij3YUgBw72iK2SnXmidbzBOeuRoZ2X+D
Miq262soS8BiESMTaM/5Du49L4k9h2o2uXiWKkU3iIUY7lN6paTVG1cRBB+5839z
ma2Omyb04Dyx/mEgyDdxL8YvfQ2imLR3lqmniBEvWwtp3pFC5U47ogd6IypEMGjB
43IGl1qbVDYgmF1nQl46CDRrXXCDsJvHn06iPQxAUMUwci/FXOwKODWoOCZk9q4o
A2wYF325QlhBFoYPAjwBgH+t66rs9WMJ7bpaBYz2F1oF3EMNJ1Iej4KJhK4jxbRl
WfFnK2l1fM84njw2phLpYxxerW7XREsOlPWzgIwM4DnvY3qjB8YLThzAW6xYuPaE
7xna6NuRTMmlQ0OhKljMRJLIsP/NCHBGTz+Ig1bc3SG5FxgY4pKw9m5MTBHuGP/x
ou/bC3kEbDVpDHV3LU8lq/u3zhfn1wjLM1auaa9XaJconpal0EfOxW2sA1Gm/3F1
e2G8QdIovYPMKzM44TkoFvjiFyBLwojwCIjMk+bH+TBCLmWrT43Nh6LTKLN49MCb
yjdVE5svPqLMdANzhoMFYPLxmHVvUaVAf6JUBTci4hRabolM6l0GjJaOL5TKeo9p
ibI/XcHJVZUXrpUJRBHT0i5iREh8s793NzdkVHS8FPFVJIWTLFNwGDPAUd7PVuiH
R/Jekn2py2sPaexAd8lN/DcNMoaP+BPhCxJuUC5PPmAz3bAFnKV83Ac7s+3EpVEG
IdDiXsJNQEtCw4zRa6Pbc91NYVpgPrhxSqXsc7NLRMV20gaI+vByL9g6zGDtgyqg
43HeUrfuSw6ZRF91CqN0jB8hPztLMs/A5pfaKQUae0S15EKRG4RPvLP2l5h9fX9x
AuRrQlYzCn0Tnqc9BFTGCE/fA2w2Ww0j9SoS0ojpsHzIz9cNGVU0rPEi3Oz0BJ0a
99Jt5wFxA8u5NOydqs4e+cQe3+fGdQjE3EvZ6wd52wim9M0Ify53SRIi4T4VIkNT
zrm6kA0jGvShGJUt8lTQJWUHod1mtyRCr1DIF914/bbTnaswWbmdPOZTVplYMY0/
sPk4aNxwnuRPTOGyyimjw9WuoPzga7odUI3HtXiEHr/W2D7Cdbxu0/IKbQ3zuWRV
fmc7z/kHoP/hro46qeK9hu7gMjugQRjYoPXQ174rPxFH5u7Ib27lPJnS4qrhNKMj
kfeIadOzirjP+D6WWyQK5OrL7GPD+8RIHF3fejv3JrNeIusXIf7Vkk6aezBPDx7N
XFCHxlL0xrbBzPqFzCcnF2wOEeVjPWoROj+bFX8lVTP4gv4bjnLuVCI+BU8u8/fV
Q7n5MTdmpgAdDS/mSUP5ejscPxefXUIf1f8CHN6YNGkuyiUMW3LHc6wavzuDlLf/
9pDJAvTSDXZfOXlNXbXOieH433GVSKQWRL9tHv6c1CFync/2w1hCdl+CO69lbaxG
o0iEjtr3C/qJaOhxdRpEHGT271k5UmOLJpnlkdOntuj7rSnEx/e2YbQYbeYycvxZ
UkIdmwP+aDvepYizCCOsT7bsJcdfVELQ3JB24zy/IOtfpnu5ofOrsyK0Eon7p5QM
ZVZDZ8SDtLIsN9EsH9AgXZeJB5rpGPC3OQeR3/1iBx8RU+Jr+3lWehwdnFN6mqhy
xWDMqB/OroiPllA3p3aN0wHouN3KFuPCkeEqakEGdqlnYM32U1fOA/aELaH25UTu
i1Rbk+XzWA8wXd4TE3DGftif9ypmSgmHN+yo9uAd335Xmt4K9f59vY6o6Yk4fcXD
OvrAIpxmj2jHQY35p2F0J6c+HLMzxz7udyx9BKi0qz753MhVvWdNLVtvsKbJ9t98
qSVdbqdGTBGNQmQVSi3+fn9voop2WNid9jLA/e0hZt4mw/6WKtTjqQL6Fn79GAmV
ySYGHqFClEWpVYLtTwstldF6G6kGB5GGCeKx721WAAe+Z9C6TWkY8+0epKjKzqaS
dp5N+eFcNvp1hm6zSaiis254FcqbXmBVusQsOA8jvTHcb5R0JlAk8s1WBbH+Fi1z
rdAp9FLN7tIug+tmFpjJxNRHeEsFFM4macU60Gr5rp0addIRiboGos83cSnIrbZc
In6VVxM0EXuJWcDkls+QmQGUl8gKO24ELBkpNb+tjoOkjeaq/hVwWQ6+ySkzLVJE
3secSoytvCjF5BnbKka65cRoFHscrFEvsfNWqRDYdF8IC6iIprRT/lxfqEgCHA4C
4UhvXUuTEk7kTbWhzptr/cQkjU81HGwY+zPI4izoJxwmfjHcsmtdbYmBTZm9pR7D
OP7cCSx/ik8F1uVjNmAz4kETXvCBtFxYq0jNd+6815rbaV7XEYnZ5m1NU/2EF3u5
5LFsq98QKxWPN+m9T+cRlpwFV+/kSmtcVZQA1KGLI53rtsWjRBLBQvFuRZ/3a7L5
W/yO0IJU+xsnLDT2GMerhQ4LAP2OMLlpz3k4fuR/QAzhjLXyTxtS/WfzewO0bPJy
Ch1HPd64aacTTn7/rZSMWigJdfQ2Bba9KSMYdqagQkpntoqVyvCufqt2rTnwbfd6
FuF4ZdsSSd6h/UCuzWb/8MUsnb9LrYjsgDeh/CHVL2wwGZFGu1pERoZbwMtTG4vd
GDANbc0RZiehlHWIcJMF0D0BSVedRUJd1Qglpx8hHL4RyZBJehyNOyXQZF/J3qRE
c5ZiHuIGxinAjbhfS1iFdIqe4EYuI533ZrAZpKVKBB3fW5YWP6aR7FxXHNPMPxYp
o626yD7FxQAR3ATmpa3F4+clVeUJp36l0qcyij5GbiBe7bNYWA9WtdSaDQJfU6a1
5ovxI+c2HnPa87ULVcTxJaKErSkdeSQB8iAw5c83cjVkhqtTuFlZvARMpTx6kYS5
wMEhnllCi7EQogEYsbPTl/RZGyFXgMYqKvCIWUxY3j3SSvHVgbrz3xqiBbvLHvJi
TiMjquFpG8WIEGnF6PespaaP6o25j9pIB+9SryNaTsXznUO/5m1HRe0Pys5DIfj4
x9OM5iklLMK4I9OSPNOKYBRBEHF/41ulxzwkXpbxuPtWbjzzGDL3osdLnL2xKurL
xMTI3AYeib1Id2VxI3m/5FYQB4wuwHIptbqM0ol+xZMyzY3BJk7a+efzdXxT742R
OktFFSg4SiMITrOo4L9Br8oTm6YTB4RyENY4kyBkNlOvxDFmbkmRW+sUfU5JzdfV
Opxf8KsgqSQf9IcXNqCTjKYOk6bybBKCVPK10wQ00Mmt4mJz3BE+Ld5+ljCFBYJy
yBf/jyYvG5yrR7UcSdK9zKNP6nfpI2swRzhSzG/djDteoy3eFq1ircTdZDkKvF1i
6iE181N1ftkVrh6Om7jg9N3v/hPRFC75442nymWJgiVG7RkTTQX/LmAtnOznpDTw
RVrEykKaD3cXiF28oPEF0lbM9J83zWU8Eus5VLcIY+4RM2BcVz14C62lY2AX0GuY
jjsBB+XfkpgPqFi2DMiZtoYriaa3ayAstnNjgZ0OCPHXjQclqgNlqGLkUVHCUfYs
kod2JfCJ9DW6JByZmLW4Zy6PtUOmtRBpqk4x6aiyr6kDblrjRexEqDCU8880MA17
DzUBWgSxfDXKsoU/9aTahjbFdccIiWf7BWGFvLJnIkgZPrqjUo3KTmBlOPBCZQ2Y
hzuNQi6Bp/wDjmysUMA/cD43rKJiqLONI7sjTtA6OST37ep8VAT3AYnT78pxARBL
YO0SYaDoie1v2dZpwAnpBGjRqgA2soKOl4NHKv/JVCYmr+LPcH6By+xkX8yfJOb8
LcRyg8uadotoQG3N/oEr9Sifi6V9hCkZ7rb+bf43Wgc7/739nLuB04MLSAr/Yyo3
IdC8Ao8XKgUf9JAsygUk+OYE7xdOywgNXZqfkUXS+lS1ubpPmxTiFoDiScB+vSJ2
NQby/QpvdJ/i2JO+6oFH6e5+iVTsUaFbFQ2XrdWSbZShi0O/1zeWKW4CXbP3tLh6
raQkyvQLeroJg/QE/3nXHX3kOVj7Yg8i1pDocyMpgJ2mO0GFT6DSyKaG0AdNzi+u
R0r9lfjbECLbW9YSMU6nxJ483JpgaDUt4hXJf4UTegRSm1eHKf4+bihrx7G60LGl
2GQG6wadQYpv3bYz2pHD9SRxrEI3EF8d6s/2FlfKkwkL8Odvt7IhoHhuMZywaHy4
Z1y9z5F0ZPh+YGClDXlU4bcYMkaHLGQ9BwyQkZ9//V2tFsM9nXZmBjgKem5ZEaTf
N5R13/DH0jex/R/8GSlvj4TTdBp/HjuO/lfgMv0owzyFqB/Gx2bMOty0bbRgC/3F
fggAfgrFHu10oze+hjGjkO+snM4imwKxj218DR8pirGNBLQwEeSK6Pv2hRqxvxkg
1iscdEY/oOuY3FKfbg996uLGgIRjWTmiEgB+aliBFBdKiTtcFd50L15HKYtiATDU
ROe3Dts4oC1DvSWx7p7QRlCZLV02gvaG3R7CcE3TXNOk3Tfn9+7oLxf/0NAsVpfp
MIeaJk5xcfEaL6tftyRzqGVHDB1Tcqag9KgzeengXbA9uJp6Nksd/46U/8FMUHvL
Nue4yWov+RwWRQvAUZgngL4MQBzb15lG9EM2ApkxKYvjnBaInYJs6rbYZ/G0JllQ
RUkY7DtGgpGYtw4PQdtLcukQs84q+6ojP1DYHQUBqQh0tbeALAeVFvCCFRrN45dF
5mLmGBo4bTU0/0dShUpf4YT6JNC2/LNbdxJxJP927AyCU+t9nj5QnMBwN0uDZWhW
lRQFCQQIU9doYrgo2QpaI0pV0tkfvlatI1MyvNImWU0zuoZT6k5rrxprClHO9kG2
iVHQLWXLiRu8jTEpiSXJMHoXY+id4k4vkOlujC6fR1TSg7HQ9ABMpEamqmPBmJvh
mkNAF/z7vnrbF+sjBj40Ej4gkug+sgIc5L4ONlntysqON/cudbbSLLEP/qc5pii1
+A9MwidkuM7fx1L1scbrGe8i99UfkQmFTgfIyuTp6erak3KZOsVIrq1Sn3TiQwP5
I7xs8ndzKFkBAvYOeYhPYoU/x7kS0bEOkFvuesrUtgxiTK5GFepGN6sUbeU+zUdX
f7MjRt7IpiOgGSrBfdmz40AvFrGLg0DF8aEU97f3h6k6dxYe6T8VP04OuBFM41Ld
od6aW8R3mTdaTh5rdqOMP4ckM3k4hOMbcEyDu1J4mctcpIZ69vpIFI0gx2co6t7b
F8ABYRZLnRWg8V3RNfmPhWvlAhg79sV8ZWaCvpPEkBWrvtyjrT1AmoPgpeJmcQIE
iT91HJ3r56tU5jNNR9pbPwSLw/Fd/6gjVHJnPGvCZA0tWxFzTTdvKiTaW9ufBZ9I
Te5v6P4lHCAdv7BMAf+r0O/2VGWDCB3Odfb0v8VpHag1H7vrwkmGKkuv8oampDdh
sjZpGmCZ13Ewy+2QmhY3isJ+vMxiwsKNjLiIW8eabKaUC1t8Ig9U8Cms8XHFJoiV
EEcLkiNHGd7FWwZGiLqe0QPGSlNenXohuIlKo6RA0FH0GbA+ye5dxzEY0p7i2S0J
cTeGTwxWMv3dMfx4qFJL+0IsDig7W7TbOhmlwol6rRLV0D3nNhmNRUAKvPQCKbsz
YeOyoj4QhhPerBZIJw0Y9AFDnsUh8cju25lz1pHaRteOCZi3nMlfthq5o2wV8VvP
UbQKsucFVlDxxN7fe+fZu87ey1s4RMooSuJa3DNm7UdKrXA/GvguTRrpOINy4zCC
Mj+5l0TNo9qDfW35hTvnaE4lhgw/HMTYoqShEQqRG8yrhShQFe7h0Pa3unQfZb2W
kYGcmCFoOEXxmqhP3KpIoUjQRNoD71vJDlflUWFPlGfiL2d15+eRRrsR3MlW1LoB
Uiw4rleSwvPCy2m3aWFi1rpaZljL7D8i7lT2n7l40yd5p/YTSWRm4+qIHCGwdYO6
wLajPLmqIOSFGvTYUPjteGQM1XtgdNZp7aFlQb4Ywo6ddBJBMUbVqkT+ijxYe35V
TOg40vdHFwcJ1hXaIs0aTd0RCZZbTe5TTfamZ7nIPPM152aW8EwW3rvsNwLpoCJI
o3KV/ZMJa+S0cLR9XHolKYap1/5DeS056odffZh+Kxy+JOfjfnRW+54KP+U5VRTR
cI//kX5vKU2x/eW7xH0ocaygD/ZF3UnzDfAnRHe4T7M39v4oJeJHRw6dmKRHzhig
8j9dXthdBlKRXyV1nhxqfGH1Yj9oC++pUnPWq+8swkHqoLkV1k5g6poZR0C3o0bj
4am1enfbiT/ch1/QsXRQohZ+3j5k6itkVp0BV6lal3oC5KnAERlQ6FoXxfk7V4fY
NLrAI81LtPuMtUDHMw/QTA6ANBWLRNPVcSq/fMCSxtdNKD3dzZ8G0kGMM2Z4T6hH
UG7Y2h7CvwZIZ/ap/ESqx6orQTMHCiUPFUwX2P3MTdVoI70EQ5DiIT+MeJklZcT7
56Jk/X5GkcX3tdpjpeTaqoHrfu9mU1W41CVukMkYceBPpJTZLfzTXVe+kfjisMxw
cG1AWcK1Aoo3RFurOLtihk6U9btDIv9+L3/JeMPYE1LXBvBiYkun4QlLoNf9awkF
l4wm96MxTqUayrXeE1/EyIjU0pokXqX1V+0b5eAd5hIhPk1sxF/iXtHFTkWFK7CL
mVEXMbISAjCuhop0GIlbibgrHy2q8aAxT/ZmG2RJRSXTfhKQa3WSMO6AOJWD3+Zg
VLaDymIf3YpPRtFtBma3ds2trHmCcuzxrFZD8SUPG+h4uX9U6nfqy8D1G7VcjT95
6ubhdvcFkkDPlXJqPevsyNrDG51Njhps5Z7yeVRblJT5pUKdFHOPg/9HNL7yaE6x
yHi7QZtJ2OapyYdKcDM7IDJjFa+YjB+39BFRVZpAWkycrBekNMUkUrhJQndordDy
7Id3+lhMdsz0fZ4S7VNnL7JvdgrumvIuEH8KxwE9jv211UDtieqDJkkB6uZYSeUC
ynK5DjCR0/YAMg6ogQbXFCvzj3Ert+QZgxldPIGB9AgykxGl15pfmEdq9vI4sTkz
oOkyvWSXxpTkIPBNJKk6e+jJUaH9Ir/RkaCYq7z/i3dAf5vBgLqxbe/Gvle/pWMU
TfuQ4PSMxmtzwdRiAjFCDE8L2AL2LWwiMbhfnlLkuO9r1p/Ua0giYl2lWQG6QbJm
iGGUEFNs8CZ0ZLO3chaDrvFWkiL0oHJM2r4Dne4+huYfmMmPDgFOk8/+93Lzpf8j
BtS6OJh9tAR//6Fn5E3ThaZahhmiJ+a0XV6XuQxSCvwuP28hLiRiCoUyd/QfUgex
7+3E48+iKb5oo4suExCkC4jVe7z1D7mJy3vY/kup0ii+DJMEMkx63J70uIYTTRco
dQVeoQ/pjzFD4nbspjIOBXc3qzFMIedap7FEL8zHAwxhhtEaqe8AKobNGTAtih6c
sKaEuMXaXZX+GvZa9NeYnIBF1XIw645eikmKCEkQQOBrllM6mY9iYeVVLU1FPWoB
PKRAH6PJ7Hh3QHz32lMS7SyfLrg6OP6ypLbZQ3VosK9wyQ5K1O08cCntoinYQy5C
2xu7Dfz8LHj5Ojw4kD30n+YxWNDZMzOD5GZYpXn773Y/tOWIxr5qrnAfy50suAEy
xuW7Zsr3PsBZPwjudIvFQWvAP01pyHG4LgZM+cWzfWG4TqRex27v8sgkgo9FF7VB
4W2vR4SRSSFfjvrX6pB2956OzsoDaXIwY0gcPNu3IbyIBNtFQY3VVwsRI0pXHtRe
JHJaYQiu/gkcRS2Gbxzj9WAZNw9ipSIIjS4TaCBckP/1DpDVbxQGwZzG5CogX1sN
nlRbsJD28eayqugIhMPEHbwn+YKUSy5mDJ7x9KQHElW55USa0jkRHrpgDhO3VYSn
cxtui9jSDqAWM/Zm0wsKIVlUpapCVvvlFhIq3B6+RTy89ZDLQ0Xw0wcFslbOBpUD
a60+5hzIqcCpHat+ydeSvoNsJcuDOInYMOH6xEHuY1B2LGVhxTNuZ+wnROapO5b8
2gIm2iNfE9mx3xTgrXuRV+g8XaXS+dVriIeLPTEiFl02+H7EInbyR9dhFoGElX1w
R3jg2+hEVr5XJMY8FmroeZIyFtAqdZnV7yjQ1mjBF0S6dOwaaC2GJMr2kGMIXKR7
gRkNVhEL10ISgwB1xnua5HXdIeBMQJw0TwKhom+lFgo2PJssabfOKf/Gg9KLIHoJ
kwI/F1WUrGcytasuHnOqG3sArA8nXZ8gxCFdad/IjeRdRlEtQR2B/9w1226Cth/b
yIlhWBoCcGdFixw1ERlxCKy5ukqFY+d3CvcJVV3RS66tMsGLMSZlFWf9v/FjHffd
6S0CZHKYm67iSN0ySr6+tWgjLty8aJXN5eoxI1SLU0woa8WpT9//P5eJG4FR5Hpz
g1EhvxV97FeJkszSMmINe1jXRSZhwdU/fY4uPf2Kz+FMs9I/VTVydUe74YDZQc8E
fwXua0X0pVxDx/r85sfcJ0RpSFZZjEZiF+sOSDjHF5bhgHuohlcM1c4Snt5dvBMw
593iEGk8rme/h2pbgpBeQP0CaDETPI75m+m1bzZMdlpsfD1I85RrHyv0g97X9mbv
3wPjE8lGgyS+3TfyI+/CQVWD87oUPYougYjaupicHZThNbtV9VyTFNrFYB00Uuf7
/AOj7povrPs7JkGgX7wOBHAHxi4etWt8gokacTyjJR2rFGaoX0Nv1VhsCyldETW7
zJvNmTANAqHomQN5wXTSwM/4UriT0kIGGuXpPdsC13yBlYdMVMYNWov3UgmvA9N6
DuI+i1J46uwUnV0R3Y+VlIhFHqOCEU/dsVuJ3SDDXiLqY7yda9Ql3g8zQXMHoumQ
Sbb/YGhjV85OZ/4RpkxOxAydZIbVY4nzDNEngUljIFXk0Dg/ltlnRTQ51flnhB5g
YZ+4MQB2lMB17GBqdHGWPeJAaxLBzvQsHIKCgAVq74iL2OdlH9li/UVNlMYpSJrZ
EEoh2sqDuXq1f6UQl+z2HDjsmmlcbJd7AzjRsGvQdg8mtkPunRb8xu22f7p5l8VK
8YNr0rSqwPxFF5uFmg8HimRq0H2tTU1TyRByt1D4ZKJfZqH/GPVk35ZS+WsOfm7e
2E6bEyOkHuafNggX/l4bMTIRanb9AxcTOk6MQy7gAk+ShM4ZdRntBF02amLq5e2s
tRQtP67j4+7uW/E9h4Fm/qkaipHg2TyR8R4gKdR3ZH09ylvlgrMcEvLaCo2AtDcp
ugmoXBwqCPmcD+qfNla3yNtl1rICXFME9iezXt3ssv3xvQRUiaQoE9bYmYaWdR+I
q+GXLb4y+qH/xvrCN4JGVrIPlgyKemf345TntQnkNj+foW44fh3ivkIZt2SDN7OW
jkDcH93mbS1wYRrrbSL4yOhwOZdm3o7B/C2iU69DK9ZlH7FmXqD4dGl3LA/SBtoK
OW74BAEqvAzHsVYGetZkoE4gYNA1G2m1WvFQN3yKV8n8bIGynOyxinNKEffRbIKB
CTKWg2B8AWjLU6GE79nzKxN5lU1JQDc+bglMIzCO8MfY2iD3+xLg2atoaCcTmJUJ
QjEt0MZMy9VZg4fqDTveJ8UQOgA4FWb4KYRDwF2JaRZny+65l3b4sZfJp7BKFPK5
jRqyZrMXEOlkryxvkgE/U60ArLY+V1bXpSlO+XgxTmQcAyWWttec4Y28McsioCne
9aPIul3aEuGoB+flUpjtWTqIX66ARc5Mf+DfKwQEBMaJGmwuIAynmEtAqsoiBpbU
Umuh9EvCcT0YMgME8EgtY4d7ZVhuhRz2NykNF+GvI7xG2FFaaIu/4Kw1Vjx8zNT/
Wi84N9y/vtY9tNaqKazdyJKpdErBOfjtb8ZVIWnVysXB8CG089db/xhxIys1PucM
4ltInj4dc/Xy+BUN/3ipii798l4OEK2bMrJ7DCPVwiRNblhr4XdUNoW4ChFxv6dz
tCEPKoXfM6EdLZD1sp4EBmXy8L7EXUa54YCuZP9htUJaRvsGwsafBA+MX8PSxeqj
j4Np5XDQ6hNxpfpzBXpy8SbIxSpFyuislBU+/cAQQRDZ+AwbO8pIHVhHmWXESl42
cQLEiaccqOYTfysDRZfpTjK/BD7QZu9rAFAAXy+mrWb6ZYcY+3rxWWT0d5GU7jhO
7hDJuRwKo4wurl+0FK3MZn/20LtEZAHeEee4wskgurIMLBeIqFTzIrUw4v6zKGkD
TgrDlPkTLIMAlg5gXGDZos8gdVIOehZp3FsnRK9Zdic2R6dsl0SEwKvBAGbj1lIt
nj8OvmLzYk8YIfLe+N3w6EkRWZJTCGqaT5tElso48apO89tJka6sySnOcwnpAgDm
jYWKIXSjyePLwpeD8xPmcdBiWOHfEfUTHl7g6a2U31w2mUS20pRMtHQsYGeXvhgD
vxbSkrz0Em03scxfnsBKqUwsdAI8xugaDvcWk80P7Q0GoyB1DzwCaEbE57DZrgKK
FRl4CiIJyiOjvsRP+sL5JH5ypCL7qneoUlQ8u8lpUPstDMMPoDhmIK1z9r9zDY8w
NDNmCmB4djl9tFwABPXOUqeIWPCBQGK3Cn7JRiUcmD/2KCy4wGL0DgzfMADa9+u0
KvaW//wqupM4kYyIyiA9Dmy0fcR3qtFMqdoYROK7UtF46TAAlJDbeXb343pnNEEV
rMxFMAiF0c1oEsLnIu1cCLVlaFrNE83k74JOfpKjXDl6LmCFj++1BjnWKksbUAF1
o84HzferXg2J9hvX5UN6BdAumIQDAaysCkPGL7951FhioDbhRORv6hRm3ai4H810
NGiRNyQfCfSkmh4sc1EwJqFxIFlNOdR1UsSkHjJOnVbfktXG7BFh0wED5IcNpUmv
rSyykPrx7Ih8hDLLwHpxKj+GIK2BqsJL3JtwNVp0SW+os8BfejbL9e2RSndIhc2q
jQzwnC9K8iZQwEEPYwqCxImYBKTeUDxYpUoCIwsccpWcRQRVgc+xJZJsEuNUyPmB
BANXqMneXuKpEINf4zNO6kNeydh6YCCkploRZDKEUfbVESV9rLlerwPehP7Hq+Bj
Df/GSfOHTm1pkBR5C8GkHgNWvifBbUGXiSxaTUFUY03gacoTUJx73WStJ7aZPOh2
jlnVXRgcPeMJS/8qM302DqL/I3a864UBDLmEZS8zjCy5fVZIOMwI70nEzvXkRGxq
ZOy7lOpCERa5QHLliDeYeUVKZBAqFHQvhXH5f4SBuP5MbmaGC1SVpNoQFDecLypj
Vn7v/K3Dkrjoy3MaZdFHDOcOTxpgozg30dQ1RXS4pn/UDhtHDmxpUpqS44HXJpW7
tIG5Z1fhHrqBC/FgpQzLH/JOwPqLW6UsxPCOeYv4hrwctriw+Rsdc2oonf/JcqsT
+c/isz7uODuw7taeCd7hKkMy1rvnSiHIpLfu7MwwlU6rs9hc8jn1CW15MM0cd6g1
z02NOsqf9ZN773v5Ll4fD3u/7wwWAbGom7QDVvftMhDsBV/hlfHt/akNngYeoiUB
Bqr5jKkznacQOB+tTf+pg/HS4AFuxFODiTUrG14IrbJJ6oq1wtF+rXRGeTJ4xRkH
O78larqrxy03I6nAoaqAHsKfCGcaAk+f8u840RRZkGdLD/FMzdJxl+8H/Qu1e0QM
K8N8pHEPZJpPY+DQJ76rvuLZnKkXVt3JbFyrwOvMlD1nyJ/gyg9iWbZPyZ+Yh9hX
+WEyDY+pNOdGmcOMRRdFjqcfRjg4XVwNrBun5oSIDPQrjGPIKtYoMEJYOI+kWqT3
nPnID5Or5kZQHr4Waw516fhNVVvXXbtojTj/otf0DzEj0ctrGqdaektB4JbYiFbf
OEwMgnWj7mwWj5bv2sF6DDax6PBMLqlhNjdwfRNR21llyKYsYJrmeIdgi0UmhPI1
xfT5Rxhz8YNc18g4UElZrSdxnnKPacdCf9Cica7ryd8A50GK9LTzo6PICga5F0HB
aQXjkeu2bVy4raDq1eoLruW3cdlwekFfVvlFU4EB5DrnOAVUnBAhH4+bSTaja4TI
T2xWuv3CqF0USoWSiA3+ac1W+47pntxMvQLvxiE8Y0p3XuHd63EsUwP1lTI82AOn
MZu0ez4VSuktNdoSLe+q4p6e5qgXfPz/wZy4HOJea0UqgkLoL0KPAS3DmT6hnsaF
M0ZBO97LqdxHwEFskHQPVpe9pcR9Wzng93UHreXIUB2L0y3tMWdg1j3zv0rpRJNa
Yf/lnOw0Rez8D1cKv2VtltpKZnLDQZPdmqUsjj65+ml38SwAT4W+/UCW+P6/S+8K
imHxDpO2ThLYQ8xBAa9QQvUL7wxH9mBhfiEQqaiCw5AGdmLW06rZ8VT51ZaVJWig
Q3pGMVDgRVZ0v6/FqTATbla9tR6FWq+4/LB7jak5uiFdXfGKr2Hp3dNmF8gjBQaS
X/2a/tDnlYvLpngZ4xrj9HdnGlbbhI0t1HYy16HSRB5BBR8nHiuazpukTYEryOTS
phT4H1q2fJVXpnzCUXBDfyzcnIjhfcEXIJvU5mLFuHilmKm9XE4ZLLTh0fPpDDNN
A2DY34pN2U9QzGCayfRlqIuCwKz7Sz2b2N7OcVGSLSLdWmnQoLJo0/mbQozlcPha
Xv9bUfLE6g18uuHBUASxnI7Plbh1BGOSH7OjcA4ljzrCCX1EFj9sPgT8hZ42vtgi
mZQsu1izRs7hRwlW8AGJrBFZaGCfvDWS+l5aVXgz831lXzsop/jbsd655+IuuAyX
lGldc8gRU6EMuwK2BvKUOD1xyka75WQwbriDPJH5GvMzjpNwRxbcdCoMan4Usn36
QSquL11cH8XQUnWVrFZSsh5BtMS7ozsCNOjXp7JQrIwI+vG6+8Cugl4atvg9bqH3
OhBaHwPtVtCNp7mJoM6sic6B0EViA2wHC3f3Xzy1fvGghbWiegXl7eVjDx6mBcz2
9B1YPmvmZMHodwNPth3XdiRmINEBdrouBVTkp6bOvJbsSj2iRW0snYvdOB75KIek
ZZmpw9J0HPi9Em99E6Iewf1f0h8n6VcH+Qi0wooFZC+T7lH2lvt4rBvmCm2Bak8m
05pPOqetp6xuNWs57HB5aGTgyMwpkwJQMSlbzdJf/3Smv0/9Af+Qluql+mYnmKZu
ZStZzo8XEWNyJrBdNbj/nCorxXwZRu7vPk6LW7+c01jKK/s9Xo4xJLgHJVmwlMGJ
4Ffn1ZSF1JgF9CuT5uCozusgmxZ9qQ5Y1NaeG9bL2DLs6+KQbz0cTJ0VzciVGUtP
aX4hyoHeSED5iEUC22g/n+bwMdQnXsJ5RC1D3qFU83kBH6Q2C1TCo+CEcKQVzqS6
Q/MNKQ7R05x/FcOIL80NPb3MLw8gjFLATZSPSASZc2sNG9ZrnuCua/4wQDP3dJfb
CPLagarGi+ocjpC6mPGbhlx7TkuzpxPwgWtRowKG/tIvrKz7ePu+PeQN0Mc0qyOM
wAmp2f1l77vrsou3rtPnLKMeLQODZ1YBp2wpTYdzbdmNFqSLPctKy/nsy8wqZYGO
xUNWw2J9ZRIPpGrGA4moVd/H3ONW9S1pg+on3FHMOQQx2K8OlosKAoAEps+6Zg+D
bxaVQvnbzsrjA43oBDXEIOCWoaV4F8AX4px+CBGeLFxH2Z8SXmnWOCGyVaJQCavr
TumMdBGQ5hXeCMum95lFKgj+UbAuwE9YZTf2QknozrFoI5VUDMJWcBW3p8h8i9xj
YmdVbfmntx0UUk7PsnP7A2eRycFxwHglgNNom7ORtvQkC/K/d+UqrzPgiOZcTiya
vetmizEubZkwxZwkfcFhHb18UQpdBsYUJBtqfnozV+zVLLCMYylJV3XoCvlPutrB
Wp5L8Ya+UtLV8FDnLuyZ7eDW1DLTtgaLdE8XucAsnC8kd5N+5L1JXGi7wmTw1DuK
HM9gmQzwXrzi+cr3fAfV7FGrXpLWXLlCWiTklSsc1xyDKYDqYkqz6paCMAVmcoxj
UCVGMVabVSN1ibCtOCH8Ml/9eNxPbiGn2DJbdtGxZdhmhZG8/3wJbmDad7YrMk+W
Gcqy/F6B18QgVZFlq1Rqb4m1z/3rREtJGxCFJ8Hi9fZFCuHQ6ntz9vwxyBZeF82B
82HeEXKU3PAGzbY0Zt8LRXXLiwM+QruPlFhFKa7rp3UUfjb2TBVs1WYtubLwbix0
Ti+U8WY7gKJVcgPG864s76DCT1MAK8mH+ACJ8a/c8tPiT4KPeSvDpffpIt5c/d1P
PKFH0BuaA/i5m3p6AKene34a/ZSaQvy2gip12g/HwggzYH+P71BvE9AkIEMppu3R
UE1askyqfgPFqKV933MMSkA9gYEfmhdPoyo1gBnsUAbLElkWG2MteQCfUduMYr28
q52Jo4zkdmRZ49PMim6Fj27GluK1sodDuneyEbT5OfMxPUsbvPrRxT9uMQQTSmyx
yM2ksR+/9XVIneMKYqLo2fuKzpnV6WVH5yAh4vKBuuor8ltntGbCJOuLqKM8Ad9v
QMMSrBiucGqG6FAtCRa/iz6mlz4n65gPPMGvlZpUucl78P31oQzM3A11xqy2/VHW
YRykhaRP5tMb9FpLvL11+J86jdq2FKDeIrjGKIdqSQSvE1gFMjOtFGp/n+iXs8Li
DK9BMq8p2mlCSCOwycnpYMzzHz9pP3B3P6JOU7KxO4xwsEaDpq2fZcB8ihdkbyqn
IwbTYdBe4/JgJoQmA3NirgykJAwFfo4qlGe3bPSLHUlHeS5E+1QuQlP41bfec3FF
c0RUEnGt9hY3dz1MEZ+nLeRQ8ZQIVAWPYzfW0ajFEhO3L/vCZGHTb925aGgUUgXQ
jSR9QS4YH6zDKfGMZeB64zVD2D4xotJI32DBh/R/9ySLGYvYxL+4iSXTqF+Ite1K
wLgB75UmcbIe0NLN3x0Rp0xsLo9gTEtrPWA/YBTn48cwswELhQ+pMQyLbyGFFXkZ
FvD6dPFGJzx6EXht0Hn+06AnyK4wVePaGM2fU9jcXUXH523LwQs92rMaWIutmsDE
QomlMU7LR+6t+A0Qj9EDYUt/sKBxZFe0xHA4ALi9KP7KAMzO0aNZ5Ti6Oj6l40aS
B6bwaljdNF4EZ6DqLLZmYV3vi/0HUXBamIArxmcmYmTsdKei0cK4sL2CKuZzTY1S
rvItmL4eprcdV7xpkYrCRChBPA3moOK8uJnkefdZ7fizlEA28h6+H33fEh0vGtyF
Lm5N/0khreVZIXHugZZnkgnR5W2N+dGzM1kj8wSFHubx8fbsPyJVP6FIkY/YL8hq
AWiG4LEyau3I3z9o9sKwhMSvbw6Es1vcK1voNbuAEmhg2qzSeYJN9HsASeNH2YKp
O0FjZiirrlbeojHx4FL9gNq1t6ATDUweCSJFInpBFU7vAfU+6WEFhbLB1IZfv65b
QCwh9TJOB4sMYj8HIw6fas7dBcxsi0foZr88MQ4+1rQMIfioyf98eWZJP0fIhu7h
xiVUO63AfP7wsgZaJ58SbVLgNGq54y09ACs32TK7YblpUDDeCehCmffC6MSGBB59
7r8ZzM8v1ro8QZQs0GSoJTrChaROuYBqcSredPIfHdXmWnxXnkxSsjJzQ8Lo85rw
wrkhxNV3A9m+p7rkdGWXR2j6hgTBa1jHHp5MfO91+cewCnafjFgIsCZhBd9nr9yi
MdBC8S/O4BrBy0qJKafNDxGNTmKDaGdwNsr5c8DL5CnbD79cuIgiGnwR31pXmnrP
I0zxammmoUVGKp3ek6lvE3ce517UhJnE9HFQ9ePqNx0vqT99WgOX2X+7lh0WFRa5
XqEE/5dZJSx46G7HJuwj4znq/qhU16gC7PSMlIxzgFCcV04tv9vpi+4hUiywVLI4
i7o/h7antIwSd8j36OkvFBxl689otWPcG7YJlnBIT9g6TfK1dyjHWKBqkU7b80H1
4lQwEzYXls/hly2759OVXCzR9pWEt5Zy0tuXSmGtiVI/3/WeEH6Ftyz8w4IqYd6n
qnEPT4xx9QqhITW+1l0bnNps2yRsv1jsgpd9B1wy6hr+xFQmtWanaXVnaYo2qKwc
27yzP6ZZA9sJkp19ISqqPviV6BVVe5GHt0bB68z1f5aEXj99UueQjH4HgXFMIjpy
GXMvp4A6hyrh7eNvECMRQPpGhD+RNa6P1OdnifU2xHrZM53HLkl3w9PYTTKxzb+o
C7KTpozd2paiLbnjlttJ60hdHGW5nSN4Xi46/4ylxJStO+z99wWXTa+UR4/NdEVf
PaX4aVZ45ykXebRPnFaC/iWitKHO7n7ab39jYEMy+Kd4zC2mXsPuhhfExhSH/hoW
i9huHmU7O3wg78drfzfDovqDRQAi1FgX5w8RPLoFgGw4CH3ez+OOL/yFta2Ty9Cx
BPxiJmyxMNgDXjNvc1pKVNoi/N9CpP5uEGIlr3lw8O2+IYIil6gdV+OGYxHNf0K1
Pu1ZEhiyjCcYh00mzrVAkH7g26dS+RDYljLhqrJN7akxlHPwx9XGJ1FIl8n2A7aI
hzZiVjmMo+veaf9OvaDRHyjY/EK3WDPCwVhiLlQ5F7pSOcu1vAhmpLpcNjciDF3e
8qe/lGqdgS/dztcxh3tAP/aI7b+7Re8LGBtT+hhBdmKgY/oUi5/Bz5bEEfMmJOB1
cwu7TJ+8qzQzKL7k+btFnrpNJR7vG1ki6kMsAF96aXLzWtfi/9QKVxNI4Rkc7Non
yg7+8/WDGiG46P0RJ1/RA/jIFn1jnKDXmGqpckGBc/k7CYEMZ6/C2fwFUadoWWSw
MImizS9vPAoOwgROkrQUHn4wRwsA/tGAWlxgobg49LvZXj4ao+ff+v6oLV7/Fec6
r8LWsgcy5kzSORaERumWKQckuUbsAyjBiGBNhdMUNsN3oPzmdUB4Mk6mfVSpoSrJ
1LJo/0L+zexn9AHk1UGH+GpTnggQXThXkFtE78N9JgT7yOKMkNZJoujepbsMblCn
y1NwYmRMfWGDtGsJbPf1Ve5LZUrWjpDcSz1fQUWbTPYm7Bg8wEiGmmfahP9/d/fZ
P3HUK5Z7GYKjYdJhXttit+7nNFZR4h9J98yw1w3oKV48BtqfFoYQ70ipTrvpA/Tu
8H4WNa6I724agtCFbcHSYVgWGFGn+LNnvlDslI0dJg/2kBbYguJtu3Nj19wlYVMX
qq4wjuZBlyqc8D1vW8RZO+5E2th5laRKYrJXAUus7SGz+qHK0cZcnAPZpRlzmQwu
1btJb+YouHB/+qg5Xw8ZIr/oiuTUYXex7fEUB/5NEWkhgLRqXU3JLwH0EO4bMRHx
QJrcd+dzzvwkbshoFx5zil/XowrebGn2lDNDuJOboNHQk+sQ/WxRzaewS2NgY5NK
sR1acKxgyJfGX8EcuBvokItUds5voHq6333zyQWMemblRsCH+EfMawQrmbltCUBQ
KDGYnnt8sKf//SdBvDcUMUsx8HOjAsij5RwSAInPbRMcd2HiOUcMlsJFEIupMiFc
YNFprSTovfI8m6k/eHw0CtCxfOSIrmCUpr0Zz04gVOIVjFezhFWEV9xSNsSQhB/O
SxEvB7/6Hl1M1b2RoxKWURMRWvF8BZ2WNCsL/YO3pdPV1PEQr/+qcgFVxG6N/oDN
7qPk40ThtrpfmN2s6M+e6ncDVhrwJHdVnyUK7oRnYNCi9a9+2JgkEzzTo0YnsIWl
U2e3thJdzzLrt7gdjZ8qY+ku1/PlIEDit3rvBm+D9uCIci7vgj+hFnn8pOb0n7xI
uYGD2F2Juafrk3KzUM1kpkjXuh1EUoXYorMvwFztUmJvQAT0isXNsHTqvxJ5hPHs
4L6n0HQ397OMOs3Mz9OOfsW0eyM2Kleik2SkQIplwxSZ27Ih99sVpZLrMhefwKlj
gl6uhR430qsYTKSFZtiFBP5oCsjXfPSoHSgIah+c/LFRSk1twrsQOItiP6FciXPB
zPAkVZ9/yh+zaz9KF6Tmz361yey7XqpZl8qyGdFLYvTJ9hSCMoB1KlQrnAVdgGcS
d2uI8h+nnHd0fAuFyrCjNmUzNmNjsUC5rXdKKFdWVYpfItBbWNy+revIXx8sGiip
Q6z6MvQS/4rGQAPc/0yCbEsfIcf1lI4mOhHO9A25+S6m/crEHW1w5EjLFsQwyM7D
M8RXIjzof/gO3EjIS4HnKZPGxi3M9T/Y5lcZc33VjtXnmpenws7MsQ4FtiRgZS/j
hyMSuhPlii1jsCMdzlTBBZBBoWqY6YAS7GrRfUSaX1/wNBYfLSv2ullPZMqq/+vG
+BEiDIDsXnDf3S9vLX+MaxdQ9ngkA1GFn0SwDQB9R0HzMKWg+ROEU4U9trqdYq+s
Jk2ntxYCZRLSi/2PHfnCy9e4ZH7/6ciIVtItFuraxQZ+YJDpjOtuATycwEf+42WZ
v14OSLCoai2NnVjOY1qKAe2s+P6geGHNx6wAESG+xzRBfwIiVI+XhT98oTcyIrAj
3MhxHIKQZxUHtkYHGGisptxXDdBLGCJYtnqgqzJQNDmBMXvnJr3qnpjdXT8bjxTu
zhhql4HU7JU6h0y0nLq3RxbT9Yh+Ybqq8LSHWEZONImiOOHegHPVSks0nTV/w3D7
cw3vlpMjTJEEXkUA4nBi9IEz4F668juHvUGv+zEdyS0Qi6R6lFaEeOu/HBijG66z
7Cz/q8xRg5GEB/8jcNG5A8ZLxpWa5EULa902fa/eKsDmdUZAQ0qw0VXOGwtK2clL
+eTK4wp+Eee+Gm1QEoywZ8vPR0H/CZIinFMl2iGU53saGaKTiF8N4vgBHkDoNpA/
MYny2rdwNDMbUv782UbLUg/CFzxhBrkvys7V5Q5t/mirZSimuwEbXPnfdhMtH8ay
LFXLJtloRbOytm8Uw9u8uKcjDgYNX7A8DB8RgvOQ6/Ijo7YixyQPjMJyjl8nYjYm
a6qkoGSKdZOjz+gXyBIuY+IwMYj1bDEvlPdiHYD4Py5jtQ6DOvFz9d9NpJSeTe51
R2DrWKjdlNJb83YP0IwI9JSjqQ9U/BdQTtl7hk23H8lxe4AJMk5RnoKI7bo/eoa4
Yg+fRCSu3yQhu/hhfhfRCkH3wy36234Dq2h18EWk2peAboK1G8R/MmLEX1LR7EVu
tvswc/Xmbp0HPvQLcgFpeReElUy/WjED0q4bvsPr+HeC0qWwESbjPSWTxLHSC4NC
FTa5BLnNsZy9VcZyC9O04OI4oRj/6PYYvdtKjFpRoPTZEb+8nNjKwy9PfmNVSujM
q6L7d9rs41yJZ2NlvsCN+N0I8aqj6OWoMvXd26qRNaiqLjpmGb9tD+fCj+ww56cq
CpHfRwllS8V+SPSSqboum79fsVO/r9Ta1bZX+e3imnWq0aSife+PkaaGaEMv5aj1
XaEytHGejV6RKVLRQnCSpkHx8fX8RLw82ET9735MyI7d7YGV1d96qJ8Gwq+nppVc
gFrppxe+3bdlFsFoVN1Bhc+TS1eqDmaubb8kR/OtFmdPYuP+TlFF0mb155LUXXDY
fT+HMp/z60Y0UbU4J8zCi0wApiutyDooshNvAuRGC+/5MnbZ2+FWHzPDFDCZTkTM
2N06khRyJW08HQ7wdl8u+6e81BZ8R1f7PWa9NwIgADpYPIqGTRPDXGu0uVyINIES
0cgsmCeURnN1a8vB7WjYrs+B1tT/nIlaLI90vMRxOSl+ffY0XqCAYc0Zn3H4O+pB
7XDWn0Ze2YThapG5nrqkVspQtnqp28jYZtGJBaCHytMNNqlLFOKZkOcKiesWO3J7
Ws2W9aeRbiUqqOvoMmLzkfC3IT1DBD1w9o2NPn2kuFerSpowrqB2r19CLyfeP5aC
LqLNNVTjWjib5b13+v9Qo7G1oaO6+Z2wO36zNzBM5o+QEh+9WTbKzfGUMMV8EVLl
dBZkIOi7nsAzN1mcs5y/1wUTsfBRuajMODcS9IlGFhNQiuxoUiycTzks79qBvK5Q
lBUIlaJ7gocJp5wEf9nGxoxm/58N+6+QOj5nT+reuqPdUSHjAY00Y11BM0zPGwey
2wJM0dnjCK6DlUnHkYX2H1fD1k2S3/Ce7hroorTFLSvWrYOf/cAI4yvQ0aRe/UKE
VWch1Sqtl2SEzq+FphS18qq5OJrnGKDEpA4J61Phtvp6xDljcr4t8W0etHiUHg8o
gUwyYlOk/SLNVHtO0g/b5m8CgWz52VxqDl8Ak/MUozho3sWeHm2JjJ8GRR61rgTR
EXC2GY4At6TL/SW9sg12QRfFkjY+StQBOZNs3JIdmCd8iHvOC1NIiZGi8i9LPGMT
6ES5NQxgH5cAJiF2WXmOejcL+DL9//y+7hbKJAZq0pTbu95ASkecq2iVYE6rZhXM
wqaBsVo6hnJpXATWXQDykQDMgDG6btsR6/s8CYb7V9h74/kVIfTMre+EymLlMK9h
HH0Ny8I/iOdWR+TFbPtGHSzSlkRWdwWft731uOUNgJ3QYGqqi5KgVhI7wkR8zNZH
ujXXACP6ubCSNjtTSXkC4TTSa/7hBxC0C9yWPypzMroUBxLBIj/7ZFwdrweSDIpg
LHRF/NIV+l9gYrTJuT6hQex/AmGbf+pCKpBTG5f9y7wCEKjYfpzzmpkaLL5uZGYv
K/23R085rKSaYmC/q7Nsozdhn4NiAGOfHTlhuGGp9R3k9cUki+braFFQG2T5mDNX
ViRLNtfyHB+z5JMeEhK+ik8zFredgulZcaYoz/mVceB2wt5IRjgLZumUz1tlOJNR
a3JgMKdoA/7PEk3JC0mQFeaVw59ie3Oducq4CisFqy+COZnqAbaUPMQFbzA/fg5x
xODzpjBDtaYETPOCwpyQtWGLXF6xJbWTFEXdCPP0L+oOyxS2RJk47A/hsbMR+Ej+
1NaRlvyJI7Wd6mdw+3HDjUhvz2EryynJLKM9OLmxhL/lVJakJ9AD6MEvZ3EqBlSA
jEBDXwL7rT4Slvz4zsCMFmfm2EohNAGv3X88qRhQoXUf3TUKayoP5AN57k496/Jq
ZRNo9fcuNw7HRhzr5uBnFwBUhRDbPg5gjaGfRYQeKs7HoWPEMjAL3z3f1F3YWhwf
ES5DmFaowfM3Lnk62YNYJArji3RTkx9+1tet12vCFNTxcf46qhN/3Ql4+4VKN3ad
8bbv5la0ix61IXo4V2y+qylpnLwC5ZYVosBoXXuY6b/RsRh5pkO4zv93ydexeaI7
sd6l0fU0LgkBPKyE0Pxe1IRbK6tCGHog3bha7nkfJolg11jlNTF8mtXxsv+/VXNN
m2Rg8ZuEF1IXE6/q7aLbgxiqzSmP+Xr+TmBBIKgKY8FeKqK/CkDkSQVtoFj4xaNf
dF6DvLY7IOxrwpVGYS0Hu1lJxax7VAGYbLDEQlzZHC8JTieuMESJP2S6gZBHURHk
ptNOhZkv259UxJJrRjlqj08MZMQQ5yvbl7rO4SRPTOaq/honWnG51yEebWauQlHw
xt9ILNr2dGcWkZy5Uurn4Q0NtYCvCjFhJ4yx6i0Z0zYMRMz4gAZaNUGq1u5xhZNC
1ZXnqkMnQPo9Xc2qaKiQMybeymr1wEivVACupfRJ3ybhepzJ+rQ0+WbyiuUo1elM
IvXQVN25/nWSHzpXCyT8zSzKW26Q48xRJGXIHDOJ4DjaMOLGxua9DopHW6o2xN/e
ytKFPp4Vn0hCqIDMcykpl8b9dmaEJNvleMVbq2VwcGBMT+EX33eroaJwmV+aCrxL
YEsNADe77mYq7bt49u0LlNFmwlcW9lX/oioy6SMydovaluS6EIExqXjg3Oh0T396
FPeYcLU55dped6qv8ptW4I9QUR6b9j+lMT8LI+HCIMtVcCzw80A2XV8i8FeeuEKU
5W9d0X53wToJCm1oQMmr7H8EtcIoHWDtFNa6RQrxaXv2iwWpyPmjWptd6zBHjkdk
xUGsgR5L5ZnkxJVJXD8DNFpPWMprNLVfqNqpRzmLwKyT7CGMVA3g6669SmDW1GnN
RbCpwf9O82/rqoDa4+NvEFjT4AYcC+3778JbMKf93p8q4QUnv/0nVHWaCqziKY8s
ujRZy1UKq0cNh4tG1ePLo7IAQ2aTMdenIjTjMxBp6AXP6b6s3mfj3L2jHloK+JVj
MOCYI1p6K90uVhuMkARRiSVf1fP0Uvm4YgWB9CHEyycZKHMxltJ3JbUTrg880zTA
PeCqaWx39IZx2GdxWg/gLC1nhgkqEwwCID0q6/7ADm/t/xhGGlGZYc1GqnxnyNs3
aZjnCfZNJlf5eC0jiBdfJE3PRhowCUvNdHMl93mwvm1Fsahkom3sF1dZtNYdBNog
t086NPjPVrXK3hpv0LWKIzxKKF5ANlyyr0v8JgondT1UgtFNFpWRIhJzYERIHMpk
Q7CCVzjg/PzK1SA88I3hldkUG3dpqNqtUbe46hPkIRuKMmE0G4MxfeBTUFsCQGjt
gDuly1gB9HpxeUO0AsIaFSufgRkxRHyrxZiLfViROGklZ4NxJcHvRE0qTRLXhQi2
sZJZdI5wOH8YsZF4XdjBYQwYkk/GzXSmSz6xgL97L1QTMYBHO9QkgFR6c39L1a0Y
HbtqwP3EBehKeOZSF9PlMc0xqFp4YRSTfO/CRAffjL2re+F4BMt1QKYigdX4VSSF
zsP+6zeWgPU/aXSWJ/bPUfD8LGqn5kISM2sPAelMOEnHPIka0F2KyHhtnLX3DHmV
lhPSQi8gl+njyNrt/+A6mqsnMvKcvorg36M9lx5KMdv/SYamIZU6y7iG2ny8O5fe
YrZumLZyUFvmli6AwtqcudeHIowqJW6bEjHLEOHc6zmBmAkHCInKzHS+V5ObijJO
yVOAkJ5CkbhwgVVzedgPPXFJUk8+kCIdpH20NdEMlnfUwOCqkvPW/7kfR4ghTj/R
d1gr8c8wzw4dSNIZcU38pn9B1PScbTC87xvNfTxxGBH39uoFNqCNLyB6pAT9rYPP
DEr4uvJtai+K38NNlP6XMt9EqVC5cYS6MRYqInGn665tgeMCJ+qlJQRiKvVpZLd2
NuqCa939pDCihu2kdvzSZQd6SdQtIxqmuvOICk4MqaKN+gsE5Ir+QkUVINIHK2oS
KABb83Z8voh50ES0kn/PUAnaGlUYvf/aBO6/M8asGrkn2OVu3JjyH1bznIiQDC9w
uLEk3Qiu3ZkylG12NJC6OrJni+pY5yDlmI9H+xOqC6cYcllBhX0FklRPNksuHLv2
W4Qfzxsd9x7QHZdwaEopt7Q8X8lKEOSPTY52PdjimXF3UOJb5dkC8Xj8OllG1b/l
oRv++vW4YrfCzAvwkSEQ2XBCtd8VSkfekt46kcPdAdX+4ljz/TRSplkOEHzRJSu0
CxQwX2uqlrklzWbcuO9szb3bV5oH9LEkjCHD+c2Lh5MRN4d3icq40GDwx+vr8roe
HM4P+8W+53TCo94qzv8nOD8bO48gIs8FDolephcpw9us2fj1YKLPB0vTaEruK+gS
X0bec78jiNd92/BWSzVQC/XVTZRyFMCa7i7whPDJ50aowRsdvmpPufL5pQNcwOoU
bYWa93uirDngA8Lq8wZTBuA/bmtJpyRXa04z4aO+DFSsW4GuIxFxEybXjfqK7SHn
9ZYCXdyLP4DxDFi9tjLoftVwDK9zovniyJPGVszH8qORqsJu0xM9e3iZmdb6xEuu
5ejllukJy3K7IIf+hE0jtrLVsvx3YfaWfjQ4TYUOfqL5pXoHFMGWwALKv6Ci36HV
I+qvZ79A+XUkdTTQgLyBleEjmJOnz6fgFZgtzd8c8ZCq6CDYLxhgL5I7aS0nzInU
CYSEedHPN2Yy1EZLtK71DWM036RCEumz3/EcdSWE+jsHf6hOFo7V24mzdPwVb1e5
1Qkmardi2AqAldClZR3VmZMnJ4g9iXxGDQMydoj6kJMhVsUr7/Y7rmq5m8zV6udW
/QZ6ciz7anN9O1Zj/HeBx8E3R2Iu4dSD8PIXvZwv/MJDBU91WAJFQIZ6IqseZd4P
DEXkAsBJzNAZ0McKiLvsI9rYP5A1lc3Lkr1aqlBsb5fqomyFdwicOmdDqxtJ8KDV
EZ6vpr6oDI9uPo5qJFIFj7nKp2sa/mLITeRojfXBO6AVwyXPS4qIORsLPsPzvNAD
HqYoZh5d74cd5YkpeHOwNONCpJR+nz0zncE6UX/CBemA1BYpK84SjwABPvMJZ5GY
CjmssggZOU3fVUO+sgtoOUqYj/9LiC7oAnNJuByUrMS2IfBAGgMnq2p0QhBIPjai
2Ntfnnfiu9KL3SLnwyhFJJR0ZWmzuDZtrkgPrpSMp/298BBVsN5ucIyGVvWJDKLZ
RcLSflo7S5UVDow/9JHxEHQPrqRtE1agt2rsSkdU7mDzFzwfO908MKhhveKj4vN2
CvG+2WKuOApshzSsksHuS6P39QSyn61yt07C08FlnDEB9aQZeZlMxT5CnihajkKr
ZZcNBx0C9YbndoQ75Kuq+y1npCbAplA71L7scipWdkLuDdtX51lhXESEt/TJODkK
hPpv5QKNs2m+JG3tMlSNKafMUMX8IwlRiCWbgHiTc0A/PJ6RKBkkjxt6GwUdVJQp
SNM6J2dp6FSpBkepeeThku4UcJG7SYX2rhZ7vDozZejqTFNbB5UCRP6vKbIZdyr3
wWxLorSsU1Kc0whDSzXmoTv5NQ3RUQUwakMJA12xoit5bkFY6tSNgmapNK8vmmxv
+mbNyuumjsBZlU0CcHHBHUMH6FtwtVk7US+rtWc9Z6JL7hosojm4gpbDE9Nfuyn8
SOuGZ5kW8Woxb6XXGfuGpnfnEtSI6JZVBBNuO6ky5+2AJDWazI0za3fg3w5mtjW6
aLIwWO/4oYmSX4eshbQ/YEWpfK3tF9CyDzr6N25YJmuJhLjytampiRaD3HIPetla
9EeekdjYqbQY1JUR1li9tbQLfrcxStH9xi5f2d4prlO4kwYabbFSBn08XP7pGw6F
cJ7So/LcSS4RBUPip7p7V3HnZhXPJuUzWk3RqMw7hfjFbKtxJbaluMU7UbFDhQxe
ym+WHefMkgr4oSbp87bjU9QoLmBObW75nouTQkAoneZt/pC+L1MfsO5wnMng4uZJ
yB7gGo6/wDYgxcTJ4ji9Srxpv/nLBBZEffBwBeogxubPQjgNYNxhYKgR6jPQ2KP0
77Wsdg/l4BqMh2tOmjuPU4kikp+5RbPLc2zmW2pYn9vWO0X4dp8fuowCUI9zNK5v
zxi+orNdiQqLQ8dhUyn6L77cGnipifARUgb8WlRVs58m3I3jWiTC77g/y45AZNBE
sg+QcV7djKioHnY31603/mVV/IiXU9+z4Oyfqanou22jY9X9Gas8Vbv1gLtju95C
4JMOV6OygtGTW+G7sCaOTi3+JnUjphQRNT2NtCWwHAh+ufNH+IT9FyP02B+Pd6Vo
G9afZ2YejrT7VQtbayDJwY5zaCa6tzgq2ZwyU4xi7zymX5U7ZIYQqEOrX4em6L01
xjcXZrvUJ6/oEJ9vlwTdiEs4QeywD6v/9u6pUoR1lprqrFaZDJ0j+VqVBJqx4buL
Aso7iG8K3DPEKQIKQyeRgvotHb4reGTh1SjrNohkXYU7HRkSJ5SBm7ZhSrqHiDRD
RWTzvV9LK11LnEBv8OD1nF36CU28g8x9dGdr3lr+sy+oLgpbHRiJ195gMSMCLTHT
7ggEIz96XMRiXOGcQKc6WTQCnIuNUjhz2UBF23uzztq7xAHndh28pwzVcy9m4cXa
SqMHafj64Yq5fddPJs0Ug9U5iPoNMHOoFNDqUL+fR1jDxLFThz/sivTi2FnSKOh9
rLN6z6ObtD5Oy5wQK+uynceWAu1w8QypvsI2AZNL/x42zJEj0ogi1AbwIPqx5+VT
wuJXw3A6dtck/RWlprmy5BhBIktcK2FagwvaUMxssYTL3fpiPXL48p5m1WJKKpLI
kyhlXFZTGN0vp2UMIdBA0aauuJTlsNWAnSqA+xfiL3Z2PUn/UwV79uZRCiyUvDL+
z7twsljH/YjWYjxSXXkXLT7iZfL5ttZtGqSolXq6SWarVcnm80nsj0xrTLELc58B
uLc7dPdzpn5EJZ9gMn8/NNuxr8R/og2aFCCmVHnxlXmbFp6F47E0hV+JG8TC0uGW
PVvhQo1dizwrRlD10SeyGldGJcToPhdaApzwkJuta8Kcp9h5DeldNnWAhPXTfrLa
GfY3T/9zGyF706YQUtyeVivw2+uRV9fCNy1/3zpK2bDl7RJGrLNGnd0yTcSQfGhT
D6tERNqJBDVFzwOfWKO1s6GszkAZAGY9S+nRDol/EvQ3DM5qFv2m1ZYXekjUlD/S
6pt2lIdWik5wU2MMY9p9T+JVptzt8Oe4TIv9y41qJAI66yxMgJi1jn2hP6YCGThN
GCXPLHesOvznKQLlBsTm6zinjhF3WqqeBTByZocCs2dlFOYpTVarqZPXhJsCBzmW
VhcNUbui00SzDa6oaHJX0/mgk7jkIYSRbHp4WqWUMRZDiixnvt+okXykoiBiAAjX
fIRFUea9Or8kzjOljGVqUDlqh0g8Oa4vLBVHRkPTS6bijfhAb9Nxp6feK2cprkvJ
VtbyU5PUF+XM8AZmnbgtWPv5t140M7xGfL3Dm+UbcBxJLNLDYDvz6g4P8SLv0lzp
I2NoqVyCAkftSHiv6EidbB0XeeT2wGm6ibQstOCOuO7/ACJ/1nSSv9wkOwKHyKQ7
EulpIGduyVDTpqewN53n23NR2ideDs4H/QBjitHjdcLDBQJ2J9bPClLNNSB6+NxY
MRjtK35HLRLZmxw4qAd24qcMitxVgCs+TpR9xLHA8GXv8WwoXLKV1tby+xaJZRLS
5EjDC2aMxCh+36R3K+bXGzoTDfVEQcYH+fJpuTo08Rq+lPNpY1fL1RUBblT30SxV
NmrQyGAAQjpQ5xNY986TQtf0fEyakF7C3hU8mD7Lh2WoQFf4g3xuuM2XzxrEbzCT
R+K9kSrUsM5y3/FKac4DWVLb235TQtgCyIRACbv7VFH+Z09rnF9e0NOA+Ne7QSfq
50W1CfYVdP/eVKwKWbtXLLTGoRrCoqpTTSs6/q3UdHPEOZSR0C+sCWJAbJ85QA9q
ndxtvPtu0DnOiGmtZOZ4Vd18SZPTvpNH0A1hr0o8YlWLqLEGbeLqHZCi50ee9AOK
zhpmr5EpOlr/ms4R3U0dgBmf20x/gy/4xislbzwAcNiQmHHiyh8WSbKwUGbtRUJl
fxKK5/WekavJQgG0rHjxbFRr+rdSIj9e8LMflrDijCC9kr285GaSJaCcnCT71ubQ
keQkESnLRemSF/xvqHG66YLOq0oKmXsjXHLMIOgJhez0X6I/SGNFlMWbNFqfpdKX
FUXHbrxPtHeSL2uoz1Vs0tYykMMZhxIxKSfHQytGR89b6gkRpUGTdRcIy1ejQ6Qz
QHMC7ZO5ExxlfJyAysHEsPZCAU432PQEcsKrJGcrjpIUl6tIEKQc9Lul5+cHVB48
RF8YzA+XT3CU89Ki39vgaVKzQjDokEnp0UuOpUlFg40PEMOWeQb14cV+2LuAXVn8
vO7HazkaxcfQAJiReaIwPg1hTZL7RlAXpquBBuGO7rVW6K7cnAIR4DAbQZbNPYS3
u6L0oU88evD1yf77ZT7IiFMEyWRR976PP22NPEBGyEYKvkfjAi5nZbFxQjWMkR2b
VwsV8v09sBbi/qNIDPIrn6ro/bRcl3W9miMDUARbRaKfYfB12yWGKtBZth1Ned3f
xcv2cVWz/JLYxqYZJQsHeM10o3SS3gSUbzX7BVVlMfSUaFx/xvH/UGPWyJ86BFMf
av8apFigDVcfVUreCBuZC/D8rATJ1ZDcsKqfGzIV+JGijDSVqbGGI4+rlXzJ6IlA
7Sxp8PCnRX+aOHWPr3/MDCHbQiEhDJLyDdixmdKMPiFmtwgUE4Mkl3HnwEqCeI4X
ASdENpo4nNCCHKGaSc6+r2TpJOp01Mj3lIxZvRpOT60CHj6up4UjXupS0EOdTzJo
QqXTA+YC+L8D2sZDhlmEmAm2VuR5AuY5ugiYb9ewPOpzSsISoRkK4HfXDJHkEVkb
L36UGnw1smN8vHJZF2bTfL53HGBy4VEtbc2ebWaT1leFVtKsYK7OrU+r8Bc+bggu
v0YxmKh2FxPHaa7Pv7mD/ciE5+vItH836dxDe+7oo+fjwZyiijL5b7oIyMyHM/u8
KB7pRWWFZ/harFw6xrTs/+HWITVefnetPmgVLveC4Eob9EZZR81A89c8YVEg6M9H
Vv0o1RBPOqiG1mmvS0vT+bbeQxMzxXMpGCeWFQPJ61ODHxuZWmSQKSf6qInae3Ug
HWkUdDuMo9I7xThpCu5KmodUJQfrv/m5IiNBLaxsnIASYCU1/ag29sgFlw/54cdn
KHViP/+xhuPYYlAqEnD7nBPrlB95r5auCr0hcxjqTuezI2dFnEohgFYpLggNB5rw
vWzT4+ohXnXO3k+7rl+wDZ/+2wlHF5AQKsdjVbFZBtV3wFCxQjRDheeD/8kQ6H1v
R6mRKOMCCIN2zfF0GbM7kBFWptUXebdhETqLSTn2we1suqOnh7LNO7ocr/pVvEwI
AoZTqocPpwvQ/FHUwB0EV/93COTBe+1AyLrvepVb/JHQ20W7utJ7VYelZdcx2iK7
IygmPULUqCoK74C8Fi92aiMaTCm9AoKDQSJHiRC9z8Pu8Y4RKfvHn/njv+NeScQM
aadTh5rO5Z/Cdw1nm5alIwtrKg/ZegSyxkYXH4RQh+/MkdYUA3cuGmBMtCuo2WGL
v516huU3kUW/Qq95TjmZRMUk2p5KnLBnHYIB94hr4hI3/avwYmvApP/iKZa9VeJX
MKYaJMgcSKEsrxTnAUNbb2wHVHSLVyeG8lJZPWhxxlvlSpjuFG9ELblQrjxmO9DL
UuZX1VI2QJGiDmkqrW9LT92ysJOSzBjT8BohmSCKYlNjHnWli8F2w4sIqlOiQCbQ
lrGi7ChatXeVa9pEnPcvqdohpiu+8c9DOnrvqhNpMVODxZZqOaVd95j9SXcPlyJQ
JmJ15t+RYmn7zf/0uXIRKygffpNrsxh7k6a98ulKim4MQeZM0GzZDO6rQJ7YascN
CEDAWwGPcebOOBZS73wLhdQTvN/BM+3/VbmX+sau19ECSfXCtyN6Z+FZ556ZxvPa
oHf0PKidXcFLs/kz+eG5kFQCQZVnPdufKwKkt9cvG+RBtP4Xi/BfJ2dqps4/3AQq
Ob95epFH6ufgfrkeham9TJqnAHpKYLE5mUH61TTsJbhgL3kXCszTw37tUx/ffW0e
Hr8qKp1H9HIVBJvp/FTeuCsq7eLga/n82P9qwZkCJBvPg37y0lzxchJhWHxmU6wB
kenDU/bTpU6rggoRWraKQmKW/FtV9gEUI7/WUpn7Vm7KmsxEQX7MVeKx7d/9Jpl6
x1KN/Mbmgb55ekWg2cIORINHo6G0yJW+ze4yXmHv4/ziok607YneK9Tye+4pKTEu
0OHSiZZEDBID0MSRzNqub5WyKauccccW33z9tdJCiuw4ryhCEne/+EPw4lBath33
MEir9HgMpmqXxK/v+MQQ55CvEauh3sBEHg9i666fLEv8mj6IggpX4zIJtZq5JgWM
OxxJMaKwWeCOLgoRgzYVhy2HB5xQcIu0s7eOFcmC8/ExazWwSwMFWklgrWaN6kmx
O/lz4QS8rRM6icH2RmUoku1GCbeRsftIpxZwqtZ7WfHd4Zwb3Tx/+WPUj4DZJHIC
zq9jymGH3D08DTkDzL+5fdlBWE/LxnEityiBhfYH/DHvJRWHgjudCQoWE9Ul2Qk7
6KZrsQ0RSpUXECtHn9Gyd1ACnkekk875vJQi/6xpyEyWgqsXZnZCGltmuDnYoolE
QFNzRDRrqUONj/KHb6cyDhkuyotGYMzxxR2waLqiiAnPIrZOgNtXjk3PE8zhTQ3Y
n0E6OQXt0hZ2ZCOEENRztpVS0MGEneQ1KyqMhKiZi5Fq6uCsVVBR6Wv6jL0nWfi5
aYUHv1EjI5xlgLjvhSjPVADZE0jOlBUyOv1ih7D4o9zQqmboxAVJSwWk791+48pL
xKRthOdG7dv/7PSZJSIzoVIO/thJaI0xiuL9pWhZXYkb1mfQvoH3VRl8I25LOlL+
GpWjnWWTWPF7vy5hlnHlkGkh8AU0JnydMmo+jqCGA5HVpN30TOM2/U0UhiJfoR2X
4TJNn8zIF09UQPlMYm89NjUswa7HV9MkPOLgGQVM25RDQfBelpoBu0v1oLzlgBo7
zb0pMlX9d+wohHZrHWGvWge3tJ+SgPSxGaEI+qbeuJKTHi9gk6gO24yLoDTon35z
4w94g9NdSKjDu+5FdSfC4Zws9Eyq96tOmExAwmCUTwTUV7PCM/Dzzy6eosetg5lb
HxkU2Hh0b2T/CJjtEcGu6BvUgEBxv0CcTYf6vZ6epet+ef3RabExOGF714+P4BPn
PbyGsu+FlEyyI3eJffJQXeRq8XVCn/OdAk6IhWwovx9dF2auS3evsWsX9iVQyszw
ZZQASW3CqZc9gvGXhGB5pNuonhX1jNOeeZBRodKWS1WRLdMCaOzhXJ3HvoBYIXiK
iX+8sJSGoq0Ffc0dV/4z5/y631bocS2qln+WnYh7ezfckyE1xnDXKLNsRRBUJ0F0
NuD0P8PvNqiqdnRw6Ww1mQOBrUGeFs6gM8rn4wAg/y7arxcCATd2SOBS7oZjVttG
ewkRsiBhu0XPy5xV/DaxoK+CqK1n8975wCgDncLsXTM7yON/vc9Pa0kgfoeOzbZ7
8U5lNbV3pMbSvKzLx5H7D1MMpDmZz+N4gPI8vLwRW8BN1nwgow2pykkcyJOvGWr5
5akTNuqLPzVjotz5wlGAw4fGmP9JYSEkXWuZjPHNnZkKRkNiBfyg4vwq1IYMCuMa
8sAYQ/WI2+TDy4M+26RUbxTFF1FvhngCwQbdTWvkJfbnI+C7y8Fyed16Hq3Y11bG
NB2QMHgYTz63hj5LxkQQ2AkTBdmcRiPFonT5DT7r0Q60YClLaV1gBbSMwOJy46xO
uX5Q7TV8BbxNYImMyYBZVuUxII4TwW8dhTMNXhvqN4YlS0ue7vZdWMYt+GqBMzPm
fTdNld6Zbuo8K5sYVt/0jiiCAnqBaEIgJ5TYVm71iHRrxHNrWDvV/+9x3qidl25g
2Vk5UkeqxvjxN0svaBbSuztsCZzfplkIxb23ZzkU72dzB4qJ5mF6zHI3bXvgcb1Z
9ZuDPEHaALxvdS8F6SewzOW4PvDGq3K4K3UXCBjCA8wUbJLHyIKM7kjlXUncAxhT
kzIYMFqeEmnubZNK7IGZlxORKvn1Qzjock8/8xR9htHdnSZSOiRAzT9rWGeK9vmf
UnegZ1MXtkSY2lKxulmnXQUyc0hxK14jUjh1mlKafaL50MRtri3UkksvvpqQbA0c
VV8z6GxhbxSA6Xi//y/7p/lOEEmlG3wGUh3E6zhjhNfdASVufRSNgS8Lrtu5Zmti
poijWmfYgetral8P4XgQizu2NRdy67ik/UGSE+h2dY5o5TXJ2XKIW4BwG90HwvyM
CDcnxF2Drm8TkKyE5C3zYjSAD+7J1S4jXrM/c1eWxRHtqraqHTWkoXEItJAyK1cX
2xlsZ15L0d6tan4PuclXIIPLTojIHT8Mxr2yS8YvAaS4VXxumsEHpXT8/DecXbVi
vrNCykIPcmx21n4drWZxvVw2KydC5fRqgKf4TYjEneXZ1bJSp1T6PjR3jN95iugd
VuNtCTLh9eGk0co8ldNf6xm+rV8tqBpRheC2bUKZFhKzWeZ12Ma4tm5ryIO+tZol
NFDXB1cIwHVSDA7qKtDZPG8sWTbWIDqVBDdjlNyrhjK4nTb/KvCm5P4IiWPWNHMy
IIRL6RpW1GleBzqhUJJx6hNDRxfkvJepiA1bXDlvzjzQ1ZoHh4v1AybB98L7WcEN
S4bL8Bx9fJy94d4ILjofEfm5u37uyvzpU8wesqH0ZiLBMDPEIMAwO3SHTqvlv2GQ
FfilQ5ptBOong7DLHvuKGmhK0a+OWU0nAZvYZcNe8Ez9Ioh2RCaznWGqIcJ3IsPt
sQoBvbdVXdGl8pNng61p7A+P7zwmbfmw2PO1gcWd4FYYs93p+7o5oKNgMSIXp6jD
0ag8Fi+SLtLv89wARn2v1V/vRxGPiRoHb3u8OGdixksu/pJ4rwbEaYzuciNQvhPG
qfP3bdNvDbPiCZ7BZnWoxCIdQj3CqYgQLseDvprMl8EON65pUBY++E283kBaJnlc
q4X5R4CWWQOKFfdGqYfd1m29OV+FJd2wtAb4KCjenx8C8u2V78PTeECvFUow7ZQ7
4kxducY/YuOQFM8ZVu48h2N9LCDzU2yfz06Oj923e9sbHqMhlYCkur0mX3yH87qk
dMwW7U3xxv8A6364QYnMtD7glrymDEfev1WMNyVL676M0Fnlm14jrn+s19iPTJGq
of8iRiXg49s1VsQP+gue41mZ49kKgYKBN+cHkBkwYum+879/6YUrs6BEvY5UmQRb
dyKrMo6ExdycQeIa7F4yvdkRWx+wrEN8mG92p2oL1SC+F91v5qMa5PZGxrY+ilwl
Sd6PwYp5pEya3QhfNZXGVbM4nn6nsTdmWGhTt0/7c6Q08GjkCDwZfRj/eTS9zrpc
gtxrzy4KXfaiHpAca4sumL5jocxi8t/XYvJDPRU14VYc4tuldj/UqRNU0RMc4Jnw
tNBWddw1Ab/izUZEVaUHf4TTU8+vlrfvUtn9qQTtQHNCkGl4Uc22qBawd2Hf8pHl
iZbhaXVy/sKnH5eq97x7z4/qYzaHyi+kWg37KKmnkDpTBTo07YMwrhBh/TCYgwEi
exVGdLwro3bFLILJeSSB+irAX7mrgqYJkjt69i8NeP1LV0+MEhVWyy2latfBx50+
xmSBFnVewSExc/eF79/f1DhKH/7E0YcuN52XCFy5oj/w7qRIuAMXYwn9srmKOGN8
ay6J2S+4g5q8OLBvVlh16EEwNnMKlEC8SRVeMTUxfxbL0MI/0HoLVB4EPZtyId2a
C0OADybvNdPbZqZVZGVCf6NZ9S+RTfC/bjiYg0Sae2Tzai0dzvS5cxSLSvrmAry9
k/PVkrIfcKx+VuAkjNNLYqjJeKbxftijBMGn5ZtrWqZ2xMj2S3y+tZxG/UYglAOM
kglwH1QzJVon1Fv5FXJIHWowqJKPboNmGqTyn67oS1sM9v6IISqaaEZdWkEjDAzr
pKXuricY5vyNN0bjJSoAIGHEN59Om2RfQSfn2iBXKic94Jol7Lle+/eWP5kRjSTY
JSMIqpxmaq3TpNUYESLemPy+KX+kwNLAzqAsWGqJUTnpX5JFwv/4HTRnzCLfxrVL
WfnxmBEPfWHSP0FFjOLDlSH0El2CFNUo1RpoqXUaORxUVlOoLEOZN6sRzPkjZToL
LXVIwql7EZvBhsvf7UPVUgvJW5hX96kNx5PyiCCuxoBYC+n6jrC68uYh1Uuo4R1K
bWnYed29ZyA+YHclMp9+THQJe6TSF8F3kmQgMl81Lz7B1Sw8PCK8GVJGu0EdMhT+
XpYCtyz3Utuy7cYbjGcGSCdMTiz6p1E98KSrFjDOyhMkeCZk0I+ikxchSMiwSZ/K
P8hc5VL5Q5xPmrzuAYWYzROiq5o6j5872KgsMysOwU7HDwYKB72jJhD3h3xFsuQD
98nRSTMlvfkfdf1zF7vW3+GofAelD/f8o00b/qgL2GB3X+Il0cng/JBsxRSRZtiu
5qiUoa+EszTMEmWXkVa3B1T4f8QpaVSXRp0w72EE/8PXPS9bJhCajHNUpdcLuEP3
HxQOxper88Cd+h9noLcRBk71PWKT6XmLaGuDDiyVhqMQp113YJR4WFUJkSrifSvB
uJ4hscqTi287slqzxC+GrB4lzQtqKnwI+5us8fPf3ExC0drxDZOXltkBr7H5oo0I
rvdJqJcNQLKZpC1ZknRk5yWhXMMeotIBY7w+GoTkx045OmiJOFku/1YYWdETFN6D
xOsvEior7MWfpEWyywXLfUQhTPvCb3YUUPLPy4LrT5/D+GbbBOAwd9SBzYPDYwbg
CBZrRxkrDcWR/zgPu7cWV2eEj+My76zPH8Bwpd4ScKk/bqQUm/WPuzBPJN0HHSTC
qWAkPAmYTXYb2miO47Wqvl5dxc+4N3kIjwYuxbpIbkcFdlHX1f3ibhoAlhrpyJ5+
GiUtq1YXloKcm5AI9rDl1vPCYxX1YCnDHn0nd3VeTCfdDW01anF1OIK8bSjwMBhl
d36eoqxKqefqnNzemmjVRKlea/F2Zra82szBMzHXYepk2g5uSingz8RgRjwVjL1E
Fa7uw/BbzVeqshMI32V4nnfQmSuq/mgvZFdXUOpoAQC5Rtha5kXezOJX9EARWREB
DwA5ALoZ7Q1eeDkOv7UhrMmbDFSxFmCViq6/DuRvv+XVGFFv64124hkM7lWOwyXk
/7NIKHHApsyvglV7ATHDuWS0jiPbip0/0wkp9d0UCDl1brYJ4Y97DulADiV68voT
Y0H707vI6M+cNUOfTIt9udxy28kVuw5eZGKI6KODMElfdnmHmByfin+pKpp53cXY
BL8PC+f6v65+jqtza+avMLfbvELwze2tKP7XYND6S1zeEfrJnJMbObBKY2jwNJkk
r4Bqw+3Ip4osvmaNLnyIZdyulWIsQArINTbvUtSkvuACw9k6RSMJ4INbnglG+JwY
nwybtI9lCs9YBd+p38oypO9MLTgMFSg0XubpKKDFFOoSInGpldtAY+OVB4zBG7Vj
Gh/KgUkHGJaS5Axf6SkGJSLQNkpYltJCMRpRIdXDxCTfrSeyThhKQDYrrUU8+Vnj
6Ou2CCGqRYppS9YSs0wRQ9kj8dSBoGfutqPl6BC8rx2oSTYV56AwK0gP6oWeE1zC
Alaa9E767tEiyCgMwEeYeHGdRISw03D+4onVchutmg4MFsGPrDo5F8WmlN8dvplY
M00NnJnw9up+RxGgz3ywcmSV68YA6CIdHHmFmNwYYkZ4M2G97gCO8G56blijmMoL
zul36PCi1m8BM9rpnU6y9fMxUTBe4xUvT84F/HSBqr72DHeEADA2lVgkpSr8jr63
X/4ui9GeA9ykAQXzAs4MOJIYHQPk5cA9lcoQwrhzLwDTwP3mniV0y1iJx7QA+iI3
hlvN81RGjkWPDhFu7Nl8EScGENFNlsP9KtoaXXzhDa9+OzCBh+qzL6/aPD+rNwkx
sHAdmg7+NUGPg2T2IjaCingzn4o9syVh78fjgG7wGW0x3bo80/S5Cr4IFfGAs+o/
rALPSdg1efkmtxlpWj3RWpVn8c3Fa4QLex4Vz80bHCoxHM8CsnHeyAgruY+G0ryH
yMB3tW1YEZ46J4bm1t9vKYQ41l4gccVcGg53ac8b7W7TLdjPFypgSJ356EqG1rRN
4wYgczjbZqqgTtnX3MygHPEhHWk0WjMSf+CwkgTO9LL7jCP0X7jc48yonwGB0Kof
L77U8q6r2JfHHsui2+OGAojdo7sOSbB3ehdJuXj7dZ3ERp9RKZa3DJPEjU1wPNUX
rQu69cuy76lOBAjIJJ1OPOmoW1yVJVwRL4A/8SEwvtEmkPZBsf2mn+9yuP+4d0nH
8e7XuVeBobiAh160Ytg4GTowlQTj1aIm2R2EK/icoQnmyrq8eifkjTwZaOhhuRT+
++IK4uSQofQ4qOu7WgFJvykcBE/q9tORclP1MIssd8JZKo4x/cp+X2NiuCzmTB+H
s/959rkwxzXvzCIapx9l2UllykrSi3sNP6zQw+hWBB7rd3j1cngV0Xv1W0fIZYMv
6inmNiZZmaa4LNEtdoTYBG1ZePq9aAqczf3iu5TA6JfKK11Y9TOtwtkuMvQzgXpt
7qsdMtE25xY+wydhtgXdJ2tr1S+vcBn+PL0WURLrHoB2HpZNUETyJYfFAbYwvMlx
TagZHLbzOR62Y9TTX3jlAkCj5d/icVKsaqv2VmkzpifCq8UDwbK+ymNb13CfRLJZ
3jxn/GWMRlVyvSy1XcNoUUOz4bMLioicwiLuiNycE3FklWctMBPOA67IepeApeGe
HK3+edkJ+HDREVTIxLI4II8zTNH9x5BNNn55OQ3s1Kf+ZLQ5h4aOocDlSh6Mfhs4
1auRZJusyr1mBFfPM2v8ePkJU9bNZT6i22gl02bt2jPOQliQ2TzzJBDSTdvtPNaL
MbSSSvvP2gZt/lOcQfW25OBcoFWbYFVnPrzUod3vMLhu+hHgmtno0n1+pbOZTM4C
EZhHGcS5t3vqdEntNJfy80PMvYW3rJyYf+7FyOiBiG7ITaTbCUon/z9KDHWftjFz
4TCv2odtYfkM0d9XfBaNTYV2hjieAmkYeIRu6FmmIH1VmGW8L4n35IMZDd7M+VC2
WpmVXwwx94XBgmkM9Nnq8VMh2N0Np+2TCcxopvqqOoOXeqpRP6IDTnFQHPOMaBtU
WFYx+wRL7+7u+oLgkNBPtgAraDE+HyW8Xw9k/YCWzq0v17TzmMuxgOSTU4skZwwX
TbdQyxUM8vkC5v3pzhTEAEbLBSLqtKUPOxsELkGCjB24b0au6QeGwoIS3BwpjVHG
h65TYs112amxqQUQhr8DqPZhwCTK/9sfMOueiCk15dXV3XePzjdzMSrWHr35vQGk
6oKBrTp3TicHpRUseP7+8EPZ2AB5W0AbR/aGuxtEMSUUvuDGJoJswpfC2G5p1vbP
3ezpdmP5bsP1WXVEf2amSe8xvoQIEGbHgv18bKeOyhEtkqQzfb/R4KfEMDejgezD
h2LeU6C5rrRAZdnFfc1zhIvUi8/DtSylKhPNDyGKUotcjNIPV4NWn5uow6DYPIqX
9uP6VxMjAoW3l00GFqTSBltSfi1BDSx2lg5hBbqnpmWx+8KSlRXpC9L1AGl33zrP
7WeGLQFvcntwcZr5hOMbW5S6XVlGZ9O432zPutcRKnWYaDQs0ZCxMVFsyI0Gk3vI
7KrWOloVIFH1PtsvM7npP7v7vHMXpoVzxfag4Diwdta9nY0PjHCsDz1APJI4Yulp
DgrqXdiNmPlz2nZlCMFDNbTFo8ns+FRjSBBrJyDn6wcr3e9RoDaEChGx8HKoP/yO
fgxkz0aVrnbNrpZhIZV3o91WJEaNQEHkQQE7ouzdD4rh4e6aCwxEYGjdCwqF5Zd+
gcHLRLEBb4DMhy3F0imjpZgWmOCfYy7Jhjv9c8l9LqzQIT0NV32PhwKYgGEPeG5P
1DLPLbu0PpRNe8YU8EZZmhlXqfaK8ocltfgVTXXAL++2dRAPhd0Deh3F4D84RCOg
2Rr+87scoyvV3FZkSkbnc6LhOfx9up0B+KCPx0UTUvhin7o8XqJ2NjGHA4ADlduc
aMQrRN4T4tplmRG7ybIJ5vbza6y/swz14ASs4v6efRzU3yriHeLfBrmPc7ooReX9
lViFcoX7pX+zita65yUqmveiCZh1SvpVFGHxAFlUColOX31+ty8FeDWQKWWJTsTM
Dq5XI/B+UEAf5iv9o8d0YzJ8q0QA0Ktv5ATPI784CsrYyWZxOEjrTECq4dHF2jfg
D7B+tEooniw0NQRxdx4YrXjZ0+QzOsTsFUYD1GL62+uQedRUKAV2J1bMEc+I90VC
fgSMC2EJqupwiZOSEtxgC4mgh8jbTzbaHy1FlbZ33Gk80zCHSxqg/OiHmSLRrqke
WA6epUtZk+f437knYljKqzxomzscKzICXxRx29KuAszY1/CU1ZLH2nAFk74M3xTz
oOPOOi+VVUW3ou8PU64H1hu6o0dr6uTvPBlK2rfPg0r6SpFlq+Ku45BP6YE6GaTU
rvqUarfq75CvLAdq+JQ8+V8vIY2kufBqE6Nir1PuX+gKpB3xVfT1wqkMnZBGwn5Z
M9zcpeLHD25rPIEnCslxNTHVDCtjqfsxS7ay5WAwVuuz8HQluWnQX6GxeztKA4gN
H0wvKVvHXi1ifDied+EyFXP0zHo+coznegJpYsex5H2lvo1MHQp8UPt7szI4ZYoy
Q7FnSe+W9g+32U18GerN9JlYex/SQt/2j9i+qgCN2bd95BayIQAehZe5sEXCiM0f
9mTEmiBDs/EHX3n416hHEEArYlYRfOaEuJXVgrpoWLB4QkqEyiBR1k/45A0VKrRk
ug6iSzFii5Zei0ZhoL/1DDJUwGzu46bIU7llWobfHH4R/h8KbqHKGPfdWdLYr7ti
+MYRWBnezNp9xyjzkqhtjLuQsRacGS9nDmP2VqaOg2kRsZ4kH3h37J5LS6DqPKBh
g0iCSrt4xtn2eU+MIdOgzRURK6XSf/xcn0OEu2RErpXxBR4dMBfF66CmxLPxzBUE
U/K4oExtRrHOYOCUbDOw7bg9r3tzm2FnRL9hhz133TImo2iF5TIAjbGWxOtnwLK+
A9PWyoFCsFjNU5l9+FiNYyManSveIjp47HNI4gcWVKcnEhCvJgCwafv3ald6FBdM
ytX2StA1HgCVTWQRW7H6MOfrJntjxScX83gNGz43qcddy29Lq9qmBUcStNajh7e1
1BaFGUKXzoQQKlVeKpkb6ssKFakqqXmOFsEdECsLZZZoCkfR/+ASqFSLzoja8ey0
Ang1+Odq3HZHNUHRp91FyWvbnzfu5Ji9I+xOF/CB88uQxJzgHTEFS6z5PMQHkvP/
KpuI0HTZM/FwGYJed1LL/8HMzVrHmyq6v7MEBQqj9ghE62TvZZ09pf6elx180gQv
Jmq9eXxTXYtRRafWV/az1Tlv2+iQ86pKctS7RbXS2vWjy3uF/PsseH7LObbtPsHj
uewR2x2T8Wf5kIdeVoQ0qhlIcL596iyvVafJaKZrMLgy2EEx9p0MejFfD/DWlKzd
QNuPA0k5+evbwMYstvDMqno8lS9iyxzZ/aoOxYI+gKWzikJGn4UctkIHvVRLAcu2
tegeevL1iW8jNHg8vUQ6VYHwXZpaN/bpiNPyExkVph76Rvf6Rfdf/vT7b7/vg3v+
84t01sbj1Dl4HY7FM5AoClgwhH3BocTyBzlE7THavtUiUQ84VG5WbNwy9E1pYINc
8an8W/oOCfyt0/ip7BHpgyoYqFPWJ6/QZWrmMqnqMbn13Iaw1Ha3ZAOIYv4NtQc5
vmDDQIs9cc04eys3xup4PDu0Q5AOzZhq60xEHNXXueNKNNNP6ns5RzhOjsn9I1ZT
Z74G/QfZHwF2LN6iS7p+nTk+PKPNdOs8uQ1LBL0LTN+O4e96XH/nhClvIjDgGD/n
GRec4+KXW65eSUlQkLb8cSKt5nrmWiZVc8KnuDhf4Ab4vHGo7PQJDgtkXmDMEz57
R4l92/k+YBmyRAuz1dEbj0ih91xGUvy4bVs5WDjKr7AXNvStrtHLRUP5dedHuC6w
cO2w/SCA+JFmGlSITBJTpDMBA2Oc+j4HZFzM5Mq5b0mahxu39qUpe7TMT7+W1AhI
AFTj2hc/XtGtIDjsjnP3f/eTs5p+4cSsaGepuKSPdqddZ5OpdFiUJ1V8aT2iXZE2
2Ems3w/gnbZGsfxrodSj+F1ObICMe5t0sSiV1GlYk7rQlGBwcYFewpP/GIfejhT2
nEn2WbAg3u/hledjwH3IHYv47DjCpullu/8DpzUMdh3ocMwPayRcNXxUzE2nqVXn
xOkEcghTLmsaLoFUHOzJyMMWNViWIzq/5oocW/9h7nyGfZESUdsIsM7QA8zMh+8i
g+/4yBqG6WnXYgSKZ19k++tEQ6vwA/1uxGwjIxsGkJzDhI6p8StBShWVozbaAvIE
du/bak9TI4SL+MSNIZtd08ZBYWcjezy4Q/3Zr2feE/iE3KH/k7pyJ05pByqr5Jdt
qKVz/3wOOGnmfuG8IEHMI8oOZf+ardPsvulgFdy+X+CyOFBiHaQNBRCyy10UpMWj
DlO8pB6J7lDpn+UWWrX/aUZ2pzbHLDvOKIZlfvElaM8QMVULOTQif1u3gUEeeOCN
pQeWuIyUvMl73EHcs5phniZSXwZKU1A2jY1g48huYK8W0UuU/f5SDgnBWjk3ACaI
Yi0dRIery+kSZoWl/ObaxVgBHTrv+jVi7X1dxehKxQNJdwnPmFpgkGA9cj9Z8DlL
z2oaLZIu4JGq/j2m3SwWPhokITSddMUn0ic7o89QGSMFzXEdws+54X25tm4f9hOT
yDY5G+llptrAHxiPbJZmU69JK1L7uUA6veBxZ1/etrUJULCQk3z1/NC7NF9PxLdJ
XvBB9W0RXu9C1DAYWpb2x1h+B21akAbi+wvQRl12d3LzmdiFlaCj51IECrwX2GUe
S7V7Le9n6RmSPM15OpdTQD0E9X//HedI2vFmOix2tQbq4/ic9ooTC0FITeismBaS
dMK8q09RyRRKqg33Qkj1D/xY1RrrUvtkp6dbm1pCGY0KAkaqaKearwycBEvoaUu2
tY95zxJLtUCbK3qP5wuKSlgruKMPLQY1ej2Y9Gtc5RXH9GsLpwxbO561MVUPlnit
FLNKszlcg02d+5NR+gEjJSFNWUFMbaFBx2iQ/EBJuHXlg6WfUJVM46wxOQfZOhn7
jUXP0Njr8doVyEPuS7vjWgkFzDALMWS1vU3zB7UW05lXyUBDisdxCJpofQmo3Y3c
Lqg1WahhpvwwvNE3vC9tGFnCk827pKrJE6hI2wqSQmlL7lWwSTgnLWNfADJ+UyD/
wZVnWAuTOsBJPEKh2vGWqxRqe0pHIaFzkpn63CxtPviCJ8us1M3MgsEXMZjya8ty
+IrVpe7OjrWBjRWkRMKV00jCMsNsCG2v7veaPjP0M/9x8uNkcKNEE5V1n4ZIw6KY
A3EnddyAKxifUTspAKk3wb7csQzVEFV7NWaUGeLldZqa5t0DWMhiQEBhcjOhpAVx
iKHXN65ul0m24NKuIYS85vuC1AK+YRAqxhvdMQ39A3GgNTmYIrdb/iCEX28M8Eht
H4nDCYQrOMK/Iis5oyKa08veL0HFTvjfppLkH56gGa+JYK8TDdBkrRA1vFQqD/ee
W5rvdSWy9HIG4s2mVQsSJChNhwRgzSJL8a3HIYwgWWixo9qccuAGJJW+tJq+FrFf
d6opPrO3zpMSs6nPxmY8pdwLwJ5Cgz2B/TX6a1AR6H2qgkvzBji8JprSbcsXbspk
z4Tq/JFeK6dL5ZjiDWEYdUfWceuNNeXLFA6mvsOI+3RJ6vXdSakAx5awy8Ncfi2j
DtA4BEElf5CrgpVg4nWJRwG3mYq78qsSjogK1BDvbxKMYz9/qW9Jr8Lu4gF7N+uw
eYh/sm39jr/zuihbSYu6P4cgMlTxKCBrHLq4eZcfg3LDvHoe0EnH6XRzlRARIN1D
Ldhvcowla4cNlSTrZjNSbo2iNSSguRoQjaZu10hFmNLPzAogtw3T6mnwWoO4btPz
IOpJU1yLHJ6Po3dl0ZRj7xctaI9GK20P1yVkx6xoce/+0PlNvIFkmGtw0RMo2BPj
PII1nEGw9JgORkGTpi0f/FjWWcsPx+b0xrlufmgby7zAcB22qSqOtQSprZaB3hgy
jfkpb+HuKlWplg6/mgH9Fk1hdsBcho1x715if6o6pb+FM/dFqWukr+D1KOnnaQrG
Y+KlNTv8Wml6Kbg/LvywF2QcufCZeXCZaxYXN7YkmiizJCHsJOaCuMtLUaMcYo9T
VV1fyFgncPS0jN3puv5fMPvSGMgF+kAkK7naAQcM+9eZC/21xALjjbZY5v+N/K44
PVGE8mtLyn6mWbvWXF1RVYpzckxC78DEmVx4fBnZ8QU5MsPRCfoVKxfAAXqqo/OQ
Wbr5RUOh5+VQmYsSdvqRQI9RW/Gi85oz9mPWM2UvEWHkasjgL00tM53I+cNcsR/5
xK+EGxLUvgc/KSMxDkuBiMfbxtcO0qNwuZN68dYA+LxAu1KAfh4vSYzPLMqLpBtS
DRHEUqo7o+PI+zLtTNyoFtXDBvm3W9tcZhz22U+9+7/Um2XYwjAwGctAOYUBy88B
BV8NlbHYqFXrS0AlMF8P1iEonrC5oCF5M9oiiLnjcZNdq5WVsjPXQewh4XDWNX1z
N8Ezs9D6EXNF7lM+r5LjahycjSbnIbdQE8MSWs+L5eaKw+Dz1aRzPxXEpHj47mBB
lvDd697KnTcvzewe4zzvIN5qpgIAvDONnbD0ObZMyy/TPFNHCc8Ef4YXHNptawHe
tljhtjfHET28h/VAH7wq+KfddXMS5fPDIrMm7utFErgSDopHoCuDWxhp75xxwCE9
ejoi8RiJzQfqR6xG+tum53/c8Wl0qVw0MKA4SuJkZry0HFzpn60VA2tbC0Js1/jP
9rz6RCK6oRg0m6PD9iZC52eB5xep0PcKWq9f72vF4FaGVE8u35zavMNzGVuMUGKh
F9PWd9H9sm2keYQsMVc0o9d7j32ByVTv+N/SoVIJfj7x2mcLYbM0wxWA6EtE/Haf
F1pFdF+IuTUWki76GhA03IFdp7gd3HvOv9o8DEe1RSVoR4NrAjTOm2apRdpAqYHw
ti3E/76eSQqH2Wbt1DmoJVhzBc3ROWrEzvXua1RZq0wpVm4yK7DBHQk3Eo67K4IA
HaSR1py1e6TKxa1+pX8tvwu9Ub4SsMhAuq8Aa1LMR5Lf1w4/hdnR4BDbYH8YBoGh
k6TjqqMXJOeFy7k6FE/p72XAkstK1LSawNOoscCl34h94/WVUrLGsxwrmUhMRjGy
AUVnAbQYzjtt+BnB9hxyywbiaO4R/P2DhJkKD1FP9sBzGjLsxsivZu4Jb3iSTD8H
xuBtGagfq5ph0PspkMHfcKHh6HdkFcqBNAjszytpLTYUJmSJNGgDuU7LUnjzVslk
GtCpiGa/R8Uis93kTDUxFlGF8+61PrSxI+hEDoODU5vVehRXfB4+H7Kb46krl+Vw
WwxslLJAnr2vq2OjooLBHYcp8RjTuXubIpZTFSGca+6oQHlqgO9PLQSEi86PgBhB
4LqF3YOeYZwk/RkA95tvoFwzNry1LQXHXiRdUHOrQF9tUDLfpN2LJsCeoZs+bNsI
85pNsK87ptVqzhwwGvk8RyWgadmydjFSwuc2SpdrlvP9yu1odP0LlD6kira2pYEe
tQY85WMedhC5935rYbS9KlDe1275MXodO5MRqEdP3a7HMO/vlugIm+vCgY9MeFbJ
A+PiaRHbau2Tzwfe+TP41ZjR0xyzjXk76Y0vhz3U1JkG8ZjlS7ncifQ/KXvBNpls
/7oQtWz4PPzYUxKAh9z3/n14Sk16+OSjwXVLEc3JmcDvLwG2EvqQl8mIBy7LQI+l
acBW09cyAphQn9FK9zqRWkc7c/xt8xjwodkMWrywKudNSB99ExkzvDvRMOvHjayt
DeASyFhQOiDe68GklbX6xzP2OQ6pboiCZACX+VyqXetB+Q7Eq1ZbaoDEvUGWGI5+
Cb8zgklpzqgUGrHYpeTljZLdglihUKAEOxq+ewLN9fSq42m1oIZjjlR7eBZm89oQ
G0UzG2ju5hzt7zMunIWVHOvZ+pKyUt99sQYI3FmLGFSLY/CsVMPP4XfKGX1ajMmR
DsP2Tz59NKDSqFkummDm5EU6xADSHbxyQJYBxv0IzyAHvD7gE51zGNdvArV0OBqm
mTUZG79s4oXelXTF5rYuxPdyKNC7AeWgRPkfGdhwTgUqgJRZNiAYQ+EmFlEY/DZx
tSYEaTNGKDOYH/P4EjdmOZ0vkarYz2o+tNn19tDOTD4GhsJe0ttHQwPCTi7jmMIW
ZEQ/+FWXC/HtFd+z2dMtojAZwfNRevpz6nf5DSuvgw2sXU9vv4JTT77uRIuI6cBJ
hL8xkdZyiW+EuMvfSeR1aBY4zHCCVsEJBhTMyT1BhHTpnkXG6iaJxdPV25W8unKT
D7/vRkph6/lODvS61PvN/Vvptb0x5F6u4Q5uAZi66q5tKKrw5+Y7TPQJ8nWqXO2U
TB4FLhChxNwQarGzToXgF9EDWdXlRsHkBRV3d9OMnjafoKKeRzVkrdzQwUuJXLOn
Fn10GCfVRLE6s6isK96H8ihQfp1HouogI+zUgGI35BsXXAI00bx+sA0XV6RIRMNF
/TRBnWs2PHHDVar5lQfbQ5ScbPLWXQb9SmgxKlmtAhkYx9fE3HAnN/WeghCLnOtP
+r+iFxZC2EAzzL2T0ErBnq9fAyuN0AEyErbwr8yruw3wa8b3JdCvrDEaHCbmszVg
kmrNhdC1rsZLqp3Km/RZx3rqU6KhA4FvTNW1rz+7Xe6i+CIFPUMs7t0fDToop7Iz
dlIBStJz2YdQQRQF2r0A+b8p9ZXCR4fxE8cqXZDpGVCceWvI9BltfoZFDl+DBgg5
WDy58oKhvPjxZiwn5lJmLDpmjon7yxjtW8oSAN2TaFTXgdl2B98bJ6T8wIGyiZsV
fx5pdPFbPtuVI3k6eG51BfbBMlF20VCApZ/ExcG3oaheLc4V1/17SqQziVG70MxC
mvbOiUeX/22HsIqRXxBN9vqGA30z9Xv7aJvOMlfmOJZ/cDrH9EOFFh/JJPSQMV74
qomM2vC7c+rJsMgXtO/dKmeX9zUFt/BHgc/K0ezJlnnkrmpcty2Ws/xmE6DfrUG0
eYDbthjBN4eQUylvQSFvOHxrS4kQFFBZH069udov5SMwboiTVa7D8YKe08gOASGH
b9Jxa8ak81LN+UqEE+H3qB0oI9+fa7ehF7ghvI7gCe9RvKdS1mIubvmi/Xln3Hri
6rJeW4IxOa/EiQF8cSLTTL/ENfej7Iotne8n2+BlTpfw2HlgJedGWEE7ghA8vDPq
KQZzENp87Cg+mh2GOrF9n6aWcdd++PxTIipDSS/dKSsoYrBJdzKTIbStTrhwVaOH
FAIsSkeA8ZjmzI2kTS369hFB+O6N6tkdvMuxY17LFd3oNEZ2LdaGNEXIzZ6lNRbM
wCgsSVnB+XveV7KGe2i1gG56v8gzMl4CKjV4/YTNAq8SPpAaqAbhPC8rSTLYD0xN
Y42IdTj82BktAnZp6yXZF9mC1Vr2aZHFhI4dNnj6j0L87Gq0IOt/iaIYnBlEcAQD
4RQJ96NsgicNkTvBwTgqEirFLLCbsjBYY8pcKqeoE2iO+CWwKDERiKI/nr5lSqb/
y+nBH9QNdxXUDa8GjeFS+OHp25A2M08ocysaBbr3la01xGh475VyksSGg0aZByUe
Vw2pVHtR1r7+CNEo9IxnAEhHf4LrdVmLJVJkt1oRMxB2mn+d+jkkQQ2w3eEBB8/J
XNR5poiDr0JEJzqd5Nx69flSgt6Oiu1EbYdHtLhc4yKNVbyFhSnn9jibz60a6XNC
WhkjpyFDXTjHZe+wg9ppmYwhoVi8QqmUUGmsRGJvx/9D/FL4WAg3Jysc9aLIi7h2
hOJxBbUIwm/3do6Zp9ElIS1cBTuBXqiUluCUxKwO+o1yguZEtjMrWf1CZvlJMRDJ
5lAMSD6Thciy6hB9yQ0LF+cxXXBESLqtpPhLPcphO6Pqho48Yst7fJaZ7mUouyPH
Q+cqRwz/YmhjgmKGeJzxCDDaGBy2iTgX+dV7IyXu+YuKQiz6r+8ItiMpNuTCOJMl
osCz4wdKGR16i/YFqgUJtGua1L0ejqK1MdewpojCfcJpdimZLUezjdwsIMDbvRQF
wQerosYavkiOoV/32sgN+CoHmn6M97OctOmxQWjl6SIJ1b61kMYilpQ3K/Zeqz98
UlMWAZe2m98d9chD0U3JSClWVSKs3CWUDy1+x5Bg00Whd4QSsGmAw6Ny/py6Fyq5
yqakXBLU40MFbTnTBDePmZvoI5RRffnJG9M3tn+RaqLTvieRkUn8eQ53QyHM/IQi
b6a+TLc32/a5qBtts8c+uIHvNnqy3H/FLojpikVSsDFzGUIEojgMlwtPgje/vDRu
svrVcipaFF7fZFPMVMeS/D2Cc9zziaZMOH9vxiID5aposP4RIfgBKLeab8HDzwLU
HgWgJ2ceGsw+3GO2Ijdig+6GeB5o1L8ee2f8qQizaqxSV18o7FRM0IsBMuKoJh3R
Ys0ZkCfYxuKsnKqrytjyoI3KFUyfQT2rx59/SpZAt0oYxx25oehT61kXKDmjB9E9
bzzVuqyj/+uM9U1+bUj5LrehDOEjm/RQdbWRe/8c6+6jz5Re6jLL5krJfQ4qn+NP
MsbnMQ+D+ijBysIDMMrDIVZ9pZ16UQ6vetrmPAM/L1/8f1HhVp09M+1ZbpTUdpGY
wUayiuYOeObyW6SPMFbnjB9s9IYJrCgnzbERnpWanhCGJxwGy0AbsSQHuYkXxqvK
Q9EKMwWNe5LnRhzj3NKwVsfMfEdm927xTk9vHjfftnuwP4mO30sEiDPpGIp40qHm
ZTZtkBfdyPUdo1TWoIcTg5cvx1TQOg5YHKrefUKarhgM3/VjiZDPv7R1Y18iKT+l
A7n/TRjtv8hP8Fl+IYNcUX6vUbqJsoquwwpw58NqDCqdC/vcIsiqzFN692yJ7N4v
kmgPcKSnGx+ZtzFak0RqZO026EusEUXdeT8EqAvQfT9vy/P+9vuVNKhKR5Szp6Qw
GsW9A+y8ISFvkFO0S0wbtgFKZaWkq4pEVyt6sagvKGdWvAzW0lv8wsIJ1SeNj4xi
BqH4aCpAUfkgL0hiBO/zP9KboQp5MJ5SZwzWKl450PHOgU/lkaxHbD7fAbWBRXWU
xeG5iMUD4SSBUPewJqvLal0OjXPq1R+1axzf+ZerkZIypjuurdCw3J3+k+vgXLoa
X8UYDtpExpGkfWrPzzOPyRb5w6YYBNexkm3G7YsKwSGiQo5SktPYEvBOp5fNyw0Z
q6E1ahb+l1kuIoMsKrSpRABcVeQcvYK39iJvfbCLnXQ/sjL9geCr8flMJ2fFHrpt
uum13nndomfAxrR3Z7oowUTPG7RVqGXvyxSyCMT4oOrFRfN+dI6ubeKMOIwu14YS
toOO9xBX5j/uXqzBx2AfRzu85WKtPBvW2PpivrSvglRlQRpES2XUHDh0/E74ztzH
DZztDFJDKOPN+Wg6fBUE8DxHj8VpToBcPU/SMdhi3EF1ojR5wr/LBmPOPx7ePWFM
0etmj/qRrKI9Aj4djt11TdIIQEIneSCspHOv8tzkgazgCSca3otxlZ982ZxoSeOA
4J6/FeGhoPK+B6kANoW4SNQhwC5fxpOgd1cvBvqhQA3Y3IQAW5hEwgE8cIXUSBii
uMS+z0tILG264zrYHrKhzZefdcshznGfh0XKo+jLnPCQYs1apes2q5Uw8V1XRlSB
sYLlO1w0eAl2+7rwOYjWtJbUunFtGemdLjBsbnzDHVqRbqCfMPHyh9rucUblO7hf
l/ncPwuKwKvTTM2hh/K81eAb6olp6RF8d5zqho+ALJ2M3Nz8E5Uw8zlAAmKiX9G2
6k+ogiEJvh7vcsF+JXaPVXOhKreKq4Pl0buLTPqYp996sXAiYW7oQJ9YzGUCone0
5dbZIH7BixH6lOcPfHwdBSRmLIn335lTIzZ6zpUUPwbfmQas9HDBCre2LnKPmc2U
pE0tXWjnoRiR3AHT5QnefjytinIolYYpJKt6IwKlwxTsHePIGMMtfprojJM5Nn8N
enIXYHpI4HJaowwMU8eOPB8HLABtywdS2viEgZgtHClrFX0MzmgCgJo2VB1uj32s
HGtd156FhyCfttE4TXjGE7OmoWOXN2bKMZdb1PXb9E/Rl+TMCVBkQGO1nOqawIhN
0yVO9ORhS/8MZWgP4fZr11ddtkTjzzX/gRH9AnEjSQPBdjfFjj1J798OTw9i1zry
3nprBWrhK7iLBEA6KIR8HpJ+QCrfoSwRFu3EmZCe/05t6mkSHALgsJIjYM25/z6C
Be2wGIeDT61PSE9veKPVlQza2B0kegoKJXrPG/RliINu2W72eGlH6MQmSjhGGi87
xxGEiRHSB/RMA52KPs5BxFwlBsBRz+1iy7aRxylP8hSjRTnH1IIoQSZf5RMfz39L
+UADdmnT0DdKbInG07rsLhLPUNzefR8nxdHeHPL4fnxYYseTLzaabgWzXgyYSpbV
H9AHx3x+gy5K1zo6Dflq68BoP2UioBc7K3XQYE0gDcb7apgdWROxu/3DrRatyDYT
3uAJhWgJqDselfSPMsSo08/HiFOlMeVHXxA+KOHi/zbJndBGKsRvRjS0STrcEQWy
jv86g9/IhPFnS0wxyZQzpXEKMSpvtTFmyAlf3riisBTStl7ousq4Ao2UdQlr9vsW
AmReFxWz6qTe/UOOGNJQWHphDGfjV/agvtAo/RZEEGOsp1FWxKSsFd48q8NSdqjV
6zjBtmCcIPGajYu4Tt+PbN3gGvsfKW7m0dba7Ys2AmaNpk0QTW6ciidD1xAsGKfW
PGbVzB3VDgpSdhuBrc3c5F/3o9OT8gTeQ/xLN8nAviyrLg98BNhKQ8IDALswH6Le
WFF+UZ2zLVJJWX9zhRCI/TCP3cT4fRxSFo0HehXsACmgx8LzGOG3VE+MphpE5um1
XBGfvofMkM9y5LN6RMG0C87phw+aqzeIVMQ149Gknq8M3LIDm6RYmCy7eBr7M2Pn
rx0bcxyl1sXK7ShVUJWWNJMYWZZ8ZEurRu8Ri033RRZuSK6zA70K9bduCstnHsyB
GJIOPXLnAwCrdGCKhJkKPJ4zap4Z0Fu+6cy8t0v6rHNUYv80+PL1gu7Qim6RL7RC
VC7OaZkxE5UTDUGTOptuyfWLtcDZA1P3nVVFTlo1XWdi69xERPXaUbEP1g3dGSJ9
0SKxSnSMsVy189T93k0HaGP01IpORzjIT38s31dUsGyM6r4h4NFogKiA1KtDSz8u
jl/1lE7/35LWWGK+S7XbUrj3OxpFl/YKmOVMkhPvHpC+HsKvuCsmozvy20vRvbSx
gvYGcmd9zvHB+EzpOx/Hmhw3tPHIaubI1L9EdugJBUs7LhtmXD/DwWcpSUBEXVz8
bKFLZLDhusQ2wIDkwwQpkDWlKdbtggJXmxmrEAaxBPwHHVvnIFNdWbRxPryUyqTm
eGIz0j3leV7/vwUnAr/01rVHbCciIjrhlS+1d6qax/wTANuFs8pn54IzvG11kcz5
FCXF0WJRBYjVAHQHSJ4AexfMnU2VHZKQ1ONhtjV6CPPf0esL0uKb+aqZB6qblQez
542eiJ5VkXhPfC2ahEbTdKiILn4BEPJjCc4mYEWubFQ7IJ7l7q0aMq0LUSm4TR10
thq4YtNuKhB5e7XRSPpJrpnXvkhPH11rV3JSM2xYu8oeyRX6DdI70cJD4TjWclaU
/oSQFmhpKhlGW+vdlP5+/gqMO7ZHgeKOsRtduzve7VmKulS//nmFvYHhCMAz/8jd
IkwJHEO8qjJ8rHgoKXINfrHhkGeWDbBMRWJQT7pU2NErXYs7HNnQvKl2VXniT0Rk
zsZ7oKJQixFZCLaYFjJxi4bl3bhUan06se428viBR9bP4iRcXNiFPftRYDM9K86m
ISpo27qlwFt10hSD2YvaWAgXTiG+RTo7APTWWGmKQawd3UGfT7enuXTZbgEQAsZr
D6O/yI1u7QLCldfwXYw4zwI8vuLwV5LDfQq1zhuUw5axIbANdV3n6d1l+vOnDqL3
VieZtifdNxkGOVGJEhecNBl1aesbIiLxzzC1NCll7ZNcdbKBisJwOQP6teuBq40S
482nhaZLrssz4AVPU7XtkFH+c01AGpeIT1oAXueI1xNkT5lltWmmxRH8oBnLPBa1
9+akfVffXs8Rl5rtxuGdTWtEA5sF0ME6FaE0BUfDq0avnwN1AIhdQUtnIM5EW9QG
Mm42yiv80SeE4ogVt1zPaQasQwoAVUmujepU80Y29rzajmHjArEy+21PlYayDKxy
V68+h9seUbxodU+vzHVGbXHvPC9I02SvExZ+aWCVlI7sUHsGBdjarIjouZObPTxb
rzDNXq+g/NkSsZhdZEWzcWd4AudwkyxeEcky32VFtkYa6ooM2vvn5aft0gdH6cR4
kUrE8NEaOqij/SlnxaVJkIeejlJRFimQyqETTU3mxP5+3KVa4jNdD3s7nvRW2WZ7
eLK33NtXFXYtv4Xu6mjns2IXgOL+Vl4lxWNBd7LfPrBPBzVS+Oh+Qa+olUBNIWHt
vImSX873CdmlDcDrRb2PiF3aVfY3fRisQUTKd8jOSxyxfKmqtmNqbb2jUutvOCkY
JLAEeSJ8TJu42sw/eRMOsIp11ddeIa7B1TBVSOB/3CqNXDwqeE56v/AU/PktUfLn
CjPQI+VYY2iMERnd1tTDG1KpqSPMWzkt7UeKtkeHaxm+Vgcvj8Ithw+7shYh/GfR
E2TfIz+tEEtLuoT5p0FHffqRje9Sh3P8HdairOQxxHzpHDXzy/HYMIC1Ej5Eu9el
nReJAzxGt2cbBHFRBrQGddQX/Te10Ju5IbI89f6KhqaS1V5vcq3GvF+Y2gYWh7V3
3M2eGDw1l7fa3QM5tY/s7yAg4Er+ut6NAwqTe5kY0puD4YrI8bxgrqqKdoel41wg
D1OF4uE4caJi+1jad3KcYaEs/aY+T4XH1amMFCprG2ltOVdgpb00SkRN2dcXjSGT
dmICLstFiHr4QCoUeFi7jMn3xpMXCilkWzTYWXWm9/2hFSLHyAe8+MFzn7ww9b6s
0G/FX0zI5CuiKLb8CgWOG1ZVrb4tyqn0sL+NhCvYWuK33A4p2Znn8SwigUwZJpK7
CoMhLbSWlriPmsi/xaD4J6NZhjzhXl37xKbqeH4D/hvGXQCx+s3oVvpyxwqbc7CG
JrUDK/3qbyZaX/mmjhifYCuuUxCuF/NafE3xuKmgApA8Sh2D8KjbJlkCqImp6hUa
0SVfLtusgFDsyqACO9EP1JMp+07pXgXYU2VYOZyMMU+p0QRSyf0K/Q112jt82zQu
h1d8npTgov+xjXBzgI9FqWj/uiAtUBNVx4EKa9h+jjn/BkVTMUpu4iN1raxKR0Vm
kmq1JUEoPD++MwhCOlp3T3TIasTtzaoYZGW4Zt0fbao1WCH74vnyS685PVwjLzD8
SH+liiWuDuMpNLkcKnXTvZ1Ur4ZC8riK77paionqRKm3NEOyBA8HyrJhcUx6/DGd
AYfHQI/A6lUqmaEwQmTwOv0QjsgGe7q262L2UQivbw1HGYZ8WdHs/WQY8j0rC0uZ
rigd1braI55HtRW41vFQOFjULS8UbD49Ilv3XCqkTOF7yoCuq1c1uMNKqpPOlYyE
JAh1aCHNh+lDBcCr6C6SuFZUrnxf6tTyrgEa7wVJMxesGOBLVlKhnjdk70dJc8eU
itPg65ittRpiQCpd+IE+w5lPGJT6F1Tg6g7UkQvcCXp56B5hWDMey2/uD+0u6ZrG
zuvMMoE336WgvrU2eNPjzJSXQpLXNNkysoqG3wDQcv5fak/B+ooVux5MOpa40MkW
bXj2250G3YVxgT6+msDYeUK2r0TtwBZv0OYHmGiOozNbCHGGCl8jiFxl5nQbSM2a
OOFu3CgT8zsz4cCffZ2hk4/jfNZi5vWWYl+00mWqXmgoSuWWJ1tg61DBFwwwrA8A
rHh82YTaA1cXUwk8IscrOIuH46Et4rCHme/NVLQvo6K6VvreepnEjksZ6zZ6KAsV
6urPY8+5gS+N/9cY9qYVgdK5+g1wIqNCq3WdOa/2kVuU3848/jPnDvv2ByBd3Lai
/97M6RJ7VmKCng2A8vY5Gw6U9ZDDkg4PUqhWeDQ6wQqNIC1KcjlKVKjVejnqh61c
jZ9U9IMf3wYhyhHqGV7fzzC7ERAkkgEpSzipgPXb2HhCnlbufN9MhPHDEUqHoSSF
6b77hggm61OGHLIPVnMfm3L89NZDbH0APrjtWbiR9ZfxdIux2w83Td/ys3YDOQs7
jh62H7nCAqP4DI3fnjIih4z1yjaCrFNuqbt2m+HJtkSxhVDW27kKBlWkEkmwmuqh
qQZOAOEEfVdnyORCvc6UcuWwe/+Gcss6zmr26COSCsAK4hzWXibundvYQbcyTaPk
ZSF9Vg/2+4G0GvcGjHCKlHID95aJrFuBFEfPJjLbHYdAeLNPpCLkrLLlPVzcEBHu
wqAtICKxA9DdaQk7IuHA/BzUWbRVDx6vdJC/WjSDHK7kWN9cDevcZufbDOI/bssb
m7oCdoQmEz2ZCkwCP8DgLBrqo4pgSwte8TnWlQu7BwF8k5JEVC/eCvnNIlyIMW5R
4kCsFZUgORV8KLmnEWG4C3uK1mN92xcDPzOZdCHvPdcgUD6Xm0TrPgEoHGvQjkxa
hGdw9URCd8xAxmS2rSxB4vAU2uDoiVi7Jkg/SgANt6ieH9YJyoR1sQZcK5G0nI72
l20L6lA8/5pBKyFpCFizYRqUzVlOjOPB7ZSWdf8uskdTAztprNiTynxHSFe23tpZ
kXYTxTUFpuAO4Y9vG45aFgonO+wP5hNtX8O2PpRqgGgU6oFk3QL37WmfmL4oM9Ca
2IHueDU68umbLAoVRgP7XKUbVKxdW0jKatl4516sp7liEBcPuQiptg7bDMxo1r5Q
b/3Acy+sa8Qib+cOEBlBHkxRwOERYd0esc0l+uts5HPGYwliMwxOGdrZvO0bwaCF
D09gfWYOEM6Ji9Mtzx7Bt+wERlrQA65A5fc4KIj+KbETyR7eF8GfmT4Rqq+ZNJ4Z
wy2ihI+bjQQie3c0xPogVVIAfE513C0eytaV9p7T+nxT7ZyISdh0ZUtN6fFsgEG5
4FQrASZ5yPJp9GQEp3bY6DieB58F8/7q1nOr6RX9+vZU1gYpC+kkiym9aiF7Um1W
zQDo37lyDS80BlBD6SLrcboag9sSGeUPpgOtzMPfBJfg2WZUsB1hgU1/o1aKkpwz
n6J1yIp6yi3ExWXrAcAknFZBhY8QZF07ySS+pTdqV8yvgCOuhRD4igKGdtLy0Q9t
s+bntIH6TuxsVCZbANAlpzEvKX7z4eDEUOXtdWP5/ctVJxoNqKoFcrZUqyimmHaU
zNVFUyYHeJT7WHtIAosNqBdM932TltCixhdHU6axcnaK047zZZ7/Orw3fbce0ynt
H2yhLcyU7XbC5efOgZFevKZa9J2G4vQZ2Tcd9EUXoTKpW/TNM9jPBybt2b248Y4L
q13Nx2WU0v6EChOaxXFAB3Wc07WnnfFrrRV8orttZarFHYf2LBMw7lkgRhy0wv/h
z8iF/X+TYsFAyiqgwBtx7YUyYcUbPhmRs4of9d0vQ8s7Tl+VOIHE3MPaIzxoWuEf
CBG00v5qr57YdGVgIEAq1J5txT+LM8IpM87dwWJp7BEjRo7g91l6e4/m1XpU3C0j
3xK3IgJqVvCJR1ll6Htl2UaiHbxxOrQQ3Sj0DunvPhBVKj41WXfpoQxlWD2pK/Dc
PldQjimvCOFuxFJO+5gLnurYaAcL7xlavFpdeCijhL6aPhu/R2qQ9iA/Wlh0weRC
qITvrvR2VoMQIFWjtIyw8++93CpMJOJoTMTHitcmojfRolKFgRZstTCKQ0wrCbld
DxwFwAm+86ydCm/Ju+q0INs1vvw8ua+x90LVSN61sdBxvP6BMD3s6yuXkqLSYxxU
MdrYFkj8YXKvuqSHW75xFSWrzWsZV2ghDmKfRHytM00OS1v0XVo6XF0F7hwRJHqA
nMkuI7FTnAbobmrzHG8kmkr0S6ZLgKwXuRgdPNK5f6tj20FE7mRfr9hcha5ycZos
D0kZCw23iLU47Z532iWkaCQoMhcrMZXenWT4FeDR5rHo6VyX9Rdowb5ikygyPEm6
wLBMplgP0nvntnPXAe0oG/ryZcgcmNXm3x2B08VL2MFYOAMCpbulV+yBbxFGiC0t
PrJKQCmOVHyTKhSHap2kPvxXrfjd7kk1GzM2Go1cGbuQVFJ5ZArK54Q2VIkGHocE
6m/jijYvkvUPqHzzlQlYqL6OfJOi8VoOm0vNUqvTZmgcqomIaSlh0R8CceZ9wrCf
jiaL9AoAQoCqmQueZICBv96mSmUuRJfjosn9ap+Huzm4MlX6wXut0RlVeSIPBoN7
U/SuPebGhZU5kTzVJRWNSf+l8+HM8gNvv0a5qbYdf7ftX4rapKe+YyDtUxaNDND2
XpaUMgm2iv0n+dMU26Mt4n2FQoTXXcz9FmSc4fkNmBjymL47izR4OJ4mKvUykRBg
ozM+kb9DQUwZ8iPG9zhJ4e1+Mm/3X9NVibLfXMCYbtj0cr+JoEqCq2FqkVGhCGb5
/74R0V8XJ0GjkbYjXU4k+8d+g2iMjhpqc5K3CqssZ5Shirp4YFsStJqc4/QKJuZO
PvHg4ibzbsobYoIh7fCmilnqU5QtFhYq9BrTQHPg2+Gvny2elKEaVb1pX+IDgvpa
M1m1SvOftcGbhX6s/5BACQN0FzIj95IOds33eh7NbIdIxRY9MwgGUr//vbbogLMd
vd2R5pPjoK8HTqqaDUVqDrnklDAA2449GeUbZ17w8S3jWY11HGtvbR/abiM3pLUO
/xbDhCh132rBN6m3JsDMCJdjIKjWB0KxWneTBzxbQVNogAcvaZD31Qaw4RbWEsQJ
McbZHNgadLxgpF+ULhUMx5xbOQN0inCIaO3vxkNn9o3S+81Ur8uk8PJ/f8NXVGkB
KdDBc2SgehRXIRRnhhIPBRtGLHw69LsZ6joYeWOQPta5xEttgL9QFNEkciBYWNZ7
JqXWd53hCTQhq4bpC7B3pU0G8V5I3iI2YDzT4PDBONTwSxzXBYQZ2Qiqp1NTFv0N
PkhDGzEXo35z9Jv74bakUYnuX28IbD/6w+mStZL4uJc7x6MeqDjPJHvXLze6LvZE
wHPGHmuDbxeLMYGty2mQ5arY8kLpBW5WMBm1fpKjzqc9+oagVozsMW4HwRmvODWe
PJoFQhMIjVA54DM2zrkA48t3INDDGD64iNym91wfwj96j0fXbi3Kd5k0SDRERm0R
L+3A5poBLWyv6WUwkOQ+op2a0IVAthaVtb+mEKPqC2ohutsD7hk8VMd9TMlg+YXs
qcPr7DVQwRVz76ktqM+odEOvXHmkepy7SS3+MuhGCIHxPRzr7DHtKGI37tL0zHuK
WqUUM9PhpREJ39LesrsKMwpXHe7otojN9k7jPFJwxIy2B+6LaiUdHQtyP3dXhAPR
2/3dEraOlLGgn/1J7bh/zXL+VppyfYR2E+yINZKo3h5K3SmP5OkvpE5PgU6aw9M/
yxz1c0r830PLfWrkrjIirYeFGdI+cUf/TE9c7qqpuoIl0qv4HhLuXXOvwr/k99pZ
wDDHwgHE8/BDxR07oX0mUAhzDWBHkSk4q66ImvUN4qT0oU0goSDS3wrCQiMWyVEU
z2PRcT7IcQhlrT4wXjfBnPWAmk3pTcZJP/jf64MDJzPcePvMDARyOjaM2FKHDLxX
dxenkObR7TsQuH+Cudrm4j5z7/1bV4Auolg8EHqkO+6DizxT20VeQTKwttvguQth
uR123VQ53Bv+1pXH5jmHVX9eGrx3vBdKX+q92uIw5mZTcY0iOwOShbwJWxzXehPb
zhG73m11k1DnmNIsubF8GjrIXRsjbGZfnEXQ3z6NOwKawqP+JQC+gMUmfsnH8lCo
HAGYkjnAlwPLu+Eg+iw45PSZl+TV9AvQCdByTgWXWP8cVux7hantcR8aAnKvQ+tY
HdWWvG2i+Tr7xK5l+G8HqfMqUuRkWjkwe+89NDpUA/aKrqw+FgLKQw6hJYvxndFF
8yyzmoMFBr6sAjzpIqvdYhq4A3qqfSyOGy4Z3CKx+TQEuspAKhNDLeqJOVC0RfIH
t0U/u9GPBUJYm1i5MehkSKyHWyFL50xNkYOrp5RBI8W4tRw4WpICNDSMIhH1hc/X
rDcPpwyBOTn3cFCSjhTGa5TuKUtFg13JUysOgmANlM73B1uajVW0xIbqXWO7KFZN
vTX6zwEksRvNPVQWNyFNEYVia1Cg3d1WBTH3nF03OyFft9LYO5XD7isVDZzlhZWI
FD0pKsgvRrnz8n/0OPglp5cqa+ds2GoOGFvpiXZDsEDxfPwW9deGB9baO+aGGXPH
maZDLJ+Kqrn5aEZULLGMfSHkiFX26WMjAQJd36dTmNFfePZPljTN0audA0i8+YCX
oBB8QzfaYhBWB08D06kTcNR1Q8iSjS+xFKxRX6GBSgA6Ktae9+HHzNKRhh61IylY
DCzTmUwUv9NwP/swpOYcOUoOGaH+JPlg/84MXMN4uFaDnGldWe8YmM0Ti76/EuAi
G3jCS0cX9N3d5nrdtZx7JBTJis/Op/jSpam8mBYq+4Xr3TZIWAm13fw8vmdx5Ar1
huQqRYDkrpASHqlcV18ItLOLjA6Z3Ym+LB87QexpHU4AOQ2846VvyjWi2S0uqIJD
xJbFAcFWxv8rJQXQs9DUEWLaWi6E5xmYXIvry0S0iDJfbnPhtWPAJg6qbm/hCVuL
hXtxteb8xxSd6+GrqBJ7Z6MZKaArancc/zIaSRP/w3Q4HjzEgGAasyF8uIJwD9An
HyBFdJtubUOlKEDj4I+ahyYj4qhiJes1LLfL96cT7eOXPzHNE4N+ETncmTf4s+oB
iK06F4xWKvOYjO8+0JWekvj80mDLxJvfNg1YJ+lpr0sllR3rRWSAGcoJ2xUiOvLX
UDJxyWFZAUUuEg7mIPZ0BdbKseEOYBq4rQSwFjum/bfshVzd+5Seez7uazemBMh1
mhDeoxNnQyDhHXA/yFqE0hSsIJpxG23AOVOO4MYvxmv+WGX3vH/XUBwfw3+2nM/b
acdTK8avSX+Ij9eqK2+jsG9wRrkgUrjkXoD32Zp6fBTm/9sH3Gs+KYY33D+KLyn4
6vGyTaPcqyS5/TZQN9ufmO9Ki++/RKG0MNHdQHtsrBEt/SyPCeq+SxQnNBYAOA+K
V/1WbkdSvsk3bxK3137rxCgYNue28HnaFVTr2gmdAQtDuAoBa1WCnKz7zDzl6SVr
kEZE+gqTzPYRb3mpHT6Bf8fwjCxlBdKnsXt6tRowI/ziJyeSNIPM04/gczv2tju4
v5gFmk+M8h7jTY9cyxMfOh40GaXJqzvShxcVg6E4UF8c090Nz/N/EqIkN+/a5qh2
LSv/ITe49BdsxwH5K/reSm1koXZCIqfJ1BsZBRClI/MLS0/qjC3Crjq+KaQYNtVs
YL42Pl1pFwHaRPhS2j0RfGaopM1x7iaQm70hS/TRJZgcO1XnaBGOD9RkicDXParJ
f9gI7P9ZJekKCWak/1lvVjIjwu4PlCaE6F5UdmYzuI1tYmVNFbHubRbMD3HKskhE
SxBbM+yny79DE1t1P5l1pfU8m056iEW3RYkAjIzcF4GCoxXJRDBeVf+XK+yWcGDS
CFrSiVSqeyyNO8VFwN05pt7hoeCB4DJycdlORXMaqegfPUXzWQLQIHh67gZlM0fL
cq8QTiBBtVUu8Sy9kSz9H8XRVtBX/bktuXXxEvFpDzCuInAcX5B4pdf4kFwkqL9a
ORwJWFdLwnV0zS8yqdgeHHvGheAKmWWqnUbkQFk5yTrCqhJcst0VGN1zLrdEyTHq
qzw/c2jW44x9zIiwr5wizitznJ1cIep6DoutQ3jiFAJiZYiJU7Cn0pdgM/003IGk
68jvk4X3VJ1jw6JRfbkKKNzV15iHqdTFvMiMhFWTSaT3BIqKm16YF3GZCJIjeITp
5rTgEGpycZZSj0oCfVCkaOZFq7Ev2Wq0Mjg8RDzztsXa7lfgqMTugT78OmzZs2k/
QLyjHe6w/HLSCUWmPwDzhWhXjtHgiM0lP/oKRr6ezgoK/L8aX4pdQU3Q2ozBF99m
SP4dCS5LZ6EP+slFm/FtvVmpLZQS/9CylJHNPEuGE2+EwdYzpzK8yvdp7Beg14y3
rGEH4a8//4eG6fm+qmGW46T02SNgPS3bY73gjsyXDhCuOsN0+OBy5daLB7P6lSz5
BN3MQTc93aKqb0S14HctqTpEYppeND8EjESifdEGGizjAxhr0Fs8kDFCfXo9jvuy
TyI3G/ujyLuNYToCugjRJmv41K58ofq01scX9P3CETO0qZMTD3P8ETpYWgCJz2N+
43T4PE54NXBN6HM0JeKgpYCnwKLleRrs7nPXx6eos6/gsfHgwiFGI6pyoyth1WGE
lA/1hdLMNuPIkyJ1dDkRZhBjow39uqhuAdhBuAJN8e46kYrk2bG4CBXKaUm1kUbi
bxhJ0PFOAxwQgwVu4vwgXnQ02FWbz2QtjU2P0IGwAdjE7VGQNAlHVJ6MfWsj7ILg
frajVrsviRBxN3LBSu9EDXh4mZW1kLa8MO+HFTB/9nKwSJP9U6ORAywhFqEd4qhE
/8kPKKSYWCCFZaLT1x8Sqf1SV7PC/59P2Y2Z4gS0yaRhTwBYJQB6sQQW2p7TQV3e
pbGz2UoAZlGb6poEsi2dWc2cJCQasXqwU0eDq5Oxx1BS2LuBhySB3tbB/6/6e6d0
q43lVSEpf+TEfGvIfLVSgkl/ZiKSagig9dQkggxjzvkU+97FPY2Q7BMLyD/Mqzk/
M39MN34Kb1kA0X3vwj483eWtDYlrB0Ae2v84mgtrukhvtGhgD5rce+Hga++g+8bS
5Yk9POHWeDyFlpOjpwVWPUBhlulyIrbb2VvvDgvpv0HfjhhHpwQr6mXpidxvCegN
jvOJ0SPPTSVcrgsksaRHGRwLrl94n84YxdZpDJG8O/qWCAqN2/PXhptoQn9S7XkP
CdtXAgRsEW0Wyak6aaeButwe1Qp4XSVqMinTJ2K3h8TWe4/yGSb4Mu/++SMSk++t
qVWh6+eoYHrdLROCmv7UBF+SeE6AykGiyjTdcZNNitEYzVXNPSxnSB+MuKvmBvzZ
TRjCeqV+/nHd9Sb9LGLs5FLEMbLrAp4y4ceyj4n6eeF9nsts7ObUEJ1YRCmFTaty
4APuNKbyt01PCvRk0C42N0bCnmPZJJFFSjOHoIjy9JIzMMq9KC+VD41BK4kcKYyl
2IZ2V7ZEiZRP4lWPVRvGlcRo90a1Vudwgf31cz9HD9MfAXtC8vLdBULH0Ip09/7O
UmF7eVQGwiYkuxi5vADp8VZ5QuYXjxYoqtSmtISJS0FGHJnvjZqoxcIKtJJrQqfB
rPRoJGTPIZOvJ0i74ndBXjJO+cVgIfrI7J9IXkIV62Lk7jjqlIHqOD1tM1AXnCAG
s8sKJHB5pAOY8B86tM/8y6FSop4q+riH+i8Cml8MhqxlpAvJwX7rjIQmZjMfSocL
pmceB+bFO9MgnC7TqFShHIQLgoMjfCNe/Is15ZkRZaBKdTcj5FetLLirhqfnB00c
Sj5ywXzzv8GVJg9lekRklDbYCxaWZtyA7YyHO5F3UR5JkP1+1P7Z7zRrTBFrGUy8
OEUobZnsM8NldgJEuiNK7ILVLHWFCyM16iUoQ/KpI1RQ7Z2M5iOGytkEGjk6Iy5I
yVGS+EjqthH8I4mSaQmBVsunyc6ThdOqG2FoijRLwLxN5wP++NUyWk68wcjsiyyP
knolLw4UN5hspJGSy1aaN4XG9zB1YYxXk+dGZblMHGYmXw7cIBbGuiCWI3LTuGJ+
jSF2Rhem3qqjKIE+BHzbcDSkBDF5zlRnGfFW9Beef/MnjgHHlYwJ5k8q9BpIHYsX
q+MF/sM0vkyQm5qfHDLBZAJbC3g5WXbTBtYUl2Wy3pCQI/cLbmK0iHVkeAPjFb5v
zc41X/mgcCb8G/x6RoPtn5SFcOZn62DU4ZOga4HfvjoXQ9e/MvreqxYhbB6ryJu7
dqVGvOXgznXHUh990Hb9Ltsxdg5xojvYXZei2ie+b5mvOe/Xqv1hXj7csfV/2J2I
uj0RQaVa/2NjJdX8Gh6XEv0MyM7/d/lAuUVeBd0oRuUY2gDR98nUEBNFSgWRMs6O
9wdDk0C0v1nZBcJUV7C96W6FC2Y/wULd6B/f4ns/Q0tcuIjL83VDDq9Swus3WaxR
M5Jl5gBy/1KAs6ZXCeZhrmY6E57fFqtfjG6pNy7YAlLK95Kx4OQfVNY55GA6Bnc7
uykinenizphydj72zJ14YCzK8ELotIlV938FlmnT/lJs8ZZT+bkIrqiQbKaYjy/8
EoXI3fNkgB7J5LR9RQd9W+xwgcARlrI6usvDH7/pBY6WRAFmA5FUIh4nYVroX8EP
WL5WbC/IMcurQ+GQxajJS7XO3sJ8mbQxiMSls+GLsEBtALedMNO2kJg4CwGYl1+S
wjmknRxa0tz3mrZV/4yvfty2O8bVWwnN72oCv7u/xWo2TahiOUlCzUZapx03Znug
JxgqwmiHbBn3N/s/kHu3NsVA2eIEkUI8g/GacyBe4kHgpiGahzU6lAAeLF7/xoXC
NziPs7PSNDR81M6Ro1GtiYgZZ2DcLZ06veXw62aNcTrviCNyHmi3LT+4oarl/rQq
2AIeKjKp3navBYXDREoIB+YtJMyFh/31IpZKvVLHsip3Go5pYB6AaXp0mdM35eMQ
+qxdsWFFH8IlRLBLqSucl1Dzoq6VkTnZAZtlD14nwRZdnVP9oVGZUvnlGhVNF8bD
VQW3+VlsyxRABNXxtMnYAv7j1aw2GtpcJpRwbQ51+q5GnMfRJXxGWA1pVcgb19RQ
xeIrt5oIrnuocCyue+XtbVJfW1XF78QCzIUJhxJBGLD6M+IvQRLd1qh4dLBAP1GQ
PlkmA7RWke7ItP6gY36BayCDGIiKF4C+hbmDO6/ABIfUS4uDM7GZ3Hz5qE7aFgqb
7TW2f4s0J/aPB/wEuBrpugv0Rglhz2Bu3cj4ahRnKcD+qV4aKAn5W1DCuTog+Fee
vAcRpRbbA9U6ttfG3wuQq9x1AD6QU1nLNomZI/ijtKmZh7SqMNA9zX1+0a9MO9vG
TmBTQdW68528ZNpDsbaUQjeVtQykckmkDLHrUqtQfBBFwCSbyoi9PHSDEtoAdTVS
npiB6jvCownqCEu4OWYdO0urqExHWTclcpuITZpMsZbDWtCPuQsXzdsLeyiNbBKz
7inFU6N8Zk2BawKvgNrP5+BsTiVXSQzkM8kan527M/9lwj8FIrmFsaafGW5G95bV
OpkHXRfiOT9hqIB807BqutZkhgdN/Xa0dE7pWS483Lyk6GUhgkzVkMuiB+Se0iNf
9fiDnxyPjX7qstdthPsM03nexTi0LxMaD8cZRapBT9nLi1j2Pq7tG4TaxOOAFpsl
UJITVBhx+homzU/cfpWO9j0rqfqwWIfmPXbq8OB0g2qUUItzfWOkmaxYfHvVSurj
dw7Z/SkptqARFof8/SwYXh2yhGyh2Nw+uUYImAodBTYIKVRyw63g3fQCbeBGATgB
t6Otu+JK0pcsJXSpC6KaJ66AcgLmq9dIQMrEwvOG26dswyq8wa9xjjaofNtZ/5yO
PNtVGv28fSTiz1YppcNSB7BzTZ3U/96Bbf3mYtjoKUMHGLQux+6EnMvYQkVYqLis
wg0q8EJ6queUFJdevGn1GVwtUUN5E0T0FRrpLm2//21YfgISLLHcHvMPeOyhwrRu
owXgfGYgGpT27xxmVhYaqGg/t8EAytn0E5I8kHOzq8Yf+MZ9wWDHbPIOOF0S8V04
D/FlmgxU82pYrMCL/VTolQXaoKqFe7WVRBsPgSMNZyooqxeaKuJ69yWoJca4wprR
sNtZT3DYkcGM3ct/C1UkTLBlq3I2NO7G2x7BJvnGlj2hKrs1Pst5Uya1soN3AxZH
z519omiHg2sfERZpBhscJNmE11Z4sQcPmvjZtGxWe2P50TW6PbpS1DePz4aVopzt
rMKfwQPIeOv8i8qH+p8fcZTxVnF9lMZ2bq3FKVZjXTQ8wt+3BhLb9VQmEfaq8oor
dVTT68WdXsNEwoAqCyAeUjBPUiY2TatEqWmHWOTS0/XwH1a/MaWRQAO+65YVjWH/
IF0W4eWMxsOeaXBVcX9YvlM9bYY47QYI9b3fer2es/iXtX3wA6ohjrttJK3e3Dzg
f5yr9PmgobwIuVlTNh14lZ1WnlPL9xOJRmi3+goHX5NT9zXUxmOpTV4UXPU6Eqii
n9l7RzJPbZyNUeWjOcjSwFII0AvCBmUzJjG2ZG67UxP4Hr+IpvofMueyxFzz1w+h
COymSj1wyR1i/M6YwxYN+uPX76D2E2BwIRs5RZhftqf+b0O2Bz/lBmdphCYsd8nr
Ih0M681qrvQyHQOBd2gtlXvh7yL8C5FUXTw2I5TQlfwK8wLQ8XG7XwpFAPtX0dgR
1noWcUiIOJED1XOaSZ4zZqYhHlprIw+LyFVAwORHduDwgoqANbPNKvkJlRM18naI
rDnr9gaKoDVwFYXCCQuTGaNV9op/BP27p+DJFIxFgTeVhDNgBkQy76CvQ1ZocGKn
stYFeYZJa/6hnbYl9i0lQ2JB6qCyQZiEsCgixD8mHi/F99DRyTpagJ5gqGvDlAgh
7lPN/xvxB0Fb+o+KxVc9EdWLfE4traj71pB4VXLDWgOIiNLINE3iK2apY+m2Bgkx
zJy+gutd2ffVHBXan5Qm6p/WvggVNE6PPoVvBX37bG7WOH0rZkYQFlzlnDniWqp6
6T0EMM7uEaUi08kspI0XNsFjTEAEBpf3Y5XiCXW5+c3Lgox+I/6A6EisewDnfcrH
ZN/1LvKIdHEQwIMqcJoSCqiCJrJ81OlUmuIcnF54BA0hX7YHCcHLmA9MK7huWn9g
7Z8O0jACdY2jSd2wDfh8XN4Rk2u2L19U//8olxz44jXTgn0MwAplV3PEo9Z15B/+
Kq9XrgI9mpOqw0PXxvMvKcoYtJez4it/vmD5gd4RCsiutF36DTZ2XqlRXlY9+1uK
g647jgzF02yGYkOUogsx26mV0N2DBtVQVegfrh0708CWSJ0XgmkRrIOEibVeWrut
LkG+zv/QiNZUp/jKB23KcEH4lgceZZGV8EGHb6IIMFKVN+VNsjrCm1B96MHHicta
fbA20Iet/btMLhRqks1X3YHTtd7u5693gWHIeJIvXfueC9qFGh4kxW4N9jPMNsbu
YT8rxIGXp4z7LP1bA/0twedonh06PDEE08YEr64hHAXVLfLUt0mOV1FjEF3alKOY
KW4LAMaVgnGXePD/O30taf3s1a/bsBHgxJKLDQGBwjXqh+W98jWTc2pasIMwwT1e
3y8WjCpjKsynR4JqAawSxWM7CV9tRfsicuP/NOIIQmIXdGUEqgllcb2HbgH79RK5
t1ZNIagRx5KBpOeh3fg2FFWTmlxNrNb3cgiuiD5ObfPRcXOAFJunvf1AOLWl7XC9
fbE5QQsUES98PfuCWAnoB37qftT7mL1gjEbNXwOXJqvMnkqcRU2Jyw1K/jhfYB5V
HLH0ELtlBTlz4hQPn0Ljzuzge9yUf2Nl6BH1ISHvQucNLRlpuEg5ehVog09akExu
O8AJT/oDZIbV4pAlxLZ3x3cx1/+w5vgQRSh/Um072Wprvj1IzaRJxxItW+lDPCh6
pjmKKzNbS1kj5PG1HIWyQKJORHyFhAxxe0a19od2DozH3/9m/E6ZKdD9HtNV5JdZ
csfyNf4n4hlN3nQ7CbXhxmXibeYa6dnPFEhq/dOvS9wNUBxIr6U7xl2bR8D/OHIt
2Z2h8KnjE24YpBSqGEHgPoZcfIO9t38usqQLO8zFY/pg88xELkQF+y7wFJARMZxF
EHvnHYNAwplcZI+St5KfZsvE7C4c0CVHCGa/i7aF82nrAQ06FFZcLsOb/hYMT4ME
ZBMNf8Ls9A3R1o8c26sA8C+sAZ80gAtQqXHjsTpMOSl3WFCiBjChfN+VzdqdXZBd
rUkN9c2LC6e48KBMNWxiH4iGrDxeN2p8HrN7OPVlpW42tbHlRCzT89K9YbL8rYPP
/BDLAkDnrxH2cIvuJxz+dNDOWfLDS7xjn53iBXYFuZTEXyhXul+xuL/2HnPYVMEx
N0O10ClsgKFEpLh55FznbZQPyJKMl1+SLsuy0dlMlvXUrZfeH52cm6KsFPSJ6Ma0
D+1iC2/ko+G9ukj+V2wqY4yZpYMPdUwr4VvjDcLf9SJIfmWkCN02C6TfMmSrfEXh
kk1Nkp4WG5Rxjeqg+pdnKRIssRXCAli3NqWoQo3Im2+gIqAvmRLbSoCpgo775V6O
lLKDrej57tuuvZN1VSWupoj54OLFxeVdNcCk88B2B/kJw7bk0zI/1qUtdUASQ3Lc
PdtZifHydK7lq4RV0oRp+L9JFhi4M7kMr4zHMhOc5QQv4juTLLVGAr0tszB06sG/
/w2+Fo0usZaG+5E5cGIOwHQJu8XrJfwptlPS0teV3WsjR2TDJd0Z41JzBqJwc04a
Dkw9MEAkIz9yqKujXCFN+KSfD+bX/w1i2BvBVqLWrZizv830Rg90Wbonyx4BScV/
TJdthExtkvj9B1YQRTWYJgThOe5+I02Clk2zXW8+8x3KdPpUQRukFW+QjASbddzH
RBeLt3/N5lsHE04M4NMo4xFqrTfT3W4F+7J6UunwLnj13/LX6++LcwKhXDiwDc2S
fC88uG681a7bavLFFM099r4xG4RVUeqWoIN7HFnbIEvSvPYO0ABFMM9EOdaOJCwW
5RinO5EAxjHk3apK+/29gG5TM7HevNq9eEOOJaxTSZWxPIkUVig6+BhjNozxSVTk
pBrcr1DefBLLbHOHKl8VuMk5AHRxmWugnORUme5QxcdLodZa6CweCQi6BFU8eipY
lfE7yEPqV1pgrB9YhLukk6YcC8+Vlmg4im0yjuFJMn9gZkEqkUTmOzMmhrgnU8VD
5X2Yk18W+YFl5SsS2kw8s/1m0IdXVpPvFWnTwmddtn1vfLaE4Aj890kQIyN9UXDk
rr6QXb9NX4nUf5xc1byEGsi78hRtmLGYtt7v/cWwmoxnWezbvWEsfk5JOXDvVgzM
aASHfXp3DmKawNJ8wExauR1C+qOel+5lVXNpOP4OqEDf6k20gUcaCUZ8CaJ2dt20
D3KFIxMJK7+iyhskMP8A0F3zbA8qjZjPwIJoAas3SGb48Yit2lq5q6c4lO78yrrC
DjLQ9zvcvWPC7jQGDhr/DNgu+4vn366WBaJcbN0eVmgJRxJ98nnXSIB268377oHr
ojK4TKNxp40UNCIURZ8+rhZVhbQTzXYbOU6otxfzz+iaWJH+Q+sPx6A5tJz+3yOH
IKVdq+MvK+2035c+X/N+spzBimf9I1fqpmM2oiCiTBeob9K9hXgZI9nCYansYwPn
RdKCKUaCvDYoQQZfXxVxMG0PICONRHrqGYZtWwMptFS8Y3RgIKVXoMEZMLzsPZWi
fwXQNOOhVD34LSVgVxCz+x3tflW4lR5tjOmpGbvHpwGj9CRq431N3GEc7AnRgcy1
xppDUS8SPcOO/gx/XL4Mrw2HGXnyZ8nktxsq3tH4q5Yfk4ZK0TMvgxMAifwJ0FT+
rI5Dkw/Vf0jgnDmSSNFyaiB4/xU054jQ6X42FVnFi/xbTdTDlM/Gb78ZF60uV7cb
i4Vv+jnRYWsWqMl6aIXKOaZuESd71PXcSLE/oY0DbdtxbST3hdTd32fXAOomgtAN
GngCvAyryvIEub26i7ZBRK1OqLXG+NYEZhK0abTLJD5EYByq7ODc2Jueen3SRiHh
8SXO6JkonpawJ/DrM4HDAh7jYBvfIW1Z6TuDyy40CJKTuj9qFLYNZ3aokkQ3oOeP
zVoEtnqE5FyHo33QlRGIbSJDKOPry7mUYunW7Mf7tkxZnnizdF/NNPcsiarWqhjk
pEGgMHNB5koG47iq8y1hKQt8fZdRSU2ImDBraZYwEUI0qcyu93BusnZqKufvDt4U
JIom6WInj0ZYBZsBubfpx+HAUUaXal/UQqjXxxDgYmrdj/hSIMcRKBXAE2cSoKhf
6yWuEO5YCfcB4jhQ3EC062AFoxdAfF2MfMCEzupidCTLzSa0K59jy6Uh3fBtpzlQ
c+JCVd6mcvzYiqCn+RkhJ+RXvP0JKFQTN+w4mwO1a7eaUi+++bQRaEFIh2eIons1
Hn6OsueNrWJ96aBKLSW4QD84XHZzhXk4tGQc+ULwjk6nxms+yg4SI99AtVpWnw0b
Q15BmlTFwNpSuz/pQuSQjQ9H0QGTJq4S5EWW32iyP/XQNmBiiQoRTfwnxWd0LL1k
YkDio5H+LGhx98hLKOwLK3qD16W3GplqlesCcKQEykRx9IVmONG+TopquRRwQ4+l
6tBjrGdXesp//YF/eL+CLJ+yFx2ZIKG/GxgGd69sVHJ02YQSulv67cm0ftDU+jVI
fQkdaky/v49eX8CuMXCqJNXzzoULf8/D0dr9S2acLLN8NSDOHARg9hu3QdKjS341
C61QDxZlp6mOSr53edgDztPTkwmBHFFjP4Y+CFbZizrQ7eBO1mt+KMusFPX1uEEd
hKnhdj7JjgAztcQvWMXWfYzzDqG3MexQncvzBzymWsN36x/jOdILIOuigFYo3XwZ
vz8ax7FhRxP5r/SRPnCKRErfriO8ZiKVb08PIfbAI5E3p6+H5Lf2wJJqak24cIds
oXuAlmT5xTKyzk0A20BmKyFhtx/1WaYtfzLO0DyeSpHmnM7QCiai8W1iDnnlqO+Q
/VTyEohOIJ74NKGMZX/lRQGd6Vhga4DchiInQ6mqJztfx+b6C0ruQEy3AYv2YWxG
cjfyTkz3gZClfYjOqy3w1kzYOhWDm2MjwSiYe6oxGtxGn8BQxFjZL7tzVgMP3xwD
bgszYgluonWR9CMWaUn1CEZBYP1oIoEDqhAe2lLM15ju0Fe8XemmT9rya9RJXcZM
OgArRUyXLZaSXxJCsJgs8fV5bZYKb1HCUyAzjHeTozD2fY1LN1gQpYQ0cEdFEsER
lEw5Xcu9eCrJEli0FPwH9PqHxejkojXxsBaMAWIY5hACUfbzPY8mNsNiCI0boQi0
oefYoR22Z6jX5RWYCUWK4UV0aVnNmpvq+ugerEE2jIOpaGYhjg1N+MPPhFMdOcbH
eCC8IaFiYC65oCBjKmPVC4tl3dlvYVor1cHVKNYYBK+RZQxAyrah7ddkZv74OGiQ
jg4r0u9no+duWhrB7/ck4t/gjnZYg0420WyJLgzmV38JmRiQSRTOChBWCBPAOo2e
n/Cmy1ZwsvznCz15AkxLBbXJj2gB1vSWHVQV1f00KLBe1oO1IThKLKNcIjVjEQn0
nAUSMEjOPoLboeuqtZbAHOC1A8c+SrGVmOUCtiqJcS0W8nikI5J1mEvg9uM9bXJw
SxkX3hMqwni2QgYracc31dFf7y/25agrAibd06CiF9y6wz49y/yAdhG8SxSHCBBv
+U+M1++A5nLYNBwmm+JOEH2d6bL9uFN2NmaiFp7Ub5MsjsVFUjnxpqhntlezzfMv
n/C5ZaUbn3x1OktFKwwy2LKXJUyuAJ9uWlfEVr16IHuWAdw7UfDWse3xob1hb+j6
X7tkhaY0Nmj+usSdCJxSVkeyEHDRSlC/3OJNNZGqORg2XECyHbKXxXIn61Qikfx6
d6uWuHz4TgoAFOyQWsdcUdJ3HeNkvmLm950p59LPSqqtXmUHFXw8eA1FPgYLC2tJ
qTfa2AfQRds7Okq4EpNw7fmchgLPlPk3NeosLNJd3ogshaMyAIT7aF21tm3ELsw1
iPXUVEEp/e416vs9TqZzdZrO6sxVFzMyYqRXMPvIxYxPojdl4vR3Qu88MON/drNM
I9GBj4ehjbwQHi49NzULMTequ5t3UvmlMS+ivwihUsnT0H7+R26+s9gTBPZS5rqZ
V3DX3/CcbS5dbA4Nwl6CCRxXdbVJECp3XoVg4ffY860zY41Ltj5k1vIOPVtN/6E5
coiQhDPoFcXDcHB81aPwRP71lsMa7yw46/xVAUR0ztcl346FEJCxIT8u3XNJSe6q
ZTZzjZYeySkyTmLTtqjzGK1+EGvIhHz14FzYjHndxAAsQXw41ihqUu50+wMBs9E3
lEsi4BD+q45kuOPJhudp0EZK6vf9DHeINdAUrzY+emLNLZTxHb1XzKdU2M8sQO4p
UF2SWi1iIaEoVN0S3E/Gk1DAVEHbNCg7wFljMsuoxHbadrYhlTqA+xofiMvaVozG
CywTrYv+d9JzT0wJnniSH2lB4kupYL6aYHzJW33NwbqV7Hj1c49PcFKE3IA/tjku
AKysCtUbEgH3bCCJGFbA8AaCcEGG6zqNNiFQXuCJHdjk8ADriOnmzVmNrivpXbjp
ZijF5flFs67XYWolg4z/RBTeQ8B3hHffqkxtj4BHLKofZ7+zj40kFWbk/rY4KX7J
Ra9zDcXA+wOP2HN3ZxEB4Nyfmw1Dnm4LS49RdJofCfAaNdIIT3rEA87WoxkF04f9
hNHWlhNcgMB3X0dTOOtfxobiG/Atd1kAIDtu/Xnb6pomDD124jh84wPrxsK6iIAF
Go9ZHWfVa5ml08as/0M8k10dckGYKseEyzmdm0VqT9DwSWW1tfsipKC0Hiht2SA1
TjnVHxZCJW+vX5ss4CfoQJLULPO4V3/LogDvAImkMFsp2hNJlCnJ+4B+FZmFQudx
zQIZiAyphr9r5FNM89ZQo62mNzorMLk1PvEGnerHqCxoRBr7wJjHJOsy93iLgah4
J+rhVSWmoAECuWxNkXG/9tqvxgjzatk+qqH9OhwU+1TFEOYkewp11KrMk/ZSOqOV
FfCwkTvbCi8fibq427uz6KfTa6p9c1YRWtDvdKwrwq2uFYw5DvvW6fFJqrvc2DcQ
gmJYPKjc1Vrfc7GnTXCRGSL6VuJaXOSQjzPNBKXBPdTIEBKrj6g6yRP2jXGGlgol
91+IrXH2ySPLy4tPvzwfoJVP+Ki1Cio9R7zeyGdMeQ/f2rdMdczqzl+DF4g7GZ7s
/cBeP2svXKIqRsTD0L4zD0fT4IFpaauNAOGu8XCKlQ2c3lOnrja8UMOpnmHPJ4W1
9FjpIbYDAkZbukc2DZiOq6aBxwFaL20DLLNQ9k3FUAuvwm/ZIiOcaN6QBLowGC5t
8d48QLEBh+QBTCLQWYStwn8xh0jJwI+eTKKqRlStG1iWxxTypCpCxMr7hoG+7fEd
5a4tAL1R4c3EuVDQHFKphguZhUJ/WJrYW7xYpazv4S2+hfY73In3qD9O96R+czxI
fRcP6zkqMOhSBQKoa6jc/8antywZzBfsEY04xRtJJmZ1BZmhwQxfFBD2EL7GF6lg
37rV/sBZDUQaGeFogQLAVjZV5QAExCGA5gjSOpbSszHsaMhpjqx0kAizZ0MMM4f0
/cC6azcfs/Vu0GXFM4JyDphIYCND2flJYewalTKkC2bGdOwLrWS/C79DOYUJvXnX
HShocxWyn+Cv7HZc5d+d0z7DO4Oq1xYzoEBWUC1ZpwEiRur6FbrPOaHL3kMwYq3Q
BXpwe5YFPudtHkGDjkZfNA4MeRJfszezw3eETS8CHbeLfOJs1oE/FGGnhtLAtJtW
BQ7YEx+4v80I8OpLU/ATyXhcHyFfHjqfyV143WA3Yev2pDx44qnfxFgjKs8qF1Ao
Q014mJPuumK820Y5x6cPpSeWi+cpCTaMr3Oyk+0pe5ekzDgfUHCdQst+QvybH0zj
Bw1VpBiqsR31Rp/sKFKx22Pdf+aXBK57M3BNmRev54mAUk1XzVUizFcnoORWHP/L
q2ekyTE6hpUVsYBsvnI1sUL/58Om9WMpn6kYPZdLcd3uYH4UIyWY1VfnQHn3qz27
YIVIKXeW6+AFo0kxDrGOwzf49PKoAne+mnJlRZgl+m8S2aV7KfiA49W0PL9DbSxe
Sh/JI+oZnePBIGLICWSOVsw0BHsVf6/NhkBH42NNNVw+fxNIC9lNWYGEJci8HOBQ
wjMGI/RKF76Eqw+dfLK80ow1xAJS6HVy5TNgNpWjeC0qXPdG1RtNhR591mLExLWl
YPHS+esbBnFFc08kg/j5cWUiCwelfY80sNc2IhgufnCaH8g/L1dtjw4UTRlz+J2e
f6paxrLHqrEwsJ4tUFmD0zCUSBnOjWILoYVMQTm22iC1M5es7gJKz1sLUZcRFIzg
7RNIb4x4jI0Kfsl9fJREkYg9fwn7mWHclJBZNT3eC7OMItCyx2Xsj3TqbCzgImFq
LFFRugJ5iaNes0Y2phBHDGrsx003/S99xx3d6tvxj4gGHNM/54rhQWC3pSeiM59h
vBEeYSNMzPif83jr6VGJw4DZR6shYaW1mmNYk634nwRs6Duh6VOHe2mDhnR8guXF
VIhHXwjn+NG9R8TSJ+cG4YRPDXC90wZAfX+6fqPDZ0Zqcdo8TQProg8MgdwyjPmN
VRPP0BSNgenxxtRopZkNAtkBoWQVhSLGo/i+cxVjy3zl0XK4tNCj59JWfAOaW6hj
X5TkeyZteWblF2Y6RvVteONuLBi/OQdiNRTPXGP3YiWlkiUlH06rC0WZ7KltbWo/
U1Hb8mjvbo8xFnlWYrLXUnlhtucv9NX6qkTa7uBK4CibndLjdLE/s12M5IlU1eK4
ciIxBQWrA6o+GwhIVlSl4FP14PLmEUcH12OdMzaV+GzpenZdRvwesb7ms34l+vYS
mZ9AJnNWQ4J92vC9LWXG8C/YmdvZ3ciVwluqD0r9WHzROChMjF74OUa7x5AuP6Z1
camzpNEq6HvRujgkaEjXPVV8yiD6LV5BfnjPBIaIyM5Cxxd0g3YQmAEpS8VIEbhc
cWx5w0k6dddh/y0ud67/7S3xR5wFntvPULtRujMhn2DX19K27GxLuAUlAI+lxvRS
iz+lDrCh26CMFcVti55Bwl8TrQPD8cMvsUFEGSmYvl8hlzSMTyqHbC1G1EqvMzwX
NW7HUj1hJBvW3PaByMbmE3uMZz22O6H099PAkxMwqaUJWaURSzJrMS4HggJz3sMj
udoC7OzraY9vAKWtxO/M7ozTIyxC8lJv/8vcp/xI0vbaPU5R/smL2zzI1ajC+lYW
VqsCB6MXY7zfWrj+QUB2ZhhYGxFbV11LBWdRR6ep0Nuy2cqw6cMgypjxpIS3ZeaJ
9OEtHVVHTpuq27/UtaSKRO8P+0WMabboiGew31k0ZVpKRMf4f6n9/OPCHZlpkeiZ
sQRTU7ZG6Z/FvqxJQzlFAzPsSnMx/cGTMxZayKBMJlQ2k5WDbVvvMaRyOVFSKFLy
WZO1iaaSaTDDzBxJBluv/Vneiwib0HDND34lxhE6pybmIDUzQjH2vLl9fASCjpss
bgv9SYXhqUtisIQ71Mh6XXCetwUlRR7RALGHh0vIEil+kDMqRbLzsonRi8Vf8RAG
R1XAT+NV1QV5ShHKf1IErukimLCphiAnGhYGpkI4lsaHOe0vYFyb/iniuZ3IqP5S
rbhXHvIbxjhBhLoIt670Dwgff/MyqJMh6sHztRdxJvIAjx1R2TzN+OSRKmRYt/sS
NH12QeHxvI+0R5H1X2VwYPrGm3Zy7GLqeHSrmSIXtvJVt4+uktOypMkqeK8B6cu2
wilIz1W08vFeuny1IC3C5mj4xNctLZCr7eM7i6Wk4ZeJl8LEXKredy/9gS7rvd5Y
Lz3UwMv7nj3MYRRAQxXSeurIs13SDfUzVToUFXQEMMG4mxyJC3RM0efNBLurW0+q
S51Gql5CWbafVgm5LCaNslflIu51PDFvlSaKZO01di5BTX7hFWjlBOMaybICQUwk
QuVFXlkSbs/T2/hb2HwyzlrjFzzCmpMyCKAdb58knxzWpi7K02szGvfRX3ZCNJvn
9OY3BWTQbFQ1QrPEGt4OPRPYXCjwcHyTxxoZgJu3/62fi/8y/7EcGugtK+4Q34TL
PFEv/oBTfkaJdlYIOtfcHQ8UziXJz/G1tPLUIOipv0RYcXdeM90FwNbVIPy+squC
osgpJjvPn1UPR8uPiXN3HMeVYTtz2GIXiSZjzrrmVtLM3TbEWV6Fkqt0dUXznfjv
qGSXzKKnmrz44jtY70JhUIOTUnoUiLEG5qkX5K2nqxzRmsRGsL5Q5LK2XsjSZ2V3
AR3DajBdBX1i1CJgL9YYTI7Fk5Tb3BxQD7GEKHNkJNHbVmfeMAb1KU7Uf/6XbskG
eqCKRFb5O9OHKd+KBEjwUW7T9JOB/tEDchZYQUlxItbNHC7f/mQXgKIE/2F/3maX
cVsc859rxZnE04eWcqrSDVwxZ97uWkd777IZLlR6KfsghxOSJFyQ4OM8Pdts5J7P
cDdPdFICb+l/EKA/mIF2XiUx6wLA4ES1L20lpl57YAcxMD2IGGw7tW/oaOEnWxC3
swCkbFUBcQ5Z+ubx3SZ9hwE6/SzaZ7OEfrDyFjVMiceKUEL1IVU8T2nNljH7M3r1
eH9gMY8Gi1OB93yUv5e/gczlZTHtOzkX/WuoU/IhvShtA1sHHR8mnTuJuOc1ChRg
9sg4zBCWEJEtzFQH66YSPnu3is7OIxcVeTzmr4nELFgdJNV11cjJcWD0GHheNGsI
ijVSDzgaKEU1evy/c9kXfgl3BlkuAD1xALvnQTHcwKnuemuwZyf2T+OxgyJizKGB
5M5j0+33/ca/7v1kNfbrOOThlM8Eowxx19et61+fxVFBMyW0lDmT+clldtlBvRiw
wr2a6E/DIW3dxVeHXvCRRrble3FH6HkxA6fgAUIFzs5pEyrdbyVdopmfPTKQiE6w
LKdYTcAtmU8pPka+Ay02rYx8w12P9Z69dtEB8BEf68LDl9FwW33fInUIBmEe2nYs
7VTuLy5TMm+hVcb2yCPWhJzvqE3FN+5yqaeCz4zmT4zsHZYOcTN1TVTG5ioKV7kB
gUfCs73/cJ+c12x3L30jsA2k6iKFau/PE4KSuUGR4J1LNCjHFgv4LRWQ82n5of70
9+KsVDrVcavbDpkVpDHasTC9btWZhw2+gYWwHKboMaguAlhNQfewSX3Qe760xMUN
DpdXnxfBFElNSfx40VZe4i6XSL+qqhz0V/+4Zp1sZbq1XVBt249SS0R9+0mkriqT
QjUPaJObLVptmla6ojpLORR+6GZftHfM8UwEFQNDPhK0CF07U7XvmNTrNunaIQb0
mVxvyVDOloaQVjbmD22dA5EmRQeFiL/RWKQ9T7lblKxKKOMmxoTf0xrgL6oUKTi5
w3A0LFdCfpGi7HeHhgKTpJsrvizrDO3uH8NoHz0o5zJi9ptE9iNlUdXImrGMCslT
8B0aB2zqh8IO/SeGdPLBcyW+CvIqIgmVPI/j/tgyzr7/k2Yx5HuYaVFvl/XTgJkO
vBktizazBRdKcRgrLEBkVAAfDsQlxtJJ4zguBQgn0Qwa0v3ZTKow5VU/StIz8fJN
2skGQOGBrgxL+4QzMehDR/fT17ka6YK70rbIwT1B615wa7VxXVnGH28eoEGc2AIA
p0A5boStFc0/uiM+3Oe6gRNrADRUZ5EdQobs3KrtKgEYXaygzIiY+dxHz85d/Td7
/RGlAS60qY418RxqCtjYoI2wiTbTAQd2C90i1zCy5L9rLAKwGF+PpRLyJHDu1Ha3
EjVKqS6LXNiOxrPrOY7Pb6Pk0e5tzKC/8JqnnltjRDpeStqhlsBg3fy8FbPQj1F9
ftc/wGcVVRnpgCSnKyedEnRISnvxANMWS5rmnIlVHYV3382UovNjku8ffoVPD2TE
Zz/lRo/vEw8CZ5H/G5JGQ/SLjEcuYksL9wfPEUD7ESD+/IsrbtBd/qV8XOULR5X6
n/K+wBBYER8hk6jj3O3uBoeVA2WBTbGC+w5m9MkvGCR4Q3tvahe14nBUZqN4yFtc
VcYjsSHUKp/eOzWe1SRs9z3Z9Tm28QuK48Da2n6GYntmJwLVH4iUDl/e+pOb1tNZ
eHlfa1gm1PU8pIsmrZBwqU8ynRnnmprt3x65fs6PKszOiSVIORfCMR5wqbwE01oJ
nMWZLnTZo4h4Hb/BiDpV/Cf3UaNmMinVeSYqtca6zu0S38/3AFc1IijygFlgfUMd
RazrRb8hzXNS1RQaFUoNNfrl+vDGk7zazCrZRq2OkudhJI4g04QgB4RrCqxKSVAB
3EeJlWrsAo6+rdbUs2bSW+0PE8PoKugnqXLP8akhZoTzjn8PDOLcv/u1XHv1VZ68
WNY/xF9FDDGLPalUWmLm0cS6pFfMWGHWe6+RfK7bqafADcFzquNjjN8e+aR7e9Gj
bpTlxwDUBOvOjHRgJpm/BV7ZV4yY00/H1RtuAtcC5KcqZsRR0HYrD580ikf2n+Vs
5NiLyJh6uZON0QUOaK3WugNrctKXeaSLGJ7jof0LvLzKmQjXuLpYFPULNKPhvYOC
9tgHhQ2LIo0OXctOULl9astiA6nPh2aw4BcHa4bwpX1E42+qdA1736jncaj0PBxD
h1oHoBhzvmTf3mXdhtjb0X15V50CN32ZR5i8nphlOgdp0/BimMj3V5OgOUSWkBNE
V3t19X3etaSjiQDPjB3ggu0psdKj9JzkHfHf+q0XstG59rUvYFOnIIKR3qh+IWao
lUM4JRMtP2DLqNs9k/1LmVtQ/YuyRYQfs0yjaDHOAQEK22EepstYoPVR9P78fSrz
ffavTTK7A5OLpBjw5jSyAJF5uJYUGn9JzhBMlz6TFyAWYkWP7BEeHGKa40ywiOg4
eefLqGZbjuRbcuCOrx9reYQJZiK+XORAmyaYZC0i6yUh41g0DxIZP1TNDwhCbE+V
HZTEXdsVtNxZA/7leIGGzqHAVEAn3Q2EQ5YLanSjbTnep6X/lUaqAPYPMcUKyQwG
h4zgJ4BOOIkpW7vqnOirkkH1pWtRQm7IlnYVXaSLH+U+izFWBYH4/Kvw8wDPORd4
CyWB5kY9q4QeWUFrGp1TDss5JHgsiL9ZFL12U7HqR2Qe1EoZToSj4S2drRbW1sZX
bppqXvF8XFRzJTnO04HdvuoF7jLMaa4ZcsEugab4QAmZmvP3oCtWe3DK/VlkRxVk
HlqsJgt61zWzmU/pMbreHAkmWQKMwXgCsAjxQaU7lVihWdn/Xm2a61spKH63I73I
Xni1HCbY/V/msiCzE9nf9K74ZtdkOWTdE9GyGg5HoGHTtLb0oP0Diq+f1l635CqE
xKan9AzmzDU7QAkryocXyYu3V+L1GIooVYsZmrVvLssofCfRMYQjpSKWP1/kLJWf
7yNhcqRuFlHGjztIt/2wiLc8+Fo5JAGUTceG+BNfCBibwKA7nfdZN4mME6AgWbMq
Af9mn/8xz/yFmJ4WiPneuB08qWYQeFTi0JIaiW6yKST4S4jcIR+7TcbwO98SwMq4
B+0dIqckFl0Aidl1TFpbKpW+ZcTkP8gW7Ca7NjWrnYl9G6NVoQswf+YWBGxovYKP
fpopCCPBbYzUujea03oiAkwVQPfkWedqpkQ36y4Z96wnpCL1jp6uXLB+sYpKmYaZ
+vZNRV8UMCBAHD6xTJ0b57248GmrK9DccSJygHCmGaYcVimam5/p7d7117qn7OJK
l9xwkWuUpwPve91CppTylb/wiCTtaKxrQlvaYmMUqxIhRKYHDW/t+ruSyPoSysGH
9phaO4X+t3wbHgCvbCB5NbJPDf8fn1PUtrxhridMddgOnwxmGIXjb5BjEYaRaoG1
Nj5FSMW6ZyR7YEhtwMkjDaL/2SMRir/g+HYYx2Hjnr1WjLy2eOgMZas3BdG7eqxZ
i0Sdr+fPv78r9lWvAILZ9ohxkZUUa3xIKpDWhiX3wPMH31j9mGIixpzkA5mUsdcW
zVk3Avc8Bb9GKwfFEsJZz30HmRaA5JXnN5ak6AKqjQxuKsSAXEkamRJbaEDLEMyx
3Xp6KOo5odRQC6DXFYl8vZTXHZI1T7B8IiLHr6X+L5AtluWgedbHxKbOr841PqTq
yP7rVaN1kN+64IBq26dukg5nKKjegpRST45KeamQctTDx6aQKiEapy1cwioMdwvT
gO0oCRifmOSQ91OrH7nEqo3vCaRVHBWLs88O77Wg+s9Lq9Gfnxi3dQys2/rEbVxC
FYv+IQX+EF5uydLFNY5d+rwApf/dkPOxLJtrd9m6+h/uvW/6POt9NMkAHLtTBK8x
vb5/S0Ma0aw99uhwXtL2SpMHizhpOq7a4CkXNwGC23PM/3h45NvBGwsOA4qc6WjF
O3peRzDJXhueCc6jPXTrRTFzjOgPhRLAlheau5/503YVLMi2u/PO/FKmjMFjWx5/
X+KiduKxqi/6gLmDKvAUNzsFK/l6w/7zQw+EsBdDRtIIqUf1lBnKSp0B6mEKBMzE
/WfAJ1y0bJwxChJO8EN031wNxtt3H1kFaSwyelt+U0DDqkrYx8JCfwfNPt7BboY6
8wVAE14NtuVSpv+eO9JRhqWAp808DQMHCd9EsHix/We1c44704sdYJyliiXbUMuM
3BB9dFSAH/wsIbHcFZAM7f14J25HmuyDAuIupQ/BtgSbCCX4JkhVvH+u6NynbxWx
YIWRu8dHrSOvuVpI08xpCA3vuM7gqK1qhx3qnluMS1CHh+t+tIbz9327B8SSCV63
/UjK7cNr54r/bR3guZoWiakFNFGr/WA6nV+UBQj1xrDh2znjHb6L/8bvMqwEU1wV
dbl0k07nthLehlxMT4zfulOZYHB45ynaj+B2Rl0xJ08xxG6qrd08ohsOSF5nWJYk
9E//+qB8BLPI5P6Dcep2rT/mkhlAIswsXLl+V+Xs3sUeFkDrpChsYxZ7PQuZ72Pd
YBeVo+UTk/Jc7s18yQjm0u221lg21QiF/YR1FvRq+afotXWFkkxeCaVFH1eVmxa+
bEDW1u4wAbMqBaZn486BaGLFZkWof1etTchfQV6jlYFYdaalOy4BdQNZ50wazyUj
zRn+4EMjUdIUBT0WyOwuqB7lbr3FacYGcgKFGy/IkuqbRTRh5jxlr1Yvpk7LQtIs
6XiFT1FCyJe4OpsqBl5ga5CfRVeZ1qPIwYq5PSDGAjLcgwPgt+4wl0287skLj6lA
V6dUZ73C8Guk5mqgISQpIxq7dN52UbVt6haJxbdOYZb9z9W57d9NlWIjpHgSHwjd
8DKI/VldBowzwlr9ORz7BIivIRv2eKdzlDafRS/1mQF2+YqrV6qJ4p5AfvrJpzf9
p55Xo//gpzNaDTb3bV0KVPUN313fYwvGYhCx0QIIdxQCWGOY3/iTNlzwma7BcrUt
YX/nk6youpn/w5xh8jcILRqb7F7OQ0KzGtsNf5ftwCFwkKthePafgsOWgHTGTxyo
qW33qXSVN3si+RTWBOHhIbX6J8CezkcjzxTBTWpfXRfLpiEnfu2rlIPsrDzvTci9
+DJQ8zMTxlHIpeY1H3AWqwCp5hYvNAwkaO/wnmYqXBVogwMVOUC46XBB2ypDdh6M
5C1bIid9/K+BxQZifib3n5S9wr2F3n/RDjqoXek3NTn4iG00dhLfl7c/Df9tGE7v
e8ZkXdJOjX5ukynPPBfin/UVrXumZ1Mr0LiMlvmnxCoGZEpIqCSJKdHepuDsR+mS
x+/2FCgxYL3B909h8M6/X75e4Vvstuefd8vd7pbn1ESXoMOv7/tA1fKTa7v6UaMm
GWg4wf2YAB5Sj2TlFWkADkS7TyA1+hCZYn1Gj0/gFnInLfCvXgtT+XKGsCAi0Yr+
9FDqAYTl6yZPSHnzXawupt1Um5dTDAgUI1L3PDub94bpxT+HTK3JC0xf7BE/SElN
BDXeHopt0cULg0WYPn7B0zHymuiEfHk+/rltaCn1ktSVdTz+fSQ4gdqYxzuE5NWe
KvUdConpN+Eq8Ql1OsWGebsFYW1ETYTbg2w11Zn6BQw+4/7WNhrNm621NWkYOPJ6
eQNIHdf8qyqY0E5Z8HVwtFP5XfOqzBnD5IOLpLrEKml6TDEbI3XJHm75BjPsCV1+
8gMTcEjPgwvW7X/YxZWt7FIyekv4o8+Ss03vrjz6ANRvIJtx7+hSG5CP29ATXxnI
UgzygHatu/DHlmExh/R1WyPPYW1O1fwRwkbIecLYMlSdfIXn9YgQqHFlXOD7j/ht
RUxdJruOnipanMKNQBdiUmenE7J+hVzsXWqrgNCbA+9xTwiCpclqdrGY+3+g0Qb9
P/d8+Qfqg8LJGYRd3jyHGbPOfoGfSIO/uqRPqQk0ucwDL5xOWqnrfybB2GYyBFXt
chEyEwTodPv9sl1n0hKl6mbw2W3JIltbt0FS423oqZkZkQVbjFp7r4xbAbi/er7h
42YNq5SFp25Ks9cFE8M7hVFz/qDt03Xa00BHbNESYU2bhPy/JHqnUTgSww1M8tPa
EDNt50Q5mZfqiOHlrjSfWF+u5jjOpKI+TCphbQvo+H8iAyKUwAGk/aRfAJBfuAMZ
zI6RUnuqli+q6YyRcPoAf2YlRvL4tQEIPv7By+YuRgthIrM7+lFysKg9trO2O74/
QxG3lXuDRoudYOjZb2Jy2s/R8gDqNuJyTJgDqK/dYPefJyLz6ZzWxVXi8JQ9ZA/x
b9QPVTZ9rpL+TfGCOjU9XpjVBZ5Y8+Rjb71nA5SEzMqFQlEUv6xfUO2mFeODssBz
f3SwI3lQwhT2qk0C9svCU+KnU20zIFgxKq9suBRWObybEPha09PXxbJj3+tk1wtt
iyc4gfxVKXpL2/RLlpu76JdYLaV8CMoRBzQCJJ5n8k/Dspi4207EGZ07FLOI8eqT
thKD/VbqqqMHAIEHVxxV+BSLjyM3XwHMP0wlQnpWoTKQtEMkQNe/HqiFQk3t9QYK
Wdngpiqh7BJYVGp9auBuDECm+K3vgkOeKC0dpN38gJ7cxk16OxLiGP0Ka/hibfjK
DLcwXb3hTou0mI/FYWc+WVcYpXhuJkyR7WlGXE9ttd0PH7L3yefoL1Nltj9hORx9
Ht2DJ1yUjnsV3G8NwV6HKs5Muq25itkRrJp3HJpBsbeZKhERwnyWoVzN5LSfXrr2
UEC1pT1pL4Dy/Sngr9bBdMCHcbvwEDnHYWR827+K7EM3tDTr41tbPOIIi2INgLZm
yeokDKfRJLC5Cpkr+XVOApb2T24SEEis7CBzjwhBG9b9DB5oSXIIOyIaj4NiVHSO
v2HewcmRK7/bWASUs6Cbwwzta5uvRYZrIJCaSXsx9E+bdaGWDLzMg8U4RmdUg21r
CQF9di5IiTN+59aLmrDaSIvdIbMBUgZ5UNPH83lzZxos7JPspeQLMeM8vM1imYae
Akg+RUj33Cm3sOcs6yS9RiZfpUBSL5Kl53OqeRztFB6y7w/QlYoiOqm5Qfh+RuSp
JglJtxsWeb7ObrsmuOTNV/ncflRLvI49D9A5oXkIcdktpfyuaQ/sOmpY5hM8i4S0
0iauD0XDkQwtUFE3MoUU4X5zdcn6rg3GZtj7hsaBSSxymYOmXsMvqimwYnOUSmec
TGXHhT4Mv42vhoI7UDUPO0P30ixqEDyVzt8l3x0zhAz95zdXmRQF2EMb35S3TPxO
FIttX0Imvfdbf4H9YKK8C5Fap6sN/zEJqQZOsMbUzeykltWZ7m40jrO708ePNQUW
80f+GV8VNcXB62nDoEUrQGmro3mj6+1ZtnH0RxuCTFfp+OI4XsfhiraMQZ9SPhpH
7a+VI/Ig9ROfbG+7Uy62aww16P4QdVjbpqmzPATbRgyklPDOOzAvveVwxYRty6Y3
K8LXGO/ISxQEGSTkGFKiVVAftysxtwOR2HfLOcafCuCwXoZA1F10T4nzpYyKiUKl
+rrRrjeHD0L4sofbMe7U86YUtEZ9kgdvTw1Hncv3pw7MoKDzB+QQTH4+e8CYaR2K
a0iuTJ5Oz7BPHgFW5Vy1He0EVCKWgdoNcBWLBqrxu6KmLGv4J/Vk0C+lzkt8kLUO
xsJbNWu6nYKeiQGeWk+LOFHY8qbNlMDfme9oVwgzpWRjX8Xe4n3xoav3SzgZxDkN
Nt2vwXlr4O4BlZQxpqTdziSoCgJL9aPCyQT+6jhP+5bcvPPmFDvO/EzEo9fOdqj0
8Rt0ICaNz7KaxkkAw8cyh6todIfnxDiDyBWP6w1Q/6Z0rbePn4af7BXxQ49OVzmS
vegj92Xsq3vdrf0fTPQ7N3/K0NqEbMD8fike7vHTK+WhJbz/z1JHDHGOvY1MRcqh
CIwEALrxuFDlvLUm/MYLqSMJVpNsRzTOdVwfFvUj5fWkPmG8Ml9MTG/eKFrgvB5b
yCL0r+HMNqz9xXzk4s4dlsmWFe7vupUCIjURlAkyUGihLln7KWNPQ+u4AWyXKcZY
z5r71A28HFAynQFriFKip25Vu29nMS5TImnv+IkelC1hsXRg0dTGPRSsbI68F0bF
nrCaHz1CfFNANAZRH9LT4ebu7U/CNV2JOIbC7NglncVKB6beqiSgce7oWVc76Pe6
6y70i0dXPGrH1rr1V2ojEqiR/Xy6g9FxPdR2VG5OpjwTCZskppDTEhfTVOzGGPrs
tnERZ27iJ/lhZgS9QFq/26B59nDDW30n9Fl3HLLR2jUcrfidHnDrjAfN4DArTWGz
7A4tPwpRztYGcDGJs3GCJp6GALKx/JN4VU6SFZAvZlqC7Hu+G0rZX6o6PN9IhcRj
9UxDKHIXnrU6xNabsc1haT+5F6YZI0JXhDKU1CDrhQnzbJwo73VCS52mbHGuV7NS
0FxqK5/GGxSD8SfbY4gDCy1+/bSNx0flaZCcoGJ8s7gG6pOky4iQa5WEen1F6sg6
Gri0b/cC2nogzzlNvazyJ3OLNqZDlNMbIPKhor5E2OKyR8noRNB6JJDlBIDlhcUk
GgF8rif2L/wkdWL/iyLKIBQdM8s3uoESM/jrCQAlzmbxlxSMk/8465lj1I6YVs6p
YFoyRTLC+g6X0VYp+h/o88WysOtUZb1J8Ef2+kyzs5vuOPa4XyUc7S7ZocpDeFJp
Y/mgQAuXfkTKtu4xcIvPG+q7VRKaVYF6wGE6MN5mx4mVZH5dfgk/kenmLv6RArxR
gSs+Lot01VP1uijsgMjofVkkq67zprs9kRdj12MqQSAnAY4cg+4iaAwVghdjCvtr
1qumd7W73BVXnThnM+v3N5EFx88cBBDdGRGCgwZ2RTBHytAl0G00ceOtVxAIthb6
ONTMIiifYL7YbY0OkE5IBFvwZ1vk8EUYVGsWBH93Gpbfmmp5krk7CajA2moTHAyl
8n8DEXRqMGLIDcZdavOrEy9fAsamB+nE/4adIINThS2ErIz/kriI1ieAZe64r+aw
/PHBQIOEjGeJRSZ+zgGmY1aeRq9zFKvP0AubJIRnWJ/sTckR0MoAIaISvNWNaNIt
N253eb8+Fz23f3vD5ISt+kzM4xcarkyMCbZBOXzfmgvHycevmyvQpRpCWqbbfovd
lQrgUjenUdds0dHpzUVlwYWKt+ON/DScg/BiBdasBskwC1RXB7GkuJc6z6LzMXSH
n1q/Hc7w5WN/4tLkGmspBitcPljtzu+NprWg3C6q4ZTbELZeFdViWhC4im+/HWux
vCwBpwSM7tXElXC7/U7n5waAaiorAm4k1PaM8JSdQnrRXaLpTiQVxcwtodA0B34G
qSqmzj2rq+FZGByy5g3+/cfrqfBgdK/NZHsHKVSnwd2eBNeZ0+sbt0lfploGrxOg
sN/sEr9vD8v0uL2ayw/WoEssAHOHbp8tNpCHL15IUq2Nq0fP1kfE6uAFkeCJ9q9Y
5SGGowVvI4dr5N/np3bGe7uep+ki4PEwMMetQjbfnGKZ3MAL5vymcJKplWjyxdlm
nmxVnpBT13SyB40vZCxUpagFGA1bJLgunXmtZluIuvIwxryQ4xSrJXfEgaP/Y/6o
wrkzAs9Zx4PF0KAMicA3gG1sxcuhC8YrCYugzcJl1C5QQjkfvCqjF/YwFhah99Qp
pBqW65PDW+rgFA4K8M6cQrDIMlw4J/DJCAh6IjcfMj50AQgwM93Me2z4vIkFzFxn
p7u41yLelYqXDoM61klZmlU3tmyDmdpFd7lvUqVetiKcYV4rqOdw9XDpEs86XOWM
5nbhN33sTG6u/XJoWRBmeoQQPGwsIOWlzSCkEojA3xO/HbDJaIdoFD28vd5pSqCs
fLXMmj8sEnGX8qSuJrjMzxRC0Xyi71rc4JE+IraaPxE0mKYzPyoDE5CG5sm72OjC
T0P+SFFjNZLgzuj1B6O5y+0zsM6qWcuYuGdO1nhhSymPaJ2K5mGrznKzZ8irJhby
j9wfAHawNekgNpk+qRlpruOFAunVfn3BmyMVpssJXTyJ4jSdTeOMzJWEYxw4AohI
DISDh9facS8p2uAMw9ZMkSTTM/MaebtCYWNC34PBLSS83gGt1eJTBZa3Llfp8nCO
IeOtaTSRvPcjjc+2Zhno9/+NiFSsNByGLttug4vOh6cOwNUyyGgVTNJ6IpYz3I8x
KaNjiui11Ddd1F21ihTsRXbDWWJl9wa5HQzu440ghPgx0abssH+GC1l4/fsKoXJA
sPdX6dGM7RXih3vav9Nvj0TlPOEDchxT5eM9+p/1GFGNkryWyMbq59LOdztIHC5p
QP+2g8oZBm25juWITRKuiKMAReXMu725+LFp6+PNOKEuz+xII7Zq4vLg/SUM8Hz2
PcymFL59NiUsAJWYvb4F9h1bNp+Lwdfa56To2w3NbB2HJI3lHDQXVagdB232SDDo
eULlqXW8J8Kgjy3THrDG0Yl0iji2QugAUYRb9132kXrIPAoWKZ71GEeAtAHGjVHo
6NENDKa9rDZC7kh31N7S+3rq6odtr+WywJCkvzAHnVaYREF8jxTodiaO3hzuNCej
K+WxfYaMfpe+EIzJxQBp371xrIsHjpKjGFuRouVXvmGgPZHwPEUv56h/gjqP/8Bf
BtfQevPviZPEvTQTkDorRcgeA0GtwVGvFuY0qfqv1ft2ug2Wc8IEUMekAzxWRs6c
WDu36VrjLY9GO8MF+nFxIMlw5P+UAv95GwjSBupFLJgTUfivruEWsk0PKLYYXvmF
TILBxYUOx0/hZlOsj5mBWoxqmbsrB1nhAzKeE/u0yy6tEq0gOL53beHxAiUz/Aem
zZTxYW18vzysAtsb/nFVtEmouE2/doxHAuaf8go+2S2Xnyqhr2I0QaUt3Y9HTTId
pNL/ECY0qAn9xO3oy1p7E3e8/tOhoZA20Y1g/Eb9aYxc3uKNNmYos6EJQTx8nzrI
JWsm+OwvP0W/IvGQktnKKof0265CZPJ3TraMdIYDvUH/UFgVXUsYLxPSWRr+VNyK
eNl8G2vBatpHKkist/DW+JbxKMi4/HQUmM+xfUPq1/T8cNtR2zlIEK95MmYhNHv4
TYdcl/4TN8lnVPMpBa4ChuS6UaUTLfMWxLn7BzLmyeMwiLFsfZRJoNrGvznm5ZFA
L/tFUmKVk+iAPUkwVTmdNVCYsBV4DOAhQthfDOAa2Y7EIxXBHu/zzKqXF+1N2MAf
L0WvFJ3avk6xRqWIOn1sr59ugooUyvA17B9+yJajQTVaIc5gdge5Jb7izCsxaSNb
nfw6xaGiGlP9xReKYF7AnJDS06J5Zf7vWww4hqTl625ie/WLKdu6BNXYZCKQxQUD
AESgzef5bJZ7tYDNBLmhwzROi5z4BQJbFfcLZujEkpG4877ziq6+8dqU4ELsadAj
KsH+HgH3N0yNuyJ4baiRWAHBgF8xVggNJTrLpVr6Io9luqdOgrU3mO4mPtV4hztf
crN2tYDdwtz4BUczmPkPueBGG0QMtauGnnieUaqdrivguVV9MCZs142kBVzkzdV6
46moiVTGuHsZLm9oqEc7DQvKk0aB2NUBMXUsretopsLv3i71lHJJe6EIa3avRPI6
WsLI8qJfmxGyv74yQl2lnOY/vtIqKaP3HV64FMYL0KWn2MU+0gMVfHmrKwq3NB8T
8s7TNLAY+XZJ+4iOuCK+RQsQfo0OIEb+7iRkNE0TzsupBiYarlpsbBCvMFN6q2zm
HgA+PVaXLJ3iOUrEl5lwzWENCfvjDBAatq2KiZ9/D3sWaYm1m5QQUJktR4aEM39S
MNBUIjJLw0ODys9/nWS5ijyvyBAVHr5yH47ftYmQT7PnrH8jaLzTiU250fNF0sW/
n2WeU1PNGeaYI1lbsH+Uh7NKtmPsfDxsybMRJcXzMQfrDsZN4rHoX49Sdtn5x3JB
HU+9cDM9Qbi9ndRMUAa5qGcMGgQIUhUjjtV58F4DEhuXjMjfjk4eFGa9GuviyHNs
mnchEN2WL35dEzrzHyE6Q/aAb530Z+Pm10KZXm4MYKTHcWVYtKRPHe05Rf9bpGdd
0jFPeQHWAV8ST1w2Q/CkaG08DteFfMgkXNJQ4Hgwx3hzEEtQFRidlFQPLsWifZAr
GqfRysVRMrJtTweC9/sQFzNy+SbIsy7afLhI3Hlq/oxnCpAWsUsM2JtZe63GY9D1
tY/jYsqL7xZIYEo3dlmHzSO5m/jZ7tAvoSPqhlM6/m7dLSVSQubRiaYkM1NpHsK1
1WgGbZHr+C27ZfHaXeQ5duSPfxWR9D3u8W0E0hwyKNN7mmXNAjZkebe84e4bCByZ
qU+4CGifX6F7dmfHNjJytfNHXvN0phTTbBvz7TaFdymLYc7bQppmkAYCr6UvMGhb
ubspYpBwKrQPosamJBGmbgEzGlLraa9VZDL62FJgOb02sj/qaW8XvD3D5UoKdiK0
WTcuWC1WoqtODvaOxyE9sEWZJuNBmsRfyH7a5lnxGL8WyqIugqo+f1OFky+NCHzR
aSRXxr2fkZQIbAgeZwx4xiLrK0SLJ9ROv7zYqV9LI730vcID/HN/FJxcMql612YL
yrzg3lKuvi5i+g1qImsmGWzEdzy/eFpAZ1MZaA21m5KNOpaE8TdrfvLdn23QNjc7
OYBoD2WYcIqDFoULetmxsiTuornDVI07ouMHsd0ZNBsObvVhK2S3sXtJbb2ZbUHw
OpqulW2oZ/BJ8IDN4CTr5MtPhADH/o3JgjCqbOlaN1At0V9wDB8crVXYBZFGyJeB
TMk83yunjH5YXCHzhC4ltUqoNVdo4ArVtBvcHNdsQ6lpach0l21ZY5B82wFCzB+/
XkB2ahujE8Kirhx7K4jCPNN6j4RQPGOwDWkuXLBF/nxNgfhji5G9f1FoRBJns7Yn
bSyUwD+C+MPZ3Z8y2LSQ77m3TwYCLBSIiEaATEONDgXgUHYg1TsOBy1fszj8poyW
oMxx9T4La4E3AuF/zJDGrYA82uJVt9VkaN1wiYh3aD7hhc7moFirsFVshjW4ir/Y
a9S9vMhFXLYP/AKXNGNTTcJ3JZM4Cxu3BEmTMgZJV1hLnHRLO/5xb5x+Uk6+GH14
JzR8fXRw7XuLAJ779p+Pjg3D6zNllV0vClOGN57d3dbq8PzEouoFdPDUVTQcg1G3
WkeUPgR4X3boWUnIwHKsrvQBqc/hKGfednMRKHg/Mav3gVnk0PBxDW/JCVcKrL/R
+0uWxgl7JjxcBpZUoHa0xo6MDOaqIYJFmPX55u/xypc6gL/5FQxitwrhE8QKUBHf
sc6Zdq8XO9+LB2xytrtRmAdbYiED90NR8jUT7k1zNGEyAq4lMsADq73qeF11bgwV
uQMYhcdF2mHDqi10/4FTSJ7epbn2KHVkC78BhABwkyRDxCiylWl+l90tEfmElkrr
z5AwjE0hpF0BTfVv7coE8TrpN5XTv2bfbX802zBE29RhJdlSeXjEDQFYAX5CRzUU
ub9Lqw9Sw8e2FS7i9G1vTSkbhOb2J3vAyWlkuIcUVGqegFXDoYEvcUZBh/HnoyTT
6cd08rGjA9pY7uAGneTNmNBVMrj/XpLLviXE/zJSFdZmTEZzyT8i5/Zlt+ouk6Ad
Wrs5XGuGH52pU7yBXRxvvN3uNyf2la7oYeXc4H/RqwYmkfNOt4Wf7aC7RQ166n7o
I2XsbqbujCzvDhmfyrX8KXC0ZyqYP0eTyuOr7HtSO9A9w6hFRfjEPwx/3j5JXwi3
FTOhO7HhXEhHeeWPFmTzflBV/a6bKWDbMR+TVsRyLW65NoDLpLTVhMExruCvbuVB
XjKOmMuoMYhecfeQq7e+2nZjC4J+7m8bJjIi3T6ndgTuPfIE0BtbREPdiawAC9di
ZwKRCoMgWJWpLlya33wimypGKDo0HujmLd8iCFr5dl+UIYIpoBbMee1adtdg2W4Y
LDfh6JfJ33Tsy0dDIVB8MIeVu/rryXv/uRD5ixopTFmc7KtNsX+SKRRicW7CaKtg
4al7pYIJy4vr0rD8YYG3Bcw+3E0mVi4+tNEKY+FtXscN+QmgqvscG8laHh6ZLF2z
wMDt7qvx989I5a+1QASdC6M6x+Zuh1DFh6BNZjeKmD09yrlngJI8YxXrBU2GDzwC
INHn3lgN0RnsQJVgCP2I/6N4vEozTaa3b29GvP7yR/YrYfxI8td31b+rmInIi5Y0
/46UeHVnk+2Cqx85OAYp+uusmfylLDdE1bT6N2FLwxSJZQD8enKvqY0uKLQbSsY9
+ePKP/AtpRAD6WqO4tWeN9bsxSJF6VsnIgjYcVMZTYJBlhOKjUuYGuTJj4+zSGJi
QARDfJLmd2py7j50dJx9I6Ceyo7I4V0wd+VQMgtMgIzg/8cZ4eAHMAI2gtt3SB1+
BoCdl/zM0riOSjryxodYs7lg2JiNjFRasamwQKJ4Bc6G/0YuMQUxGFfb6LRCScxO
SB+IMZgH2KM/2PdZWdOrju0QHkxO/mG83Lq8GE/jWEofhOqxtcFHGhlbuSIPeBjt
VQWwGVoD9e4xnPlildpN8DtUApGC1V+MseMhkct9z6PJ3VfMjr427YODpyypq6M1
2gGJqgY4U+48CzHowH6mOs2n0uPPWNJUoxqFqRTFvvE5bVEg44A0Gv3eBFwDGOH+
5FRn5RMzYeI0SGSD5PLgsGmhSKEdtsixCY9lXoyA9apkmuoAx+MrsJTC2W4iEOtd
viQIUmpkKHSd0mb3oYxGr8wXy8EFcFzKkV2Q6znw/M2r0fmYsEFi0ZQ629Z0FeAa
sAg5eR2gBEw+UoiFeDT9Nwj5DX/cheZxjo1lmHhArCpg8lpiHycGnrKg+Cz1/0qs
XSoHpar2qNZ7DyALIgmrsgFMMcjSDjG6lAqAznAC06Ia7r/8UhbyQRo8xGR0FFQX
FrKSR4AzcF7jXoVhyA09kO1lztRWQlMBdWfPFICzGKgqMXMt6l9JxJI5RjbuTLtP
xtGEPyIPkAXbZ+VJEkDLQorzrvYxL31sZMuI/jT89R7LdWYDlYzynaVMeKgGRGgx
yBNh02pFHiFqr0p7Diq/PjVuhaveT0BzmcW+mB+qG/fSzIKoOll5PIjJt57BRfms
GKW4Dis6oyg0S/XMln73+fw8HNBoGZrrqMdduZ1QPEnQWyu8ARcQVPZzdUNbzz1B
GcbVi9Hwe9CE/m0DGEAGFqVHoL3dE72AyjlJ1263X/068+sf8a777RbbegBt3sWv
oO9nSYOBOUQCjTsbzwDx5BSMyOoO+8tQPoFsGtLbYOw8xn84zX2Xpa/t+Ug+eGXV
dd+1pyuKnQ7bx20WRhTa2pk1m65bmi5BuBQqLhKP9YAS8udR45pd7wqTdCAJqD2t
AoweseX3/n+WAGUTfuQw+Al2xs0zfAwGL8yPwFbm7VZGQmP2oeWjSBtbukE0PqSh
z1Sk9/JoU5MWGsIcDdbHwJPNqlAVgl85OyQDsHuxySDdzJZTuQ79OVDbiCWpMn8s
BIfey4NXkhdxpCiJP2VFq5qyCzLVrAkZMLmLtN7ena8Ffw+BnYO+0Fe15NjOMWv2
W/B4E/Sjh9uEv3utyABsyfKac7V39trwMYTbpmQberTy5vcMMrz+7JWL5AYcoFFa
ZZ4aCMCmqIrgtQ9YkUZRNrkGpxYJMvMld4v1iR8n+lwusf2ohGFeV4r4agJx8Tdg
iDefrn5uq5J26E0KoYaBjA+1fgHKAL5SdKLBNEPFVw0byVWRa55P1zVD76Ypvcvp
4PYVeqa0cQzuqSImE4pIJOcteyrFR3UF1BePS50U3oymXpNtTITgYIy8H9IJyu/z
q883rpGvPUI0PQ9+vT/9TG6rBaYd4dVNx+25BbeFo7Ug8xQPVZNVh/gT/0hCdHBA
TFYQxuPPL/848Ka0GsArZtDSKPbVYipY89VDTnAXkRc+9rixsVmwCjF8dEgCECxx
9OET1psYaDbFLOUxUnR6DGizjTEiJG1e9+D4jB9CcWuH8E420y3UMeeeZZuGL2mY
tS3KYtvcaI78x95HjLoK7CmFoWyYr3mHk/mmfj3H1mE53gsout/k57lprqHjj6EV
uoJdF6S9Sgr24QNvWSyq1i6CsWmjrY5PwBpSGEhRPVb9ejQEEmCcuwHFSu+vR1rd
gXfVw4Rq18zxXZrEhDaFXPRaTNBfZKm2InpTQ5SJiXwKNa6i9BqKOQTT72gUd1tU
xX0vrlqZmXW2DOK6Kp31+Sv3aTfo8Bev1VBj9OWrSexby4skST6xb2FenpRb/Bgp
cbIYVHmVVUFISrSDIt+MMHWOfGcs30K01LZQRQ/SvlRout5asuZcU8HTi5WV4ehE
XfBwhcWKnL/o6ncNh0XXw0tpct9+Ju71cVNnmWU+iGNUalwdd7ZOEW7Np12VA3BW
9rbtLlZQ7XGHv7vAxs7SRPnSlYlW1mNjL9PsDLSN6v2hcNnnhUzzb8phgr0bfoZ4
PbgJKPUHwZFHMjaBtx9YjtLzXYUs/5YnFuzQNkpbz8UPyZAo7/CQqBxVOaJcQPSc
3Fp+Jjalb4jdSLfbAY7YaJ4/TORAZTXGVIgLlo0T/OFjo6e9OX2WgjlMI68wlEZ6
w7R9UBrOkTaQzVXHfeeD3n5mOhaFzJeE4w1LHT+u6wEBmnGj/FlKxTx02fbFanY1
BPzde2UuSfbk0MEeu9E0yiL4U6kYb5eM7dDN2UH/WEZuGiquDGrP8yFoIrolIjX/
ANwwLhrkeQG4IS9jIc9B6YfJRwyfyACBZq/4uZbDYcdiJVWEw3JycE6yLZzPhRPH
VMVmLE6zdsclEFr5eNNuW4DwtR0A7kmJmlNyNT7npa4OeCLti3/sf7hPrfp1GOEF
LmZF+GDdWQh7PWgmdAEtw2Xt/HHbv8DzftOQPVtKP3B5LJjm/ncaMOwfF42UKAtp
PbcVq3pfpKhcy1tQ4QNe7DkzNLuEDSw2b/ALp0hQUOypN01cjKXcPcEp/GIXIorc
+dsvidcnP6QBUQucuuUbDviSXgG4IfCZ6CctgueuB59k3WtM8kP8lnf/fMYOEy9c
keqGlk6upunf3dVOVzVCMtQBtCA4spBXofZr6WkqCYwSLyqoPjLk+z2jgUED9PDr
9QqYLwxpDyzYwp4ZY9oIBqxRmEu7pHvm+r+Zrvc0tZlrxVCXwRmjDMl3hcpB8Cp2
3DbJuRSj9bQx8LXQ2rW2/JrnRrgGtfYIRhX1owXJrU3ij+CEBVdD/Gd6zgpmTU3m
1/kxjizfEcjbIoNP/WnUWzo/bIPq1ODHlOXjyVeSCVhVcZBhqe7y1gBYoxQQnlcK
RAv+DzD4NHyLcMOsdCNGfODe5raLOWzMrQ9N/YERo1Ygg00wWgZ2sqAs109Ox95O
3sTXj0LSiM49IjWc2hAjdQAx/Plr3KrTfl3kNQiAKo20x68qXBKuSt5qHwPPa6vQ
EvixZt0yin6V63354a55ofPcopOEOlw4SGLMIUacUL0WPO/4k3F47M/9g74TAHQH
zdchsset77evX8DXk2KT4UKzHLo9LtG0d9T6u/eCqb2kr+YyN/QUnaRUTkx4OQIL
l+vG4PIiQSlRA//xMJzmJ0oRXRFIQhw3QEwhKQrlCFv20eNXUTXaxZQ9DdImz+VT
st++kKoxTEjPLseOOUtYBwR0HjXmTmugp8kmL0xb2gUwQACZSlKTaJa/TjZUhR1G
480Z3LDfB7FdJd4ITwloj49fWXO2z4B4PnKldYbGXiv1j3pHcylgLe+eDdGsdYJM
eK18z0drJH8U0hA8YwQYHnsvOd2WbswdA5dy2eulwMxc5UV5IdWEzoQg4Lm5XcIl
r6POYotLZa93TtwrseNrr9t42IMJDqC8WROJBWqa/ID+jPf8hjW7zFxBHyBByZnT
TaKzE21aF+BUOjizS1IlNSp89s6OdeROPQRM9Pj0oswPqeRcr2qxSigaIxjMv2L1
uYXGVdH5G3Y2CdL+zTTfuh1icReIWK2jqep33Hxdpnk1RtuTIu5GvYZ5CKfYrBtI
YanuIN1h5yjPn/VRR7ZE+l0RP4OAhnE+nLoiUlubpYsyjZ2eQezysp9XB5cdekoQ
oKo5BNrkZZh0gAmd5xX5BItllMAZYOmF7h5XKv/Tok0cjh6rS5Or+3H39w7XHdWG
bPNqrmHc/AeIbBca40bPNmsY+nOd1Gk7L5ayQxCytxKXua5LsmV14UDJhk34CZyJ
uYPBzEOB4OIoAeO9Y0d/2RlW5YiT+V+eUTzYQ4uYstsBH6zqsLiZcru6jAkhb81A
ouXrxA+FQ79hDmwrv8FX9lr/PCEcsvyMfDiE+e/whRKABCyrpPZGncLu3GGZkUxK
hiQvNdocA0SeWm6iFLT/OuQLG6OYvnjXy7Xh8+++SgKIs7+pg2kxJz7kWzcnhIZ6
rQIpM4SnbX5gJGfPDG8IQ/qA5sGc0GzsuPs2klIdiKWC/P4XL2F/i1tfaocXMebU
sdwJc8fGQvozy4s38oQXFVV2XYvTrQGcnBkq1QWOaFqLQwVdrHD5D8dGYnZBODpq
2uDu+uoS5cbs9fs4gZo/cc25fASZ5AQHqokikJXSK2UXn693WhKLkJCupvgAZvks
Mq6Siv8WleExz7bJ2FeQLlUE/eWqMBCv0rmGGqpCqye9GzHvPdocwlGmrdcW0UEo
/4XR7tUU5bqzZ9c8q49F3p/ecAFpk7Hs+SC4IZseNH5j5KQ0yS0cAWu/gYz3eTee
u00QWOL47ifcoa76Pxn+IshogsE84qlBh/oJOC9RfHqB+gOXnbBdjDhqx3hQdMbJ
i3Axx7V/UZIBmkL1X+ssALgF/3PfDcrjfzo6paW1SVqvsChehT5624FJIdbuMp9O
6peGllYawoa+psZ9ePNCgKu45kS6DFnVGB1XsMA92MiSEChGbvn10zOqFXl9DRdD
oTmz/FXKB6cryFpJMdu5+Exupq7Yedfy37CqAucNDRygKL32HXxIyOQYhhnUIlTu
JNQ4L4lmu4LTvVibBWaaEhgNFpK3xQ1F5Ac9Br6qLZvnjMAGrIaGbBlCkj42GwG/
eoAqWofrquqfosTkiyN5Xc2CMD+VBLUPuOUcUCoRVes8EeqtECCX9y58oXeVvlWc
HgAre0ssxISrU8tACqOfrJn2Tb7bDn+Cuk//cferwwJnAOqo25+WBSevC/Z14NZh
9W85Z1B6vEhRcNv8zPij8/zNF1NHsJRUHCxnSeQIjworJ6jW5vfJYFiq2KbClLtq
kNGsAwkICN9qT8jIhFVHv15Ofscg6lfOdEVYdTGc+OlMbqSBBilDCIIxQ4GRKhQ8
ypOgVdXLKPONs2k1QOJ1t1TSmdmo+4maNAFTog+1iCXtmLhSMws3tLquiqtQntIV
brLDk6O4ZpK7tFgCFhOH4UmOzYfItLh/nsjVh1HJwi77Z8f5+qcM/k/IyiPj/7HH
ZT48JZXYsIGRxhhRO9SCtO1Zp+Ujjf3O8Bu0TEb4eoNEcioxj0azZ5Wi/UIdkPPs
LsF+YLjQfnQgTyZCqX3/O+ixglMreB6RZwdcEB14nLJQywOkxjQITAL+tu5lpsQz
KrCBlwoDOLjxmq+McOT5HSBDpwXPPU2R0aSj+NRneUEXeLRfchdr68Qc6/J6D2OS
jfPpuu39kuo+z706sWkUckBqtaby+g9kmUEKUFlRUG/343PSPt4M3za+g2lXdekR
jEE0pp/MV200/MXqSpbubCaXbZrFj+UX+5J3qix+y+AgfJU6HDhn7Htj1dibqLI4
5FetuNLF+PeU6xow0QqQPpxgp/1Iymnc53kvQmKtizHFdiTAV00zzGVM/exAlBjZ
cadizHSZMIT76ERg9qNT4l3aNuPHbzWWwA1NjrfxZubl6nKGzDp47AN5PVYJF4xw
cOrZ9ixI+6VrP82oIopNaQ+zILexnIRPS72LlsBFaRynPT76UPJG6FAUC3ovan1e
osqMkUxmUSoKccC5zaYf8t7BRZTAhkYIwYUx4eK6haE2MnS6PSCb92N2zC9qkZx0
hJEkcxqJDtpWO0DrFyiPMQRSj64UmoyXxIQLWJ+vhbaLgmLZQgrzqAZ7Mww1GEuO
yO05WftycEb0lC9PDQVC/QObwsJLF7wwC15A11Ki0YT11aQg6ErRLNS3oXPEXOB+
qlM1QRuBhYbnMIZ+C6LdhKxg8wTJiwik0XQftGcXbq1OVPM8DhqV+KPBNPvHiY1M
RZ3op55+kxYmSHtZ0p3+VXaluuAq2wZdTtzFSt42C8H5su8mH/ZVaUscGfEwB5rf
aANt9uN7ounwo/n8UawVPXSzZ0o/oSDePQbrfP7U6TDTU2XAwLvjzpgVmskgM0vA
FqUXOuxT/lFNR/CmEPYqvupwTmHjQVC/S4IFKgA5/OzovC1SLbe7tnHBezvPHzdG
1Tr1YuwPwVn3q9U5dbpvW2kZK2XBRcjqyofgQZ+CfgSSC9t3CLThcE+QyOECaEZb
6CrCK/aoHsSWtB3CP7wnXQhUIFB1idCPoImYqBNTMYYBhCxCr/HzOWHzYlQqBT6Z
DnUEj1mMw1qwFtpRw/WRy/I4lzjr4pkWffUdldrJlxW/3IwdKmWcBH0v+6MlVGji
Z9tpQ12AyXH5xTtmZxbGTjI+CfqcRdTlVlGHl7vWnDmZXKijUt6pPdi2w3hFqZ21
eZIxoANPH9IO7QnQSggNNmHU7THX7PLaSv5SqZ3AkV6r/jPSYhA8CjBevA1XveDq
mnKJp9Pdit1/Bb7gvdLhEfRJiNCYacGPC5nM93uzKgCen4nmUWvE4LkNBECJDh7G
lbYn/RTdBkTLf1OUtyc0N5atLdCcbxZww+Q3UR1lrHkPjeMBjFwW1VrSayaKVJ0n
dnhRsn9Y7EvUvh7hIZQHsJc3Xh77XALOCZf+9trCtLvRqCEbpPZPuXPaiTxsH/Eg
IJoE6AvAmVK4QEl22FwbY5VNsm6iXFlhEgd+ndJWKlN+SFYyj3JkFsTKDL6Q8QbC
mIOXGmQ7fu09WT41w6rJ8VLKLo/I1ClyRvIIgxYQMIZ9ICyD+W605EPXKN7FAy15
B9FMWXHJrtCL9ZQP1YtnSpBOjOdfVwqCZiziZAtQGKVNSNiUl5zklCJiSKVjeqTr
OTiKmMeTlhqZxHzVuD6Bdl7LGTBLn7lpyTAN4v842yE/xKBmVGJ3SnuKL9cnxv1O
E/M30BcsI5oOQvNWmqUysdGp3+V2FGih7oiUZApMBG516gFAwnwvCR4Mm/8co+1K
8YiPfgPq1K/o3gd2RiVNReNCl2t+ssqdpogtDRFKbOBgLfonc0TY/zI+rwD4gwDM
rpOYP0QstdOORfyIZjgEyMrpozkhvTG+HrN3RZgkykLYckXazaHi+pG35C5fz2zl
be5G6MRfFxiFIcROPhaofbkk4UHCCj7rE1zJxxh/WKj1TBr23LVTskIZiSA1axuo
N51QMiUO11tlBD2wjj1oVCuqteBRJxsODnd4kO/Q9vo91B8WBmU8FfXGbU2/hjxN
i9hNouZdiJymql8xysslIB2zCrsH3/LlJyqmomu6ECBWErzBJZ/jd00U3La8NZJH
6Uj5vXAsi7yZUya5nATQlHA/1dQIGqFLvkiiLMO9inVHhbrwTcN8VVNEA70fjVEl
7UD8OGg7qrdxAVh9EVn7JSQBls874HTB0nvhxXvGq9q06dEfzrPLCMX9/PzC7+fa
cuoAbo/5urQfbw7t9m1P4Rgzx0t43isu5xA1+DkXijvq3TbLK17nNc9wBQMiDFAo
87uYqMhmqglBD3DwljuGvoz2WswS1S+t65U7KgQBmupfQVKgcLVb1u4tOQ5sLiE2
5CEfCM8ZAY0kjmB4sNxR68DWiLFYUxTlQVhbzHIPPSZnYGcTX9KBf15yBgNQRW+4
t6j8ikkYc3P6uCLhoSjqfHnvGcD+++Sunnagc/1Sq3S5syOuMFG350jMaW1SCs7T
tLMa6O/gUdp9iDxcIgJuYLpHhJ9iIlKLollI1ukaJ6k90Fgg4vQU38BBLxDWxSs5
12QDWWgsibEQJu4zEi6aiAq2zYW1eojESNk8kxRA6h894AneLfG9XUUW50YX0LWp
p+5D+Zww5he1aJUI6CZ9JsxHiZma13kXk4cxduCjMpWN3L8d7ay1IvIS9HrtmxU+
NCL2dI2Bk+cBsLNT+wHs4CdKpRR7FU0JfZDLsogVHwJFr4v516xrDClffF7qlc7R
3PIlWEx57MTFN4ZoS4L8KF29a25yhd/QfCoP55KN9wxP8Ohqgww+U+g/U0+gjEzR
34LXgb3evH/NVLMh3Q66Hziwi+gk3hTIRfqavGE3uI3cQanVOIV2EmFJ9aztCjxl
SiO+Rtl9JQe7W4h6lanQ/NIcnlRaiNAsCoWdlhybBtIthy7zvFoJa2zAOjzJN5U5
rkzn6WhsnzjYcOMK4gbP9VA+GUoSeLeI9JbxoaGhq5C4nMzsTELlePYDcgXksjYE
3CJAUjVx7OhLouDWrvfjAw9zCsd3jEzyShs/tDMR5ggjs0i9/SJ2/cPsf1YbM2T3
Qruo1sUNzF4SAHn8VdLX18B0WkPwhloImAqDxsvD44F8+z+8VBUL8vfSz2BU7tLE
DY1U1fJHe+oHN6ZAiAzONbYk6PY+BejNOULSzT5OAH+08KJq0MtDOsrmfzDHUTX4
yKhdtZPD/1RfFVzobuC6BMAdFgoSZl0lDH5BnWk/ARWbPdUfNQXopVUROIYtZnm6
AuzSSIWTJeuvAOEvcfzdMNHW4y4GgacGkcNExhBhHyjK5unbJq30HdSkzRE5OWAj
stwOppaLA7GWod8vCICZwXXhJBhNeyBRT84u/ZLmo2Z7msaw+ydTSVro/0t2povA
ynn5fUC/hxYCK9bRb6OdbtexWYLh7NfX2LiTiXOzdrUH/3eF+Ev4PaqGZ4sHJwe7
+EupLN4gDZmf3N0hOuhw1jQ1J77PdnmoOdrP8wZXlOEVVt/5jFB+R01AWlDDhk8H
vVQDq5pl3StTUSfxgWF9HyTQO4wpVgHjcKfLdTms6UWVmtK8qLtEzRIusvEV/GT1
jjZ16K3acF4o7RG63v+knJNxBnKAU87B8yGbtHboA7ygf+Ynv5HKZF6dJo4PHYWu
cI+kW+F7UtlekjSZ8Ai0TU036Z+tewYX2fncGRcvcSJOjCKcuDngKcx3zV4YfD3t
JHNQzyC2z7gDOKZFBSS7F2yZDIucJ4wpxZ8GgsYJlSxmHXzpnCwVrUeOUd7pJFYF
qEKDWns3ixSYVhivLwhE817HdlM/xZTymCJWUD640T2vnKwRtLSxT7hJ+9nWk0pY
K/RJJHBkejum6ModYFCKYHbwjLMU7mOxoU8nhmhsZJs6ZdgsQZ9WLMdEry8YO51c
gsqcJH+lvf5YoGka4rfURf4PbBHpDCcESzzkfc9SKrj+Nc+zt2nY0LwV8qNHrNHk
2YttjHiyNKZYzx03jqzP1Qr3PaFXbY61YXqkBBKE6gvJeyA2cuKuswWIhjti0S89
eOpRlKtOTJkHZh1jzl4iQlGiFzp2m6xYKSckz+oEikD8YRwGv7aKQU/wYo2vBoG0
9CgQ/YbXI1C2Xcz+wtaYZMQF3m9PA6mZakb0uuwyYkKkoGj96EbqG1xz4OI0oXU9
8dXjCAmtdckpaFVAj96Ma2nQm2SvR/n4Wa5tMH4fkIPu7y8AUPHBELYXuHgHo2Gv
fpDGozSBt5nD7bpnfULIaTU/arfevs3nl9exuHFDLP+QkMifWgtDZ9ZrQyKqaiXx
lqrdUQVPlvuT8SJ0P/wOZw8XLBSncVMeWrWp/LGUsbMIyDZNCEZ8MOvQJUw0FNn5
yx30kpAwF2h6ZX7nU8i+623eZle6obVGJdJgwV3ZKqOgI2B26kmBZ04K5PDnBpcM
qnKiUovthcDLKybID1nDQtDQlZ27bewxHD8UaYKCu6egcM3YBbdeFnt+TICILX4N
enoAnivuSW2J1zA5xiu5OuwngOfjJMYlVAyFzdaebsQj4IKpqW4PU4ICZu5IJEb9
e10zBT/XoG2zAPGAmQ0RCXt0fxnpUuvPXe/vQwnlWd5NrndUEPJcvgAE+ZL71lJS
9KN3zl8Ix19J7r0ecwychxJFW2ZDpbqyg9xiWIlQ2UWmhAGk43+j19VY3OkDAac/
q9jlQ3rUZ4xmF2KyqC6eCEuiG+u+g/EzexvCBeAhFIoTAw3V4Q+TAkO2Qx4vVUrX
FDCaWnmn18mByKIBKdbA73vErhsE+X21b0iaTTEyZR5h/z37Vx4oc2IS34rIP+a+
Vju7Q0bP4E9lumLeLm8xInKNmYRrQGQDLAOIXZDLCQ26kFNVlHIGvYkR6Dd/N8m5
vvjC8RuHhnQ+i6FSyQuMvNdiEgFVvkx8zd0mcLFg17Fgh0pAaS6/wPO7cnzHps+n
7d7jkOOoR7w637LaJJyrfZ0buJJlfdJ+Dfo95+L0vOs7nfbopMukCighpsmAPkeq
0ZFv2AJXSUxx5ktChyHT/XRSeXfkZ+fiC9rVrYvHkeZ7tIBU1E0K+IqVf2/Olp+F
wadGY/jlbK+Hb/aHq2dVB0hbfcbIyE+xfNsTgKUCfHSF6JBcmQPyvLcP6SftpIXd
gSYwM3bREaovWqb1NgtN3n+ne7DIMAG0Pyc0OKwBd/g1gwtf/U++IRF+fAtnL6F4
uR/3oCflKJdfC22Bc0Fz1xlGky1kFBZG6KyVGkbKFOQrVv6m1LIzr1rfmIAntOgu
W+GJmIWsI7D/CX7xqCMoLwz8n2i+GxdG3ZMbsb24pvzC46G/yNtbnIUqU/S3mxa7
ulcz8u8msK35sWqxiBfN2SG+OshVXAE9D4zT7HnRb5YM1qCmS/P6lbBHB9Wx33/p
IzOcafk8EEbSHWjqL2uy2gJCeQCQjDYMk0ZJ9wkGCtN/KxVMi+w8K8GPkpEhPzKT
ngRAO0OCZjJxlPXNlgKF0nWFC1tXXnfcBEntU6H6Kr3Kkt7nGlkR2sqfQ1h9d9ho
JgymbHiSRynUtadU+icgmBIvwdCfU4kyoxEKyVb1Rew5RZTGjmmu4KxNtjKgMf7I
OGAsqP5NcG/vPtLoCZUZH2SBWn9E/YhTUwoPWvY81L+W7EPOiTzy0EwVRG8upMfs
bjfSOx89tlRoLfqNq4DajfFRFuhValsjilAGr1Rw8YyP9bjBSICdTChzYAvbH6ts
+xD5Za7urb5cMA4hP8F/TuA1CaOQAM7aXO+aDFIfEwkXbOnA/L5/nd/G0WEJLQEO
k2JxUCTV6WvZwSoK02+d9g2y2RWHbt3y49aiCefNlzFb615ERrxqr0q0qYvp6EhJ
MxiSNDRqS3gtZqyW4JGwPhbWqHxIufFZX+6mRr/8H3gCdwLHjrIJ17wgEruePXLl
TTL6mXZ9gfiZMG+xKZO+BmysrhtqD27zx7YY0MZcjTs0HxMoX9yxFrqhgXrlSLB3
W0+7lNgMxEtUAcJ2J6iCy9xi+OUIspogOFJhJkV6hlytBdG3Er8p8J86w8Mbklkx
DIh9AGEoUIpFLppUa3MMa+xgQyV0D/mRkHq5fuBbE75g9YLOoaUqt9FNzImS2x4V
nACPP+F+WetXg7UQxHRcEe5amDl93AMmw9bNaLoDSwqgxB7cWcUVkBTmK2NLRtND
Oj2TiNUpdwB7oa++Kkq4jGlQmhE8E02LAFPh0ygczLvHJoHmprZO/mXxrr53uGAC
05rLgw9vR0FkwPbGf2Q5soqDWnrc0NlslXO/haUhLm9cZblZDXO9LVqpr13MDxUp
lQqEcrV/jBskrDthUuCslELSrROA2CVdLjQ4yStTGirOch208AJFL52Bq1BRi7U3
dc10EzQ02DBI+66hHhuCNcwC7kzqDIwrClP5NhtKAX8mlX0ZNsut4cpMgHLc+SUL
1knbhO5lAdCdcWDufU2sPWH43akCir4XzL5aeflbUECsqi96hlTHtnas6GodTs5o
8vbi55IV18s2CAdTe2qZSjaPkNYN/i1h9znqXuQIcNDmXQ/3/YeJgKomVxDwIc7q
ppvyFT3m4uwcxWu2qS0hh/RQYgpo1YLAGGv0d0Yo/OaWATPfQRxS4qR8TrCppM5N
q1RC4n9vzM/u61ePeut0ekLGaWvuMTv8x+h/Pg6EtrXHnL8i12y8JQU3QxjhNsy/
EhNoucHVVxDWT0VbSj18xenQjqcl67nuP4LuNqlAXsTSceh0nNBrM3qUW08aJeW4
PzMW1GpCRcVeiaP+MPb/vXaYwlMEdhXLEBXJrPRSxuonAAamo8y5jVEEbGAGijoh
xN4uIA7EL7wtQqe4xYifX+1/Fjv8hW/AcgUS52dBugdnkva+Od75H/1WutrHUjDK
WeIbfsvkhX6OSt802kU5MHg0zfnm6GkWgxTWfWgAHOdOS35vgzStA7BXepMe0Hcv
8nOJ4yhf291Y2yVpZeu9vstTjCWuR0UNUEQBEfYOTCV7elRPTIEj8VEO9ZyA8p4Q
ybymEThvSqlOtAa2ucB4GvrG0F5zyKSAUs81bOJIikY8lfoYqz13sDpZQkgVyFhp
k/4QdFS09z1HTwvaYAFAVe2KjEJlZzWf8WsWT/xsqnfvb18uaoghDmmYPj1mhmXz
4kdaBS8/S8+rbRVeEHaWcYo/H5CtcmDFFsC3nBZR7N6VdTq+pm/iedeB+CSX2GQm
+Nf1o1aQPlfNtjCNvWp0xJN4Km6FacofTb3EPGe1Sd9o7j9UVNPfrEUsaWskILyG
6CwQRYESIK8nmOm8PNcw9fGIS5BU4c1EfXo+2xXSPXHxB3OQ4L1qiTEFZ07Uw3Md
iGNB/uEvZnMgFfFmQbrwUWkV48UdhXW/vRivQu2BrTuB3NA5dqInEF8ECvKv6/ix
hj1s3nyJpATx7dTb9o5N3QiIUjFF1KHvyVbse1v984FGM3BWBe5t5uC9zO0WFhcC
cQMmjfGkPI4mM8cPYn+p+AdwrsNqKhPFAlUQaavYWA8y8kJ0bNX9PVa5WpKEUjno
0o8UTgzlf2OuR7dfegbmBgwtbTioCLOVQy2yA0DZnE5UHCB9OPWH1+tm5m3v9rDf
QEHb3uyvknP5o3EsQO1P9BaETPpyEQ+8T1jgIU+AIdZcs6fDVaLgzJkARbDgcUfs
D5qqpCpX+4RPRStHIs8z1uNYTubHEYdHf58KuIQJoWlemix8PGnYJXALQWocKytV
c/5VBNWmB8PnElBJ6wfXimSjt73Xi4Zn6Qq3UdTzqRtOP8uxxnPWcLPn8KoSlCKC
la5fxn22Z9YaekwyD/ptB2VG4cHdPxIggxd1C8jybRXt5FthUy2dj2XCvf6My66+
yYu2HGrndLOlvp421BAPUL8W072jwks5GtZqDVPsII0dHv13L+WARcanrPj0h2Jm
ypf1C0tOG0c+K09LXqVooW3c+DtBrYxZzslUxSEEKzBT/d5hTPqV1J/x8WFeSgoa
Jd2xhXXCJoOGHu/kjWBN3I5n9TZ/n0CuHH6frQbghT0mZX8IMXJ/Al+YTe3OPdDV
EY9/AgD7z1E3QiH0HWDvgiP2kRT8rtQuzYPU7IF5g0lTuYqOPFnESQ7aLmPpJ8LX
9B98ZxxlEdv3pxPBcNg+MQTdeBFmeGzyrMUbjQOIcFh6thAtRTHKJRAGW5E1r7eG
ZbDq2sjHgFyaI07R8EyKmCPe29wFIoh9Zc6qKVltYa81YjG+tobBwHqTQn7zgicS
tOeLwlsgj3r3JsJykDZ29lSiSuC4upkqVpeA1JUuuCQIGglLmZHMlz0EW0oH7gxx
TOdA0o7ugLgCsmrvYusegwHM1A6NpRSlXG8LEB/eQNZgbkkcCqZDaK2LhjQLrWoD
394AGf0aNoczpGVUtZ/VweNTTz72Qrkmcf0t1cdYPkgS+kYrDPexOxIBPEP8GMYw
QXMm18BAyv+EtuU5G+idy3BAaiYyAtLPcTU4x1seJ858ZAscDC6mkGE61WXw/LYu
DwrAyfHRQ7G4eff7bY7d9NS76eLjDLvxP3QslzgRG36QCLQRBFVWJjxfQ/mNhiDm
WC3J2HX8raknUdGSyqBfiJJGGSCXIYTnU+mt9Ap2ojoOZx0Sxj4CK9pzvfbWer4+
F2ttMn3VZRFw8wp32X+GnQ2j0u9RcKS63adVaq2nioLuDIt34hrqU4VPYVS8MAzr
9ClAUuZVW4dQcbURHgDuFywTBJqvINnHJVmuCYDAwNegOKfldpx48qxMq+XYNj0A
0ChSyPdMdoVlh9v7eBV44rxZZoQuKwxkezznamR7Y3I+caTvF1ToiWqgpuOyM0Sm
11NX9jNU6D+E4qzctXTpeRKizIdYxtLmC6ftuFjOSq5yHEWDEFFoziH/dil8kudT
d6ABiKDhXxW7IoMzSx83hr3wrhhX1PXrGTUYUBcgHYpFJwul7j+EMb0iqTh3Kq7F
p1Mb/J4vILn0VvDRc/7ObKbGjtLqtG5UbSuZe6C1pqcHMFik5anLiow3ucdGUPU2
LoyyVqvUuj8iVKme5oMehSmzwrNungtcGGrS2WdrWOzu0Du5k7R5eq2ywfV2A7+X
+rtIdJf+P1i9lgegsmZiJ8wNfX0lBwUm0BTYt6uEUzO8MGhSVCdqm5WgzIriFune
8jd+SCxqPT3KBmTo7be5KdYyLHSXHOJL/it3pUb0ODp8r9bdP3mBszNOEC9HZQ3U
6GdMiE5ohuU78LTI4/qVRAmYpAvN/kxejuGRjYvsDMS7wvJ1HYvrD45tfBYKPhlg
LFXrlcUVfXbis84k2hnrKk3EAAUZANzvVf4VyHr7vfTEl3sySdXOMcXg9w0XgXSd
CiFJCJxNRl21pFGFReZnUNzh6uwqG9tB0edvWVhx9Ct6bINbrTBgXCdgMmV3EA1D
UGzGOfqjs4pO9zUVVcfwBsUSr476u8IAxMkC/x96PxryEXpws1RoOoLP+62jD2eG
m38k9AJHgu//c2/ss4535B4+8ATpqofSb14SEiuxOpR+9P1hRz8xLToJ5meaOzVu
MvRCHzpAfoJGJNeZ+p8t7cmlGEXU7liTy69qB+6ApOibRecaWWnfUL4KoOYiBxj8
JT3+fEsiYWwGBAHpSScE1EbeV5jQH3TGl72pYbVTpOs0X1vIGUO00RE12GRIv1F1
CZitIncn7M4DDSUzIWmnDsOjCX2GNOYjRBaR7UqN3V1pHnfuEf+ka3NW3YqnzuP4
duZ9NcQuW7cC1RphHGKo5v/Xd91GKKkkYvK3TyK5djAMFh781tLMfUT9X3oFUdnI
idf2/x5CLkuEUdUSEzB0IWVmr74t32zydCtoEA3oRbBm05DXt9NxLvbWqXn1+N27
OhpiVRMeWqC8wz6iA9EzTyreSEOKSmAG2j66RuHjWTP2RrYjndbiPonRJKpR8P4q
eC39bXa89X2QShdqeZQ9ndZbCWDuVO3WgR94Sol6CmQFJGwvz329+jKqPIDo+yW7
aX3oDtu3Pu52HdGZWpD52nJUpy44Oy9h7vXKyInSMN53z48Forqz+wiOT6ilOOAk
MA9Xiv9lvf+PdQJxYfW77FUmsgo0WggIyMprSE340zLLxOlw4VBOhzH70lznxPjI
vab2CeJAZQwJcDKz37IFBmrFiMH4ZPkcNQFmOGyX1uLxm3i2HsWB2PfkurJ2k4w5
PMnxAV4q58LNusLqxWvXavMbRRWfQNWNFr7H8DySKLYvuEyOniTAUjkNZpwhpaPC
WWMHWGkXaZ/KJOahauuQKq6tZJrOc4gTN3nUo06DfIAtlR8Ot5G47YjS07B2dybk
meALJ5nE2x4XmoAflydVtlI/4YqVrqEpIDPoUGTBWwuHEeoBxbWJEVFjLT7BORb4
XiTTCTv5/vPDNJ1w5H2yO4UkZ3QYZbF1dBKOAniAovCI6GVnN7u7wKc4U5yXEmL4
+7Hyq4T5RD97JqxolGMGm+oWgCiyPfJKmtIPEvT1CXmzTEEsPxblm1XIy8+MGG+D
lg2CcST3MD9DRzAY4Eo/xNrjwyCbqtWTUV1lCI79ngjJXtCBPtSxJFGMT/Bn0+5i
4Cn/EcPpBHeihI5W3w6l7H8u7vmUaoWEHEk+UvIrRFOkAarkO/Q+YW4jzCszzg5Z
YwfJIfsdNOpEkIe6Ngrr1JPZNErI77gxJs6BALjjuKEYn/wbHEVBrIBOPamzx71V
9LiG0xXrZRdEgsh+WOb7UX9LrSiZizquPGxFizysQJUI4dANI+CzXTqWmebn1NBe
RbnNsqENd+DneKHgJ4hTMxwsfx8+hdeCYejd0uuUw90M5AmtQh5awAzLgw8V5RsI
+9pXUx7hlVBhhL9Wu5dKuBCdpgxMslLfQpS6iEpErYOD0k/t1DPfIhEeRDtu/P3u
Y2tpLadLi9DB6db2Ef7uPb6FYuNR4WzINdTQbZOZ8S06WqyjeMxk5bJU4wvUhLv0
RCtl5b4xVU9paVmMzMcubwlgVRBbk0I91AsQ8LGQFXfNGdqHXfCxZ+k8sJHvDQOL
QTUfnhnwMdsELhvfLbMn0B2BFlg2GmBrp+vSCxNddeOym0DkkSNSQ/7SA+uouH9B
HBzl7/pso7vu11CHxXrcK5+wC+0ayJnh+slIR+l23C75jyQLaYyht2PpQg2Q+nUr
02S6T8lBIgNhIWgEUN/bQambCnX2hvZjR5n8kllX51FABR4O6vnOoNiR7Yw8ECrn
RZ9r+Uzh8kfSZv238tDHG6/gXtZiiqc5m5DNrKLzt+s3i6HuTNu1j2SWlY2vL3fe
ZnOjgvp78hdtMxHMXbiZQ3LY5uB2kDjbzoitom/EE24DoNcGHX7zBJPJDmWK3LPq
NRuP4lNj9ZWvsNsxwULtMioionFV1Yq/V3F9967nKfJOng53eHIaeal/5wrmVQtL
llfbOBZuwR7Ro9lbgssnuZiRfAcxfjIQD+vlsdrMwpvXznE78ZDC1459dpH9oWt9
65L6ofkBGm/6/B/s1amW+wgRNeGME1jePV+ba0Hhb6craVS7o1l6qocuFRfsW/5c
52+/OHDM/mLszuCmACv6ZaBguFoydKCVKuvfkfz2ZIvbr3fw+Ztg/ccAidTZWvkE
uE2DZ66sMeTsQW/RXjg7TukPaxNJbxEoQV+L0aq7lazelhDS+/fLtJEcmkkH4Hm1
z0tf8fJsxxA59ffF83ynUxFqhwh6XK5SDnWtCyLltOnped8lsEIMhBjrJKcv6Yns
7cBkAln6unMHV6uiQivevyRdO4NouR8ThCVIiC3zS17Hq9Fj9yXnICm0GGtLzXzP
ZvYKhYWI+BvYe611HkHrML8l2Lhc3aXoHK1r+gzjXHF7zPgQVY067t/vMO18y1jT
/RUUKLJxK5okr15hnZMk21hP/E0IFcxxWzfsXTGqwqQmeb7EWr3tSQlkS03752wE
gQ/KNdQmiVU/aL28Qyn8ykCs4YDsIU4sdM2aAQ4J/wzN8KNTw5zfxgZyRvyY/wnf
Eaubrwk+zqB61q6BlYdgQVemKJLvExSYq9cZ2uvw8UBJBFaBThV6jJIs+DpOx/wf
kidmSP6Tmlj8UbyOVwFLLhXu39cPT15FDILGe5lp3oYV1YLPpk2tQ+82DGOP/8Tg
M9DdDshMUs+vzkQKxQhNeTRktOTFjDDqZP5pftm5d7F4XqBuX4tnN6Ra7JUtIo7j
anF+mO4d7tqA3P/tQieAefeg4Ctkl+8IIfmvnagZUryNWYymXMzG/v2sSBDbhoUR
QQG/bTojxNIBv7p2K2xXddeX+kc6hnMwZSDFbUGwOwnrX8n230lQv4W3xs8FJ6hm
e6Hdq4h2D3t60VFFPTywBgAeOn8ggVUqRCamTRv5nUvnueoVMMF9RwH6Tx8XoKbB
m5d1aFGBsJJNdfHflo6daZ//UI3twaDXyQGQ/mDFLHILOUvlkvz3SKYuAn6GRRMD
OtWIazXgK58qyIL7w52ztX+XoIMfvIDs7CIJk4iZF1EWwen6gRlksLUVKquwU1Nw
nXlZ3O9ucCuWVEQRfO35/ox301z5O1BqvQfS7C11Uyp+s9q7jpih5hruZWZTtg0t
7kFyPYEBN7WLtK+DdY9GM+S7tqGRDZiXi7kT0BUhttnON4PV3r9NbIbvnXOodPwL
AktnZCPCc+8pdwwvsAvGDUXggl6Zx5LgeisEwwxv2bSZyW54sBUZe2ma8p5lh2eu
usAQA239juSrTqE5pNWRjN4SM83DcLVCY61qtienKJONcXmMpZE45Erxi/0CR3tq
PZhN5eOhIbxsfnsfgSh7xmLPX628oeEzmwMBmSb3iXbRI9c1N7UhUlSO6PFD+nGm
Eg5ICgvEtZ6qWerg3q0woz6j8VJYnkvU5/uJnSZt6CnaxKSM9FrWPPoDbhrSf/6I
1tUyqeXZYnfOQ7NBfyBw3Z9GbkkunyopcRI6mdsWTxqlrzGyVfV6WvoFy6cF6Gse
WSEOYXGkhjPpsD1anRUzDuwd88f2DaAn+AhQe7M+nxba/OTW9oZ2I9E7W3XA/cMC
kv+zRhmR8rXbYPIuOe2jylHnKeLOEtEcX/OhWpBnwdYJYIorBWnpGkplpMUN8SYh
X7rfUQagxcVbIOff+5ROrqdHiNDwQUK39g3aZ0+SLzoJ6yptpGmLbatWoC8U1itz
WhPFcAhuKKK+wYj3Uz008GIdSCTGaFLoSHReHEo6iRf6Qxr5bUwmVx9/lOPTUBSX
xFrzwk1IAHOWu8Lxo0tDAp7hdzQzj1416pDL4Irzk4bnomRR3+f4hDU+MFBZWpQJ
w6691Volbj6mo756NMHahXIH/irOF4H0xEQ2NQZWjLI+oW9RdFYu/hqBUWAamkan
u7mVJbAgW/zr4I+n42kWC47/BEtxXtuTvoaxthldaaRRK3sydTMwtG6fE2Wg11X2
3+T7HbAzQrc8Eor3a6ad3LagHOzkNJ1l+hSHA9ZREpn5dMhSlOv6HDzgiTFhSwPY
YT8OCIOxCUDdCzMmBVFNJMrJUIVOQVtu2goVuyXQKAhqVyfgU5ZdnIDzgqwj4IEA
GwHyTL+mpgDBnJnFyyhrQaZtFzZCcmD8u6PrpKk/mnqlZW8ZXDmm33UXxnlF1KwW
dntafqHd9+KBIt8nCtrZomn32cwkv4fzzgzUsDGOUBOfB4X3ahDi7CZassVYK2Lu
lGnsJIo0uNoy2RucUH6H98rt1A13r8Wc6Gnd7eWKiVFHRnBY/6UllAmLx72zfqe2
WWDnqgEdV4pp+FEHSJ4DcUBOI2yNajjQgwJMHJx46e0ncEfbg+K0anX7yv20Hr+X
jZjzI2dmuio51tJ8V8vqrwhans5NFMUneNdetOSBR26iLCFjSfcQsCjMHhUnJZB0
diSHR1TNH3CLfOF+S1zlLtAGbnXp9LxJByXxlv1ga3ILDkCutqL0jeHRlFmnnwJ1
C2ONC3sMzFXKtnFkNS3ywNEzHVdqJGyQ0qgjBlh/wwH0NDd8U3GqTJgppcFSP6AH
NmVRXnz0ix1EgFbnIuKuFtpMYRnjyALRsCsq7wliSMoOmsUy5776BIgrfJiN5QYg
KSnm+g8ccxyfcc1miDdnHhrhSt4u0ZC4Fn+5KZD+Hq/X6eC0BGcYvhWoLa/UziwL
YAQoI5B49s0kCQSZqxRsYzuFUkvKOVBH8HYlvTLD1aa0tMFoKVgoAi5eIqqhfMme
Cp1Q9R8naIJFqQH7npaM7Um6VOSmekAaCDVTaFu0o/BfiRF+32zhNFrpBA2hx7QI
C373xVSRndFcRJlUnQ14cOcuUvyUE81eWZcy7YvWpBDlHw+6CneCeP3JOMmCEYwr
Sdqy+Q02fqnoSNI/LtLvaXuUpecE70Lr9U6DQ9m+mARVIfbfJi0gxlBTOv6bSByt
hE2pHij+N63z1HcoijVWBCPXBG0VEShoRVRNZqVPbzBeP9DsJaQBaDjfYXYyWpsO
i23rgY7WzxnF2Ty4zxbZu3/N9uz1QPzUAGkZPlYgR0DdnI1ZHzfxXhDCFkXgwwsP
+pQ+9xty9nA6bZ3cCGG9N7/q+y66o3B7eO1fYEQdWumLivTzq1yQUczrgG2hKvc/
4qqNgiFmONuycOxbU1Ad+xrxuQd0E1AdYS+ri1VukjdPiyfyc01Tf5mTnK/CCqu4
iw9KTnXjt1xrHponrTWWZGq/HPK8GrYRa4zhyOnVPKJMgGJrjDDnZpB3eY2FpgMX
eTJ/nXstO9bzkXm5hFtsw3MjQqWsqUuXQ/jAnhaJyxWFF9TqoeyIC7i7P4OLWgD2
TF+0DnWZtvQBs4059gxlhNrc4fOM2i08QN5yro1X1IV1iNQyKQkye31FLcT+gTfW
AKavpUdV2ieF+PIMOTpQ3Crq6LKrWf909jpOssTwQ0HbEmj5vVyzHrjH+d8ESiha
1vjcrreHBMm0QRMbpAOFK9/abePrneZV/i+qY4u3bM0h/FLjd0JJRfgQzEtUWzau
4sWktZSeImwMYPcYtgplW6aGkIOCkQwS6V94CjCUQcnQItfE15j2YTe4UV0OgQql
0lu08EtTLhQL/FQXOUrh1ZBH5U1ZBKsyowZpQ2Fq8DsexeyLCdWqdiZ9KiBln8KS
dFUbG2VwulLf+k1GINnAvAaXoDAF25daGDtD3Yj+1reVJ0nOuo7cXB3ispx+FUM5
8J3i/W62LeyRLIBeDUzrPMo8LJXXUN9a7ecysl1KLL/11jqHJrrxZDNdqIk4RZOs
wIlQbcEVBY13OTHkbUfyTqKwZdF0v9jje2dbErr+E+UHuUCEFn8g/taBLNwn58NW
66UV6wm2S3WpHlGLRb8nGN/Fsn1nDw6atUg2AoyyYRDfVeeMh84WDM8kQX2J9Iia
7tMNbDfMjyv0WocncF3I/8QvvLnItchiyMvLA8WxtJCEBBSF9e9C6nX/fqaO/lwr
iZaSxi8o55NGAqtEWwQ11DNHGIXLW37GekAEeJRw6r9C8Fwu0TgbqjWk4s8Y47Iz
GcYDCfzLX1O/OPjxl4N/lWMrHnBB9o4Tc0fwVyMcXi9CpoaN1n6pnjh1qhcwvqii
qoDf1GfhwFsF1VTOhwywvdXIYW0I15qFr22jvKIb2P9PsVtm76zfHLqmNQn50dqH
0wBOkdoOjGEAxyj14NL+AJ791WV6wGl03h9FZAuggMpTZhI8fx+sb79oW2QtNcNb
pn6ZIT9f0yUuDZIr8vlLTMJFDJQviQDb+U7ZshiLNtvvrq0tvRlxbnKNykA5Tk0J
3iUbE6Yl8c0n6PxLy/WKFYBs10uB/a2TLJ+pLhb6cDT8rIGHJselTQjzpNs+JIRw
DLNaUyhlj5vmrD2lg7KOJeYhPOTXPI3jYHiXTgSbx5sgc2i4cgbguqRuC6950C3j
XF88hA0yfdpVKI5oZEnBrB5LmSVdcmVtEEkaV6IUA98GLindXeUjNJOomhgR0E0i
WS3jpnf60eDj0NruOQj8F982L9LaweMzw2fSIy1ugzpBEL/oBCVe4lnYO5PJanV4
zwutO13sRq6zagM/EJrzgfTy/BnbOgUbCW22IoC61iFH8MjxWlB+R96iSw7mfcH7
eGheYOpcZNB93kUyz1PX842jLGI1MiM1nnc1CSbNYnGmyUMI/tH513vBQe4abubr
uxAcLgHM/FS5JZqBaub1azzyoJI7R77iXND85+D0gRk6IpaWm83A7m2mlnoU22j7
9byjvVcaPLKK2hD3fnM1BuarAe3pHG3+ut21YaBP8jQmAA1IDDoOX7LVLV7M6AXx
HUWpnbMxlYybjOV5wXBRJV+FbjlvGfAan6mHisYi1ZP4qv2V8vuGdmjkdPaX+hft
SI/QISR6ugPSryTiZ4PsqCYz9cqqOTOxxGG5/myad1mblXxHLZj3h0f4BO4bmOks
PKfj/yKsAYB6mtOEG3G7XC9oQSHcFsv7QM+89KJ7E7M2c/N4yiB/O+sjtiRcwpPK
gHUr7RGhklmiO2mwDPfZ6nWYaPM1nMUZU8j3BwAboOyResgzI/+jES8ejPADo/Cc
okivgpCJMuUkUJlyYOB3OUkO5SqxQ8yhcGzNlbIjrxH/je+uTggNUFoU8DMbxjFm
tY/TKsMPZI1X33kl35UFJsOr/X8l+odQR5IM4GSDPHhqt0Vr1J4NitcUTvoU5oJy
GU1NtwZkoIYj9+dpMN/mapgMUjY//ojQklWDY0StXWLF5N0f5OEBHgfEeCfhXLOw
ag3unTJVrSbILE1QM8Gmsi6hSFymKlv5S4t+BUsYZVYPiqelwZAUZ29ShkaHoirE
gXwvOTCk67DktxsAmEiq3odqccg96eX6wqvIIoxn0V/L4rM0kH9MnmUrIHXbf4wH
2giAWxlHwKgZcILizEoOGKZbSTKqvU7bu7MhAeee//KCJRI6siCoL+apP/ikhuQZ
5hmX2Ax5CsaUEIvNEwJ1HoJ+MZKdjZllEFZW9fleo5J9m8edhfdBSCWJOkeRfNiP
czvm4AeAQSFVjoXp4z/bM2xhikIhYmYUJhZjYbDosX54zQUgVauvpMGQY6R9gdfO
JtWsDBKC3txhEee0/O3+K0GFFtvnzOiuHYSI+OgKcMd/ilgkDp52O0faKcxj1yrN
bN4AwRg7O91q66MEIGQz2/+GVH7hNOQdfwDRsK1X6cnsIjDLyGYBfyA7P4uX0VUI
wll0FbSqEbFN/99L0eY4r1rUyWktK2LRtjBgFYTxbSLb69Yzhww75ieVZveWwy4S
fWmNZvWPNrvZVqqvfpxEokWlUDB8gNmpW+X01JcwFXTdcyxfA7HMkYYSd4LGfQ+q
Z8kbHz6DFJzQELqQ0ohvwpe74HJ+/zJ/gTzWaXg4vd8H6/k8K3V8/t3qz9piSNFF
mzS5HaxAi3t0Egwo+pij6ch6AontBGFsH8atc2HgmmQvcFS3KxOTryPp1vUEAPR9
saFZW7r/Cay5E9284cbrdn32piiP1G1GnSA5TIB3tdpDZFkpSUuoybmrJkcubyAB
dOPnh0cInGPnd1vWYv2DivEaN8HSIwtJPXDF3pdaMhogKzHyTCkIa3QY2ayFyjSC
ZwsS4+OgP68zRubXETec0KDrCzruvs1s9reWZ7dJaLjX3AZuz2r1FM1r1NXHhtOp
u82Z6ARpGe4qepqHOepAij5zjtTuEJ5PR8e0se8zpI57DP58CXhKY5nNNCstQpR7
FOJnUzF9urOvLBA1HKsJxWO4lZAI1rF1S+R0XtF7BMo8vy2tkbQtjmoV7yvd0/HK
nMOPZsBsdtMvcFAext9pjrXxaT4rZWHFsqBE/IacsaStk5PFhxuuDnfO98KhgOfJ
ibBy4yKu9OQ7W3twOobRGZyZz4wHu7OpN+SdJTjnL2CRpultpdpEhW2EHmrBsUpl
C24dRtJtXxQ7Vk71mtFZjZxCvd/6Jd19kvCo0Womzi18Ws7NRj62D4du5bFBk+VH
llOjbTWLQFDOF9UlG9WH8nXtlV5luW5N4lTujw9W941+VPoF1RbMc85Mq0KpACQP
Y4GcvfkZSEgROP3uakhiEVfrRcm+5kBfBuQEbsfymw89gy4qMVGZ+be3RHmqfBtF
dNCgqTaZ7p+E5KjcXRxpXHfMOW2vwHEgIrkcNuTv8i3we8VFDExCBVsxH/I1+R8D
nKqkwpFRN/11Ju3rKTg2xyqVsFNHskJlOFC+jxaT6v8S2v2c6wmtFIng1dzeBIRN
nuZ+AVgtBX3wJ6fcka7w0Wrz76Mc38zkLEbsJy4sB/9JV7adrPGaBZODZNysUiR4
cgjSfs8ptdEBoheqhGH/Ql1BJEgfa+zHGuq4YnHhNNgupc8VmxR1Yaadj2I/CDQ/
lAlZopNllqLJixmaczo6LQ5xObM56AtmIIp9Z3tot8SdTlW5Iuqs9YWuYMbM/dql
QdkhuQ+TEnfirZIZ9nPQ54a84pOUH1zHQyijXskaKTG7Ih2M6vQY0gcMcEp0m9um
29EleoI9FNtbUFoRT6Oha41xs3A3xRu+QGqSHCmwfE6roAhesWm3YF0bTf/23uxU
e0jpdNXaZ3ciNfptKZp9xc2/9lJFozxrGFnBuo22ivsx1fBvJCNcE1EHzal/1jod
31xFgeFALuU6okwVf3ThU9ipRWE3NUGSC784kuQN9UcONU+jz/a5VVz2n7uumSQv
lfxZFvoiU/UwueXlgS/lorr8F0BInltspxkeZVLZUofgc7w0YhSAv0IR9jjDGwIA
frH1mWHFU0Xcgi5FO06kZrshbN9qvzCuufSS8ZklO69nrcAAR6S67LPm5ZUXoM6s
F2c7zT8NZ61Ch1XlhnEkw/QM1zP7Sn6zim/9LKtPI3b6PqgZAzxcMLgC3OUZAPYC
mgDpJ8vxhysX2VdbEWrKCHttUYvySPPyJ1a8DoOtv8PY92KhfPU8GRFyoYHmDIYT
ui7D7WQyY/W4y/CHB+QIfoyBZe+g8RsicE+L7TdwcfUAQ3ytKC94mfuItSCFD5Hz
HWqomiN6THmTHKte94FXg7bA1ePNlBLei5Q2Zq/wSMD/MI938XXY+44Jf1i0jDLN
rVoZ0z4dqVDj8QsIe7feUFfiLR0gdXDnXLz36WdoFHnxGDxNZKEOzK1ZYFMAwMP7
QIBu/cBlysp2HVgmyLQtWMr+YzF4LsrDlO4jNJC3yLGLSu9M6JtHRQSnsubAn+pb
IZAmwneTJeThEwStaZz1Cyf/P0ByGGqgvfhv9gFfNUkIdZHDxgcmk9gHCBxEjbhz
uWfqETOQAtG2/IIOlOkLmrwnI2f/pc09fiVcp0RaKYVlBcczH5I38KOfmpOfH7sE
uQqH6BhxYy2LIOBeaEoInxql7gkqCVKPimQ2c5S/QSJy4oCBqFsUf8ZWyNAwEkL3
WmDEhu9vvTMQpeZk6jmOYu+Chk0PXqoMFN3hhL3hiTonst9d3lLdK6h0MiCXI0o4
jbj4nQni9Ds/F+I8SRe0KeIkos+GS8o14d+BCXe7aEjH035H15NL+7XO2ATNOmlm
NtInfTX6EOMcKqToat20mj2wz4R9zd6/48sjnsNlIiEcTFM+cw0KQ05Mf/OfZg58
AJpvFTZNiSRgX+oZm8DvUU9aaj3cLADkoN7htYvE2xR3y8s9JRp0f97f4o5/FBBD
CZGcRl6PyvdRpgeyKyqRhs2jGMFctbhe3m6lhJULvZlWmIM4Zy60kKsc/dyOoyvk
nBFrFn1JbPztAezUi3lFOJN78i0LMy5LFL49dnEobrcJbZ8kGVkaXiJI88G/f5ut
7UAaXBlV1bd46rIOTkGnrdiNC3jpW6nE9gP7XAIxsq/Iab/qyZ1E1qCZpleMs9Qc
5a/Wlc4Zg3vWnnKsmudL7p/s/jlsGOqs1mfvahdtkFJoL54VjOWojgZEPUFHCXXD
s1+ROo+7JAgJ9cE/VkrQW7M3ReVhcm1jo7rz53WxrF3Oi4Nj33FP8nSC5H81PgNX
s3y+BfEVcDW3TgWfRGRVdBwStHNUGieDdIdMs1ErJTRRZ93v6bpuEq66u6zgEztR
SdM8NxuJ0j30zMP8mxBQs9IQ0YLuJEYWykJlDLCwF9h7tXK/BwbDQl93ojztnmjg
38NnGqQfHE/oI+KQ3QdyHcFQsIB4SyvjhGQ02ewl+S1THlg/Q8wB0eLezwZ/496p
1c8/yYtc3N3nPmiQomBvCbKh+UsH1IkJ7s9eT0y8qYDL/9jO9dkjDSmC33OYTkui
NiHW4izkkwez8oXX7X59iKT30J2kfdfr37IAHO9qoJuW/r1DWv2Wq19bXzBVr97u
UAZaJ9iQGpbx9HQ80ZWeVWz9tjLmtuwswRYhnudYRXoRH8KxDWt8nGFFO+QQKJ4z
nVumBfzIYDOpahORjjwhzpbDjqHGOlw5EW6JzK3XAFdK/8iKHBZKrCiJ+Huf4A91
UKwzXESgFFsrFshMPRiOTFY8dHmhcfQ0zzjvmQOiPssJOlnWv+wJImp4ZE/IBdKx
JunGS6OBuIbWFb7hQot05PW7dKkkxR2Un1SWZZ1YIbBBNGoZSpLDuTx4+tRXvcC1
FcbqJK3i/hYHHAw5uumCFJACkneVLQKhBVCYeHu1+bBUagfMWq3oDEjQ2DMLMheA
S0I1BFhlZKibvNDJSUoBC6HHUnGXN8aa/xiLYDrW/S+abP1U+2j9oZ6/0m0z47Bc
q/Vk96Q5CfALUFesvAjo4LQQR0WbZIRDkIJZgRVc/3LoT2uG4dTfzUy2coAWB7c7
92OTXwnYZHFm2VPgIfUbnGql0k7G8Cgw7q2wtVLCMB1Ii69Ish184g35HfVnlBnM
P2a96P0qNY1xpRU5iN+Fse09csjkQe+cshZlq4e7oQCQCGxLUABIv0fArhViN6u4
6zPaC7EDoLRpqcW8m6Rb7rlu8NaL7A2VgzXQWxF3cANd9rC1s/gG8Gz7g5Zhh/ul
dvIOAPNaRKiqRBBQ17tEEkk2N06yYlAcxm7m4wuO4O4ltA3WZgqaw5oL05IsfKdh
peD/5Ci8DYVIIJPupqyiL9UaheXcU43JSeokk8QDNlMVgKjUD4HIbAmxbjzoMf1L
+JpV3hMdsO8SpK8iKkYrOg/Bq17N4xTeFP61SIntjRxZDFjsYgSWOLX9o5h67Aar
HcznuXbiNKZCJfvg/y7M/oKjhTh8bp7nKKeme+gU5duawnos3RcDUDIURZpP/Uqz
YJ96pKrn4/C+UCqmVjQyBsw1i2mOYzdlN+GhStIJSdgM6RGtRWreelCJtP3LGti7
caRhylQm/glu0sCvI3TklMyWdnx8uttL4fmrZzmiYZCIENvyhjFdHWi31WrraLs9
oY8tMXVI2bt8qf5VeTO/Ql29lN+TCAGtdWiPvVdIfXu6aIy+JXbX7OYFmCqGDwEw
o5ZiAi9lZ7LGcDTrWMJBSy84obC0/j6avEaVTTqkt/ibftLbdU8SbfRWjGX7fv5G
kxaVkRFrn0A2G6xg7CbYUU6pr9OKDblXXFLdbQG/AVFjqUvzPiA2ZIbb0cMWqXhy
MsTmwIaImJ8qS1nw7T/1WzqB8AbLmR05sF2NqJkWIc3BNXZac0vt3ev8d1gB3rwH
1ghTQIFc10tS3Uv9hjROFu3DJ9rLKVOteel+b9LIH0Cj63fxA986lyb/c/lCLrLC
w99La1xxRfuL00KCgHZ4NApepu3mEPsMFAYAiJcreQeX6Gjr1q6SV+viHc9Cy+eM
qklOjG7yVoVmDklfnkLCEO/6w+V80sTOduHbSeLYA1CnTvzaqGACNKg5JHurNaY2
Re5v9cQbtvm2pcVuNq+DFeD6QMS29qIecJw0RT6kgKoDaOdlPmuMsYi8ueO8/GL0
32kCfFt3OddwJ6LKeTn/NUR4+DGt6dlQ/WrWLGWQl344K6o8sPRofIdWWWGGb2E7
aa0ewYRxfInG7aAjY5Hg1fi4qetsBUvS9rYseA1EmIIVAoy+c0RyfLY1F7QhBYVy
APhphuwlqR0h2BQYz0fZN+L5Zd+7EzHnBdLMIuJAiTV9NPBgPbcn4/g3bziZT/6Y
YPMQ4jVq8v/2oPcLVCwzhJRDT2LuG8StWG3O0P+WEMIrrDLR5/8VA3FS2u4OuMa5
EEhGlTBztRJZ7K+VOI3Of+JFF/J+iIptcHHXuUCvXN7g9ffB4tmkqCJox79foAa2
ivZgL1/EjMomEtz4J0JL0olXyTQzy3ZjQJZVdnJwoRk+D9oSFTBo45mwFLhDwxOw
W7oR1IcZSgTH6PMFaMjDARPIZBZY/cAozLDgM3jUw2r0fGV+LVO/8JS+xMiqAB/R
uW5WHz223l3kgM6EJeMIEDFpUrlvaTxJhxVxJ6PPwezo6LJHABSUXRhv+HceP/cb
G49TVSE+AQYuSfqmpyHMpvtCsrbf6/8E1muge9cPGF14c7aGJd3NB0o4YwGpiiS5
VtPyzuGFB6WC4dVW6UNl4cfw/YgZ2+okj9/KtDfrW4Bi7fwVVCaREpjVzViBQpB/
QkW9ROW749M9MmMTFB9uHn9eyXtUvLcsT5okkZtpNW+1mOYDq61yr8JBoYG6yZx5
P6J/qjrcDwkKl5aGvevIkuL62hnL1JkjFNC9sIvN6lgNNHsTnWTQs66fw0zN5gJk
yb9/M36uuDPL+1FuJ55Dm/5ZIkiW+z1WAUCOPKY/a0Pf/sH45ipG11XSMHwgIxAh
woNU9dyHJ6cOiXSmZFd4x8oWlKheV94dlAdCJgXFpG3ucDMlVjkOYBeo/UT7NO6M
6leiy2eX1VkkpPxTFLJLQBkEDhZ+d1Wg9k81lzSo5GDYDwovrgnbBQ5WlxfCvJlJ
iG+TkaE3BM456K6U46q/QeuZ5/7SKXQlSPsqjnd/H8LVQt0kTxp+/EbzV6YSoWek
N356hBMsFAV/n/tV38k/72zRtTLH/vVWbY+n/9b/KNpsL8T4GXvdcbIAAQncGoYc
e/pq6gLuyfasgWVgqASKvFVcv3o98GqgqTI6g9rPEwVDXrtydqR+mT5NbWjqUjhz
7xEV1JuWdQ1sL86CvLMozoxy/JPTe3iD/me5qR+ZTLB0L/u7rK6aQps16mGofbHR
HrQ+g1ys6otNA3mLaWYzvtzPWmrbb0PiJUbMYFcuzACVwSK+LZd1ueF9TKHACMqB
F41InDqknkKnk7GouQR29vYOJQJjTKq2da2N0KZjHVq82yybJk35c5GOOxt/53Te
g4v1BbjUC1RFKkovNMvKTMNVKpNmO+w5E5mv3PlmEFdmobZzEiNU8i8jD8K+6xkv
AdqNr+r18XLxQTf9xtiUE/z4n44zR9fjlaibh5B4uMi3r7tCtFldYqeXHjkQm+HO
3QsBBbE5A8tYeLCyr7PCAQNNYZNzT0Hh3+PipwGvdPt4amzHSMaTBK6ktSUlyvMD
ZI+26hBWD9gi48Sp6/QTQSH8t5eR1suvYtIqH/tDvZjTmrWYB0gd26xxC7uA3it9
mhDZGUXS54AlTNa548JC3GPOg4kMkhrhQy4dae2oCHTml8lzrN6d1gvBgHCVGO4a
HQkJPpuoeYlDUNQTUQe57paKV/bpu6HCnPNe4bLsz3184bdkBn7ZsvW9L88Kl3F/
r2W5ayy4P70kPw+UcRymAv52yMPtIs/FHGAxSdFspyzHWd2Uc25ypIPgguNhR/Pv
4f0utIdwkOf7P1ZAx/EEcXpxFDriRtuTUDaXF4DnN0H0lmv9Tu/FCqomCZm5Hk7O
SZGmh9dgqVVcqQkvoLLO+tTSpJpA+av0FfCriKLjfI1/N9rkI5bo/lV8ng9P+gAP
WLfTCwqe6cEiGEcdnnrhUDsbbR+kAj2HePby60FDOaK5HvEhY3fVZforZx6A1YDn
Jtc8OSZUhFMm0Uxpqjg753GK65KhstmHcAAadCm/E7CDMwgvyqTLcBTUSbGo8AHv
ECXwH7SduF47ZnO80CbSCl6JDpMiQQSdywEiMW+rZwvtWX+bRV8GmoUYva7mXHzX
+F2FvqJpqI/B3PsBKRBdqo6aZACa4f92aIWfmCSYXVeq7rIkHOO5b0/bGqIYALte
q9R/AKo9ts8brK8IwVyZlAJTxXXQoqRRZ/zhG2iCvR4CIVYwF1pWevdBiuI8LBjp
5x+S4Oxv6ZUWnSjrn6gvoByJR2gnKuq110xl1eJBaSemNZeAMZgpfI0w6YX0K2aX
G68OsF+yLrBxVMeolSPi/OQD7PjGzYYLo7JHA6Uuv+gL6F0nMZEksHpe3trMJF+9
njgu70JHGZ/tpXB/9pF60Hw3C4RAKXRY41+1oLLwzWjKMmY81PUtmpNKQIPwRzYc
PeG6ZuhvGxCFapC/i0lVlPSsvQuNL2gPe8skiLCqcLhxEWbt83k+DFaVmKd7rxvu
63teIpvblWC7T8elfoXUVl4tPEIAx+R2t2Jz4RZAwlerZwtly/Tq/a/+6QlEv2tH
CKYdDua1UxJzEo7s3R9CzXjWNJVpMJ2mv/EWptvdaOWOtGRZioceUp9IJLXNkt87
aO/8Cm/HSzhqW3oSx62+EFGAfQF3ma0hKbv0/ZH327gBk9PLutvRFQ0O0f3eFcPH
ial0dlADTXyYeZOYLhw4Q088sVmAOokghSxmbj70w+wrNIvigYc8t4wr7zNQg80c
ttw1Dj1xRLxnUrQm23O7/EOvOBqW6a4de1Ki9Th5D/4CwzR0tbbqJ1DWMdrD6c+A
y7YStKHTyRvVVQHChhMuKoj45K/3UrJVk9xqJ89F4sdJTRr/D4OaKjTRf+xDA9hL
joIjVkNUHxvDSA2fOS/kxCLCia0rDnzQTe1CR+sAxX00d03h7GIjsBGc9+XS/3Up
Edh5gyIr84yP43BBz+9sK27dCJUaELcdp9Nri0Qig1htyMpHGoufzPjWW46PjgGz
zZmXM3Vj/B7LlzeLd71g1bKGLP8RRErjgBR+gCMZ8vfrPJSGHTEavKYz6+29FOQ6
/nUQtw9cBlEY2Y3+W42jIB15XWT0qFGSIOJ+GnR1NuMa72TQOpp5vyEniSqfgG9+
sZIA5az8hQHlbGcvOceUUq+t1QzfCFJnSTLU5zlokIhRIhB/HZk9khI48raMgeM8
f66y+tY09Hsmt8flE9Jtk247KSDGikkM0eawkis+KvMPwHldg4o6KzzibzpNJUdU
B47CKeP4ILmBuvJsIDL3LcCafqx0jFwriOjeMkEQvy2xR4JEs7wD6jj3OW1pcaNR
5Q5aadl2Au+2nw7FnvaRs5WjspKmxj8U18mkVZv0IbzorhScFhaTtc2N50YGNJOX
5So4OO9mOCudfCGtwKpRywu3tYNK+/g8rH1oxwnoMUNgNwPw79uBQjts7ffrx2GX
x2CFyOXNKaOgOfiEHgZ0GZXeiubKTwtj4J77KnOQYDnkmZDYTQv0ZHx7eSXdZeri
3b1+eN8uIKu7XpE23wVpqAlWPIma+c2K79uwe81YGhaxtFtrzFazP53rkR3Y4fO2
LxBm0uc3go612AGgMEx/iAvUxFi5ymmlxlRkqSpa8IYXWs7ktuLJIVHcNX88O4bH
Xh+yHA/VqI3sXNNvvD/gKvQLC+rlkbGXVs67RC8qC3SdvEd9mKUDO7pO/3ppWB/l
yRAktTolurUwIjymqqWCWtD4LJRn9b8jM1ZuW9NMVbHzYXCJo7FLUDA1VYrrdlM2
t0q1wJG418lEE79xpLPo//QFGEgSPTLSjOswqTzGWRjPAdeLkbDN8Y5/8HIk7JQ2
fv5YxAEPrdP6ZJt0R8o+zpud0S1TTWSXRvaT41ZOROKmcx/LWbKpx/UUN4e2+h5f
jXMzoz8CnztsMrHR/4IQgAXNqL9wAeJZOhXu/KcM9rW6P15NlisVuq8UPO1RmuTy
PyANIV5QeEXolzDxzaF/xE2YMmMeJ8LL7jING+ox0wl2Et37ofh1izfEbUn9AQHG
YjC9OiJTjQZ+xaVST7VKh72cUUpA+O0Yp+OXgUF4BKfak5apIMQaete9HgOmJetB
p7Hpe41KJN97HKBFYEJSOLfRM2YdMZOFGnSFG25M8obXayVAhKtKqjD0IadO8Fzs
s6jMZT+xULx47eB7YVzl+q5VHTulHSn6cHm6PfqJjqpoWJV1Gs4oCmECWtgbPYX+
/oO22kAgwdKrj+ybSbN34jXEoWz8gdM1USQ5BH8kNnvcKGBj44aL0CgeCb4MiAtp
hRlKAMxbl8ukvRdp++0/j+E9b8CS0qgj+3EtP82txV2fZUio+GHja4Mpz2hYspEk
z/wXGCnbLofyUhv2RRHe7w8zFY1C1grA0sCt3SSQFXw/YL4Z0zWRpl0UV2HBrHEf
5aq+3DWoRLb5261co3jrAuD/fUQG74OIGZ4JNAkV6BxOHrv3UCqNczRfOp9hfPHl
lY7kfY4aIPfr0oiofd+BKhY9aky1XIiEXZclcLc5oCaVtIKI2AvfkMgxwzB8JRot
l2keWpxeTHWgoNl0Pqc+NCYWNuppex6EJtwNkHsZYhby4LD2pgBOe9rW2USg6mZr
6Oy8sro++/FMvHLq6cCGRBSmp+jmkUviDwtRr1k9GWHfnTBYCD/04ehVN2kzqiwG
mlnK3VtPwiDvD6beOmcqjF0VAbixspk5eSNXmbI3aKt9LcQU4HrZ1TTXLmSwQUox
MX6OOuFO00xobeqKFG997zZVUtBUoj8KG2FHNsX7YJyENfBhSw+xo3NGhRbN8U4h
1wIG2jxtosb65Gr73+F9r45pj35FlackdHS6QsuNrm8msv0WSElHoFTALGZsgW9B
MusN34uO/fpG6rbKc5l8ll5/5om5r0EHplC0GUD0tIgmO9QsFE/tPQqEWsvbXSFf
YYuLBj/+TVb91C+C9d9Kevb8EPAwEdriwgqgFf4jeTQ/0P2o2dUy+q5YapeRf5wM
JeJJtVYJ1rL7YTqVKCh8xmPerdS349cQaEPofBnhHszMCVFRc0jYeX+uUij/2keC
8kmJzvUcFyQvG/oLOwNu3HnWTf3TmcmxdHiU+hLtS3CxUiw+gzO0IwHQKS/Nzvw9
/GrP4NHP4TO/DV1hyyz+5/PmSPlfzz/PBGbQhR13fdZ2KwfD/Dc/RYifzeyVYw2t
Ejw5Vmxx74BXn+EzgdFXr72RDGLMzHyJo2sg5r1y/3JycWGR5KGmHPrxZ42ycKVD
JszaEB8rh6Gm4LqpSy7LDIPu/sy2pXAc6DUVVdOp405vyc+SBKsvasen2gvBS0ky
tJlWPO/7BNG3ntruuvxj66beN/BTZbi/lbTBaEA/tZ2e9NMpNPcf7oJ/opJw8CeR
AL90Y9B4FtugN2zfGIAg7M5lcLNzYx+cZFHbbqTuDd+6DLfFcrCrPQJX3Y1lF0j0
Kyrxgme/XpXcVl4FUPpi3c4mW8bvAAiMpNJM8mX+LnFB4KKuY/C8Js0fT2JABx9V
asdhZDAmwYprUlNxWHKOATwiGLHZpBPMaAHbTXoZtOEohoOsBHz3K5Wskv4871fU
q5kYtQ94qKjpMBm/geXbNo+TxqFyiS/dG3mmCqIEF2sSOEVGenjWXF5V5zV/lAw0
b4/8vRNLEHa6621K2845/cqymZ2MfOEbjNeHT9cIG3MMdp4cFdTGCV02lnT7oCTQ
NDAK1T2wQtkPcIzcX/0LV559iN9YT4vt/bmy063v2cXBb/U7Z6/lbZGEcbkZAbOv
ZLIBmeM6c81gv+/xutGVnpDVj/G1Dnv19efNJXUbMeFOXWy/QqeU9tfb8jQoOixO
glHFqbWKJA+ybYJtHO9iIlVad1a5hkuymTPyaIu2WqbcuMdZPg6ORxxH2bnJn1Wm
2hm5KCiXdjwSDsgv0AH79hZ6XhS7615aifnQitBcGMljXoggMPK7HIMR3yuucZeD
oxIVYYnpwzn3vAj4AYruxo8VTtPjeuKw90nsf4ssDb699II64GXhr3tdQ0BhGg0/
y95k8pLSRynaP7Hkj9cjrOWie8/d4JU6Gl6Sihv23V43X9B+WhUVrhWHLVnIdQDz
Gtcf/CY7yqIfdjvW2gn43t0bk6KhRnAXXXmKoNFTQlMZJz1c6vBmOUPpSYbN6tXs
Kb2VjptQG9DLVp2IcgDsY/g9ns/ExxNh/dqR0+nuLIs9aIIvX5L+pkgkiQc0ztnG
Xift05xrSGNOigOwpkwd2CvjHJw4FfF8a+0e5HORdSsOvrqShfdSeJUBv0NLR1z5
nevfG0nUu6Mi4/XHLzPAx9uPZa6bYLcxGm13XYfW1QjwP5RKSYIrS+CwNUnS7XrL
HmBlURg5XxE8AqUxCFifpoEjEHKEX8tGfNBXDWmQliNwzp6tvlRKcMesyPOeT3Vp
WO4cxk1HNHzJquh22RlZJxnDV/34k/i05lEjr/zNlKJEsfaBXLLKK7y+TrMCwjV/
JFkEldWYtxvBdvvgWiWW2ptstw8wASggGpkZAAGPWHM1ed1Pv0dsd2ajcj29bb9p
soK5vnHxBO5BOPlz7M97AyeQ0S81qazTixDC7T+C38sue/vKodkdvQJlypJ0zm+T
j94Nrq0MEPHSb8cGurckXRQxXh7PrADreN8EsZTaxOupXNaKyfhOrpUr4Sqc1vAK
Nxn9eJGVb9mlHiUd+VSdWnCOmc1PFRCyYiA2v3qPisc3GHePrzO7HVuAkOb/En7R
mGJYljYZcNXMSWvpCzB6L3+9KyAI2j1/wKmIzTxYHUr90kqwkjLPSkjOntCYnmCi
DNR03EuHBIkkintEI6ZluFegynO7/wntGEbebAit4enMsD+pzsl99ldkXlrU5Jqu
Bwdand9wH3WlYeXhDaKmH8tIx9ViAViEwLYHV5mwwTYnqOmWv3hPztc8IwVGFVy3
TM8fTLZSwsY/M8N0gllHBAzF47Z1fYAsms0MDvpEZs2hANX8FGPT2K1x/+vdKpgZ
AuDuBHFWmpU0RZniWm6SX9mUKKCgk35o/kojTxAJ5GFFj3xixlM2xG5U/hBtnO3L
67V+hZu0FcknZBST1i/TR0QpPFoP9SnERJya4MtZzgQ4vXFYBBsjJFauHXPsuia6
o5KFlanDy4L37EiCzUdqbkgp+MNsP13g8cVTWOz03UJnDUc06tNeHMK22i0hDW0a
+JejYZ+C3BTWlltLVNwonxtxyi/8JA9FiKYUyp7HwwyZmIJuP5RBcBLvqRv9mGHy
1yINwWyN/JZNPoD6yOy7uuTAjRkmvkLP6QsOHjP/yOPDnBVEQQrVdWKVIwJNcseW
MVxpYZJgS8qckMS/2Ekus/uyoaKVZEbIr5Y1ylFwo1XvvUCUD1tOAPrLpGATaMwa
apmFX8oo9Djich2MARd+y3evVdmSIBU6nSm75O1M6c66DFprZus/GBe7XVrdm9le
o83oiIaPtle7yocNMYQe8+FABcnNEGIdibR5sxY/3BfDPAWujRffHOuO/W/mS2BF
JyOwQlFVEyDR/UWXh7NRjFk4q4PHpvvKcWe1HfhEs3I7/0rX6oCYEDrJnTWJwYNa
dxEyH6h5Sq/C4niyrs3aa7sUGHyfVBTdXP16Nfi1obS/Ei+UbBpABJ8p9js3s90B
cpzZb87GkUO4vdORSUA1wcmupqhxrwudSVWZ7jatrBP5gNOzL/iHPuiQb8U4hoVh
60p8Om2uIzL5+4rOjLnr8SsY14O6Mzh1sQ+OvG9eLDn/Zh3Oq5owwCD06NYVyQeZ
jdA6GYNhSTv95bJ3e+23m7PnSWjMELgysuRx5IwmLg/JcL0ykI9ey6YvDf448lfK
JHIj+NqI+pcdl1AYIUMoYNcUaOxUuvKBd6P+VVyRpssoX4OcvGVe33GzFeuPZPay
KlKez9PRXpARLLLub0TtJbXPF8gKZECdaIZ/5jdfkHCitDN2M3xqltLILTC2SIKx
dRDcfmYRKfg0GzrwYCYUjUk6bKrC1EmlzIE+9vCE5tD0ZIV9wkfVIf+gLdYluzdO
RHzmq39NKrn54RY/hLdwyquCoUA8PudKzYqJlUps2b/hCRzS1aDVh1PmRxyKjyeZ
fp0xlexj4sgmZLFvgiGInrSWygiSIIW4Al4P7SoWiFoYN0nushZIkcIlXiqlORf7
fZo3nkChVS+RC26ixek8+kp8GbkEcLlSldmDr5IL8kMAS5oFD2hOcwfLiu/DoFf9
bvQFejTVcQ45fCmtci38j1KmRQFZsswTX/azIqR0oBwoaQbuR993K1riH3HAiXUM
Sx2cBHeStVKOToVCZkXLGlR2zrwXdNflbu2LIlzAAqQgzXlUvWZoUsDFgwzHXDo9
st1AzmPA5nbEq0CHos3+bbOq8aDtBSJj4NvRl1VZ7Bf8U7FnEDxFoSZi6oIa94wQ
WWTObA0kXWPzGio56aILFEgoedErd/Y6Vp4GoTcj95oP7gu9GqewPvj0E2JECW/S
92LdKdXJnK9/TEeL+CWTo17sxy2NA3JbYmT3Uz/5q5vBfbeUiP0clTiDrqZEvCoH
EpqKBpgkz1yMul4uAoIjhEDYd4VbbAKs0TynGz+CHhRTfq/uWNmSDR/w082zUhId
4THlhD1pfstYZZv99+CkLbsUKxH1zWSLwGOMddD8/0TtD+tfCrlNNQxtLFJ29TH+
YSU/nGmo7ysu/Qu2kwOJeCJNXrLSo34JaL1hMOB+5fA6FCeJHWZxLbMLqIfAJRO3
nzpWeVt0wLxxRCU4jOp4nKk7psCwk0rROIbI8BrE96J5OfSQ/IoSKFJz7hU0BRHT
TVA8Vai+QupZP+Z936Xr6S4l0PLBvDH1fWx9JPLxD0/8YVl1cILd9NdSYYbI3L3H
mg/YMq/ZzEc0Lj3EHuHQcIHrfse4BEVUJzyg178wlrN0s5nC3Ai+H9eJkYdI2VyT
tfF4eZUDn4gH8TnPfInqMjTFM8bj83dHzT5MkPGvcBJ9aBCmWkfKEX8HVdGZpS3X
qQUaQDB3v3dFYD+CeE/yBTBNuHs9T/NGVkwUEdssNcsR6IdbIburcYlu4EZKsRBz
DTxAognSB/Z2NhLZWRuiL3hE7Deop6SUihqLeGAZ/PMTvJSue8btlsuRxnJlgRWK
1MkUTWGJmbsiw5sDwWbtrtwhN1UhRDDk7DRMyypQmD2ezHiM1VzKGPakERuVD4TQ
bni6n6AdvhD8vv9Rx/XuBBgKPxTpRNWNsrxDEgmq8ke77eYu1FF6oHTjKH46ohn5
GCpQPGIYRPZxY9s/lD8zUTbbJPqE5WLxlm/hWoxFcZzwReCzP1irITiUGsSW/pB1
HTYJM655IXEerVtFtNv5DkfLRJxz/zbUG/Aox4Gr0iT2O017apuTHHQm93fdXSpP
ksHnzAQtKAMYR2J7y3llEmccCrxQ1h6Gr0eMOKA57+C1Vaa+AwFI1vKq5+h0M10v
fDWSGdmQpOMCaVbJMVfCE62uFHllsrOBZfLZQ3zwQMC1UY/VNg6LT3dGorFLgT9E
Jt/CjoIOUdJZJyw2V6wPkSPnf4Wh+b63ajnNFwENgSbypFgb85HR6B3hJopZit4a
yUL4cwUXpvbA708hgFMavSE4xPSTpFAaPPY1M+GOu5dZpJ5ydyf5tYv/eWgJlaFx
gYVVbxASoSuNQt9qo+IWUAixuVKMsDDS+LyH/GcPkVYviIDZnwGCUTRs87Oc81Kf
Vc96Gnu8Qgr+W8iQGtkcAvv57wJ3O9bxCcG3uLm0qQlyaMvfq5JWMhhOqvjcVSLB
1+TQ5OQ/22uX6SqR0W06HNcD5XWxlw9MFSRBwoirpi1sLjc+WfFjKZbw8J/6rxHf
yTanJAmm2tYxax4h0WiI63w3pgpWHmFYAC+ZkePAuJWV39A9+KScKeYYiezaWDg4
gDV1Q3jnKitejd2PawLR3KuIYOmWkHAjQ/XunrBLldHPkLKAvzZEO+0lmkWrPOfJ
J/3T14hA/gvLyC1cMeZCEHBHmSYnVu/q9J6XSLIRIcUQ2PTwI4jHlCxJUnhCZFsP
bvijZh0OUEVoi598R637Hle4jkPuyDOyXebApHfPs3iT9HDT1tQrHQbgqMx9ojSS
r9+Eu5X9AxbJRGDrsli/3sUCVujLCc1XiqvdSwivccOsL1hZwjKmLcM19/CenYMX
3ITIqBjYUD1mG0M2JgixR1cw7ZHMMQpYr682mUgMAol2Kyypb6iU2IL110rt0xY3
6dQ2f6wMgPVTSNUEzB3/d7WGRV2lBdfe3UB0500vIKvlYmqZrKyOIIe6NNePkOHJ
PeVAAdIkG/ndAGO7DbplMGhA2Dd1sS9VrgLPKfO9FvKnTPjvRJau+rHqMgoYRVQV
33OaFXd3SCLKTHXtUX+FnJ5RjzrGxU61xmzDOsUlM0hciyLMWpjxmGcQja6Kb2BR
Y8P0c7naqnTgokOI+v0Ogu04FZQV+cfgg5jBggvyMZvq3vd3HoeBcHWNReYEZ8bP
/liOF9IgIKg1OQejn+QVdCVj/O7/1qZwVn9M8/hrttlcTzUAidu+HEE9MfWpcxkS
3BXSpbW10GE327BWAdNpMz6mBJfF99wnYgD8procEiz5qLZzXpKrx9yuMYiECbyg
nuSsCh6ZiyAXFB/gbAevjZrq4EJEqlkvrtKa5ewTR7/Aq66MjdfQHcpMjwdkiwsP
D4AbQUYgMXTYBNxUOmK7Or9PSaLDtU1mP15dxfkYLldtnsr7kdQtK1FPFiV66+bL
iVDjD1BIhHiGGP12qmIoQpzPIdKAJdw8qXQNI0Awt1PdVoIY4XkH4S4QNWLBa+0/
TJl1/2fRnHZHQWjG605NBMHUs90oXTyrMg+AvUbTae23+awsJrngwaaPPNhjdDYN
2x3LtRz1p6xmHDaAYXyZn4zmT7+gRExUNz2Ky3SoqNZxfWKOMN51AZOo/Z/gIWmb
i1hG+sGCvZuNMZdURLQGtZ7MuOTylrExFyj9evHy6N3Bq4vr3t3SvisTR3ivqQAH
Oexyr8+hRmbPz+peukVOB0MEfFsFOLLOjf7ZiqGpAuNU8UVzrgDoGrHml8/QqG04
tG/CRDGzc4zXiKD0MjMZJlHW21AP6MYRtdoeyJrwmXVHyRHHQ2Suwwkhp7MGPJUN
78Yj1z9gQT3sZ1Kfla4woti2666jCbE3E9LBSeVhmGQnfooBBLuCDAUv2oUWYLJo
30CZXuWnMWgOostDsNWZf2gqQSbfFZRoCIb2xp6Qx5i9kyW3MHaPI0bREGw/TuF9
cupFtaEs7gA41cpaSTmjr02YpuN8rsE45uVUhf3K/aTPFDu/pKjGERkb+QdV3RI7
G6ijCgjngfoD1Re6oSzRUXlmbBtf0fr2Hljmg4t62uDdJ6ap5A7W7Wn+lt+uChIp
KrjeE+gkX/oRh84Zxm5cff0b0jQrq1CRT9CAHg7qd4m/eT3qI5x6jddkGXQhm4J+
mc0CoSLZZakungozftTwfk3p4/VAvMVC3D19V9TLRKc3SjzBQceYP3hYXtdQYzHT
MQYaS3IMpfs06V5PsIRdyT6of8+99NuuAJ+EACzeaefJ7JW3QEdzvk8zLKvEctX+
B7HS9XhhEf/Si25C6JTSj95sdo1P/O/VMrMuYtRmAJxGsjRd+xwH08ON6CEOfWe0
nv7dgxJuM4LkY2vZHKJ9eWwO7Dkvbkes4Mif1rNAc4ECWGT/B73fkWumKCZOJjgq
vxyVnGb9l9fbTenwjClzPRd+WR0g71oBUET9YI2Da5IlrC61IQL61YOPsp2XUHiH
VDkbsUJQ4iDtd+BOZR5IuC9Y5Ba0Ja7fmkaGjI4MJms0d9jVXa09gYUwMqkw9QvT
Ovw3y6eo+AArwfjXJ/OpGyc7J0AgUsU15FCRMn919sNYAINkRWiCCSObxQM8cZcj
/K8ua5bBdUM7WwD1a3E5uD5k/05oKSaXVufEO+1wn676YMetFR75wvEV9xV1qiR8
zp6j0aj2YgDD/EEBnYv9CKT+k8XRx0kdyh+UGj0qOOE6RQuvmSqwW9lACCs4s97K
qHaaN5FsPgWse/FXBGEXrQS+2wYLnu7xzLGQqhGMzTyFFl2lnFlarvFTIvfUxv89
UvEMTlsGvdqXQpBEkb2MfwA1qfIQqIPhtK3PxYnHRhcqzWb8kRPDm1RcydJArZZH
ibVYYW5JWJUt3ilMuZeLRlHVIKzfR0z4+L1OotHNoDYo2nm3ExXaJIXMuGXur9Um
ChSn/n/sB3SlAUt54VFHKnXfzGrxRwMpoaYr3ighBW0C7NszGE+0Ag47HR/q4utb
fJ4nGzkkbWIAQMx3oHAVio6AjazUofRHKo3hukPFfJf69csRr7A9hdDYbLoMfQq6
GRFqHjzDmJJ2y9glKvOvf5INewUVxh6pfRpK+cEcn+VylyWO5PFWI1F8KoUDr6wK
nOZF2YzGjikJoOmgs5pHUxbB/+g+oGdUhwSzcwTic4bSTC/QkLb3TKUx+/ZOnM89
z3tetOSDav3gkU7dlpdMfy3yvUQ9GlITWt0J/WCRLprtaRRi+27fL4pe3KTWSqvA
dSg4dS3sfWMIXIFhtnLn4gSIIhHq6p86nY7gmlkSf0yRKTDZ5p+dkYZ9t0or+X9F
mJ/QI39muuppuHTk/co5TvsNWhVeqgyqUYywomeYWBEpE0NGv0i+qsaXHuy7Sj6t
kH9ixwqUkZBlyWrWjDS2shdH/6ZKXJbQ5G1RWr4yRO4J6LiwLLajeunygFdNvEuh
ZVcBZW2/wGRkgBIjZ0DYdZ5sdp+wjnlQen7C3z/rZMKp7s7SyQvTAyltgDQ5EHX3
ugw+Rah142kfSJGyHkRochzjsp2B++Fqj/8JfH5/3aHzvv1vjezvrsvtySEPdVy7
i/mT43c9751GOAVZCo4n8H1O0i24d41Vfs2LUzZVFd2R7T+3xEO3BPIRDSIF1PDy
P12qUxFQO4W81+E0sUsRc9Z71hiBH7hgqSsmmqPfUdVZADJapyn7oThjN0BT4PnT
oc9EsZ6TBxZz8W6zkmc5NGiFRJI69fpOtXCFtFplICEX5FRNrjOd9h7q4O1b7d5U
Gd9RkpCpSg5u8eI6n5h2jiksgIky4bzKzPLkQrHQCcQeH6rIEkIM6DOcYvMRUsh1
5qzXjB/u7JkG/iiRetjuxcxPYQ1t7xM8/0OcDDo/+bVkYpALeVWqRiv+6v2fbUhK
fQqzefIM31qQrexO0glypAKZSTzMTZxBpN1duga5TZi+2YnAW8BPe4FOp3HYJLxy
kR6bYhRHBzm46RGtm0LxG5hYk66R2ZwWKV8d17WRvj7NIz7K0hGKjFt0g5iZmHwy
JynzbmWRiAEuypVK/T0AD3d4cbp5CF/x4p1JXMCCTRmpm5flF8E2DTkkKXEXKwJB
S/cj1+WFDTSAjW6xvvRLuL1bzhgfOz89QTSh6JOPpzIPt4J9S8VNFVbte5TIKMeQ
znbcbqGtRXhoV3wnwjX2HlR6wT/GD7sEoDiejeRlBRczFuAf8cgpk0EDNuhS3H6R
WacU4x1nl4Zhamv3zv8MeragvP1vz6aibladXZ9rhAoxE9zEKC3tT31q/12OYIl9
th1WwTU6warofWtxljbX8+QDT4jQebdeX4Gb/+sMBkgw5awUTRbyiqALqfhBR0Gy
DuFV+Q/X/RV+iSa0F2p0mfYxvd3tVmhbrYWIJVsdGPWj+HQ7CH/MJP9zQWs7pD/b
U0GvvP/p2+GpXb30WVEGwlUGpLn1ppGOClZQ0C6kJLiucUtq9Ave8oyRcK90ixLx
RcXiVRt60hV2eDSxITpMOf+ZuyzTRCVOPlq80qvZKKZUOycs3Gwc3FZBY74zqKVt
ZuZccFhD5Pm2uDE0jqMYlnND/l/87aZdSG8Jxww2EbAbnFlDJZ9mLhdtc7EeaNAb
cQaops1rdZI4Edp6n1ydrvZrWkzNtGIW7ETFt4/1azcJ2vrgkqdJbsCtM9GrJZmj
ZvZ3opQHyGipRz2saDnyTlW7btdlJU4tQVUo6KX9wnEeffgFoGHmq7PIehC3AWjK
rbIWCRA6nmt1uxiPEEpc38DrOQ+Z3Qkqy0uCZOgrl3gdHr6E0RMyBdW6P4evNU/t
MVA88iEIT2bSdYu5f+aUWllmRjLhWtXqNAEuioF4p84/fDnRh4VnzEAC8RZlnfEZ
/crq5018R5OuqO9iXKeEQIZOZtTXEKF4g/T+6tzDWjrvNzGJakKMd3MoqaxYpGC6
/4TuWZ8HZVKgFoSiHTjIaIio5SFf2D46/nbve/8m6Dn97sp6WvFFvMBYhl2noDwV
me5vlRq8XwB10Md3C4mTByEYEgI7RWYQDAQSa+qQmar7/mdmYxiiJasW8G4usqPt
YDBDD9d5+0vsJMcuYiR5X1PJrsS00InaNFNckRaujpnWat/zKd/b0qKoqaXBqXGa
WAs+5ZddJQAad/tJR3cC2j1RkPlcuD8a9r23kdexB/xTGWvcSJn9AlovX+ALinuN
VJCD9vQdZTLEjJwH/i+cUfVHrEhwzbL2TWIZzW99xbzy5Zj2bQJL9soBahDPAhak
eXyix7BER+9pLs5SdVEosPvND+C59wIEmuVaEBRGP3SjgJrPAjIvX91oZIxk/Ysc
5p8H31LHyo49bRJ9pNivdKJ6FLHrvRxLYJq5ecuBYixF1PZD7bOhv2BOniajWKWl
6I9eKVRu7kybsBXdpYLMt13zvXYwY9+BhgwPAueRzUKdKH2rTtdP+6gh7wLtzDvO
K+7K4AddmLNdfszwwDPLP96MPrpijO85QLVY/86fhRhsk+tu++ZcZldVbNz0Ix0H
dKKJp9YWW8uNYIXVNSWNRGZ5WGPUPjqN1rsXaul6FGvM04GMtM4BVsUx3IW3Tx+k
4OCyHzuLq89wcrAzUIDYQchkNZL55b2cMbtYHhktHOqQdWnrJa00OpNWdxgdg1cn
F/o2M/kA8xc6w5V8amPr4nMdBaej9OKmfnH83GF4RFOzXwdlDZf7oaq+zYukb4TP
2tMhx8gWy4sXkJi6CEBCjkflAitfT1srdyZJCYBHpXMEDWXjkN6NvDEn2d8zW65g
wPKK+xyPXbGyTDhSMYWylJCiR1Lhjm2Jo8/2VjsWYgxy3/Enba2SRp6mrhXbijv1
xLa6hZ0h5LLJOPCEyOlkoSYng1OXK1+LGc8VuliKqQd+MrZERSS8y0rfKJ61FTVG
1+HaE0QCLIlnirknf7rdYax5m8qZTmjzWfSaYRC2MXNAUSNWyCylKkA21P2sKMz8
t+4fHjLw9+KN9HK13x0BkoaSCAOc6fyiK582lfeoRLJ1dqU3dz/aRk3RY1PM1pg8
TECccQIWOtox57PONCAbHcrsB4c9hL974K3wLhEa8A8CvAx8BbdxkhrqxJfDLhLL
sAbcdR+//d35P6Bz2PQE/jFQZtVM2t8Aj0ofcstPjHq93VZhAf4oaAHWEjLH9ddN
SHmb94kT2Rhb541IvCCJ7KM9msi8lWFEU1KOGBNRK9Q0FJbzt80R435Rw/GiGOWo
8EaKflWJyuT0T+YD7Mom8FLVFwYC+YoqXu3ReGC3KtTt2B1oaeW3Uf7wAFDIpZjp
SbKxDG3N+trP/hGugpiiVsG1mDvE1C2rvF77LW3a/DOgOeiY2x+Ho6h3Q0Pis8Yx
+ldkHCVbdXJivR3sxr8XeAlt+IaKmMDe00mnOeekE+lCk39vtGphIPdpc7nNLoNe
hGt87TKfBGCMkxgDwvPzX4G4/NvFGDwRKsguIyVQQEPWqWtF5NE6VXpnWN456r5L
JwppF659BoiJt8397vC0xo7SsfeGYB4YQ+INCJrqR5ft8k9VVRL0emMXGUhOg5zL
bv3c8A5OVYVNrhzMjf5EA3ktZ5JFMAsEuS4XttpBI63FnGioxoJvAoD2cALdXH7l
qDFa4m6tqlUKmer7tUyMkDEUmdT3h8g/mDvvOHLBBQ+A+FV32adkKNMZQT8S5yQm
/QJIjnG28tiiQvQQ3an6G9AnexAehQQf7i/Xu0A55qDUS7Jf6zdL251/OX1CWRgV
ZFWtr+25YtYxRT7fny2ksSC8KuClvqRpuby+Wz2ZqFXqg3JKAsvBh2DM7UAclX+T
bfJ6IRqkSEefMMPRAqFIqst3zW5lrcqY5Sw011DCvdkkbhkw66LlA5kKxTYCLdvo
fIp+ZWHr8bCV8EVarIUxZUBAjIASsmr3j5ouGZ+YcriaqBTN7EutwCrHsI5zO/ki
AVRN4hOwGsmjQsJCtr61M5QK4FegG6YMh3fWzDoPF40Hja0438gZfn7yjweMRLfV
a3Mn9yQdHH54s40BkRkbq6QSWBS+8in6dthKhklNbQEOh1h2/fSVo9EazWftdm3F
ByNWkJPq/X0+yxtmyebvTWSQNvbSab8HI7IbAlsydpMGrP1wuBRZTKbPpBGvU6lw
aJtDi1AN0xUV+WSXY1rnL5lfyWEWn5CnxOhj3Am+3fQpRs9L54oYnimiPSaxjITn
uUglislHA+w1X4Og3+owohrtoMtLAGYmLw8N/UwZ0fsZEeEVcK+Sl7CB7OMLAPFI
01LFxVSK/bL75A/H60ij3jM4tD+7O3qfpxf5JBDKKvCJQ8c+ZVLqObH/TOQvkdLr
Ubbb07ZDUsk8kkalZHoR3bz0yMGDg9YjcfxqgJl2PvqhFflCjvLYfxqtMJzWlH3D
pamu0+8mlZfLapc4pYixRTk2cPViYvvw1Sncaj9Kku3eyG59Rc99VVkczsyh+1hw
+m29i41gkD91vXGwTtrvSs3eQ2R5XkgWttf82hmuaxJFEbz2LvGPnerv8qxOusag
BeO82/Qur6iX07zS9kBXm0zATSrSZOMDOX9x+aZG7ymS8D0nrg4zfvYvpRq5m99l
RXimWSyaY4v+gIC5fQKxivS9TakYZ9/ZAEfb5Jg5uPOdAdk/SmmYuhgq5DxseGyo
YNG3Jbv/QQ8M+EvPkHP3oL0qLIvBYUCDX6/O69/bBDrvwbycG+VQi9Lc0zV1UeiZ
Snlbzi+1W35kr15MSFuU675xHu+Kq4mxiQ4khmN53l+GswH1lcMKGJy0BCrR+2yx
kZx7M2jcdl5rEFOgks7+ya0ks2D0LHr2z3iWdCrMgXaFlaUP4RzuJxG6Vs5DGGXj
E0xUJYQ1byCf+YAE/RfJrq6iMM3JD2QaaDOdAqc5KRZdJoRbVtRULTQHUT+7gJZg
5ZHcjV8dG9Ifo+6vfHiip3ddNxKYmJ+jMWRr7F+zGwosLDyE/ElvxtG+CuCnPAFs
RqhWyTlQF9iwqmLQ08a+0hCt1jM15xyUvFYfa20vxt4VcRLC/zU9F5ANBkAGx+Kd
XLoQzCpaiz27GEZkx5KvFRBSMpvyfkj0zc+06AHJ9e8/IBLT/rR985z7f4/15W6l
szwSVqpq30LJk+VuZj5MaG4W3IG28u4GNBJcd7JG/1NdgHao3Qz/4/JR0BHko+8E
gZa/xh6aOG0h1qIyEs14B0+obLaYiel/Agz3xwZ8+jnNjm1pib7zg/ez9DqiKNdV
cHQIgEpD12EzTTwksVzvYlWcyz0h1fIeqeN0R1Aqu9pgGP27rWEjL6hksxv9Akv+
O1fX4P+XLLl9DeP0lIkkNYcJh7TFoA8szESiTEBC3Jl2hwu5zwXepgkNr/XU6dHO
WBp7PwtiumwYQ9egfosIehEWug75RB4pLAQ9uA3krhbYJyKSJ8MWk0Mil9djkQNP
g7vX4F8fEm5av29tSHKDlaIJ5fOamIqW4Vw6N+NuyWlDetbV/vV+qfp98IPfGxH8
JXGxFQX3DEYFSUDZovATnTREcxHJgZMGyQTEFnbEsX50sLHOipVlo4P4y8z8lWuG
1EWauEjufEl/r1CqgX5lwz9cyN25cDPDyWBWrWfaniBRkBXUIBAmfaaDVxVEjPM/
MasKlmNaCS1IB5Yw/TeK5ii4+UY+we7p7ua5A8ilH0ruJCFSr3u0TCEy0vQ4RFFc
qqFgh3L3rfMTVMggGdfbNLLRwqXutSemD3AFpNpIa6MiQZWriBFvdb4hflxaEWG4
vCQf08ary+A5/93WnNpKAo9nPcpxCw0qMmev/PDKzTDpXB+otMQTk65Y85tdNn6f
WkVR6B+fIRxKCFkCbCo3Bf9DCk/QGOIAt3N/KRPxaUPPKNFvfAKI8sBvzLhQXEF5
YsjzHwHlDlh2nA9e9ytr7rg0vIoGpe7IvY/1tNapZYH18gf6O7Ho88nEcdZQdzHW
UmIkR80Ax6Eo6gmcJeGckxt/62f2j6JsoBPScPkLYYYtv2O8AiqnnFX7WLTeotox
DA43Z6K8R6eQxdV86f2C+qQGBKE4JNFEWmVR7Ouse5wBftIIFyl+tswH+lMeiCX6
npbUv5VU5LVXP95/lOrc6aPUMpSIyROhKO1TdCaY+0YfIHIdQC1WkJi2fKlKu/Fe
cLT6AiOUKNs88eo5fm5ncbiF/nPf3Itt0CG6cVJ0VB7EL96x2TsL4Npi9/ILmwN0
7PXzrxe8+gjTJFRxC4AzF7uqIY5qHObIs9rFDtGLGuGfjPHtKevWNjBAchCYfLOJ
60ikUDnbwPe8RxPlMfwFSgxufwLPDPVdWd7zGqCocA3qfnNrAn96aOPdulQCAyiH
XL8gyG79WJNu6BNpkktyEUFrl/MF5LSYqmLyWRH0RofjqeLZhN9jKXnuIoTEFU49
2jI5VbMWQvO5geGWpAuSj/czbrCPNuUELsVHY1c52ZESKh/kYlFN3WLlSOpAEL9B
c03Y02GMUO50TWv8Idgwa1q/TFBimOcf/5tb1OpuHRZsoglObJZZZvRDz2svC8AE
rOxfNZ1OQsBqiPxmdvrU4ns1BYlW75j2Dy6FxpE5DmL8NDlBw5/2wZYl31WDYxTW
lhK7ucPEJlsVcMwDXeHX0inuUXLpZ/1m9GbeSUnTioGpdLvyV/nLpT+VBM7Ji9ro
SEcbt/SJB1oNGRZnpIIV1DNT+/FqMF2KbDbDvX/4k2na/rj2o6kT4CzkjkrjpIp2
BeyFwC7wnHV9Gp30WpzLF4WudyLhJyGvGXrsO5TUePLi/bR+fuac48f5DJmk+9Xf
7qAIBVqvaIthRtcy0qLLy2uE/eE1MH2c6BStMZYb2YdN0GGASCv4iJNQvBdX/l75
+/d4akN3VRBuZDK7uhXBo1pzIrf1lYM3hpWNzDwZP4GAts0nB1NQUmvVGZB17WTw
goSyyG19mGNkcckHpzze+ZXeP/NRjibUyCHptPkAMRLk9wG32ClEjREHQL5Ap4EO
mNQLLqazQHjc74C6N95jfed9OfeFMfDTUDT3Ub/EgY0Dy3PXbQbG9Jfv+Ch+eyzI
/vp/KXldVS5IadPY9OtGtTsFQoU2Yf7USW+eitksWGKH4604FutQJV+QqEoGhpmx
L1nUYM15eWlUKGRzezRpYUMIj+jXSDsY82alkvi/m3ZoUHDZqeu1QrTONXmAd2Wb
FWYiPhG/NZLVZIhXc5osRnwEPIyqzWm5EXqWYCpdsyl/22PAyg+p/Wl6aeP6a3OP
q3A7HVBD9tl//yMwxTdkkfhbvJwla+pU9JRS57VLuBn6eevY/BZ5NZthTYlgrNQW
5JdV63t0vCaic/E5AsZmZqKMbsLVGGGvMfn7Betq5Lu+JHfAxy3MVbMbg1kOo993
0v+gU47JiJQ4uBCnV1oZ29zJF7CK8vUL16DrQGnusb7e+IKJqP08hno2HIwOjheN
47rtW6qUaAVUIKZNSGL/eawOf5NE/tcO0CxCRI6BV8x4A72Bgc7BOd6cWcYaAz9C
5meDyi6UL3s1kL8r8+DwYFXfAOnliUndcPYoUdRNHHriugLsWvjnOcaQgP6KoV6H
tClbD0P6Pj7uFQ0sLHVllyiIdY1k3xu2BsU867OCbtIkyknrtfkf047E+F2WlKwW
cy1bp2Lkje888pCfKk8131i2BXiVs9kK4VOqPof7u/IPsn0Q+Iw176IbY1+k/D+3
xJJSMeOhnfPNO1UpZ3KXFvzgXoCsn+qGk4zfWnzDoMGXCeDlijkeYDkVQZcEUNCh
E8d3eBQy+RlA7NvGB5g64nvRusS6MwARboBm1H/G2UcLcJYjl4jSSAEIZK1cXi14
ga6xUv9ngQkrxjeJ5P/lYyAdsNcPo9/Bqs9dYX+7dT9bxdfix15Wtlo3C9u67QMj
DnF/+sY86UZAp85zsdgGOr6JXkQCp1GafNlN0k9+4lSCy7dZMGqOONFJriXB4T0k
7JHrfH8xaUiKmS2Y1cOdmH/tYdTyyn7R38m4Ebqpb49YlDcvYhXsCV1tLrYWC1Hk
+ZyCrMfXoLPNbpzUfw6+3611Vm+O68dhjw3CddH34rcKOnkeMuh5GPMk2pgdbKMi
8NMkeJE9VPtlxRpdqZHeQq5xftJMtkxTHUsME/57RHy82xd2SvKXRuZnJpWuDehw
ITkwiR67i3ykF7+nENdVYW5hFHW+F83Gs0px2JL1T5LAls2orlBikB1it61WDMPP
PK+2kWxzjdgSgjdNJ818aTIn38Oy4l53DMadBfqzNz+5OLrJLx3K5qfvaGAir4Qj
47b5JLOP6M7Mmy1UxAF523jBbNuuRNhjQTfthVbIgCECEM4QkejRkn1f+vLVcA+C
e8aTDDSgbKmWp4AoK9x/fCVPGT/ACNG08+yuKbXg2HmK0vUJjlwbF2ZwxAa27CWU
MaBdSlHe/P6a9YaoTd5w/UvgLwLOR3qllptVDK+ZUQola+k3abROPfj7oSKdydSQ
MDsq/krJsn5IhRernU6yvXlDXdQWdirqLhjYC2u74Cb34ZGtOGEXb59jCzyrqteX
UwgB8C1hczuGeGTqy5Xzf/TbqzWBPCxurj39svMyInu2QIlxpRRkJpQPzZoX52+q
j+XdQrkN7r2xj5jF3d3JxRQhW++4pKb+b8s0a9ZYthQpIDNTRxgboE1tgE11kVZy
v71ZpsLs/Wzta3P85nV2BYuhHofRSUVyoRpCeXAc99EU2HSXFQUM9K+pV4IbYxeO
Z8AkrCG342070DxHYa1gz/1d39JWjPtTz0CL9VwLjpozJmbvxMG6H+4EuR24F1Ew
ORR/fEOvKTmZcazzjvuDTQHTU3Jq/gvivZir25jDG0AkUtwSm8SMp6Z9we7FqwNh
urwvF/Ipq/RJ+5bBzZubGy/W3isc0PT2KDlX3PmJEFjHnc37wq1isZx9yp9yRkzf
wH8eT3ZAGoZBMGgs8X2RSEdCSRfv8R8Th55XX/Mo+HQQbd+5JyVT0XzBSvs3/TtA
TmGPqIR76yNOWWzJ1290orZ8WJyf55+CVRa2u3gxeHD8IlhFUpfNf86aWhn1r2xo
MDz42pcFGtyS2ecBZG9HG0sSBNOA9c9DqOqOYBo2+oTGWmm4NVp+eF5E7xnZU7qg
R9sELQmgb9FwwXbbuFGqrQpM6/eLHBmfmawz/Bk46J03Go4fB5tuFDSn7/HS7PlK
yMChGrRKL3e07BMuQOl3VaxTfaIUCzJa7jGY2gKc6Horx6hm76OJoNuSk2vV/Blp
Rfos++E1kYWVxRgB8CfrJdYgpvR2+5wx3V/F5PzNl8WZqyyWeTKgCBFIf3oaYZDa
c58fwSYiINM562yOt1Iq/dn72UiNkjm8TcpDaVmkZVjxsTqibmrPL0B6ZLQmFIw0
jTnmp8iBSrz2i34aiYaWduTQYsXhvJJpcsCk1pcIppb6dKRbnvELnfDgsM/5M9eZ
OCUpmAtF4pi41++gZ2SenBQzkWU63rTLdef0d0HwxbeQGsxXbAmjuALZ4K8tQpDu
JCXfKcEEd0ZRjVLq2X2zcQm+lk0dddHpCy2D5BlN8MH9Ab6zbUdytllWSFi5jv5D
osKgYMoLY7uB8YUuNFdxulTNnDEqdaFNlMpf4bvR4rrxAimuN1pODt2W/hc932dN
uiN57FsrNDRg9tOEbxyBDD58CkJQLWThA2ntjMO6nTQ+4swEkSOGIaaclWaVyMMq
cz0xwT6AQ/bhBu/O2rvDR0mdEtP+JF8NJvG7bcTxXrk40KqBuVpDvtZxJ7xD00iv
EYJ9c5TL5Seei/rIRkr1oG4ByRMx/cFj6fh2g4PyRX7IZi6EeuxK3O/2nq2tAqIp
VeF3vrXIsXt2FXvd2SvcfbBBrCmtPrsYzsgKaIuZ/1V7h3HS9jYQSsRLgni5W3JO
FAYEQHmIqEKAUsSF/H+sWMnFjHv3XzSVOnrmat78vlOfWUZj6amiwkghhSCRyikl
xFnFWbwUE/DFJDrwur09VjlT7bP+w6rnbTxnZ5ALiy99ViL605opFIJLDsCsuA+g
Io7IM4afCoM6sv4UUgtaL+jS+6iI7Hh7z0x2fOXlsjzsldu9mm/EMt+3D2YiYxqe
etbr4WqBQRTkZyOJCtuEmd193lNJC/jUL3kpV9q4aCtD1t9aZNv32KCWXr2BLGyP
2Oq8IJPS6HTAvE4TwdLweRQyWS7Q6FmfunsRoXnY3aRxnVnPLHedkvGQtoYhyPY4
gquTt/6Md1tG8UwLLBVKBAkCG69njrf1wGCwO1gRoUweRp9rz3HAURSh0I9IqOAy
tHhRBUYYJ2JLOaZ7Ps/a6pKTIUV0Ics7WLGWvT6/GmnWdMIdAIfXaWQjjyMTftgN
gpOHlCHLKRg0DIzeTghfL+a8a9i3ctnUWMOyC+Hrjv9aO2yDCbn6FdLQLMGhT9sv
MaUWA78FTmc6ht2dmPgybfbxUUlZc1JIBAz5SG/EmBXSexEPkJ5DCrZo6gwlGqxM
gpV4CQ0Eb/KxIVfxHljrE/iv4WxIkc8MR4uuCOJ5BcT3Z3vamm7bu42jH1b7vFjR
0J0wP6e90cMUn7dWSkPMSj+8Olm8lMoADM4Dxg1NQ4ed20WbKWilNIKsu0NV3XjD
+LhORGwERdFWATnDzIRkRmymmlWFlw89S+78hS8M0KFuWuL7hd6rxe4OkzFYsWmh
67CG9kT1S08SUzSDhBcqxDbCmUbJDi2/K6tbCRn2OV2b3zGNThCw/My/QmykbG3x
F/LfCjuP9HS6FvnwwFYA/o7MRRPEGrq9+HEWqLCnKw5Jbhdkg0mnGUum9FB+4un1
BHMp3OICT+CXZkIery0Dxjq665M3qYCdzvw7TEMk7t4TEtM73GGzfkqz/2rrJzaT
vfH5Rp2b6ZqPIKVgg63WwpvKFb/itNB3ucY5gu7rLQcOdxif4bONd+e2I1NLB6PI
sCwcGsdq9aq+3CCDvmDM4WgUVMvrHowFrOdgAmbkp/e3iPQGAddeIkyeoZ74pWIJ
NUKqo5noUHgBTYefmsDtSCRrWiL9p6CeGgZ39v0khFNw/fzNzzXKdW9+n9P8al12
MpkD6NGY7W1u1oLL4ephW1HarFb2wpn+PfzjfiUCUSR5w6sWxDquGE4Ww4g7NGDd
av2QjW01uu940QRIab4Afck4u1vSoKATXlUlpKaAoWL1VZHm2vy+vdn7yOGfryuZ
xxsizVmMYIxl++HW3Hq/Jbn9BiP3mG3kIzlp+KHl7WFIv0NROqiVtFkXY8yX1St2
gtqqpLc2t1KRdB52jO0zEzKP572y69g5CPF4pEgsbRVhSdXj86ydE2PueXGXsVK2
uUpNoNzVw0IRUSHmShd5jHlEUWQQ965uVGjsBaQaun4CODr0YrcXuydNkcSUheWa
2W1SaVbwYPL2zBEoC29mvKRsiGeWj0Fq5e9fA6Y1fik8Z2XIV40f7zbl56oQzWiw
yVY9jyHb7oVOSQBfdmeNea59Q63rGoOIz+kVVpADe9QOitsjUmIKlzfg3luMrS1s
GQ0HLxDEzDvTF0dLB4fN5ZSaAlxwRn6VeBq8R7UsRG6dKRCzUqubBq5gR8RyVIXD
6PhBWXKi2VknRTMTS0imhE63Hz7YQKkjA9OtyS4E9rs66HpYhS8Z25ga+91hGavA
UItUZHMPM/BNqxTvdxSl5pFgNgY0q0Q3R8pyzsUP2fOStyZ9103Cc/PJ20OOHe7g
cqtSFXP8gtQAGarCQQfFoF8lcvgUcMgNmbf2fMLUmIWHQgMf/UUUknZdsDmIzFuy
6bMJdY/l3TmH8nE1vtGq8R4D4qdPg+bf6MIJHqzPZ47GTuvfIbYCB6TM0TN+a4fV
udUvmQuMAvpBpgi6y4WBNmviHwjk4jZjSArlIAp//ATH6fVoKyEYTwIuChRF5qcg
dbc0fRKtHR+xi3DXSuahDuiExGlw7bgd0i0P0neY7VE65S6mBAnfBG9ao2bWatM+
/uP2NVxn1YBohcDHmiVO5fWPWTx9XpqZlG1s8G2QJaMxqOAxLYisz8Q1fVaLDJfD
Xi00GUmwyLTEi/1EEXzEg2em+cVkBJI7QLmJbUAfpcG2/hJmlqYwh+VjcPZj35CK
hL0puxmhEhj59fsEyN4mmmmpydi0rPDuufThuDsYGPnjZ12pXYIPAXacYdlLHVYS
BJenJUc6o9zF8wS6F4O9kkaYJ9IIgprjGUxZezuVjinjGamMqk2Rq3+Kq80zGxJy
tWBbTcBxpZttbjTAsGee4hMGmh14TB6c63oz3HPfxVzeCf6qp5/iibnQf3xaS7Ou
68Mc1mpHxDGFzjBro9To68PV/+FnhVCczZZ2wdXFX/EDTzz1CYY4KpGumAUrMWe8
eHNVl2/PCinBVRbKKf75vNIAAvtXwyNo4DwkfZi1+JhwucoaADvAADNYNAJMbPeY
Et6lbCKhE03RZwkXF6+ADW1piLhdcW15qSvIo1CAKBaMnjRHG6YOZP8wjFL7LVu6
tCYR4e+/hdaysvRd3h1rHI8K082i8QB4viDTMyQGkDJxkrIRVTgCXYcA8GBvCem1
Oq1korS3WYBYllvpcaLvEA2MPvVuCZy8LhLtQzU9tacZ8dbTEC4omqQiOKePwKvV
t2/wNkNtsU9Q4a+aJXBo4wy1Tfw62KHihBV2AeLSlNrab9qhRWhMTJgtI0bVBSIt
XBuf1GpV3JUjSY4+9V+vsnzLKVU7LRYAJ/gbQ60RyO4yaKNwYCJU6oDG4ng9lQFj
oizfEh28RvF+KeGuQvT4hWas+Ef+HuHehh5jxkZOfiiEk4u56zXDkd4/a4Yybbw0
t1WP7wCFZ5O9OxksDliKJBZWQiQqSD29BGthUxXLCJtMNOXCmU0yJ8M3VDgmMxUn
o2pYa440e7u/vTP3TMl4BhQBNzPjItJFwypwAtHGK8i50FXm5fWWer3MLwQsk7X/
yW3wvYkbFWnJZA8sbf9EmO8iB0FtvQRv80bxRvJOX8Kec3sVawNCtuO6ODkDxdCG
6LYRvUzaWBJHb9kA+upaVeApCQentd6wQQeCuLaolE41p7e/rQ0+hjRDymZhjKUZ
QLer6LrNPgDmmMI98+e97b6j846GjYffTB2osWfv5cWZPSRaTwgXB7ATYzG6A6DX
h2q8U9mUM6IL1/bIvMIrRgcibE+01L5uAq+TV6MhYh+82WVzmyYQYowaZA/11rC9
n9eLtC1LrRzrdSRbJ91a89/lnVc1KYtNPFg6AKty55HSjmwoPbZ/VKUfRQRO5UPM
6kfK3wN97et4/01VmgqDAxO91zGkk9WOI2r10RJI1r/8Rdf/LhDr6leNet1Y2Gji
n3tykQg5psUs28flsZWlEFBTFaC+oTpWEkyW8/+q1KYKvSDul4ga4DMd2kiPiHPY
2NLJG//b3PPnl+jmimiFURWQ4kxB+XmS8AXs+9T41JkhawSrfEODg18k9aicMY1I
KzME9da7VtSF8RAz3cQFgzMJSOqFCrCvH0KcJsJELFGXkuj7kEfz0yADXtZfwYko
/Nb572PtyzPpfaLbkMtAU4wcgC2KvnmmRwnZOT7oyNUxPbt9dOMI10AFLCtK8qeY
eHH8CFNAXz7Zw2kgruwJmhUT1nqoHX65s5xcM7VbdR9NGyOI+uEUpEZoHOXltFrr
BWoaA5tEBWlHCpQri5E37e9DJlgmhFRGX5iOSF3DcU9Cp9P+A3KPs5GO0wP/OrPu
Qp1Ar/tVlkRBKrPAuwm6D/h0NEfCeGvNZN0+ToZOcE40fuskVpQZCqgqDsAyq0dj
C4+PgjYKWJE4nifZn+fh9jLdN8yqDT2nui5Q07FukjH+J/rlX8tlpVJ8/A17radg
PEZQJOQtMvb/nW2cV+LdPs36MOUrY01N1T9z3vPUjbHRn5+PwRJ6XyXt35du/b4U
KCDRaCuWE6qkc4ZC/W+mjFtW0D2Kcqr1XT0T4OVz+0BMWKuBj4Xmfs7lREk1QQi0
vt5wPkt+F+u5SrRkDeEWDxl6jieCwXgqG8JB8pRV4oK6wfrKdW/RTW47f0b9D3A4
SP+06tOtwjY4UPVoGmvdM2sEOsNMgxhX8lKvVzq5GY/gEjE/Yg/LLyLky080ygck
kg0VuGmjXa5rPlmQTm70LPUewb9hpOz+ULIY/vr95PKHWU6aICh1M8Bvs3LOIMwH
hifQrKQ95di29FKcJjamkY8kRKLJKj/Z49uVidrHhqsK2z0JePT/zywc/ew30B6P
fBQd996h/mTxbqcpkiMOJFtocw66fmSMDodWZSaWSDXZT1X8iAWSx3lWK/iFflPW
TT4qaYm4IWNix2CU5iVGPcqIuYgB16S5W/jHO/b6WQmse91LFLQFCApUPIAZ5yD9
FKJZxsj3knDdhDItVgwtMsdhBKz7VsrQPePHtpjD6eHHIWR//ihfIzjHQ/230K8B
ZIvNRxvXrWkuhi8lLHbB83tAq165t8cFy0fkviYmdWbr0uY1oDdNpUxlNqCQLZxk
n7FSFspdUnMTeoUyCNMsJMtrGd9Yh1w9fNSVaMtpOnh3odLCHzvSsJimDLD6E2Fu
iKn6M+Ek3RB0pSobRaAiVW2ho1h5r0GUY1Ht6AYM/wwpSfnNf7Lpxr3kkjWUy9Qd
6+S6P88z+G1DfqHCahCAtGroD+YrjWGqVBA9r+ieuHeRIAfoeN+5ghgDj9RbPEvs
AT5/Ln2C7OXz8Tu/063nQ6nRue+XKsVP7symivxbOvqJOdYa2Mu8aIgQV3HBsKI0
BlN8Yfi0KAfRsNiXFIdjZFzn8ixgNGxGGy8AtzkUPDSEWZzwprAB87wUZFzxlnCk
i9lFFyib31TNhxKfLxdZQj2pMdKbhE/u5y8SbfNAYJmfRzM/ga2BbZ/CiWca5Iem
VdmkFzqaq1vK7DnfowdmvmY6i4nPAWKtBrmY+6ItmSqs3HBxY+Xl/uSChthRoQzZ
GcEDHEusn2cOcB/eBjDL/7Qmv0gkVu4oOM/4rtZaEVPqSy2OaWDgWzlJgEPd/07Y
Jpgk8QvJ0POESC0kidRnHd3l7aBDEHK3/zw9tCwTbjNtYMrxbAWgzV/ki4XzbGYa
qWOUOIjn6E6zkbgIzXm4y4xkHV+x1ljzCHr2jkj8rNHCyV/1jiR39Q0SDwqmct6q
7JYjLKBd0gL1jMrBo6gJOmp/I0nvpkF/eU/cNCXZFwqRW7IT1xhD9edKUwrEpjY8
xXZsJq+G+Sp1REIgkm3icC4QITE/F/BtOytTINZspSgsSo0Ovqmac4dYWYYhi5Oi
5VMHxaDrsfmPbX54S2jbWMa41ZXUA4XtEPQVxW7XMmIxaUYJsXRrZAA6y/4ziwVL
5u99oY57j2/Kcb2Qv5srnIrFX5A0ZAvP1EhzJOGjfg4NYVwojUlCAXZJFR+CZnf6
wRtElkmdLLQC0scuS7tkROuFOgtuUJ1+H7frOD8GgD1xXJ7ICvwK1P7KW5avWthM
kh6ks5khYHmk9zaglWHplxQpqqYSAWc0/r2AP5YRcnnJBI0ZkyAtNNb1FpkzMoon
2Fj0sCwacGWsigEb3ToJ8dwuPA3JDSpJjYCxBhiPUOFfwZpGsBAWu7+9XmmjpMw0
n/14zsBC40eEdnVUSQxHnVW8MsPIn0vSw9ZSzw5Tje3u9p7auhW4/0QtJfmvpvHy
++P84buXYecsqgR3vcKvUOQFTQ/uSpVwIrSJkOJcp/b7uVFV0CUW9emXbarLC5CF
5QhxmqsYrRsN0Ob+0zJWsjrHfgdZyJ2otU+FxC/vMfoqR9wJkzckj1kaHZnxw/55
TzB5wCuhEGtIGTC0iRA5fUZSl9qn0cMFB+/ZMhxV1Rd+rV16JURZjhsfQkZo3/KT
esNECHFKkwiRPE8U3Vj/LeM0cD66lmazhkiVE0CITANMFicgtE887ZOOJP2P03Hi
cXrvlpnvmbOq3h7fZzNtMs3e1fEDzZ8i+RbKkSXbxL51Q4Ug2lImMGTfZ24zoD65
zKCriu8Q9qLkr+wFHeDdtv3IwxSeZyULy/4eXe/ozgwfBrg2zIOwv4Wcq9jRdWit
7h/k9aAJs4QGq0C0fUm1uxgJ1OekHZqmAtXD+Vm3hwYmNhp8G4j1TMhiob9CZJj9
iIcCbePDlgHxEJE2RUaAXxv8R/sCixd9iedrNHpWn91GjKTt3Z2aJ1fXLoYB1XMr
rWxW4vszzVuzuqeMmHqUvut+lDuW9NdUgOempV0OJhxAL4GrE3t6aMELL63cXwEG
keY5jr7fxuzn46F2uhnTFIiSGltNIVwGzKha14HA1aMCmGdpMsIHFxQkOjb/mPRc
pXQZygnuywdHjysxTMCmRaqlooUgYIvoyhNZtHx/tqHJ00nlGGpJMXcV2QspfIQB
v+Wy5+gzQOo7ijMRU9ktwWEyQCG7cn1l7ejwT4PYOmda4VLnvbXupUpFvLOAO3dP
uz0nZQBbsCKOU65VTUiXqX9UYnx5sXvm1lWT2ujBRvz9sh4RkT+rib5HhpP50s49
z/mrgqG8y2WAr9d/Iozs0NsTnp2cwX2xxJIYWRJgmrwoJ/e7fk48Jwbst51nt7wd
oTgpccC5C4UEi8dWKjchl3L1QNOn/Rc5x8MN11TVwCxDQYy8wF85ACkv1BnSEHn9
1A174A8d/eGRYWCVh/YJiTv405/sPVS+r4GkULUPtEixGUPrBfAdKs7MXZyGtp2a
y3KxZPr6HZtqNzLU2MhROOiyI9PWyP72mR4XfwAMr07/qq1E+O4UWQ3jYGHzf+ze
W1feapWBZn0TdCHvDxEJfr26uIUIXJsazdepalqg+YojVZ3Qkz18jA8fgZLDO/61
a7tiS9MSS03TKqAOX5lrerDzsgfg35SrF/l/4xQfTEkTIpHxb0uxMrPC/+Dyn9wA
3Vx/UP7zHcOY12nJ9eCqr9hJmhHCwaAJTp21dQODOU2JDdhKNaF8jFn17DVRkEvY
0CXj3hmS/BdzZLpbGQS5jqokPlcXmu7eNitPskCTkhM4WfzQg1ld8652Y7+gKQMu
UnKpvzloaVmgyjs3uTVc0cydDCv4VfCoxcexHzo99/pUM5u/95uqpsHUqvOQBNMp
f9NlylPGY2OQ0/nhbjotFzZKoczU1qvg8lKj5uLMb2rCV9Uf+3Ol7T48Ne/pAw6r
HJBz7sz2nkl2AIkmRhgePK3W3N8FKlek9nBbkn2UMlcjjduRNHpE2bMeiPvVTE9E
guQDkZDznFxE9IJjH3CsBZxQGkrMqgYDUyxFS4B7nJY3ukHEb9G/nP0Ns9oRYz0B
BlQ50dirVg9QhCKNvuoVpe+R7Qx1SYHwPTaH5xVt4O0bwbnZFssLaOaPINgdyXPO
WSZGWAGK21HhK7L0ih8UyG/64PfXGeGumFCzbK5sSBBLyPS4BNz3pRg1d2QXx5Fr
aA/LZZzOdlPxQaLpK0K5Z1Uwn+0+aI60FAnF+XoT6pW94U4Bn0Z69En4drNI8LDi
nSwLvDlwUM3tg54SPoPYnndz8DIA4uOZuXB88KzHptjLEgRq8F0NirXKQkGXP/Y0
ibTC7NfggRZAaOMd4j9IUqiqBEyUK6MNnOe011/O0tx0AxmquBLDEt7aP9tgPxXB
ZWlzGG+INCUCyeBm32xkO+RZfVyYulGtBPppULDOCCgMGVkdGE/PUMnpxYIe4aC7
OzFWbbYfN+H0tle93kBibvYqGLkqdNQm4GDYXPb6Dns2L1Ne2wY8x3nMggL2VnxX
DhoKeDPpqayvxj3iTaDeJykZS0+jc/yjsPmqpkD4KfpRmb4bVk2libpSsgbLFK7P
ir18bsHQlG933b8ohvEX8N7m70dVAvd8Y6ipr8OvALUY+MuE8tYPy+I0o8jCNp9L
KbKdnm+H96DoMGyrF1V/OxOA8EkDydMMNWymKRaOPaZJeyH2WeDd0r+8WhwSUJYl
EBvR9mVr/bxGyLejNQN8YBy8Bd+PtFwBbw+FfRTxmaUrKSQDOBdZrRwEQHQnB1DX
iXEe8cUrAi7Nrq5P8SjpafL69wQZ2JL1M7iYO0Tyq/11+rcfdoBNgUQDgTpK3kk5
MJereUOuvxvX8nuVfm1D+f5clOKXPGNFYTIhj40SJDgPytc6EK4o1FFgltqQKBVG
1sJNJ7CHFyW08d/HEMXyZeCJs467z+9wQvwc+yJIWo+9mE2l1wtAxJhKHXxlzrLE
Em8roR//gjEPZe7bPyEG857/tB7ItBeVfIqReX1LPEjwK/xHU2oOPa+R2IdFxi3+
mIgRADi7bjwlhobJ3nWiCiLoffyg9WDrkOIgmEmI1OOqWnd/Gcomw1gPqSvH38eG
Gi3WDhwJnCmPpGBtrVArhVfpinEO4w7ZES6C5GZiWx/hBQeeGJy81N+pnOzOrwPU
fBOZqFsGc7vR3mwpXuiIxQDCo5Qb3AsibfZTgCsYR0tGXNaizhhi/68r0KAuaAkm
LmlJw4dNdpikvDsm9ZjbZlwbG7Bwhx51ngQocZ9khqg9CYNAnnvQR8AXuIhZMHdK
IEXu3NiUg7v1kI2NvZ8Eb2Chn6PXEZMGAr3lb3mA5Y0OaRm/NChyECw/O7JAGOw8
LSKccsx3V2m8GLzL+OHBeOBEFjVDdTLz20hLlEyRpYIfvVAbhku1rEHBpx9Pa3D9
TW0MjRfEix5zVYLuXM9TbptwKNsa9Pcfh2rMWhd3/LwyGkyJNoliqD3cfmy5itaT
0YR1trYtX2sLDYYqJ0bgFTzshNdE0XoVLuT96COHxwImA9Ct3JbeqVXgllUGzr/G
j3+iLrBSLfR2X9znNseSFTtGL+V4nH8vCKqbndpjAocXwzlePrV7CxmGzmWa26pf
A+bDAikwIUw+aBZCFyp6gPBkVfq1FLjobE8AURL7vBwuxVbjpHmFvPIYWbFYZrUc
+3b9kGbr2B6fT/oonQeSYjd9Z3/k9nOj1k3E52LexB08ZCvr4dLU6b7WW55cEF3J
REsBHv4Uk1CsbtkxUTMgcxrWwgAHRdjmBpSuFcFYtFlJBrLy1l2zIkmevQB95kuU
n25FVOAxZty0BhTJf5CRPaMrSyz1Tvx1z2cvNXxsb/JzLWXvrmNb8XHEnZLF6pJu
16skKmHM45kji+PgM0Qit1dOskyge8ZtrZLEpvRy8xTQQHoU46NHuipncf668Lyv
AYFQGCGLP6OO8HGpMj3Rax/nIt05jwJny0fRiXD/KUBKn2+8CSDDnl0QnWLFe/vs
Xxli9lC/R58QKkJvSVvFOcWdefcqrRzne65HdhvR9gcb3YkkF3ubxDWADhkiCv+k
vTbq1cFUa1E8IFsZ0H4QrV4OjkL3Qh3CtnNhoEY7PMmZuVRpTS2cKqnsRzTKyTRJ
yWw5OFydiWt0M3hEHMB42VGPWNnp6tlCh1oN3t0u4LhJNOhN0AD8WnvrYK63UWIY
hT7eO1uvPQypICEa7Xfg4Tmyz5ptmFatJPK7miNUbkV/Kr2VU6qFGkG23PQb412a
CaUscJZ/Riy5HfPUjSU+B76YlR+U61uoyik3kTyHMx1xJ+I+cVsMS2bEI6SeKbW3
vc/N4xEle12FM7p7tXwnQ+ZlqYDzgtop6XDJs0eNtz73taTWDcE9FsrUNTfUghcG
2LsvQwJgLmeW4SAXVjLYAEcKSOcGlKSIY83qD7ZJTGBrGokazdXTmr2SZSpZ7EGF
HmHiAAkjqYW3WXnP7zADlcFHFbD80TIKtiLtU5QJQgGgtGEpgxpwjJhXRv3OC3Yd
eoS4QQOCWsALpSjxFe48D61a0UkXXhvGe6qHsemXB16iFUux3yxJkE2k9fdpWdKJ
XO58IXS66ATdEtoGgFBuC81aciQ3OckUnmhKek/ip62D5b6noy07aG1kqyJeuAzZ
oq3+7YjyCgMzL8TQPSb9/fKdHc8WfpELQqPvlotfDfjBfTjCrRxcND8hSddqCL1/
BmdXqZ65YV7KrN1gfv82HnutGsm2akHNGCE9wEOrrYP1pS3locb2C6ij3yfTSEdl
VR9EkYYEI5zrnLgrGyT78xVSZD5IGp6stfloW1KTNByw94/YqyC/lyGM8ZalbnhG
pfds3oyUGXmvSQ0Z+Be1EBoXWeYO8ndUCxczLqIZqxw4qNva9+SV6z4d8Bw3xVAb
TmmkOYH3mzVurb8qa/0BgZ8KWIg7JcbukViAzShvNXioLOL2gTelAwXmjc8LgXB+
ulIzRfEJ7oNpIig53OtzOjic+CWXjsA4I5AnVOemEA5lXVMDEGZt1LTEGUx00hr2
UPZmON+O38MCkudFFOf/F+hsjHtKsFq4ZctpteDiojkQ+SmnHmjXuLBXNUSgJWxs
5oRySwMWGDwrBifUnQw++dDcTtvBp9t+wtcmEkg7gEN4u4QLOYaLsaYCQ1Iq+txC
vIykY8puC5aC74nThZzyJdbi5EP1AUBJcy9ZMKrBm0E1K7UEQLhZhszRCNd8KXfN
7JPwkVWIQhxwrLemihLYafnvPX0FTrFZxBjun9afzwi5BmDutrbWaEDn68g8Yev+
Z039L8OyqN/ODxQnb37Wxa30PiG+PG7uQWq7feQ5NomdFGsyK4Ei0Raa0wWmYHwD
pevdfrXpDh3fTiLBD2OEeFIv9XSWLvplOTI2Ne373geOMXmTGfZSnxJpuFlpo9Pv
rvaUjY+2LJMkvcFiYIptj08VZo6JC508vHc+PEJUDb5qZCDY/tX95S5Hs0hULrFH
tEdE1brVeuMrhYrSwbpdhphcUY1jgVw3b6XAdxthAPMbXooj+INz1LZDFgEM+IBK
sZJmmotaT5rmsO6trx5X9KH3K4az96u7Q9Fh8iiD5OYjGcx6ok7Ohz+JMb13l4n3
KbmEH3YcWiXXt7loG9CnVYsXIBHkvDoCiCylaHNJhSXYOS0IxBKdoq0MCGzo1MO8
ZTImHDvl+1gvHAgmYxWYoVvKX+xg5NSiTwvPgBdK0+/ruo+NOdgvU34dhZhOc8vn
+erIsgFtmtcThYE3YaXAqyORT6NtcSQFLL9zC0yL8/R3dRl0hTpc+qNH2hL1A+AX
PMWFEr3o5OAY+pUEPUEdmpPFTR5sxIQCG8h6sdaBYpNhxpXyUBaxVyePaazjth60
ur/mAJuZQerRqsxk0ueN62s/5RPz/yES4w9FX1kC8+K3bcplkjFD+fiWSqCdj/La
uRMkAdfzRF50N0lo+obpjh6CgK9P16Vxwbf4wjDgFkGuOfxMygPKCJvbHKirltfU
IIXC2qqZ1IlFAnDDYrLT1cY8w5UT5qIFP3BWadRxqcpxdEqK8Z4XDCGAnsu5WiwQ
To0g1/OlqxLiDtGkfhl6iE0nz4pAcDnovF2azlHlGiKdwaxq8xY7OqKJf1kA3tyc
5Q04e64s9Ik5rNndj+3qF3/B9GENsGLUWDmWIuC1u6Q+mED+OGh0rJAW3EHsaiK6
4Ea1DSN2JnNGNQZfSyKS+Uaz4WOfgpOhRSizo3/yydZ9S1E3nbK1/WNm4gZrGXbN
7F9mXFMSg8T8/K5YpmONhIXgf2ZF+7H9f3WGRSaeo/RLYFHntA6m28gs5feMVGWE
fcSIl73iqqZAzzFNWEBY3PvKIZhzspHZ9gy4yMwkjZFjyvOq0McLcn+bCIAxQ23q
U81NaIekFT9+IqU0ZUkevK0KUGVjwuR9qApj5UFZ0ZpP1ukVt2iO6UKAvHo8T75y
jJxy6YcMCPEQdS3zFnLHYg8s3hiPM2hwTcaokdlFXmq1oucmm3FJcv3O/x9O9F7u
xW0ohzUs233L9AQK3Xwt5b+shDgCqGCaEL4RT/1jMU5w62QqLItQPxwl8KkBeCt0
lkv9+bm2ESK5l53iFXIfiKEfaMqYlVfE4G1cRLdvuOVNreuC0lKKBwKMfcD7RAQF
211z1SxlStNRHDky8097o5ISLTG6B+NDbu4KAlWuNtyzcFS3UEc82RwL13XpkxvW
wqt91X5EItxDiwe4Hwrtm4TsuXCBGrVA43GKKSdl3AWNCtr/y2KKOT/YAVVjuOAL
wIEFAQM28vIgPy4Qw5OTBXqfuVBSuXbolsRKAnBHRDdW7DgMn8+XGmoHMfUSLyRP
gdpNkj1tt1/Mwl3Gq8Lkl2GdvEiigds69oLfOHEIa90ISUNthd6Ux5kAERm8jt+r
83NQ9QnJd8Hl5gI3fFTkUypa0hvcdG2QqxzLJ5TjCVlt0khF/ox7J7Jbkqrj8v8z
HFHptTUBF2C7WqiqWcboElnE5trh4LMeojAnLNiUAm2EfmRIz5MDPUoqP6EOgFh6
cmF6LChA2evEEqexigj8TIMLfnmyQUshIs+4dLASzjiLpotmOsVHoAJtAshB8lwW
ME2TkwvEoN6FaqmykElYXQJaG1gTe8PgLsSc/hkacsv2N+uQL13TYJPtDv+dlrZM
Gcv0Pt8IksPUOWzokH5J13c2+j1pU91/CCSwyIVgaVfZ6TDzeTm9vahpbkMebdbV
RFkafQ3gd5yLHkSMfc5L05UJ3dFGhd+3MwPH9wdBaw9VVeniV0taNmA1mHZKyHf9
RJmWF6CHGW++L/mqtcpWIHqao4kVczSYyeLM8RQyDCF10ycDrotacpuipya+vh+/
4zfZOjLhrm6g0PHiosyfsB/Euw6o9cvvzBVsl/coeCmt543GFxtZWlbrPTWfxffV
wJZaEPLEY7DIPRTGyL+XPmATDKXgaMGUPPst/f3RI8pkw3ykQCrxUbsS6ERmdmOc
xwQFOv+9ielf6k0KsTC+2Lp3b29OpHF/XCWaOpZfbyA7jGKF+/SfpkrXEua23Nm5
OYP3l4c2zn22VNqH7oqvO5ewfFgMB9fmFQ30BWAtV6tZJi5ZXNmzLvj3MN1aPgeK
8+aqG5VxkPZM58XE5+RgPOx+mxUr6dj+Bj/jT7FWGV+MPVgQBvZw/32Bt+rfLGKF
bppN/Lzotqft/2RK4r4bW9aiLECnXbe6J0dllINPLEFEPcyIkHOL42gdXrbvyMoX
SZ4GUJEnvfT2NMGEupyfPrB73TY3FeBTcSScDq/7so4Mo91XurPiLyrjESAxQxUP
pxYj2Iw36MDGafSP0RI8Z3pOfhrzOCGfPRRKLWMe7ZsNieyoPYTwlB5bWJQPWX/C
/qHdlZVZgtLC4NtUn5wp9P1oWAYIodYJJ000fGruAa27FvC5w6IVDrlDUX9J601Z
f2Byqgp3BFVF+LylQeVBI9dnrucaUYpG7D/RqCfWUgp9jM29y8gsOOrfzbeZTyp9
T1TdBFwdldgbsT9/477fa6G8kKXpEEweMeBKLCh6Ob6j/XGNOGfkfwklFmQvD43N
qg6YnPfXlo28lMf5ob6gpk/e2fqH9Z8B2u7ViZBndoL/rGH8U94vFu0G8cr9NGdB
pRPRVNPY2OKblm0uQ7FHkKlSiNYIQfSk8DDSbZqo75FvpvUaxsOqtVVvguKD2qyX
YXKDF60V5DamTKdk71y2nnh0LifUbEeqIownB8D1OqY0g0dxAxXaW4lJm3GQzGG5
P5yzTWwfoYVdqmGbw5mMpfSZvypSgNyboWwKgwyVIO/I+u3IqManVIy9N67YlHTp
RAFQrDuOZLPaMBFrCmBmSFdZ++gCtbfGjLbuL+DXaDRgreoPqtnrapJM/vZuaMwO
tmK4o21ycuM986M6NLUDA0AZsyvb8tdcawUYhtP3Mwqbq+YpEo77Uxvc+zgYXxso
QV8wGvX18uAj4bmsiBJfP0a/rHZW2TCHKLeIyNXZtwadJWFg4m7ua234ITTOMuPA
jOUVOXjqOxEdvoROndhJPe2NPEsy2ZnwXXUgKuryWT1Svh97PZoUI3jwol11SNfb
oZKyi2ybp6C7d7K2BMmdcpmUdEvyjM7TzugbDWr2AtOZMvElfXEfeoN7HpfgoxBY
183wgbu7KwQtsG3ZkZh6vmYWHNven3ZFezDErqBurkPYnExA0ELZjkQz/o62QN94
Msb0T0/oG5yXbzIdrPhjbvwS541jZqHIHRcnDP9mhVwAghmFRL/uqxmEvMumUuhr
c7dlaKVzaZFWURVdhK0TUesj0l73ReAV0WWw9N/WS8zPed6FrtRA7ZCDBt3iDuoY
emkFepaDS6wvg2qtdaVYg3GCVhIDs1IU7sFNfELtnNgvsT1mKIMfmzDCa6NsovLp
Ki34SW7kc9lUhRu+6LEQYUTj4KNFR4+o9dUkH3nmTT4OKMti2Xd7yM1fssfnqLd2
gN4lCwwHbLdhfE1aMPUDvbSHXokTe7IHWNUOtVdm5H0PdFN8lJ9RbPJsI5WTrI16
/zlwf6pzic5hli1mIeteN+kdOjLAauOqj77Z7gQTbnln0iH0xmK/CCkpe5QZvWGl
yl1H+Ay3BewHYRtK/UQgiQQjtS8azcBv48hjnnAtitV48qQ6DO9B8THdOeSPfaY/
UEuzS1uOFSbVXs9QJZj3XhFkLn2Z75pt4+EC4O/0m8DCQXcUbgASpt77XyDvV/0g
lhgXvZxC1dsusN8Tfm7VkbxAwIX1azByqiiXUa50WCUiiqw60otTOVUDpATIPr8d
AFgCdLRWcOoLvcZRTTd2sSVZEfiy3bClbscgICLZRmtWc8C7hEx/WnPX+uUMemM3
p8bf8RuJmRHIQ5BuzKTtLCetA3QioGtpErUpkP16scS8u+baiTp2Ux89SeHyExof
yjjZm3CSmXQpJU4IaxYZYmErfw5Wmot55gNICwNwoiJKvJJTqWxqmgwY67531d1d
tZSsm4ZG6rnqF8K5mbkYbY8Q1b2AyG+s7e/t2bbmqJUv7xUOgHytG81E0ObgAlUv
KJjAcLEnV8mdB9qjB71FAyjn7VLGkuvInwdx3F+fatTci6egBgGjmPlCuWikNAsq
6A7NHN7DFZx24f53dQQpl4X6Vy5/xMrb4PFNUojFpf9i6wfEfsEfzsOCl+g2Q6DY
M29t0I86/3e7pDlb1QPmKSMnQKpv6+xARLZjtDtcKU0YZpf/x6iPuBCLFARAFfm6
TUjYMc3lEXelresALj7/8RGZxSNP95iBO54aunrjHRapqeMNrzvfE38TMFo/9LWf
YD1TtwQVwSipp2bTl0kX8blLC1BjJJnMiTMD0yV0czourmrDYM+WIcVjlGuWItLX
0wYhXRqyxcOZTQ7VScz2lq0apzxY9NcItKKbej33l9+Z3lFvzEWlgrwletYK7URc
snD4Q4t5ngvLHonerkb3rTKBFXQsK3Tgfz2UqIpnzbO4yce+tkA/rUHoCegUzJOr
1PK7pjuN1Bcbyu+p8w3sxrHt6X9GPtYUjuVHSi1op+EWsjtq//wSKL8ZwzKqWcJ0
Y8lgY0VWcl9e+FQSN8n55U7kpgmwtvtoPzBNe2PxPzgiDTa98TCFvQHHtkHBODwi
IZKgM8TniTh4XsE7InQqmMkNk0zKsqtv2L8gLvaGmSAeRY5TvYo2Ot0ZjxIs9O9v
tK4TF2bPoU+lDqNIrqLeecvWCBvtmkAbB2KDFIPvvzIRYSSV1G1wpEglPW/Ksqox
ZUD/tc/ncX9elMEsVPJF/YC7+RTIgm0v2avmYwxJfuMAo7joXOG1zOACB/ktRasX
3gdrVH5Wz9WwM1x7CXCY0izbNmGd9J42pB8XbOPD9bPG23rVJZzVeAuhaCKsCkWZ
6j4k0yo4G0mXA3Y1/z7rBOlFtXhv6kkTtY3NPiXChHvwc1FiCT9bhFYIfRJ9SSjd
9Dhry7/ecKsuP3LegiUYx6CRohn3IKQl5FeEwfwasvPzzbyG7MbBhnRwySFgrzAL
FnUA3j/LDKhODYGsnIOQXo0DxWrhvRz1zcEGKHe42Fh4qvZhGchR0YDQqtxBA6BY
FdQXCy6HkRczouB7HahVg9rEhAKpJwoGKYBsHoEX/tsajlf8fZxR2l9r57nk8dta
gaVwiLv6A6fPioBt15Yih7r67vnlZD4wGRQEzXZVlwXq9bmoOOwjQboMxQvFCIJF
j/a+Uq/170S3J48t5yIrBVI+6K2MQrSgei1fRWf9VejrbL7KLn7/UZnig7CThVpy
VB74DQUXgY1b5xFPThwc0ypPyfBduVzi77SqTT8iZmOh/MO9E6JQRSHx5+xN9ufb
g6PpNuVsVO+4CwWWSLg4k9+yeYKQtmMuDVfnqPzAXdFDUXe7VHQBM2KLHR3JWk+W
UgFDaf6xJvTCb9zU9vesZMSRiS72uFyIKfWnsayB6SOpdFXAmFSQYo/apRfsAKwF
S3dN7/1iPal4lzebssgGaltp8xBrfzFeVr0cw2yO3H3OLgOIK8Gwnba9hUq2Pdu0
nSTACPTHELbt//p+AOTp/FdWjwuZXAmaw/mL/OsrQB+Glhkih9rhTQjMHj1z7gBi
INkmWDrjKUNoIQZTklqWFz+aHWy3eMxm/EYdRdgCEq1cbIZwZDTpDo8qpXPuYnSL
MHSvHYqEiCDjoXsy/gvv44qvP893qVF9Yb7o0esTrrP6I5A6g7gKN3MCGQjpeOTZ
hVxbPnY4YNFF7cwkVmljWIxmlO1WDQUbOJr2uTQ8cJKE+Xu6mRA2+xwE9UYqeLv+
af9o+sqiBgY4kbtbIY0gY0pPog01q/bwnIrJlRDNu/ugQZq0peSkE6XHjUTj4RVY
nrsLaZkxPYdOHbL0+1e7Zwjx7yNMzyvqQ+4lxzmVtOkfzWnmxsH5p8Hvy9ncJRdy
CQButpQtDBeaKaJnUzHnENZ7gC7DDk79QV7uI1RCn8VuoKCOFFA3Y0e4UEez+Mho
MbAU/mwZGEhM40/sQqxAU9VmFpx4RViBEPA7W1HtK+XfoMWSmh/5V/TOEfy0jDcj
BdJd/hvSt+rOGx7WDkXW+PYETx7yM2uoQXW4CNbYegfj7Ixq6H0UES10vhnog8FF
OsQ3vjNn6gzemx7qO5u3/JaUh6Une0rlX9VOMEsXMsXy3+X94Wr3GpOfeIws++AX
0Dnb/FJ/CXxCB+qzx6QpkFnUDrvYMp1MrGzBRCuzPp5/hGFngtEYfTGS6nGmLR+3
Vf/9pO9/ex898hqZu/RypJNxaFA16eTOumPay2vpI+hsL0PnZIIMeWTIziNQ/KSl
oDeY15srxSquD2qVBJ7SCx/uvXxlMf2P+3bLcfqgnpezLSmU21g3DHimjZC3kA3q
b3oSvTFTgeSw1HoiTNeIX1I7lAnHGQgSVlsItkzvyqTobzDwi52nmKoqsHe/iW9U
4fb4o5L7hxCflfOHRpz6ry5Pd2ok6MQvXM3VAQQ3tW2rzTqlifRGVmQH8u6kfvUY
QCXdmMGwhOONVU5MNqUYCTjwSVYNM5uUwXf1+BAV5MEBi9QNK2TpDDIE/KKUmEeZ
L7SqTzDV71CtV3EjI7+8kEMjHF3kbEzQ859qE28zsQka1FFsAW2JKWIDnv7AZIwT
YvaT3jvHQzOh/5RxB7Tpif8ZRw0L/y0g02KX7tocz+oLK6NPg52W09KEh8LxjT/U
x5SjkiS94k1uwIGHBLgQS7f5U0yjzm0GxBNT+5mxfTUlAplbfHitwzu2Wjvyd6Hl
wx3QCCHrqnzReLQJqz4P2fsmwlVX6vrGvN/gcrWfXX/Cg8JY2kjrYAK6hYvbAcry
0+I2hS144taTiqJpeQcrJgFgu1hfooWOSLWEbdy3R4RDlHJTXfbKF6JIFJQnl66L
Uz0vvbJDD8NOS2wBKgektlLN8O6udI3pRQF6BIgsAQ8/fUyAfnZvUnMXWqOg7nxo
P2FqYxWCskqO5XnLOWMaf1Ul+2GdrwgtGvOIPWdB8eGs0/SSKQeVCvx5J8O4rZ8b
yoIb6UIdt86G2H3rwkq/nkdyoMpqCsPuAhTzal9+dYij5QghS/+xlV8V1J0JPdyj
WBpDN/Z5hh2EQ4aeYbvFmXJf/YyIjicbzolCCmZ46f4+ZKjTbJNn1De5BQi/CtrL
ePdKToTwitd2aXvZGIQbHZFIAnXTrqvFfPGb18jgwysj9A1jEiO4JcgMVst7fj0g
+P4ab6JRJXIxgQiMAnaM8HrTt4VXQnl6LQQgG3Q7cykKYEkzWvLej258O0YfiucX
CgiYI7Q8YvaQBKBty5+5Qkrq8oK+UCQlO/Pv3FQkK6l5HJ4SBt0g+F/TqGcXDoNB
+EKM6oA8sQMoSyJecdNWa1VQTaGo2w4Q7/Pa0Mlldvw1JP5hlQCSW+JE2Tg19nk3
Bn0F8RNnOocK8MdV2/iqIsuOtSXXlkc+gALH2uis5etDQg9iqGz6TJWxn+VuLaAK
ikEWq38owuby/LUdel7eZAGztFbpBwjaeucYXpjzSd6iAD5sD31zSSKBnzeepycO
srEohdLF4i4BUKgQPlJoiMmkdXb+1UIpHW07cUb9ECLKVDtQqP3mAbSphqHHN172
5DTnFVLFD6ACkme04Xo1p+dR/gVvFatY5Cb38Gz3goUhKRdjRGe/ruN+25LDs95J
XDSFXeI4BqT/vTOdgzqYca6HFgLlMC4R0x7ZWOjjLyt+i4wQbrfTS//PgMGciCKS
g8MfFX68cQ1pgF++/6YLOpzRJvDlg/mzmrpr9Q2sEcjNYUpznZHtgC1EemDfWqbP
yv9lzU6r7cnevt+W1z5EVo/qYmrBlVkCHmilC6zqwzq0M3YrqGXC2mMMvD/MGYtU
lPXl5xSwts0nW2vqcI8sMLA0XpphUs7qqW3AhxaPJQNgVhm7JncKcU4XJSGouzEz
2AO7grNWp611DwCrkxwGrHvgjUYZlzA5NpCNv2/n5hYE42AhjCdJK2c8J6VaPao6
wx86X/dI2LgR+9dUgOBz8uACo8BmfILK+subD/+GhXiAUVcrvxjAkt79MQQA6JCa
KZ+xr1wUb8DPwmRpVRDaZAifw2wLvZ6PtgxlaykdEmHRYfYtwAD5HKFS/qcucoVH
R09KoHlUVO3AHJpct6Y1OTSmyTi/6wJGL8L/fZO0B7dxpmyJqZTg1a4mlJRq678B
oY4spUaRH1aesh8SIGYQgzTOlpOOz9IhuyTGaD8IJqGV8z3DS8xhxvXZFLaUlOEK
TybpWL0unJMR3pKpxx1WonG16kEAabOSnzHoxOc/WYM7KIqhs4RwxJg3sKGDg+8O
y4IqrDhwj/uAWxAdrdUwCO3XDr82LQyG5JwsbgYCZEaWP54hTF44VFZQ+E3kQq2k
jPij/7fQ52svTXBtv2/RJZAUliaMguH1+jFQ/EMEfB6mlFbqJgSjMS1EHOSFUf6Y
Au9yxpNWlJMHLC/Wze659TUyXQl3dD4F2fRlUvRZBhU0GoIwDcqJPz542qWvTnei
9z4UKDdzJv/dN0VVSV1YyYbuTnDIvmG+WLegnn3gDE1lgkXMDBjXw2zAFOsy/I60
UVWgr5nhHkXAo91sq5mqG/1aYunqyIyaF8R8ixZ69UBEflVLRewjEiLto2Tmlks6
QNPtt3uoky2aLEs/W8XwmuoZLbJOp7bOngbSCWITe7JQ9u7+VoE5UXyxnfjnW5BF
6rRDtCJAr3HlLrK5H10Xf5e7JwMpzI91dd1+bYW+YzH3Cwd4EW19Yn0Vxdi7I5Ub
j1Rw+mYYRtejiSoOzqjkFK+gBiFjpphjLIhPLSx1huiNy5gNa9kabPOQAqWGn368
y+4Rp57h4FictXa4p0jPZG5xtGjqpTsGGHRLpHc4mjMJSQH5Ry6KXQ7g8kHOiq1y
PayM1E7lHYiDv6+3p5SqjBUD4V3P0OSCMa6g29tD7XmvBcG6SGH743TxAqq89nRa
6IiZ0nvfUzdDsGeaFO5sJkT1c9PNSMboCbL8tndl5szpIwukfzG7aQYWz5Srk8ek
47WqVQpsVyg/S3Ne723VcWUenzTRMDoQD4k3WFyK/29dWmi2krzjhcpuFODmu8VU
CnD1QWt8eMJkAe1LvNHsIgrvgLs1vvJVxweLblJvFeiZ+AqufJOIg9+nOpglEI0W
R6IhLYWVouExwO9ZjPqeWZD70KJx7RU8eKS/TlM3QsInfFQ+8ZDgC0AxNMkQXos1
y4vTepSDwnUW/R79bc3agiAZH/XAmeZsf3fBGC8p3+1uEwHXzDCo6B7zi9NRcFtD
elwKCGN9FsXYLrQvR7dKfcngF4tTHIt8eUhs0tESMVWfsVV5Tr008sSO0kXDbRN0
crbw6KpvSsF4Uk5vhofWibAMZrL50IP9aXGDkPRjpQNE1bnhoxeCJ2ISr1vbEfh9
/3WObM64rmI5QRpmoGkfjdg3pHN5c5EO7yM8tSjDewAVXdLHBcDcyuln1JzQBYzo
ZTI9f8UVlfnjoE0KubysuPjPausGHAyGrYar1n1OTC9OFQd2cijuUIcyZV4zBNt+
U8lZfUtfc2UMDuFEhYFzbArCjE02R92jA5Yv5eCb6PdQSaZbEFQ+BycrkFZVKjFt
GiM02UJ2qKrTT5OUGpWd7VZbElLGtRX8tx5uSy4AVatvM6dvi0oTPXM2dE77RWzl
8xtdAb+nOUzCO2d4zYRynmYjOM+PA7PcOkb68nrcGvOq3/3Nph8+Gbb6m0MWS03K
g+Wo1wba4YyayMLwB2jfrxdZvNm0p8ni+Hni97LkhFTPkYkzFSK8tBvTkZOMyFjX
VRkU1fDX2dBgBczCyRpy2dO5F7GCpiD0qBYlgsoqkPrvl7lolGJnQm4hYr7YH+hD
FHxCeRzIekqtR7+WpBQdOHPrgJfAH3wdTQKxGLtzJ6FpvoG2q2giZumE52ALd8bn
BnaLOSploy9TjAEk5+Wc3D3Cfm8M4K6lHOE32a/smyoWssKKXSqhs14JAqYUJ0Qt
CnDNG/QEth5fySLSpe3YAv8dQOuJGYk0MAc6goimg93yBBmQWcvHCMzrJu4hQpzB
baiZqCP+ZEEg8k/UpY9ZIclLymWuD/OcYIqA63WisNNfcYAQWH0cvJ8N5pD9HtwB
qI/u50uUpn87pWif7BTrfOGw3RFcLALFBYpfVKBMncRJvmhtj2Qs8mkvAh2Fjc0M
lC7vpUxbnKLe/ofAzlIQfZLzigi/udv/hW+8qC4kWvGvpWCB6DNVKxO0BudDWqtD
zdJZO8+oY0Zt7q8s9isVDNs3VVow/tbPjNbi5fiE/nyCZCMQWKpZJcUHlk7fclco
oSbUgFqXm81QtpS7bTVqIwMcz8gfNInY8EEiiMKU6IpiA20xHVnGsk7oyIBFB44l
r93lBf8tkUJwNYSRYrsLY/5587+UiozvZ1uSFUyK5sgRG8aZ+pjyDkHiI23QAVJA
maYmkYpSPm3H49g492/n3P7KsdJVu5wWpJKm7ZUCZGe9x7qZTSfCDTabUhR5CBPm
XL2Sc9HCH7FJinnxTMwgiNjcH3i7ETYUL2bL3gkk3LR5xCQWXZWS+5w/NOHmwAgp
fCQaljXuG8n39oNhBRui94Rm5eClZ6alhsFl4GypeyEzzHDxAIyZvb9H8rOS07Td
V31c+G0g1IXfsuhFMrzv9BEqD29hZRYBPV8b9cwk3Oanv5D8XUDdKfXEyapS9Tzq
B04mACvFryNxF/OKeHFZIGbYYiB9jo5lAXjd5Dn7oADpBdYUOFtVZFYxlfAw3pRl
oVh9XYAGf7A6jJpsuTxCBzBo412+Z1DPJnkropZdV08AyPBXgMphxZCVjOVfJ/XY
mNR7eoT9DwgvsTaWpv917sHyKYbA0Aqegqabw0lwLVelLLVjkkDkfnSeoMi2+Ro5
1NvmFPJv8UvvLIa6GGPbohuKXDUnuMCJZq8yj+uhka8nKqLOFxiL/j0gQcdTVPvk
XT5PYMrjcQA3kDlYvB5/OFSrzfD/ZuM0wrX+XMIjl5llJH1uyTFiGinryZRPYcTF
Z4xeCpLcxTa+4Bvlpq2GYui56Qq6IXmz/KYxHY3edUstx3X62xNE8/NZQLPy98Zo
E1oK1TzxRfNFjKNzy/ARygmMKj09YU7+qiN8KcBdufnEaTJl7cVVpxKh2kI3afNP
xjY0UpcvoTbjGYM0bYCdwTSAZlNkSDfCGvd3BlPqc8/TzcQPQBvT2b67t/N4dgF1
WABHh3DtyN39fBAife4QDjSthgh9Wm4zxt7ACof0DcBP4m/nbX7Ju+K5uyHz1JHU
y7liREJ0mRKEHtwIKUl1imYCBi1LKO3Ly1+VK7XB/V0kC8Gopd7BneWAaxFrxGYU
8dbrfD1L6+s2sde6UeH4C6/e+O/t3E6cxlDpkDtGzQHBn9DI/Zt7Ikz+SKj3V5Vv
ywFCD3LBApMIhJHhC3wtfx5rbssx8l36Y7wytqXqk08w9XQX8X0e1N+OymKRRtcc
UnaE2w6lbhha7cxrcVP+oDxRFxDjt6vKCP4b/8SIt1BJZpBOEeNDAhRd7ut8Ydwd
1vpj251U6G1zNECuGynno4RKHPr1K/C+WXh+9j4XMzI/+SCuGDxM5Yyywe0WYN54
vm1EdDW8jgr+vu939hbmEY3eP6x3w7fS2OhQ8hsO5Xeo74nmhOz99bS07HCD+5VL
Oau88K5KtU7Bz0dQU7CEu7ixjnyypNnv0GMGwunE7nH62Yphm4B2KzDdv92BifD1
Gm3IPQ8kGsj8+cqZQwcvaulLUX5wZ6s5fYIDwPCe6yVERcWRAua+X+SGKuUId9Oz
QgrUeA3+463OxnFDBZc63aQ26ytpGEmc280zy1TOK1Jt6Lu4ghGYi2gS6Mhbz6mi
vPXEkizX2uwZiquX2PSTecFMglcxu8ZM85MyR3DF+ZnX61vco24rFpKkkKiQ/iuH
Z8S/x2ZiPMQq5qBVdqJJwEFwWsmyUUG3TudRpg8+nffB2sRymYs3zdaQc/oG/a82
cTEnG47zk97lvIXSfo7iuucqLgcbOmkBcdy7alEhndR+LuRgK1tXQ7OPMd7er0dc
uSQL1CdZwK3izmX8vVDMd2OAMDQQ2MS40z9OJ/m1Zra2IcKLhNQahTJ73rbO3ob2
zP0RdE6R6H4lDYXnXaVi4Ll1IVlDsMsHkB78ET9wxg18FwjuwkmCiNsXNZK/R37X
AQfyTckOsMInoCN6Mw0ohqqOUea1iLgK4QbV0uasNNt8yf6T11vufTEiRi4p3ecE
uiKLMg+MeP4ckVghBhbEtxMYmD6mrip5wDbCp8+HRV4PJQSH29CO2/NuJQwC6Jhr
YrvQ9FTZAZTX30X/93znXOz1o7LqLPs0ECJDrVd0NTg1TlKARUNPLgXj363uKUAU
y2CMYmOtCkxB1LcwdGAzKg1++RIuYy9E0dOUU3AQDGvQgfllRJ4UDSgNTnkyigWe
VTkkpmrK7MNkF6OZgMUezOpFuNIx/lAuaAQ7Qb6FMK7bTu7Cant7QRG9XAZaLiA0
dlFdD9ZDbiz7xtJyKKx6LJfJK4Ty+HSppFgEgFI/UlJ5ljsl1MxeO12Hk9013J9h
SOEfAdR/RblJMO+azYL9tLxO2Leohk7NOqRcuAhlOqf+ICFkU6cvMYa//Vp4HHaI
R8zZhdpwlzIq6ZBtXNsByC+otucer3bvmQhzKJK/9iD6DQvsgr05w1HLQQslKhH3
3Kt3rHbLX3y4D7jQkhXGoAMbduoyl/dISp+MGpdZiV8xmcDKy/9lMk/wX+rCpPu7
he2eOsuza0tGJLLOZH33ZrQsfP33TGssHfFH1fPdOb2Cz7VXO0TNNxeXZwN6S0wq
vryPltsjdo5/KKrEfpvBcnoeTaFOuo6oGbMOLKrzvRk+uUOAjtGiB614nrmCYtfK
g2VITVcfJuJjylw0VUYrTV8Go6SbdE8BWolGNLHw27P5F99Io+80Ze/YR/XKunQW
o2yB7nkkvqDKxDrJvaDBLz4U4d+QuuZ1BT3YE7gt0CpthZ2mzQ08ZgvD5YpVZpXY
2wPKYVr8C8bdqIhrT8dALJE9d+/OgjFpmaSJ+6r+ngloEhISOWlycgYRn1Kmv1bm
fGQKmPXDj3e7bCmAGSSo3B12ji+vUQ66NpyeAb73QX3R2e/KtAAVIFzr8tBOG1Iv
rzb4HvlUG0BWDOdma3FwppJfFpAT9Jm7QqT6DjI9FjgCzI/vNyK+4t7V0li1b8Fb
uoKbtB/SkjENRX8heESr1jgQcwcN2Qwlp9G6/iFpfPeWH7mCXWgJE4h6vXQ4lg/c
Fl38psoCs9QwchoD+o3uWTUNpYXbiazvHCkIIKA+i+BvtOyKfNvydLUjIV4W9oUw
zqWUH+jtDu3NRJeiHXzJHiqqh8kiMIh25H7WpfX4q58PfTbjzEAHQHyoq+M7Nwb5
MAmTk6zPy/3BWqa6tQLoj3kOf8oEx4wiFvqywoBN98Aze6cPKoHbo8e2W6d/BTeF
txQTwWeDm9UvpqRSFRaaCOUUgv5xqRsWSNJylI7jBSvxrs2w6gpSZxJ7CltLrBJ0
6f9C7C4L6FKOdCDlymiHlHz3tVl7h2qOQmmXXLufunbw8Qt0Oy2ZJpr0SWiiMkYq
XiQWoTCHlo/AKoFYbnAloUmtupRu82FzGm89P/GQDs6i/I8aq1UgQoUlqCjx2Tbw
DpHlXKmc/cXxrGPCGmhxXu0xui5KsQQILj+CrW2IEjwaLxNLIpPPE9TUa4j/+511
Dp95HK7Wzmqu1S4NeVlYFMK6YJ5HBvKrBmMEfupUWL9pLzRW8bDgqJT0NiavpMow
8hYY+/E0VMcaFY4tgMWvj+JqH6Li3D+5dW86hSYC8UpMlLPS0H8V1g7iB0Gx176v
sOBznBcRS7thKRyq46u4ZrJyH4JjG3VeEp9aJRJ/svByVEiTm20FdtsshbcL4TtA
83lh2IrucQp6Zm9ApJh6kRGWYlzXYSwt7ZeYtr3Av/QDlYNBzv0T4+qfB0qMSCCL
Z5fLtP9ZiGKJzmfYuyJFYLsR6bQbvc9+fzhnbBCEU5nhHO6mOcvwbLPWry70BbJM
VCJ2jOMTWqpwYXGwoolXLLugFK9hPPlmuOijpMt9h3kXtSAJ7HpAp4grE/YLmIhu
M/mOQdA3e97tPxrP6SUs4bHz0fEzxX+18OPPl+4SbIhavSrom9UDLPvLdZoV+H8G
CpJDAlYzq21uK+/OgKRRVi8JvxaQvbG9UWF2qJwNy0Ujl8Ioe1Pp72700xY4z95t
msPKUjxyRMdHlqAHR6Vq3Tf/1lB8vVQnTXmgzWU1I0JpxOTyYYdUs9f2yqaxFf9C
ldyCq9e3i73HDD1CqADRTNM9eFc0YikzIWmdLbxVIAiQ0VhzgJwYhbIJ6JDrR85X
9TiqyPY5+sLtV4Av079mBbkuaXBvrH7ahjSXf2f7Psxk+OsMP3CB85tNh5LZzN7S
KyWmY/nUEOo/n6dF08akEZXWoUu2fdBV8KFAFGG7s7tp9sI5ZrdRlAaM4Xirk28E
Ks2DkkCxoFJidM9IRl9E5fjDCS4gCUQUyQYk71nWqlOfj30i83UE3G9+WWjNA0iz
r+IF/0pdXmISmpX9pDk9scS9fNE87tbVhUDJdDSS0ZDRCb9KAm6lvkDWu9WpNpDE
l6TuSCfeCjO/8MOktzOZSuaN0K1qVXNrDWu61V3pDO2KFM+dTGYGP/nDBpV4S8GX
wCgDU3cPaqJw1CEJKU3zM1jFDu5bK9HjWSxqOkfkWECh05rRJYfZKxL4gbBQkZdQ
cJ493nU2KO4XNloc8FELZdN4hk5x5H1g1SfI/5xZG43Dh2wbILNofszyeyvfJOm4
wj98E1iO1H+D31ISnsC8Eqqj+Tp3PFrVzQXGSK8t6oS59k+RJ2oHHTjzMm3h36/L
YX3LjFUI4amTBc7fsilPEZrDFf1nzledPDg2aKnHEEPtlfW3/0oWrtVYFT6Z35Ai
04pXcQR/xt1Ajhv5gUeJZdPCwtwQ1kos4WqQFqEUln3IDDAoGKU4DhsEcAI0dS3G
cWOUcNNk6RdjjhPUYpukEOGFlRsAckQ62410fXfr8FDe7cpKiPBV+qC8e+jikBae
ibY0iHYNKGuEzyBPkJWOK4rIhW+AOaKNNcUAu0C+GX6Pjj5pWdIKKg+cKLYgKK/E
CbVqn8zbB8nWtMk6VtR/+f6ZzUlWv5Zvg2pzcYI3b5lYT+Gnk8ARMqCSvF4SY18J
SFp3xOJxUdzuX9UsYIL/3yHDYhbnqJk6S033n7l4buVOFl0/TBBQdiYyjoYsTtE/
kzpUF3PrzJGcrAhkqcXFNQnxZB4vIeWcyLupJixrCs/mGr3LFPNUIUGfcQ4uT/zp
pYy2m6H8s4IwdZ5Qb/yEZZHl7NHX2IkdHoSd6F5hpTsJ7rSj1XUaHKD+ZiBabuY0
opLOjJninz/UWQJcCnXnrVf1sKL0uU2ZMEyHxGZRumPXRok+epSGswD3sV4D49xM
nn1GlqGPUQlxMDtkayEvf10kTCSUA5DgBYgunDKDu0qWADF07WiMwUaJcHav088S
ztPipEczFkWhhNhC/x8e6YpNpfEaOg76UjGgtmKsC8XY+Tj34eFDGdvxVHvunnyC
6UlDm7aZ8afKJSXBjj+dHT/XdSH2/c6Xiie7EfLYEa7f3LsJ+9ooo32kEfggE0Ft
XTuNvhgwPe4FK+xTjnwcYssDGLSUTFSKUKg08jnveoWgD68IoV10AvNP03xuyY+X
Uyghag+9jqXWuXRKVam9kmv6+FeStXpr/V+A/6y1xw0ZtCLy0v3gcqGro7HXcMYJ
FMlRCZUAsOlgmiLEXuMeSvWrA1bfghJshyYCmrJ+OBEqIBPz9RqrFvQqsIRs6Qp/
RUuH7veyIFPtfpPTbruk9s1/goULYDiNNh3QC8sjblV27WAsNtWJUhWHOqv5l3u8
OlyE70v6SAKIBsz4vNa5IhMV5+4GkYtykDfuL//UL/tq8vz8CmNRaw/NzGoOCosB
eJBdYTuvuNRLmtfvphNEIRbtPcNB6equx/1Qt70526i6ELKEpOS7a6hugz4QsY1x
U00g+g8zBcVu263+AGwiXX4tbxqyWR2sDvqwCJEvwVA//clDYqptxBN0nzWcf0/m
y/+E1t9147eXIQK3uSLslL83qvXGImWEjfGZgnUs2r3bNBu2kdeAZlJs+JqE0J2p
4VHr/ZubIhnPSBKVrE3OWQRuTjCUulmJqBBopubiNK7faHxmkgwGIsEQygsWbiQP
FaDC3bG6LDcQmgAgYdsvslvoM7zKVdDJxo+zMCYWm+V5b+9u1X4jLzp3+wJeBnB7
Zm2DwVYfrh+FEDbcO2/rmmw3gEOA5GWkOkA+gdYqGwf06di2zUY2XEwxsRVZVBH4
wKbYONsMUWr4jiL360sr5E+vX1mrkWDok6iQQR9xBWUEy2OFpi6soUgBiGhyUp38
JSTQM9iZzluoaI6TrdTa2F4l0M9oXWfJCTp0te/JOboOwxCaBqDp0E5ycCazRS9h
yFAwV5nSfm4xc4YQg5/NZyHtSXHqcGsK+jekRIGS4yuzncsj69/f+zQOvgbmzNQu
RjkuHEPwUEKXMBVN1yJgJKW3WNVJvY/ZU7HGTLsnGOjmlkpd8BRs9jhoig+mGnjh
GDjXvoR/UmIOQ49/SX70GbPvKATL6g6QPWgHJ0lI86HC8T+Umuo3kakieY5CJBxd
2YluSZ1QRE1VELEtCCfQ9fTT4HajGj04SufNYAv2h0QymKNR8Gs9yuy7Htt4kS7c
9M11ST427gRyZdPYjaicW1a4YrxWlICQZw0emQhBTCgxvX+9vW3FJzypXon6h89A
LDd2wyZG4211IQ6Y1n0UjlVkjvnrP0rjb8O5fPHYi8RzvKHwSaHMWELEf2XFlZFi
PuevW0U47BfxkWlEaFmwKZBOXekFxiW2sp2mly5mYdt9EudO8fC9EnB3fOgAR6Ve
DU/bmPxwE2IPUqklniGl4iEwtQtZ+NIP+2B57mWJG/2CuiPmU/ElVReS5NOcbZ+9
UTPZDzamOWYa0LqXbjR1wJsZoRyBx0FxPQnEv6mvnA1oJrmuzzInYoijTDC9VujU
nUUZHxTZ+GywQsOJ1F0Jy4QDphOm4P1jWHfpZMHxZiY/BTVTm+Ghug1uJkAcugz+
GKq3oFFlwPByjCz7pZKS8PPdnM7U+QWu7SVJ+ltN0g9P1mJHCdGZCmCAckY0ESSP
LlWeC/ExKVH93DkjBenbI2/fJMaSgjXP4rGocN9enDd2MWmerN9HBz7JtnBiy5YB
JNANlm/9Zkt0kolZsxUIry3PHq1QU4hG1Zh9k8kkWWgEtL7UnVbrJ1jfxfdw7Qes
heN9iS8J3Ey6q33H0Uy2w7Q2L5Am5aqqMakUyHSo1KngcFbJZFr4vk86qMCb77x1
Il/qWnRkS58PYPlUoNunTXzr6ons1j9bQVu1soDRwWL6YsNI/uws/RzZx+qHnMho
8Dns2h3X3/fAONQ0q6V+BZSMz18SwsdveG0fks/2r8NX++3IMKEdj+U1OeKsM4xH
Uye9t4usvA8T7Gqpfoq+PIM1DtTMCKBkFgMYVcgH8GLhgd/wUfQAPJ39hGskIqcz
EyfLRuK4nEFkO/FCpjayubhjnF7f5lnD0pdtlvQjGzF7wNOyVSNZlOI9NRpqIFeF
co5RJWElEDbNFJY7aaH5Ry4JLKxl+Ps8r0ndYsCL15QhdFlZbxxXudYqSijTmyk9
Rq50R4dixD4v9DIx4hiijgaLW3b4mzIRa073RMfeBL64Ihgmz523WigAJNj60ngd
2D6opbkL5lxRXXgbVGh3Zi8DxOHSD9OafZbVCJv3UzAya/wZ8twTDJ/jbDKh8MCM
UPzYFsfd+jri/BuDqbTUB/zJlO4MnsGaznZHwXRiidIJoTqYT/3e4SsSM+UVXJ6C
lNxHC1DMG3YiCY5G3n8rLggrslhkTvbbX+B3Qpru3X9VP6+hDIKEDJbm15qFYrFy
jSeK9i1BhGf03wJfH9X+j6N9B0QnpmEnGbs7Tp4pl9HJfP0dA2UqUDZggI0NuIK5
eGlGpHFO1EXcJ8jQwfhn5bV6Swd0nQR5znAkh6E23cBRvibO1xgF+meSG95LmqS5
TOhobLNR1T/U5F34We7KNqIT3yhLx3iCbsE+lX1HSHk3FcGd5lsOwn2InCDOk7cy
E9Z7DrqHFogs1wo/FqtdPHClFMq2DmGobly6A20BRqnOj2kI3/hc7/fPEaMF8M0r
q5ze5/VD1jLoYAJfLRzKe6ACSNElynWsBzwc9KRssARxsNxBri+oXFPJzfvcZRJM
PIxZRMVJIOt3cWlSpjwdYMAeohD3sL7r5snh1jXT1PwolPCnp2ExUT2j2mc+VGB8
LaMWiGRHItQ0k60mRZoT1wtaNVKdiVNb/964G2pZuiwxbMmNrinLEV+7+gLahTNZ
7EQ675Upx6ceD5B37pwjK/uRTKlgRDni8EPJ11Ba/sJRbVuEckhh+MSMXbJhhXA6
6vqDK+3opmLdDQMXMiPhqgxbHahvJaK6A7J3QlgFw3a/kqyKdb8R/XoPi/TXh3pL
WQg11xq2WA0JdMkXy+v/f2cGBRGhHIb22ZxOM4n6u/BWwtIn3AjwXxCzigEwQ1cH
4joTfDWC6nYjl4m2a5ObU6EfJv1NoAGEEMPg+lHnkPK/dxG4oXZ7pWZYJK3iefIk
ULmhP376JT0+uVO+Gll9DNQSIdliRL6VcCR6QmhCaqL9Yhrq5ygQ59rq+yomaBhH
Fk5kBL74r71cm6rKArkfTo0j96h3Z3G2HU7BLKm1hiQVKogoiYguRWyZS6X2Q4Cc
H5OaKcn3sYAe+qld9jvbpOyZMK+1fCxys2KXFlvYFo7etgfvLbLnCjFwKz7bsR19
YqSMk+QxJo+Eng9RzbmTZBntlYe0YYG3lrr3hIhjpzzKErVxVqTUCxML2wHMeupN
BtAsvRHv8z1F7OY4ruxoDSnSpLM2Mne2CDdtcC1V/pEN0FFR+ulZeeNi2xZcGzXA
SI8RCZrvP+8KSsHHhnJGnHrumd8OUsiMTa1PYzd7T4uPmhLZPtevyOBo6oKjWXKK
mJe2LnaoSX7YcXWfZ3t/Wl+UnzXw182f67fayVFbpfmHCKBA3HTUdHu8yB/0r2mt
RkmhTiuUgtL761az3N82tTaF1L6VUpu1kzEnfrvo0Vc6mWIeSubRSGTdPWnDxVuE
L5ponSNOE/QwvJCRVem1IAS713e2rTzJDqCNEC5kEptWu++aUETB08o3B6Ul4A78
SMg+k1dVj8ahVNez6G7glcA832LaB+c8whviBhSVwSjDMX5/Ezu+dsT0+rs2FHe0
CGUfqTsou5fD2PogMG0XFeND+OpNB/JUnNzOzFlb91jfZe9xPHPOvjZyf9qQv08w
wR7St0YKB/qmKne1bo6XqLeLnjnTVjVy3iUpXGwiElVvNtDEp3FFy9cLuwwIPedr
FCA6d1HUCiaWFxuZONOO76Ue+wG4t7ZBvonZzacOJxsxPpnRiCOnWqWIMogWSEJv
tC13U/haDTPjve6fBeI6l5rDzGugosP04ibz/UE6yCSXgIMx4TADmoyCtUZEoHFs
w+F9AcYHr972L6GoIvoRrBFRa818dpA1YBnerMrEBarc9lpc1fpXMSEbev/bwcG+
v/v0FpXXYnx2XzK2yzn1PGeSlshyUV6imrQghOjFhNU271B2Q2ApjNkSqPyR1QHV
qV3ADn9IEEAzXVUJf1O0DX3GijANZHwo1qdU/ROvAwf5QTjr1tAtQXTQfu9jNxit
9zOtOq2r2FNEAnGEt0+eLTzErW3khRFnu75MTH1KPOHRaUWeVgEKb+mD53OYO25G
CK+Sbk2agfUK4EJLhwZZLy9V/GjBnJvLUWX3vCprpUbiyCB6Cgh0lQWCgaZm+EIj
Y/skLzsbvuGeckwskqEetA4TF7LVdPFaDiTa/AE3pMy7ouTFOLHZofCHSDKosVsQ
8va/v913bvNk0i10OGba3y2WYx0S04dP8I+hT9wY3lA9UKASmHYJQke20ua/DZXD
xqPEPNqRReTggSS8nT8wdQzzoJoYas3AEO7WXS2v72LyIooVArrjfe5njRkdBOe2
8BABRF1OeUZXGhChZQ04WryXmDCZaImO0KQqpOwvPNxKhkWCJTRJNPQ43RX5i1GE
zn0AhcwkKe/3xUM4TERC+dm9/KykXhItjY4Jh/rM8ywLdrkdk2rTTClS0qkNIrue
DY5yn24WgY0Tpp82jMZqK+I4fD0hLnD+wLtMMC5fVgT/QYWWre7dw9mVKGQh4gOl
EFlqHP24+aRxsxQO801xzbzvhdbaTra5vIcE1OtQ4/swNcUzMkE9xv3Y/upVllCT
Z+5ibJziZVG7VF/kdLfLu86w+0cS+ILjQvaYB3WG3nvorpmayp0CJNQh887D8KtX
Wf9zHMiHlaAWpEMcR1+eKPPFb+dUPrgOQGXgixYqw/Oq4RW/pgM1m/tKzlDzaJHs
HQX5TyxnqFLfB7Y5NsKkbuwr7MAL12+FelQDbGKiXlQw8CWkYex8oSRDJsxClYYj
rptFof/X9v+K4oSQ2d5a5aCW5kpFdBtEsYWcf2oNCSvzb7XFz+ANPBV+zUl5HVOs
TIgZ/XZKXITS+fXuyk5g+Ok/A0Qz/IIB6oVNIGJuzFi//bcPxRCtE2frL4/IscT1
+uM2AF6c2nH1Wb5kKezWCk3reHWHjme0xGU1qZ/yj6i58NJpL8YxI/gusFdJRd0O
t33KaLJYvzaazPWVmtfRqWXMQ7OENN+Cqz9TgKxUs6Sa7+ycHAr1UYYVq+L3wX1j
paBHI/qKVdihBy5FSkuhINoxEpJFYOjf+TFGpP8rSFalLb5Yp7toCvhrciEeZa2b
EQjxmI0CkEK0U38P5NvUnoIiS5xsmqqed7SwkBqP31VhwN3lAoWB9ZI7Npxs9mQC
JC2A/OhnEApVdAgO64hPlUu6AFSkc7wQKBO04Ge+rry4fPxCCcx8HoGB4hrNSqS3
QkzvFH/V3YMaZ/XSHBpqfmJMIbz2TI/fpaZ+jQL7zyFP3dpe5/FLFIhcKN9c6q0W
6HqmPz7cTna4NkeyRHRXRvJRJmPlLM/mGkESkKMB67GIoStIjdm4sZVmcxsd3j48
pVPt+4FGUmMR1BZCzC9TxPCZSNXINuOSYbu9F2FtoB8gi54/DtBgyrEEUSHZKsW+
mXHv/tK7TB/8ZBpai6bnjgBWXXqhoF0zMX6mhKzkV8NItewekp+PJYkP0WUkosJ2
TrniY/qF7F8mMffN34kY1GS1lWU9i1cmbYrKwLswMDzORxBcLAvR3QioLZpJqpRP
6yq6c8LNbmslSaRbF7DFgFQYcfNvFfZG1726F2Aj7liIPfEIAP6dUiBAN7Cfg6Z4
S2enUP5eWFQccg7cg4Cup0nXcuS5MmmWhGFmcHkIuy/1BjCjmvQUMXu33OlkHTZi
kP5SZqSc0T+J5K2w8sgU9DxjIZ+OBhQPhodtco+ORNF1Wo9m9/LPP7QxtLJNBiOI
MsD1k9Du9E5xyxoFTzmHj6m1vX6nkyhzkwa/nHzdPdxv/xdIyYiOpGajVYUjqcoY
LcjHULKn9mteRiksi0qnPc/DmttHhsDCiNrVaWTJTM9UZoFyyx5hD6shK4TFddLa
g3RPOFnMn0mMRp55D/IzgVK4J0vSpzCxzZ+bhLVpLImLVarO4uIxhzRTiREJmsHI
EuAkLCy1YfEkaZPHMcmcME+HuunABzT1XRbhzEy2sxdnLLMZ5j+WQAAZKj/fQ3kp
6WIPzHeLJuLV9nXzY+t70TuSR1eUN7P2WrzBXpTbbtS/bZAFLSoHGPCHw3a2D1hY
FdAm3Rqv2uRUBhEKe25FWmhzm/v58xwJeHE4SK7szIZ8v1l6Jlaz97W+NhWowvgw
oHLMZHzGWdgmNNeHVLv7aVjm+Aayn4hWC7JhMa5EfhIEP4obypvCSW5nMt2n3dOL
76xInKUsMyCFVzZfkCHW9IwOs4cDwa8uZq1dmDZOexymedTos+WAciVlQbXVFLkf
sxuuCurqNFjmvE0u5pFtSCdI4VV4gajQNkPaDws++V2XsueR8Sb/CP2sfGD608C2
/P1N9ZnRhpDKxCTQPYQrAnJbioX//eRsNg4cHD7qoQddOmBC6jKQfmpughG4MS7k
9ToJSxAZ9cYpZRLyt8oID6EYj0xFkSGtJEXEC1vb485FtuaYRtymJSFcAvKQeK2Q
/4LDt3OFkiQ5SkVJ6KWqPe0VLTxxah1R7QwsIidLKMRKgmYXWmJSV5oqwHmdeXyw
CgltPo3qjl4toe9QbdiJ2EHd+TQhPwDSvfZ6+SqTFTCBaSEP8QlMjXLyyQmC8W/v
3W3NMyUD408UoyWMM9p2CEYwUzitliRtD2nSdc7DfEZ34+TT7rUisnpNBZ/xYyy4
2aqVW9KhiOoQwHUiOzW8TQlY5/qdTXDL2IeR/akZaJ6tJnQu+eP9Cm4vWncYUy9p
cA+n/sb0xW7na3gyNEJnBNp818lOs0HL9BSTWODUaLrK81K5lv8Q+t0hYNZJdKFc
gLg4mCykoMupOZBcIIXumgemMVKGjfZRjyb22udUwYHlu0elDrX5mpxiL/RJYGTZ
QgBk3s+4L5ihG8rla9Me68YYIT5L19QnAqnwf+327kqxwP2otoWmkpM3mtlUGfee
Zg13zJJuNvEP8mrr6sDz0GRBiINvneubzdiZMVW3BzDwk0nGxooQg7k5rtFkVzor
V6unTZWxxRS4eEIWACdpGNUhIUcv5+0RPcf7QxWcK36BZHl/hjgk6ST9pEAXWV1E
zKk5IvTUn2+xrO0zM7RdvR0cNoFXQuuNgPPA2raq2L38K7/TQYR79d4KepoWntp8
Gp5Sd5dwkHvuqg/jQSVRWzMCqnIhLpw+VKsNjXjMCYZQopViR58dPNRKoioYNUgX
2wtdEu6Yb2YPhM3PLwX3ZuJDLxxNtLLrLzKkvG9tuQSlGmyeIp5365fsVIfwYjwq
Hor8HtRiOGt/VPAQb4uDJO0/Ez4KrAnSLw4tiXw2Fx+9mpfg7xN3MhDyP95Bmw+3
AQig2glLJasI6MdsESwnqULkuK0ls/xva2cMOHGnXRzl8EmPa3L7/wSuV4kYJl8A
vu4+6WIQLlmjEMY8zxLsMlT0fZzB94gPtfVqlRGoCWSL2Xjc9BXb3xse+Os2IwKY
AqN0CA5Hayr0I89K8+WciKpbqhWLVOoFW2qlYMvfX4qjD3sVfPEziKI4u8uk33sA
pGi26T6A+VVxnx3OddqqxkHYRhkUeMf/J47w+ZqEkcMvEOkZ2Jo3klVUahpJDzWj
jA8JCw+uoWzoFlgno9nHWR9wvXnuEDWuoXpHvmi30bXNiJ2fRvis7cUdl1NIuv27
qB4pBxEfuNHPWOP6+l0fZuqjfDGPgkX1VD+4fVxV7PIssXzzedoeQrQ1zumc50ST
wPkQ+n0sgcUDqvi8mbz1FpxKCTWc3V/UubcWmfDOw73VjUz5OZVtuj9ZhQxx2rnf
T6h5+G0zqSyGALZSdEyO83IXeaWQCf57pmzctYTgZCUN4mL9QhkgPt3JGufJps1J
931NXaQ9wt1DWICER7WRgrvolrio71TCLxu4euWRy45kgJ4HF6sb8ECI4BM/XYLd
dIcGCPffVSJmRpRiKxrYlg1Xek8y2k10OfB5ZMjoqIwQnwrmHC3gDYzuFhpzA7kH
UWPmP0tIeKkRr+CN/x4/Qq0DK3n8KgAejIPNDNyhSIqaIxP/KFE9GaF32xj3yxxh
Q893widtmtOPUrgu3FzaLg4d6P5UPmqxrELIjuvLjM3PPJwAKkajRI1j/hKo9OpF
L5bZN/p0IyfXkkteVv9h5rFGGoi0Wlu+V6no7DzpG6Yk/Qtz3JgTgGjedGDAbB+m
khgkJhc4yyccTkpraKts9MsWSJn98A0qli7RhobWmq2t/sk34/4uk9dZ+VIOv6mP
31hkau3rymnQrkYURFVPoRK9YCSdORpYvZhuk0U8j/WEJNiHi0eyYTCElOZ9BBPR
Jy4PLAY5x1i2ByRGjHOg+Iw0tncaIdbIl1M0VOv827gegvppRhYVnlXQnWxjpVe3
peIZoV4pc4KPkXxKMNDv9KwrLemWOCFtQjhYguIvkaJoIoCsnhhgQLKYHVRUNiS0
G891n9qOP9WRsG4+VdTbZfnxLxhMxUeqmyyJktRsXdPbbg9HScqSi25pU05TP1nL
lJkLbsunDVEBrep5W7XssImYX842pOypkPYcwxpLofhnSCGNFDYK3ke4e8fGl3WP
5AKyZ0FYbNgbarZ4FgGbhEmjVj2JOIpOyzasYgtY2/mHxOFs3KhAksH8qjYPRmmB
aLftDLqFlli1jhfYEvEIU7fQcPZlwcAyTEXWrnTArNZgxUAhAKagvxXY2geb3zlu
Mp6rbWilFs2KoiSQFT7ghBeutMbp0a3BXNsxjr+kyLVeDf7FOzC2mkLz6pLOSEFw
Ggrugc9KF/+vIlLsQQ9OFMzx3BMTt1p+eMCkXiefRram267Kve/ZUp54YUJyGr1s
hBize+hrb6vnDJvVLjJD9lSdxixtyW7khcBP29m+gaNkOsJqeqo1tGLdsDvPdPMA
V9tXq46SadFFSPEj2CPerfyoEnkhVShhVcaB5/T5Ap10J1eCajSw8U2u1nqazR13
Oxdv7W7dagrd0WF1vQIUhdwGWDWPupqsJkyq0d8KnVI35gyQYybprucfnd33c+er
0s6UJMKmtvYLvlfVNEl9iBSnW6io9zy6bZ74iGS0tPPQpGdMgoVC6xgeytzmLDF0
V7KrNW8HiNATjZybbViXQRW7UUP200vOEFOjXVM9bs2dq9RFQjgYqTLHrs8G/EOg
Hyo9kv4reIqK+X/ycC1CgFOF7fL9gJQDNalqPymhmTuloFZT9WCqksiJCEZwVk4p
gSKdqrhSUB/8NgKPTlCpQdeWi6mY/GNzduj6hwIQ64v4+CnAhA3/Rshppr7QdFtV
ikcTLGOiC4YvRtBZI3edCcuxWNsUEWtMUVsPsGcV8qWT3LYcQkW1j8lM2XXUT+FT
bJm/tu+vKSx5xN48w6KsHHiJDd5chOcazpq1aKz6HbQDaaVeKEqNRB+RiScjCmer
UrEiYloY/E8npTlnl232tk7mv1fhEPj/xinkkwm4Lvi8yqi+mnrMSQ7RMQwcjumX
vTGmafFfWUjQJZgnbBWKPqRqKnsOAcy1UxAXIVw8/Hkzr8sqwjnoib7NESgyfqM0
5n/rAvFASA7wK9kmx2sblTftdm9viQWgwXokybVY2PjQUkDVR1pdipXmyNQyKrqI
/oNjYTceG9cl+7hbJ/YDaI2rjaOYtdGInzl0vj1WbnK5TCH0+RgaOHOVEIMoL0zE
23ZQaKbHEj4zyyduMLQrNJkI02/qT7pAJnupMiB0dhOMSKcfsY3IonYLCrHkMEUZ
gdXD++5DLQHLQbmW3VSWZ5zIUkLXz7t0hXGEwh0C8TANnIXgm5y+3N2SQjpLq5Ia
6+GvFTGrnnC6pXOtwlNkdyBBg7YEQ0zzlyUfTYsh7AhR2ePuoLD7ozhw2ZwFUAyV
0ZckWczfxp+ARpMn9hja8FpvXMl/BZUynqKWFXuSZ+eyQQAl73pstCCuqHyhTaVy
kWVKbWPajfuB2kgobHT1pW2Fl3hfC0s6imEO8q6YADtoUDKu/qda5SM3owGgPCXI
jIUW9ntd8FxrrgrHoTnbkQJkrxKz44ftrcbY1PqyQpbBg0v2xri34dlAlIUmhGJu
poOf6OqSwxIhbxke4bS9p2pw/TnvhlPTb+N865zT74E9HiWngVSqs6PtUeLJCPLi
A2P0hEWmvXOyAW3gbzMN0xI4+/Avpe75LNY0vWirB1NrWx0x26HrkW0a2DAsoBRA
NJ+NL7MpVLWU1LxOXsoIi+ZNuCASr4jutHOC2P42FFeh6nF/ZzOEEga9j6kGM7BA
Mb3qpiPB7Fl75/SdkZIxHf63TwrpxQhe8u5KHlKdwsTwY5ESGKIDz49QhQA2g29H
4Dth7lWLIkfBtXz6NWTZ4oBm4HLgu6VANB6mNCaqehAxM/JsDbEae+WENAiOY4SU
ciUf3FsaPTWU4lzWUdnXS8MGYxn6pWkchPZG9bvl0YXl2FcB9CPvnTHoCHVC5N9O
8KXeKGU979tUe373MdL3KTcumxJNRY2yOhtZYt+P61M/eG8dwRmad55N6gH9YpWU
D4cSBHcydut7NRKIVvjYgehUsYg3zAtFWXe+Zyq3sV/8nRqtH9zM5S2jVWQXLctc
Ayy9+OSM6h6f5wB4/pmle22gpKKnmsnd3x1i4CDWRvs9HMb2dYR86A4Ad9l2cg6/
BgEOxytY2Q7z65OzrDMtCbW8iqQj2J95kcraEXo9gYQyusRllF6t+4xj5jIZRgVH
BzwUlUa8OTQXTiaCs/2wg7gzfF8OlcYel7sszOwQ+UmRN7yPgzBUM2PrFsAkuIi0
mxm59Q3CzVG6XZvlOUwnIxXlVCuJwhjnC7RwmeooQZRZ1Dj1iSII5kMK4qs3pK3X
qHZjpoUBK51LXb0mLnA8usy86dWUqAKX8GpeqQjw+q9jdJ4PRxYOFqCpI4n9Fas7
+BSaV0nllqThPURezfZtnAKmJZrhGCX5VKKRgM4GjJEnfKKfeT/RjsM2FGHciKxx
5RmJIqBQCRqpCgGYSbmWfT3YpKnJRo6YAEIn2RNo2nFIQYSSurwrGRKC6Ol0mY+i
DZ8p48tyq28SAP6ZiFW9UbIHTp4sVX3FckhSVgkfftCoAxiFly2jJWulLOtx4axZ
dgcof+zk8mMuj7tr5HiLjeOvFRmDENHEfiCVweFZG0UN2HzGmP7Dxw5LfH+Y1d7W
nQvt+kG0R8LY5yXpqIz8kdooxZlR5bkxB82+l74xA1Q0NFq2xXSSY3LN+WonjFm3
3mGC0EcpW+MHvktcBpkzCwywsh184JwumJW6TjxJARlp+d0k61fO7adg5ZrdwQ0G
0BJqIuDHqWBcgqY6oTd+E6DOiv6XOrBZljLNXjlrX9dj8tVZQ6Y57jxszpF/hdis
7tWPBTqtZkFc/2e9TNmZggKUPj3K0us8n9yrTlJT5cae1/C0bdQ6BklbWHFYnw9J
giUyIp76xuVvLrz/VqCw6s1vRjevECwTYByzmp6TqH2uhucyMZRwsndBetNAZU6o
uca+Cu6l2I6+HGKvSSQYhlQTOwAqNsy1iPIOxKakQeLyh1lumzCTe5QihqC5eIuE
puXE51Eu7wFnDStbsaeTEwSXtJAd2Dx7wh0WQWRTBeJ/Pjua05KF2+9Hmh26pfSK
BqHVtEj5aQefn3qHyOv4j0cs3cYRe45jPqCDu5ez0To7PfOHVMIihncd/zqNYy8e
OTJgSgStjCEZLn+JMrZSaDPsSsHuX+BII2O1SpQZKMKPL49CX3LLFsXalGvLZGwJ
98fys7D3yGRc4ON9EKuEQ1CHyExeQcq4KTnGqXaGOUrR/jRlhZYiYfISpXwuyAeT
2SSafoTG/jHZ6Gm9MbkYUF//ehFQqPHp/GbwDt6GLmwPxBR+QdAPY2r11JKJgPa7
ITw3moCievD7NYbyjQYgIRUx0eK3qtxSwMOdLhai/u2ohgqINmpAqRG7dlIej+Gb
2lMWcaaCYAp/xthsl7+fQY84ZA+r9Du9F5scPfTNDz6DXY20C4UNmMcJh/RnnN+1
25qULU8tr2BzQ0jzS6D8jwSbeaa/Q2EDJc9i47tSkqJ5GKRUG6ieAckKvk5umpEY
d3c+hK8lU5Ym5GvJ5u9hkdXEz/wNI6U9QmefAXaxZIJVg65sJ6K2DYPP+DvpYkl4
rxouItrizIdsNVkciTMK+kHBqkvgQ2ZByWPcSIHwQ9GU565muUe0szS3jegfJDv8
+/d6vjoOlYvWoaBiP8TAXlH1wwmn77G5z4p+u1shIWhQlpmBtNV5nsbDug0S/toT
5L9Xef+pZ0t0uCPPaBnhV84H779Xec+XRRTjJ+ov84Fkprco+wIUjWyJ3J9kxByV
FCISuYpgnzML5VZ51QNxOuUgvW52PJO2SsiHMzrUop1oupMxBktE2MsEJfDKVlQT
W7nVmj3s867EcWG0fAePbQ6H00mQIbpqPRVMfumBnEuO1rD+Od4IHeTTcFtqHrdc
zW6IddEdrBspGhiVB5lIQROjAgoFLANyGvZnVEaZ7tBacNm7MmKwgOFd0t7CsVHA
cvJSn+sz7wKC33Iccfg28bwimEtmPtoNIpjahkehZt6pHPMPXfPHY6Psjw9z/Q00
1zZIV9SUTz6sTZLsdDdYpGelOBpfR6Ooei99Ba3gMfAuzUYhsxgLE6petwi2B+70
/71u/bVJBJ/JAco8cfnV2MIN9MzBxeGi+kePzkApjbzOTOHrxU4UPchA7QKkhZ8c
ZgJgLV0mu6In1gCyd+X5pkyN7CRUI+TcmnppifcBrsxWpU6uiIa9n759f+pbCHww
6LtvIEeOWGlO+mHWoYhauw81Of4xzYDPGEPgYjQiEL4FZm7CkDC0CbFPHlNTg/B4
AWNMH0hrlR/ROowF3WV32eMIyEluq+SqRM+Ix2mT3e3cOU/9b9z+JnC4d7AGFE6t
TDAQUpA/ukyj6iicH03Ab/AbaAFEMpuVOGfpwsWPVgF1kVPL1FLSrNud3qUeZj1n
PnUW0nnIvFyGH4KU62JsKfhQwbScu3lTCXQkkd9Nd/4je8FD1F1R4lxKtMlQDs5n
i7c8GIrRkd73Iv5F29t2WMHF7l9EiVE1X7T6lmtStizl0+WBGGBlyNWNGtheZqO6
GNH2uPqeZ7vZAz2Msg53HbV+W05MsIdGm63lz61iCYwAmPW4RlpNIUbXf9BIz/w1
v0Gk4qni9qbG2tjt9c7xD/+ZlWh464GP+0fBxJi+ziSYyq6e+XcYqsmycEyh7g3E
SXNtO0iW6zVgC1qyntiinuJvIay6cvhNZABhe+ZaMo4Dq+sDi5AGQ15EOtHvctI6
yjntBWgfmROHqeYjbpZTVrdkguQjQrrhfAhJ2QoM+1hUOOlUB2JChp3dyEYufsxt
8+X09BdcEhb1v4Nbo9slicp/qQnQUPmasD69IM34UT2y3WaFBQovUqoc1mD4eHQ7
2qQY/puWN2l2ntUEZJSv4jbg9HYllACUspj6JxjQmcEm+e2vJ6tmK3Es/FavgigW
T7E4BYoX2g6x+UwjEjlg9acct+1chaR6OgSlm4gZc+TzCuyjt/AmHECYsOzLaYkr
DZVfJ48lAG28ocAmvS0/UP5mEQ21XwUK+EUnv/gZ1HL4cs51fiIM//bOnJXNo3XS
j1tvzI0cWBnJQGPwXje68BYXtTwOYhY/T0qvD0koX6LqxEXuccTxBxVyF126kkO4
p/WFYSxaLC+wvDF8ponzsarVk+rtrc47ji/OOIe/DGbypjpDS7MNS9uZNHKKxMwy
vMQGYCK7luvwOyCk0OW73lJ6h5Nh8ZqoAV9ZTewFGe0a81dA3OLv7aW4V+1lJMa2
wiVaVgmHvGn4pc7ZQ6nq0j25At1DvG/SriD2NBEVGKS3cX+hkq9zqwsLYiPrg6PC
Yhp4aSjX9ZBi7g5g3HKMybToJY0qGtPRHT6dCIkG3aS9ClnLWGhrnaGEKQXISGIb
cbNw1Me6mmeN/4ZbwGe2FgDe5zb7A7A6+oaMwN/EOZ9UU/hUB9XLKRtLkQUMEbmc
wF7wV2UFDuXbWIjZOxeCGAaAVsNXRILWkMRo4zeWD6QDHNPMIMcu/rCagbkapoUR
rEYQdTd59XSZvK6j6GXFJZ7iJqHHW2Ux6H+qCaW626slI64wsNuamhD5AexMj2kR
n0zKi90qz4oxfZXZzmzfpxqIoWzKb0JAuZ6xtNiIdGMYx23wWXf5VYfaHKHfF/We
8H5ZLlgJ8Rlw0jJM0o91qTfeF44Ffk2mHt0OiXjdpT6Hfl3Qd2Is0rhrFFV6/WC/
tPSZXt3BBhEWuo5Z4/ag5Od3NoyQpHt4xHdhtOjR5qtZ47tKYllTJtsDOGHKJQ9f
CIK5/Ian8olVNcRUaa2MhcKj4wi+Jo1F/IPW1pclMDheLz8YDuW3R+MVZKAaV7gq
2JwnRtwSZaXsRCzMcRE7mbywSe+aOi67Ze9sxmZ9u5uODw1Lo9XxSFDtqmsYGyDe
1pbEvMoMZOZ2c/2N1SPcyDZybBw+rwyOXBCRpvjkGb9Qcp9eKzWXrQTnZp2dS8TL
nUhR2EHjSHjzSTciwSPUTM90emqwQXGfkEUiJ0wwxVuhkVW1ZwfVtYyd2maqVcxE
kYkQkwZgJF3MzpgPnYlN0yvnhXRwkigQC1q8yh2x5/ZibJ9BgJv36mbNvpoLjsKB
jBmItf72nyg3aoY37IHn3cRCEHdT9plFCUnluMqt98Aq/+pOpY9VUQI9YXi5iXW/
ehOE8GAJ4mfEnIFiRna9XDXs0V5jPWVh3+cmZvnse2pwkbDpeAIGTa3cAkxWkzxH
4F4kzCHZOKxHLcullthQuexHIdg6doGpfeEPckHt2XiXhOmNXeWFKMfvGi8oi58L
U/v6iLKPeg/tCCmeUDqbqXslXfVdCxke3t6lR+Z7HYIKLvwcTkUHfGAnPcK0Fobt
YCwFMETtasrGT2gGXvKAbLC0+M84e2G14JA4ypmYigFfNM7oo+1wR+WmiMOfr8mG
TtD3j2xa8GRYWQ+VPFnoFNkddvN9YopzZe1Mta9y717AbIvG4GTg68zC2Cc73t0x
DM+GXygYZsy9oWbjSEH6W2TWaVUdoxPywfeEX2dWTz8C4/p8VY5dzkTOucl6fIl2
a/vKC9JLM7vbiGSeaMEnQqMBpLKIZInuhSAF627/eO4Z11YS9VTyOXYIJ1bnb0xy
mYFhxsM06YDVW/CsQDEx/p8/HbsUZTGjejeUXHE01qG3eqwDGlIGpwWIj2Bwq2hY
KkFH8Tm166WcpkBSpoWPfARPP3Az+KtoHybjUl105sCth3GR7MQF5o/rLsS8abKZ
/4I/YOWbud+XQkKlqdJNntcxXD3CTGMmsLAg4/un6mMQBmKHkIbtZNaPSQxGhwQO
OQpTHfsZpZs/E1q1ZkD/HdwAFxyFLXdWpLYZIlI+txobJGJ5sYXMbUUYr4KZ92As
q61z8rLLw8jIz7vw5KQ5eeKRNqC3p9z2TLmhWVrwtWxzdWNmsy9/o4S9iy+Co5zz
9/jvmWwUmM+bEllS06Jn6P3kbc/sLu/D5GziXZQaTQ0qrukIRIIN0aFIqE5/5Pyo
OW06sxxSXfuV75lCYZU0dH0Af6S0dXOy7ei4nkDxXqllNJtieu3ngdYtd+I2VMXD
b8HFgsVJM+lBcrvGdtycnuU96sqWcY6r2ru/TuT/VGw/ok2e/UPVI9/66ndH81Bj
xWK9zlpWVCP6QccwZ+1qRQWQDVtiGATsV7xcZ4dcawtHzvgRZIwXPcRWOvTsgW4i
K5Q7hRTZk51cPPgvPqq8MUBEb0C9jHuEBbs0YDblkiZfba48kpfbZ8d8THNead9q
oahlpFSRHqO7WPvJu65X1qmPFH6n+p5AG7YFVjZ91U2jxcvTaV7GCZY51KW6YoH6
i+nOf7z1frkFVMmWy1gNgbqZfzZxsupenksLUmcLjBirfWy/rO+H/c/J9Ym/Kz8I
1x5FgeArvKh/x9GIK6sjZKAH3Vu4PygDQmtY6tPG+DLMwNa7c1S6CjqPRwfM1J/I
oDpiTEAtLua9+bBWbXMHdBuRH2zQ/JDpmMIu0vbERr6Rij7cFyR0aypuDPASQNV4
VsHilnSBbHWldq07YKlkSNeP+q5IOjOGIo7dGjDgfPkHMEsecBeI6W9LFozbES/N
2gx1TchFoJqPMPQiziTMshnzH+RPMjcIlj+nyF8mwQS2ro0nAF5Cbqx0PPI7M9Qg
5gcTFiAYVlM29vLV4UxhV8neafiF/hcqr4WfqmjM5AG1MnELiKjv8zoiaA3TCBGt
deX+lHMqHxtgihAbi2jYCHsLnqZvkKf0MHL9LYruzl9+6jgYEoPJwVYjirvIMuG6
GaUPn4z4EuYwrbafcDC6u09dNrsMfL3T7o1JpgmXRUpY/1imOZ4ljphSAc75w7Ej
eyV1/FDEvEHPD3nelRzZ/k8ayH2Lju7Qjq98DQ7oqPxMaQ7pAs9mmF4i+d2mCjNe
2QU9fTEa2ycGL2Uq3Dy4YoP6dPMkcnBL0v4KkwlYoWb7EyZkk4MFMsJJmiDFzPCO
gbsfvZSjEpzVhanUL/OrlER6V4KlVVX85bc/cJD9kPKEacBr6phJPdgluY5p3XNz
0DQFF8EdRJkbCDNkmHRfSLKNt0A1ydRyGjytrTB5vcjlsF6b3X0Z2T1NjJhmuztw
ryC4Pk3t3OtzlIRn96Ic1ZYVG1dMLemc6FspwRH5rxlhtTtrMn7EuFAg2mV0TN3t
5m/rnucRrB3Q965lS/q3xrAs7nHdBGCVrkGN8j+vulyW7u6Le4XdguyA81Z8xS9M
Dd1lvs0mUukSUww9W1F93oTNvFtEdgNyRRSxIduBrQwzGcEaLn7RYH9fAa2Sr5Tr
DtaFJ1QJGUhekLnHeCvXYr/8LNC6ruyTWUKk/EnmnENTL8T7724vNbGVDL0j2fGJ
RjgUd6xq1Yqa6JeKZPoPipXSC2hee8EBrIB5qfUYdC+4GFCJIAq6OT7dyZbVHKA/
Hb3k8DnxJMB3mzehtlqn1T90aOQTuuoZfIrscsqlRydi9qWyOizg1SgdGFgkbyO9
ianaRMum76BHsqVU4LLTVgcYxyJrVdfSzMr7rdTZhs9YhrxKVDEOSKsw2kqMwy8s
gWltPFA9QWLzGvxdH8OFNqBlcUb3BHyRHV39FK+kV8V+c1mIBZABxJ7Hmfp7an6M
KnI03E0TicO+XUlWmeXr8S4/Go3fjdzooeSLzhg3dPI8cV80ZEQ4oJwaUPgOex6u
7RChyOQn81SeboAEf3rCjROiC+fvauae5LknvnAuUiCWKF+jMbo/K1K5sFwVndnY
4sup8DpVf+gVeIAMPGvIopZPpK09zYiCX8rjKtsFexxLbrtYCMZ2oVeMi3SR/fJX
tsVPGzVaH7U2TCH7Kgl5SYDduCF6B/bVPRsw3gpqwWTbauCvSc4cquaTEL5VoGHG
5KQSvO7PO1lhieNYoOSHGSAC6OH89pjkTeHJqnghg5r5iZ43YXq7Ncq9HSnbwp94
mK7q5zWiHEDowNIfapYuIM+/Tc5Z8pk29CK/bH0vo5bbXhf5Evfpzi/zUcOIH8Yx
Qx5+2h8iP3Jy2r2eKeY1rhwDVoUmVVLmCaYlB0xoW+S/YLvApGmr0LqKwEqxI+GY
jIrBcob+IPN0I74Iz/afoKKoTmgN+Y4n35mvE/JKwtGyEWYuyiWrMPpDtUWYYocB
nfP2U+wy5041IgBSSWL8KWYUzy2PYNpTYb0cOJ1zrpBdv/tvJIZpaftlLuafm8Lq
IwPbflxpCE914P9VlNYtuZC7MHHEpK3WYEwURcE4FZ1bzfLZkoHuL3lNWS84uxDL
1ag0h9p+O2LOndmY/hyGcKfPlLxochr+du/G1nQAVlYBDxQFXauKbgzl9F72didu
Py8ARnGQ0H8U/QYyWzBrQItW0lvbbtBfMnMBI0BGczgj/BDggZbuNBtVGoWQWNW8
QnpirJ5FvMWo0VpPasuqtLEANgLjTZW65fN78XklvosuuyQIKA0yiVGNBWcroVQz
NgdJ3y3GveRt/A0Sou6HlWBG/U2avPumQVhoG9WhWdjRo1Y1saEDxwxO6Mw3eToS
D8SwLQXqKtLA53+AWdtzGiFTftKKYIGBzoAV6qwto3fI+yJWu0cuvVJA8ze5fcmW
6BZGRd1FiN+qfN1EtzVVeCm7i3IQYhhx2P04qBSOtcd3xabXTYmrBitsyDE925yV
M/H1qIy1DRuDA4nSraiwF9XQ7tRvDysyfHdHsWWsK8JZd8pqNXuqBB7YxDgtWHcU
MeR6EJK/7e8Krfgtp5jA2S9fkHtzT1pYhnBPphdKsmmgkWYEd8r/10uO13OLK7Dc
+2yxJc5MMQZzfQo0U5HU9gmT+T2peo8ZKNkI1K6jl5kWi9ZIlj7bp+5sF9Tf96pZ
Z0cw0dcwcs8RVOZdnehcDfzZsQYYqUVUKqolablicKuTKmoj9FP7wboldsK4g8Dt
jzUU3g/VyjMEi+MQNX9gkiQC2Asf4jcvutLqL++WQqqiiyqCgNDeJ+cPQAgdgK5X
HEe6eNFUqxdm7z1yEsb0/BhS32q2wAvQyptiOWtn0TxEvkJwsqsey9a/0DcR6iQ0
ZmaDEiHtDow8NeAFseZvXbN6n3HyiNo5uRu5xo8QQspqM3iIKYc8w7Gwz4kA/UhE
lma6WkFzUSVLElHr0EmS832neRsZrNxSiQ/dVeBcqgcikkp5Qza/T3Flb2onggjq
kGDkJsgHNCG8cSN20Qv6Fi59XGeBi1HyR18KCQ1ZrM43/toFAFuz+MiAw923VxaX
ClC/sElkeSEE0g0+AGCJe5gxhHofVmfTqN29hhCwZ1WpkKv14PkKGOtr5ZlOoFez
O7FULeL5GO+0XXTWd4BMnxDSKQWQleGZ3zjldZo8mKYe+nIaVwtYK0Z48sCCkgXZ
OGJw+eTwD+TLhS63SGgOAUN4lNNOUuK9+zLmWyq/mzB5uTb1BboF6EKwTUmvkNbN
Bld9wmf9kTwDzzPRut4K8Av6dMdxoacXPzWmKV0Pt5/HkcIldV48wabKC126Qq1V
NGruBLfvi36QuwsBdEU556fbwowTGmJDzZB7MHSKrZy1gbDY2Uf/0n51lF7ThYB1
2tWIWzFvd6h7r77ZdYYZMw7AORkzGErBo02Vk01yb0mnPtPh+UxM8679Jj3PEP6w
bEhu0gNj775+8M+b6QrCazG09TqMa8LEmt+9uJn2hVwwzkSEDjZ9nmbP9nYkxkxp
HsjRE5Q/5EvGOyaH44awKmx0x/ooMbQDUUyc6sTVex9ORWU8r/CD9O9/bCcgTHnG
/cla3TrVO5X3wkTz/S4OY6fjKWaxDOxiOuLXFRm27nv4SFPOD9FnkfGvrJQPtzKU
Luj8XmqQ1fnHjas8zP9Zq4vpM1kWj25HO77lF2CZ0My1Hl2pyjiHDNrVDDi3nWxM
pTrQlIkbzylJ6NwQhnx92Y6RvlLpHN4einoH8CX7jokEtzQolYkydhay3+J35Z4q
YA/i0GajLy4/o6oH+aHNT0NI+r8H6f8EEeKD5D0AI1u4QHsVlKqOPGQLPv51saNh
i/F/DUqiDmEfQwEGpuFimEGG+HPvsArxCSyR+FMs8bML8zksjtNcY/SAF3wD+N0x
R1ly3SLIRWQo9Pk1wBbj+YVQRLDra1I96uEio1c5tguG9Djc7IkZnrXYNBJraUxd
ysXobCwFNiLaXr37lABT+Cz9WDlaF8DxiOUnuczZVQM9IydkKCp8yCx5u8NzH2En
O9hFKgHWElGjln1nlJwSIhkEUh9dxXU1HuzvARxiVZCxnrll2iT4th4cN7z4Hm8+
bB7Mb1OPSjClEjjgzrogNXFqwCR9wvU1wB4+k8/2smQmIx/01SqQkiHB6dqiZTLS
W8qbROSHp+dwkwUKpe4UE19qVa40xqu9T7F5f/o7dNcF7Z6NFdfT/9sOMnnqi2OR
g3+YXlkW8f6XYjfvOnhSfVG+7RANP1TZP9yVb0m7paCjfMZthWL0xruxbBbNV6dI
6Ll5DzrTI1jloAhg20Yzqc6SympWz3LbRDOvvAKozJG/mzJiKNHs8aAK9cxF33xo
k2gXMVJl3Q/ET2m4n/hkBTGYKH6WROAXCWznnHzHH+mKxAkyrbLdHzEkMUUVzUVw
RbcrYU5l1w1RLXIfUK2jp8mk1a2dvl5Gk9UkL2EIq6itlaBno2fBUuUnDfAaTNsF
nqgOSSNVNtncu0UUBLyMFguoyBkylqcZHPMFNRhhn0l7RrRBvwciNSE928tvsNrv
wiSofq5foDa4v+E4QmPqw1Jx/dAnlnlSrnvLtfykjMblhdVYnfwZEPrFWzejTzxI
Zo9JHTXu+flcwzz/Erz11i/w1kR7CzAmEmZt6ovOE7hnKEuwgT/dmdi2H+iexUCj
oC6PHQBCw13MQwD8llPp+ifq3G++wgdVGD72rStf3OVwoRtVKMizLC79oj59Ov3z
XomjLhdX5XSSHk5QdYxo1wch3bKtA8tgd+Rn89DmrTVg9ozsPEk8APBc/sbDq4S4
nzRdjjg8eSsbKZbRvX4hwuCixdCHcAnlSYzJ+p/S0A4w54FBUScljg2VWtfC9Db7
FjwuoR3XxuTbA+NpKnsFXb2aioY0rZJFplpd8Ag5o1pk4psrTV30wftnBJkw47/J
QFiwdzXCapinN2zaS20TYzEBbUflw5stKuMHkmpOqT6MNe/Ih5bR0RMHmNwl0uXe
DrmfHvs/PsFE7zp8GxKPlVEvDzkNqNyXPa4wZtvMgUT+xcq3z6fQlv3B7VRi1T18
f0sWUoFGXretnrrbA0zILkJjAldukdIp9wnyPIIWybkLsiR9Ud4CzvAcjjvh4Fud
n8JO9sS22r/n/otNLfpAPx50gP1IKBp1T7+ia8QcViGEC0yLU6FLwExZi2EjCZtr
lDGG5SFxOWH+xG4lyu50aa67obfDNPvnQhM182kKJ5oHh9DFXIMFOmYy+MOkGk19
nQ9M1OVYJ8ezylcy7JvPftX0AwLSEq1OQN1EQuygDlfvhIJuxDH+oHH5KHYtOUR/
2zimFgyRg0rgkfedQRhK5W7/pyFoiT9ugAeK10JqrXxzfsgrEa4YQqiaZt+ywJhw
GKNwJLsAt6I5uUTcJy0TUEy2WXzbbiyRZZ8G/C8LTdPhQdd9wg3N1cU/BrgTRnoC
AkqdxRLROoqYgDBjXXFF/ytzySqcZhkqqr6h68H2hVvSEPSWPhynHQWPczsU4BWu
p8l8bnP6Dn/7LvSSnnWiTGB4g2QWTsquREiNc3IRg1jZsno7p0ABHYxZ9TSeokOE
IjWFgy6hMqOntS09PkSiCZJeIpgY8QrmU1F+A43lAhLJPcyY1Uk+Y1h6SvNIJvRg
/Hen0xSnyzA4wWL5Y+NG3ngyf7PfuWbPNMSKIlZMlayY/4fA0x9QYsmzT2WOU/TX
zOhUXb2zJlhZDCX8uW3pOgD51RuRiXRe5jSrQGlM/ZrlTh7LdwaNvHJ6xB19x8U8
/2TXQQeU/BD12l58T8/+zFFYtMJtC3plJDXQjVHTrYtTBH0bbEKKNo2E1zTnINlP
niIzzNWTZpHiLsY/RSey2KTC09D8zRTP7pTiEzKDWRLUu0e+Wyhro9pRZBB+wIlo
dPJGWBHLQj1xOAW4vjPohM+ZgkPhLmrMkAV7vrOZbDkkYS0GOrp6KF37+bDMlzcD
zRgBAwTa1aJj30KybZuWBIj78jtb5OhmyoURF4KK4Cf81WYB0PkNgTn2sRJPgt88
kKt2oqBd7HKYaZGgX6S0bsazTjLzLxi2/JRCZcZ6IOIsTFUjnhTCBWtnKPBEYZ2k
GtI1uklQchOQ4o/IcnV0FqRSaHHkAgjwch58Y1ONQKUlMVKXU9dDb1iUC8cudpgc
UNbRRrhgAMt2nYWm0KH4b3oHOxngx0uzexvp0JPtGO2XoGLU5BQkZMycwxIr67yc
xHQjRjA00ewsPj5xKNsqA4b0kYJeropAt9Hugjex0hrfVW0Bvr8wVb2Ln7HOp8kO
ZnoXzVUKH9ACaf/42NzWjDLQwwdeEuFIs6Vb3seI5u8tkRoP+UEZPrCbOAlpf+ic
zt3p7cZX6EfSLRlMP89xLzXrF/tNZaWgZJL49K9m36HnWe8Rebt0d93ViUQqzpnE
cipiAmxInJoyJny/d0apoOw+ykIOm7aTwIDctVLt1L0zhcfQxTifFGipgTJxEOwT
ozAdlMh0xRn6TVGam6RJ5EEhXcS5MGtxwadijZHm4xD2InrY2Vyw4UkYCaYubgrD
oZ0ql+pw9LgMD4owNEAbMym2KKvnSvmK3pzpMzX/DpB7pqMM1bzw2ASgUnRI9bEk
vWAyxNFmr0oVupNtTp1Hv7B9wfRatr6g8JlkAt9XzZbyALJKbXRqDTTC7BvLuIu5
Whi8l+kvxap5xIVxB1RgT8jiYMQUFfc2nl3ELyDn2H5MlaDnA8z0iy8UjiQd2QmF
YRZCa98WEKuuMAqu3bup/dn5OuvKfK5/QFY1EWGwlcIY340KPZmaHi5PiHVLuWp+
oAaYRyeN3QK/QcnIN9b8c5sMUc5BO4wpOiEm9BEKICyRBbz2QbxRCDYhUT5t/23b
YhPZKTwTeBrVZrBUHR66/8Sp1DBzRQ+/5gmiOOWhdZVOGe9vpeMMU1n7jPfoTnl1
VQF2t93G2y1B1D8OSUKoUAqjpMkdK0BuFDb6ox80JlKNm3pAw7vu96mpi6eyzWkb
cKbTTG7hTiMpw8nvSu4BpyjdZpTOcdL+mQzb/4ofgztLRLcMxnAgRlzq3PgdBaj8
usMPmf0oFM/AQx/++2mrUs4LI0551O4LPFj8Ca/otOTP6CEenDtfa4yDs724/IM5
LCIWxgR3xg2cFOeoq1GnvNKVnByvvsNG4tfU5vNZID7ojAYfjomPb0CWcQpUkNKU
ZNaIlR0Eggnjwnd84fkh9LEGKzYhj/ATDxcVR4N4D0qmCx8mhHKZM+df0An89F3l
Hejw9iOSi92/CEWZHrG4N5+mBMBphNcmQPDR+U13TL/LOYpjTp1zX40IVk+RCvrV
Ht4YUjnOiQSA7ZviwwIbvo8MSYIw1qgFTeO/nnyLbvU66FE4nY4PkpBGfiElqUi+
iwV98zgMUdY0z81/TjqDjZhlrKInI2nzc9OdOi9XlIJ1I++TIzsSp0pLNsjq33/D
kNpr8w+K1HpBjnPdVqoEVDVrLl6yYWz2VvcOPPxIF09XR49LX6yZ8XcKcL1W2k6a
MSALIhCj38q/a8lXKpfUdiVx0QoU2w/Ic4bFs/xFdwCkuRpIY4gL0HHylu9rr+6/
8qGxhQroLg64vNlADq2ckysQclj1+wod9pBsyfGD++7a3TPwBsSIjhT6pM5fwQs/
DtkYkSU26K9f40gz+36UHgkktFWxxL8FtZ7dUZO7Gib1TGnG2QHu+vwkTbvSmtZC
j4dgGfeJLPyZY1qQtAZoSRLAxuifJAVEcBSNXcHgE7kRgBXf3FFdH+Ef0+NGOve7
Mbf1UNxBfW1TRG1dH0SDrgIJOCGeGZh/faqV/TIUPcbaXcW6dkOGrCkr5hDzvF0k
UJommgjVpZeWIhzWLQi/PavemZzYOUGLuYFok85yv3YvnFgCxSmTKKXXWgKJLKPv
gadINfV2P0PZZBo2Bs737U6ZK+Va+R9ODcMdizntHTY38WGsla79+FDgK5fM2Cgz
I6+Gz7IrxpZitbvaYDHu2hdeABmPgiKuVqeVb34C2rSXtUiyURSRid8WYdTU/OzV
oz8cgyuI/svvoqDH/GqDZMUd420hyMf0Z6NdkxwaFkYsHjK5UJhEaiPW9aOZBDmA
KdJu8RFDlZKjUF93fvk2ZSnWMdUCVxOACsUTBbffukqg6K0GMIoo3sP5WjJzRDIy
mvxGb4btV3Gk/Ep+nMg9Ekq4MRH9vYOlcAVHzrPHOOA50YR2t8jcpL1kkspp4rMn
ckut+UNKn42T7g7ob30MXVo4IKgT0M+L2xSUqh1xg2OiuspynzFSy0IqgSCwtMG/
bBfmH/LPzZnX5I0BUMK73APj/IObYWVasN8Er2yyVHWKkhFgP/u1xo9sj/Loii+x
TfZpI1XqhPhliSkFGAuuWp0vCAdTW49QSHqrmHM1857UFW11TBq1YRc1P+I/R90O
Qw9r/iq9jZV7xPasVuAShYLiQjuwC5av9PCGhDqN50fMo4z623aXmwgcjt9hmnRK
ogvGibstNUOTaAmxEnPZLKpKCslr10l1Xyv5YfhpMpKYu5ikehMHOwaH9WJCRogL
H3/lFDnoPRcGENLOkoFeB2M1u2cJarPUgUkZpLvTpzZVIUhGc6tYko/eRhfPKKWD
KoCHrFh20hkWHLVFQE/5g6nuqPSmDislf7H8ldguAoTUc7DlE/d6obch/1T5Jamt
22YF9sLDpffmV4PiwsG2R0S9h1OD5hmBNM15nMq/ErMekCsl5F8X9zaIK/DSjBJw
1c5EBt14G/OKizIcyQYtwr0TrNXxYzTzGiezS9GiIYttJeeCLu30XYDzwYLbf+gj
AdVbm40OYzaId9RKUe8c60Wd7wh/MsfwR7Jmf+W2P4bepj127HeSSeoLe4SgzeMx
e5IgnJ7pDwWBhvg6a9Bi1nk3dJqvlkUCL2kTgqgN+zw6xEsR5f3tOz7Zntynh57n
t895xLYLV4NaYTZd7XrjEyiFuYR6ZJs0va8eGtoCryrgQHbJZjDejRlCkAyxOXOf
zkFbFXGSa4Zyo/ZYi+ar+1LQ7s8DQYNai2VKEK9VB/BIOEdOQadNMzp1+hipHonS
qbtqBmzWYLyyqbZOt1SkBWXlOGhJkG9GTP6DrqpPioR1EQqI6CpbkZJFXCy15qGj
Nnmgze8LBVDCozMrSfCtZZ5lwPMxSjwLgAMe9BLEg63CqLmXTzRkC6q2aS+9+V6Z
GdbndBLDzansVYE8kH3jYLXtt5WXCqntVE9GrkSUvbhVBI6CTI6RYBlyn0jOE2nh
PjnN+01qsok9OnfUe7wzCRd1gdK5JJo8HNyose1OgouJvSZHHKmTp3obUtySkRb/
hvEaEi5+PiQkBVAQ91yNGmrXMUIh/zmuc/fhxIdxtGlPLJQG54UUVV6Ix6svyTsO
D09tSWKPr/2CpI6F6VUbnoMaQj/ypya74fgpAmEvgV57nJv/JpiFFuEs3nJAUtMg
11c35kANcDgBQN2KNMWO38bzNg9/Vl+X7k1H76wnwj7W/KQ3goi/32LrRzkXbSab
UatF2ZSEBy70EMvSXSQPTK6Wsadw9sR8vf2cGQ1BRipuALW27ocXLRkXiBmQb1NV
j4ccMZ99BrgExbTe3zCKGJGGGSsD3CM+xVbYcixN8t017D/16FCat1nq8pYSXg20
pPLNBSI+hP76rdQrsZoIIw5iLReYsl+0OqkbCL5x2nXY37TnWWgOmo5IjIWzbsPz
zUvxQAfktAX26KEyHnmBbGIuubZcoqAo26oN66bnpPi+9cMwKq5LWHjNiYGvynah
e+RoJcUM7uw7CKqcuNCsGuZj8+BHOGwaiWbNE4bLnbxUD66YH1jCyCUesvi33SVz
KGkeLnI+Qstv+1nUBb056qzZxzTg4JOhVipQlGoz8JarYTQ9Tktle3HsN8VtKOYN
c/+ySgr1FMxqxMWZ0Ozz2q4aQDNF3ghd2WdpqiaR6i6+dfBkjQobpask/re8lgNH
2EvYVpZJux1VvgTVY1B4mVcUIHR7Oz3Tq4/IMpm/BoRuO27192mYZUNy+cmW0ku6
8kCSV1v/bTsLJy6ceE/fWXk3+mQCNuc9ahsq0aQ4NMNZ6X40Hr+SeJyyEGq9nx2I
LZTfYbhUY+mz299s7xaEScgVtfdDdR00dfXLjLqZIaptuLM2MggZ5sCIGeHdNgZ8
yNYqE6mXGgSVWus871hmEjXbqTEWq44hVIDB0avLQ4a2u0HE60UN8e/2CNCLOSi3
UvCrkGzXg+3Zjf/kbiWWsEI6GvKLWug/xCvHb0ttan5DC+NQ5ws7dB1kg8TMp1zv
TjpXxJhy+O0zvf0pVIkUK/4dzyRO1NkipfOtRPFTSjtLfkb8braNrw1tkYqb0hwD
2otSFPc2mdvqvkqR7Ni5iN0upUiVrEtqininvRd0gMxCvHf2965S9Fu6XMFe8ZsF
YFlp0FbAZGyKPkcPV4fpJfKAT9CtOFuP3I82O+/+TkP/1vcl66h4h/hi9105RQJp
DiGfqSUgMtijIwyAMGK8YPpchmYliBm9sFjplltV9QnTWINGgmWdanhpj47OBL47
lx2GOI7qk93xWujHMB1IXzxHDD6SYLqkcWA3XaNw4R0usjsAYXguo3LQAFMWtBDV
c6xbts8cPFho6M3LvETDoI+GfVJHNULq4sWvoyzQ8ScW5/p8jvS7UFq0ksmnA8Lq
6D/vWUZsnXk1bE1Z54Kc7870qZVM3zMS0cj+UMpEnJXkOnSgoXZh2dPGb2Z8TQpf
mCa2k2V16vmRJdCT4fpTXQ5z9hPwEHjZ+EkCs+ybWFOCUsAuiwcL1gBMCrc92xcy
PHx5laNXnjGmvQjsy/HY8E9POmPUXjnLssEMVg97NAfag95lsnTaFdRDFynBzPsF
LBS+ihcmrcNr33T898UbVU2Ep0dmLrfgGtVVaV5SgPlNd+Q6zZWN1CRbK7MHFR1u
Lom5SUtHho9RJJGOs0O4yoWre8HKHFepCKg1JahawceEZAlCiT8xdL9CN5OhYHbC
8UkAoMhFja6W06kLa0UEyA/qj7cZLPrHA3Kd4lxP8z9dFM2HY2k8mBpuMnrcxW4Q
ylHPJRfp9F0HTMcOiIPgbvXhpJKPQutRTodUCu0755WvMb0xp8qPuvgY475kM+WA
hfjfRuWJ7gSJgDsZSF4Dw1YuO63RF7rfDhN2ajo22DW4NiXm1p6pzs0ZqE0EAkre
kSurhvxokCUy5kq/dOLO5ReIwYYDb9oWJ9n67Hz/p5s+9HpnWgnz6Va73lp4pAE1
UJ50RbgM44IMZGksigHSsw1TMFxD/xzia4FaAbpwzmqzqRshwif5hBg2qQWJvNHv
UAPfbeOKjc9nrVyjh1ZQuyQ+mT8Rf/HcoNpIFjWNSD8td0siMYAp90q9TRKeu1pg
JkkIE8JtmYpABQRLwgLgWcu+s5PF9fgvY77umLyfmyuxaSpPoc3t5QD7RMLghrlf
ducRvGkkkon9K0O8FM/Q7w8GmBdJM79lIShoX/FO2cPUiSgvYQPO9npUJXKqqAeS
3brQl48qs/mOaMTjmYtHImQzG/vl2UYJjEhRqQ38dkbDpvRH2fUYPKl2+chQ4nIx
Tz3Ln1OEDL6e7WS9Nr1ixlNOMlRD0LW+QjetCb2V/1CJ4DDbbsK5DwxkkiMq321K
xPJECOP/CBMsyLYB9AGSv52AmMehh3tyOHF+jOHWXWhlUNlH+BTBr/Sn/FVsLjrq
86FNHAUI3DyNxaocP33A5D1ku+6rPGYLNIaI7NFSpT7TSDWcXyRkbvu5XEGVdMDN
McKYPUTfWwWyYuRE8Hx9j34SwFvXbwuLTnno+NXwT5IJqp0K5MskfkZj0Zax/w3i
8Bqk/cZQcQgSd3UmLMWMbeo2WoBPPIiDRrltHcT8q5y0vEa1tjiKkFX5qM7LZc3b
pIsaqsS2atqiETPppg/KqaxfM6ob09Z4DmBi44JtTjaPvOFTFr/3280jMlfFDa4l
MNxZs5+EmJt6UmgR4WW50zXaEuTDWiPR0Z4c0QYPRaf9oeckOZ1BVuB0vNcTIYXW
Po/FNBClgsK00bpalJpmq8s2u+wTHi40gDz2kW8ZxO+rGbjs0IfcIG9J8T1mNfdo
G7nk8Uma6nHm7VKABgBs+TU+H7XTYHBFnv0OOZsGvPdY4f1kUqOhaVK8ypLdQlDn
1WT8Oa3DpDBvxMj3yHVCNk0y6oTrNNAX9qcd12WXsnpVRC+c41heGV5LhjysvP52
APhO5QFje3pEA+R8I1Yl3P6ekIPhAtRDqcxnjO+5HFCE/ktG89BCCICYkGCHth26
Z4gOdX9IJTBiS/2rLqJrJaDG+husuwJYrq7EScUtoHXiukXpry2cyjmLf8+Mcl8P
kkxm/BJKNQ1k5lEwBDqiRaivUmrAERNtH2+QXStbmtqKCx8eaPfUEUJO4ZhQkBE7
zw+lbcu6EyAkZ+NOzLZ2vgt3pDLK52HjukLu0/j8Z5JH4/EJhP1yiTyQMaE5RM1I
BEna38qB3Bhtg1zwcTB6O2Ztir8pcxie/pEUSxOvZu7GsaI7W5zbt9JaLP9dlL6J
9QjXJWRB5AKhMq5xuATR132m5xqMXLxID4wx86xfozaU4CnwI8iKBOCi8BIzLOms
XE9VkqqTneus7xeZu9u74eMVaG9v1MH7Q6AHuMl0NA4JWXhZbNMA1VRZsFozCshE
rOje2AfrCn8UasIQxRPc9h4Paw/Plpy7H9ZrbTTQrPsWKd8c7E/KLZLh6GaVUSWl
SXSyterkC5ykb+7+8XoPd5oGZrzZHCbuDSAoKGp+5U0G6vVFuta5gD148O7PSgbX
8J+/FI326CuI6oi+g39YTT38ES7ghOHWi1Va7XPAbbZoU1jNyGibMTeIDS3Yhe3U
c+wlJ0a2jJIVSN0fIdq8RDLR/PtY052VToxVcRtjWQ0FeFw4wMd505G3ASH/wOLR
V2a1d+GetGbdo9FOjj58ONsimWTfmfSEEGInwetuSpuyh+56JYLjHwnoU7Rrb/80
bevhbM3mi1zn/W2c2zxtRSGR8kn/rgXXFKozGdzA8JSHRUfLVwMIxQi2AFmQPbcb
PST3IaTVVysB2KFwte8cG+as0+dE8XUfuA2YXWLMWadt0KOZbtUoRX/H70Mztvmj
3x8UkXJuDA5ChAEnBvRpvYKy0XqEuR6rtGCU1A1h3fm/FHPC2fyy4f8yy1ti2olG
u13sWUQrcdzqll0sqcnCoo90IIt+b5BZbfUtMlU09z7ba6UmprO81padvD2K/35Z
QKAC3hTMeJIWy+jDe7Y8hZZhoZk/KhuMT46QfEt45D6o5Wvs89Zckx99WBh2+6JL
y+LYXpJtqO4g3QCTD4bjoF0xXVpy/hi1MZHDZfc6egWS/xm+QnZ6X1chm2CZW4Wx
iFkjV1SQe4msqMagaUguXm7+00Qrl11d9yhuANBQ55Jpc3nTt4cLn1FGa/gJX+hw
Q4wTvEnBObUyy4GTBZu+XlFgUGZ7Yb0DWRca4YzfZ7jPwIVRo7r32l6ZuNx7vXNW
dNnJCNn5xYzqEUwenZ7lWOxC2WhDbpOsptT9xO2hwGyzREjM6lBESTlQpobxEZUr
8kvEF5EXQse0HFaiqF3dN3DSuHY3H9cSIJrt/10dVMG5qeR1RO/131FUFzsvy5Bu
nj4DSDoMTNGd0wM9sOO9cnury1Ysjij1B1d72eDeyyqDaus5pQTeq9Tx5csGbXSl
GDkrbef1YoaVsLV9vJNSlMcZM2pv07wta1NqbQlMyloj7h8sAG56ek+Z5GE5KkPa
fCW0y4jG7T843UomCIsZt3AW6K6vxNsfNy2QDAEJpbSSaxi9IvfzNfRX+kxWO9R8
YKOxc4dI2R94mwNwZyx4ljaK5FU03CPyq79IXm0BVOJA7dR54dZ/IYwXqafAZXBe
BkMtHJF8MTP/ClDObWy5w5M6po+2DuyCTMRSV/X0oo1i3ENwCpXvqVXvKsMCS4aP
QGwqZfXroNpJj8/I7tEod0KJJCZpo2QdoDs4l2QdR6iH14ZYMQQ1yR+TKeVhpCph
aTMuMrA5nmLo0lS6pPzYjgmIWSr4ogR/1QXedE1Rxqo8dr8PwN95yckOUiUiPQF5
xpK6C52YXTQTKK8x6JxjsmLlHdM87ZYRwEUg7fd47LxS+u5S9+Pndb1xlAaPo8Ka
rVhLgR1Q79pXuzuEgnEjGBpktpDEi+EHG6qh+gyOBDpHkJKwn/E+d6tbDAEil/3g
bfJG6YLkkt3BCvZezfd2Xf/fqgamvoYv2pf5/PiD4C1VTdS2A7fOS8l2Fz1gmmUD
IOXwqloncgl+lvlJDoiVtJfuh1SV6D1DYQY1/z6TugHT8OA7hOgsMlXZcRuMXXIg
SNLg0l2+Pry+OJnzTxP41VE6gE+wz577+HbQzTKduTl/tZDgbqNnFyaL/9OIWZjT
QJahoGjKcvtuFwEC0X3OxchKzEFYcT8EytTM71hyKoHOg5E6WtnIzUtpVEh06U96
eFS9kmK+fxNKL1kZWkSDiMEIsBbGW2h7a3xIM2/iVL9PMkaOcmHXf7IAC6dzCl/J
0fUGSZgzCStVlpp5uJLsBH18BmJb3I7n76012WxEogBlbHHU34cTcIs4GL2ATOvN
Xwx9ZIpPUVKt+RGwEWFEuQK3x2g4yZXui6jYki0t7fMRsHRIJAflpO9rQ0NB5L9f
covea9KCQqzGnEMAeB/iwTQD5aX2z1X4Q8dVQfXYc46paErAzdvHqoOvSkVsIRoX
KjnYWXPmAIfZ0yBdRMgnZR17oPhfNqsCFnKbfOF03t5m6MzDncZrfOl6VzgHcG1o
En0Ic5Uaf2tQ4K34bBHQAZxQkIhh+cduMEfttGr3Suj+i1xUkoJV0f/OLmoDQAvO
3+wkPseaNfPySGdVf2RTnQ8/A+HG2iq+zUvdg7tLDIpUNlu77O506bZ2vUKRhSAO
8CuWwMTu64I6fTB/2a21lg8fHa4T9EMX3D+CrwCCOTOxH/OuNL6wfasJTe/It5a6
gDtnN5vRfREsKrnhlH1ZUvsNDB23r1I9GGUklMohREOBZrKUwD/vPSvEit4UxzrZ
iJDQ/R6hfq/rZ3VI0Tlnc9qwttnf+C1VdIZ8/My0i0ejS/YdQ5OBKH4gh7rTrO6/
BSKe6Tqvhy8QJkg/Uco6cN1DZHl639NbDCX5I4IByAV+ZneRQt63EX8Q8ZtEt9F+
DPIz0gYowQs65ESdjuiMDg25hHcufwgmYai6Zw1HkytskNmG5i8GIPZ/FE475h5h
+d8vMVEDxmw1KcKIfWn7/BwVkrUZVOtuRelR0gi5yhPzBDoak1GJi96n8uMB0oXV
guW0O5OihLCdYybzL9MfpNkr6YNLfu2BVJI/NA7UYY0CoBU0nuZ9TR5czWRtV/P9
5YwYrg7b/7xyrFA6kR1xhyQkVvmUQoawdYfbN5rWzIbqbkwFnEp5uPVGap7OnkLM
6WSHIMbxkB4Dyff9E7b8u6YVPEsZI6MAqB9j2afbe+5OM5v09d71EXN9eO/65dYA
4+0SIyWWOV2KUPYIDUV/uta28rTssTnvwAI/voUFEAY1umVP3oHY+PuJU+J/oI8f
eZObvLqh8teyhEUAncqHMIypGjkPJmWKdVph7HoQ+EPXVzoHlbOlx/S82deqf9fB
GVfLhDlYqmoDmCj0vPt1I1lseAV816Djvan5b1iVx4QbSpXKxvKS46HaRswduS4F
csXpjFcYX5mZFUs3MeGimzVyegnlevo/HuZ8gXg8ezfe09ki/gqlvwaWw3tM1Y5H
D2PWRCtALX4aPgFgsYI0ReznQyO+DURZgs2xfzPQNypYFckNZnISVWExnl+nzYBW
zQ8XSF+DXjHhy7RStDuXGEA3+75lfKfyDz6xUofcKbjwDUcQZ9dLAZ69JVIJB/fi
DMcB/Z+qQZoAmxP5mUx8BfwOU5U+DXm3SPnbFs58n8xsEx9Xd7YajJJpLD638kkM
h1ll/VP0san5Rx7iOgvX2sWmjk1btg/1GIcsW4KttrDlWbt3bqhhDnF4YD9U9za7
UKQ43UWKhzTxGMwgvj2pOmgsYsvYrnCoRqO03kjlgzHDkUemP0blH2265PxGtoWr
DPhdHJ1dERungfMgz4T2nYldvsMCuW0IG91fMEqJAZElUEnmMm5wDKXR64CABEik
wju3H5BgOArdFqgtZyHhWQ8V6ddIMc3bVj2GjcaWwnAROikAZRP0Pbdc71vRcgFT
cmU/QSxCrPuaFiej2ALmXGdZ7KHkvrOIP2tJucC2bg3/hxSTLr0ku3/PZKfl6V8D
IXgf5cm+vmbV5NETLwGxoOZgxltwI/gSMI/p2TwLVaSfTgVgEusZq478U3k/pvcK
N0+NsvqS3OWzA3XzEeuO7qfdPd405bBvzUGRQ0ag1yg3QRT2Mslhmjts1/c6cDPk
o17TwmwVjThGEcwKvkrnlZvKA/Vei/nDmZvS0fTkgCebbpqSNClVLyyqgVeTv0mX
tNYAh5P0T93Oy6Sg+Ja1nxT2KgiIx+PSdjOMpngJk9d82Y5FSKQilkXY4CmBeCc+
ZvznKXJY/Fd2kAHgH1nqoeAAmtGqsn0CtP/1/tp8AOTO5bzwC/VkDC1GC37b/Pno
NPYQvhQxQfPz5qej3kmePm9b4FUrcL9VR9H0TaHBLYjHc0U3sIdj5PtWdjM3TBfq
gm/tejUX1nLqS+aUtNp2+InWtO679m3Y31WkFZA3EqzoB4jdUInrv0qZRa5KLh3t
flushFxdsA/nXsiM/EDITtSPQrV47K4iGtGHupC+/KDIb8WJtqIQK5G47xMXiFsk
rjUq0eTHFwA2OHeIAP35lbXqubnd2yrvMKjadNavhwyTfp/fZ8x63YzQZCui4gbc
ARb0RiBUDt3Z61E0gmxUeQD5lPZt2KoTUP70FfZQkKqbSKh1s6ZBhhZxfAOLbXZ/
Ypk6E0INT/aJrhZ/dlighMl7uZ0fXhzWiVMA4e3tdiCnSb5sFmMPidU3pefYWduX
xZLBdF+wXAFKmRsN1rRAAY7dmp80SV7oOWcqNcGyWqlgMVqqLnNFXBDykk779etZ
XRfpDYACt/DokJblnNX/vujYMhMpdkhhAs37gwsTuihiQpNJsjAAcmKYvbtmuaOA
ilJmgPYuV0QXPTLbriWbR7aJuH78lWC7ifzgz6otui/tl4UHZF2vfOSK2lMQkNpM
ZBu3j7N8jpmMOcTmdlS8BVIwvodGSE5RMB4GZtggwFmawXWgbGCl6QcP0m5lzBGp
pZHmfcaqGwrACyBzCKy4eJkC6WBTQQ9RiymE1r3xkb8X5noEzt5grp3yW4liuixW
mmvRMT6UZ7F89YTYd7f/mjRpHJkeH1HFMEW+4VvP3s34Se84ZTzpqCy8RDu240KZ
r0z6LVT0qmHhwfzea75FxCwhCwQdjMjUkOaekm4Q9Jjtc0IjRI9K67BWFb0mmUsC
ZOGhHF0Kqfk/+2bzxWhZT43jaCif/k3SpX/mrJ4I0i5QtnC/J1Pne5ueODEBbHUP
zp0dDA0TmTd4c1MRSoIJSx/FX0XiiDORW8Wb/yLd191GBCQ0HLvS9jqbEPhknyS9
YCbLL98pDIraOAFToMOratpOpkZm6WGyYvT+xiEf9zpqTBlaX19NHiVgSDJd6tAm
wQqRMmjQVBbNFngho6ly7I24dWo9hgjzEtUYbpqy42cZ0SvQoAHuPhOi98fWzuS8
wARGwxvrWTbZdcxEmGhxY5MfgcWX8893p0iqQDtSZCcLcfZj7Czo92qZEYArf4b5
RNocOzznif15XY59YxKuRspESDKA+Ud32Vksx5qEBS3rCcq6nsjdIzPmTAeJPe/s
YhA5F+x+8DrJAUFfM8weQuDtfjiQbAvykAllm4cmu4RTIliJbtI/uPODjC41DcWv
qt6YHsZbjXLFXeI4wMGTyj0uCDA0M03x3Wd+57IC0NO0LMFm7oa8HTRtOyFtfNT8
nsrFA5mPA2IRE4qIZippWFg/+KNtBtp8RjENpfm4YTbMGFaCcPz4nUJkjZGv6pE+
DVPJtVqfnr7MTrrbWnVxWmCiGceN4zlcloUbAZ/6MA7AV0w5dqyyWpJC3h3SO1dW
XnUY5zd3Ksd/swB4+Aiz/J9+BetHLhaHRiMaIvmvZ3MwEr3io89fbmJXhbIEEdXN
mFRet0Iao2FHQ7JIw4Kp+98XcrutK4K/jqIqiaG5Iy3I5sv8Fdrai1YO24qeQDFE
j4Qtr0HI12VLQZA2RYZtPAhiSSutFD8jLv/yOZ4FwKgotOmpEkBZMGlRbpPFEe+H
VHqBw9Qlh1ZOCaV8F4RraOARnwxBcqdeOxayAvDS1fb/hc/eGhEl+VugpEZ8pCEJ
5VmuA6Sz2XtvaTbYs4xR/tzki1uaPtAsysX7+NmJjTA4ch+yVKopHllsHFoLCqBE
02J5tgk/XMSvS1igxEIX8F16Q47pFuPJwt1jOZzeKSjof0hh8Xq3jNDlhmK58fpA
ylwIpVzxyQCVitgpOEs5l1U6z5EV50kAm0zcIl+0IZ/EW8XCsOWEsNgpKbEqtauL
77qq2jdeQeTZ+dFtPZ1KqKrGAytlf0sAh/mZtR+7A157YLSUsUbslg15X2I+1525
6Ld9LJbi4Ohu1tgeXCPjobcfG+PSNdHViZ0X/YZNWXBAik3e+5xbxTJfN6ucsYaY
fHTmQlpt6aWD7vewVCIS3iA+SI8N6TzwL8UIgNW4fyimFVoLVwJMGOLRdRfYPJPB
hxtRjbzOV4DAqTQe82QDsjlJThF0AIq6uziXDPEiWoSD7MUFbv1frbINzJTeTCaG
W7XTLuRtpiUfvjmJC2cqbSgp+lxkFY+z/ymAUaMhbH7sYzazJAXUXrWQOy4dSgOB
20iWrwm4Ly/2ArByutF6Z6xkw42y5l+JmaAATJkhN1q+mQap/3ocA4Qn3f+MUaFr
ZkeHq4peNFtSYHbPKXzYIoQjQamfI3fsRjzxNiRMACDIAsiPbpzM67K9Lfye0Glh
fJAcDdBn9IpZ8FHCWn4VlQueBmTn2pQwfuFf24QU7+/DlMZbkDObGgpeZwQciMKd
SRhdTQ2RQJYVR/PS9r8Ufj3eour+Hupj6QjxWChLXUm4t7HPqvexMReqF+8jhNPI
FX1edWuPHW9HhKkP5nxya8OFMnMrHgkUOg4lVkKrhl6PPIrDRsxpEsSqRCwS5OJA
+NHqrflV0c05Fbxq3cXfDN1Xe+hBUt2gP/iAIOc7cQSoKezLZslkLJzAn7+ER6wT
zXmVGyOBOIaWGgeQ2aHmnfMWCNuF7TvkVNfTfKO5Hov6/M8jcl8a6OsOGrlUrVUD
mSCtfPFEUULK2V5Vvd7KiRYTBK3GLOmr8LkSMWIMcHB76NR/xskkBAkxKGOemrTc
9Umb7z3YcFe1BRvajXrNJjKPavrBh+ZRx7HzGr3f0z8vsHyxPk5cRJLtBm5xPpHT
wNT6IYd9fk1GwVqolum8HNDhIvTYYNVn6m++3Jt6YfF8yLiv5gN69tccu8KxtDks
SBM7+jOFT61ez/HUbeyu24cSU3Z4d67up6e1dNa2vGISCtx432KoQMRYsVzMt377
hZp+5Ab28qOK5NFnw6AVO9nA1V3vYvCDoNHD+vcFi09FZnFuxBOx9EIxqkCgGzES
HrkpM8C7CQ6Cf8hCpwshzutAua4B3VTATGDeSmRMCbdmRwzf5VNdpeNNEl3il7a3
Czzt9mc5MvYWEJWWHMlzz9NKecJzjD9N+8DybJ9faVss7qGuQwXFhpZpYlkmKr5q
tSGAV6hkEO4SBXlMJfyHlVhyuRpB7fs+bvihAZ11LaGgu68JckaPtNHhjEQ16Yxt
xOQ+mFMoA9wrJ14G3QN32dFGZuCvz8ev06nNfj1hfUGFWJjhQ0MfnRMNDgIqj7+T
0tQrtYvauvzHYW44/hsa+Q1UZ6ECC5EWF6zEZnpy1yax+TvjmdGgasieWnydL8XU
TypCICfYlRDUEbkZ8iMcB6D8vg3SJTLkFV+GtR1S2tUKx+w8wjZmEuDwWyf5aHC0
6dGN9O4tgWfHK2kUv0ymATIKeO5RcS/dBYpv4gIy8uIC6dGZrS3sUTqbSbOOO39/
zsh4/eTkKj/BxHJ9zCtCdJUcPW481uH+wwom1JqH4U/QaWf94eCQ570N+Egxa135
dGrMANtfdR9OA3ygFFutAdVQHu4iDmduBhvVGlZpeSdrRmVd6DIEeaqtwCS4fOpo
RDCmACs8eprNsoygLQN2dAoB2lNLzQF+53z5H62jq/8Zs8ZTT5HLnpZf8AMhafLg
GM0PnynPs9Dru2S6Qad8ecShB6utznOkZh0CSbW4d1rOprc4cBfqKtINJmqTFy9l
BZCCIS2Z7ee4VSEVvsekjtgVxWueUuzSc72pUkMgorv/TA/MgedU1pHclcsVurPI
Ri7GcwCBCb7RWOlqXLU7RRAt0EfE7leEDk7Ck8M87fAciJS5TTCWF/J3w3h/A8SU
ZoMqKtZcAOEOzJX19lSNnXe7Sy0o6uBZX9LSIpBD73dJHmWMUv8wdxw0wMwUhJay
2h5Knf27DMGo0w6uc5+LrFz/EoX7ph9t+QKIKlnCVDxAy1w4xKCehgWU2jnIYkJ5
xao85PpF697CqiFc63MkPqzJ61PPcGDb0NAAD2KAeDSajl5dgNR8MUVuKVE+2gxg
bKGf9HITv1i05tlxZ4YrvwqwoztC7c+42bHV8d2oPHlwjXczcPd7M4NJAJancPty
qCprLDzd3bUOlpolwBkoMSmg5BsdcJ3Tbs4ZaKehqSU0b3IHXLxMhIgt2HOCtz1v
IvSEydOgTyC+D/RyExEYi0csHxgYId9qnuSHAMC1MjzfgfnQtdRIvG3i+9uEHbE5
0hwxN11/BYi3MZVuTYfIeur4zRn5/KYkKc1x1e1YniAkWOoA4EpMvR+gpe36RIh6
yur4eDlCLyi7bZ3Lhp1GxIYXbVn8QLn4on2XeJsFRISMQsEed3qSCjaGV6ykOMVu
PU+XslW3vuiOC09dx1VUluAkP5z5LtSvKbRcfJdBpjeapO8XiFdXbFkMmHiNqbDv
pqcu9EdjlEBkiNitjAK32d/I5L/Zou9BI0kVrqJ9bR8AN19lcPbOOgXakU8f3iOK
am5CdhPFe4JXe2BA7jHyDbHyHDxpXVSXR+2fSLtyW5xfNpeZo0km1ByeBAnrMYgU
cmyYrbYSe2x1ZgSQ4lWmgn2x0vAYzk0FEb3q1pN4FMchgsn1SukQhe7KQVLPakpq
yOPjjuGcYjBAKBC9/XCvP+mUmAdUd+fgzIg0y+h2TljZOSdQAQA5xbCti6DBHZqM
ooDWQmDL469jxP+JxZO9ZoQUOVtqyIDmQp5tfuKmgQGUJtlWZxkj6niTcmJG/6Aw
n4pKpb70DnGuWU0rycihSih7Xe5f5petJiYCpc5/pMfBLYRpgBJ8vMfBulLR94u/
uhHLLjh5GT4i/GzL5R/8zkFuLS683hBr3sPG9NA0gLsp4AVVdHVxkziWRWNgCPBB
gbiq5ATS1d5rDj/5ov/DNcnz9uG3UnuA9s+9IJG4rpjEUeThWsl1ad3dYc4BU94m
mxKxEm4wqDTknTZ1EY5XOC/A88Egn226Gsf2caP+a/k+3Z0JyHCJQZd2ysiLVPHc
SEamnWv8LeX2HH0fWAc+R0Z0KZjZJSV77eSgAm0qvqelGEg3Mvk4buL04v3QuiM6
gOEbLzIpWbpete3igf8isigR3R5LwT1tb4exGdDW0iFCqA8AFTwOpPFen2Db2OuC
DVbAv7UDr3mQ+PgtfWvMu0qUgYol2/kAb1XBHBxFQwEVXvrbdDzN3YyR3pkZrrM8
vtQZCGcMrKtAWOIrTehi+PHq/YlqZN/UeaOTLK9QObPfvSFLumpk0jT3/KX306bW
w/jlg9nTozNwn3ilToSUMqAE3UTniVE3WKzYL3HrmM0BIbyRxFkBJZRz/38HlO1z
6ytKsAQi7Uk8aU/gKbSZzHCVdr3sGeKB9uKUKLNXqD9eXHCAZPSrY1wDSQzOk6MB
e/ALwfn3Sfg+7gpVJGgy14plbpYDDZxCiig2JEjGH97eyPFnlGxdOVxlYpbM4tNj
zNQW9o4th1iO+St/F0sJ2sgC+ZrCB6SxLsQBc2EhMW/SD21TpIni4PDPeRiQmo8j
ntiQmmyP/K6hB1jEmxAVED/1gmCTEdqxC1QYGeV7VSGB+PnjPYm4pNujXk+yYfiv
Ou3yFmd1aNIvTJRXwG8XzJd34GdPEJ5T6zr87/3d9/2Z3KVImA+4059YzwdapW54
erJXdKnmMIGdGCYg3a+aXIYXse9b8nnvpihLyjmZ7UQfWYUq4pcSAMm6urxADxi/
4lvpVDUFzic4MiExX2Dl4ytv10dBohaRldJ4Zl8Jz0U6orvhEz3F3V7xaWt01ADj
3OO7atiOYcX9GRXXOagwzBUeJi/+Zh/iKOAUGOJkiCmXtTFlSAa+pxceOfO5w6+L
0m4vFtf1wT+AzGJ1kjVP6LilNVYKYbavCmImMwd5UCMi/98MIgASjVugcMVezoqB
Ymj9ukReq++9C/BVvo9/aAuv6nrpP4OMvGuJ8d2g2/AROxJTGXScMNLkpZm1HxIb
5Yl05BmNfglEh3iEuEZJyeNoi/bHlOQZk3HLGfcNpOVVCm68fx6zLR2ub6Smg2yz
+uufcHnSb5sYLfiTCsiPVLF9NITgaTMoBubWhZdWM/TLQ0lpW91Q7ed0Ip5m3dk+
5TADXks5vYHTjHDH+y2xc4wrvIMl+fT70mdIADTcngFB3XhS6JBMsyYRA24CkRxt
m6C1TPmNLWOzQnTCGvmCkjoxSlcJECT2uNhuBiXDVMMU2ad7eyrMXFiCsYxACuyO
Hcce/lL4IhYmQyV8zM4rFkSfgj5p0SpKxHevrZ64ux8LjaSIPyO9uIy+92AWmrfp
vmAOmxGuupYmkfSlcOVZzBhU8W8ZZoAw29e2dGibzzq6zQ3U0PnVFcT89ljB0exK
M56u2zMg6Ya3NRVhJ069zFy2FORZVZlxph9eUx5nJOPIOGCY/3mFmylg273/liLQ
Ra05kqYJ3siLJtL2cGF2k1YbGqEN6nlzJn0SNSLr+uO6eQFNwM3Hi2AE1gyxUg29
Oa81sCIGrR3xm8sypchR8P1w9r/6Turry5r8LOMOSIgeuyVtxwjMjcgrCHEdnMqI
Daeuebq6bgBAhCeXx9rtQzOW5MT4MHWVi7xRnmDluPe8nrdI4dBm8392qZL5Rcu9
82V+EbxXLlOowxxC1paiwD7U2ua4maafoilV76/h3FRs7yNua0i4wuO709htAjvu
mAnq0Rufo555XEAqTgR+YioGooP+4nxomfpGItKQ+Z1OeMjwiy3aRD9dUbDjzGnp
D2th5F2G9GSGCNQC733qqA5cGXUe3744BLNh9W+vivKT0fsUrIISGZzFYBN/+fVB
xWgk2+Gh2hoqhbkkznToX+vLRncwsnAQmEH6CTej+BH8yKCM7AyzCNw/zkXdFMCS
UHv6ZFYNaWM5rSGctf3Fmr6yA5v6dVIxoSxpNZ3ZfNrYE/pXaH2lX0srHsGFDT6i
8RrZufTkVJgjkjn/8Qt6E8jWIo2KRy2OvUAaKrxWscvuCL821QLSWWmIG/hVeD7q
ZWzw+X5+fArIfZcRzhsvHZOfZPiKMGSWM2T90vj6++mSttLzMDW+19OLWBsf7dL5
lLpkfC6H68QbCIec2LSVdPwqfdQjXGwpeTEHA2poj6F4BonTZ78V8diqVom66W44
cjZuOXevBFARGDsa7jLcP1mTBUG9rBsKOPHMuM974lXzewS+3XF9TjjsD3sYGtD/
BPh84ReWQ6evcWUeuR2eI9zzTd9RADIFPJkgR5zdteCTzUE+HQml0HKM120vtg6x
ntpmLuosAqCUhbRQVt9GVRUS3eaLbAsZ6oUa2IndtXsdMCWYSdr6LTLi4ZvRjttG
K5yXaeH0qqU8W0dvpQ+wznll4Oha/t7Pi0xeT8HtgTKKs2i1cL9xTzM7L5LI/raq
MvkIcA0ZR24I+9LReE/y9sHxai2+bpm9FyQhBX1NLpB2Uim5MkmsgWLqsPY9Q5Tq
J3UZrce84G7e2BM0kBVNj2IUti8Q75och02z9rnARDW/PHRD6RNS++bOzOQkPeFp
wJKP85j8JSDmD0ZNsG5526GHa2lQnIdvgQjEpFm6nfnE3pO2k+hPGlLELOSjcOe8
I8RfgwHNjdUW62UrAZveEKyNGC9PpeyzVcBLxyCNPE5dZTzgAZUFwXLxEcOm8HY9
rio3c1YDpriSuWHYvdBuMsQp4l32RbEt8jFlpinaYxs/fFw525u3sCxsQCgNpSfg
uIgbvrC4Ss0WjbjglOxj3ZJudnJF8Xe15C1lRVKVWLPKaY71ewVqRhh9d1SK/tVb
7syhqxHScp1E21uw+vFd8x925B/oS07nXacIJ0PwOY8sF+0P6DcPu5jX8LouzUY4
7iNz/WiEKXhX6oxj1ab4HSYSKXUYglnU5y3xYm3dA6MCKIn83KeA6f4pOt7SPJFt
XnLIrUsUPsl/SOiBwn7nuuQ1CwSxljhfZxe/D0twRxft1gwqDN6/eEBfdYE0EuW7
HTWkSIAOr6VhIX+HvxedS/M27KYJZ5KLSwsXbTgwPeHQ3SHafAMTi67Aq1EV29Mv
5CFIreG3oHr5OPPQK2ETKg6qM/HmAf6HPbKbY1Dyox6SjlqpvYrAnHlewER2igwQ
Vli+YQMepXU+f1+QK1jVwRfPQgXmq5mu3HhnYyAryB0VtYxHPFF8SEgwwjuC188l
TS/UDY1HdyTcsCDhgLFf1QVQipN7SshHyMPJk9n2uzcXAKK6W9I/a8L9A7ke76dW
2l+0FZ9wAR7/T4tog0xKbJNn+nwc4wu6wKN2bB7fLpTmdyCtS2VpHJlFOkYjvxs4
zi86b1GKsm60d0/Iv8sL31OIFem/pcWLqv4ebC2EGKRv2Q9OXVMD1SxXE/s7jEVE
kegVb13mmALFsmwK4Ym+9W72fKcAF8f2lHMWHuM8eV5RbqRKEomjL4HyDGeglLcw
wOOIVYeMaJerc+oS0p2vWMWm5TK+lXXGAAgDNWYu5cjGcCXgwIuTqIFi1h5mSiuS
+ieDmYEKSIN9+pVYPggw1RAnxA+NbUgTJPwEyP2NssSZfpX2NAjaJ4tS8GP5bU4Q
4NkCugRgmipW1u9VitBGCxfJ8tD1iA6a63YYNApnae+tf6pYSxMUJdt4OaNlYAu3
O1tsj/YiwMsvnH+ltACsKhHL5/71Wc0uwJa8g6A7e6JfCvf1flycba6iDgGFesxt
e6bhaKXCI3E0ecCTEKLjqlgrT8AWb30rVvhNV5qqLXQAJhS4SivMiyTRkq2y72DY
/UkKfteQsC23FyuMGsN2F8G0UIKGLNWAn8CerOS/Bdfhx9BT+AMrWETVJ9N/e8uf
JTIkL4Yw8cOW6JCd64z1DFe8N64Qf+kyzQnk9HHmg4Ej7Jf67GwW4/tM+/Tv1O2O
OiXbkC4dk9di0gWyGjGkskHLdE8hPvzH4qIwgPmy0YklbTMblRH0f4Zirxx1b1lG
ltwwjFOnNSG1mGBNFkFiLeXr71KsUj8e2IhJFjijNPNMwlxd7lHwevrfoy64e3G5
veHdOwso4n+nSZmmZgfgIIPTULbTGr+l5n53fSQ0pz3LyQg4BrzhZuJ3OmKGHVx7
LPX22WMfpAoCe5WyqjZhkyi4CLL5PHdUn3EEdrBAxvsL8+7iBdmwjyjwClj92MmR
TtG6c5zSWZBYv1o+XZOLdX09BzOYFNvC2pY9d2fPXgukdG3haY8kkh4je0Vvu5h8
spfhYnWz8DKKB+9dSvP7/UVRMHsKrVky875xX6XZ2bx1iR/Q+eZb2SJPVIZDN17V
qPvvXxQ+V9Uu9N+Y6MubinYp2fjjSzLA+bDn6CM2JpvDHSqAZ5+8SqM/MO2VKpoc
IHFw/obgfg9Xt9J7QhhvL+GrYdO4zO9wRocQhUb6isr7u8InzxqOv2WIAkqTkgJS
/THzFhjrQHgcQt7akN4IGuY667slv1GDvwKsLHJkP+AxuGNGfP4SZqvHFSRJenyD
f/Sn6+la1a5SjcyvjRWQB+hILKK5xSwglmvYWq8GARbQYWkn825ZOm0hxQ9SuyRC
cdboLoJPYUP0krelXQdULxFvFtZIH5RLGIeiJ55FKAnsIo5oFcVxcsaKfWtwUdja
LMsx6p0a8R+c4xLRW/iOAWtcL8az+GEbJ1KpMFpZ+m84O4Y2zJz8bbHJrMUBnv72
zrD1ayPJIDfmASVkmw99w2L5qzs/a+QOCl8yx1a3VNDt1ZRl/6EKFN8D0H89Ie2+
ZLXu9fy7lwZtUGLHSNvbr3q56KbX8n0AJmoBM6E3drOAoF6v+UhX7EC139EEOo9U
7QWy64mX9Cdwowcdn6sABJGFVRDDGqr+q5jSOC++PoI/45GYGOoYWOAsFqX9mkxG
17lg6ve1G53W3/mlVd6ja9QBEnFn2vacLoJ7rnGjJkRhOnkn5MiDs1/P7INVAvQr
2PNBBuGTZ0yT730/U/dnMGD9oOmK6AobS6EJBH4cSCXH+dYtyrnQCx4Zb9wllxUe
y5XXs+n9hFnD54Ydk1pcqA4sqVEeaGqcxSJ5briuzTaBfYeNOMkpaTf6raL1YzF1
NctscYjGUCvZ5CF3fPtq0wR71huzNSBkMoa4K16YkBdOAzvYt7EWHMaQjhVCyC6k
7a9gI15a7dJkiJLgSm7a9fMsAl/THx8MFMGZ4LNqNeLcEv+C4zd53IqQzQmF7mc/
brWmbZBJYDmA/W91E/WanMODuJpMw/1XTrzCdKU66ZblVUdi7f+KNZrTe6Ej4m9b
PrpV1onCLVGtFcmVcmqtFxsB0Zxb209AjZbSuXtw5bGNvnPlU8f6B5n3qLGaAxcv
jpPM9g9SwGXEJYs50uvJkqfSPuQvDv2GTmR5+E29hfol7Xa0tjjuHrSmkBqZq0AT
rXxpwjk21JtvZm9Ju5LwrTAy204SI2yba1110GFXvZ1cF2US+46JVjooOvSGuMdU
c5u9Eh9WbH/2E4kKhsITVKENtPMQBGFi/EL3mZpeUm43vzKhg04r9e8ZQ0lWiO3x
XlLkro6AhPyXShPlq4O6ZqwwxxmN9GTfkvNty0FnkSSOCxRt3gknnoCY0gpBmBjK
EkCQoij/OiZZccxlvoWRqxkrVmD9IkeEO59TWXN7z1fZkvxahwtx3LJOCSS5F8Nv
bA96oSenGUfo9/Ew6uTO4oPNmiOjX+tHsh3TwxAuYcaM0JJFJRw79j0C9dLbuTzv
MBxnm9A5TmRnEiCTUUUgVm0lO664kCWsdM0WVN4cVn/PnOHR8avpzNaE19q7uP2N
LCBt/bUF1eFPX25pORy7D7JgFe221Fxx4B538PHtJiejX5BpbGvTzLm0g0UtGQjC
g8qVjGa3Y54j3eJeSDuI7eK+iPYkovxGIweSfmNA5JCoeXe3JrWLrSAR48MVqT49
Cb7GxouQpRrGfiUeQugxy4gmkHn4tEVWslDTFhh1ZmdIdVpjZE5ks6cWDkzoFoq0
r2iOd7mDvY8ihbtUhoVcyy4j4EBwssXGkkO6TW6q6wVO4q2kjqJXjNwhNvlfyHmY
uPsDyFdmbLwVn7ymesSb5YYMr6XY7b0Y2pS98RzTWumBfdlhbjvZ6cptAMt1PJrL
Pm1leUhwSJEPbPTkqCRyGg7A93niYsZ9ppR2e0APmYYFBUMX3QmF9UG5ReF36a1n
3ybYhHVTO6uAqgA0JjXa03XI13GxUatSMJHKHGQJxVLSqtM7m/L6iXxSinjh2Srp
ZY4Qp9cbB0iIKZxGAURoyL421bCOG0LeiuxhXJ7A8Dad3vL+MoOocZcACbDpy/Sf
jYo8t/57ZP2P0Yy1qzasQ0VCZbm+hxsLL592gcVpv4cTIF0xEwdprMSnw9SmentZ
Evqpm2mcrSsO0R+7JoVGKtONyGCQTf6My+0muLwlJO5QDmdNgUvZ8qHB7m7sQplH
WBQdPe++3M2aZcRYlk2own5Y2hCLdPyNkr+IoYhoKSS4B8QIBAZVN1h/ffaqVTSO
5+p80O+l1hHB3GNrulj3KtyqEZ1W8R2gv8rkyydBw2d6Wmx7ywEYCgij4w2yndF3
+G9dWimpxZIkbWz0yr2ysPcWZrxC938hnXI8xhyaMse8axyth6H1FY9yOGLnKSn1
vpy1qd2OR18gbf0ZoYsPIxjXkJUt9AYlyy7yBNsLl/3KpcqmDbZyEBQkIB7UTlPM
x/R8wbS4N4reCxPdInL5mMinbJYjsYMwk0M1zOpofflvDDvVRwwD4p4RzPNjUmUx
uQtWqsovn92IKPMapXH/j7urTqnqPjqx6RzFsLF2fgFgj8GpD0vle0kMGz9usHUW
KhwmJUZQ1iIVw6r/yJC7DDBgJabPi0u/SVQ92EU/Mu2hqBjm1Ac1Tn2npKw1eoaE
9iScG2zZ0gsueiO0jcMd4VNb6TbEpkJapgt96rQicqe2kY3VKQDDZfpv5ur+soEx
W9i3gSOXNCeHpmHzNsyDRb9//w8uz+3n9rVSrUmBJsR2tHX2xMFQHD0pn/QKhp5n
blRHnfIP1lwU6RgZWDQhvxsIp6Ib033Q67FjdHAzgAx7t/mHgjRqKFWQkGT/L3yY
e/uBiDTJpkPtm8+K9QUbpn0w8r8Dkz+JkERd4wAbYbUNCneFHJinNgW99jYS7YO+
kqB+ZGG+cnEF56883u2hzPwONZaBRFOP6DkOWnoxoDEuHbUjyS5osTWTkhK3dW6r
H1/Lp2CvjUCd94qScmHMSIJn7WC39dp+xcmc9CVD5mIYn8SbVpMnXSsjFv3SAiHl
UYi6QT3xHfqjYG8DKyoozueOfiQiMZofyogD0VIzDsyVQjlWgzjrJJ5JmKspJQMv
+V2fvhL4FI2aZFtLNY2NPrCyb6HBSaF38VqoItpLMa7A1QyEisSvnjCR2szwqJvA
B08mvPxUO1JX1Qwnm5aOJLjsQ1xW2LapTpRp3iXBmPuxeV25WLMKk1sJ7OEz5NDU
oAPd1bosi6HJK0oYu+SSEFGwHgTUfJIwlFeMUbxHqf3BrLz/brM26i48rFmqS7M7
7D1S7go/CK+ct1sQ/CX3iHcvODUwW3gosMYca14xfQLh5k0a4IBBSel7+iGHFnzC
67LrT1FTldnqm2bwVddJgox9AsF+5CmsyuTjMu456qV0KCL7YTUuC+DwrwIDLu62
/GZkJaRYBselrwvxp0bzfVodqFTOebPKonbDa2CPArDV2tJVK+Pdzg5o33Frzlse
ysdYuyUbQI1elLQHsdTrzuGd3TBzMe4KXuaNTd9erkSNJJF10+8sAwFRaycDdk8X
ouOV/r/4ckvK5xa/VDN6mJ65jkRFrPhhp8kWmIdQwe/cNF/EyyA6xpd/Ukeh+bg3
CJoSQYyaE3kQlbA+fZosfSh7H6mdLumjMY53zsgftwSIK2jf/pofZqRS+oE66I4c
coTiZUKME47/yBoHMUTFQ0mZJSaiCRZxJz3lNKd+t4SJkcifd1m14vV+lhr82sur
BNG7ox1ph/XqNJ7z9viaeAj8X4hnBr6f7E5ljfGxNLxObOScGoBmnPtWI79T82iZ
ImwsCHsSgIx169V7nzLlExVZJk2h/hWNrRQFyq48KXVtNoJoJC/QBsG7tLkFOa50
7zB1Cu8OCsRFWMXcua2A68MQzzKhIUfdNgBYwvldXk5LYCIG70qbYDBDFY2XjBsd
6EX8G6ZfFsidqLxXTqF3/I8xCsy9zuq3Seize1TP70sl2brAzSmz1mMrBi+bVomA
W7YL/9f0JARYtkSrBilZSMV2vDOpDTrjz1nV5YBVheSIQZDvssC/f7TPXrEVWEdJ
oI4HNF/2yV2eQ+CixXXnoYwOwmQhfjpxMFfPQwnpoqS/vLOf/mUkoucbmO8xBqzH
VtdSS/0k63f2UYlVmB90YeQZwjVeOKXonCciU6nW1cC2AJpPZOjN5XrlvCqanYXK
0pqKo8/1OuYg8RgFYSPp5Y0ErdA5Z4eg2QtpiicrDRk4wBlYHcDUXif1YwtB7qE4
U3DeR0/ClZnRUZuBQxY0+8CktBh92HyXnDxQVjAMzeZAG/unFJK42kPa2MWPrF9O
b7ryBdzZxwLq+BX9ALguU/HWOSPq6xIr1MoMKqdpRwdBk3u9jrFsBLEiNR+HxSsg
nJIAu+JQay7G2qrnHtVGWiTKZJXDvyZ5weQe90mapr1g2oZ+pp5Qcp+atSaSiYc0
DlJAsumWO1BYJbM9fcvmhpONuVS1YKokzUwlQ2efsubZT6TIrfurQuOqp6CmFLZ+
30DcVuiWU/AM71Y9f8Ck+vezLCLrqvjV9jGLv6gb69e8iXerCa7+tQsl/cCwDZLT
cfrwIaJqhd6+9Y4YmxhoqvtJ9Y92ZhH+wubRtpRreemM+i6b4P/W7AXEI+QvkNLC
0MPgFK4PxauT7pb+Gy94AH78lMqd9Vo4z6HW8SZ+3nBL7zrfJ6N6RLGEoCeWHwwP
ZrzYjSpOVu/Danm0I82aFF3aKhAl2TNmfQ38jp5ivuUtPj+BGJkcc3DizoeUPWZD
EyLsJunG6bPV9ZJyFw2mIUwjnEP+v0clyf72FO4L1rVgRhoPCZgyPrOAbiZszA0e
agYFCL3aJUGqUy31oS8IA3LDkUMAasjWXZ1c0L9W948fGsqBE3JxkCW5R3AQYTew
xYshXZVwhZS4OfigIQBNSfB3+iaHYHvPAHI9/Tu8z/WNaHmUPbqgDuqtu84ERFin
TJTMM8lnijpZueVaoDepTnZ3V7d5kRTuaSuPy1qiobXT2IdQufAcdnJv/LZEw8xj
uuIT95RzJq8pqiqUyvemP7rudtBYpB91HPf4WwblWXSF3NvLmEWFBFq/Z/37IwB4
2MnqwHzXZeNqQuGk0NbNf3NiID9f1kPFPrpQALoDoBDqt7VAyhhvfbrXUkbJmFeg
udBUOOc/bvB16hln+1Cu9zGrKVliqwaikFIUFIJdACfr7G85ixxCfxTkavJzgJxZ
ffEFKg5CnSt/D2tX2F9B+VHC6dNrZnyAAchDGlq0BvFwrEpat1/DkdOKA8zK/rem
BSmVgGnZ4K7iu0N9VSVxUN8hWewlC8qOeCFSwlqts0Yr3/sy62vE2JtfDjQg9NKw
yzTphwWbR8zkVeugJQ59nSan791skSE928BEOWSNzCSuPFsRKhLJaErl6j+NNYtw
v2sRi7befuR13QrPHefsw2XoJQiGAPuRIgylgYoqf1LhCYpIDrwxflFpwV8YwIVB
g1amUrB2tW95xFsOW6ugoURN4kObkMWPDwJR7JphspoE6fG19cLxOgv6u2N/DEzn
PA5Is5/iBePNwwpl2opqfYfdaNmCE2YYETD5EJgoWTYA1aae+c2J3yMehHHVaFFM
hr4dK4lNvY84ayBvLk/GrJ5F/U29qGWRuCwCYeX3gwzWG7K6YHGhb0wjQRBqU1Ah
awO5KazPnyDLsDGrenS0PHf1jtWw45h/pA2O6SGXqHDLkbLInYdbruNdTTBK2Adg
lY/9XiXm/tiXbM6sMf/iDT0237JKJIqaVPG2hyxthfcoQhdh6OXdLlJz3TOY7HDc
OzphLEcZm76W7qrchtbEMZck48oNeDWzGuDUzsL8RxKiETHdrJhlfuvdp3r4426K
r3/JTcakOEcjpDgTu1L1tQLtM4Svw0To85DVucAoP9mG4XTqhBmkYSFl8yi3fOfl
aQiejMEQ1uz5TxZn3GnSMA/vgf221avRcQx6xJzo6h48RebMjfVicbPOQizuWJc0
mcnfqsvJfHPaNiUNYXa76p6FXflM2XMBsX59JKq9D4ZM0wE1x0CANW/vl/402MzM
RX6XYClf8EFfitrXOZ+st630UesIcOCizIJqK4u2vCD4mU/CnTHBUSIKXjEUvNtS
lT8HgdoGwn5zI+agIPJNuFfT8HvNPqqdD4nPKywDFzC0Io101RDSFTfC18SgV9fi
myEufxc0zZlyWSEJ8cOXvjBQ9rS+8xNTqdJJ3Ard1zPitS1dIVRRW7DK19rTObz2
sW8AtxhSUpsVUyQVXY2d3vH4LbPJ1MdgOxzUkuMpNESPxI/IiLlDqIDf/ygMhqgp
e4HX3i5Gy2RQgrQ6YAuWBJrZ99QAxvXbf978so+YCq5YTJ+qj9iqQCogdmn1TWcC
veq2vnOYF+LTzFjITngQwK2KDmg4NoHsW4BGiwscACZTkabFfIw3Ege5FeOoYU+G
lrE9lBvQ3Q494k78Cl+5YUpHugWVniO5x2TLqQx1Qx9n03HjkGA4tzOxZR+9hhBF
rpR+Ww89npuMeav83BEOXgbnGZzeg7SeEMDjmeyNms+f7EvJIIeRr98SKLhdJgSE
BAbq7h6wZYvw6A5G8vnS/1PFk15r+GoiVrJDrVwIWPuCEW1DfL7GcRsPY9RjbuEj
LjxwZhxtkCvVQ458pVglaF5igFfrUfc7leANukMh6ekJ0F+3/qQM4Dnm1ddphGc5
3zHin7KT2KoWBbwYBoKUAYD30KufgapbyF09PMKyVOEXwFcLLsb9aipHa1Lib710
SPF0VBqqwNkVsL1mz6ZkIr1CQlCHVRX3Ogx7aOniwS+xQ23mTt1uwCGy4ujaB+VB
KiOtr0tJ2GVmd5WiMtVyslbmNHVVfxpn3CnOPTp/mSJTCAl9LpDvcuAiCIj1Rn5t
yTijnJWI0tsYz0cm9hk429BBHDx/ckxF5OdyEMcH6wh/yEzIvlyohySKhUfBKsLy
bMsgHkp4H+2w9i+t7wDepvJ5A0LRKxCLHJ09wYggfVY0PNUWA+1ALjNZOSG+Na80
DhZ7KrU3Ufnk8QJ0jqh3S+O47usVGoUhDRpmuBrGhk9S7E/5LWy/RAWCwJAX9QGP
brv02fRBPijxwRqWbwG5oZXhoKySE13hl3KT9askvuBohrLL630g76nuo8fQUsNk
agyP9348JgcNqQDm7/RsEVuzWWErvlsYJWAGExqCJSbTe5iUcwq9Mqi126tiNYcC
QfJxlVi6hYy3Ca8kUvxuCtrb+oPLE4Kg9f+Z/6lXB0N2juxYe2oHGxegsWh2VLkN
r8uVPNG3KIMpbbAtI9Q7qWze8puMiWLXlxRKwwoHhuiVUr6Ne6Fj4xi7YLh2csai
P41ZapLZX38gJ7U8DITJ2RBO0W1mE3CcYX2oaevfiIkee69Q7r5X7A5u3xZpyOG4
3cfJKU53BsKzknE4n+WkPm1y6whM5YVo2xTkjEuRu+nB+h3RLfH2bRj8R7Isogzi
Ofr9rDQtMoAOdsuv/6vUR3ib4hjX+pllGSVGxydbuNMbauyyWWnQkB30v2JErPxf
lK42Km3KMhDPKEt+AezFKJcUJvLH6D4Lb/wX1hMPnfLaFdKxCF/0SuCB+g7blDDz
wl9AMPz0R+W3X+C4/U0I3rHK9mtDq29gg/G+CobG5YJUBFpfjphL3KIgepEfqRgI
BqdY2yewG87U8oPgQp5rnltInHazszNAejyfVoMbvG2w5Zb+AuXpRJCKf4H510iF
/sxdjjwRl2v5YgimWnHUpXP6ckNUj2d+WQcwhJbfjZ38fn/8v5cgXj/a0kX1BViI
hoYQfK9FT3kb/teKhaIDDHoFoZjsx+j21+dTwUKv1pSujj+2X4MRD05TyR9RyfBv
vau1F/iIeSnVWo0MkMucidCe2pwm2PGGH7rRcazuvraL1vf2l4D3BBwovXeAdThT
xQH5Rh6s7fM4WdF/7vnEaJgwjqunjIBjgWoZ34/6OxM15Gnyn2LNaXluoNYCGXkn
dkQtgh9KvRpcE1wdGahPpNN92njnSJfzaTq2VuH04+gC4l/lWq14WY+81qYpECX0
Nh9E8Yh0aojET4lnLwxDT3idFmbnexlCHShU0eOfsUQ6qqiut7vW8LF9btG205zb
G0oH/hKEExcwem59aqGhmuy19XGpkJrS/UrWZ3/hqu+/JdghPeqJaAakJPD8ENr8
43nN05BhNWRFAn8VI+Ma75uLYyqIuEnZEPjhZg8SB2xdZ+8vHXCTI4XP53R1dmZD
KLnvEoM3SHcld8dkg7Qe9iycDYZ50PQEwxTNwuFIf93QdtaKM5M3DrsLET0mN8L6
LMikvIzfOt1Nyp30doUznTZgNsJhf320WQOrPGIajNpq8CJEwrBhZAKfaQsPeqXr
bWJH3GW1RFQucnrB8FJZZuw4TB5sHGJjGA9RHIK1Y1GJt/XR9VfjnaAiMQy22l3X
oR6kPToeE3gf/x3mGr/5guR2PbsBSRdqUcuL45i+hfcy3a4w5XmxfRVG/9ghYKR5
jcPFEtsBQx2Pjnz4NiwLmfZlnCFG1yEFkFwhWEX8cH0j17OVUzO+pwDzouNcMxVa
nZ9oQukzeWUL+oqpSU62DC+VhFHEKW2BO9YkqUSKRTUwyHwZJHURosPsAchBr0zv
MnQAEFmkSTYRU1sv3He/5NYHWNmC1G3+CNry7quEMOCSJd+YTLtVO90Lw2ML+EOH
tI7fySlRxxqoqvnRfy7TlzG6FzC539EKMXqhx8DB99UzeJ78FNujFEO3LI7o1uzl
BaMw1OIJMg61fGsMxtoAkmdia9xpb7dDgUgcfg+23i1gy0kuzKolD3JRdV6Bk9Dz
sUJRSIgf4PmYcAzm/Aquf+kd3cuC4guvIA9GXY7X6hOt9YGwYkQoZkBSQDuxoEN+
3rBfbo/LjUJJQkY6GU+zKnXUcuGukEfDPdYeYEz+FdSgiHhTHVEbu72SjcNoSJNh
qHhtMUFWgoqx5zL4j6SpNia5iKerkbNTHXS6eXArxPdpclPwJKdbj+5vPTsTJ4Ye
3NXfnAgarwP8oLL7Y9fbCWHlY6AX+RcqQaqJxFnjRjDij5C2KwZ64QT9vMTKL/w4
wso29jqKWW2T2IYAKj4vDxfPmFT0Rw5IH+xP+Bja9gEgTW8ZiJa6ZZjb22lTpUre
jdU5ueALiJrxGlrFiAAKNSiaLH/zKppwwnVrpwBzsuNedABRMEXi8+s4H6lq8xPO
zkf+7HCpxrXWTEkfqJaManF34l3ar+5HxOCDBQnqShrHmU/KFtqYYatN7c6omyM4
2Hj9iL586sgtvSYdnGMYMSfmifu30ushV6r5t9B54x11h1nLfE52DRWM/Su4aGVK
y9uiFfCfhIKUBmDfiruMybzBVDPOeufuvtzkSwUVQeAODwIILBP3KiSZrinVw+dX
3MjpkG/wskuEaADtAN7NXg78BX/O3HOlh3+JvLXQMD3oLTMNFxd4fYYrIqi9hY3w
eKphm3G+r0U7K+y9W9rlCwKFAJJ8zxyYOv7EhXL4W8n+XrkTY75GIRbqdN3nCVQK
kB3whP4t/61aG7GKAD7Dm7wIZXEHfHlIZaTURaFaEHldrwPmCMgO1Hjqe/QvALF7
Wvx1wPo4S1lQGj0Pmb9hMNbYGZUy5H2oWqkk/NiwgDE5f0vyTLQX7AGiDiXK48rf
WV2VMu5cssZ1WgoQl7n4WYyXUb2fd0q56r6STnNKuezS1LqSL9+8VAfXtt5CDlZX
Dz96GvxbGKGnXjkTcEevu+gAe+t4W28uSUUNvNX9jxEL93gcYs8ZUAwN+v8kvDBx
WicvlXINMooZ1WmtiTrzWSgyZQBx1C4r9GgFuTg+zUh7HkILnYK/5RcsHKTeb0gf
c1gKOQp1vkNoASZ6ZEHC0Rb9ft+ITleFtrJWHcpR2TRs3zonhk63nDHJJegNsxt5
5Sr7Ow2TuPal0ana1lomkO8FfG18FLQVKAILqt0vj1djaMPI2ZQrCR2e9kAYjrb8
ENC45DJyr5atTr3zWZLwa+mCAO01VuLnWyoyXqsNuRiLI8vYgTJg7megqOHm6CPI
37WY6ZTG1o1l6CBVd1tl95c2wLAQTwvpl0YnFUZFaHyMlBWiwybYAkd6WzV2yrmb
OW1VHmBwwyVnFUVvYK6ksMLIDv3gG6hNhyawkRxDN99WsWVYodMG7TLdfbl5J9z9
/J+MOf4WlA15m2siFUIXC2J0gRDqCHQe6dVucQCCi/5p/ogXewhYHXJBDQEEdsZ5
z4CLq0/6/gyUBS8asDmcUHnSrh5EtfXLAUiU0AjaM4l7zKMTOxwivE7tIyD2tRnw
pgCWtjawycFmaTyz1v7u72RAJ9aPkdnG3tjYqw73LFzffxv+CLpQWNnFOZ/R0tMC
nk9AczkSB5+OqZRM+L3bslMRgxnv15iYO0gY/5ehZJVVgpJJD2WHYZyIYe/N6X01
xgIwEgTtRY0DUvYBuJ3yYQY3KBhLEOtbemffPJ4thdsapxu+VI+TtaB1sYGMUfz6
6o0ScgKZsLZMQorxl9p16DLLm7ziXPx4DE5bwBO0XACCUkOkStUPanGa952liOxY
FcI2Gkg2HWQMKbv9nWs8E+yRI3uc4KjxSpcbnj6tTv+1LutDTdxIB5fwMKWZOT4K
m1eql4r/AVl94VB9/yz19P4h8ePTZe80+0UIAbxiUESsVRKz09eNinbghqdm+HrU
MzLFCTxo5G6gkExs9XaYvpvWD1DeWfC/GCGX0/sX11MjxykuJP3EmKI/9Nc8mWdE
NlypxxNDaohDK5ck44GLG+yjnzUCyRjmTVu5vJLbWkMbTHuCTEzu6YFFtUkrRq4y
XWbqOe25pzy7kCXCP7bhZyPD6lBfa4gKrHVVD8YE2uugSSDzk1HYSCIoHu9f3LGd
roJSppzqMbCVe01Smkm8Nch1OkD6JwsklAWEn7ApsVJ6O5RDrU/gKV88M0m+jhfB
9RsGUVGYBj7A9sqrdHeFXvkfOfkln7rUI/Yam6tLPXnmSrjoHzbhtEYy6g5/oqik
nx2ND3G57Mdd9+qx+wv2+5+et8DjNOJw/cciyXZybbcs155e07Mnk5z1a90shS/C
FN6EojJsyuwtYZbUKSnbSb+YjcR1iF1bM4yMXtkHIW6vMnlkJAN8xFyY81a0ndt6
7fWNQXyTKDaNxz+V5jWTiwYkgUDLi1aBELIIvslU90xMP4YSSw6zyxGpN6CdQGSz
uBHYCPSBvaou6nyz9ZrdBLFbsqGP+V3JjoqARTM4J6V0OvkhuE7+X+H4QqeFb2x0
vfb3yf38HlLB/YHkxZryQep2tJaZPIbpHAZb4FpE17/0kRzBYNJ22HMYW88MuqMs
obXwVJ501+wHNM70LGT+dzN+Wh8VslqtQdVUvmcQLdulN9MmScZ3tAqeY1UmG37b
W84UJYR5twOmsgbB6iJOf8uWcFOEadBnUHjw3d0Kk9yKpc6myM+nIBmkXYVsvGuC
f/wC12ArVyPyNc5oumXTtnoB5qVyzkEPK5e5tTloRM62fYV5a36BRT2Ixh3r4Rt0
d7kpEJoWs0va33BxLx29pAx0zMtE/y96YSwk2R3x1pJvZ2OUcmdOcoZ1lhxpZ8PC
Elp3DoIUMWE+8V6Mm5z2+RApKX91qJ3Lj5NbUTIFweQiTpKelxiHumM9XJdvQPw/
qY4XVmBRxuEZDh1tWBmQJ7tW5ZXbLTfunL7UFj9PYiKE2Y2mr8fe8zeVsVoTPMfw
CJi1nLnLAbCfdoX2R6DfwSoszxXA2kZixS+DP4YB2B53CaTEHeaQCqShtlyi/f7d
3ITpuVGcdF4vck5uReRZDKpA7o3GpcVpJ+nrL3jezRw/q3il/E+Rt7FlBoMk2IQ3
uMLWR/oaJPPtdNNtz2NVYUlFSO64cRwby+UqY6DY20llHp2WYWxitaLWEVTILrHZ
F3Emrgk7j/bXGwOIEiPGevECsQqUONuYHLODVE9volowkvdDKTgyNHEvn3LjANM2
/n8AVeHrEykBGRPVi28+RFFZtCB7/nmy5/GuBQVg/WK7grHkZwDQn18cBYJHF2Ae
bKWzw0Ya0PxblAdBS86DtPyGjRck9kPK+SlJVSJC8ya1JsoEQC7A827y0i0vJuu6
iPrgp/ZZMbxIANX04wJRhoE2aeH7hg66IdV86l9CVhRwieW0TkOWCWfahspeTodQ
SCm+lGfwq/om/cZzEdW7v2w6t3cIbqxEKOGsIsRld8noqHYK7dtwORDBw+rPEoiP
pQNVSP3OrA/+CqUxIMPtwgsjsmdjNpF6AEMPmagLdjPrfNfya4p+BdQCUoXKcWmf
9vf5WOOxpZEsmjMx9DGFXEX3gAHtMCEsczR+15o1L/zlw0tPOwPucEJAb96F3xnF
XQ2efQ7AA2ZRLnOeIntVyb0j+WeuXDFcDtml/qrsvtXykJ6H+qbcDtc4FekqEvQi
BvsAeOcnzaf8lxdhh+8IRvlvFstPPWT+nPrB+dKpYApNrQlqwMz+JBML0A76/Aql
Z2G1ukZ/FL+JCbPlxD/3XYS8pvJCyiLeJsf7yxSkBe8S+9K8jWv3FjzdN+Xs+qr+
javYDw4VLeH7Armh4nbMD5Pg1Qecr4M/KVhXexUFxgSU5JQsYMvQZJYbH59Zul87
SZvmF3AGIT/Wj/fMRGMyGCAX/YBttgNXJHVOoFowHGt5JBDyX8QQreReUYEd2ixz
cdGeAtPPoUkapvcz5jgXObxwxbxyvmp6PJsCTx7jeodN4z7tarSpCrUM6S5m0WjD
KsDW25Izw+Ai1sEOfm3LCqtI6htE3ml/62rWVPJqSkuXu2UOPou2hrccwZ5NPHjD
JAjvna8UL3DDPBswix+fkfepVZL2vOxXLv5aIIkM1PLgyqTdhCez444cvfCj3pxX
W1b7SZx/JYzMA5a0Z0MDE7lCem+W3h8hVJgd2vPH1qvEQM9EkLICzIGBavPJ1e+5
ZKIGaJeJUasOlOxMPjDy4HHBeGWsL+IaK1FQjBdOR8TmgvdGnDZ/yJ9MOQpwWIo5
f9wp0J6jkeuJdGMoJB6Nmirrqsqh1bevBgMDbLKYOct106C0vGCx3qPClfExLSbo
84POJ//nt1iqfVCzfI5yMMB8edkVN3i9JbbG4e5/pCWB5lm0ApbQFEzbOk2LlbRM
0ffXtoEmmWNNBNk+Jkn4ehojWglA2ioDw/f3/FZntXd7tboSnwwZpgfBjBqXM8fx
IVJmf1ngx5baBlJb+va4FDl7im8paEExqyMLJeUaH9LJuJDjm8MUhS7JlNwUU4JU
RVI5NJHxJ/vW+aFPyVVG/HPE1/0BQDT16pZexMDMGNWpH2ZjRkqSE4aO3aYfv7cb
MlNLDk77FHuT9xqAa7rqysSplkZJNSpwXZMQd92OL8DueeHWJzRtfiq0OBiDD0EQ
cF0hCHQPiUm+0ydZzP5Lqf0QG813J8aeSBbn3RqoEm6+ntw59JupQQPUX3vfsS/M
hsU87z2eHjCl1BHiVK0SANXU9lLrMAo9rVQsLkzUAWUDf8oqtoibee+qQeqf+Gdj
F0StJ/lzqMC6ZIZH6GW5bcU9mP7RMqGqJ9PD9BbM6ynNvZuihXINkQctlnqQpc6m
cvI5c03AxsU5hbnhb5sulc7JVFsBshikOn82sE9AK4yOI+pi/6U329I+oXQ7yX81
6BYmbYFq7X7vAIJ+xWN0UYrmtAl0THSJxHtcTE9lKg+hGpwL7qhbr1kzWllaJYuh
aD+SaTBQvuiXONuX054rmBfJ9Hs5NJaukBZVdacy08/9+5Nrde4FF40E9mP9FFnr
Wj19XazdK81qSkfNR7T4Wi4t2iTxbAucD3duzZNSSde/gBfFUwJd2EryDLX2O7eP
aPFAGQQ84vSOiDL5kVPd09elnEpcFcpOeb6FcxWZfvjHLodBx5ZPBQNmZ3FWO0tI
o4EFI77W+FcFF4XDUfUK4vmB9cjBPUBnI/ovqLfAnUUnjcG/xJb6MW4LX/zNTKbK
8gABJoqtwuLBjkwta5frLEPjYsEdrRL5zcAiBw/6ZdsmI9psgeOjBZAQBz9BCp7P
l9E6sZbXZRcgFAfBuycHmo+KLQluQy4viuFZo3cYVIsg5hb1mFWxpXpe+15/Onuu
bcaHxrjFMLB71RWSOsob7NYFEEqGop64Z5yrajWfOjrYeA0olcTh5ENXBiA7YsQo
jmsljIh7pY96r3RPLs0E7tU8Xh0l7ctEYrg3sFjB+P69W3MzuXfRfT5Y1uF+ufSo
XYOJXopwC6MrQWXvHGVaPE3yF8pxWBkp7XgvfrbeC5oJ8l1hnbSKGmBh2o7h6+5e
IkGZIXUxpEsY0uFPaWpageq/0/vcMDReoQzA346AROUDUNeeVff2EXV+X+M2ragN
CyrVDWAPfbjWH5+VjpS+BysdCHMq4ezamuOqzvJTwvgqlXiuNwcs4vvXrutXDn1M
v2Tht5TDCo/Dobov+O6ObLFJMbaaSyghFPhLTN/pzkP4ppiYXcl8ZMzFi9q8HDO7
B3kTbUsaRe5d9yetBFZiiF0nY6y4ujDEI//EF2eC8orUqTFLO/XGj4fmkemZKfll
b7sudd2JKCJva4Z0lMucL2uXgnmFTPybIh8MODeCQGfRjGdUUMtF/7BwDhwXeot4
o5Lmby1FP2s7jx9ej32YSDh11woHy6wZuesdVpFZC0+H6N/XyubWNHtNQWP//4Mt
fKOOXGa06IIKKuuIm5M3lniACKrldSxRGw//V7raHCyqFYncFhQGxrhV+hoKyaDq
oQTj/Tn2YyJ6dj/IubVTpVimODZAAi89QSTj+MZQRfxze9XyCt7HI8fDSJeyfGFi
+G+Va4CbCMBuLh0yNDoK8oUg6fUfUQjIRQmsDo0XmH8DWcdpqgUQcuEUnx7/JC7w
CeDF4FOmpmV4qq12FxLCBRx5FZjyVynq3ZoDMc1s5H9wNfE9EqobMwGgk9pwEtcZ
UDDajB3PiK4mHWOj5vjYs+W0GPaS2wR82noS8D9mJP/VjY22g1Kny3H6xC+f6vz1
lWQUhX6FwjZdNjQRjIeMqpP4IP9BxMYDZhV59POk/r92tm1uvyO4wjwUGyru2OVA
zZgO/j/7dKhxpWbRqOLwBr2sJyFbQqQO1JJAHlxsjgCoT4F6RjUYUI1I08XmFBi7
0nbAr+8k2umkt9lpU6lLmS9uZGeWn7m+sEgOetOs3pNiiiQtnS3XkZtop24iPD9H
FOGH5hmqbnjp7JJvbMgrCL2jCpqa9YbgB+oAaABN2WkvDwlZ0LPLhhRyHkARWQ4V
eHPI3Pgoc58NqsZPUdJvXAzt1Ra5DG7kruyXyevRuAakSI0H++LDraAb4Z12QYm1
+fOjlfttEEq8gFTevVBK4F4yS0p0VcvmHJXRiZte30hcMnYEvyy6/Fq0JFJgCzpp
CmN3MZ3ghcu3zGeKAPlfl/AnogmPjZz+eRVFF0j/Z3IQy7QPIPLN47z2nMpbGgwj
lCXtEX2erpIo7zyT/tC0G19hSTFJ3pWCS0VoJg8Ql98x6uZRZEshkYM4KeguxuE3
pf+Y4nyUdXCwtBPmOyt+9WWY10dJc+zPs1b0yq3FFgHRibXWOi4Rmcy/JI1lAgx4
MCsZEENmTCIxjdzKL2Tf38e4jqqnVOLGkDUVHUHpa3WDNl0v7LeMKV/c2sdc5fd0
TLTuceZUVYedOlwSntHItAeuhL8LI1aB2zrTqlA9G9Kxr3OjIWwZJtyvg1iUcI8H
52dW7Ox9C4kYTKLVzVBaSOkiywIfzZ+w35kk3ZplXTIggt1u3nb7DlO59D0xQjPo
z8lyAIbdHLfUzMleabHraFV34YvGLezp00/KkmUIGoDjw++N8mK9lbBALEC10nCO
crPgCb3Mxv0hjnO7dj5AjVc1a4+xQ/C++obB5PT8PY0ja5v1rkDVKsw6JZdmmxz6
1ei4o2nE4SCjL2qpCQCFTmwOYmK8nnFxT0s6tTdPnaXRmA0ckg7HsbNJo56MlHKL
sdWk2VDv0TmMue5NN+PxcusqGKGJpQjhC4vsoE1+r+Xo5rstBZ3KG/cFSnPZ4w/0
sv4MQVRF18bSRK1nbj36oe4D34uELEkwU8+7DXEDCEu685ITnRuhJ/csP0NrtSf7
ga+Mi8FD01yi3vVqvjYzqa6EzDP2cmgXzARfGSjWCfWdWILFnTPrxYbuvOesq+hM
BRegPZPedleA1yW4oE91h1dz4W2vG2ayRpsqR5vBfJaODZoI6lZxXPronR8fNI2g
EK8BqgcKah1QUDhcqiJfPsWCuPRoVu2ckKBnShtf2+lzsboU5pZzYdLPUkrEOFJe
ILtgn/Jo9gAffIuWOgWipIKoDT7kgdeaJ/N/wiVeDpFZK3tIC3+WiS9rpRIOdRIU
7yNfyfNdw0RshqlBqx09t+TajdXlsHB4b21NK4T9vE1L5PpFURDKXfPdXAZ+W3OO
z/3eh6dViUOt/3G04Sw9Yioijec++F3sqemW+EPrzgLTnNInKgwTg3oXVpvAtMRn
SSaA5SIT591sAbfbBFGlu7eZSg+zm9IPY2IFq3EPlTC+pKIMC4mgn36rBHcG1O0i
lG+wLrn4Cnz567VC56xhnfr0v1pY+Ilj5xF+uirXAiHQg91tvxheYQHuU5n4Hz5I
ahv7/F0opvhnyCW3+2vDWX234muvkhmxyiuFLJ4O58DBy5CLogGMfb9lH9gTRYq0
WM4BMjEpnrfgy6MprXsnzCK/ccbjSYRpaMCQAKkabareDoV1FmxLyfnG2rxIQ/ts
7LqYOc8/73IJpIszu8GWPb53KJnBk8PR7F/oYdlgWvyRgkt5YjYkQccNEcoXVQZA
SixD/xQX9jxcfmMDXQYcBxY6l/UsBmJ/2C+gK1s8kr12digbrkfwYPV4Ry9nozyf
Q73TDWnpHaymquDY7A+dRqW+OPOXJCYg9/c7lrttS77fOJILPxavhwXYjdeQeZPx
j/4GvveDcV/5tLdRVJx5t0xOoJyivg76jsVcodsqS/5fQhuO54qLFy5wxj8DoOSf
02PcvDhHxi3uoUstwVD8fw70T38CvhVvmyirmFlCkPeLTMiqGBVfhGfNGd25bObu
0FohTatbK+rbK3oNKlPm0cMHK1QiTzs6H7jF/Dz0XaL7rPzauIU5zwQV6O9mEdAW
pRxtWZeUEueqXmZgrIPs4DnRQT4U1XPwXKgryisol5XUJ9nkFsw2n6OHjJDwQv/6
EVAtp7xOcvDSOiknL8/DRALwZKvyKkMSekbTtAveeOMIX4ap+79z8XNa/YDzKpSZ
F/QYN5XKpOfkq2yhIxzfXEUZWWs1NGS5qgTrS+bzCYv0VQppA6uPdB81N5/y1dvd
otXbQABekuYEkJG9ppP8ZnT9YmaY4/Fo0Kup9Gy1Q88qZNTGVh5QovartRzYD5+W
wst5AC4PGHmrSClliW1L/q/PCgVHy2emX/lu6pVPZZ2JxicW4yKihJwET/lfve8C
ZUwCFeIzHnwu2NgCEWF8+d4fYjD5BBWasXhy/FrSA5k+7eBQbVW2O38kGp1mdL2r
iIJo7q7Pi01DsbignXiLWGfsbFHmcAkswusb4WqbDLVfXimA+UbmJttuLo/Kgk5/
qYfWZWnl6vewNnf/Rp6KuccjhlKHBbEqClqHBCOfUn2Y8Djg6beAN6o4JtJo2+gk
+H5YC3hmZwbLPKREWfWgW6lr15/loHDehpMz4MU3Np3zQIp7/GCnhrdje9iGEtex
+E+nfNDktC9LBRxtJHuCuZ26x7kJLJsASlaRoqy4ZpQ59+bjJTLXg6EUDz9WpJsy
3DajTMmZTnUoiojcxXEjix2IfpZG9I/MBUH7f39qbZiYs8WJu25GsdT2WtUU4keA
1Jes61BWPBF7R1H/rcGeRNm33CT+NghK832BkGKiRodcM0qVgFjf703lRD2/sE5f
fL4MmJnw6ZIeTGNEPbvh72sDpwqS7KxhkJaBrC8bHTtIl4ps5Yef8dREXDPcVuKF
tUC5CpIkYrdx5MmYnrvTBtfWLNxObXuerVlyLUp07SQtWWy2GQ4TCJELhy6hrw/w
8tY+7PnEsoikQraw/t0m2FYIVmu85iXwplEQBcT50psBjuQYMJUQWinYjDLcBnGh
4+iwMWnYee2Ucu7eohAPU0P3cEziK5kBjFnAXsAA92KHAsGqAztjxsvycN+IxTtx
Qhnh79J/k+b9QoxBv9ykU/uEk+0odNh39fewH0yJXhbwPGvJwQvPakWg4MF5pxRZ
jTAPkJsP17J94jwQy6hQinaUbTGyGITj0AfUQ+74rNL9YLZpYvS9FofncblbUDnr
M35cbh9s6CdBzBFE/3uuULbZ4OsEMRMcvxmOjCR4OgPn1SbJgeRN24qeZkfh0LsE
9BVJ/osWM3/EhVpi8ACYfQDsXo9aMzaUz/Mtig7CoXe73eNPoYS0u8tiP7eBjnYg
IETFYw1YkBeqgpAokdSFCTUO0+HbqdMlyCxGyzEjcq3eGzfxxLOI5VRGwvNJVB4J
SLVS/9mDw5dlc7Nwgo5WTGHKWd2m01Z5sXYHLeFsDlXRjZGNu276EXda1xg2g/Wk
0j1gEEayH0QrPmMV2aB+9wdRdCWUXc5+gIznEAMkifDtImMmit3p6s0v/GgzZ/gT
EiwM1GaJSQqCY16xLkqP37yfB2KgAupllAcyrHohBpe178uZmHElKQePgtCisaGj
TiNX6Lj+qTTEiZzMhnqomsqQjyHtheUJyqnkqamPg9GKMWVsEqfP+AMkrW7G48I8
DbGj8tOKlkSx/3Kom6a1iT+0GQF7UZ+aJzyTaHKCpdLRS85lG4zcqR35ij67VNIf
zxd1PF5zL0tYAmJSkuOlpyrCGWXIF5CMQ0esEJREvL2+Rwf+a2A9RT4pTQLr1WPK
QyZBBzqvjpyKKpgpyZKQb17NILJ5Fd1VS2ycWWLjJKvj98ktRYECjAeM9EaXQg4U
rl+YcMW3o6/naO4Xa/hHhdpt2PTRofJPEpiK42ZLeL5UrJl8FFDF2iE7JlkwSWSu
RSw9duVVOpL5MGVfKOYlFw8SJrHJR0/LFEqBm5nknF6RzPhDbJZae79hSj+3HyCc
c38LRPsT3YxAxj1hqRFBnGF+MzsRNZ7o+SGP7G47zW9NM+1QnIFOZzSUvN39x1oj
OhVJgTx0ujomZa+4tgn6QCjNNXAQY8Rx2WsIL2k+xpi1R/ah85N5ht+LfUNoLAVC
wJlrxzs8I2SkzOmB92hzLQqNDMXHx/kuEyb1xSHzcsHrgZ5RtXRrC1zbjiFkldeN
0FOOP52VSBg8kXoXXMHXwGVz5Xj6ArBlw9+Yvp1LQgsAFkGDmyfTeEojbUS6eCmI
OrM8/mwD5Hha39r+qDVcWu2slzOfgJ8sQcYjI0nrB4xUpzjlBwpgnzgBUEqhrYE6
3PWew1Ge4soI1EE1H7q/82C2AV8Pygfs5KGyRJfxZhECuILQteEWAsFj3/aY8YSt
O5sel5Gv+LA2W2TZiv015m2I2XQluC4iWPAWbZ/GEt3ujzd/wJrTNSxpu1ZJMbu3
KOMbX5D+3bZEcuzYSnc1bMEdakSoBbBxgluTBrtKWu00ldup0cv8KIDXiDK4pvwD
y3CbmgTVodEM6RZ/m/55jM/vNXDlCEVbRKXCDJN4yfnj8e3j4kG8qyvJCI+TrOQz
+PtzeL7YUJ66EhzpzSKE6pD1jPzjlE85fdjsUQJxI42vjhn/ZEIEG145IekHAvyG
BE/j5dwSgHPmGOpEWzkPDj+FyFMZrP+fBh/o5mafY6wXGoGkRJNKRliMC4YjAsBV
rjxDK38ABhL9VpJa70SPzl8s7jsWotfJiV6rDcqMLETy8P7npNIdfnIdDzrbn9gI
jNWc4G4IgSsVsaG8N0OkbLqYH7l3tYeQ7jnkfarEd7nAZWi3h0/ZoWkwya9E9IqJ
HR1WWz++ozREvlgqRT5eDAkF5V9Uc2xvJZyxbOLH0AzMxrchEK4OuBPCSgfKBZpY
5z0vpHgXDo23LSxWAEImrpaZcqrLkoIZOCJmrPpzYU1ls7s3tuovCw57GQC+KSV0
n03iodDTJNL5bQcdoEFZWzVy4WUBKe7D+mOLVIrhuxsNMR6Fkw+zNHwO9yiTa/C9
yvsKUosEWxHdswk2Og/w+wArkXQoW/IszM9eaucihrxKMTxL2kbP/FDyvRWVd/oc
2TB3SmOJK8mQgV88ANTDOtLirG3PFOrcXQHio2mAJLag6Wf8yYQ+Y461XsZEh82I
W7NQ+Q8yDn91OJJ4Ax2p4bQd4khWei7J2zWNOdpVJiJ0+p3UWmsaaNElE36SGq1t
gFNC9XbuJcozLx+fhyFhvJFeMRoDAUhiSPUdAVuQeTU6jZgNu9wpH1fZ0bQABcso
elbtGY4VXE4njAHyfyG9nXblXe9y0Vim5A+jHjIqF88Kw2BHEnc1NeaTY6VrZi64
qgjw3VAYOmobgq1LxSP70evXMZbeiPinyQArruoXoFWLsMRzySEvfotWWMh2uk+N
AMTsU1WlvfaKdNxmalMJk6SF4GpkOTAa6nEEiv48lJW0xCKB6u73b3QJ3+4BHC98
wo59TXvjxIqGGkq3TBUwGvUGRO6bOMYWxlH/D+8+Y5CklxdUuyz9HHavof5Q5+n7
zy2r7EAp0gCAAMn40CDukppLnWBbVhqRWxpOSq08ApOBHBtENZj+x+hjA+O/duxW
8A6dPKMxjJPCf5dLotCR4WeyOsoBHnfCNRtZj7QHZj8I9vsePqYHkUXbjCjgB7iD
YeqR+EUVCTFddmTrKjZmTUbdRjCwYMMpGsDVjoeAIu4sV6IC58kCcLpKEMKWcfdl
ZFsrrUw/tGOgCgbtj3LNzXkclDpuNfBJSrJd3F8wxvKhF2N/74m4i+4TySl5dCKr
ZPYSx6iV34pNtRaqCyZMoMuEOtuuqv8NfrsQhOYbFLDV7hoArE3sDSXrAZvdHx6Q
CqbaiZwvFQ+2Gjih98b4t5JbrzAbMYxPdPuyObuNOEexIdCBK+WhkWc0bbY6lzMv
AS0OchsuMFVYXpi0Ut3OQjmqqmvatm8mzeO5PZg/yNIBvQVPcrzcGD/EzrladYjZ
TeyrHf/f+mDJuqV5www/WWzBR5CwkKjOO+K5t29zd80zSNOQlkWyjm3ivtlZifOH
03Izqp/6QQy7WFQLwWwN4LE2DG5LinGs+kxlk7YvzqVdxToc+zYhxvt0Nus10EH+
+O45z8JtNeBE3sg2gR2VUhy5QLWoC5Ld9njvkdTAwWhc8TMHJ2aqI//QvBE6l8lO
8SJZFVPybW/xjf9lB76n88pTYw1gnvK2BQt1VDXUOFQdX+MTL3kRmN+aOHlQLtRp
NQuqXYRgUSW53Of2nDtw2UlvnJNXZMQPIdpGPRCKNyPNMz9ssxsgxEUPe0iC/jaL
osrc5jviWWDjPXIswL0+Y+LOLCfyN6F/sekwICvXBKgXyXIBFoxpOFV3IaIHKOxi
KVrQ/pkgLRsvBzwdjzQjYuXJnYyPbxHn69apreSSS2KE31moHVRr+0sl47E9IUs5
8veYLtVD8fNfuyPbJHbeHp13Kqt7uEbFMqJB5tDlmHYXu1D/TGelaHt0wg6X060L
D2RwajN48RcPQbpOMAj1UoLjCDt8S5acDnMT3Vd1cf+3FL8BTdgu/Cm13KiTsNip
vPVj4mMxvLYSnbSZIhGSN+P+eV3yB5V6NzWD4lQoCqtkKGf4LEc0IzZNn6B0G2ON
gNr9GF3CHC+h0MeuVRfCB3qoS+gQpcTVcgUZBb7EpTr97cWfuZu2pIShkCvFUhnM
sJgiIZ1sPoZQ7k31pTHRT9ZdIBzF+7cjJPe3ZHLto+BpGe6w7xLUcnvZlMSc+gv+
/H0llds0C2kMV2vjF7dVS/7pOOMDXbTPS4NFScp25gZNIRsWhyWKfqOLEiL7afYu
LNGTB4XIpTQ+XTQks/iuFtyZltzYbQpwLERVZcxfODghxNfMeHVBlsMjK/H04BTP
/wadlooB1if2trDEMyfld646KzpRFDgx7KVYDoYY/k1UdwyoaWFYOVEZB5hSs5Xt
MxyOrUdQnSzE1+yTgWcQyb++/Al3FwX1NSxrZHMbsOEPvy9e9k6pJgJKGUliDSCv
nbbY0gYMSZC5RwUS5SMCA06hr8gIhwjC/n+Z9bZWLrbj9xiufyA1TRz151qUK7ri
YORVMxZ+Ca+st8OerHQnJPBrPOK0TTxgq1LiVbiCAWfM25PZRn9F5nZ9pRRYVcWi
KahcbW7jEaVTmoWNp4KMleGZ0IcRl9QQP2EeSa1wu5yOHKFH6ZnVVNv8dCsR1Xc4
ph0FiKZUB/dHe7R8hncSL8F3jh38u2vYWL+3/6RsQlJYuBBTwDlS5DI9106No71U
cA+QwnsqkzDSG45MrLH4HNabZUyne/tKjAggiX91jd8U1oqM4iJfpNgq3YWQffQN
yimCig21tCUCxuwpykrAbHeiMOXSxjuVmpxUN5wVM4w7f6vfF120JY20cP264dWY
ytRjm8GH9VhmT36CZVcF7d71bODrKQ6ZBEoK2JGPhKfEMKWYxjGIwQDGvChSR1pW
NKNWTeeplYf8Gj8KYxZhxit1bgbN3wMiN54/WdO0jQx2a2L/bEtw4FH65ETCCdax
hi2mV1xMyWnWRfXWDh5R4HQ+o4VwAZoOhPY6PwB4fVCqol6r4UCw65fGfG0/IPYs
bQAMnGeCJm+G0vEzZmZZ4XmPnlzjCbTWpPQlddOtRIoKpdg47rXA5t0un/DAazN8
6XPRSCUg82cHD/QsUhNd55djawmXRs8s/bsTdaqTWn/QE8twvhAeQlYp+Vl72mmC
CFcNRD9s4FqFzcdHY1MJuU1ESvlMnqzN+9Svsv4eQIZcfefvNnu/aj6PE2W0I0Dz
tNwtrqy3BJpnmjI1pXSzSf+fLkYbnp43N4VTzYrU7fVqgPqIiIgC3+a8bEImFOlo
KKnZJGAx7VjLiWRaTY19VNfnRDXcB4OPK79fJqggyobJECRXSSgXNAsKJAawEZ/q
mhATxmaAodc+cz1uP7S5XCpVvA3XE5abOC0R3/OXxx6UqbwJeF7/IaeZxnc3FFa7
eYbMdpGeWSkCyyYOyYng/M6E2bcvSclUx5UDd5oCZ82xUH21aRbkrsL3F2QVzhnp
at0OXqVMXgjQ3wSho6em4g2wN2RRJ9QBMT190voY8FF+FgHwJwmt9V+M4aPaoEgu
nuYjfvYUz90/EhYfm270ZLrYciHJE2cdf3qN5txoa8JYEaMwaWgNXYKqtLoCU+IK
UFqeERTaATs8Sc+xytGmki6/Bopd04moBBjGQAjzPMtXA0Lohq2t7xvpMbiBzqkk
CWeobKlQxoL+Gse3epFvgfhNZDsc9MmXr+UESCrMJDibdwffEMksK4uPLfAA9chK
zsDog/zrG05hbASfeAfnzt5GTyK9GkOaZn1dCOLG8vhnMN18LNYHZOFeSidUwzLb
Dl96C3XujX65Or17ig51WpMx7nShewJW8j1KIe9SyOe6Q7yz6mHiMRP6DLPLX0qp
Rq3bGfv+gq29OKwFG7URXGKgeBRAz72uuZDFqCWqB6wGpMf1QcoJiyeObek8BPBw
Y7DHaJM28dTMBK1BkPrBTeJUeerIK6SJGZ8p2V+7imi3PZqbY4pksRlHVeABIjB5
Yv+KS4g1mqIcM0SS0t+2ovz5n8/rV1k3hHXxeKOsnCC+DMeor5nCw77+US2JFDMj
LaSGd+/gZwZmzsONWnKJBikUFL24wmIXhCvLR5U8wyttO2RLOHQJCGGJAkXXoShx
AQtNjV0PwJrQl9m1rf10RZ3Ufm8COFO7wTrh72SiOyDDfm5Fqwv9Zh4PBpGvzFjb
A53ask3RHo3PXktMB6lrs3Yz8G/kvyFE/n0j7+Kofn95Q8rTDpdcuwcnJk+7DD0W
3vzlOP+e8L24luC3MyPqmyiQaJMg4S0Sqx3upDoK8fPZtylJmHiDJsNRaLRbNNEy
t/Ip6/Rx5913/hiU5tpRq1y9NKcDXoiJQnXdiVBj2+dmpbx0V2z0NZBq5U7kL0nf
HaiDI8PuDf/EMKCcrKL4RVeluTGjfxEpsOCWNNzFJYdk1cwWfQZuUXrolAiPoKy5
w8uu6VpS/dtsz+uVAiTPmS5BdS8aMdq7bqZuOKnm4U7f3XY+11QHQMyqchJ+/sqp
O4BMxPZGqKydeuMEvJ5pgSP9NVLLL4cJVuQHoIiA+WbTTFB/SfR64Q6seFpsP5kI
OCaZ+REgCEdfOtZmb39AfG9MY40IwqT/RINVgaA/Oe8YXdShIbMb4nyuxKaML655
XnoGrW737kw5T5dRLMtcmBekTEcdH64Jfw0hEEFyWkZmOBmYR5CYat5HRo3qE4CF
1KBU62wM5DBsGlznVjWKPeIiGME6noEKBPIassgP8SsbyfJDKuTLHvQZk1nUnHaw
FtjHBFlgf5P46YfmghW74mg0W/Jdmj0qlIVTBDlIlm5evb3/ruHs6dHbUiQdnIs4
w0cMdtZPnYJ8fQK/X5hYJFq50SXQv7jKUjS1rXYxD6xqKx1esLKj7TK1TGmep+Y+
oSBlkOzRMEb1pwi8FgvjgfbNTu9HyZO77H7EmeoeJWqzHkggAsFmcuTCwqPO/+x5
c7kYJh2WrkeKkteERsoRf91jGoPrLu0KQHawKRMBWfu43pi95769gwtUjL4yLd3/
7A4DBStbdK3P53sq0NSPUB+x4fwyfrN2e1wz/WU4yJwqb4BuvAFOjU6ZOdfB656A
E3nq56armFShwjMkQ70b7LFtZ6sIB9hsndcFjlqkEdK7QZZHCmhVwWQgB9w3KmKn
Tlo1qQpN1CKZ3lqyKXvJAbDnkt488v8oD49n1nS4lo+cyvjJYyUhuf+XxomDhgC8
M8HzUcATiedjXRRkD3mgUf1xEwVMB9/NbKag5Vx960evMCLQZjojDpr+N3xLFlyg
73VKMIToFSvlrSc6h/pX8M6129tfS7Zpv0kumGyaXE9RH/V7jd49yL77su6uRsiJ
NhmR49gcbP6xe7mKLiRtV9iDd+oExW3UiJ/61aXjc8+0Usv0DtFGnME9wFYIzMHd
eTEXQ1TuczbuTkjkaqIBfBSB/Wj5kA3pg4pdU5x8KBXkRQYiPpAbDGP8xgcjfb3w
68dWYY36ADBr5AKAss8jR1SjmmpgBi8Z7LZvplsVpPaZW9MG99Iw6uw0u2477uEC
g18Kl005ha+E2egOqTkR9z3ZeLy/WPicZEGOVBah2hbd2+WjBQxDMMVZQMEPdftj
AHfqcdO5v0ASJ849Z4BbhloYzDAuYUjrQO4/ifeEWzoaOtQ94+t5P0PXXUIW1+Pp
moa4XGmJ/0PHTtkxTa1E9GsVO/JSILQWUlQSQ2pUkwMNH4WkmF/VVZU4Uq/+GXim
vRZXvvnFCTD7iuvuad68mkBDfjSI8ZahL1zXs5G2R6StiaC4VjjWk5BtKeuj/KA1
xUDwQFJ9Kq/m2YYoSiTWy3frRnYLgP8hwvFclgO0WpXq5CYlap48Pb43Wc0HjDuM
A8ms87Q9DM9I0XWAbnd2Jm7HfRJA0WSV/hhmMGX7zX1HdjMmtDd28QLy8txHlQ1f
xpXyKEVf/ZbOLbMVr0TUtZZgpqAFQ2cZJzh3IFoRRgVLBxf4STLWVbgNsyWHALia
XQsL5a+gRZmCiVvdBgmirb5ybe5i89Gojdyc+kbzsCeZoT6UWlc37rW6fs6lGiYL
MMdmai8UUj9FRFMXd7iJm/glxqfaHTEF1FvqVOd7tLk6UKCaZ1emx9FeX7UskXfN
2Wj/ywazkBeh/xBN0iNT9+HZ0WZ9r6ne6SbyCTVZxbWLt/J70U2BubTEhf7Bhbul
TXwe4Vz8Fyma/h9DovUBryv7HnnTsmY2IUr1KvK/nBfWSx88PQXDVbxwki2SkZaT
xIvFbdl1GTW4WrWCDS8vtIo99A8BqZlG1EnaPxTr7Xz3x+s2xLLXdQdd9lJe0UkV
iwbYYwU8mKEzO7tj9F4nXL/uXUuF97ALeupjTSQEqPdJShSAyDPBFsTvkg86lvOj
xqgiBF3F7QDSwonD6s7jnrv9HmRguJwT3UOd9q6lLw7Y5gotwsxFz7C1wu6g6Eaq
u29mv4I0Cb8e+I9L8O2zXYUbkInrozTJn7H5FFLWS3SIrD7XbBjKAzp6xGXeAhdo
OwroNvw7u0IaWGNAaFOsNSC9fS9f3sEKIiUqm7OTxiPLU0J56eZ3YK3iatkQOT3Y
lM1DhqL6hTJfw4BbDzTg4jSXEGSFF4e3kLEu2pzQ7v9C/Cc39mBkU/ClriREGdWP
COGG+HAtW+sZi195XKChBqpDQEQ7fvt89JPNd2Vmkghnx9lcjFfXDys7scEDPntL
dVjcVHEcPRgk2RNFf1VpeR3F8ynm4rnSVOrjIWSuuBJVX1HtlcVigc3Edc2RNjcR
lBEdgeccliO4GRfLnhk4Bmz+u40Yslg3vycduB52BcDuXAXmOmnVPbxCflpv+HbC
hLA8LJf8AsrayeIkke21JjlpuSHRH4MAKJOrNZwIMmY1Mrsk/B2r+7AmUbwQ1T4G
gW9lUM77crLKoi81KTl787+hWf4Q8ukHyvlXHNFuLqzeOqvEiGbAF/vPXGtQT9WI
g87maAlV9OhzsRG9ydMNHkAHbwLfp5om03VzeX9C2BttpqS1ntm7LbhjAOlEKgj5
/DUVDJKxWR3rGayhvRA5Rd2lCq2BzqWYnlAAiBYlrHRUCUhaB6tkpDr/Z/wCYLE/
0Bl+udIVyBadNaQhDRQHemhc3oiHEbb+z/Y0nU2Q3Ga/N5AKuKSX4E64/DtMTG9C
bf2Nkv6XLZyo+IVYCJMZrlPs8KLXmkr2bp2FkZoWAS76ZIJ6dXTWatSDNfg0Z+D7
EmROM/vY+OlojXU7O+vylQbquxuPoZqTj+NB5e0iz820d1MujguDeteSEj+AMdQq
mS58vd1SJQzeA5TXMWnCazQMPWEBgSAtWS5dkjwU+hDCXLNwSbBSUrPGmgTUpIoL
cAmpc4LQP2e7BuvGjOkSzDFDC3uB6JhTWZctwFvlJo5aLDoj9Bb2hEUz30G1FMFy
Zmdf6dNp95UDsTuJ7QWKzQJS2GOjJVyiM7NvBhrBsE6hfE/BVd/2ZWF+mkYkrsFd
1eJHnXbwlhk5DDtPgrPIUSzxz12Dq4Ee+cH6gnlY16UtQuPIqSizWwCdxPlXVind
yAtU9fAjUneryyDDCwM09y6u6sCDlqTER87rfIOfOhg6bx82rUrz1jevEkdxknyt
maG21OXd825M74LczDo8X9Giho0c2DicadeXYZdGGVspuiyuzP8wIfguDW0QZrRh
OcCUR6E4u6gUU46wSS0WdYV6ufO69hTJ4Nea05wcOg9yx/YWydNR1Xl2xjynW4OE
YCbkty50zU5HP2dhGlUYeU1rIxOKrILjq9RbFoeM+INKynjcS7HGiSomjgHiLKS9
i7FsS2QU2Duo2/eHmxI7e3bwKPb384msFcw2MzrM28Z7riD/H/LLOHSmHlOdyHuh
MTnK7M7aD0GU0LqTu8RfRtYnAQkuzPJYyzZuuGYk4R2wUL/H0nfDcN+RotKvA3hE
VMJEJvNIz0sHlgNHOJLQC0jLbJwYHbO/elPMTSUj2SNeNYGjWjo5TmNWpcTH/L5h
s/UvQnTVbR/l3lP20F03hj0vkSrzIlD1biIYsufNcvCQyD3M2k4cEk6w3X7mqHaG
vVvUhD3PX/3amb6nsjXjqtJ2T2YP0c7oitlAC07m+U40DLVOsgcdNPcSYIEHZRo7
R7OSwXX+bLNF48fhVZKHAc6Ii6zK/498eolFOlByHsJdzN/J5zfZGOrZ1hC0KLZg
rW8r8UlKU4KaxRe4q2O22/1wWxyQ0Rt2s0IfxRvIVhvqgwZJsGaR6oH13djMfJsh
QQrVcBb7VQ0eH0IjEt17/MgieStw325/npSnmf0D2laze0F+pAQgvrCoiWU84Qcj
QGHXcwBhZWogjZBTgofsJCQUGKc4HSirWdF1whDO8LoF3HNaI3kingSZ2aPCz37g
/vxaoadKEHAc+NNGwNa9WCSVRA9VqKrpk2Xd1SKqqXmAJt6SXYJHONtnPWWrY/Dr
+3dqBKOgtsWCGOMTVRWo87QqLUwzzWiKM7m0rHtKfbNVsm7LbLoT7eJHS0cXN5t8
ci4YIGHjsnCs9bKASvRFsBT+5QwLwnskNqNRqodeVnMYSWl0V1XJDVkz1BTlMFJn
zo1PLXx++msKpKYEtaRxgY8f6DrclbOboU/6kWcfRsxmCHnc+1ioqHJY988mE/sZ
csTMYbVS1etgNFD536ys0stM9Nd8PmNONZeKR1GeQXuM+EJdAyDCXl1kW6uauiF6
eWHzjlC+WtEsQ7fPbjq3+eBF1/3qEYEFHEnG/6DzUtuteQw9kkk9LunnJI164Vac
BXijVYi5wjCmFfg4QfhgXpPO5BZaCXzUwOwSKLUKcvGQpLxPhZrGsA6C/uXIDWL/
Yd/O9SZr7kgAA1u7Op3D7a+PiGVQAawuweOzBKq2/1mrR6qgO+7zBEvwf28o7UM4
qtzIn0PBV3LnYIsY5rlGTcfP6n3UjFEI6e7da9Mn2H3BlWj87qWAfzQEYI7MBWki
lwB9VEPGX1fJjqSMjU9FX98PxvC3S6Qy7rztcT4qxfTXYebCpd2/wR8/kEUVP1+B
sKG3SjH9LKBhR1Yvwq5vErZzhifXYmDtyWa6KZ/dR91VHYQQFJg20RiALPakQ+hv
TMZ4uX3+/EKqSMu4wB/pgTCIHOP6Uckn4BcO3uqYsbbHQRmLMS6GB71PuWPWf/JH
0/iVn67O9R8Fv3XXJfGqFRHEivCLFXbVVO1DH0yQWhN920lV0SE5mk3dVw2igrVa
Tc/6BBzWHyhQfBMoHsPIsK/AFUAdwxSa4ozexZi50OOl5W3hD2I6wP8++a+ks9RW
30LhBfpH/sMPqB6aweUoTxiVL5NCLbEdBa62PAJuZ+poB3Bkp/EPAGRNughz4+xe
xlg0kjnXYGdK9oO4pKvUlBE5KQ0Pcq9I5DfWoGxjDxBvJIJgSzEOFPHeMNMbrUBq
HT33I4U+/dfvZ9zdacb021wH2A8lDkjKJcEaylZbogUBgbVlGRfXUpzGopmX8ch5
KYUTPokVZ7iU60eb5MEYZYuwmZpZivotTKtoTqRySEzQGyAxzXSm/TbFBfIHHHWB
YG/hFwFj6CPZCYw2I5SG1iBM2TfW+d33Ab0jmsNQ2FQydvkD+wBTAWjNwZCZL+IK
4nn7NfZwft+E3xcqfUNa0xbeJmZYgogBRJ1nH7GmO+L9QQH5wYw0vGu5lakBqsay
jkECe0y8j+725GDrQ6tub4DKb24G9g4sxNcmYIdhOnzgoGB3kIgpOwV1dCgQ4A++
ncyx+iMKKnyhv9zxq5fOSyS+Prg94DfXVWv/pTl0ijbCH36XLZp3JJqRplHk7tnm
1FauaxVRaFVaLwzmsCxZjTlpf1g9s6KchaP2xaNRc2+WxccrX3+5OB+E06VaTlT+
sZgLOo6VXF6jIqcDvi7qApuPlTSVRsuqjnj9jztOH9Wd950uXA+ErINh+oPODTjI
5iW9RK4y9YmFjGSF8iRjiyFnYYcNESFo96fExJSrHpI5AdLUK32ZOUiPB3HyWG8U
EBpfxqrVVryVaSooTKpyYcVXhS+P5E56nYk90ZFUp7b39FIIM/GQWqo/McehBbfU
V/M0uION1Ic68rz1YiQ+VqTuiRjrScTKbJlKvqhDdYMh53Zv0qUPAf6Km7ui6NfQ
2FojNSODz/D3D4varfmBhrRgMZx15/BylOZKB0NG2W2w4vs+Oq776gwkATJjHYNm
TI94yx2Z2OBK6HiV6xxVMQnd5xncsrpruSu9vMvhmPpnIXcEPaSkHROnBNjCvsoF
ETuVGw+XfKPZdsaz+vgrmkhPIpvEoVR3dJYoSn51UV1JgnpR/gPX55+kGVCOITT2
OF1WgMxY8QZH6BMkRUJkWJPOxblG7h5OGYlsQWRVlq4OSV57uefIgXVXe2e/SD4q
h8IjaQXr4LyXhnVTAhBCfAm3aQFlFYr9607q41/2LMU0O8eqOyr/6/NOdjzY4TSZ
s37epEpxWCc+ojWr1rChyIQQdiEuGzD5GcZrmIogn01q1cUGdLVIqU7lmClDUwnT
bkI/HbtnQzTLcMIaJ9fK5YZW6S/Bzjd0TK4KQmAoVCFm1cLCK1KEvs6jupCp7jpT
bhTNF3vbBpXjE743AP6vo0O143fowCP9zU+7DgNEw/vdy3l102eRzwCzrwjM+UY9
iJPL7ccjUNgC7pb/5lbKaSTIr/iniXHJLHEMjrpCU1fNMk5NHGh4GffN9NEjLfMl
seM+XxISH2f3ijgWdrch3q9u0YqYIQhG2XoHvX8EgqXrkeWUgcijAL6drfTEjEyU
DfviyFFhY+pEPqcbEiNQ2vnK8W5fkCEc+N0Co9DOszjUr/VEr15VqhfSD2iN5ovy
JEV+aM3sr0FhWOTo/x8FPRxrUadQhdaz3BQf9ozzciJHjes6wfJeW8D5VH7xC+na
kABWeah6lhPW1r2Q0vThpaqBG0vnDxti2e6O69EhIh2KBvYJaYrnaulIHRkeDLks
hLa4nVkQImULFush+oAvoRz/TWtJQZTY9czAdaCCQ7tZrEEX8CW4XuDzgBEa8+W9
ONMW6zC7KYKMorBhfId3gjPTshBjglVtUITFmBail53zZMH1kANTSMO93wGSUw+L
xCElnaaau+yEGrzrKOHcWW8RmRHwD86v1YXqK9P6tRMWAineJVY2W+Vo1voWp9gr
eNXU5+6JIoxB2wji5tcliwL3mdJZ1LvUc3BALi9GVpzbcdA4bY5P/OEgvzs+sOYf
wT95YyWZgMRDpXqtWCsX6btsL7McV1ufIKr/6+MZjR63oEodIhfqM7GED5Y0IPcU
JFeBnNi1QS+GRuGf8WU8muQqQPGvIEG62ZTqZ4sJMV1o2QgJivL1Quimy28u+dGw
MJXIyJL5HM+otM/0lOnz/L03xrilbP3JWsKL8P8NhPAW0PcOZnjXgnxswGpNxdOD
eZO+iMRSPjCqCvdgsHPdwaN4Z4q7No3v/M6lWyFg/cV9lukJaxl2DTN78DGyBkP0
oEZtA9NPcj70fK/IpweFvGdFmzpVwWlv2btsd2Bd59uiY0oATGKnkNbk88x1oOF9
KAijaGbrU+Y2uGCS50uGvgFeFbVaRJb69EgQmLEXTIL8o4k3PdcA7CcJUfnxAMFw
OyXjUcWRxXjCM40UdMtyky/xFdq3eaaKNCaeDEqU2ODOhpX96YXQcDCoF3TPl0lw
fPqty4XhU+smNFumSjXhSxtg6Uh0o79L0V+zpUW7vOkQuZNoxIYM1+fmBe5uX6Xv
hXYqQQgCVH9wpfq6mILF9Y7AxZ65GS5IRJDb6OAmeDXw27QRBujn3q5Db9tA0euw
/D+mFN5PXfTyxBRiEnzDiWlHhguc81N5Yo3sKfmIfNsvxtI8SWMbPdUVEKHEtLWA
zahY62t0zmhP3Zh+i+qAjAZzL5OdAckwDKfiVjrErUJSc6tMQIu+IKswwRYnRZEg
Iaz+5WkzPoFrRJBHspKAHXbGxVpU+qtgwN4mX7j59BL41/MKm/RkGhvMbfI7+Ii8
HZv53y0TtFMIq6Udv6w6/rUQxn63WyVRoMb7Mo2QO/AAW3oBmrS8nS+K3ynRKbOZ
D623qm4mFBS0M791Td24ziqEi5891ebwTeKj3BCsX05ctB17h7cgNdo8RMIep9Aw
5DgJ8jY7I9ZxpXAysMljOSZxAD4EoueDXBLh1nj1tNmRz01idnwEr4kbjV5BhPtC
Ns1m2QNQO9ufytot5V4oVMqfi6hfbwgDVobRCp0QMS7EwttxpThIIaEe2eg5YRlP
ZVBDVoY+Fk4QImxVBHPH6vnO8a1JsZOizExb/DLfsaHHtc++AaBeOY92xfd2X9qT
rZuJwSaY7QtC8Mc239ZIdxii84rgWQblvBfLU3NCMP3DzH/JPCrUyZHWm0eLOfqE
09Hwztdf5izVkU6lg5sci9RMYQtLobEASWBsQbVAnVVV+3Ao/01T0P5ObkOBSJGW
lQs1CkiNrqYrquJYN/iabqRwMF5FJ6l8O+Uf1o1ZUw8WFm/HFAP958HqFb2DxRkk
77fXbSLbGPIlWTNSAtME0vWuFPkHYaDaZVsCNvcpDRPUYQ+z2/jRib2awko36Yyj
W2dc0rD/cRw9///l3LM4O6w0qi4CgijVvI81f0zuvE2eoGC1EsAaNHZR6CW4DWe8
0Llf4UaEMLHKmhp99E/u+ic09I58d1oAuJJI75IfvMdfWM+N1+JP4WlQL3UHCmRF
ufgR56QUhnzEwvqrW1j1bu5zV39gm8Ky2mrkQiKc7qO3wdtXq7rV4sfFgjRETJ8N
pnb2yLZdkoT25r5TFt3HPEdrzSVY20MCVkoWj+se/vD9rprlr/wy/0tucbmQmpdi
1USkXbOiKgsX5NkWyz+Gnbw0kyuSBC7vuVONCgW6a2awAoAw9oeyG7mMrgS64DNd
wljdoPLi3kAOWlj/YFTOKi+x+UP9koJeBCzmeeOT7gvL2PR46buCwub54QZ5YcuI
zq4qMyI9BHK0ogDqrTNefrnwl3iD44X96wy4iHapljsx0FyG5yKHKpP6eEbrnCSc
3hA6VrHrkkEi1nPcFtwkIwUvphgQBdXkPArPsoo1mTADG8f8ZoiJfYH/Qz91GfAp
8j2e+o6b3sc+aYENEfGvbylk6CVt6gOj4TIklSGd1XF5YLEFhlwIEXSRFTMTbjds
pCh8dDMjmKaJxv5DrOC022rinaYxwo+Y0BJ26htE0J39m5upSYg27SvhbFVTUILw
+VQlQhzXI7eFOwp7RR/FVO3avHG8/NwgxVq9MUlQg+BgUt1uoXDSi0fKebHy/Fv2
4gdsqyvGiwiNXMAs8o/z+G3WBTxXbNRvEp9p+x0Bi6+V3yQztQhF4q7sOgkCCAHx
HcpU9nAj2tf4j8onp/MH8R+zvJ+Ra9obwI7Djm8smh5x/tRVL2G7VX7GXgj2Ch3z
V5NotGgCEXOXzEwawIueDqi+vmmc3Dj+EjhPgES7KLJ/idCkCOmac0Klg2RkLR6F
NMUqKKdZgLcGH86ES0FbcjYeSrYi3wfFNHi5c0YRBb4Mc3Y+k2FOveGJgWnje0cw
YM52kl/jJKKzC+sdbq9yvRBuZW0dfdfGvKqx1Hy31M6IGj7grwB5SHu2OGf8b0/H
gJDk0w0fvwnDYMZYPu7k68InNuGQVV6gdD2et/2iKvrkXWKd7ZPBKbPhd+pgajlb
uncasmov70ovkEcU7ptCJ1QXK9s7h/ElnmHpON6OUpiWkJPjaP2xHrgfCg2SE17s
YngY7Ai7Ut+q4eesY0yzDe72XrFOccVW7mWIxAiWeOasdPpjuGX+55syAwfYkZaN
diQATD/PPgx8TO0nKIUo2qipSnau6XQQZGw1qI1QdX3eGcikSqmRE60NCjc+iFCv
st5J4H+wzEqdpyaDRhHWY7qAkaiWqhMNR7MSGfcizmHNys9paQUT4EAPxthCUyhe
wH36+WPK+Id6aXvKGaXqrPcmworQpjgUg7FoYWr9CXOSlhOUMMntpvOxAlwMVA8i
8V8tzQJ7Bc4fL2GIbFszz7UQs0QGcDy2HRaCJwn81biElxlqzKhwGgdRvedTPOyB
vIzK5sU/LfaR0fmtJ7dLi3591sA3VEgu66rkWnNqj33qrWCab7w9G5JdPNodt7md
XA8CP0Jia2Ds0gaAkfUMcwdmIRfLgEPuG5woYzEBmKrLfLhrzjSPdZ4Hd0ik/pcm
pF4vr9PYKwOHhbXfWgIBr12yRTqRFppVL0LO9SwRBHwXnZLlW2/vbbqL0MdnG+Re
6fBEqqKqsfYqzfzVHpQrlpUOqKsk1LRZ7DIAU8z6Cu459XfgPQBghtmRWjdUuBEu
tRzPYEsERoCQ+rc1Zga++rqEIOmg/LmdM98uehfWxydNRQez/UuCU12Rc2LpEX4w
+EhCtImM06kar/iBH1PZwQsg7Q4YaZnmmTZKrZVnMYSlSbv9XkUIoO6YYQcYpcwS
EFfUhZ0a1dMu4JWrZR2gJPD6AfWe1/NaZexR/qVUeFWg8W0LevnaOGz+7JJx7T8j
9HY0cN/Ovbpw19i9tMC+gopN7RFO6fVooXjUAmBDqBTideSYC0bCov6cEZoN4Z+L
4C+6+7mKA2HzlW+Qqvaw7NCQ64TnkhTNYGNExpDY51fY+lo4j8S6GSN/eLCs0Vms
bMqrxGexl43yHis/9dIonLRrauNFeYBG4+4PFkefWzv2Um7Yw7KYy7a1FmpmNNX4
QADbfMsFT0TDgl3Wb/UJzhxLBtFD3gIDWJ5foKUhKWcjCLxaq0u91DE5Jj0ZfrCq
QjJ7p+Hbt6n7Tp5dCOqBQ1UR57Scx2UggIOm/JjNiHmCnysIIx/zjrLoQicnWla2
qh2i2sRhhI7y446g/SwBrt6nRlAIUzyh+RvP4AgB5LY2LZJKiYMrby8G81aViD0T
z4v2BLxbPZ6oVA/WomfFx/3asOv3YilOfjYOFvh4una5pvGBtvsCpNTsTPCDmjtv
TJzGLZVKnfelZbFrWHu2hcq0R8gHTqgrSerY8urqlBcWJZyuI7XANe3CPYcS4Hbn
jlm+6mFsx1NJ6cOHZIJ4eVXh9KrskeBbLA0xkaXmD7JL8IbycNS5rUaDF8zqnN5Y
5jrwnDFsoZM/ushIbPdOvNH82V/SbFb+r+8dPYaVRelUeSNoP4SKS9odExuGNW3k
m0lPPWIuoquri0MRZp4oaSN5QQfFUGHu02QlcNTnK0593A3zI2AU3eTwgf7zuz7A
CohOzFixTx3gkndvpySVe5l9lz5PZt6NgEAer6Ibjzx3mKPWAw255CcJE92Qv8dj
6Aalcd7EyDYOKXrF8ntjSiB6fNon4RLpFmdklTA/f04CLuH4JZBjCP8phRFStKjL
9jIsXJoM7Z8RfZI8XKHvaOdBzojUK2/jP5iPIOBkSkrwcMX0K4ga40xvngoJJyyg
nvnCv7WMPN7k1RIdE7bGaQ1qOg7ekDUl7mVGsQrJ9cwuC5KnDnUjJyaI1OZcyXv0
3ZJqwACmkiUarSLhF32P7DyXTL9Xp1PJ0ruR2aewMyHISCUEVkkVGghgE0EX5hva
YnN1NmEJvoYEox9MfAVLqrceG8p47cecnrfWSm1vf62vNqfOZ642nn5NGPkATRam
guiizPSqhLgino9E/rltUIgPdQVES5EsfQgZB7n5bItLx2edkVtpF6TQD/Sh7qzy
UmXIYHU0o2hlzubBW9jFHxSNp2fzUf44IirMg7CReLLyL2NiqXUh/mgQZW1AWRYZ
QnAhYaKhpyduYQLWn+djt+hIknPounIlyCxcdTn8VvAtuloXDXRIGPCkhsdJTmsZ
ln2aAmHMn6cJXbSQeCvXBje1pWJpCBSmghGt43viHCDtijvUguOVX2aTUMw3Q5T4
Cw9sKXMIsi04BUcU6D8Hrs1e2z1uQVLETip8D22RiZdEdNCjrGU+F6pX8CsqeExQ
tJpV0ApGl0jsxjiBSbqESKBFbjCAtVB5KgbnRGRVJ8ZFm5e3OtF02NoCMPPd0v/1
VcWsJ+e6fTC167Ik7SloQ2ccYiSNqsEGWjjYh7m+wKREJmsgNKwixl7SqwW5XWyO
aj8SNNR5Eh8Ky47Fd/CB0s6G4xR6aMP+VgQP6b79SomNNQDRSK6nOk4MID2UF4sJ
wEy7asEvQUic17x7ayaGcznuykYvuJ47bZCHzBfuXGrHHq0dh7XuOrE295h+8v1r
SenywY9NSN9LO3uYuuD86qH5yHBf1JNtrkMvsfBmzRKsSY/sWMIek5YTH3LB1XRD
Z2lx8A+5hPEzshoW3/rGayIngaH8EdPTQQy4FHvzrzN0XYmmblxWcs4VrcHhVl02
IXu79FhwSMNcqk5bz7DSm6KXcCWO2fTuPXBKueDsnvah1pubWVylJpV6b+BI+h6W
i714VRqol8N+uLc131PF32wUe+XRTg8TevwPeQPKGfKV9NLiaCp/iYIVkGpNUhC4
mv2fVcJkWopqousqZZEvEf5JQ/uvey4toX0yOkdCNEZcsGm43v2bxyS5Kfocy3Q+
S8iWaQXf/uDu5j7d3OIbpUIABpaXFaIqUJucoo1sVGeK8eupKYUY8/o+PQToZGPi
mbIX8JeZdqrh+FWhr2HmEoLv8YP2rj+t05oxaDlrTi7Ny/9jjlmrvsAf4uF6Vo1G
lD71ge0utAK8I4V9dsSDAEWxyDfCjnSsCjOssSEJnn9RfNvdNxnWPV63XfllyKJG
j4/QlXkSYPY8NFodKtYyStfLLRt1X+53t5vIPu7FV4EszeGQCf2QWSXlOkiQ46gQ
hinzUeMviCT49eW9AfHaD0aKRRYj2qSRUYMoJXm1TUpUFTLQn7F7KP0ubUC4DM2h
idmvI0gtNKW0IMiGFMm0bTv0jaCYeE01PBnjxjkZXtSuEqYFaRmKwHhR/iOsH5pP
20Sm+ZPzddN2yKnJTGblrnsWNd3lw27AzgHVRHWjS575+iHt5YEwEF0IjFaxAYJw
Z59FqmgLeQptGqyL/4MxOGxb4GHu+uc567yXCKsnjYPCK8Oh8zU9K8Lr94L01apD
aAzsauxIRxPM3QYUMTXkx389pp4LtSlJlMgLPsoXbV472z4+rTJzN6Yt3tNhniSN
iTdTaI69ri4zTc5F76m5pH/t8NshzmoWXPsZIjthIJBIwir40qIxkJS+OrflUJwI
4iIepTYT79C/FjHh004XBBrFAphvIpZtmvZNlqizxQ5nui+/zHOKEbYYSxN3sY2P
zEWkrcLdh9WIQZXI2m1qSYMkgxQXU5eREDGhT3ccZVaZ8Dhn5tm37snRAuPFhujO
4yJVnww/dbQTM3E7dGPRbV/Dm7j1kiusgQi0xSTyziH0OCP2Sv96nxLtm5l/fP+D
sKwtXMwEDtYRPE0BCyyoqkeuYjw2rMN1krzbW5ZvReooXx//gWrVHA93ldf1VfWN
wD35ZqQQVbIOD3qF9POCJj3nY3EKSV+VteaaZlZw4RdNt90e5JJgVEGTG693uT2G
74tzQvzYlrxTg3EJucRo/sOiFRbvfeeOON4E7LGr00tZgsqr8kp3XpnwQUfGeC1J
kYpNxzaF4HSnuLcX/dAHRPwDspDh73GGznNb+zvBXbmcWGoa15neNU8iE/9xderP
ybBm3iPpJUtor+5K0UfdMtlpCdQ8dbo/E5p8hwVQ6052jQ2IxXEwe2fxMdGqsI0/
9ZgtSAxwB8pT6Sq4qksotgRNDjTvp6tcjaMlZiZIVO/x3gLd4lGy9foB6sKmxC6p
RYZ4Bb1r4tsHAg29GnfbS+n9quIHM3NkdCSgaj0sxnortiQ8EU7+InKtXxr0OXF4
nBZn9OxuOcfjOULPDCc+a4UN7jDiXnRqjq6ohWfkOgRdrM71rhqiEk03wIGMf8Wl
r+DeAaOERRnBV8t1grSCXOLAJ11ZyUA+OT/cCmTxCCOhGTl7m1fF43TMY6g/PPmW
RuFM0CKO+Ugn3usMX+Zeh1Z+LF1CZP9pde0Qo6AWQsxzLabxuJbN+FMyvK2StJXU
1DAqd/R344BGYvzMFctDmjSC/+JhynREha1ed+F5ep/ieC9ovRakJ0/T5CpyPyUQ
ynPV7Prpce18FYHeS22ijme8yx6dlT4K4yj8qZriOqKkKelmgoaL/9n2OSvQau6L
lywMcU2VOusKnB+KJoDYVcz6ds9gSIahZeGmwJwGND+BdXRzD6fgOQhX2VxgPd7M
18lJS82xwg5LjsNL7uRcIGwX6zrfdTKBMWD1E0h/VhaHR5TBy8PbSLb4LDmyMqfO
0rGTcGE785LMRL3ZmuW0he42nPLwk1rYkPIKfIDwmBZOVaJ/OtTjoBN/B2Gn1gYF
lc8Knbh2U42gll3fC/NByUEnOH0S9rn8E+E+hJSiqOmHJk1pP4ej96ZeSQU1Es32
zC1FZjDiXq5WViWhJRPnoXqR8sbD96AZ51ICAuJMYhf8dVtDpa2eVY1dMEr+b+wu
NC079R+sb9Enzky7v9yLvajUNc+RXr9vz1qBinG/5Tse+huTOt4V8/3aqOGhfZDw
ND96c1gnVxrO3wRFc8qMC+afHnUTT2PDYH7j+NQjrfkb6tIxMAWzLuEebCFE8d29
fU4Zx5QTZf/1Ynydr0udSSd46pA2BTDzLJfMchPJgF8AHu7VO4kMb9r+4/STlKkj
WPDm7hEdRrbh0bO9ZGV9wWFdVk6QCAhdkEpW75xyh9dMI10XhmBxI8pxyVDYjrnJ
T9K4NYagUo3KqD4t748QR4H1BSX7wcGEl9LwvQN+mBRpcstAMsGRMG2ASD8ST2Lw
yYrLSCyjb5HhUqqd7lv1gspfvjpM1EFp2V2kme6Gk5ED+3T0cfwWNMfRlNUIxgMd
YzjRPcbdSIM9By67oZIS9/nv+JqFpJdNmWNq6gnKGBjbDPMJ6ygQk6OZ00uqZQO8
9+aGKVk0SqiuurQ9yiWr8+3taGYIAY7YnJwUdnKkTJpuHsjP03PmLBPD8rp7HRDx
J80o3KdWXtwmNeNR483h4OfDtjIwjkwkBJbJhtopo6PoxZofJ+HBHSkBX/BmEq1U
nK93ewdfjRGCiZ60rDz1ZEb7Ky86Z61s2lWMDKX1MFpvzEj2lLu9aPqd+bjc3TBs
Uv04Q+w9JQTcY3/2ZkeYoCPchmB0Rrm5EeDAzCcXW4gBBwPxqBTpbVxLoO7NgfsI
ld1YCxdY6Azn41+12W4VVzgKT0/wNPRRDOlZ5CS2oXRuN9QME32jEHOVou+VVlP6
OjHJEiGb+zocJWpbEgad4P8qmVMR1VlC0NMWPT7wsUIiAmKBuFOk4H2gte3aD1IL
/gi20eYKo9sA95AxUWQt8uobwrROxmMTuh0Te8xUaBULBgYVSg5K92/GLwBN1BGn
kQHnPjhcUqjGswsCRaAl4CYY+ta3M6ZJQnKsv9OEtM673eY4op17pvklfuok7aFu
C/uWqeqTbAE5gJ11697h5x7BuJa4NdAJW25FOlZT+SuZw1o3dT3IKZzeTKQPuKPP
QGtKo9PsEe7bkm6FLWZH1VNFw4NcmybwyVtcTP/RozKnSSb82u2IfVF31XpksScE
CfQHOZVRgUxELSk23fzMGX1Ttun7SphkB56ZjRzGG+5PbatVdfJV42Ll/4XPhxv5
YeJEFORzYrY6CXOruaLe9nm6hbaNAmO6qqJw4uuiJzgdlxXQQHu6rsmGG6HK6JVT
NGY0TDydk5msut0X5lc0W9ywVaLFPQB0Xf4fW6H6YNcFj0VbBuIQ1hnip+qEKnQM
4IDSBEW2uyRezoWlYXBYEbUQAkfP6IQsYIBPbKWsAN9TsOxOcFJRESKfRZZ378ay
kpXbXryvmXDq5qfI0zmSzzFZCIWrJPiuamZTosZ2MSisOp09yX0PxdktrtQcLrXR
cvkNwj1TAobn8QZaV9l3HQuXOSbww2Pw3Jups/eoKr3Of0cEg88t3bwUM/DVIyR+
rrwUCc/9QOSCKn34tAZL4ahvRvxASIwD7EI8DD91Rg/BSFFRZjKyMs0wiNJQL08G
bnmHHwA2U94ZziyBVBFLz2qKtcCicc14oVXkzF4ySsWhj/iGt23nBLgnx9kFPE9X
/t2tj7fgsJYjXAwIX2wDT8vhJALCNQ1Bt6/5zYiiGwXDFYcSpR+oV96PTXOUXk+3
xlNKdj55e7hDbWw88nlxBi3vy+xC7JE2LXTfQnUVPvA7GvL0/twxOgzz8OqgqK+v
v2TDG80V7zn7+4zlR5lGQl8QR7pakS7QnlK63T1SfpyJnLame6H0wUvgvCy7TWf9
DZJ0IQdNJmnX2i4Qs/U1X0s0al1IZ1w6BSlT2GV6SGYizTBmGxeTTihobsJ93TqW
ZNlMUB5CWcn6yCBiRAnlk1gAq5ae0/M+mhY1odaytdg5hpDhTq6xvg3XOhmsqrCx
O6bfOanCM01zH7Dy9yYnuKdeLMGefmwOJFnqXS0FYlDJmXebF+I/6/63a9YW33R6
TNbFVqbv860TUlwC76a3iQ0sMv3w4nmxpk/zVGk1vIVWisqqzs5wAUwIQI8s02Sd
R+dJvJUpHaZnwuzefyJhaDsL6T1Pik1+kW+Rm9Wpl8dTcqgGqFtGple9e4N1BVJ5
FNdWrhMtp3a4m9j7kXNmlOaVb7ywpobN5py2VUBBvAFaLRZhDvYzDhIzPB97v/Wd
nLeqWkuv+tneOuaXSxzIfiGvC3e8+z6NiT9qpoj1lkHyhh4ccEhMN/fELBWzLhSA
5ej7Nkvl1yde0kqsbNQZO3uVPoGISRvYU8as8EnRJn3/o7WI8oEY7SCzVubIPu8a
pZMjoT6ZCXRZ+LKAMWUSlabpYM8/PbyeMdndYvp9gIEtA/QjapQMkXfY0sPz8RJc
+dULTQ7IncPA1A0w8ZusbYLdaS56EA+hpd962rTybuOdUXGUn6hdpPoBItmgRGXY
o9J7k6mMLFsCfBL8nooCPUyI5plmEbZsUZOfTRgQ/sXpgMWJ2LfJu/SH1QGcTvJ8
VMIeit740kqZctKOgL1tywltcfeYo1LYYpaLP3RyF409ctTKBlaRJXblTC5PrAyl
qXwhsHPfSoxnbwF6VOrf4gd3kRnMe9MHK7K+9orH8jBPh0OXJSYm3uZf9oHFAxQF
FLBBHXjOY17nUbOQF5ci6PgmApS8fehxQ1S7VDXcNU/GX5MN9VOnR6u0/zAV2zJi
PWEI85v2pmxlTGhUM9A4zRH6QgFp4RO4WD4c2ZFS34bByjzX3obmTjgVRXaYsiJ/
5nKfNqLcM+6hZIHoG0GZXFxsC2FOHMlwmdXyYMQhrT6UDr9j9fpn7gVxTq2dysdQ
0EMfam4Y3qN1XwJURR1CD23il9taqJBVttJZAOi36j/7o0jjALKRhtzC4Z3rMR8V
vZnRdqMK52pnQuGh6cAF0LyC1Z7us7tupA89u+Xgv3LkJLoKCHYsVotyRmf0j/7r
4Fm3o49gYgv40qdaNib4k7DngZg3v0iebzpzSnMZXppOhZUOv5pu/qMU1cADv3SN
12bz7gKF5Vf3OmRDcAZwW1TUbXjtaZBbu7gunOg7F5rL87+/K2d2QmDhOQIsbcHv
bkLH5oajRBJjcsyrZOkqHcPi4E3MFIkKJas5bUVBCi8x0Zxj6NT2aWUMOy3BfX5D
hRlotAqWi/SH4t5cwoAWh1wlrqbVS40iiR+KdntWXyAoGDbwW2r5yXHF26nbvtLl
KYIekk8NSverGNOecb2u3de/3BhSDZSiTKjWqfmeZuK92g7sQPSanFN2g8rNldJ0
yCiOjWsyGgwVwdbklb/JuljEobDx8TedsLpSkv0KPpUurBt6amdkSfRZ4HivA2Bs
jL9ANoYf1hikp9ks/zPYem/vqvbIuB8REEMlEk2UX69ws1ngdyn8gJm9dwuNKdSI
vY5fbCFVaRRTffKDdDpz1e0r5YwieDLm8CQxYZK3MKhif972zC2u+QhEwAf5U0bv
A88+/nNdU5rgLrrFsnCbFnx2xTioKaMxZTW6HIdDHIuz4iVetntm/ibZAQ9Squo5
05WMMqkrHS4/+9N8g3mnl719barI7NHgMNHDZwdx9OmwKlkrCDtjL/SulHFH9R3L
q3u8Tr3aTnJFQDexEMiiWyTvjRmjugSEaGPjcytgsqwwXVkp0faz43U6T0aOlAwg
OeoouF1sb0NGllIOOUblh2nDcKhrP+xka1uXHUw/dLp3k7f12suVa4muphSfbmBt
4Nym94itU3Ur3f3M2GFXJ/tAVlAffsU/2qYIpVzmAnRU/s8Eic3mFGLw09Frk0gA
tVTpUfA5aQ0vT+fsgggsng8SJh88k8y5eFUnJuIaWBsVCbqLh63lFq/KT+Fh8gwv
tD+ye1n07cid6+cXpnnY80OZ0arXZVFLx4WMfDbT++P1TIGjRgJ+eeXrOhblA9CR
RfsN/nSOi4Y0jHcW8CG2NCJca3KfbXHKXmWfESkP3HBI7W8BWKWhU+tFssgoduVK
EI4QHQnEm/FGnkBqau+0a9lqTtZDaf9UTt2yvpYyQdWSV/H81Sk4y2i8948acvKJ
9fQ919dUyCXobV3Uya127DfIux7NxgDy6CbwyrubQeR6SmOmy5rn+wHsEc1wZLMk
1dMQZ0FYyqtp1qkR1GpdbE3AY+tQH65a6vJwUgY0ZifkgGB94FeyRVzqgEcRa+Mf
6Muzi8y9lfpbJJoCzT1fxfnSe/J8joMB2Ei61XFng8WKQayv232yxJiPiqGklP71
BfZqA08Um9OQXCcuRNoWIK/+srDaYDU5RdQtS8s+1Q+XQRgiETOE61zdFZqj/wWI
NSHJwIayZaiharfhNY6mB+Ot1iFKDOCWaq8/iybMWo62gt9TOH0Z5JMZ7bxFNVEk
286DB17b8wn6fBxTNyY+ZQMQbJ4i8/xWoc1oiJYVA8aANrEKrVYUdJUd+c42s+HS
1crmzGlytRJtiNtDceScYqQ73H7CvjuqMqlPm9nf0rZjmIRIedxD+kuUjN01ufmH
rLPHsA8x0Rw1eII25RSXNxqxbxRjAp7arHWOxZOVrXbseD11WpiWMlMc786QKxWD
YDv8UmAlp5LTsindSGcUX8JgphszWoROeq9CMKRWTCfb2aEDERZ8e39in+7qOrqu
VJccAFz0xe1Mpl9Z3/7p7h3SKM+R0z+GXoReEaGPcrNh0dp9C8iV5CsG8ITp7+zT
TzxumO9hTpuDZ1AXa2RnQKhjRc8DAMFin/71ZaMP+TpOfGbKmQK2V5vZPQJzRMYF
tBeTpnlo6rMh3JDytrc5HUmwr/7zxVCHinG/HtaDB+YKZkZHT9psAz4YpRCZQgiT
2aGkc5oonSwyGwUrjOn1svtz5M7jH8VlCZh1usKnzNnwwHm5odh0Kdx/RCOfz68S
1JhwW1dwzT3En8L8IAHOzyvZgv8rEmyL49BpgtQD3rpdfB3/SbSztsUH+Wcm5iwb
BWBMNsMv1lciSgvTooqcHtCXHrx+E+68oaYrvnOwB20trMN0/k5PBUWsQhSX7WYN
UFguqoqPaFm3oFbZtNGs/PjFJ/ldZ7Gf6WqQjFe+1Lf2cIovQl8BZEGWy/V9wFzm
9dXRTqgURJHDSUGuNT7aZLq7n32ecKAXPDxCDApPKeUNaXf27kUPtFp2UpSnR3u3
j0AXLUC+GvtVafsmE0sPCOq8R8ZxyPRfnlC2ltWcPFUFjpTq8i+u3PklA+AB2XEb
tWFYsGkyWiCtN08qRRpaSNzhWL32rB+BY9v4680eWXJv1XIq0RVm8qNetE79nq78
ZU8u65VrJT5VkZexn56/CQtBuINrZkqrwjRXO1xY4IUCtoXwc/pXkyDh2r+UmCZ+
lZZVIhQrAwK+SNkVpO7WNMYCMpGkYVqCqw8a/iC4LllMWAkFDOwoSydTZ5OHWZRq
9QloV3qtw2IvQogbbsIBB/5DXgP9CSjcJ4SS4Ook/lAkCBVPq7/lvi84Hnl7Ltke
cmTUZYUqdE1art1+B0Umi+d5SnIloNyUNylMgQSbhI0WqvF7bjILzHmYa67hcCvK
R+UtjdZhD8Z70xBMlKHCpMb12Jm5djUWwJ9K4fwP7SF7VnfClcEXpMauCGwGMKqz
HbKLaYgbZbo9vcjWJItsj9vwMyaTfe5jU7J3tjx+Rbt801RECs/o94aXgMsPNNEu
cOCsJ7DYtzrsYCY+pF+uDNfaU9xWkiXou6Gx2RTzVfqQT+gfsLIo8hfsP12bKM6g
REDrrJ08H3iAGWKtIFWP0+gSSRXHQ/G79R6OEtpceQRvOkkCDlCBADmUCbBfMlFg
YyOhdEwO6LugxXX+A8Hu7rlE8SPyin43txgndoas1T1OsRnm7yztz/ETAiajbiJW
D2eTtMoE7czmz7RQor+19Qhaz15tfNt1LcFfGZqOj2rg+l0bLDrL+lnRND1iAfSy
AOOy8Dec2F845g0imBOsjArHRvAfRBjTJSkQCzLosV+6Y3ShV968RY1jkVweUcUh
QxsFJanWJCPapdhkyh59YnkrAR5uUXoBsQ6OGQ2jEQhL5y6IwdhjPog4XKTd6ir/
ph9BUMttZlsCpGayZn/NR+oqw0Qh815Xszs+aGCdV/NZ13U7Mm4n1PxXiyh8FU8K
v/3krKYWjVNIsgeRHfoiXGLagIfr+LsNQHNXBWluxknrBMamHCvI4CgkqQT9MxIS
6HNgbyiakpQDIXdhlhUmETPNdzK2XaCNtkkE7TEmAGwUYAlDaLPUYaWFM+IvJ0ae
oHH0RcpwiZVJ+F8yC1Htbu1ZFAVRX8Xzy/fNDBrBB6lXM1yPbgug33JeO4/tfWrU
wXCZXrWkDGXkSuQcRJN/rj26miXeOJNTgxO3cr1iKNNqgCsQV5fkXhc0agd0tU+S
pvPZFHUkTa6Je1H/1iUC7FNjX82klLHSo5/gskzUrIDFhI2yimfHIdTtT+Wbcb5H
s+BCXT5ZWZsjxCZZUKeO2rmDYMFdlCseQ5v/ztw/C2260rl1wVGyStJM8iVztq9c
zB6j06nbJ69MF4kGT7DJzMmJEsgb+vjoyFOWzz+o4vkFzU8t3myucJDPmdDKkNBG
+m4YBJVOOKO+6oos2thX5Bh/7MkX0+u3Io5uEON6vY9Yeftwl5NKQ9/VejaIdjrQ
RHFx4cH8FT9728rRmPW7LJQcOji3/D/reYz4CWqb1S0V0G1O1AVxSdPZHkWPq3JC
x9hCRLr5oqKWseNpGEEVEZGGhekP6gld/pB7HqWM52CaoMJIOBve82yB3McZEf64
i5F6pkIuPFRTjjBsUEb8WR4fNOUWzk/cz2mtGhXTtJxMacaQx85lq1IHkFqBqFLT
C7fWXfad4tK5a5FXVPfYXjwY33CXAOF2382FiqkFJdXv73Jkmdy/Av0pBVqgEX60
iaFyvRorFIuACUThH+4jq6ZGTcerCffmbLFSsMZXbcLwRFVyarsOak4TNDhChTWg
PYgMGcpiCnY9fpg8EVztDLg8C1f7X0RZ6XQViJsAr/BA8j5mwJmvpzbbMEZSM3Z9
qL0qisxh2aEb4dJq1roou89LKY1hyagpYobkn218MTNt24gYjhmqdM2ekGP0zeJH
gu1IEgzWKkPn/01+t28FHTLAqR8DConuFu8ClUrNHGjQbUWXMAZa27EEjnb7Ajfn
fzxwMIbjO4VLuDg4hWcROqEWbirk+p+yXsmaQ77rEcTorvu+1cH2k9YWgQ5Eqr89
ObVpjf4YnXRjSK2mgrSwv514P/LkUOBTqCOEA0UcPoi1AYtmPSCW/UmJT6PNlWbf
Erw3EO0AFjNf4gxbmq7QZ801SVk2UBi3XZzeIx53JjM4UQA8/cyvK0XDsgterVF3
cD5d4LKXEpaNVVgabrWqzEWHhKQWQtkZToQv7KXfSIH8BaHlKG4UGbSuxH/gj3XU
EG3s5ii9WDgQzTNi1AZTCsho14nhxfGSnaIC5nfvaRK8re5sSKR/bBDq+LFUwmrE
UbXRIyjo1QGaTPvQ+hYLlFmHup5VFeZR2up1Q7FFL5wDGsr4VdWkOYm5jrAArQZl
xfeutvr3aVs/Nt2g1RJCHq3pCV78h94qC1+qUbf50EbECFc/fliALNUU3d05829O
gGUOnoh5U3G18QHCAMnJsEdbqBmMekAwS0hYx8AaM5+SkYZocOkXJSMKqDdDHi+H
Ol7YNlx/vcqmmoQxA64mfb1iPjPb7tsSEM4BIfmfCRfb7rqJKOE6J3i0scos52cW
tDboOhf/sMt8dqQlYLjCXma0zP4dkAR0e0+SCFVt3rNwO4enrH0UJg8I1+YaJ0HZ
Ve/kuUvDyKl26oG7vOA0heRgzfHJH+a2YzH1RUg7eA5PBvbcYS7g8aZKNdLkaEpN
oU17bXom2EdBwrdhQxfRbRzN5ckL9s6oUF2zlNIglINJF80Lr/iKjC58+CM7v6rr
T6vaYqxGgicIXIUJNHaAZXb1jvMaIkE5mHJhe9oqhzQy+5UBFeUUMOQ19aHeWEB2
qGxTKRuyw9mu/GvneqvWvLzDl8RRhSoBatw5NoqeqHrxdFP8KoCnwQg7Jk/xJae6
bGO8/nA2/iHlGraFkasC9UYxIPkeKXfWblAl+oGLOQ/9Rafrv8dkn5BDyw6EAALm
2ZixN+UrBS/wqPTo+g7SAiT17rOSBqHfSF8eRWWKgjCZ9EWS3J8T3munk7wa21Ef
NPCEIRe594HGSzxTlwVbWPLvueIWirjjGfvdexA7qzONJ6jhJOoLM9dtGCZXVO2r
c44T40An0nHms9RrdfbIGH2sO7DgfEheBl3slqhXVIaLms22r3dZb2rL3L1URxwg
A0o/Fep7oPF9dUtL79E5TqSyjSTyek4wWIVgcCBXLcEOQJOFb5R1alZoUiuYDv5h
pMHj/+j84qMk/uZfisIg+iFUfwVuyuzxak7VWFLTY9z9YtlQUSH+8RS8+/2UCT1i
C3N1B2qmzJoXNA9muNUuZAt1r4Kl0hxwrkCBoQGf2io37evb1LjYOY7Pn97UEZXw
zbc3m0kGJ18rPWDlFJ18fL4/PvSaG/U94qjnuwXQAviOljECG6SFEwh/+3AgSAbK
pKdUoitV8hoJfcOjjsvpA6c+4ewhVZW+UywN4dqfLDWl1ip/+lFY9kXmO0lRvFgK
1vwZJxr+wV6mLYDZwpPd+Nz6EdEAJVMyG0R2YbP44WrURxocs5fkVzxhx8tt90hU
86fIvX71KdCBl8s8oVUvlpet19KoGwnf8qpLsvq+NAzE7e0TSxf/ZB9Fnhg2WrD5
JAOUewBwSDdvq+cAM9DTggY0Nay0rZtrIudZe4jh+NIct0eq6oHqlbS3rQ7NdTYS
lhgwOtXR34njNWvvMPEFs2pULz7qgzj5ZvyOZO7aQ8Mhm3vmiRP+CVqUVqSUO/4M
rKAkaybmNNgz/d6y3I8Kilh21K5k93gWcSEb73aAQH23SHpUjrjJ9qCplgmqmFWY
8K5qiHw1MsghJT7tNLzrtpZSroE6S6M4DjQ1Cg+VVYNrBCTpyX21aBdtuUakSejr
2houpoQl6zJlZFp4AaAW2mFrqiIhive4yB1DWBwN/eA1HK6Sqr+wFXWA9bWMhXaR
eSbVVNuOwcB1CKEEb7ep1enHkkfWB/zDuLWP3hP9O6lEkZ96BDBAOc76RR3u0sNg
8TKhmpPltkqR/JDad4YgXHzIr7/gsrOUf8TOTKrnToZw/V2AgvkdAis53vytwzMY
r1lnKdtqbrVT7gq8fOiRYDezX7nR841tobeIw4CJGBgH1pu9F1VnTmqb5lSc8pEx
pdw807tFWFvmWf2Lh1czXHpixzcggpOMPyPX/62wjQc9wK5bzUSNJjxzW930FvGo
Q5uCHAOOqROnUSWahDGmy8/05XZkN1rOgq4llzUEkIxSYouGPJ///Fw2g1tDdqlc
9ineolQcw5L/uZyXTggh26Kywn32gzcTS64zFBzpcVCv1bpHDDHud+1S0RYAGDJ0
q0BVE02ykWAxhyDQ51oi/Mb9ln1fIQ39LSEKAJ3sRGQZOchwc2HXpJ6h8JW0WdT2
u9LKcT/2ax0ircN1o4il5YYgit//MDTq1P0zQD7tO9CY1ggTi5Zpe/OmJ0YQ7pW6
BT0jzJ6oeYalpBIxUuQB6xe8q0lEvDbZragG4jz7vRHEv+R2rhPhHoD/E+/bgV1L
hHRmF+JUFSmY4H4HvV0XyyBrgsIu5wGSfuleh0wrPokgFsl05NDgUzKBP8cO61c1
Uep9rMJ8phkLT5Mww2bKuPRHpbvOOPbZia3+Uz2iw6WIv/XW5pZt+zWq9pqyeBvU
T1vev23XkwPUQErTfcaK8ZV4in1QwmwdFOIp404MDNR/EMHFtzJSDTcuGmPYIM47
szoyLpjVWpucihRZ0QE0HwEooqyODilzI9Y3SKGmDw7/QipVi1dcqD4EpjJIo2WJ
RvSHIZdiMsqXkHgNkDUuDYX6hGKgVHpGmyex86AiSEtoThokV00KHzvb3FUqSY0U
6rNsbf0P46aQTSca8cb37zHzNMt+jfc5doZC77Bq6w64LfwUhUZAXqtftlIw7o/x
1f7Zt0vm+NzLjGGevjXRgk5vjE7gtdEtmpVjHqibmgrxQujMFzIT5uvd+kAJTjJa
MTeZvkXF4IXUWhGq7ricz3NBTWyfoiILa4vcXQ3XZs8mO5P5yH74Exky68nC4aqD
aLgYOuK1BTMurWC/68AzMPJyUa8VwlQqGTcOfnUS4dqvvZ2PBwxepNdd8vbH8xTU
mKtU3KXaY/A3UfzH3Wo65lPg4B7r//dhSqFbQMEnCnCQpt37misCZ7L3sDtY5v5A
K7FUITE1H//aIhJVBDj8S0jKGivJd6dtEXM/iBn28XXQqxEFYFwhChb8zSnHq73w
SL4QyYGj5fllqzNyB6ETHgvP6Jg0gUZa+n/s6vi5yskKfEhyMkRYWC9/IIc53evV
YBQ8Y5Fw6h+0z3aiuYQXNY8dGSAkQfNRzi6k9lm6nwGKuwN+ziGAGsPh74+OMvvT
g2w6MLseYRRyeaz2cLLJjNfM/VNQAH/qiEL9ipFc7DTHKbLo2lQgUs3p9iL+jJhG
nt+q7GF/Yns3y1YpHiPnU+BTMpEiC34iY4fVlhSa5a6+J7An/aYfSUnoe44vloKK
wRvyRfIjsijL/0xCO2LsQKNFPHP2TW3ki+tq4WOUAygfYL6cj+tZ1hmGlDxKxcHp
0Fo87rWz/xuOfsjS6wxNzABcktdAHuvG+iOJv8SLQK0l7vUgcWyh30mhwtpB+OdT
lGkEC6Cm3eRR5tbgnob1oZehd+YvJ0ae+X4eLQUVk/fbPt0vm8WND8l9LNt0B6Bp
zqnA2gxn3dER7IYhGEPcIOuocaBznZOe2fCriYyvZ+VrNQla7A1Lj5aaQngEBshm
OCsCGXiwQ1m/Pj2e+yPu4WsoO7PqFzcxeItk5SKpxPS39ctL4k1kWI5t0Qc2i5+G
9Qvb/2OENJQbutdLlaeoCTl9aNL0KVqGyPdm4fjlQOdGCnFvfu0XL8Ir0T56vCS7
viVUhrDk1/ur3DbaVpr4RrWZFV5nDiOLsjOX8w/vILAjG8RlsFE4ZUEhzMM7J3SH
k4b4N8IaL5+9qV5X1XL7CaqWwKtmZfBqXezMM1zmlWszR6Uekq1khM/SVzqLtH01
rxCR9I9gtc/cuYQcgljeAfWKymIl6FSWgMYmbSDJReBO8rBnN8ETbEpTQcl1f9Kj
FQFIxD2viC5Vs6hajYqe+gZc3Lls6qEguJSWcr/BAvgOYqbv0lqNqIqSEWqnVaGu
LLQ5g4XOLrPb3Y+VqZzH0uPgULBXPI5aw6syhrC9+9XmLVl8JDhmz8OEx6pSO1SE
AcGzGJfXIqoAu6WeeYlRfvmbW0XPOdUe2+FvF/twxOxO/hhdgMu3NBGtAV7TCsbN
69eonHf41IEExAaad5dUqLnky+Gk8BgA3iQJxjO7W5yn4liPQDeWthQuVoM4jjF7
g8luZJTr6VTWrSjwLuHYVMWiLAiO+Ay+tKdmOA/plwzzUZ+ISTBkaryWo0fScFsT
/6QgBP22qkoJIw/K25iCkDJ/y9Tv1oel3oOmEuZOlSCi7qILifPl8Tu68kA1AnBA
3HH556DgdSyn+25Acqz09zK2wkI5xJL46qf5eGJ4JNCHBL6I8NUOlDYVR+RpVeex
iEi4tOlrP7KciSCXTJxmYcDfMA02kC8EtU4hBV94vOTPUHavp9XDjruyqyZKRjvt
/eSWYia+rtP6wjnxNetfMxU0Id8itJ4sRWiu3fXq4U0p4H2xQ5ab4rPYYXrBAP4I
Kv9/GFT7LorM/AGckdwnPVlNtz22cYZOHQCXX8DncpdgaKTc8rZ9Q3qEp6boIX4l
nORJPEuK+ri7AAKeMTcxZ19ESKRId8PVcfcipyaIOLI4XwzjhCCvgSyQp9A5yvxE
PdI2FaPx0WTdCI5JVMf7PsTKpNjHgHZZxGFYQ64aJm5/q4+zUNtSc7jzZtODn6GT
3Bwbdb0lH8hJj8XmDmtqLl5ewJA6rZ0GHWGon1ZKwuVi0UOmObRrmpLrudL+jFI/
e8TvICgjF0Medwl+R6noGXpY2dgTe5k3mSw5XfCCcSHhsEm+owGuxM52NK+DrA8j
sMkWPE7mRrDD3nMILQvkLHXAknEk7Q33iHCYVZVGwGBhH/SwVr3dIF4S05E6xH2q
1GNYrsef3ZUKQhT0i5ThggMk1aZGw+fzv/b5JwzvUhQuVq8Jn6et4ouly5RKJ2FU
VQkI7FWB+DX94zX8AP4vRx+BNsOayxmJDkdt2nLrS1CWO3ZF5vQnYCPNCP774iz9
ndZ0P03C0GQjqnwgQybj/CRWeB/FAE7sIoZlZLjHmiLWQpiEnmeIgoJc45Vuh9TI
O+6yzkYzIefG5WwVqN9AhRNr0YN+vO735P2Fu5t+L8XcALGwJbIRTO6Qrk2XDZo2
BHBjsaYCqpRKd8RtXgtCa0j0nv58XOCv2d3c/g/IvTENYLX91vPyUy3ezASLeLG8
b+vmRo8HMWNRs0Wb1OLrLo1l9+WmrBGoH4ENdA3aAwhlmbBb7j4Pz8ogwMCJpRec
dR4gomYooztLI/WXEx2dduKFZHfzZAlvM8iNxdjOkT1j58m0PRybUQvtrsiuNrP3
kC08Z0KtXb09XMXCqC0/jsoRYpmz8xUL3eWrBMm+kNc06Sx5s/J8phESLCWI2b2i
igUNrISH5ex/xgqekGReogEQKUHljAcGDzEPABE7LsvcK72fyH70zxPvZ+u3fWBu
Gd+WVzzwDDOERzJ0SWfw+oCqZgRbnYeE3GdVAuB6Vemik81ekrQ6Q2SGzmu3dr/7
7jSSUjYWR8QGJUFs3SkCcGqRNNKJPiIdo9MLHJl60c8A4O4nUbSqnMWTFB2a/+SX
v2TLhsWtSmQzHgSgK/FLHQejqtk2eZYvvh5uH/EL7n1DzvU+nMeHopJSsId79c58
zd1U4iTxqexJBTTp3aXmCGPvftxE6/EiTAwBbyvhZsu0wPDrx3chqb3T1yvyVLmc
30nI0WERha0GfHba5kw2jWBwpKmWeDV+T7GoyNeELKWROQLT1ljdeYg/eGG0IfLD
LlNDE2QgXIAhveumN06TTBUcy0IFoSl5nvK8EzWdABx1Jm+m52qH4hEiA8GMd+hT
pqGqwkTb5FPysjwlpB1vZBHJMGQDcvqbntB6IJYdiSzDuhmISZK4K6MsHXzoFPkG
92+6g3KUYk3MqWCJ/LU56jtrmhsByKcYWrHe5UMRhOltAuS11AX4r6xutcToeFbZ
DGyHMx0YztZze77vEEfrUoeArMc4IHh7TttW4fraEARx8gXusbcN2LbEN2gY+alI
rIqAldXVfE/mRP+39Xaz4AGVpbh/9RoJh94Cgx2u1cmqWsbCoYrXRz6Cba+Oceir
xl8xocxEJrHK/ZJQOn/O5V3momdrZIGOwW0D+GskAmJrZlgI85wxndgd1was6EHH
dn5fn8OJPjlA9XsTzOvZXHd5QNPnRasInICaw1yQZALcU2QcWjz7+uoAqwzgZg6a
wzJaL7HN7uM644an2E0ACc/alHXKPCDV0RZtx85KtX/STFxWYbIg1s4UxKEmksqJ
i9o6tSeuzjiOF6x+pZDnXeiULKHsCBABpxn/0vAvFQ3bdpqygN+aIhF23LBkAqdS
bXCDRhwAdvzx26wwgIJ6wO/km82Bbug5F1Nf3EmefWauJdC2KpeRWo92m70NhYer
9itxCX++IOE7/n0nmbFFdKD7uK91mTUNWs0U4y9w5SaVUvm2bNuvWF/tcWZsXg/U
2Qm9wyZFrcmaTe+ynDg2GvDtj9AWA2wRuVmTOzhhbiMKAqE1JY/Hk+zadkz5w/I/
NAjVVj8yQpHDx9w5SeFABjtBnblLM1XIV0vHrWoCucgheCSdmYb8qACIqWTCj74t
9xWNFyJHN36/N8oGD31tVx8+oHGQpNCMDsjprJR2xfThsk7QCnGMAM4TeQEvh8U4
zvbCopRG9UmVdiVFYx2RdiAE95ewj9vOkPEnuK9cTvQ+On1fU/IZmU3F5aFYytAz
jvmWpZu/mFT76Ka6/0glgpFS8FjnQyeDgRJowrGp2DMc5aVDV3blVsA7a0DZXjtM
02XUgGKDUXEZCJ0nOLs6LfE7o19luIdPoqFN85lOZc+vzmfOuRveS81Fr9foO5Ou
yTtdK1Lk8KZVddHdvB0jsE+EdSlU5PIDSnbUw9N+q4X9qWUQ4Qf2wk56dQdLm/jj
4HwGgYCgtjqLdfWBBsVbGST1QQ0TOfp+sTaNw7ZrAtpOsooM1siF3YpXbu81/wvf
qJYz0/ShCXU5rJXe5Kz9DOAU2w3vZI4OoaDv8psx2G88+NRwW0lwKNIYgzxzS+or
rRbPgo+lg6fDxgDOxiPVfyMeotmnFT9nU6wtHfRb3T5XayMONymYJBzHZSfEOwqX
qmymeFQsnP6uTb3+PnzERPv045QbYxhluFTfbe7cQKqX7w0PGLwI3V7JOOutqMPv
cQuJMA4Nzm/4w3vi2cgCslBBE+jJ5I4SgUrzTRCh5GNgjjYUjqbwlSCutIKM7OAO
y6IZdYwLtS2MF9EcK68avCOX/MEtgLdFML6BOMQGyEXbMJnuz03VvrAquiVWRzOM
AODnUkilPQFpLlRhovat1XY9bh9Xaf/KX16cZA4mYZfFpQeyaGi4viGPfaQRL5sg
GHgRDWxzBP36x6Qr7R+BBj3Z+RgpgRMlHVxte1pGMTo7phMZJmbWdcvRIILwbv0p
yAXFmS+Ufk5f5QuKdcRcCweqijjhY9MHS2NxLhtlDZlXV77HV8I24eHvj+EblzaM
/5J8BBjwaJUuQg93gH+tK5fBnCfONJvmTcnVEdlq/I1/4WVn7jn/ojO6JNEeZlRD
hKq6BzYLKJuUIQnCCX09zHjZPr+crMOX4oz3haj6YXRAnZXVbIbWYA4XG/56sNBU
QhaRqqwgZrMQsA+c9Nsy9bACyPl+9wCgDgaFy5VHtf7dxZjZiIDEo6Wm2qtgM1ox
UNUgnYy9iAwSky1w+DC75BXAF7164qxiqKx8NelClnS6uJCzTmNmXiO9orFRGOcO
jlkOnY6rLndohKhVrd1UyQi0JPuFsx3N5PvOtB3+L31OQ7pMjPOOrwIo8t4X7uwc
GHOFUHvP9YzbDxoAR5c7DlarDUdyB8j8Blyozcqygs+w9snWAzdLc9kCjLFuMFvh
xeBVwQ295dXu/+EEYGuUTNdqMmB5whtQ66o8TcYEKwvLY13ZaDMsezlDi9H/02ge
aKj1Ow1YJk0E2gGcxZb/KFoGx56J7UBYl/agbPoeIkuG4H5J3c7pOzhshuqlY5ZW
rrIy8yMpGdefmrflQ4fEKeN3I0s1xNkk7Vy8lipG0b6WBTf6WtcYMOaIoYR6YCA5
xlRMuBIDP2THocx+kkmmSeOZLVOGfaub5Zlw0JsSaUF8j2DxKjRaW5V570RQ9laa
ymZ70YOpKcrK1U16yzc/oLAOxEdFf5axxcBzeKJIJ4ZzYEzafHXbsVWfCZDidCMq
yQI4Y2oTMKcbx90HPOnXDHRLH1HFuIs+bnwixtb4EFqHW5HmNXMT8EDeLUfHUIQ0
I9VZ/g4eias/3DohVlD7nxBbgnaXfF5P5yEM9iPtGarkXtx6hun6KXIG03LLPzZV
aQEaXJaOlIKTGjh7oQoET2eq6cIyBS1rlLGpff+JnpHuzealJqquT2wEaBoNNaIH
5jphR8uucKf5fRi22VG1CnzRji4YEm+dHRG2VmfbtFMU9PBxbEDETlPbpmiwd7oy
0W+gf84odP8nVTtqW1VuH1thiGNMCOTSGScyYte+ky1WR8LlOcfIFLh6xGCA34j7
3SjLmvSd0q3nbezcK+t4RuxsgRzZX8JCTl2V7kM4fJ27mkOaPKJwSfN22hrY6kSl
5c4VjlalW3uvFFHkVFMi9ud3h2qa5RRaULiC9eMGh68uYzx2cx4gcR72/3IvUYxl
DWI/BO/IXE/6FYTrjVvWjVltmDAZ8teX0P7bT3okucJUMNubTzsvMg6GnhVJZY/H
mW2201rvyso1qKzhXmOJBHyacB3R3nF+6o+dGmUYA8063SNrdhvMTXKa2a9LTvR7
97rm0kofFGs9jaWap//SRMzcgWxzsRk3oybpwvXGSDqfG+gRk//Rlf70gM5Gbhal
W2NSMP247fw62eUg6dxnaWa+UJ6rTK9QudgY0aBW2ELBqxdAanzvLfpmJbQID7UM
q+xKbnecUrehTLxC/2SHZI8WwcJ+Um2YQ1wTffo98DfQUXWU/ig7JyOpKAdi1ie3
7NTrc4sRO4qU/gW9lQpZKv2/2zPbwv5Kzm2BAl7jP2PocwXdk7nQYDJPyrKXMEpI
hIqtMbefwMp7VAzO2D/ZmmJgTbu7yMe1rpdv/yf9+onKqwlPy0ZmWprZGxYJD8W7
kIYhMqUbFzoNnmqgo1ds/+7BZXNCTtj811zB4hW7tnd4BaiLY6sWEtnlkyiNWwN6
9atEwg1TaSDiGzicBgZnW5eFGYFWXKjXoOK4Kum+8E/dMpk7W8L6Z25rbHC9lutV
cG+UY87Q0lYIJ1rX7YrLlGnooAbRwxf/714dUax9a/rzCPkASMwRr4RFJy0HTBOs
d0L3qUCdu0d3vqcczGETtdVNL0P1kwauotrU4WpPwmOYejn1UcTWiM31eqDp8FLJ
L9inNQiWYrgKcMVlAqNhzNiZDWJhPdgYojf66bCs6gqRWDHyKkkYh4LiRuU8NcsB
oDN1pjKDtmFCezIqIOiX6pQxk+nXKt/PS8PccbBi07/TdLLKRznV5r1U8q58cmaJ
zQIXgbt9TfH1puUE+M/uRAuekJOg0IMexLLhch8P/p1GOHOSClBQxrbQ/+UFO/CS
lP4kcbFRiT3/v/lCKRNLM+Nc2pC+md3R0GUTBjP/kAJE6M9EPpjBuCSFBKT4s4Tm
meduWsZwyQ0Wi8AU2NY4qQyToLDTfB3OPTSbYsDetWOzpehvQbOdqP3NTqwJ8dn1
+OCgt8UuygcmK/0m4TN8iiH0pqxRyebnwqFipLozDL1FS9kaFeZJWmbE06HNK12J
Iug2HjyijoMdA7JtylWnLnNoWHkG5Kg/zKTVBmcPio2RVOn1693S2bQA6L6yaFuD
8M8QZfYDSv1HA99r+0S672ifyQx+zFYPTIb9rrZRIiwrQ/nc7/gz6/bPDqNYNnzA
IE4i7M3ocd3c9u/mR3q1K+hbL4sMx5m00VkriKS2DAfWrskufHYdOXB+MtUm4/Oz
j3tgqlL4QFFu8PYmC/VUFbssnm0+8msT2pnV5Cd7Xry4rEcwZRHmT0GhqzOx6tKM
lRTGmm62RLsecivaia7PiClzsx/Fn2nZ+GPbAz9Mmulf8UK5MBBeQhNsPrSOdxDy
166Xdps/wJ2RNfQiF/Gfl1UnZ2YcbpTYI3T3oG9r7yQ3lMyC3myJvAqL+i5WG5jC
WgbZRiOe5F8MfJQ+ZagZcNIvpnugOlcrRgpk9YHN2+P/eLyqno4CmxIbPU3UJsi+
Neg/jBB9K9xZHZfvEuFrbcFQMsU6Lp7eo8O6W9yM5H47JklLnJM9Z1NvDc0T0yws
35y/odHnmDV31/9tmktMIoOzV+URjyZXyXcxAdni6E5m1/XdwSODBY4es1ftQ3R6
p4Kc53XGk1y1P7ZTVZP5IElY4zAr0efQPT4/C8n0vrIsqn2WkOIFdCrDNufZz3xx
2oHa5+Ecl+vIlrj+rCLFrsmt3VFHZC5rHzlBJMFVbg0SVwaprwWe3eWAWWCx9Jmn
blIrodPyqFZOyGoDcJ9TV6nhMlzpalpdhZRWe9EDUPtLe1YgJNRH+XbAUzDv9O6I
vNG5Xis8XaK+bfEYrkD2D+SZjJfB9Hi0yVOuksyRb17mqxmQgOW9G0CUddMgmgWJ
9tK8Ckw1jRuj5yb4ash4K3ZWv/LQGn862sJSRF/AIn5du8eAGH9f7lUkCvck35Tq
Hk7bfeAK7Qfr0O06AzGMzSCuwO0RejNajsvcxVxAfQzRRWSTqYaXRfRxXaD5Cn6g
kF0VXU42lfjbCkkhLXr5UzFkn29XKM+BX3U8xUQoEAAHu4g0QMZK6c6qvJUGiAYG
shp1BqYsVdkK1DOMOHzd8m0uM/qdO/cWPGx6vkPFEeXLT/Ej7L7IdAjayDyDVKgy
WdJ4iuYe8dWdrzw4q0xXltNs2B7PdPN6CfQiWjOdehPemqAjtXPG/Jy1REunZtnd
wbNuQJpY5SqfaPsEbNb4qwmxEGAy5bR6S5YgG+g5QV/Bq4fz3IzTRKG8ZOrGjyfc
3S6vl0EgGsmzEvOa+6khqWclg8XDN7yn0u5dVbfbqYJomyrcCrGiHYe4kT4WJB1n
h6s81ELyZl6+WRb1/2hPDTNgk7ilpf4JHmzW+Km6DTh7dCLb+UwrqgCfWnyYQtnK
a06Nb+Bxy4al53kKzaWXCpWlM8OKFjWp1GeBnJSyZNBjO6lp2I7B/kDETPtNm4x+
hj4xLLwWG6igL/bZSw1Xab79k1+3Y9MgC9Au4U+V5ZpPOJxzIOS0wE82qf5R8E6/
hFM8cJ1aVuPSNIXUZeWbdhiAW2XhGXuB6czDr/gcQNSoMC8BLYtn0XAbLG3bLj8A
DVkH7jBtmHZ/gsaLMK7awOqzSeZIPotOZ4TOGy6UeQpL3cz8YL8YXdzJv4dkPwU5
db/XWPhzS1Gqz6Z2l2/3K7sfgxfPSjIoJGsD++mmToPpVZYM7Lh/mTmswGkjTViw
02t9ejbedNMOuBUOaDb7V0Amte73KlgWtLUKgZ4BUNPGmic9XFGyhQaGVniX7gtZ
54W2eY8utProGRMYMtcYmSFTnTjyfzAu3OlqhOOBsBtI2LXkAWegDsWWFATQAbvI
z6e0T5IPgNuycA6H3Z0TU414ROl1WvKqd2Dqo0pqeyUmbwkouT4/GXn84S+biMZs
UaaB0lcsBsvpAl4BiZCBPa8485NWY01FRDlxrWDQTnwpIYQO6olpEPFEZ0ULehYd
EVx07GvVhp6qMQ2m+gcLMM63fOHjF6t19cHSASvJpmGYah4Lzx4eH6l1+nUViJ3X
1HkhJUfGruj0vGX81vXLDU2zUZoC7sDdp6u4QmoX8y8WAdyLPxltIm8oW3W3DTur
/7+3Y7Adqmpqn3nVX1mImBs4v0x8RH9u5w2Tk4Z+otSzQiRCTzxe3aJimpU+fsuP
P+I4eTfV7EH1gx/NQLbRX3NAZC+fOqIuPMCidTwsmf81m1Ih47ErZJT9qP9bHwFd
87/0z3fKcA7QFFj5CfwbIZ9WscncQ5ifqSn8+qgE/v6d/HwukkLDVfpL6mCnlkH8
msWbFN/4ZtXFxEB2SORs721clgMsrJ93F0y2c3totFrpujo0AFA5K4iGRwmIHxNO
QHg1raUI9DxjDamuOeROHphB/yVrJFcuCHDVSYAtX/MtQDD15Q+xdzNLNjml4R5u
qNiJyczeD9yfgr0BVWiyszrlGA/5AbhY/CeeGcWAzl5eUv0x66CaSv3IHiBrCx4N
mL9NZ862JlaOWUsIGXPdA9GlWoUd/9+xi9FTlp1MJjPvaoyD4ypnqN3nYKCpVuk7
v1YQmPFuKvCYeyqMYr5HNIp1vOjV6vfiDejA3Czp1VqK2XYXl43z0c82DyIs5JIw
0PMWlvbMT8Lpi+IwZ3zYxmNwWffC4IamswCE8jO/viTsz3Bc3W4mCLSyKX4UVfe1
rvfEng4n81LmCNhlE2eqKfhchKs/4UuvYE7YYJ5zcpKha4dTdqEeKjwqq7XG6eIR
Pi0qfhWaJnvTDvxCg+P6uTSEdHUdV21hkxUjK1jr/eKDK/+L4I8Dm81NYGPQNnH+
f6nt1jH+9tozbnPJGuVlQkP28nMB5sGaWq4jsoyPni39rcq+VQM4hPta40NlyEYD
4Q1r1G92hizkCh94tdL3By+gLdnlvOOrBPbGkusaMChSALGp33MAo11DMsiO6o7x
B0KDK53Ids2WwF3RBCWZ5TOT5D0L6AzGicO9YkmJSbKNNL2QD8HIRrL29pGjrILf
TMFklf2gAzvC8FwGOVpmq25p7JHgpAdvVW/VJiWvB3ba3k+jr66y/22CYuYd1ZOZ
PQdRpSgCn2CJv4fr6r3dHNBRIm/hHKqIamUa5WAuVeqHRQihnKsI3u3LkdixpQzQ
idthM0c+BzRQWq9UyBvCgp57Wh9iabfkmJ5I1gxNHpJJZCbSNXhXNo8sid63ugC7
W2tb0emdj4peoAuqTleUAgBZK5+qkqfPpX8teUFOE6k7Q0Jr8ZQiQ6JE9Hp1NRpG
L/I0ccGKqaSvuMOGi+kUcESkbUqzT2So3U6k7CR5XTTlXy50bb2H48OU9jqn5u+v
22Lp8F8L/teZQMfMpRvei7KBhjtrrG9pwbt06FARO1U9lZU+XpN9KZDGSbFkE1NH
/AGcbDeN7m1uFllsDl/dcaTQZKuCKWbTsAwxjDUMEmf9D6wm2y7i3qowSZq+iF/o
c0ScanbqrALFfBbPHUD6Y1DtT4TCbato6nLR0LwMEb5+C353rMluEMOL1gasGqU0
4BGekjCPF22eoY3OcPahX4VDEYnXfow5BbONFnzZEhRXdIWAvqM2SJq+gOuzhEIz
47AnuirB+ClSrTw14oTHkX0AuHrBQ+iIFZVO7EanlytZfG2l6Dlhd2EQrZqgqjBq
DU8dlci1vfplaGpbUr91yavPaUg/zludjkM4/wehHcXBNv5xj6CIpRrvAokEsqET
vsV5TwBQQbg05UA2swdvdjwrp4ZYYQMKSa7oKyC5dIt6wQjHlT3z6Tr1Mo+mdR3L
vHRtkkrE5ppuoHjl4y4A2spy4Q6bJPvVA1f6/S0qDv17+d4rLJi3n64JiPaLXqhw
WDo1Tf9Qa78Nz2081uqRfTsdfXDYGRddzi2xqokWz9shVPXqQ9D48Jl+b0YkxGw4
rMUt0ngXnid99NVFmMhU4p3yBM9B4+wOe7+HBpb2MhtwWKA1hKyfOLC5EWWlweKv
pmlPlEhCbQMCy+Tx7n/UXptizyrFKy4ZjJqv2jKq4SrEF2sJrBzEpLRPM0TttpaN
Zcu1JPOhWEeq6cljfEJWpLX8YsdPxr59y/mm/chcTtw3hIfjkPeNf8GZRrzyiYxd
/bjBobrOG4BPKYEEiUu7SocRiHCOOz3mpSAY8V8ou/cpyZZdMoniK8nO59r2u/hG
eLun0GA9UVa60+tFGx7Z+K6TGNUuGF4Su/yFwoqRwdbqeAK5eRKPLtMfvaSeF9Cl
vuv85NprVPL0wU5hyjk8CC91s4p2pW2Ckp3LWoLoGvL20QDzooC1rA1pC7Q54LzD
76bTuz7ByzemBl0jit5lvO/bBrxYm9O0/Hl8gmyAt0r4OeyTKqeATRPghz4wjDmv
hSR6o6I7RmK9nRGqROI/5rvKVLEZjv0NTU2z6RplyNo52t+wc0b6Rq/Rrdj5kV5O
zXFNTwZRaIGXTRq5EdaPchty55nXHAYVOxLEriesqZbACKJSFgmHuBedEU7aaHGk
wzIAZ03GwCDhi4m1dc/1y8YnvjxN51HHlxnGdEmqbWyrKv8hYDhp1gPRlyzzfu/x
IVvcs7d0DRWBCUamZLEyM+RB/+gWV+EnJKOrNpE9x4M/QjrHpitatji0lfEJyn4+
jVbrDKbhGde6Stw8pNnFLaqSCU6UnCfNC1iTGvETR4qm4tw18WN3qCHJ36p2eRSN
1OGrGxa5h2bAbe/oVkE1s6arSgoK3q07JhV5l0VKwyMNH+NJhHAsnfJ8DzwE91j/
lOKUOnXgMEWXLUt7Oiauhsi9orex60sQBRyy6BY6Y5PLJMYDxpzZAMiPVQ+0aJXb
FlUCng20EWDnEd/aY3qGR1ubs6X0QntIwffCQUWOh+Vo0S/MKWmrfVZA5toZ/nzu
YYBmRTlkBA1SIqwglEnh+C1P8/D6t4RAfl8cKcfBw1qrfPJnDQp4q/we1btLzXAR
Q8E+NsDc2mM5RftLk5/exnUAUuPldzlNcJIbjQE5fmLARn4SOxCrSaFh5xLy/D8+
trbbj3hKiPGuY07q+OqMGcRtVq2/Ore/KtzARdyebzf8yRn3h9ujnMGGV/qxghnd
xVhAtyaBPpcwmQjbNPT1Whw+4Bnyhlk4cgWg2n1bWMck0Tpdo2BS7LZS53dkbb99
xIl3CsUdjq7/+w9DNz+BtiD3UAA8E6LD3AqtAKPQ885gKEPyS2aNPuEfsKoE1JD9
i62KiANyeO/M9ZATRIJLnm7fznV3l0nui6sRgB7kKxkw/2iYQpA+DjDaUk1srPTK
bXwDBBiugnv+nYg71AefGdUkrNJ8g7Yz0tsmZsXSdELz3mbogG2WheUgbw4eI4Bc
jQX4E/kc0X8xor3VzGXl13QlwFKz9xmufme85jgBogw4QMrdyxhBAXhNmAFZysy3
MeXZku0WfIfFsECz2dyvqDU2wYCfxr2ux5nNHQhv2Pe22PAaisvT2Jag3rJDpySX
jKdxwHrqecKxJBCP4d8jbtdOx/BwbBx7d/I8JHnzSuhIVOIgZ8AvNk5qBInsLBTo
Sa5E2Rfp/hlRh0wMXJvERnikKo33TELZhwkcU/+yJmMkgsHLOqzU/b1leEAWwWHD
U9vN5wSae1vKFIz0LH6q+TTgf/g02mXojB0qNr2Q1C6rz5/1HVi3qeI1waS2EQCl
NWmg3AOK+ifo/M7/HxXtS1P+VJqKaqLhfmloOSgxvv9NBDPFiTlUPYE5pGE7n9Uy
WVDDg229RAPU0gBFuQsmc1GjVbbhAQm0+E5crSDbuSXpHdXBxXCk5nTbGm/m3+JB
I1O4NMVoANWLgYYKZen+B85z6IPErvHzb7putvIJfmV9183kKvmV6MbGOhVOpvti
OfMHeO16lyod9oAEXKklgvVJX3DEyf6wVn3ffLx8VZApZJ4ERLLk2arrE2EclbhF
o1teZEH+giR96Wpn+0pwbVMch/EC8JhQqM244U1fpQJbgYR/rbM7xCd0JoPd/bTy
vB5PQA1qDubK7w18rRcHG34N3ul9bBKVGd8Op8As6swFSpQCLTLc4kCGA57xZ++f
fzpF75RIkIuQ2GEpz3x92d6IKFiL16DdypTh6VLepwoMaoZXXo7bHbVS2mdozrKN
G4giaP5p9iz6NaKV+xVH1EDkweDLutRUs9tX+qDJRRrAJvCBzDdIsCJhz5hi3Iqj
hTZRHklp405HUERC1eWDFHlpY8Lz1RmW4D2LyJJUO5wzkR00Ku1gbihG7maSxbpj
RT6W+vDXCa5HmCQLYOfKo93eCveHfM6jlGQOrQI1nBCGba8ELUGXTj3w6RSE2eDD
ICjNPlPZBkk7VeE1HhwLpBo6Sk8FccrhoW2o31gebfTcF+WOXT1cBGdqedkftT/e
MXup5iMnJsUAaM4LyiN1VpBoWdZxxiVQdGYeEaJSGDHOJ5SR14dZ+/VumqoucRzt
J3ERqGYUTdyxl7heSyfkOBLTKpuLAdLSD2kncvOGfb2PjJOihjH51NoL5PHdNzNt
B6hzprNhLcSeTId2QlgdAroVe+ErLkZE+xBIneiEODdv4PMxDFxL/eOrPXxgmYAO
t6Lpnwostf1/ktHzf6cObUGpYRAhmr6oHcL/xsPtHecanOOERZLM7DN1YD9OPKyQ
+RVcogT2Zy7hplUOJFaRAT/vuuGmO44jsUCl6QbqGr8co6ntABBG71iGhWX8Fagb
7JGB0aYXRq0FJUidqW85YHArGDhGB9tnlhah/gXrdjw/njxmzZtmDL7I/bsiCHJG
eF984jlqIS6r8J9mzTJv97Cn7ZkMxBlalF9TTlF1+PBiVdiYaokB2iZUs+lhmJ1I
cM2cj1P80y8DDpYR3nwZBPMX+r3FwLjyyJ/N5asSKGMZbbaAf0gDJ0X13guHoyn9
xnpq+nUZ++MKeRVugs0XmBE0rzOZkb5KoP6aJDr5cfXbpp0xipwNn2fn7IL9UpRi
/kI6iOXJTaXbsnyvn7prfJWkrnXEjS+CtsQ5NaECP9SYs0h+g5bvbvQjCMlZ0WyT
K9WfwldC4hoLL1ATepvzaGhzN0igbAkC9gC5ATNS/qzHX8mm0rSRS0oInJYxZJ9J
dis05bQnPQihjDDNlOxGeo3X+CNiz6JSa5NjB09jpces6l9yxXyg1E4fNHkpd0zo
snE7bpaR7nTyNFzT1Qh3tnhBDMxSr/8qm5IqE3dKqGxqVwLuZmDQE7tzuzuR80mv
I94gXaGTqDYTWVJ2103VKVM+SdFVobhlxXfkEdWfT9R1oW2clqrVVVAtZ1Vlsf7i
ufoSFWElWj7AeNHdf6BmkAnifUK1Rao3G8r3bSzLi4oOUCtPgCqstX+bs8w1cdK6
B4U5picheBng66aJnMDcbqxT7f7PEV4kQAWhGUDMBmj1vH+cm8h7NICLGSUPruvf
+kxgkis8zHkZGhDCqXSCc5JsfVwHb8YyQ4ccKO/Z+f1XHjQHNyaROga1Ok0Z8HL1
yeZeV4QFwrmg6pSUOBjCo41ZfKKat7dfdsVnkw8Le3zwFG6D2uVuENvlMJcDN5Zl
xybCIAmxN5ekgxfWzQmiBTDcDemvn5J5CEsul3wPo2ehzPzBfgx46jJTErzGcKjM
GQ7u265XrBOXOn8DY7E2yY1WqZVHSZrHAYlkmnz1lINzORhLdnfLRltqF7B82GWn
/NomFtjNuqkg1HVFLNf6BK9TsEwkF2yYVcpU40FkLEuORJHXh7alGt0FN9/dHGb1
79jRXNPZjqbabv8+WFoskCmx+FIFsZKhYY9cej2mPkdj8gUw7gH0KPxzD3I42swp
Pnu4Q1E+zZc1co65BdVYw7K/vuZ/ad24tLmLvxrExm+KxwRc0OBmyJQwOaq+p2jZ
3Qb3GBU4xosAXVLNtcYkALIum42AWS6uglB6lt/cNujvwc/ME5IdOZdzuNuWVOiz
zAeC3sEFJlddLNg7v+8OOFYgXSy4m/1g2N5B+1NhjlYHEWW7973LreNKwcBATqNB
CPueFhJ/YSa88xNe7Xil4oksvvJ/w6+XUpY/xt77kJIImoD0jwO0xe/fFaciKnf9
rROj/W4RP8oxUg768vryGQcivZdMypga1SJjtPD9sGLXkhap7mz9QjZYTlKY8jrX
257uzo/fLX2LZGCl3fJgiJ0YaWwBHcPJazJ3dnN9XBV/n70SEAUTADnbEEbIIhSg
M+2c/qQq5BDW454fVB01kPrjcapx0K2jlYGPUY9G8v20TVG8GTVDlPXun5OiwJ7k
txRRxjRK+4B+PaxWArdtSFxvWuWf2P4UV+bombnKmc8L0DX9/uwswBvqS+r3bTHC
dbbXw/0i0Eckl60pQ+dhyvrnozCzxAQwcJ51Sag8xaUR9mgODSEISMtVQb4wsXBy
N2//s9zj46bcxKzDn6GaJsxLVaQ9PWJZSN4gzWgqwuYi0lYl72tr37COmEG9G9TC
mF4L1+3QZ5gbzI5i1JvNdeVGHtKfz1dtijzY1yJcOfbyaRLDIK3OqeWZbYmYH1bw
UAxbcUQMKzEM9YrQJ9mt4kK0mp1l8jsc9jFznkKvFLl9qNLsJTmWJT5/0STcpEsa
YYvVIkdBb2ZShAR7idSvcSrai1y5wK5qiZrucLPgxzHTVQtjdoPsLsGiHTvDk327
N83B2N31hVgVbAN2GLCPS/z+3eJksPaGzs6FcrUv/1rgKIFYV4uYHvDPH3qo4MpH
0ZlsHG1JXV0CKTMCku08VrP1LrA8p1LPrQCy9G4vvhkRnVszwHKWjRAQRrq1SCyl
BUVzNabCBPaDsGKOCU+rJgqeG9IIWW4j1k0c532fvXN8TOgaEjnJ31FW4jIvF/9t
sLzo0mFQALU8Q7JlhyKeDoOpYzfGHswbXf9mcrd68h6QAIAMkLPlSnrFhejDD69n
bnzF+MwEeDRHe6VuW0NnEer0Jm3aec6LRQKwQKyFrrtIytl+vVVPehH6W5ya5eXX
D861mytsJA58cnYQU0EAeohXBIzAfe+QSzfMQth9XosdQljuzPZ5rUwdIYIbklmh
v97deSmZZzxZOWWtibYaMvgzOoFy0PyF7hnqCT2wQ96F4XYuwxE7sN+9GvrmzurQ
ycZvf+PGnWCJFYWWok5qOEr2oxQ2vKt1i7xu8dB+wltVLzlKacBCE+Wb68bMrW4Q
3La27vDDfoq4WESmO2Au77jfDNU/R840JpUfcvofbBhgCnY8ks7uqQcNq/uYT3sS
llSrQOuC7s2V0MFhbvqiZlc6EJK9GpMbl7lg42NAsrcpSm3SwB/LFDIBwifAvkj9
rbviVxfGbHVgD78hacWaFy/gDq5p9zxwmDL0nF4rKsJOMlyXL/DvysUClU1q+d3D
m0dwuxPhCkx0Kz/6baCT/vvqwjI54h5Nw2jGdxmsqJff07fYsABnZX0YksHikTER
P2U2wFhlY1l7bcXQAb1CH+VT7z1RToTVBLYagX3BvlRfTiRHXIq+GFJgK81BSyNW
V8ovqp2dOtvhaipXteGUUXIk+KyJaptqVpneGMoJDQoWay5t4L6d8iR2Q7W7h//d
JoQ3XRhHAK6mq7aEZPR7PVo7JXmidzlB3bWo5YsKqzF3GS135ZaeMGd/sSRbVmLg
Z59yL7eJ2U6leTCx/skNBe0ihxqDPD8G6sxgYnF4JDvb5rK3eS5mh46J18vfKTLU
GqYY0zo/5dnbaQZSyyfg/ozgM85Pg1hyE4GlKlEhHMbk1Lub/cIH+oB5dV0lpNxk
89i9HRBWlU21k9m5KUeWPTpf6J5mSoMrf3QA308FTlTFj88WIaDbalukgUf4V3rx
uDg7mPnYh8pMxZWTgpbB3U8hFnopcSV6Y1FCSs5wUQpLJyDeMm5I1d/F51WaOYCh
jFpF8Q/jRN7ovlKt9CAymnfllLCPcURKk7g6MOPHPpJpy+8Y8bP5ExlUN0MZTrGY
OSy+TlrCLhizrcO3kOg5BXd37Vd4d6gB2ptn+MUJZzRb6P94Z+ayWkwW+mjBR4Mn
/Z8huCmv3LEs8dIVgRNKK83y/IbJTTszW+WU/eJF2qhB/KYqzJylmhwLN5ZBsNen
IC7QORkjlZXSTJAwO4qvmUBlgJclu8Q4uBj1Yl+910heAuQPQ4DgBEmO9NIsUpdj
XdqxQcIVxOZRa7PYiuqPvlDO1+b9kd330YgCdlHKr15eNlWePoWhtQpP94g1YTwE
lDhQd0YFqLnZbn9ruRGQc29Q4i9AyZi2cZp7FKl4VNht0JMRmbCbeWB48JqWWMFs
uSbjzwcx5JYJYtO/WPKnFoAqks5Ef4FBoJeNr4sJlAmCGwPLcl5ZsvMkUI/rZ59K
06IyvxDGx7ZSsXdj1pQQ/nrU/0Ea790zfXAcEIQ4n27FWIyedPIzrCafrfaJzfwj
3uDJa0NSO+dXFt5UNLzn5zjDFuZRqZ+c6RunyWodo8+IAq30CMUmh88L6PWRt7qi
l/Bkc1zl9KJDfSSuBIQMnySrbSskeJXHyQEO/TQk3Kf1b4a+v9KN1ni1q3An7avM
XMfiofWAxXssL/Y3mrDPVK6ItpX5ukgPCYOj2dY/jzHBwtrhIPR/YfFAr6weQdtE
1bAPidW+vJx1AJ6FMPAbTivUSpT7OunkqH/zxry6DTLBb8CKgiACCAx+Lf+QqpWZ
cYa7VOq1JHyVZyDkrx2S85wp3h7U/4kA3YSuAfAFWZRXL4Sb0I9QTeCFzHVIz1zf
q/OhxcL5zzVAujBuvdX49bwAzsa+XP1wf51fZwW9sBE+tlxHQAdwMLYggBAb/sVs
8VS2JxQDlvY1855mYL5k7LcyM9VqiVNkBK0R5Nb4AjwgYWBhQDSeZjOVF7oPnq8U
+TeTxOHAn9FsaaSt10FGG533QMHUfD664xe/I8O9mtAJZAq9Ag2JR5obBBjFspti
Y6r9sFsqoSyebVwi1nh3m6aafgDOcAVqBPaRAZX6CwiIpPrLCk3dEWK9sUX+GU5B
NntJZUJ23xZYMwm9IsZrMEcUbyokp7V7GiMqdRwS6bq6sGh3Zj+UH8/bsjMbplmZ
EbQF31mfRCIh8HKst16wZDmDTGtodGx3GYTqlsu6E8bY8g5U56bqPJZ83BIu6hu2
S9AOImKggy610C7IbIut1TDCeu2Kj4PEpzxQ7GN+DdG0PMcsPQMmGKExgc4MR1YS
jDv38H+3wBLMbdiqLY9XzyceH2t4p+NWaj4hPYkpIBOlnevuVcmMAT+pqXLSZXIG
+SYUCYI6+BZGtka96YmEo6gWcwMqNxikgMVmXC1CxwyPyrRohFRj7I89EK2wHtX0
AKp/LyihOUP4igTuv7FQmCzG6uGMNk96kkiXIoOLDred+Mu2tMTosYyCc/xgdLm8
x/KvlMP+G9t/fjKsWBO0focEgJueh/7vs/l6+G15TNsjHkW8JeX49HjUFbW0wH1a
DchFF7Icbue28MyN8lwnuy6DKszu4/mxxvRM1HYA+N2587xYZMPgYlHpmM9wG8Iw
501Vc+/XQUm+cGG8E49jYyUQefzF0kM36adlhQDr0xt/HFdnHYZf7KhefI3XNu9t
1cXkOnnC9Mkbisj5HxgdHg9gJ7HJEb/GaT3Z6nV7ddljqRXJcck+Z4UXHG5IH6U4
ODcqRaaxTZZVZh4d5qGa4E+pI9hfJi8ikyfuePz0UibRXROjUcZ9e4fbTWM4m34X
lV5LOoT5qgiGcmxpk/xARpebfGp+6vrT5+lt9VZW1hVgnoyUbSzAAoyQbKJ9LETn
Z97jS04SJ8rS/YAFAo5Zh9nWBF+yo7bZ/abrAzsYEehLF1Jap44b97sHp6jEn7Bq
94QV2tNguDkhkcqlm1N8JS6/k6hxlTN7kGLHaTGyLZ5zmI+K39q1Fu6Ac3B+o1jy
R306RmklNHF8zapr+kxBOxOOeM6qWXKcihqvVqaxjfdGO/tkuRau0HmF08qIcmNC
+ixdQFFQDEZf/0e18/2YYkK824IbtRDvVJUeqewKmqbCNn7hygHMoVRujIc5wlJQ
b4HvakzsgG1wi1NuMlXGZrFqORW9n49004/USdSBGyPNup8rTaJPmoUB+crMCB4H
oaz43+UNIdxk1lBkoyU7WlVOMr65CPW1ezq7dDpdrcwNDSEZWiEGwfGNH4StXjdi
ZE++o1yRJLaCX2GwZfo9UXJCWHptZrSfUAjmWlkdHSaBC50tzan7yiupQKs+xgiW
cQsFxcYT0GVBO60KTvc5NmgktRKf/bKOIldS6xQZi6lvHni+mkV5mGf5nKzcRHnW
4HSFObW/z27tJcCN1oH/aq3SgYggQ2rbfZpcDpe+7Xk6rP1nDGcmARVxk88AZVhI
FKRWbTAhcdV1SkukdM4Cwwp29P0lHy0OcOr8SiZOz21wg/J0hZTlJVanAj3NiQnh
pLNXE+vMBuajbZRTCmM+EGMSu2AYYGJhsFnnpyRHlDi7RHwOg3ALlsGPVEfoFB3C
DgvrRt4g7YkHgWNyIPAlmgLQ+DRsXhj2sJ8/0AYSEy2g3AE39+ap0iipB6Yo+V/p
LUqy1f77tWvqOuTW5hXkWVpOnKQTeU29OnHQqtqGn3SwDaZVzh4leG2RB7z7VfS7
M2ZiZ94xbZ/iR6Moqg92xUWJnzU/K2Ysruue0IC8Bej2rojTaoGuytQ4vUkRM+R5
M2it+TlxY3Yv1vECoVDH8JYz5an8cALAdfZLHb8HlQk9XUUQLVOmhnSTNBPOH+W2
C9bvokQjLZ1OM0ahUiO8fapc1BAaHCixap7IijLl5I1NNA5b0QlBsPe/hRFwLnL8
nyGicVKdSxsLNK0AQ3p5GTskVvmvDKq9Z/LMx3bRPlcMm6g6QWD1ayGxyOJCNRQG
lV3f45VGfyzECBJmTbOZN9NYRVOaFNqMwKLc66EMsGyYID+gkgp2el1Lgebh67Ht
g2tjJtq8Ez0R5dXI0CrGVttsuy1LHGEKh+CgHpn4HlGOX7JP7zZoJ2KSPlhDeGm+
R3hBf2CH5ZPHqVImq4SP+I7lpoXm6R7v4EOgRJi5+7a5VNJ4dWnjmDEnkpgUTT1V
BVSIZEGu+eReYwN/gJ3T2OnYAs1jHxcuzZdfgu5iwMryGOeyuaWPaHE5A+bNNIOf
dSuty3R2lelkMi6Hl+FfpTaFkjiQWEHbHhm2nDV76cZWLje8L71hrm/C9eq3ZM9g
x/qYiBhwiGPcH5lSpIAeYiQ06DIe/56GvNwuQHcPewBOfmX0qqYmz3/fyZ1PuAB/
s+6Y2SKiOJ0ox9PAYwtac68Eh8nYVEbE8zvEdcbDns2NH93SfbQ5RjV3XHk9i9iO
WXSYudOwx/cy+zsmMJ3HKoDNo5JBpQwThd1VGfTE8Z+nwVkgAXZwJHE78iGDJ9um
nwen6HRDaRDkVPQSwlJrSv9WJ+aGXTQUOhUUzUuuatj0xIxWbIHucwM2WLTJjl1e
hbp/Bu3J0koF0j7OivUn09DJyY8khNGMlSDjH0kDouDYyW34Kw42otmZHC5uqydh
iTlaars3mpKLtAAR0rqLxEAIMR8xtdrYXbFH46e0eaOT/O5s8EC+gIRCVu3XxfRv
1j7YlfI5gYOArNiTjacR0GTSuk8NtaElw9e7EvftSnAeeimCefqI8OAGBKEq+Mo6
IWb+S9DQQMtCQZFDeEVdthIcJaQRFRGJcboNDQjzBJrIdUQRcFb8/zhHNUe76pRh
ml52sthi8uaApycfNfYOi2tJvTiDkPO86pk42qSaAI1b5B3LF94xkB8bo2CndLq+
TaUUQ3DFIh5dRcaVSA5xc5wo4PWooJ/iDwBPhg9dHUh45Csa/v+TQ7C8tHSfy7fV
D/BO6lkG3MXCkiS2B0PUka/VcVw8O/dsfCBbMuxHWTUenggar55ssVYWEHQ2Pl3b
wgXr5FQy+flverFdBM/F0Wu4ltjLfGlaeinXz/Y+hpeIZvArtNwW6qyzomMwlJ55
WYwixGIWPaHWBzDDcwmsnxtHj/YkWZ0Vt5t+g5jD/1kPRxBvewQxrI2GKE7nFZj8
2BiM4AsoreVfRIgMhVPKwtBLviyWZnrQP1lUQVINLurX+Av5JM97rK7oXygn4tVG
hN5NujdPVxG4/XHrhn3UUokADX5xu5ONbLuHhgKjIruENuWehDL6xTBTds6okAPL
7t5i9AogsP4Rt6fLtJtjx4CilABIVYLYIOA9Od6L7/tpRpZpP9oPeLhtiyJ/xnWR
6E1OhxFyzaTvh180Bbxy9UogAWQaYwTXsmtzWccwaZ+FbZ5KbeeHIPuLGbhYmvsZ
mK1HY4M2QmOni5QXkE6gU2+voNZsfHFTT1gJUt63+7Gdj/+pzIF4Ua+zGL1NPVAd
2uhQreeOxBCgByD3hwXpgfKhKARFkPlPKcyc1rrN8bNYb5CC/eMF5/qTCCS7mhGG
mvxwPO8CvW9czV/3S64cm8HAO47pEM0Kq27BLlg1h4ogx52JPkFiSbVzBK4TMIrt
TPRDjc7uE+AfA3Okf65oA+aqXWcqaUeyWLu3nFja+BKUvaY3M9VqDQ4QSZJ9qd1m
lJrLVLCY6pbSmppvgVeJrADDKRrNe0gErIMy3coM13qSqeT0v6ahcCxDSVOPfCXW
+dQWbrsDWxZEeL913mtWrVlJu+ZwQXcZTgQrf15xCZLSjEIo9rDne8Lt708n4dp4
3Uke/bkVkm7P5mLVfVLgF2bG+SVhwtmdWBR939NCjW2otY4WY51N0JMvFhPXPCuP
HzZeSIDN+iMDJJAws714yeTTIPJCKzdLgu2AE+ixFJUtbmvguyysDGfDT9sBwxmc
cxTTJgWjTiGGbP2dRXG6RKN1x4gW/USLAjToD1o0fBaW6wvQz4HnxGyuSUvN0nwa
JQkDr8w/hoEUvoD6dSDCRN/TeIRs2FLLUDKgR+HjlmAw0ialwRaXxO3zbKW217Cy
r6NpHFWHKU5erMSPbZ7JCybLw7yDllCGhv2JMx9UmIk8WJrvybZk0yTqsf220w57
4DcDGGePgLGd/T/cIlp57a6A+rzACH6h36l/USgFyPxsb9XwBqYPFtUEmkAkxn62
I63fLH4NnPqRGo9jI2BXFG0VehuZIcxh/tse+LJ5nDi4DbtUuaGQSYXNOiOFazXK
nJP9+YiyatFCuPe5KP9baPEgkwXpcR5O/DXvnmgvMl9GhkMOqciLQFPuhhTSydFG
TEgrno4ScGZnWpFaznzmOa2CB+Iu7TsVxC5wlCUMtKeyavtOA6FRwP6R5FHIiDnh
fnMrdrlpyPPJcbLI3kd/CVlRj4EwxPazv/+9jM+ugbmspTVfbbQvj72XXzHTE82c
7HTWDnVHbxQA7QHVespihUpsIW9wM3ZFZurApdaWMgE/n9OAriVHPcBZXS+EC8iw
61wju9G0v0QXh/gb77fH6LBVTVxZh3QtuSY2WtK7CeCiNZ8Rngn9JQ2G4vCCoQVz
GnE07unnZ/AF6pcOdI1CRkivej6P9G+gIRyhRNw3BEtO/Lv+zkPHdBCeuGfrFwF+
8weJ7FpQzbhbKJJyGsq/8jYzcPWalQHB+VQiRXt/kLrjd8TuecbjxpKwY4TEYrZn
GpbqNGCKwT0TkxHkWqfs1giBJiIDedc3zsFfanKC/+k1GMAvTOrUd3D6jaxKA4Qi
NumTVIF5bzBqlv+b1zhr242BAYphI9j95ZZEL4L+t0PdFyTXA8A05SlS1tUqpWrP
69wJBLhwWjnfoHc3fyJcwZLGWswA0yxgMhCJk/y445Qndg2EFGLveDThDP82Tx1u
PfI3C4M8asoU9/nuhg9CrdPL1Ti28wJBCIUcj/ArmJ37dLo+fTrvboe2/GzcxjBS
uowmG6A92l+in9MlXfexu2wr3Dk6Yh17/PtHRBDIDvEe+5QO0ZyGr9uPe3krSqsh
+DlP/F67p6R/20CE6GKz24miycgY1y42q3d9CHuhtdV2nnBtutZbVWF4SOZxhQEw
VBQxfzewqWfsYc1O0u+TyL0hqEBxWMj1V1yKiZ5wUFydqQi3WI9a6uPV/2erdap9
Eaj7Lf3WISxOxOghd/520BY8f56fuaKO5gFP97xiDn3bQZju6HpKcFjXi7ERjXNH
vclAHt3jeGyi6gXyTpWdz8sza5NYW0c4CKrcvxnGxt5PJsLUmZrGe6OhWpaJsPXH
TbQ8RzZwQlXuNWFKugK0b7kvFTbi4uBPFMgUhPSg3eUyMLfZEaOgM8nG5mOTS6Tb
y3DyD+0o8BeLLFT7PjupFX2kVpZzSJQscokT7DKqJqVHf8fjtvX7tEExtZWXOoWz
4m1gexkU02XKzPEkB8vQGkNHOg3Xry+fPu1Isge5TtNC3ZAjo68aqWPDHEl/Xosy
N1Jq5ci7tqrt6A8vAm4UBpUf2iDKyXN4D//dumAA2TpGTVhroQZ9cjOXwxiC7XRh
mbjwZU3qWxIp0PqCf+FPHkowJltlULmeThI1qJJEyLhyUjvopsUJ8gwelONsBo3/
/GBfR9YgSQhfXYxCgPl7WnMmchMW1QEb/UZ96QKh74p+IikE4qpa/l8A87yJqIWU
rwCM3JDiv5q30IXse3ilyUE+/3EA/2dAsTrUfBZWvQ3Ttedr00sMsW3+RhIBOXGi
stMUthvaicqGQveL3NsgBcm2+y+m9fF47UTqclMNQJLZGs6OZyQJoqb2jmqtA3uX
NVPMcHX2TKlCD6Qj9MeUkWs1CkIhL4+s4xagGRdasElKKB+OqQF4UrOqxEdiueqH
0n4+vZnKUGOZSIOE1C3kIKAwxfCYipyZnfQj3/t2sihobjedFHUDKmI+q4HQPk6m
KIG+pqtOT99MAjwv5lCz54GXXnQkKsMX/NFjDkTxJs3rozo76yE7/2pd4p3v/COw
OtsNHDIvsZ4G3nYx04HE+6BT1cp6JcI43ipjC2Wv7+M+JzfwCtu+fqOG+1CcXtfm
bnsLd5ba5LT8z2K0wjIXN6uJWx6CSP4xPQSF0e1gKkhPtC7PnaaCCMDKB7N0OlEH
XtczpYfVtAJSPsTAt2nZ7DjqwjyQzZS0GbCC8IkfJtMM6rDJSxa0mWo7H7eZU794
UhpXJ5gtdY1c2Cq3fbdksGGX3Tow3Y+ykp99lZh1eXWpZFDXXZ1gGzqDNCGFz5K7
FsU/0QfV6fkh+QgA+N913vMnHyE6aMzSlJZ5klYkqJgaQaFNKHFR/I1BLIkmuR2H
9Yxl2/sJz1jAcNpuN/34aw6sPICJh/XHGBkkfBrUlxtAdUuA0E3u71qEiEOVl57c
yebn37FsN6WiZqGqkrvCqJ0r/5fGXhYJ08kvKiWf4GRx0M0EooB+QjGVz+YydGmS
IR8V7+K3J1R7Tyktbsvs1W1IJqmhMnMdS72SiL9cNlISgwS0f7n+hbCADS58A08n
nx/74F8CUNgzJX78crDAG+llqhVu3swzNCBdv8Lo1HDBhBLJ20A40+P6aaeDVacL
xOrmWSTeEfpsXLWGyI5Xug6mkLhhWZW1jNbT3pSFtaXWnDU0cQQ11x9nfbmUW1tg
QVIyhj960uHszVcMEd3qCuqtrbdgdSPV5EQfmFlFkJMTHyHt0TP/n9UGyfqNlJdX
/2Rg+PmOrlmVUpS9JrYpcZq+44hOavVPAuP1AVhyfv1aoW8S8jsZp/R0KSLZ3LtN
pmM+7ybgp9skO14d3EvrXBmI4fyGZbV6+F/AmReQ4NOxoOVIf3CReReSChvz6NkH
qyvEtak6Ck0BYNguHu1+kkMJTZocG0pOFivatYK8i0N9zmXbIKcLvCdSQfGe8Y5O
TlaI3sCGkL4lMwJkdF10FzKCQQm27LBiougy3U9ZG+gxSk81ssR99sFk9xswNiIh
LkuNO+gA3PI44ixMuSwQ/MNyxTAVDCZAEqzK1aRpMG5TOw/FJaRvfaas8/Of17cz
b5s4JlmUO74evtrOWGo8qrP9jhp4ZlBi6YP8bdXzbW8FbR+aP7GYZGmcoIEijSyk
Dy/ZTCYK/dZT2sGfDyDSScr1E/NQRX8gaWLxatcfjGNJGWeZUJ8RFJedaMFQMjGG
jjOZNApAS4QL5i4dwqdSCaglOpVgA5S2o3agRp1w10tPBpuHYsnNPN5om3lkBNh+
axrtts+fKLmjKKcR7IRpPtykEiAoXZDIKPvh0uDmoWHsMxf6EuZtcNIUpr5M0IkG
Bg6oGl7vWirPpM7TnATg7znckXArx83FsYnHIpZZvS6w/Eb163U119rA6qSld6WE
PQWEDy0XBC2E5Nr5AIp9bhLNW7QQXqPmbwBKfg0+ozaddL1YUY93UhthEB8iLJ5y
Knj63djQ+gQyPilJuHCi7IwF938XOITKdjvx17zI8giHZXgh12/5rNVWdqnAQ9FI
LR+UuXazN1P5D45lTq1xPB7oX+lOjWGai7jgiP1f80P3buv6PZoc7AWWM6KtFeiy
kEDQdJUt/wnLmQy0ueaGFEHQb21iC7/m8+Io9MNQlF+fzYkEAe+25UNDPLGDw4y6
8kQKRLmEfWq29v7ZYkrfHye9dGTCJrpnEX6cq2Lunhk6tWHIeD4UH50aRjntFslD
Xp2pQ9wuW0hCQemism+EGuIS7wjiaoxSw/evFvcNhrIqI2NM3Z05wYJXr9GTKqHV
P1nIz82JOoYLDBfWuIJuZOPqUINjme2WpMPYsA/LXy5aIa3eaTr4OiDcPD6lPrMc
4XXhRM7A/4jqq9Uqg0KeLxD5Dk6j6bzFeEzJGd6q+lG9j9UIkHbZUChxEsHQE6K3
tvaRbWGq4oWGxeEx6J2euhk9fQC1KtrozPLce26hJz+Leptd1OGwI9hSqC7Pm44B
ZU3q60ukQj7NLSKHTHz6a0gNCO4CuF8oVERjHBMaYOMjZ6ow375nO3J+Ulv7AuuX
UqxIPYeYFLKT9wj1q/EX8YsM1Uils8rG0VMDU8nYdXPF3ZvD9wKW1yjRJBhfciZr
RsCAiYRGCRyblUaT7tL9G4uJIPL+Zfk1RfkbeJwiO8ZrOXwh3Y/B6ZPFYFQ9B4bk
YcQUyxfQCV3KarT/L03YM6RTVe6thYwCh5K5xAoA73gxfpPge0CmfEpHQX/wouva
d2yr5Kj9F5uVKQZ2MprKJPGCXUcdTI4am19VusMr4wZUA5F84gky+hDxhT2/IYtB
PXj2UldF9wY4zygX4m5it69ZsR+Tw4dqnPnYlcHBOSqmNuLUktKOjZKiknLuAgrp
g8tY3Cy7W91qIpcHko/BI1lGN8tft4Q15jAZ4w4AkQnhUS77dSw6tiUgCbydxKxJ
oLO516Vye1ma7YtzFr1cGB9jbrcjhC0ZtJYfoO1XryZLPbwaI103MPNSTDYwmnG9
ro5XdkF0BZJyKHXTctRQmpYvNzUl4ySmXIxHVkSi/1i5vXEm8wkgvGzcarYBl3Gb
iAWJ1htPYXrd9iRvB87V+roXqvceRXjDt7BLTl9bnNLQLqNdeM61XgEUFtwm61ZQ
ohaVgFmeY4Mzi8cb+IascbIRYsfq2Vv6uOtXI6PGx8UNvY9BNvP6c9Hkfr3NWn+Y
tAOy/v+GCAq01k4BeouyznPdUFJQBHexgBpHG7l7TpBeGA5kGP0v1yXPmcRYboQK
LMlU2K+erqRrZDyOtgXFF0QuWAGX2Hu67y5sz2HyVvZsiXzgCjZyojyj7Gc1fiuu
LeNUcZ0Csi45JFvIEoaKjSzgflWK7iwOkI0qAwO/GiHOwUNfejB94cC8RwqX5LQw
f1o4xtGsBQ78lE3g0RiJoaw7XUSknMv5EVUB7BVoIzzYvIRMwCJ6qAoejw3nUMsQ
qBBAgp9c+FDnDz0Dt9xV2tpXcHCLlalFB5onb64yhc7dAeZXKNyEH85pKIBdFu5N
IVQpplq4P92Tr47FlXqITHf0C3PbQGKVovkrN5R3rlDBV2j9irmOYH2xuoA7OvwV
ikz0OH9ypUQldZp/Gr05muUN83n+YQMf8yKMglqUvpagAmWkqPyzDCqEkk70e99Z
tCbmPAmkNcWFCGzDpPBlEUIjLw3XoWLSIIzxKfwz0g1yK3fm/anpsVSVumqimNT6
DmrAIQpDXvMEKRp6UjdIIO0udngy5zIRvM9aZTnMsZVE+6g/Uxl7j9WY2Z479bdY
rx6DzRI5CYmZb9gG1X6i1PnV/JBroQ9TNrV594UJQZIK2RhHaj5yC138itMj6Myy
Ai5I+irEkB1Rg1iN8t+G5g1BKjypigIYVsK4yWC0gNt3vN4Zv4yLIieXtlYSzPzu
rhakXYi6dhGstnqL821EMlOuQ8K2d5OFD+F5AxPRX9mMeug4uqdX550I9YWQQ/Yo
oPm//tv6Pw2/VWjEXasfdt9K3jgp46tY3h2v0Y7Vomh9NpSL+wzzSIumQSM28byg
DSd/frt16hq3tJ7RwHneGg6SaRaqR2eO/G4mAAN5IalvsIcnmL0iYzMSRrn7xYN7
wcdECgbx3Tyg3ZmLpYHOfdlQ39qyFxPmdnD6pITqQbVyHMCUP7UHyu9AVUJOhpV/
pT2G8N0FIx3wkTodHNvUM1LRe8xEsOS+o/QuLVdus2nh/wflb6FRgCEb0eemGTI+
FotFxQWfIL26MpeML4aej9q/aEB3Qnx7mFsCT0QgIaUO9ZiTjriJGdeOfHU1Q/JM
LVVNtekRgQPnNHXbXONyJ5+5F7A8UKg2Hf3Z2ROPrITsMFoVZLhRDSbZDb2Vi2eC
11BzRhJJjga5qLUjj1JDPCwq+vUcHl+gQqSasXSJgQzgPEW+CKjDJzaLPH0EE0kX
rLKPUNIl5uWj2Z+DjH+ng0ZRRKGAWgbnbXQg0GVTnm0i9j9D0Ai2hQRP+ixNl+UZ
MRf1XHSDlOAOq7ByOjtDbtnk6yMMZutkBS/rIxYE8tVzDTQlrVz3hamzcMipevRq
ZjXpGUl1SlyIqNCHWU/IxuOyBQEe5TR2WrRrh+HV7Gnct4sp/+6krxSuu8r4PtGT
82ek/zFsiAeN6FcY8uEyxurzq+slrmnv4Vlvji0L3CbVMYLnlDY6GgscTQglfpys
4fFCW/ePDCCZrRi36zUtpV+HC8w6mJLqfpkzUxwWx4Z9gebPUDsOHWBXTTHfhOL7
qm9GthHF3TqKNymMX7XaIvzjkM3fBBGzjHS4Nx+d3+EgmarOaD234QTPKZ2lOYdn
IsJs0whjIugq5hAmfwA/6vnfY3hm8TUOMmjD/fO+IV1fJVxqkP1y+8WtApNIYXqg
B3bL0dfyM3awaJp418onaHc2mW51gXCcoHtq5HbPByfxXTMXfB6st+CN97BTRAs6
6hcAE4QbXqh/fQ+EYOIyLjPQqCtYfL0j+0mdukRXMR5L1H39DYW7LueX6LRQldW8
hOt6rvOaMRzz5Rud2MYOBudQF0MnFpin/O9dNcPaCgDNZahX3+f3yt0n1E+OXAdd
esDbRZz1VLSDDJn6iM/JWNJV7nZOLj4ExJRF199XK9CqLlOgoZvECBKlZmMpRbf5
ZFMmxCw/aUuA7D5UZRd+IG/JOtD4KMe1oBMrlh7balvgjN9R15ZBqcouxkwMz9GB
r+sVtBCBBYUIAA0CrBkscsE1eQo1vaJaJDeKDEcCQsqYPZQuLdeWfsg8o0riCnDD
v/i1Dg/JjYVgjjlN+aZWUvCrusblhp2VzwfpPBIcuCqe2NeqhgfyNLTk915bYlTP
HHndI2cSGr8IJ0+RvH10qRP+VZpUN2CI4Btl4UCNFXUFg/iLxeNwA2aJE7cyba/7
g+E2YOak/5bN9/sqP0HXaoDVUvpu4IcjTJfZ5YqcQMSo3unNksr3hXwzgVklq6We
cLqynGssXulgo3UMhMsrj+5Jk7MCOkhVhk+A3StgK3NagOWFJ9a4qw6BctvFzSIj
mAanvcX6r77+pc/ZbBm7/KSBybUrFZCb7wawMBOgqhigUFW+bQoAnyU7fE5gLC5M
GZzvZnMlg3S5+DL/q3GtwZ2ETaIyLOoWx8qx3obV/xkpTTZOrRTUgC2ufxOUTxcf
IRAJvdBrF+3zFkONCkN+hInvog8KbMY4oYXXSCKgM9lLGZB8h0RwiIUsQWyGGQkc
fmkzkC1+NW37vVIhCxgeyQOC0zhi3GKhhrG+Oqa6MwO46yis3VfPZQkjP9wxjggs
BGiPSptbgD3QnXEQ4W5JqsPcDar5hW92jKkAwHmG9fHLKk6oW+tIDsyvLd2nqqw/
bD3uBuYZAjFg2cJKyejEtUwa4J0EaPooyNzZeIR5njP2TxeWEX4fK0Od7qIUHBEq
i7QB1FbwWL1Ncc9AGaKgKt2AFhWhFfKcsl/72ZZHYIFl01AXqo59DEZ+bPUpAUh2
9Zr2jMlHrG8tvsXqioCihHG0B6rWSCbvfG2PU12mmAywo4uIh2YdLpOGxAX8ypev
ptxNjy6Pi0AHbc8/dF4E5/oJFUJy9pkXNatgpDRrepmai0p2Pa0flNDgQNctxnDp
lBSdZRCmaThYeTNWWFysMl5bwU857smMIK0Is1rebzKIYrciAHyUwTrDHefNCJNM
xXnfJ0Z7mhPU/11vADfT+f97vy0u9mH76G6VwvJtOGQIoh5RtQBOCALkq0TYSBdx
UuwUYG0UTemyTS/6V16X3L4vdxdP9d3RverLSac66np6r4ppMXa/x5WZ+5PND25P
4HdVqTH0QTe3cIZa3UL/hyfEVmefxLEqorBC+zTyb7ds04dI+Gz2MG7rrjgYEP+s
W82r5LXlBB0MOUTUJmqnv7tB4l6Qxf7ST04Ju9CWx0gQw2ZQl8CpeNI/Xbm0a69/
pL38H8xpi0lFyzF5dimDHB+Dq0Ro/1vW7rSDQeFt7eAs2o7xUsQART811sH4Na21
d70yXF/KqfzgE7uAtCdHryfhRP2FnVH+b3j7vo7VZrxiDCME40rskJdETaK/o55b
1cg3/QyNVkdP37SCpTspiCU52xQXoL7RRF14BlNjgl0KCt3XD7NDastmBytzwyB/
FkJT+6uXun+G86wa++Fr/xgSfTH3MDwQKyRaFy35gUIaMZHYF40LmkgcveVuUCLo
vBCjxujrMsY/nMIs8MZU7Bt7tMgisI5qAmksqlW+EfVDaTWV9D01KOPA99c6aVSR
ztbDZ8PYaUqA2j3LHHnywLukHFuQz0XOKKMxQHrakkokfJgnGe8BW574P+7pAYbd
lcyti1HLUvqvCfeUvFJkurQIitb8mnoiwtYdjr7sphI99M9AzU85hgy8poGyxJju
lgTNSUBNZrzuWx0zE++J7i/+3roOP1g0Qlt+zRlhMUqkQCANpGQRCGGk28va4Gor
G4xPRFhrXyMqpAcGLNHb7BMGmB2bhM9Ov+wuGs9BuJXX++Z0VjIVORIbdkUvUPyR
CPX/F8vL6INdOFs/TpSm++q0k9FT3mpA3sLZLYTHN10GvitqsJ3WWwFJqmFVt0Ne
YE1hOyLdyUyTXYQPYQMIq448/z9GYPNoRreWWgij5EID5B9QK0+hlT9Z7mcKg3A3
t3pydCGlBnDG5ppH+Lo4Y3x9FGFD71JrpdgSD1Z4VF6vcCzSErSO+vYqRJfZ6XKI
W+dwuk+Z9NTH3D+u0b8t2IbfcZ2eW7kt20bs8rF4QYAjyQGxNLEhnHwOjPKcubtv
K+NR+5RvDuFUk7uawzu2IKWyVik3pBcjEPyDTDqSG+y7zvgtg8PfccchJBXA1bgr
2ZCeY+jCbjQ8EiqUmtO6UR5lGMm+/VJTJw8NfTIv/SI5wsZQoduc1WY6rFoo3h3/
Q+Sp2wf6K9nv3pQ+JIYF/NErMpkDF6nIiJzpgX5uQ2Niy/aR6RiCJDSK/WpLqixh
8BR6Idl0Rb2tSQflboY2LF8gjsZa6f1f5kz/TEclXPoE5hPq/aKHr3TtYRB9atfD
zFgm8J1ydooQ3cy4cP20fxM+YQSOWfIEmavt7YuqiF7RPs165aQ081ybIK5eyiV0
5JwO7es4OFTNeBafkEjSL1ma50w+OrAm0GBBhBU2BVZ4BPpqSqGPhiXwL10m1SGB
2E6FmlaUoOIIgNFZ0a+/0GvsZtVKmCL3Vudg4K9BuXyMA0nWz5O0+CEve5lRrcPr
jJ/5ZaubajuXIkfu5FAAauLuQq0wlnQWX/12k+UiW0p0Pdyq/6zELSC2vgJyo4T3
aiCO7sYaH80R45U6pbiZ041lU7Q4Y4pFiUzZbl4BY7VNGXkKb5AIReOYdo9bCZpV
ymgTHp9+5vLaMNlNC4cykDZhYhx0YSQ2fbXGPpsHcey+6ubaJ4AYmLOWRz5PhIAa
X3ORH1t2yf5ghnlL5EyoDOfoRsqPVXJLwFFlXpOk/Y+kjeK7sC/7T2LQz/LIm5Y/
gjLCxAlZtUEmi9ElByiVb19pTpRd4NGc/LnHRWPiBicQMqwUr430DM+/3tuZLvHZ
bcOiwNRGVvniSlrn3MwKK2gqBAtpGG291tWmh23rGbwaJN9U81P2pjy2/hiNcq/m
ucyb4fEE4mV2NnaI4r0AYtStkPTjPYNpOScC6gIYFvJHcjOQnG2yttnS+fGVEo6n
iQzabNIGUY1JkKUQwFD4HUsQz9B+7J8LAwRgtUMcYX8xZIn0hmriNF1fu35os5ZT
+0ze3Spi6J1KbiPPh/b/gVdQ2VccAWtXC4w7bE7/XPnjhjPQDgxO8WVgwpOX3TyY
U3acIG9KsOpon4+Me/Hbkdom7lYRasg+JJ6GbW6jCWoSpt7aD6NYrQElpyIuIqke
KPs7rjv93dRjKhXdpo+kSoFXJJPGXf4zsXSL0kjng023v5tXdZdtsAoqbReXsTXs
ksr/cJl2JgT12npXiSELQcjk7FzdCMbseINzKdA2+twHNb6DlGO8fbIGgb9r1965
gEU1N7wPiji2tzQp6hMEFzGrulv8j95BFox4m+ZqrXqIxGhmYnRNkKl5iOtqLFuD
blZuyY1hTVWoULJc91aHTE/dSc7s4xNc7e2nXv1gcpdVo9lwklXNaBHwiHfyeaL8
345VVoXqsWjdB+DecUEbZl2rdZ5WrLs3nYD8ncDJHXaWV1SyqQSvxDSNk3CRzC87
poUlo5/bsfB45q/Y+g/iaqC7LnGg0NSbYWdtous/xDj54IaeF4+FIuKp5tx15Apg
0+BTJA7/4/k59/0UPKuZPrncIeiUSFWWO7Ma4V8jOzFeApmr4+WLxyhBJkPE6FnN
5UUHNZFFBIUzzE32MdwdY2Aw08ch3DRpimSFHvLPASfzd9qf3U44W1cjsB9c67od
6mWTWnpLrgjw46oXUk6n/4U1vtWx2b7Kk/wzUK40Weh/LJ3pWqKcDoV3KnU+14+q
DAxgOfRkZnj7EacuXhefhDldE6liMm4+ShogBjMO1uavvn5p03uTTouCf0LmDCkJ
zasQGKEqS+2dHuew5nwfrUhPOl39tspU4SskqnSmU9/gvl7ENMky7SPiwW4Non8z
JO26SQHU5OLvkSmP4OtqYxeRxe1hulalUy1osYYUkq64on8f84Fg+aYVgNeRSMi5
0XQTgX4KxA6ig92a4poKEMRBdquGNKnESca6IhWQwSZYitwvl9a+IZBygg58++Ts
04cfyFFdVcWffxA2vUkpRD08bIlONAnlfLYi41bV3DH4wtX5CcN5cVLwGiHkKslx
PCIKzeMCH/lZ8+o210M3uuXJs0VD8EidqmIUSROSQFj7nS2KWElAHo1ZRWNB572I
Oy+OUWgGf5ny3f+eGr6HR5mctQvmG6RxgPAU/mxPmnTIih4QN8uwsh6PCHWtLZMY
kM9LbHZvg/IUsRLpH4HF+yT+70GGjctug8bLzLNq2mu+CBCP7O3b5zfR1de0yz9p
+NnHDo4U9WCE/WvXaJT9qJT6l74TuejtH4UX971cwj/uz1tj+Vxn1/WLpBHIyQIA
pJYdy7twKumQSJPfYKVpfphjoXjWTWg6vIOxO5w0qslXKaVzlO00YGSf51/41qp0
qA7bK+TW1kjLkoe3tUuylxzTU1r1PaRYcvFN0VRR31CRQGtahNq+N6RgusNYL///
ptPvOeT01zZ2rDRuwHPbYdJ9qkjpt4I7Ls0/nvX/vuy1Sa/mb2sTZAKfCh1LmPgk
uUBD5Jh+ucaHZUuguZGmvSVpvX2k8nzQMKw/Byyfth9gdGOeIQXruyhHUYfbbqb2
Q2yg83EgStDr1O/d2sGr50TMD8K9B5q8dWt/3RDgt31Ks0mX7gKe/Hl1uOahECe0
LgUAi1ED99ydLHx/+LCQG+yVuCWnhJ6PYzLv5XBKXgf0PXBhH1+4kDwuEsU1wh2z
RKE08XjLg6yz3q1D9aMT2S2kchAalsvAbSI8DwTQZX1IJKeJ62ypVxQbpYAzFxfk
8z6hkDNc99ybi/6WE0a3yFisEYaIYcxz5F/lMECECbewmdXFs4XkNmBc1guD/Gmq
cIu4F0tmhhxtC5KZ2BueK3uCquslCmcaWBTFf59wUPo77BQxrEeJ3S8h5xg9sMAp
NQqnaWUyAe9Cq0hVXoxbEAl+Y/6QsIUpM7rSsIV1r/xApO96epdS7lH+J91oy0FF
NxjxtIs4cuF5+3wACLu0joEKhdmhfRvhZdpueyrLEo3/pNY1FDqwRmOU15vNNvDB
N7q0d4GTkQdKxP+Ozam2aYXgQXpRmisBB35Vx4c74AVhPKV9UU5QGFUdK1afXTci
Z9H25lsyCLEs2KnWEsKglsoDrc3ddoS86ilHspsM5FOdM9Ckbvic/oZL/rt2HAmX
//Vfk7N/3dAKQYJ7tD1ZUgON/LoW6yJxU3FSHGtQV1W13+BLMbyqS17cJXosZrlp
wsCmSBzDgBx7z9bBGGq6W8hx9n+pQlD4efVi6YesD2thvZexi2Gi77NOg3meK3xv
Xk0o73TbukYLtIMoa/zgNDfWTrciIEXINjhh1DXGiiidUWj5LyZb22w14m3ndcq7
79M+GD9Wz8mvxSpU79Kth+Tod6qk41IvghpnVAVBXwUZhV0YpstBuiCRhG6ZeZu3
2nBEUq45y6eKwFW1AgUHnVnqc/dFZt3L1y/yuHXP04C4i42QBV4wstVneZGgx/HI
f0ycEUrlLQ0U5ZaBuI+eCSkZ0HqWSTbb7ZFzvtmwyayRwqlIvJJDe5gZlKCrwZjK
fcvByo+k4hGewg4y3RfZrLnD6IuL1abWgpiqpdzL/4+GtgwTBLZJAGfHzZU2R7rr
RDoUQ5ulkJEHQhzwHaFAFIoMNwYqlg8mi5fhCdvQNZa5dzgDXGDzwmyWaIArWWvn
yBcPo8rJUCBCsezbj49d8RqCpjePEMduyJawlhYldJ7bBFIlqdfWLR1JHcUdPyO1
vlEy8e/51K9BeHxFkbzYxH08K1epIb04rVdsGBXjC2IN2yMNjGmzTR4cO9Md7cvN
cfPI89WuE+G3U2ynQI4vLtzhPC+ZqfcC4ZvfztHxWZtIXuKmd2hihozzjHZ2EJeD
brMg82YBdmaVEe9+Td8c50lTLnSxD9kW5ZOtnRSeR0HYhCkTUHLRKM9Lo8PsKcHl
JIBDzTG2aSosJlCK/pKxc37n4atthIil/R2rtR8MzMZF8n3K0h4EJRJ+oHxNWkfT
GO0/mQAlwwwEvorlzT7Y0A4YNHznyRwPrQra7jf+pXtxqrk03Q+nNZ0R1tRdlzBV
wVq2QNMVwssnLXfXXeZQgF/LaLshoboDZDb3ys+R1MpzRjQIJA/MilQJr7IvqjOa
vhnz1H1kCnfUtkKg1ZuijNnxrJs2hrZ3XU9gRANV+df4dpF5gbLZs0Xxy2ZzFpIg
wPKlVjjAwFplMsMn5OXLI4/+YZW3OlTJU8rM+DRWhiWjQSC4SvZZQC2EMtKl2epH
rLpH1Cq5K8uw3+U4H9oK2Wa47erBIraDW7e6kO44RKu7IjppGsCgxtHigzoClXzJ
Ul4R6r4cAg3w9u7FTzxsv2DYdt/ZmUC21ArequyEgxBfStebObiSHHUZ4UyCXdYL
05pTYoQXtv6yLepbhs4lGVd34mw7FsXkSy75kprelx++NM4GxnQqKgwrb+cn65yK
vNaDD+jHRY+myYVzWmBHngo1dL47zQs/NyqZoFECIlMiyqa8U16ouIfRBZJRiP9h
kw3EdZdcLLZ900P6px53w7Z+kuOxjqE4BPMqJR8cwnSU2NvI807gCQAFT/4hqXYa
tY+XxxgY2k9gBF9nK+TkoraGG7VRJtN96GJ0lIw7oBKKXnhbLgF2BitQFs7+mMeI
I8DbnemPad5WUVXmgFpmqieXh+se9QxB0R7VdlROOJT2e/6L29ew733Q3Enc2Yr0
0XxvY1XRJMfcV67JNeGobxKv09dGHBkfvqg5CzLWdZqSb/Cib85dVmVlWgv4AQSb
uYwS5SwVeoej493qExJBnwFrZlyY+IyGcnpFSG+ZWTOVrKjGbkbIMLMe03cQQaS7
N1zPWmLGC0kACUhQM+tRYD9zix+f9Ycihj0oG1C71x2LMEbNyXMIiuocXGGlM0fV
L54EmFkcJlPgm5mQs9s8nhrCEGvvc6RE2nUqKXq1b0eri9cXpNfTc3PuDKH9VyHa
WTU5tx7hb3/26cnw2VHi5uNHxHF1eYl5wGdAs+ofvURxj0PN1JVotCS45+PIMur6
OXLBKWhGHZIw1Tqjawc8lQPpsyKPuyC6On37S+lb6Jz64t1lT3QExVQUgcPZRNT5
S+6V6fCHqABLdqs8de3jqg0wibn0EVtCy6WtsXFY1EmN/w3FFuSww9sZpQY5CC9d
gooPzADIM3WFv5LaCd8TaG2h1AV4Cqsy9kESCvh0LlWgbO+BK5PSWIWDs6FGd8y9
3TYLRndPL4TH//tQVXSCH0/3JDHkyOkemUN5sA5L+TmHspC6FY2NhOKYxB8eXqQr
Dfryaqhi8U1042iD7vFvEI3ns8kZcYD+6KewTkWnySwmlrc4AujlLchA/Sj0zv+j
kAZXszc+MGNyT+7WUizNdJ+gphFHwH7K3mEuLJWkrUbDStMTk3CJ1ZfiZsZ4NeoP
Ly7PiI2YgXuvHy8gQCOGAeesypqRIVcDt1DyWPVTPpvNvtjc36GZQyAG6b5VIpDS
oFOiNQ0zNvwP1EnCKQV63XLj0qVRRTLb0/CfCU1K2sVmESpIlSVpJ3uQJ81SSGUP
Uqtcenq/ccrAa2TlP3iruTNSpe+hCsiTU1ixfZRkQocYFsHKQXQ8IMgT1seFrPbx
uM4aVqs5DQhpZHU0cgkBhGMTM/LE954jkhg9h6bZ91Bf1ty4Bl86U9ZSyKF1CBLA
gHj6TVf+EWeEXj4NYmzFkgH2m/2j8cXZCUycXhr2D/g792h9HeciPYERGD3D4Cn2
vk6sv/91UxCSZo5wjjAlfBMzLI6kx1w7zY295D8Lj9OEqNrhqklz/jugLC4dIxez
dLHzSh+t5/KLpMPGR4lK9CrRRZ0qwrilI1chSuXguQP0YuiHhJWUojV057aeTzlc
JrUDzUeQzMMUHKufqLy3eLksKlw+Oyz0/aue0c1YQTOLs9ifqvSKpFEFu2ymWdYK
sZX+fe6rVbwPhbatTFSmDGaMDAIikCgNn+g8S7cfazz7SymO9ntym/WWPnNYN77O
n1+VpUQN2fyo4RrCkEPyayHvXa9wu8j31p2qYzMEBm42vfwzchWZz9GBY8WIhcrq
DibLzMLA2m3mUt5oa7ScqolANOD97ZhHcBFuPHztYBgYsRcsDrtMvLLUh3HLlhdQ
nzKH2mhrBmNeWYn13XyB5nED9QH/tdF0/CZfF2NAMicsP+S2pFg62U9kn1cK6cq+
SkKeR2So5YXcq81dvt+DIYf+zgbhgr8A4I0ODcO1OlaV9yuFAK3Ox2ysyfEb2IJN
xV+cYI3W4K2F8S45QqYxIpZqp2t+++BxaJYElUpwLlyshK4BAKJPJcXr4lpyKRel
jvrxffbctupi10+8tV6LF0x3dKk0/w7fUXVvA/YHT9GIi2YwbBJJa9u8VQeNjhm9
r0GR3CjuIuobfjw5tuR8u3uX7Hl1f40SDx4EnKCv/Mr5fL9zDpyBcNHKGIVYzjom
6JGtIDdZbsrc7GFrw5u/YIlLpS4nZ7I1C4q6RN40pLvFTqjBOJWPKb41gem1IJ0e
Xt705awW643LZnvzaCHd7vlIVljpnUjwK2wcL9j+tgfTntBkRs1oQX/ld6yO3bVQ
NevnhYjjM+fka18NBc5ynLNJcmpZPysI1+6VDF06cRANZgTk33M42whbCiiCD1Sm
51BWokSNqsYBBaAaLciMk634iTdoH/UiYkvfOxHF5OI3oxxb7CwtP3g35idrGGW+
Vso0j7mkyLU/B/1Vj/4/X9v0jJImBcB0xu9J+SQD9GuoeGaLXkyTWZnBvvi9UxTE
ob5xUgG9G0RUSKZ5vIe8yjpmT7tNmqtCq67ZGesiI2K8ZZegfzPF7MlMoCQyGKST
XVvLGqElzU8dxGDWIH1KaArhf/QdXUnVSXAKrbynAcrfT4e+/SRJRnPwDZPQsP6H
su6I504dQc1SeASS8Gon45lMgLAeKw/dBR9bWQb+cuiGMUhew1H0l7iutvyiBIIm
YWM+JABy6DZXM+acZAkvgs0A3KXE/s9YM6Hv3epfO8ctMrQKFtphHxDLow3bRcbC
AKYkB6iXa4SDzcix4GEBoQDfA1GZYz6ilK9i62GFeXKBQso/GS2fuuDw97eGlhVj
zSS/Jko6xEgT6ROBY3Qcmc54bAC/76LGTZiakMrv3x5rz2SMtNU8lk8izQpu5tiC
QClss7TcGMY2b5Rn3bCg3isrS9DF7DDZquTzF70OkelukXkpvZtzQ1YBodkgbw6V
NTKz+n7kGAmSshhqIosnXT9pDLqih2fbjw4dnOxgNWik4BAuivsb0aVmiKdSdDbl
TyGuf1hyPCh1sgXee7p9Bu1kv91rq43jM264V7uR3KVRLYBt1Jkv5pB4OKh5OTmi
4R3UxFX6St6coI9UPQjd+ZIJfkBftogJzIqkZH991P7g067W7y+JpVQpWWK2TNBW
moOS9IjiaSzPF7o4h7sUmTM9Hr597pE9c4tc9mLsmTGKiCQ46Lt2wLVdsBvDhnEr
sa7IHnOtG93LnS1eddAeCWAYrzlQgs4vPfz1IndlZ1Lz4NT2g1dMyt+cCfFR1P3d
XC7Zf+nTtl3dRuW4Fi6QWHmqiwAEDIsj1cny+uszrqpPReHZQe8wd8UUn3RrfrfH
yKID7lksIpHReUkK12LR3OI/pXRLh6C5smCC4ZEsihvDi4t6B6va+gAa28Tc5Kol
dcVp9cA15ImuVMVXqAj59PdhjBZiPeJVzG0V6oPMnIeQi7bF25kflqv6yRvtDIWp
Y8a45HK4VWYFVko4jKZrE4NNkZkHnAEjIn3AqLPgRs+QgtWUz3LRrFDJyE7hS44E
xkE8W3enKwfjD+qzOGPUwMLK3BFbGoAm2U1kD0xLvQ/WUgvmHw+r1bgqWjIL69Vq
A5ezB8vGw4ON0hQYWq720hA/2q0YooqHWVYWK414gdnBdhu82aJS3OIDIHKysEzT
ujXJJFwGc8wD2NMxYnLEjmn2+fs8FWoMqq2ur+ycV30zJ6/50S6brHeavXpyaILo
qfKd0Co4AqsZrecCUr/Kzl6Cl/pbkavIJh8QjmLYPX7NXsHZVjsVgWLZWDhZtyDM
tyI2/PLv7b9k2HKnNB+REQ5Jaw9M074PiBi9kSxSRVOlcOzd4iti0tSfgTTtrKFk
DFnFeGR0AwJvYIQf7BYVJx+mSliWsYikt7F+TxigJvRuuHY3hLB5RwES/pKW0y1z
f4b8NE2fuj1XypKmdWvQeKVu675KeMzTvhYnSbbigq/dAR8yMkTYGacimKSePaYr
L9dy9JRlFVVBC3gHQDQGPJsCOuQu0hkDaJw1g0dqyRWSKw1qA+56xdjGSHwLSzBd
gPf1G3cuRsYL6kTacQqW0llmk6fd7PBdANMkxk/KECg/DxVjMBFVXtX1NmMw9EQx
rRaJY0LQjT/m1tjy/YGvwu2Uf0JmdqbRu+MJ9TniGknpasDajMXk+JhlOFzJ64Bt
KFQVSlp8CEny8+EywfPfQOZt+gJKHZcxF5h/KOzTysb2bNOEuUBO2RKX9OQ0RXkX
2t/WrpEx8rRYi7kgb+FaC8ELEOkWbxMdF3oHeRS830mBFmpCVernhF9AbTvdetRr
ELvjHACKE9RchaJXqL7RKvrHUOYMq0MX7b9zzwo6mFkXQLnujrysCNkInLKE2mr1
eKss73cyHjartHrN5T7LyFzX+SwITei1glFAwoksZ+5O1Ayi4zK6RQ/Kcw5/gP9K
jh5x04+4YBn0MMF/T1J2o/ZHnvWmBlPppl5pZppmKCsaYXNskXboW7rc74vcL+BB
CuKtU1tNooF1c6viotVF2UWF4eJcxSJ/JHgCHiFENgXKwe3jWMJVDj2jK5+mcEDR
WAjlKDXJ88fveskgfhqvz/A7oSsSP4+1u5YNS3WSt/aXU/9OqZn6+FAo/Kl30YYr
oQk1ReDwJQfyzoyztSfS84cptHSRv+81ukP1RS/RbGpM7BoI93A/OcB0XR+GukO4
R843t5nPxRvjycZgQOZcofZD4cwYoBcG2GUfIl5Sd5mXrVXIahlhgUUcTne61DTx
xo1pgQ5PHX24nP1c0LA9CB90qi0GqXeFaKBcdoKBm7LNgOcTLWXfnzF44XIkHjVb
Ke/mxtacxS5mizRPsTiM5oAXPp8XZWJq2tqmKjQWGKtUfZUjVuEJYF6YEY+AFXnC
y9zM2ElRg6DKSB/5iwGBREykMqWmqUXqSBVIW6zkKJDcyBqe99O6+SYUZFNjsm8M
zgITKzg5CJOVATnMZwe5dJUMDyzNaoqFw9LaFDGnaBbrVzGcEfnYOfoO3ZTiaHer
b2xrWJd3Hsg8hpBPDUHXiWnc7QTx38jJTjDKCQzN+epuUnunLD0gTUhW6vvrjZ12
T4/hgNvaRLkarhxqOiePAJ/9tbiHMZCW/iqfRI8fPw1SUHPGY8JEhB0SLuOEILTh
FYe1oAtW6fAG3KL6Ji+wxdSfKWLumLYLxw+tHaPLhyd0xN6bIJt5X8Hb9acu+ZPD
LI7DKvrmcslLeDysSsLyPYRsC/qbjbkZi6jWHsTB/DhOyMvrwqyPYi66SLG/ep3d
/Gxgdly7A9pBPCKPUZEBFFia0znn2lDzWFG7uiBzzeY5DS2vXJsmAcPcCU79CMck
ybLCQ+kXyfvxvWMYVNfLduoxd7ji7Ga5g88/d0DsWJfCxugIjMjJSP6a8fmlexXJ
jI0MMra5tRAOOq87T9816hB5fDjvqKUVPFYbvL8hXIqlpvSMJNJEaWgxxvHwPeSf
XSpakcgWhL+AvzaotQYgMAHPmMMzYyf5SI/6LFSqLN1SbG/Cxg4PmpqZeTfjC8Xr
6STf+qs/Y1MuMPFbN/L54i5Qty3L9E2LK2ymV51bog8VU87eGT57K6P0ECrJOI+O
6Gpgvs9mB56MAB4Lt4j/NuELsiLhZPYNGZKHf6W/9J9IjPOL7AA+mthqXStzzF6K
p8X+2NwHT2D3dlYj/BYA1jcLSU7/dNww4bGtlZRZZfw3mJxh5yx9/yAjxe+vTUQF
dEPCs3n9fzi7XtlxUGM9HRlBPJJ3NFqBvAMfLA91wAWqaXcEg659qLZHy5vYDHmO
FwcEgYlrMpkIonPpYJN1fX4vNIWC1wG65ES0ro0jg5K+t7Q3Pjt1Lu4jL03GOKFP
pYW6fUB1lrrsi6WdZE9aHqo0pNgQT92QbbWW5j7gHll67TeNEA/Jx9YwVTlzZdDh
i9/pd9pVxxY/hNOI0/0tfMo/uCou7jDu+peBk99+8zam5v/hy1aroXvNw4oEVKTm
LAXC75wB9YOCwOwdfsCC7RGThpLsklaNRm3uFh6f5PCzEiHmHn1p81yuFr48Jd4V
uw5NV8vpcrGfRKQ5HQAyQc6PpudSxIwm5vZ8mv0l6FTvjW5y+SK731uLCW8ODZ/M
pc+lt/KpCluIbEl0wtMyaMxSfLmm7DYCR/mfkZ7O8lXzn1grX0p21IOT25Rnh5E7
XMr9K+eBS0s+2V9Vou3ZdP4Ej0dSZloHS5xC2h7/gYBzDFJrk9Z0RNR9600NHFyo
YyHklkh82Wpsr7UZHk0SJGcHdvX+OJ+ilM4ayzBHdT+JwuLUPiOVqJbOmhfOBAu5
kex6wiFHjU3o8LmJqW7vYePuGz/KO+Hj7Z+QTbBcE9Gv1X4F+fwx9Hs/xImh09PA
dkhUn2SqgNNXNDWkl/vm8OuKSBAlSyXoegHQcSmPm/IIRJeBcjZ4SocFkMQPu04d
E4zHjjc+h8ywZQEBIVlBlWLwrrFEVBCSO2vjYoJrKkICYI0u9eO0cw1mvKnUdOlg
VFWhZFORH4ON0BcZWJAsrgGWj+HcA3lfggrknSw7WjJwH6GyHk4cyEptIYmHS/0L
gaDUY39YUKpZ1AyX0kQ+Hz4ZDMofnxtBZDTOMVbuJNgSwxRD58SHHd77lCHCox41
FUbSv8J65sgyA6rdXhebHl3TG0DRjcf6py6tGg5mxU6U97+sBylEP20ID57yVR8l
JXoHk1TqPGGWLTegDwU+QIr75uzf2KoksZZTdafUtOqcbXCQUHDV525xBv39Wi4C
FbzzZmN//tr8RagAu64WecqX0ldAcJUWizmG6G3B1fuSODVTutX5XBL/d0GF0xUV
4Gp/a/MsczLhUXIxoN2Ms1AkinIREQ25fIhJ5zpQFkLSp6uY10n/SrLqRaaOMwFM
XZoigflqQ7HsuDBtjWWxTfwO60URwYHcEeWzZGm5mpd2f5BPmG58rhBfbiFk4Q+t
vhx+veFfow/IFT/Yr+dRNXnVUEHJ+gmblHbJh9X3LFCVqmMdEUwLrAM2A2+Qce1Q
sgwBYdhYNbFm72wjLYPP873zXBJ1rpj12u37dlHejadSLYaBt0fGgkieNVbThK6P
zmLSacFxQ5P867K5f2s2SdFrfQJX/G3WpX//YFZ8VU3o5q6q2W6P1L/AdTdfIQXE
+ckuIk3EsbBF4I7JTQt1XNKMin4nMof8VSkxBDhtW9UCLICyBbCWFxAVBjC3mVpP
6VdFLo0okNDB/utiZNQVcJQv46Lh7qQ70DV94iHh/Fb91S95PprnS3FattI1+/+L
+4MwbTskMk+ys9UfAiCEJZxHtggWKSl5RLU9h51dSVCIAXiXYlskBLUSrq/QjvCd
1MdKt1pgQtt3EKsOXpAQYXp3C+25LZA9rxsvV0AsE05m1mXWmZ8srgcnRHdD/NyY
66qQEW5sIxG0O1Chwunut0UbC/QT0hwEvLxQ/is9NQiux81wvyxT7q8egrCJol9D
SQACCozTCM+U02LIQEPpZ2sopPUtoHjQBrvPs12cCxUBimvwnNMQZy+CPiDgWIN4
XuJk0jrhyjx79VMIgbvECpoNqd1za0gEnQTCpy6A5lYMnqQ14OmWoD6QRIakCUnQ
RKuMR7+uU+txkGI2TLDdm/WzU/fLKgAz7utRmGGb9v9DZ/S72nnUeAk4zZ8E5rtQ
w7ghnWfp3BGuSobSAHNgW5T5Q6Q58qklQvhfx9oI+5Ta9ndF8N+jwEf6LgQnHqbB
klnHZXVxNDDUK9rVPPBVwc77wHZIwcFOyDvRBAe9D7QwSVAw7EBMT2vFrRacWKT/
zQn+FSbI0Eer9a5NTdXKpJhbDZl7z2LkBiOQwz/ltJwsUwwoID8raA+zRq6uRK3f
r1mP4m1Ilt+S8F8xbY215OMkiSChOkhS50qAhxE90dqdpYkGERSqQeYll3wbW1K5
jh3Nt2XlQUobhayTbU4kTjLHxWDdCMD3wYTl1aXpTII1OqLfS+jVFs5zeGtklqS9
WVFGKOuaXklStJZ/8Ca8CmBZ6SMwUZpXl8zCJsh2H2XZT24nZ/nLXW/rjqFemHdX
xLdB5RhG5+6MY53UdX+CZcgSm4OcSxknzhVqVYvlyDiCp/YEa960qqpykSqr8QAa
zhK0CZ9VbHUdcxdsUSuJfAcLJjJMHTNuDgWEqLK6H5svuTEV4d30vPmGW0cYpsth
AN1ZIYgdqh7cCd/uXxcMbtApXYwYB7Jnk61+3xexWXH2z728EORAP/2te2yPE73o
Jh/55FMeH/ANW3YL6Rz+q0Tq8Q+FDy9XYTuEIwmWrmNHwkfmceFV30WSsW4s0xGr
YxEtQkq9BVx0i7n0KcpcNHcAWxOPgSe9aTTKHH/ZHN0hPDNlXYwDjawPn42FM2M9
MvjhLOfLTZBrDQt4mjffvwlyGJ8+7vORss8mKcEDQUm5Q3egN9EaSE18Hc7x5i8X
rOn3oadr7aIlm5F6QM2/i6d8lHKnHsPdHpKMX4a1oFLdDKPLtq2G8dC03eiJI3KA
2X1QNpbzZRBqHXEh5xArGZtOjK/YOfKzQ4FVWzwoHKnjJfGcJyCsM2AkE597m38T
/CtRUez9OGMrdD7hcwIqPmtFqovd30FYSIEC8P6hQxC7icBEZwwSYFT6mKPVEZ1j
/eA3GedQUSOPA6QtleHcGvzqYdKsZSYpi7be6EZkTSiX2qaC7DGk0B43Q/gYXJEc
vebMrCh1JLZOYXRaXL+qGhr/7xr9tnn+c15Gt2iYS1e+dNblHWUyQiy+bEyahSS5
g5Mo9oKc74GXaL4vIZHZ/Zz9UJjiAWmWmcdI32cC7JNJO9DpPc6GZr0BkK5gCJPq
jViKWPDQuH4UN3Vy3uAUeiuyEhMqrpoJP5caxhS7WWULT7GeRNlb4At/S1cEkRsN
ucyLBFDLCfxksycqjRTVxqlEWa0aGpsurM1FHLakE+QRLrMxuGX1IuQRZnbStNUn
OKMRC/zbgTALjqeJ+bYq37Tz/Wo43lgj8S4JVgdAcob5Fyx5Pw+8xrqkzDqDIFlo
ng4D222Hz9GHMMD+K3Dfif/+8SykxaEmWiqH9WFKzdObYVml6v3AnLDxOwR55JWI
N1jRRoZWFDOK3Ae1c58vbB6g/8tzUSkwMomzHFqom9FnHpfUQuj1FWGdNH9z9xdf
DOH1r02w4MTgty+fLScMgSIQzHQs17blIOfqlcHZJPdKu1vdGOoLvqJ5OaOqxCUY
bWgqEMEjWBSW//ohg3iDbBwTVtHeY1B9eKriuPIJodx74m/hUDtYyX1DcSQ83wQk
3KjzLd/U7HQGWOcfrfqnMr1RNPmIj60xKa9M1wJ3iHC4d44vTkvKOEPZHKUxhWrx
qv6l6S7qYYK+85+StK1YvH/sUwP4f2YYgmEq6pi6V+5ntCADzfhOCI14I5Ri1xnt
qDK5kKcPgcdbnfu9Zd++5cVxlgjMlJgsRvMgn3Alh/lwWzGRW9memy4YHMsq8kBG
UUGJxmZHi/GoRPU27yUeAvKcF3QUzlw80jauRGPwAQhWcE3jeHRBFXufq07w2fh1
PmIx+e25B4ujL6mlLZoy9AW/2yYzdmdD1++a5YVjqcqRDNaOCd2eVze6qBs56Fwj
1So0Wx/WPHMmG1sakDVPiwvZs1cFqPiP1b/ZsSetm+xbv7uiEKXyeN9v7fwuhi3X
lMfvT7ceAKS8bw2VlGgSXBpqU37Mfi1EGgbrle11aB7qg/LpNmjkMMSxrOgyoHic
cHnY9lKHdCBKO4ZV/ZooHxfSVw3Pa5aiZXtyCWPYJ0g3igaxkXvN/wwYTcabxsBL
+E2KwqKZEaMOgDDmy8JFkqGnOho2fQnE9fqN3z7v/tBriNBqf/E3ZiJMl8rJQxYx
kY6IyKupnDpZzInzSi0mkCnCNVZoyKF1vXDHk+Rjg9kwHFY76KmSzexuBe/pT7KP
XdQk335Bt93jEHoDUvtRQSJ1Vfmtd4eaSo47CzC1lLB6FwNXEkbPREne5+zJg0ZX
yHGeBf7xfsF3G/bjuyHuNoXi5siFBbIQmiqFHBzWSfhB6+7k089ozl5k3mD+ZSAL
xNSaSuVA/BoSWPcwT4yTavjOsIJlvmUOQmwz0MqZeVCSxs7QlXxErd9569IdoTmN
atteqssTPD0Y1QbUr98gW1m2BxcHhBgV9IybdfdTTBOFOsrHyhjayxJAwz7lR/Cc
n17CjfAQbwEwuhzqAA42P2b5/mzgPodd3AuMUv+K4lMB3vxfz8NmjBUdpjeuR28h
TlrAzeGNFIALqlEAjy/CfTPkqjvT+zRtocKl69viJLU2d15yVUWMfN58+d23S731
9RGodOSk7Tav3jAkF5Q1+oqWHlF+HwOXAIGqOAZxIUIECQnM0BDY0lIwpdyG9NvJ
D2UFnWWJ8qdHvndmVONzAMZOMemHSpArvk9oxgvCyHGRJ9S22aMFLFE36dvJeE8g
Pk9rVTx1H9kuUQOcAwAsmqF7W5zSRQ208O999HWSfJAgZtf1eAB0yE57UmQypLq1
pb+FVrH8vrKmTogj+lnBBXmb0oChpIX0CGgC70iuliOVtIXeIA2YMnx+gbkLMuJ2
WUHvPR7ZVZ2ypsSAQ0UAqiNsCOLc1vcEFaXjwnxfXoVCiZjXLTWhswgXU6q9HBNU
AmKQQYaA74ilL92ouqb7vE35uTrGvZ8+VLoLeUurq1cYYmT4l0WORStv9D6Tejf9
crrTWZDnwkBMUT7uhxbTQ8fpibY113Tur18T+skabFrqeYGdkQEXORCQ49THGRBm
hRjAo/E22L+M1mXHlPxfglroYKE3s7pC1OKf465/JNXZUJ2z/ovX503uBD6wtvov
zMeJz6tHEcBiNZyvctS7LPJx5DMYW7Mr9cs05qGlErRAk031ino0Mwd1WIm6a/fm
KMXnIBFSzltUELl4kXQQCY0yyNFYv4d3CP4Xwd5TmF8kZcnf2dqsarqlPY6AEKRz
+Wj/MjcsElXpRKfPB8EFW3yim1pfFI0pBUZdI6fIsgQDpCr4/llHlEajP1NDCeUG
ixEQAoGeApSmbBjwi3UYrDN12KDNoKoScwh1O9AaYmaGMMdefmudl/cedB8g0Hch
lbHG48mc3pjX1wFxO4QOo7QdEgmIx5kTe9VSHQYTlVtx8VJY0ATkOjE6nV3bDrOg
F0nk/cAiwcqTRo6Je0Oco77NFIREroPVi82qm8eV6O3eVS6j20Sc3S0Edw33RZvy
8lEdiI8MoqMf38Cy0zkRVgmG5kAhSaRaOD3y4hnAZpsseKVHUZ+2RBIYBkxpYWTS
YRTrLNASEY/XgxQrUtr73BSBC3NIiPi70yixcwGZBvWDv8VOyAYguZX7K6NBuCLR
VCtkazLmGst5ne5nVI6oULVH6APmuLm+sdsSsrHCBW5YLZJNJcUOJ5BEBaJs09OK
2ck7SCiN66J4nxbmO8lXEzRXRGgkWET/+82VEY7/evQjyrMgkSAxOCrFTGgmdhOA
t+rPMkPbquwx4l3zCxRzD20+vrclxBZnEJfIM6t4QsI96COJ/ZQz1dIj2ohcP4b9
Xh6yTxqgUOMSGhYyVZJuKXyq3OPty9AKrZQeHSvAbkNE1Qvyif47co3FFytKwoUK
Pdj43rl22S2NhYPtPlLL3g+/RX+oHUEUx/pL5dZpBjfa7jHXrspQRfP0G4lWxXFf
qpWMCSWyFsshWhx5/SoKM+v6SuYwgLdwgVb4Ws+jgX/9528yJTIVtg4BINm9nCN+
HobNO4WK/pdkJW0Cp37+3ooUq6H7Fbi9rVz+UOrQE0xiDfBkoxLqqhGUXq8W9u9g
ZwpaE7O/uEVFIkUnQgA8FJPzf1Ulo75VDTLRw6gJ5j+Ig9J//1/MJp0Z/QhojTe4
+pwN8u99tBO49IW07LD1JAB8WnLRNRZzlTOuXAkBsPc5SyULwu/byaFWgDeqB4Dx
qOUtSTVHX53btbD3oiPYTOZVGSaeEQSYhGe8w+qXWmnXJJQJNj8/h1TmBw8BdoKK
Qxq9TRE0hXNe6xVqzU4GsOwKFl9tmXkoO6BwMCQkhTuL+1SsWWtgQ57GE/TVwFCE
bHus0F8rCUy1sv9pkdrs3VPQzAeXQZjgeD5u6oSP9laltgYohk88YYg5x4YYpGZn
WjFyNysodicUMYblwylUBVH5+EKm60itn53ikJFzPszGuAKT+JakthayBDJ9QCKI
Oc/d2tRADm4MIi6N7GoUxg5Li0OUu2qWAd8ivnnzHHUMUR+d5G33JbfM3rYo7axl
sHOCTk9zpW3kJtuGG+NhawZBlTI/zG440tpSBn8s1MPlxmHPLtkTHJ8eOnpjM97Y
t/dDz3bteHYWN8C0nYh2JvFB4z/24UC7mkoFxzAXslHkFnjAZBPZJIFW0LWs3mss
TsLM9+ap7zmnHCWPDDPt24DuB5Oieh8LSJEvucEHJiIegRKI9UkkM0XSWzjv9m2X
QuPtI9Ka+0tUO1A0pFayFYVw4pOgpBj/atCMZ2XprImikgfSdGsmz7vPuHVyuNSq
5m/usVE063bgcrwy1jZ/ZwdowtDSJdIbm3+1W9Jw2RQH74hZKT4AJcysD4rKu137
W6TDx2FZa6bRYIZvS3Bk1LTe2B3KXboUPO6ecPpC+cDlTMYsHvgHYCSIP5aRnbUN
X/BurKxqjyJsfSRob/ayqTyUCf/F8L4TeiUkKVs34Ej42+NhVXa03LPTKHzXNhlJ
u+nM0zQW8wcCQP2hSHXYQKsneythhiV99cxOziRG6STtqRm0SIPvzm02L9vzZ6EM
oSeFt4NKakDQQDYFYNHUgWwQfmilxIpCdNAKFCJXYeww+ONouIVFpaE8kcheKSoV
636rikCRciNeH0ElhbofmTyUY5gR7xAMVE7Encjo53h8/3s1eDmYd0qRDvdcPV43
yolBsslVxXNFAtuzZDxnhCN47g0SHVl8QpKOxuwtMYpnMPbdAsZlzZC8JlHVHqpV
uu7aPDyEscWLXO7BJNZ/DyM3p8R24Im68Gu44UX/6lkj2SbbvDzloKVN/Ja3y0+6
xiRMTiG8meUwCyiIblKkiDPm9E9d7NLh0ltTIF4ecn0HQimmKKEkybEjgsa/7LHt
KhNISWwO4YHR+V6qdKwYgoTh2G3nAYMR/xICjSyFaBAprRCKMGIlAOKF8IPInrZl
7weomUqA9QR0XGGjGtB/Z+hMD2+rKuXMvQUwvovvRqB5/fFwh37bGT5kEHn85ee9
bdrDKHoauS7QCYo4SxVSrsrkMQnlay6L7GK0fqVO9eBhSaM8O+BeNEvfoqd1zLdf
EixN7pa7TmC6LvBqjFKA4w544aOhpSmCD8i6SKad73dH5D0vW+LJg8u17G/sRzVt
5FQt5/kZ7M3YFj4LyM3ILZ4cHInh7TwvAmVotuNv7fg8tcXw48CH/NxUJKgurdP2
cHlV4zCFJ7ADtdGrFwdKRwrNKUidd9AjJXGK2jFkNvMCS2GNJQkwuRY0vk9UwP8J
WFNN/19eQCiYWZkYVvQuxigyXCAEW7uikF7bRpfQ8pWtNlb8F0c21dnbEs/f0f67
Z/fVvXwfyG9vCspP1JkJsJQcG/IKGP8BnCcMJ0cAKg92K2fpjZ+68trQzXhXcsOn
UODucGKY67y0N7zaUmlZgwIKft8GKYJkvksIh3dT/0pdX7WnjaBiumukQLyfSPQ0
9U6lw0ndun56OH9GzdVg+kuNndoLqxbL+gpbWuN8ZinzhK/5cArJxtHcgYKOQS1D
kztCfxXFy6AeCFNq5Phy3eLe6MkKI7KQ1gPcWYocQB3nJOubr1qCaWucTzaUFNAl
4i7QuEDISRP7PtJIduMycIxNJp7LmfW4r1WIWdYYvbmI4XkB3TvwmMaaPHFDW8Uc
Ioa8GH4gKchuEzdB0q0wZLlhb7qS1QAISI0bEuSlrbaOJae2Nk7RHJFnMlVScySA
QXgZ1yBi5k98tO37HEEVKFGNJiee0oeibl3Xf3lJlIjz8QmctkhB8ndtJHvJvTF2
+n1d4y/E+LQNbOnHmGgqRIeQTAi+94m6sHiCSKtDFw6tRDE6BBpJdpRsC4E94b+n
4arVRuyHDVspJ+bWF4nOVgk+HT4uvqeapQLiYqD7SmXxX/6ZcIm84x9bIn7FcQ0R
THr2FGxIAKYFtSpRUHerCfZv/H3ccm4oi5T9kmZZk0VFSz9DiB6/tciAvGh1OvFi
kPNFt7dUzX5pdAq983ouN6QxTD+7ZndhlhnapyCJrhC1DvK/3jcE9fL0DNITvKiz
rKIttPc0PsuzDNHPXIfic1kJgdhNRjr1HPsOhVhde9UZh0745L820+mw8A8UaiMh
8inL0+HtReIlpWNaYkikwdl9oamKQm1AF7pMcPEspZYtZDSQyeNRVahUy4HZCDxg
vYAWbGE198riWIxLyI1IElSJFzAobi3Q7tymurJKt1hB1ZTuA2TcYfjI558X+jor
4Eelm16l0qWf+V2zihveajme2N8nArGZq4M4EuFgXd8M+CEB/U/r/EC3btORRomf
38ttCJOMZ9wDYDkdJb4g2CCrHpa5W40LF4rwQ2AkZRb2E067zneOYBU8iZc+m0Od
Z/sFvgzMeBSaP2lJd39x4Q656RbERWC4FuLFfyqAbjTSYTZMItGsv94//egtalPX
gT5Vfty7Vtvmn2uh3uBjc2vTUROaNIymSHJdGKPdt85IzHC0mpEl6nNad8nvN089
fvInEFHI8FQgxCkGieXkao5Sd1xeQQyeJkk5RTvHHLJfXayhguMG1eu4tiwIVasd
9wMUs0CwieIF1dWo6bv/vxVkL798ITto1+2Dp14e/X9A4NeeSBeYKB4oetkZhSFX
loqocvgulfBHn1EBegQ2zutILqRK8qRNfaXOAuZ3nOStx0wuDn5J37uviFjvDiTv
TlLoVhKvSajfuBCjzePi86PRH5vPDhl/9u/qrDXKvD3wYSxcVsZfaBFS6nUNXrp5
pe35OfYmRu7addCSg4xoL+YjqOeMlzJend2qmOVmD7D4wBXijqex4GVVEYmCtRWk
kBdy43qsEzwScavJ9o43htxIr8FRK5EphZEV3zQqM/wsBnn5wK3SPufZmnB8VwSO
cu6gzt44OBSjND60K+RKb1dI2jDW55cRfl8+JZnU1q7MZoF9lbx5Z41b8I2418pC
43Ru7aIgUBG1T3CDhAvKq5ZP45vmUZ1+aN8aJ8AIXDLCgTywWlxVXQxE/QVLYSdr
tZr8f528QW0meSsueDYIKBwJHenzPJyWu+UjySM8xnGqh3AabWKhiRCQ8TRck7Fq
yt6/sCIMEqYyhlFsd/mj32Ep9qctaZziEkGjNkq/VC5BLOFX4/xeTAlgvx2KKn7x
RQieek9vMaWi/P74Ds0ts1QuO5P0tUpTyBw/uGbSMtW9bBgM9dmU12nE8rI/kJkI
daV3h9576AZNmW/vu53bLb5+AZObkNDOT75yW03aNBhWM7dQ0QS5NuwHtuw5HqBP
kbpe+0P6JhBijt4UjPBZk7kGvmoyjiVCQ4gK6RrfA5I0Jb1bAPIRMvMKOplck3mJ
/MaH8hqelWWe3HhJDj0DFHbw01dDP8SQNAol1tGxMaB3QQ3ofwWVZWz15GoyXas6
tftXjEe5LpkTmzHiYx1spwb7snI7NEPeiWITn2mLig00iOwSEy6LKGK9KYtUlGr5
C5UQUMGRCc303HeDwdBqSBKCnzGlKekGmQ4ZpMqH+0FCxk+I58MDI1SMuI+5Xd4e
0ZWOS4ApDV1kp3oqUdSjNPJPBDrYu4+lVwXgvMaXbrFgvPkn1QJG7Wx6I2qm1EN8
2fwYftceR+fKIquOrHJ7PgnICcHxY6w/tckcG413nTVfVFth3bKt/nDdZiC5PK+4
joITqppdT83AutE/kHpG0UAI0WF9lhvCnEwzOV8QxljedThSTTqgRmYcuK7Ga42t
95MpYrK5QlIWlLN9O3d2m+AWLtSAJKcWTDfCoGCTHP0Pbxt3wytywwfzMwe2E0zO
IlIjpv5/xS6bQYcVkqkK7nsYuxLLSsIfVuLVeUlk/ytf4aF88A08UisH0mcZVU+e
UBu7jQaReSbWMDMXhQuhEbtV6jlwydle2Ue11mFCJVU8FuSofH63vW3l6+uHZbdt
ZdmA28LzRixV/0HclUguJrAYdPa9Ik33nOI2TsQOEa7oCAepXUW9sylXL5hXOW7w
Yf0Hrmsr3rVIIR70YcDBc4+/V4W8StQzv0Uxt0UdQXzOlbhmFdN05MknNvF0WwZl
xWOa0FJc8gA76aSwzFQKJjaFpLLsnRRmnfus4NGS5jsAQXw1f51PyZURqegOefNU
NgvsVB72N1dl6oV6JH07nfPraFUQ1vNqkozxFidcLelkrk0nj6LjHmNQV1Ooq8f5
KFAMvsTAum8WaWXOCABKp8P2ZT/2c2z53MeuWGstXKaIEagVlcDQEB7b15eGp04L
+1zWK7jtRmZcM7a8gTNDIMMG3/AbzjoAp0I4N2BxH+ckpfP/q/lZYicQZwHiMJRK
n5+lkkpp8CKm90zH7vRLpljotmVxjPmWycbuYqiJCE4LZ3x1u1SXi8Z9pUwMbK+i
k52W8LVF+1mwRitSDS4Lq7clttBgj12rbNrG9Erezaj580xF8hON4lboPYJQmnsA
yaZ+ILLI/svp9zfQ6XhOrSlvZmoTS8NPTY7VGxLIZvHwfAhay/pbzwrEgbv4K4Cv
iTR4TrkLEEk1jcxqaxcgVpUTHuGF+GXNX+7flHFzDeK9jSg7WEQDWi5LExgk2aM9
iHsQL1mbRzD6eEl3HHDzIwvpwFz4YiBBFI1S9/IFYexfsWdC2UM1aJpynOrP9dCW
0WzqePUrq8Djnu6dg+DcZHdcY25fEjanihhurY9HGnNfb4Yf35axPUfqtAXh7a5K
ebIJlO3/130kXOsdXLFlUUyRDQYlph5tkG3SW2qbhTk0KHBEVKp4ZZ2ziLtLQ3ta
FYFukHwzmhfQ3OLloMXixRZhkDUlExUznsLaUHYcvDrWXUlRXs92zEkNNRz228eV
bC9Y1S6SjhAWyG5THAun5aRxuMTZgRbw5dtI8lRrRCLYjI0lH9ex+GwidhfnsYx4
UCYRJfwvSau2zLF9tnv1+e40w2K4qfgKVPb8BMXQBa5Hf7HmSiX0mJE2l/JrCdK+
mCNJhLlbyT24nVjoKOEJnfj2DSWMdcJsLjWNRdgre4rU4qs3nSOndh4bQMwmB7eO
yxlgyzG2mzyfx6iCHRc/kecxhdOYVQIYCECji05ITRAXIDqHAkSx81MlpbqBzlVE
990L/OLelarjLYwn86RUHK92drj2HL0OTYMelfRDQj+JsQ6iYwZ/c7mqxlHdOwCY
Ax9X/4pICIdiB0XuVLr1nxlWVTRpaLsjXwNhY3ku9J1VaN/nM079Puri5BK5GWa1
zseePsgG4N7Hy1EzZmihrP3Z+pIFFKqHxhYW8QXl6hvFDrJ/UyMZgER36RRcyzut
chjp/pnRfW5rKYj+qrOB4UiBBB8qVSsYumtzvGvnhNqQ1eQAjtNQvop9J+mz+M2F
D3ArC5nryCE1OYvhLfjbGCl/DjtEfWU7uWx5m2+KZLMjubNO7WFP8tDrZb5v4viN
Qk02YAIpRgVE8LNu+sGwfbVUKXuYBiAZQgxFluzfryAdMsTFl+Kh21nFSZ7h8Zwo
CSxQT/C/6p1QzWWbGViayi2GveiXBfvDRfQbiBNJ6xgbATz1xJA/6agj89f6tRex
vllMCiGOoutcJYapH8GZu/Z4Ycxe/LW/zQXRqFhebYZ6x8rZDWwzs28dCyhA8fuM
Qd0tcWKltJ+f4VjMuUA6pDfQ2af4aDVk60GJ6VZFgDDHWabUEc4v3RTcsYJO3Hrl
hz6l9xeog3eYnF1nUh70j4z9uTeRCGNKoR5BX82jpI6AGbHJDoL+gxy52uUBc3H7
3hNjHszZ7vwA3AYM4pKNk75WoKy3k0OcTaXHnm0e34AjkkeOXSC6IFKtq7MXMuDo
AmdCjrDOzhUrmLyKafQjCqI0R3k1u4EiRTBFKlujYqq3suZnq8KNpKLO7wIBIQax
X8i9Ua4/TmSMYpmx5w64pl5exJHAEEiwC9gfvxclBBE3+nKkXrq66pGhiYdFA7FI
k4LaNNSKUGjfqq40VlQWwD69Rs4Ll5DKwTseedfE0j4yCAYT5DlA7Wk7zcr5ysTm
gw6SlyHAnjdM2lGMbwX1qo8nx6OPfE0F3LCHxcAUD8URcIhrNNTJVAEKX97QKoL3
scf8aDtKW4YeB1z4k2b5pgj/vbkfIP4rkC/xvSgUkhEH1gPAQkOVsNXqYii9iWfd
+RzbmEGoasBRziP9mITiqgDmpop2TZGzDEpx/Ib8OtDDwO0gqnLz0BSF0G34mqSh
DSCpYflBu63iNxQ4dxSJzq2LtPPrF4IxtfmdeDGJun2hVI7cDkjxe/YzoHKveeeV
sCI2BkRj1508GqjASDw6XsUgdCW/bsyyMR+sSGGg8BD+szpcfsro6sZJfYsrM82h
Zj7FwAoZGEAo5DBrNfGSJfltGleoMBSDvMtsv/M6VcQsad5Kk9fFDbmEyX2UUOGG
aj4KtIicm1YssN/8TIYdDngn5BbeVuKPMAjNB6Uk+KvsMjzFwSfI7U8LyO64upah
XOVAoEMYTcc17diHUNwQYWMEMvv12JmQfQC6GKU3SBbGxvfudbQmVk0rItte5b1C
NDERyBXB2aectqY2pxyUkIWymIw4LjMMy7JFZpWvRExos3Zm6nUJHfG0FfWBw/ck
KMckbBbetsKcoHOn2Hl1X8SRPGMEfP/ip5C1N5I2Si2ux1+EHAMNRSn28gIOa9gJ
vYplseRpTZSyj7wsFuqQKdrNS9VWU0T23ZdKDUNWXm4c93pp04Q3imZy9NXpXp7s
AQIa4a9N8di6BteYvKdiYuHiez4zq6Q3QkyeZFKBxkyQf3qCBr5ilJqnaAyf8SsT
p5hljmIm89d7gxOoXi4mUw4Rn0YWzFbHcsGRrqpL4i84j+LOXcxPC2Gf1hEcG9oq
n1JmRbJLW0g0D45PsSjFIc+ms2y1zGACwZYwD7PXY24WwtcE1hMqO2qMFhMaO7tF
gPzxG4PiiybqaDOLR0IbYjkYEre5VOT/uHrUw0UVl9Ur8VGmVuYuz83vmrpRu4Ot
csA+T8d/FBeX4jvL+MldgLzSPwCJXAcr+pWa4r3tLkfVt7LV6QqTXsacjr2foJ4W
NRB4KNkSgX5qCOTrl0M2woIaxLeWcHMoPHHByVp8sSqKgXuupuz5s1AqwKihn9u5
8r3EF2qMou32Yf3KHOo7oqQxUa16SebuD9oG3v3R1jUDR98m5wfdDSbYH2FtFrFF
kQZjBw3XomwVLgOCLSgE57Nr2O1riJpU3gwjwkZt+QE1d32e4wvMQ0OSgwL8NqQ+
J26LSuk8FYimgfi0xG3C+ugFlMJpWbl06dju5otsrOASVeJ3GeUloOhVx1TAZ9Gb
dSHmKB4C4rQZzegm2drNvnzaWlF2bpRE8oulsgKvb/N4Cjol/jueIhdTTVDT5vgu
n3OHh9IIzv/0ihknXw+F+Vsh23SpiKkt70bL3TbSOMkwm1fvWwKkFQ+kCydZ2s5T
dW9FL5MetKywLoFmRJkptSKMUVj4N9guUzXWhFGTfhabdipBmE5a2k4pWFNwSiLw
fypvibzNAcNsEWz/h8wYiapVvXCLprlP8n6mtvWDYDbnuyT/0b9EeS4xnK9UtV7r
vLlZnd+xBvJmZUskbvz4QX82zGegQ6tmlTdVK2vtKGYZ2DLR7hHsOr1w4SQObv2e
rupD51jkRQ3KmnnPOrohtH/tyWbl6Q1kP9XtJ2DzN/64mvoPJ8eI4cBWYTTUnYyw
116jy5jQN/iWWQCDhUs6YX2NZfvPiAGJJnL8Zg+ZgKUd8rtR1hkeJ36nf1EMgZyb
4GQvI9dM5pFIz1Swahf5RWaa6mNd0dKg70WnLU9rAWYAU/VEnm8aVcCSt/PHGQK3
bhEfEnHg+P/uEREk2O7orus+eTxGhGGYiMbHwdCkA4MU/9IDB4AuN3jMw8UQ5wog
nUpn0+OY5TSRH9E6nwzCI7qonsfFXyADjhTa9xjF8HvZazE24ZjCqKVPrIrihZKE
WfMDQPansJ+32Dj0H90HIyF++LkDcIJMsMYB/ekLYdKQg/dLiCGZ3eXml9S4bmWm
X4vDvtM7IhYO0mIDAXSwY0rIcS52NwCsP+Bn62QbIqYyvhOfLRS061bpKuevQPiA
Y3HvYkYU2LGb4yJV7kmdcomqd+ZbV3Oe60RPdpAkiLjm4CRNRhJ2xrLUj71LNHZx
ik8sdT7pAh+og3YAi5r7OqodsOUa6m3LFdVMG8hUl0QT6GrCYShUD0cISTzFTuAO
1Lm9W0JDQp6I0JU5V7jnNpP3vbsKW8ljc8SH6XrBsFI2qmbEnCtFrZN6TWfNFvcz
y4y5K5okp0b2nZsIuItDzpv5L/CioDZ3nTJvAmKEY9+fQ5k639aIMEicAoLMUgDr
4T6MIpKQchHtu1wAO2KT5Inlv3GDKHS+0mn+sxv/igT3xtJOoPLf1NCZQ+oVXGAL
FoHFpxSTPOW0fr79t6XHwD9Qrdw7u53np91x8MMbfFGSr9+ezdN9LV/rq3MfZaH0
7E80v01N2CzaqzchoVUEVmc9K/o3Ef8LLNSNblCI0P9ZhEL8DEhc/Q6lAwAdsvtS
6yu5gTkLnpRROGIc45MuAZwuWvE5NEhrtGFh9AMioYJqTr6Z+1Ee/KNAjPe6a7ir
M8oyFHyiorwP1dKe/bAMl1V2Zx+7qhPSpQKrXi97n513evwa9p66ZZswlVbp67TJ
QQaPp6QKYmQGkDA9krJZH9vBrJystUZ8lZ6/oC6W4WzFJRdMfqKXTyK7e2aZUVT1
W8EGUMF+CDNfnONtN6lYQhHJG9Hm8lGP6GefNyizJGZc8Shzae47s/zZAOfPInce
oWEdBK259y3jZn9L+g4zwAkZSKEbMBoK1zCxs8prgBoSQpVcu4DpCFCW0TyKPKgC
bugJayZF0giDqOXfVzh8Hb3GXs55GOGz4rumL/7RIlcOnGX+3SCbgOPikegRPCx1
R2t6dZaBsVaoyXY7bHn1zOnxywdDGzpH4kpOtuGc3qkTfpG/9TTtU3b56dIKo2cp
BsxjzV9DmgZPhzSGrWYq/mhKQhqm7kVst8ceM5WdQ499CVRNqllVF+CIwhntjV5A
+bOZO6FfabyPH4yrkr4UxrMC+92/8rMfdoMkt7WflxdQWJav9y2tobejiyWsvyGk
srKY1XUZ4RzmDfkQ/ZQPr7YixDD7ELQhr3KfWr+LaaKs/z3r8v01+1pQgF3aLcEM
aG9aGNnUAslt3hWZTY3oBjk+6mqJQEAb7RzSB4tTzONa5rh1I2YGY3wWqc/FUdrc
qPr5ZjBwRBZ1O64YMJ1qtRSAGnCQZhyTpG6T61dZT4WxRe/8z7w/AtDLAGQm6EqN
T+c3j0FVPmht+6P1yrtVxYekPJX0xGqw+Ze0OFsShYJhH6CHvgW+69JCRtdXuw7e
dqNAxINMNDaNeoghar9dtZ9j+ADZZOoAIYC+diAiuaAfEovC7VW1tlrgKYvIuCmc
0kNK32eaIxk6NwRVHQaxrYYuRfqK5mTOk7eZa62+sWpFPrvj1VADOyKkl0mHyH0/
MJGeggWIZIN5SKMBdTAAMDs3FUVaQH64H9/jQe8LSfvyckPNirKK+/SGEfNgSwlx
yeyyEDcMJKfLfLi66OrBXwQeX05hcg8lgfkTQyVGpM0zD9zPi486R62Fd5pTWzd4
iYYGkCgQE+8k28EToMoOl9NUnv3lLbdvZm89lEJqRkG/Z7rMVHg0fVqPWpHeQPHB
74rZ1H6yGbnrrF82xDZWs4aZm2QHdlyr/+GtgEiQDo9VzcuanrYUF5Nhb3+GgiEn
QGNC+c78YkRFldToHFP8rvSK/T1Ks9IzNrgBxRzi1NmIo+FoooVXaVOUUIGQjOpc
w+DaWk04EXAWB9BdTIw/h3Ua0GLWDYZP2iacTOJbZsj6DGlalnLjDLQ89TyztgPZ
z0yoZbwSR0POHyJyC3NyfeBlR5ngq2EP3wEGnXhIMmjWRWrkNA2HXpC8e0Nbgq3e
ZiFERzDfXw/UNjW9DOoDR4cIoTSHSe2+n4hcg7bpZJL/QehAHXNFEBJJ3vq3AZ2u
19TlE3rEW2CQ8H9jyRxfFkQVMrthOYPvZ6OPXdWLFhpSJpWBbCf7T7SA6vBcCzVo
qqZDi3OOiyiBr37bmzH/Wja0CemmdbwjT5AW1OrjCUEWxBa3LxKY+1C6LnqDZ7Yw
G3BSx0heuWOBBUXiPXijXdZdCtOUb48hJaLRY5Z14LgDAeMvwY4fOuFb6c66dysw
EWFbOjJcOI5J1jXHrGD5YUA8wo884+PRnzwHzRp+pm0X7xVebIwJHkYdF/bF7uBM
0vB7+fnP0oPCvzVFmVK28sEsS8hpcqTMZSQ5ydczmigQaLcoo05Qt+EiHmUOiBWB
BxWrkrqFw/MEc2rpky5sgAgw56PzMNtkX9M7jiMGABPOl/JHJomv8GOwNuZXXDiJ
A8hR5xoVFcN1/jTwoWDL5SJnc/gU25z1KBjkfMI8jIwc9elYkI+UQ8hR1KvNzd26
+jBUJH2dTMeEzBTRAzOU7f8Khd5SVBtcF8V7BLb8pP6koQxFiih/2bryHt8mi1SO
y/FrMZTFx5+TvjwvQU/F3l7cmAx1WMCR6d0oDozALLtcjIgHLvZPe9y+RmVV1FU0
dP+kXX9EUXp6+sRlY9IVu6atESqflf1KpAubpUbXV5Ym0ygQNsfF+FMCAH/WtBfy
hzUldoaUNXHzNy8TwNzHGNNb8eU82lZhzbt2OceikZW1KvI+Fce7BOt481jS5eQ6
N/gweEb/EZ0ybnO1QnA64mQecUIZb0epm8ctBvBt3UP7d8sGZjbZRtYAmmdpjFLg
WkLzpJAAw474r3pCnM6h2w0y0f6yew3uvW65V7NOhBWVUciKZFt0MNBjJ9a5k/vu
2Qa97KvW7XUBx3j3S+LqCY3JOJgwST/jlyo/asDPgVJ7tIh3eHXDECtjMMn66FG2
/H+6s30z+eMW3GW00dtWDckjq1JnTpLFp8WePQ3QXxjfLXG+VYYyYjX/l/DcyXyb
oLn9QSa9cv8Wucxs91vKfmHykyAzXRoqOhlUtPDvDXD8BhCY3I7wOBz22wxT5TmR
awPwYq96HxZiya1LuHCbOYIe7N5ZOFQA0JJIm38QHAy9HqAgo/qyDhYDo8pjVpBS
wybFTtADLfzo5DQOHi8+Edv4v75Sul4+vrfgNdEP0M9PWoRK30ai2ALD23DXck4T
/gVLMkk4JAsCmZub2iD9rH1cyEBxwAwhEVQMwTfh/FQ36onngXdkdzX2p2mO/wRy
v17LRo++yRZnQhT1I1iGIsgLy36XgaNVb450qtqbZhXZzzlY6Mww5jWJIKD8fmiA
QKlr0Y8wnW003WExkUeZhjP27aLu4MYpWvqEEIwUCsoJ77XOTOuw0fyXnrF2Oxd1
nX6Agon23sENbAM3P0MKe/R11xbcEAJgJQXcSgxqFfU4iIqkCpsXw4gcwcZT1RGr
UNYGOK/XMMRhPEuIFDro7yRCopA2oYGq/yquR0O3K9n7KLy1S41XouBFLvGeuDKn
6oZBY8LTgQCshrTxLTy93DikMK2/tiqySYMDkFSVOIyqTCjvlIq7FIChvYHNie9R
gmjIaPCtIJRnR2xIJ/X4bqqQAQM1yk/kAeK+DTpYiDh/68SdfCZo0bECu4Fq1M32
0AnbHiu03jU7Ue77reTobAQOfZsEAleMXGpmqdRlhLdfx7U5YX1QUi3ieGqKI4nt
6y3jRV/+2M7IBc1mM8o84WurhnUsluKC207JQ9a0yjuSO7FL7BLFPpLo+nnYQ8Ff
DM0mEQBa57DpAkZI/My7TW8H3T2byMplRnSmtMuNjVUzdckyJpueV7H4WtDH3eEs
fU/ch+AEdFp7f+kUqzpmnz3OcwVxTfQcWGMMiXJa1JRIaDDhAHe0poLnFqrygSaD
cupGEEBxBEYniFN3seArO6m9pG4OTFtbwN6YockQQyz7FejXyVMzj1I4MrTqLF6b
nqMZx3AhE6d1Sk0yg/w3CBHCIu0NteJoXeYS45TxV06+8QXwibyTV/Ss6XXdiyxp
lNdqC3ZdVcKF3lk9rJPeDD8tfnkHNfr4BKKhrPKzRyeLf05D4cXNCJgxvC05FvnH
koUxr+CsUU0gh9I/U9YiLhkWMNUlO0g/+rPqqxH3+c0Wgb1jjZ4vrVPX4KO8Tqig
7wf0dXF2dbpM88OMx11Pa5Aqe0hNrvsxrJr0Ml9nJ/nN2EGVwWE/o5X+v/6tlNd7
RC7QGzMMS75GhC74AGsfupQ/9hH06GdHXZLaFqQ00fminkC4r6DBsptb0ChkXwvs
FpiRsXK03W31F+ecsJgUqsx7t6RSy6LqXdG1tAsh9F24BzmaMogyP6l2RZ5l/X+w
omGF4mBLaLKzBcexzuhk5BanQywUlykcDjXGdeDKHRRe2bdiqFCYR8AYqr5FoCYQ
P1YiyS065ExwTWaPZ4GvDPHcK0tg/vWrYympevvHD+KPIENsBLTWS+0yE6KRez4d
70N87Hj/hobhC+FUZV+jBwPWdA4VP97xPnFAXFImlxWOHe4sOti1PCkQahtls5Rr
IkE+lOb5Sqog6KgT9e5TJmg5QsCMxzv0bjA+ocFo9zT2O3N6mU8bya0s035EeQuy
XiGcR2I+xbtLa+kZGDunhrPpmZVF9Mcl4jcQViaFi289FRRXla381i7TNEOB3qmP
D1XKRYnxj6rpCgXF9OkSpJKn98AoAt3l9G7+uSu1Qe4CVjbmG7SgLK3avNo0Gdsf
RwnvcxPrNyFw64+AzMInw+8FPd1nAwpLaeQC2yulI2Htku/vp/j9F+pYoTkQfbK6
Z0H/f/7oOyahzSMmmcJhosG7O1iz0i4Eat9tFSXo0PdLUBnpuwbhsfK4AFTW9u5Q
nqal1T2VBKXho3dO4pOe0qI8iFjYKdDD9bJ/youTzWW3kW4+3vyE6bir13IRap2V
L6IoB7N+8Bd61eVNGSnViI06gw8p+SFgL6Z1if3uybyRqvFbKa0BnVCMsk8Zho25
NQUK8xDOn7qOeu/1UVhXBUdKvXlixkVhg+JTf6Hj31Kqy+eUsbGD/829zz3jUh++
VB8UH1tB97Bc7gC7LJtgqSOiH+PJUZ3i1lGM+F0zwblL+L3wb+zoUGD+uoHOEDT2
JQks759R3snhdjTlPvdcLuMYqAu55TxAY+HwvYhjq/J+XYDkFdrvVphrc19Jrgme
t6CMO5zfph0iAsH95fEAPp7zA/nqsiBF0E+QyRequT9ErQAVYpAL4sK9tm2lNct7
JAluuqzXC0OHAs2czWTOM0RMLZT4v+diB6bTvJ/rT8DcjyPr9b6Po1WKucD3pWv2
HxdlWyxd8K5CzkJ7xiAZkIrrNOiAU1RMYQ7nurtd3YgBr9SprnG7cviQ/rFYzLMZ
utoo7jSlbQ8TsrLa78H9qHZKFGzYewcDQs0aG6avD1V5QwqXwyoOSqtxt+tazD+U
tjEZiR/960P+ooTkddLTOI8c3JURoRjIBJ1OZuTDBTnV2IbeXNquyMf1qLrnr4z+
vnpLhFLdWIV7/s94jZbR8xDj95qJZVinF9HgzY2X2zbezLlQLT17BkSubfaPhUQ+
4sC3IMOsKTDvHHhPhkjSXIwJ7Zg0ZQm9vlLmbKybT5VxVsP5jEmxctocZpaEboxM
GUQGi0NWw5LLq7c1trvGA2UAG9AYEWaNpgJz3MLRcNYdGu/OjtuIKXZUH9vWvrUQ
kKiDJUr/+cu3HmxgtO/2Lp6TVD3PfqJGgDdkcRts7A+5eWs6cy0NcOFqbZlgyzey
7u0epHxUJcDCPnyZBrFFI3hdDBUyH7ExJ/0/p3ipJk1MsrGEoNfEcckslXWvPrAp
kANt4E16jG6hb/okmK28/3QN5zL8z1OdcCbqD0J9Wj9NNf8vl2mDAA9bvHCmSoWS
mcqMLXNdHrSNRWXGriD2eC4QTxL9srZEV6vuLc72Oft4btWVUVpr3MiWlYzuheMu
evBchj2y1USR2/OHAwCIQfio40KMwbbGMluDUEeGZyL30Imwow/CymfYNe54CYxe
S95AU8vNiRd7pNCHkK3vxw5eh7OtoVkdUVR/tPowsW5xHVkARVeGD1nB0GJVbZ2o
4bwMuj+kUdsczdWJYM4ENFBjx0v4KTrvTa/qa38nE5tINjM8UAY5o6XB6P3fl4/t
autzXRLe0+XEbYd1J/ysYrkufuLKDvSlyP4mjfdgXIKw3oHETWgTChP9kR7e7/KH
WjQg5NYfA6pwXmpFUO/21DezWrxph6dFm+/H7iySleo7c+vhmaaRLYS7T5hGXVlr
EbFECaHQzDdb53wbCQmnPC8HRm7wAT+m78MPSQPKY3fMvpzUjzMVbB7iK5h3wb9a
aP61gV2/Ji1wWRS+NbhHBssK6XVBl67S3KN2gJDSNMLca6VHdkElmw/Q3jeTmKqc
8vp8aXuU7TYCHPuumrOzm5HX9iYFQG0s6P4ltWND8bbaItsQSekwKlWm7eD5a/xx
JfqoFceFnXLbc89FhfTTevcwR0CKEZMm52AsZ0NP2XMGBq5dZyrsmSiaAfwph0Xo
BbvUIbwrpWhCLodZ1nljc2cyEXFerr6S8/68vlcTvKtGIeJh8PZKamk0RIZGaXS2
6FZLVbBA5rRfLznTzR95EKkJIbsT7u7x6FxeVI7344DBYADysAYr5av+fEKW2osF
vXgT3tuUtj+DY3HKxdfwQsGr0jmg0MbLiuhR/XbJlaBnCLc/ncuRido2rXpjuU4Q
eorRwEL2SkBZ/1ni+yxpneuVhXMjPsgzDgeMHLy6OPJRe5HR6J7+4CS7Kr6lMMKi
/yfmpqSzzTyr5QSWRBM5PMh0w4tn5dHUeHPHsGwEMtHPAOcOZ4gzYXaaKAExaqDM
99VPyRW0DnTywq5WVj6qR0vU6dkOpe7mE3VpWiEDhhdRIuwZF8TBxoTuvpzr/rRG
LBsnBZRenarG1IMqeFMwXrVmshMK0uJDrWpvSBx5ml7eXjRnCMS0IZ+m349+QKU9
zp7n701TCjHomP96/iRSd2U8xRiomN+UzZNCrU2RJ6WE1KvBSHdrSfxXiR35R4Pg
WSxuqrIQi2SF+y4UbQETEYGJLd1GMndb13ve6nFrQbmd3WYXVusaWSmJtzu/BaP6
+fyE/nBXo5qXwxOTz75gnag741tQYN8EjpPe6u1vHhnqji+SVh8Cr6VFdGzOtTfC
KTUxtJ0e7JCigbFE9cQTS1/KMR/59eTn3nomSU18DNjgmNxSW9eu7++O8T+gAbOD
xmHU3V/lmEKBVbqQsVaDSZeBun2aVm1eAeOl43fLhjVqVFowRFOZCxvLZkrhXLkA
ZL6GKdiBb7NzdYlMHhYlAoSrmOhV20K3h0vyhKf0UvPm5YPQggRH4jRc3657yiIO
XsHNEN2IUtPvni5eRb/7OwKqvudJnpQo8Q0GMEuMS2HdEAEVyA0QEq1VFCPgjT9r
+54XryoMuzbFraaA1XuLiRB/VAxyh5oYXyrGA4NwYV1nXMbQoKvQSKc51tEcLxcK
73LcrpL9s7L2aS5hRMmeagGljPCDME3geIgaepOzUZFHzRpRTipKDQCQEPyPWwwh
HhXGLNndfWxyOvjfRyM6WdW+V66yOimfWC9GUJKXgG7bumdoFPhFIfN+VJIowYwk
HrtfPbpjkwfyGUqcLsDdQyslr39whErLbqI2mAvL3pe5RrAt2MqKnO9jvXqB2A45
wiYokrbewep9973Ah40cBN2ui504mqRYQ/P8JOrCcqlXJVFeD2mDZrJKBZnJ8NJ0
7FyMYwGHBwA7xJDhXMsa0Ajoy/ecK16Y4aDqroiBsZB9NPN4UPQ2gB8IMU707813
bMXQGXjjbm7me5+qI7366OSosEkg68gFAaPhS6T7gs/B6DKZIl/JfsdBQKCNjnUc
q8TFxjb1qudmmD0Vw9QgD2LtSvODwP9seU48iob1XIyW+OPWexN84RwSjjru0drI
j1GW976IxGVVVSvuzXXOfgxKuL6yFpVcADuXDyxNLGq7XNw6Kq60mdbvEAaTDvkA
zZoG1nhng5+3UZ7xatur1Vo3GfF/mg/5p5XaiZwnr2oWL8SC1Lr+mDY3hwQwlXEZ
9NlBk3oAxhi757sncYB8qR0+8rcZFtKI+8gTzxeCDoSQQR52a2d5tDE+tvMf9IYs
vu8cEbtLp2BS9Hhigf7tkePgYKVLzA1nZk+XfA4WFEbYazVQCgO2HXI8I3F/U5HR
pFoc4i55BlxPO73HjzJdrH0JrQCklAr54/Bnj1pbVVOecUFfpYwOzxVLk5zRYnc+
QgIrgTLUphce/gBg0a74cDQETSyH+dVQ6+0U7o5X0q35A/bUfvv5IRO+/cB0M6qq
dqegErDAjdTrBBALLGoPLV1UQVNUhCJL8RYSwgmnTXpcypPADWyoTX44T7Aydrku
xr9ehR901nAM+gAgIVT8yF1/3b3bXSC1TsemQsUOAa3YhLCC5icZ2lX3G9fkcKAH
A66lCSAgCc7STB56pb6CG0KbCF9n8iBGnmg0pDzjDfMkDvGYB/sbJJ66aK5eh8QT
+P+J1WNJ89bOybBT8IPJYDJSsQDyKxk8wRXCrU5S4GY5INkDIB3ywyrlDzoJuDd/
QUnLIIhd93UX83UyIV94o3lWM6pe45gMnpe27MQY2f38Wt8MmxrYxGRrlxRuKPvh
iCYFhPVcLRko6pNWrZcaFcFB/J82URZPhViK2qHwWV28bj4XL6TVPSfJkLUyKZJJ
pmbO1vDkJWQpUbOkt54dYPY4W7kRc6/Gxs+RrGe6TBx450Ayhn12sDHfzN/G9CNR
hUT3BfWu455qZaRtRIM2m9FVSlCq6qC1xRA3RCX5DbMNXxkcRKxERaqeiQwOk2l3
HXZ/+lF38p9CcYzZECamgJqWUpphSx1k9tPEgPEERWRrHipbuAgMtS5uRI84qFBQ
2S+TFpszJVngq6KxNYjSVwJjr4ASals/NW7h5IDZX4HFBA7l4j7ZqmgS7oY0XeUx
i0YViTT+cz1iSB5+pCK+W24rry3D6FcMHiCxHdbHySgD0GYsJ4dWV3y3az2RkgD7
o8X9ed+8X34uO2TymNQ4DfdEmrbaFGFU5i3ft+h9QlGjKBq8vjUlasCX0YphMyVz
+EFWWTevL6s7BZp/ICVChAjg6w++cuTCxKBEpLqKrXl1rk1vQp/6cSdTFOvbD9/h
XmSlMuZyvnwFljnAe2pGn8ykOIMvWxvBZzlWog/9cMfd/EzyMfNPLEIkb0QjRo6G
SbUmQWND8TTZjqliqPOopQ7bMTwaUhPqrHdIpgoTj2x/FYOdL2pq1f3D+zCJucfg
J3wOxKjdGcXQrdsrWlNr827lvUWJIYrSgXpIy3tm7MZ84WwqQACFt4dkDDOg1pT4
RObfBumZO5RQFsfDutPHICMyJZejLrxM5DzmQl60XRcsv7k/KKG8QLTygDBhJceX
EMaDy557qg/HrERJ4tUr3XTzH9RzyjmHIjboPDDoCw3I2PjbKeYIC4S6BVa8iP60
jGLOBOKOQDfdV+jxH9FSfUI9TPSj0oY79Jsnz0r+F602FpKY7e3LgD9JKD4R4VsA
UAvUAm34r2UzJjyHXFJfCil8gL+bcvU4gLYmR+Z1e4qrb6jBpAEMikFd7f0x0pif
wJpS6Y7wFIfCpSAyu8Qgcli+/h0hUIy4Pu3XsMUZA/Dq8vNURIRwxi7VV1/zlyjO
CgiYZNybgdu1v0HOHJuTTYLTAxhYbvz+U6elUKUgRsvozqiFEwWdwwxA5CAjNegk
XWobPKuGbKGHUDAvU1h+FuNyYB4GQjJ1/eqeBQoUIXVE0F0vYgCHhuccmBgO5nND
9CtuF6i9Mi3IbGpDHecHcvWh11qHkCEwdMXmqOeZdhshDrcRSzXBXHu7At2jQL0d
t+M0J1IogvW6+bqgcGUECOGvh3aw0Y53w+LQX5jIecrJN67J+N1jt5nY6RDqUq0v
TY9/M27QmM5E8qXuAlqSzjYsAOOb7+OGcr8Hd11cQwLY0COGEJ1ILf2jbO3BOZoV
8X04SkiCo/5rck+qgQUetjkDcBPVVuDOOZ8/58bb3O8hK3HojfyXYDyrUPAErqIK
M//Jci85j4bsXlNdbRjIwKkxgb+XidCVp4cDMLDusWQ6ioo4e525tpwmdN59nVju
JeGMxu2lEgnUdHaxrtk+gwAgoLQ177JFGRxEDfF4nYpZHBcrIhL9spTpK1VEONhz
BPeCqzSjHOqlCf3ZbWw9nrmzVj/ef+zaNu595r8z2vlzLAql6HmiSKN0FnHwrfpa
8kxH1rdTASGDFqqX6GhfODF7BAYCpUBty48mzTihQvK3qK2gByoMtL5ECNnZ8uSN
VJjDVzFBTVnywgC9t7cxmfPZNn9Y6DlSPT8OPtx6udt93XEpwRJrkq4ZaTSarCBS
w9uKXu/5yMuR+ehSJMQXaCKXWQWeKVYXDB6KSaF6kGioNymZHlASytfPqWv4FDWk
JqxwOTZqAC1unj3I3/ZbVYpWsmL7cuPLJGtTbeG+KCQ4O4twBshHdzq2CkMmkVz7
NVl97weVlB/c1+5kjfxJg/NMcwee+alLesxkGuoIDJNouhiHlhmItP233sc0yL5T
jyMWKQVd3Fm8DplyjF8U5gtHysB/KNmeRRLuS2M0N9EyfHtNoed5wJf2BREHh44z
3YhWicqjOqntXiTFyV5zZzEQbBn4TXDvNQe6Mt+5tFtk8E7AcGqbq5+aV17FV4GL
OGc+IhdNHeOrNAq39t2RnZtb2oJVXQPcb7V1x+p1P548CPjpYd8KUYFWaHwAhjgN
jmenG44TtvZTbKaVR5djFwgrCYeZ6mrBqKqc4xPbIxv1Gk6tdDqBMhGJxPn1+zhF
ujhNGPVonbtpu6KA3Ggn7ZqTZ8b5tts4eRo99i4+slFAiRRmejPc7OyhzlmZoa90
bHa1FaflMbI5PnVVJdMruzPGBKUXchnN3dEeJlO4AmCPNp1TyPdcN+Pn1sJG12zM
nk8wSoaMBnKz6TVQGJZNfGk2YmRkqJ7jvUhest4nKHARxC5SufmjpERbSza0MjqJ
WwORhnc/UQavQ9VYjKyti1GnM1xw5f2VPULp3c8ewc4s9YVx0esuCLneRsr41Q1B
boxpxE43AqgtmUwc54calVBoUOXppVWcNif3GFSfMvQF33SnG/6s+T3CCErfqL3a
XTnhDNQ/9/tAhNhmr6uF5IgRYEcyoLfe9Eb6F9/R4Sgf3v7Jj/Gsi6Ta47afjjmQ
RlYrLs1uFpY2rVBrrVwCGtKfjdcI1/g8jc50Xt6oYQJN+sjK08mQjx8z430x128P
/dpuomx+jg+adKOAVqk9XfKqp+rOMnnoaSyM4YHEjMEeg336tSoUT3T/agbVCkNj
n/IM/ZS7xs7d4rbSSvpSLsTpEF5h7Bom1zeLp4in4NesWiupBe6JYMSEc0l6DYuW
sFYjbPrwsFLvAad/kUHCxODipEBc7RUciSu5udHnvYdBIqe/dmaSd6EnJINkb2U6
aOmZSvKVHV0Q5BwWRlsoxmBOlr5fKw8Y8BJyRJaNtpSsyPRhGzjXeSmQcKljB7+a
iaf7As9+GJSHXW1RYZvhnVpheELGYsdCdNZ3lq5YmMXw9lsAS+pMcmcEFTpT9a3k
v5ZpGJ4Gmwuom4Z3BG2+TuQ4xM6wyEqhw5QDbU5X8LiHh+YthrMIwAiNBzd6gMmX
Js3fQnzY0acYTA4ZrHpOdmriwk62RuOEnFQ4TWVgurBOqjCjgR213JRZ7EyXLPNi
exB+aiICNsX0ySjAkxISebz1pyOAohnI3XC0DCRmRUiDIHSxfTuMA+UheNhNts0+
/H3S+xTdNRNtZNeukXqXF26EpYpiguPw9XDQSrJHcpB0p1CeKCsJW28p6J+rLUhB
E3NpUXbvuneZKca+4CnH0eWIKnB5bGH9wwQjmIrgxyVe+e8KFT+Ixlop9w3plb7I
sEcSY3E5T09hIBsF5NfBJbbHc7q5hmqsTZGnBFYSc8ooErtkp1b2CDB2L8CO8v+o
x3ZoZd2DJBUQnAvHg01n2NOYoMdj4aTnl6REkPq6dXTG7DimzsUcSasgSE2goWmz
RuAIfqODh4pIBdgOaMyzMBEWwhq+VP0lRhQigrh69M41402rk0Ie6rWeVAoqHRXb
QF2IpTbeXg77qOjm4e5PKHYRNxwUrCBiNLVD4C6pdH5VSTuHWRLADtKZMl6G5TLt
phON7iOzSri4X33tXew2i/gpAbs+nrOq+fSLT/vycPuT4Zt8RyIgDTJUIe5fELil
dZDV7f40Qn33oZPBi3l/taYuua9bokm/tXCEBUpY87PvGdlYGUwFaGKWuMEIGzcz
euld0F7g97iiwj49sn1W5O5LVha72vig+kk7mP2c/e2aF2blcqepw5Aap7hGJv/Y
oqH/zhR81rEOGbfv8eF74Mn+0khAlFEvCUxQjzOZWZh42i+sf0IqLd9Z8G+SXJXV
EZhXzt1ipXhLzirbh+Pf74+Nv8n3tVp7qDLOuoLxbm9qjCiqgAqA1u5sqPuxocRe
S3jCGKGEtvMuUCeZA9vGt1c1ySEIlO31HdFAFsjKCpNlxmGRHxiJ36q/ydwFV10i
PTTWM9OlpjYZOFPfwTT3Ug23b6WUt5hOmWY5AzrQ+kg3h6Hq/5i801D73rCamSiS
HHLOl8hXLCxdUzKMxRVyoZGTL1PYnihG5pIN7M9uo+VdZnb+VsCAQaRp9C6RzJCL
DWibceZ1Ib/zdESmwFpmcUsO9nMVNfn4yEAV4TsgqoQeTebBP+jScVYwLq3sfAJD
lTzIpbX+AYnCzfnRzuRJI13ASFE7CnqwoRwlpHo+JJM7R/VYMl5zak5WCA5F5yuA
1jMwLP8XnkP+Uzg8x1WavJf+gfKZtmi16RQI0x8x3LfqzDfZucFwEnNxYw7HRENJ
rv0KVo9eEAKEMAIrXtzbr6JqHv/W3/hl9KtEbcEKdZ2Quxprnf/xO3rFUbfp5KyO
X7ZpoaxdEkPuQHavrimG2mb6B3mc0CNlfP4a5nkqjqSUa2b8+YyGYd6I5l+2ji9/
LSDHX8huk1O4zoATJx9q4ttHvMXbLzfs0ch/gymuP7au+gZ+GVAzn8uhs9ec1Q7a
NYFwztGyaHQN+zCUhX+2PivT66P7EwFWRYy00zoU+XabBcQ8tE70hVWKHP6GI+6v
iWLumjbsIrPRzcMCXOuy6BcbmepEnM9qAv8VkuqQWaDSWNit8qneI06VVvI1yyuy
6kthY5+7TnanuRTfjd0bIZfgX5BwN5ybhOzNmYy0Hq0v+t46jNWpQ58D3axj6ERZ
012j6vLGbVb/MS2QAzq8o8Ja5U131Ltj88SAk6NCGSn814HpokBqI64Ym3qa7ROO
S5+bUC4NUErQQpd1nC0+rjZLeES0vdA/lZt5G5+TxBSCpFdZtY90q6hA22EyptW3
9dUwl/68kGwe8GKIWCN4NabvNBkXtmaKH4iRMwHHsJEyS19ltvQ58iTAKyivYd0X
MOSkCBoJfry2aZeWU1p9WaclefXth242JNJHUI1mYdF5pgJy176x4M0bAHsQp1JR
G9YZJCrBiYwYt01nS29S5CYvAGlds1cHXiS1nVxbI/YKMTDwJsKLrelNxxfdvisv
cce5KOXQk1sGW97PxrL7I5rp4r2i7kNeblz563QrpWaSb5ccuaM+ANeZQklSOKxx
JXYCaWDripg4S9vNkymrW6C2q6puWxW4ZCuogeQtNssoaCqctPv+Evcq41lEvuov
MpkZiIFM0jWiFZpawAFmAP80iwZHtp9swzD6VYIYMOhf3tnnRjr93qqnhjhWsvn0
M43kjze46VB5O0o8s6a9j1j4TvYdCl4X/aMQkr+vwZYAuwCdNxiWdMFXZ9XkxcoR
IsVPU25+cYA8QI1HpNt9dgcsK7hQOJzIm6IWYYDNTn+YWsQyJAT4hl3KObGedQik
tGEhMRPufwmpqooedCPSjXdkAOlDWEF/XMAHNya7VSbwp6xiXgfvu1UyNRqtZmcw
42OGoPiTX0Y302JYzRJskv18VYTDSBG2n/NomYMK+II8QYuK4OUYfo+JYA9D8yyf
GqGRO037RsH31ZVFhsNbL/Kg8uncLOEMN9Jqhv5HQ4RJq1+X3NKfPcJGEqQk0i9n
ZNk6q07N+qUzmMDpI6quGM9XV7gTd8UATMLXEqhnELJAz6HgTX+Dd99Iqn5xR8cS
yuO3BgElVUty/gKL6j19qwZTm2EsRuRejc/uCrCIxeqUDAKglpgvdv7bIUPXLmWS
pgoDW1nQkKohzDTVwNSMXsVkeiXBaNKNHPWd+NkL0rwOP4vyt1gSV8PM4l+SJakQ
bI2zSxWaqaoNRdDcpxi7T5QEmJnlmvDMWURudIWJEDRYlbs/PzAqI/3XPYEojOWL
XCVT9Ga2ZUj2D7mxyBOLw9vN7/dmvfDs4Z1Q6bf4KtRNV9b7l3ABzo6QaOfoxwEi
ZYy25vrkQc0DRFOMCT+nMtUcByhHQIN0UP+TkoHu8pNg+Qse+DAMNk8hAUzVqUvC
E7hS0UjLWWYr9ZHyuvkCCs4x1spXmiz9OmUC3/icv1RUlDLr3Zj75OM0ZsX2wIpB
T2DyXjAhiQkiJnaljLwEB9HP8onO4NhpPscQ9GzIm+nXynlOf7oPjuJU4Cb9x4Os
osqAYFywnBYVgRfYogMzWN8Ia60PEiB/d5PLOyOc67L9us/EavVcZCnWEkhDl8en
5PlK6bcD3sgREaY6y5ZlsrMUTCsjcz5syi+jNQSiTzepEebZyiG9Cdl0h9UM+FT0
UdeKrM3DRl8dX3RL5ZD0Fa7MkmBSSQaxg7aHZgGfkcdwkoyEfe1XfvI69B98DJCX
vXT8YcdXisQiqRLoe0Grl2BEYTE9nFHRQIJ3LJjnXUZNolYmNDhUYv2wcg5js8CC
D6rwaZacaE08aSVsuC2zTRd+ojDRA/H1FoxPPOY7vGfZCD4Dag/dHahDzwo0oFx0
t6t+SCnMdXv5iwL3kbR3xrHHDUASHL078l46MTYAW71Ez4vNzvr+fS0uJrxqxE5y
XQ7w/4v4llVXMwgHB/qlZreK0tPv4/jNgzgJFGfnukz5G3aOFYqaUJUET9e8ECDa
nTAO4OI/SdRADD62Mg8rsOI9neN0IiGS7smRyhfF4siQrBLcNX8HuEZ8vqSZ2dXf
CQ2/s5vSFIy+2xb7hxHeeiUaRxwHhk1OaUHHcwougSXc8gtvGMlUSm99evQToFfa
A++WfzNeiVLB3zeILdj5Ovm5lGO5edfhrCa4ZbqYRKyEOHXJtrFux91JxJ1THUgp
Fk8sz+ss7d+bYYnpxMEEO3oSBz2cNpKigIOpIDdzB+qwXMxA04Vih/HvjIrw5gCl
VcCoMvVUvw7IrVfC7dBNyYYJ1ng+1WMVLge4Ty00qV7K8eHpFtKZU+Ctj6YjgmX7
U3+q48SWw5d9uBoArEFV5htQhQ3IB2BI9y7coHl6dkzlfM5p7fE0p478hWT4eoCW
Y+PknywSCmQDT1BYOU0+BZ9ODlvkwg7CjcEyEd7d5f2YoHhZ6YLmwNuxVt3EHEen
FyxV1wkBVjIIUUdoGvs9PYhfc9qZxPTUMfCD273aJ+idOBjmplftsRM+e7Ix300h
h5UVjANVBdNrXk8r88cJw1vd5i59pWO1myicg8fsSO02XDIKJLYg8bWdeKGHQW73
qAj26cbJ2dbsX1zoWwgTpOT56+TT7ndCFedFSde7uFIEA0An796gahbhW86JdwES
bIb77AZXppz/xNAHbMARq/8CjgcRDJ48LJ7/t/iU0lA4Jtsmpwl7h/6fwUAsdQop
iCihCTFl82lESsL1jxaVvCNUETrLPHQQUj+jGUcRP/a2SIjcmlIbrTUlMFKgjmxJ
ZLFgqZIdFqlB9ih4eXN9FcgBUX4H4ezBBC7j2L/KDXYDT22UDtQYuPJWBQvcF7T7
kq1MVJyeCkgbBosNkx4NmzfxgjYSICT/tDJI+X722nRZz3q1pPy1FnjjMTri1WiW
LUh458vMjnxmISrWBoWVBfRlO31f21LQ5AOsbmYalAKHUMzsOOyTTblSgzw7xuaM
B3EB20+Q+rP8Dj7YUjUyi4weTgGswNMYYsmX69L3D1dtp+gTWUidJY1eJWFmpQiJ
pvCbg2mTdVeid+VLCMsTE1iDT8/Ne96/WaaJLqAuCCqUBCQMKQrFowPMwILdKEGl
a7GraYIXgc9mzXA4DktmE8R7YDKkpF2t1jN6UosfqkXRojeRlFWQwVvHFtAzo3mO
iwtGXdZst9PO3sSrqFbmilLkYZycV391ROszLx109CZBY9pFd44j5bStdTEGyClE
yvD6igTBnsjK5zX/Cu3HSa3MjmamZOVjg5nY3CCuI84iLd7PIyNKpwIPVkeKe6pL
XLiQCnkin2lxC2/1lHusmJk53a9QgO+67mHmPPzm2DLeIZriEyMTLZ0GUh7At9F3
9o9CIDe7v0l86ZrvgkA+u+/w3PfC8GpudtS4mjvtNFhS+t3qzXkhLuxzY7k4ZEG7
13xmmwGNs3B6rTXmweJN9MlfvSCHiPUx1piy6V6sIrc5L5iyDWzlvuNjFGYdB+Po
k8DODo9MKXcMEkY3FShKmq/0EO1G59KI0WzOWK+thukbT3DhEyl/xxXxp1dU5Pdd
gD3ad8X6uekbP5KooIT/JaUQgDc3kUMK82u8lafoSALpeqoe/4PvYreIwvvqjlyq
p+1WEUMhVxH1ceuE/Osg74i9wYR4CFH6XmzNQ/pI27/xe6hsi1xhEAqtJgq/8HBk
Jj8Kbnv5ZnxByg5vQyNxkW529DPlwQY1NLxKQARGj4qj77fgo+k2wD+zHvBHDhcm
zcMwkNHTXf+fESvqfwkrXRHQFcpm6tKoFUOehohuUYjOgrEDZotT20E3q8eR4/bj
E62LEjFZyPx0Nw+SlWnjxzsjNNoMFhdH0LNwjDiYySCKigqsAoFDg+MHOpntYLMW
aKqFD1MdFaORWHrBDzLcyRMm7WR2mPwMofRTKo+hZEzfXqXkHVff+Z4L14rNNnrZ
48HojQSe0A1uBd1ulmJBPVxuMKW/OetIWndNJd5e+iLwEjOfdQNDwQySXNq8htYc
Em7bVMjzVeMaImuuGGvZ/MurXUXK0qsXbPnShA2oQBMlCVlAwN4f8u7dOVhBgjuz
WbYz4D9JDKvJQlTS1vS0QW4aUAsVGmT0FqppyoeUSC1mc82gOVZRQC+NHHLDuBQu
oyxIb1A+4Rp9V35ogPhdjg7/VrSShHK1xnToH3TiUR4ZHbt9Th/pIZ4/wdbdTVH7
pcodvgT81G7LrX1Wtlks7enH/MCQ+QvMpUtYYE3KeGOyTNRybvz699TRMTVnTNFR
QGIKUX5No6xZfGeBD7b4LMcEo880INwRzLjIn5Rqw5raM5lOqrUFTg4zH1qhVce3
wIW5+ORotf3630hzKsylsh0k/OrMG1IVD3i8bFMeHpLtqhXKgfgWxPae9WaLzZXM
houX94VrUtsZKVFOGwQOtJrpt9WILGZYzcrcJADEcg+Bru8r/+uy2JvwAy0A7dgi
cx5hdM1CHTi09pd3LAKG2wHIWA1B5IyTf6AFO3gVaYRbzWPQ3iSRuPtrujVjnUp7
bKJUjmFMPDJo8NPzQwbifZgVVexVfPoOKY+qDR7UsHJzaGRxzjqY0RY1tDU+Axj8
lxniiCVkGNpX+bzOkO8/9OCQOqrAeMimRUyXYHzCMbf00Q4xAILrZ2vdOrI//hyZ
y50sOZH7pxNA+TM+x4YS2V/vZJRQxgEwl+GKMqVa0q2/qODLmOjVggHfWBXUj97n
AMCZMtFrKTdHd9FaFt56DrbYi6AKmF7VIsn9LtmReEFtERnRzmqkfjN8p50LvTYX
WQdpM/QpZqUsqqg1LevpuVKJ2ThEoV+eROhQ3+pmO62lEE2ZiO9HEHn+2xSCscg4
m7RoxkZY6G2EhRjrEdPLFelyPiajb83crqYNPmTEkXa3yl2VM39TEliDfWrdA9Tt
guyBaQ1SkObDofClIi9ARvOMJphZ6bYt0QourH5h2BbPP0B/T1qczBH2g61FWpp9
t7mdgfNeFYfpYGqzDt+VADv3VK3PDd0RX4lHTRtRDTziQtNBILf2Qkyvgb/CkTK6
9jUgXJ1sipsaY3Z5aLumC/e0bf/FS8uWVJdfuEOwXGnBI//i0M8nd2sRRzu0yLi+
4VUnzjZrlD/3rZYNVIAc3DUVcmWLjOLxGmT2oKcpARautWmCRjhBBRzzBEGooxg+
/30+aLtkAFBvBjhSmm9kLBGKztE1TH9/iF8xHXqNERYO8//hgyH8j/oKXqGGdYRS
yCz0tVp5byTwEmvR/s4778w0SbH2OJ01Aue9vj+WJl4Qu97jtT1QOUZ6UU9iAt7N
Nw0n3Uwq0STO8rKoSgJMpudNF8plW9ikBXTMGone5wmY6dLt3DAsUA5ZxQ2n5Gi1
wMw8iNmckpFL4GBt3RcAkeacKqTD06OlYAguS1jbIxJsjAfBvLI3TYWJrl+5YPTa
e/bylUMUJZBzAviZG1fLY7/nU1ClccZbQVlLlhK3gFU7+dyhOrdQXFZd7ZHl+GXA
aSLIX0v3L4H4cFXHOsuKjifnvgDu9Rj/H/Klry/QCvmDRrCs3Io9KJl7zKCttrlp
ZzJyM8kwAG3OBeysUJwmFTf//TughUbnD0EIt5bGvfvBJ+K4i5CHb01wirFVSiVp
V524jqf+FjsFQ+yGkYH3czBEfwPDolH27LzdXTF0NQAfMVVKGwNdl/7nuoLWtzX+
rG09eWSQI9Uabitncvb6pggXZIuj6dIZsdoQfM9AnKTONWJOw35DxgfUkKAYQP3x
VQ+R2huI5seV+DscEoaNULuAWWBYuHBAMKvGWHJ6tNkqzyTgrkK+dl5r+OBmmoyc
OTrFCV6NdTRDOc/Gd+mnaKlPHi70HSRmyMv55UCwcAIhzrTT+hAyGLDjbjp/3o9q
l/QpFzkd19n4Wu4lM2h6gcRd7DJjBY7wyedQyYQr2pA3re7LMCFAp/Q6p9UefG70
6RFI1GCepeBGe5okv/xk7lqX0pfv0UqHCUHnkvkNU3bVveYyaK1X1jdy+Oq3qiJx
yf096MzTNus5nMRYfQWgCw5vHDZktWesp5qk6N7s3rz6HuvLo25ehWl1bXHEPGcm
9Uk9VsdHs5LPzXEv5zkA9yjs2BnnJ75UoDrij58sw3G3AOCzYXgj94JziJUVYk09
W6oE32GFiMZeID0C/ni36rve0d0okfFcDpeMWy/DwhyM3wOs9j5znVEH68JmOhpH
su7+p8bDd50I5KlSdCIbJ/ddiXq3Gnt2Fzmv9qGFdr3bqv3UbiehWPIO9DJK5g24
kPM4tw0fn7jqREx74Iqeja5kwzjMiB+2s6CMMrPP870heY4SNo4jzXpfINEsjzs/
X/bpbyqRhT7xYe0XH8rSO8p+9Clil3yYSfO+najKogxqy7bYRSzG0MS79dRKeCfl
oE/MywBRAQld07FaJ8iX+XPx8iSpfPBfMIdrlInBMLZTMOUD7dlAW1lpL+2uwwTF
fHA/GxtG/BuAI3EsHkbm9jqf3XzUbKmMya9sjfxYoqimUjXBP/+4z6gsSZmzjIat
1qDUaTGB+Fo4yOaS9WzDFgDXoMvcc7IUjez79cLk6V14aLNIhM1E3AYXfPzRQOv2
3PH5QZREQLW1+TzZ/vSHlVSWr5sLf2vnQ6xCNQHMIcIaeKPOaui0UZlXDY72Tzvj
exz07wdCzPY9orClHXNuoyk8NmYS4+UfkpQdzP6XWk0UmzXdTpPQXp7tMpeo54UJ
rDOR8YH0mMKlU0GiwMAQrgxuemH5yJ8ePZwbeK840bgbDzKue+Tgzv4mtNtU5PHe
fw1oerkTjQLRK3nB6LUFfeZ6Y2HQD23bBYDMTp3CaxgklNpZKtAHvFE+avCTwTcc
QwuEvS1Ot6MVWQx3lfoZJulhDG5BfemY8/RfoBjANlazp2GnRPyxGG1B+wqCtwQ+
V7bejOlyKw1FjIYM49SHnw69jP0YS0n1Uns9PQ/B8GPQVh312bFvOq34T485kppS
nYtR4UJclefuYqik17L+kPq51b3ULY+hR4yxcVtp1K/vXj2tvIBR2Bhg/xqyANzd
gBaOiPnvqIGjm0cUx0QfBbgM5gIST3XWJNj/0jfrrbUC+a7/EK99YXgweN9i3TsZ
Z04QRX709sZm0yexdGodRq4i94984oWl7Af+NBQm8i3Q6GoxUtCqEH9UGyuSB+qQ
75VzMH2fXrYgmSBT+TDYSvNd8J0at4/cMwrCd4P7vvO5dfZRY+Y015ITTVZ3Wq7h
xIqbVCdQmjcCEGlyfKnD3xlgMHqzGVOVdM8oXcI5aKSx7vfK08ZYqVEUajjUpnGA
xbnF1Zk2d22u3IFGWFb/ePowyAxvV0mrhhjZ+TXBy+sAmpmrp1BmA5otOAaVwCay
sLzO/TNBLvprEmU0FmDgFgYWSVGW/aiWPMJuDnsRfOiTx+yi29Sh7wWn9/y7Th7V
Af4ajTiVyMSSS93qjhEVdEo9+4I21oiLSaHe8cDtFXpSvaPzaRbWzWVgteVC4u7C
ov64ZQWyJBTW/AhkkPnz6ax3nD32sPDKJ/jnnajUR0P6p8ejj1czWslWxOk29c00
u+tKq/fgpYOWL//eShKAdswjj8IS/gcr1R/7kWyIo++mqmPlJPJixFNOKZcbb537
54rmA/LMpiJ6kV2+g9iIcnApZfvPhhXm4/dp4C+tBYYr3YKBMYlAk7PtTKtvlDCu
b/ROYghfesakqYGUrKXZqAzwidf+Q58TuZH1T+rssAqrWOUdZB5S/fQMFRttbIwS
Houdyercvz9hgTMVDuz8xA4pU4BcKZ7PI8yCCsl+GweURgIoUX1wQ4wCnDLcbJMv
127wpU6zB9R2BWLEBjbAFKa8f2PZ7A2ThiGWmTfUFcjw5VZkroaDEtAaaZzX8T8V
aXYgChjLrjjOcG6yaihiDBPj5xy1zf0AKX3UM0SwVKSinp9WVgX7xF+nyUxDRSrF
lvy1MGb3L5hcpedjdIgpFZPoTkiJy8+HYpRO6RD79kY29WX0XxtRPASP8rMSbD+P
dePkt0HHpmdkpXw8NrR3pj37iUvCJxCgd9kdo/6JIZyCLn0KGjjbKVE+iGpVJFhb
nJqXO5+SHCYtXFkOimPEkOUcSE7pW6zJzIdm+nVwq2dssTOSHlSx1le18VOrBtOs
YhSKeJ0AI/fuTBmipbKgQIMZ8xy66R5/55KkZw0ClTnd3z7bvqCzWEFvzRxB79Ea
YQ+nb+w/JGkLsCJE5V/k/YZ9FI+VYV24Yn8WCRhj/JBQVbUVw6rI4CsuUlE+fWML
1HJDguRGgEylyVHd/SYWYX11PYxtRkSZcg3+FQ3u7mB/zen5JdHosEg3/t1W2q/y
IvRcNDg0pifNwPd5dzp0Ytu5uowTs+hOMusEjfmcVSkHynHkXwZYoFC7uIhWjJAN
HBdGcK73gdZNWBM3sFjI1RzCqquZmkFDn8YU1v0luzrDBlWoOnOb7SknW2bhxans
PeJc0Jmr4BWs1zVfhyy4t3+sveJ7ZhxT3cpNm6MwG5nQB691NQy+qkxB9Nee1FN0
T48FRtR5X5jlxo2EObXmjGir46+VzOy7n+lOHz1ShoMQtALQjcYyFEpYqH5pbBnv
fBdyy7c6Lsxo8krxGvVlXyWFejVQ/zqMCFfrOc0fVFA/TfVBTPK9vvWdIJHki32r
xRyfXCo2EvcczN8RaQho02vyoVIGv59WuDq66+cJd5ibeWzrpZD2vvMcnDQbj5ER
O8ww+zM/mGSsmJFpII2lN4bZ6PFKCuVD1fhmoVeAjWngnAjdz5Z3wU864e2ctqTE
FLKKQx8UeVgkT8//9Qel40mtjsjt+PZSFVjQNig96Pp9fR9Qj5UcANR/tOb07OGV
ZMP422rU0qi+BeHo0CDTkEBCNEdJR8tR8NsavQi5ndgpJW05boa0+++JSK/XOZ+Z
9mt2fIvkfaSA/9uAV71MYCL+zqxyX0Q6lQ28k2Kjqo6PLNN/vT8jWbPg4MfLax5g
9OHbl1SnHt5ITU9NIEw+oodz49bMbKY1Zm593OWTQcaP3+nmqkQjrAgPnpNJfVUH
LK7ALZ+NMtG5tMNTxpfWVFnukX2josoT5RsuNhLktevWYpKLQYAa+jqLN2JelUYL
IgAJhtujl0UBO2rzj4GB9PWj4v3eE9s+rYPcMkoQJq5zltYfo0nKdYXmt3IOeOW4
Bx3HgcTfnlz66xIAx2wOoekm0F7BXI2cieLz7u4+xhGUrw40BP1IbZ7P9tha1uiJ
Wd8LO3kCDTca55kJBfJG8oTr84h7ThnG8ilDElLtiXcjEebr32fVAw1VcDJZvAPD
a7JA6xBf3veLzl4W0kARviEd123K0GezoC+tjo5EotEBbjzSZPi0IZJ4ij4OWX8L
HNnW62SPf3y/12vpVFJhUT9B19oJs47iGjKGZw4PYYmz1OdWyxLUhxeWcf9N6GLg
CnJhXpeZQhnSmLGVNkrd4L15IjB4kPldWwiGyi1/PdPIie4zMv+Y4K468o1ZuJWj
oAryjsBV91dZI4DNl+fSNz2bHRkELq7z4eZw08QFxIAcaUqE2XaOTez3xOgEFpyE
0uqD0xChqQpYDAt1aQhvCg5jkH71I59m3wLNyn2rKjUxnAy6BRW1oH8HIHIrzd9p
gR4o2SpUV/bnE72OSurGZnVeXeSvFq28m2jdETF8L+Ib3HjHbN9XCOO7uhX1dyMM
M8LHn/vit4TwDlrdDe3rGcekR657FWQcQqXnBbXPypkXEtSzbAsVSDirr+xfB0Uc
j8f9hQY8tY8lWaJLqA02JJJ/19UWZmYtHsVskBYWAILt/O3W8WkNHS+kt5d2ZlLu
PuI03tm8nCaBAEoX/xAupD1q7MlhSHefsaKaecUmhIDlUxB1WSdEqjeIlHl0TA5i
q4fvfJtww9aDFQr2gyPl+z57vXLcHoUmKzDpiY8VeQU3qbpg2LHYk7DF10yugtE/
W6vqXt0fRRbuDAjmHtpN+B8lujbPTt+vD/UuqnX4z8JDlQaedkQU2L9AC+aSmwBl
MXgd5eBGOEeYQorTRgPyynO4eoz7MKdWxeJTceug//gPv1DeIdS8ZW4b+s7QNLVH
dQOn8y43OrSbrWrVH2fEshKnbbZVL0FPawQXT5ZKUaVg1Wys7RklzR/vVPFK1opY
R1oAwFMNcDnkqRZWla14iABIi1uHzK/U8O0Oks0kBiULleIH0pIfnkvmh0w4UVo4
4mkD4CaHGRnT9wfe8LDBg79dQza5/iJdQB1T5JdXRkSGnC/xPqQQmdk3UZ5ASrD4
z1xv7zkvdBitTglBxqWzR6qukjmAnQ+Aa8zYYXOYPJIQKf0EU0L6KhpsBxorhCZL
ycmWXU+mIhRv7xJU/qmsKCMztli4WftIdzaAsEtVdZGmOpSgh2BxjouDyC0N4WAH
Bx4vPe3Wkb/rNKs/HCxBLPsA+RXsoNh9TCfC5AYwUa5ztwHzixQ2b6eE8JIWZHSD
sOOMZ59Dz/sKF9iMyjbgySIOUNPUNWcbS8wBLT8+/8e3uBwa1RzebbM346ADS76m
ZZoG4PfpQsxFbI6jKoi7QCrqEnZ6s0Lg28megCUyWVspdpUtS/luVCkXzp04iFXz
S2nXhs263QDG08fvazgL8YZKNjcsf37UykIRp+0YnidTFUuFD46j4N3YE67NDPwI
eomauXuyxx7C1KW2j5qVKeS03ItEvGmeAu58IkAsRWlrPrw9KGjnU105V4Mi0gps
BryIksdecMQk/kytH2omgqMTBjCwWGOfzLOutSovZDvUuBO4bsS0jeGwzZP5D75+
CqaVNzooN311RSQeBTs58u1P0BXbxRq+AH13H5Swmn2vnzGSLfT2IAgQG1m+25T2
WCYHEVwRm5vKg+/uqS6iscONFAyunSZe+E4Ueha/HdslLFKQ2cU7gYqpPL0jO5wx
M/Bv3OH6O/IY0XF4jFyxI5zTkXuIEBY58kUKyM8RhuDhwMYi1/jQ9LNYgWLzQcEI
OppttkMUYc5phBCP0t83BksXKrRewkM/HXH21HAA4cVw5gAa5Vb11oPvRr2JBkHb
jF4z3MCipJXY8FLMihFsZwOsmN6IWDYVHWk9vjUQAas8eAZcOYJjgE7WlPEDNLhs
yw9VTZdLxAec1RESpqVNuH/qJ98nuInSRYPoGSHpQueNlvBVC3nCaZot3NUf5Ahj
zGBVPJzZBu5XUcecaTbTWFGu6XKIrya7JPtS++KZInOF3qyNKyeERpmybmoF7jdB
e2zFdjZXOjBJaGB9Z/7Zoei+XcIvToK9ymg9iy1tFpqf3Yg130Gx3y3lw8/4i7es
Q6MEhP5rTVPgVaYcDKuN+rLDBVTkgMYVegEraC/nFlcARN6D0NPZOlJZQUo5uAvI
UO5m6MZwOgTpMFfuG8dIwV0Bv9B/pQ74ymkPrrmQtuQefr7LnZrqimzh1mpADni8
p7M+Y17DnEPZa6xAqotWyvsjzY7pOwJI+P82jlWjICBcskKBMobgkWLeO7bV307Q
C0YPMvqb0yRTW8BwSdB5uW5dwe6onpG6WTHN0Im+mFFae8PW+uCk1+go0SNTUqMU
8LJUdaH8CX1EF2TZn21maN+axkuiaTPo1lu5ghNypfNjHJbVoFkX8vBLHN6OWmvO
kOPqDGB6IEMUBgb22lV4KaJEu1ngk/aZR8PMbzZGetYS0yA3ralCQf6aO/agVRgh
2YzdJte/YZrcaHwWoAjr3DeswlYlXmeVWFWCyw8GUccKKXP11SPkCzNynPmvo8E7
niYBFC/n0ZAd084g/5wTikZRUHuIGtkj+M4WIFmmk96iitvvMkST1vhhDJPZ95/0
k2P+ayNpSOiF47eZgFoJrvFS995DQ/BJhhtFhHmi+fDdFXIMdkb2gCf3Qu+Fi0i5
HN3Oh8sVznQC+iGR6ThIeNvbN7ljwwbmr5/X29wZVtrWDTbYUIYFKBHOsl+X2cF7
3cB9pF2F4F4ZrE/GK4nQGMqDN6LsSJvZxc7vdXj6BhR2EsHFAwwUgIg7q0KrJz7A
RM7FYq0JVytdSC5XQMSVZGIcvnRc13ceEsyACt/VP0f2AhgyZH19qk6pUm9rDVGP
tTSZrpE+8TiOT4EHwZcyK5ynoTZZCDgddFx+VHdIefhaEurGeWSV5ArcdNr7ByuN
3o8EYM0NbhCHn8Fx/z6BeqKOxUb989oM6ZgD+mhHU9DzV7T1hY2yxj8G5MqTPwGG
fS8H3SEPlL3UpmkjTriXBshPI6kEdYCS6OTJ1YOgpDqYpGR3b4SuAdc4TEbpKk+Z
ix1kiDuhUkUGGKGf4NjiJRXmPjxXopvQzw9bFdzCULcj7PN5KqzCCGb+/Xi4Ti22
gfoZzPie6b3fT767QExKPVtoPSfKxMvpjwq3BjIZ01HYLpVtUAkpMqHOUyUwnKhJ
GrSlovr/aLShxIvmBxas0Bh502vwclJEqPUqemsUqq5d6iq4EEIJDNNw163kK8Us
QQJoBoYPj/jO1koFwpSvGdNDI7B27BoGHrXg94PwJeISRB44X7wnu+Su6THvApOZ
rsYhQZ3PYwc88XVV2iKkJTlRJ2ZzjLWJ2c394gc5YbxPWt8xe7iysfr7FLrpWv7X
rM5n7dWTwlB9u67l8r4lULd6nssUlhFLwNNA85GyqgBpUkAnbmoJimZPn8g96nte
mf/ESZcTGFeHcvqi/wvhTCJFYRa3/M+zfaE/Ye8zKQxXNHz5CggmbrGEVtOTi0Y2
iBHRSNiAdz4eveBDz5VrJa9ZpKn7QRli5GZXrSb5tb/X+JqiPnM2LtBkzJlgtevz
eez/tKTBDO/7OGH4DG820wd9JidHQOqJ0XO/GXn2SqNQk2JR84kNPrg90KTy2dxF
JK5B7kvwMCA/GZXc+LOHgZQTL6/oBdQ+xc5zcIfc2d+cT7OyU2athRn9SwZfO5ee
W/cX6TskvfLHaRz4acQVlSqUWGo4T/9/a727j42oQx1/yR5uSYIxqD62wi2xMc0i
gBA90nJ+89Q8QRLdJvHb5r3ffx3npTHlRdqY/fDimpHdeK1Iga0WSpEaDEHAGvmr
aGRqHwA2KyLXrC5GHyepBNwNheqmFA79HIAjVzFjdDYd38bU/lNSMUpmI8d8Why4
hDdofaxuo7TXvEvw1TeGBofjvl9nH2q2QOJBeunSg6Pr8t2I2MXYZmV+yjqUzJQP
jnlvcvQoC0HpxferliGBi0Tm+iAAv1BB0E8ZMfJ0Jtg+Q4aVbGFOfhCm8vCNW0xL
5u0hcH8TjSw5VYFC/08mqZK0jQlSiXIOhQKD+b8BY61ZtuZlBX+mG10JCQ0csNXv
Sxd5fpP70VxUJMpWUV4CHCW569vNnBdZtehdqWDkr7HP3FG1MyCPyrRB2buK/KKQ
1vorSCkPzmJ+sHc6GjRFhpOir+5VtlfIw1t/+wejBD3wAGpqg5E2X88zkVqDvN6s
8C7ijOlH56t/JZw3b4CBBhpGa9aUs+UjGC21oFERLALjYJ2u9XBD1cbJaXo7mrq4
dMUXGmp04tf3kEDwX09e8pUExaq3j/MeRXcjCCNVAmprc8IRqb5xOVd2PrFJ09Iy
imNma8AV/hRl4uZj2LMyl929+5NmmJTmmMOj0ykdH+fTOJcL02m+L1HVPsj0QmHT
Mnim3U8cAHPlzEUhsR9odMp31Z/65PIjYPkQfhTROroUt24FdZOxJ+/KBWZRZZR7
zdSQm5bzo8HGlD1iLCO2GqTvJLFAs/oSsV04b0S7o1UDfB1LtqTD2ZQ/vpDHJMNB
UWZRL2yaOZ7CjTglBvtw/H+AMwbWO//G59xrXi2dM4hFoNLfnRIbIVC7IqKJKOMZ
M5PKafkz8baIAohADMKE/ZA7XJM9t77oJd9X4hI41TmuLr0YJaqqhtLRY30+yPAV
N4MylL2Ny11W50hOr6unn2QhjB/4OLfNNhTBiw9pNYJvnm40Gz+Iy6Emoo+0dHY+
PVfVfOrlLq4U/OnQpx25R54lrJ5pU7mYdJ8YZ7EcTzWi+BzU5N7n8i46lPVRTGte
ZjfM5fRHyMxq/InZOKGQPIFoSLa9nmsDQ0HzJRYZdySq4Pli0U6SeKTB/XrVksNo
6myFKaPJ7zkI0KamQCO+Evr8Ld/tAuiQZe2W6/EmpE0XGgRuLGltQq14rTifhaep
4BtVXmIq3ZNTQIVk3xkfv3okMUpbka4lT/lsQQ+gB6ExKyA9o2c7hb3THGa+Y54Z
GyGTwEJBfO8FwDsWP36hp/aO/ANW3oxH6qUFm8Dz3Q+NTFmHm5dmKDJlxM9zoRTa
HlhZtDFBNpFBw4e2ce9NoIzhLm2uEczsWbxnbWp/QwoxUM+uLtX1qFMsAYZLQ/bq
W8NX6H4HKN+y5cHnihUXPpSz9a9FeGgVc+bqQqU+p5Od4TUMoeUTAqJsUZjxiNoo
eDY33qcqE4w9DEIDHN246hAxNX5suBCpPWb0wi+Z1skQ4WijevEzlaKUDwt1dXHm
uksde+Q/yNlPX/HpR2PFAClMoQta2Vr1yjj1aW1b4mSEumx4L/8z3DSFpATEOEFG
M/JvmG2dF+d+FneD7s6RtttQHWJ6ajTpned8698SFj2h7fdpgNBW64XrwJKNrdRE
kB3o8bIj5mkv/bbTqc/q9ixIt/I8Eb0b9oyqBJrsNGohtw0obP2H4+9JzxHL7YiX
Gl9TAN0nRRZhwKd1Po8kgIDCzlgbReQU9LCoFzW1NCOWJE2QAQs6DCqHhXTxFG4M
A5nSwU68m8bjFv86jGtpjkhiNjql0nvkDfjG4WWUlTC17ZJ7P+PBpjdgD07uFg2X
6AIkH8Y2+3j/8q8ph84rYb63UxMR1mX/MHzafp+NeApGzOyTT6qgZLpXEaXALyuB
nR2btoJh89+UqJTIpm9WWiDzQAsnHkSKvPBUP6yNnCzN+wo7H3ouvMNtfajF/yrk
yOH0NG4ryzPonm7bk40Tzv4IKvcxuvbh51ixWHYJZ7V8U8TToxd/PLW/tcoZgFHC
69uy10EUKPZ5WFK9sb9eidoUfXJqtj6ZV/rCZ1TP6UgFcckR+vAzvAHKN7ftlJgI
SlKnm4BZLYG6phM5Owx5SnKmrxO5ta1rqMf5R9+imX/TWA2M1Gd6tM6NATsL0x5s
TlPPwEJBHtBWKGdYgbfyQ4dR0FjIHA8JAYANBHLfB3U+r8zgZm9fB/nJvv7HsXy9
wHkbIHi1IRYP99752c8CWinMWkX+RVigKH8GRzFKngg4oB1inuPT4XQu4Vj5/rgj
8OyR6ZaIbjM6MtHbs4IHCLOLrkKODg9pJPIGogB4CJVB1KW0wHd0hgXky26QKI6L
T5+rxe0VT+gYdrmJW40IfMpWxse6yWt3XtNsTyVLdcUpToTAnHxo2cq8wVHxKrn2
TE1Z5L8MMZJ9z5iqF86c1fvGzF92ndBUiD7aXrBjZ0wTKV3dAj50wPEkqIvyFztw
B/4izX/5CkV4lXjwUJOG7UK6xOE7ABqON5KIxG7HBIqBnoVIbvYgV/N/uzO9YN1u
lriHbkiQVjBEfcaJhFpb9Z0JTLyOs6Jywv59ji4Xg/YE26Ms2Om5ahka7xbhR2Vm
oLPFgeaznRN8MoEl7mkF3I3ezRz8MzUyrbv7WbWeC/d0f3yTPXoy6J0UDNXC/3Yg
AlNGamkcfOHp1o/IrVfLxTDMze2YN7TdZ9eYMnGnsn4+DoBjkjh/MnD17GZEppyn
xvBTMTRQZhTQ1zRpEx/bBaK79IN4v+69tMeEVW7U4fiXx5mbvC2kLOeDLf/gJGyB
Nn4NCqDHYbGl/awTIXSp4ottaaQXkw4ogitse6DpXLdQ3t+XN8R6cWnQI+eretPa
Lc9ffdqWMHGwMTvUnzLUzAieiE98Un9kZMqX/aEu2jsa3FSUyFfPwaFNEQD5dRba
2GYBIg8C/UynO2JsTv/vbTf7MzbepqTO7bdJMS76Y8Sk7rekCOw44qTGoLwZVrO3
/Wj5aUUSLm9NdE2uFA/2/JbkxHaehLUuMjaL/EGGVX2lCP0n6+zM4kOgq+dOC3AB
3loT+Ejl6RYcohqio/ntOm4Kq7o6O927/essMs022MaR9wmV5jP6FJFrpBpxWSAs
jzIS+cyui4WIv43BhBpe73n2YnAS8nY/ICB50y9TdxbWnGQYbj6YxxWLVJntBF1/
CsPX5iJciTh71qlpItFqxe2IiW3ERaUSUmqB5b5DvBX0gRbrq54wmJx0L7WGNuxU
8345KVckT+m30KmPJkbJDs7+S7eBvoFBGapUmX8+kkuf5gF/j7M1rf2gLLLidadT
n8oj7tcpfcgOY+dE2RmTZCysE+lj5a41+RLshEtiRN2rdsTngkBpoJgMi8obH6C5
32YFQxE1VlelBinRvS7CqJuAb+4WYec/ENwhFW181CSYIL3Z2ih0FPGy/1IYbKsy
6CfNHLbALeFizDPzS+JClWECEoshumzhbd42VZkC9yOLaH+F0oo9vku+JemIp1+2
Fuf00SRRec0C3ATIMaBfY49t5VQEXwi3GYfxeTJPNR0POkNipt9jcsZcr5NeT/hn
50QSA++5HAMTC/pkgRbwCwaWAe9JM9pq2LKZ0cVuNU0IpqjluOWVgZ6eB8p/WBk0
Mo230A4j5OKDeC8KsdLShF7grA3O/EJiaekMVxUx8IbQf/kxCFNd2TjtCSeEh8fQ
dVrz1Dqxb7OxBRwZYCYCf16NoUruiZuXwVTL+jiQAkhtS9oBw64MKQlDTn+UmF0v
E6r3YT++6X2+QSo+tVvAa15zM0FoLfZNUIK2oWroIsj8MjqUMTnxkiz5VAsCXFd3
yDvJGXDq3C76rulL+Fy1ircSLgeyfK9eGSX0+1Nq8JMSu+vfUcaMkNVfk9pQ20U9
Ya7m8EZ4H+M1J+EPAuq35WnCZsF8LcjdqX9qFcwtKVv+U+FYiG+gA13v5yl3ipen
r795YLFBHzYc+cgchD77cZJ+Oavt8XVMmYLL/7WODJ0+/g3UmfKyOtX1E0uyZViU
PKoQKy/6P6rrszXxYOUxAh/WFk3kuFuM/PYD/McRsPA0Od08e2s12phzex8SUBKv
nEAhA4CRhOHQjxtWJjULdto44vA1xypf8FnO15MpRby8xZw8oGqKByymDD7s06t1
qwx3bTxPFgztcU99ZAtNPvnwGLLvwxhblNv3Y/3bDPbWCYIDnM8SmsrynR/MxdGa
3svmaSd17tbNSV7nO8fx7btMC8fSAkJjth2M4yPDaJd030fZNO10Dp2r0WftbkP3
F/sBuCJtIJ/6LZukEFZY6YJ25KjL/gYpt7fQQYJ51Bd5cDgdKduoFc6vU5+Nua7a
c6PYvKairBOHSMNqMS13u5SoBqpb6KlsY8M1Qpr1ZAtPJVYS4FG6Lj8HFw5CRKM0
WutoZlX1CmH9UX+KfSmr1fSyI2muzz01P079i88JuKjldvXGlKzEkLDBMZvtozC0
Xehe82F1fkh/f9BHzvU2jyLL6kA+ji0eTV7Ecwdy0NHzVQM+SIfmzllZN2VJZUsx
Qn2U7pl974apIQUXtgCBrd+uSQnvihT7TfRsuEfnEllX8QpXb93kAw4q1ToprNTk
fcJxqDTk5urtjcBX+st1I8qc25YyTSzYr5cMfaEJBtVsYvxFDnmY9ZTjlB4icdk6
ZHkPpf6Tdlg3KQWR4eHxosKhBK63BGtVMDSZclqcYvn6hLXXKkc7fiQIrvvSyrt9
ovEgR5SP4gWP/+QmqFhFi598ARfd1DIG8Nk16OxwFPPetBAutXY/JP7DsDFG/6bQ
qQbbjD8WYs3dm7NO7mjMxV9aZPs9nNIesmDsPayVeLhU0u86Q9m8X292YVvwRA6L
UOldNJzSff6cP8Onll+rDuVphC8aqM1IARNgJI8lA9eg4K0GA5Zb58WeLyLthfhl
GWv75YpYE4+CXyUIzyVw0tCAYAJDclwQ0mt0EevxBY5MjcWI0qPsPE+mAWk5i4P0
KD6kO+rtAVClzif/5N9THIRWHuPa3RKPfVqeRRW5i36cjGBbhJ2uzjWPlkU3THmD
d/L3x9pfsv/u+KW9D5XSEOXhe1P1djWE6wEYKo5Lwd/UbMLB7B3aJYYGnWU8rwQO
HNtqBuIuvCIEQ/1ImklgcoR2glfKZqXxRB+yFbm4mWlW9ttfufHHg6UUeaJgN/3C
ZeUc5MsAeUZ8kfC5xuuK24G6JDxC4R0XdgAWvlwilmt2KUhucIHzVziCYgq2CzMf
qhr8lzv7gXTvCzgDpdZvH8gzjQOpyUJy6wGQLsh/3MngvE9/WK2W5ZByszeP4NiJ
bX0U29W+cOtrHoFoSntW+N1LKYMK2l6I6P3mJqp1i02fRO4lmAvTsv1MdHuNZ4Rp
D0U/C/fjmQD8H48tZ7r2mOxbV6HDNVBSM6n8kXobHMpmswH0iMD481dpAAOpk3Ys
rXP5nvxMgAmRG2x7Abg2TMQ2eMOIRNgb67RvineFRO0CL56aHB3eiUPKeTC0bA2O
Jj2fP9oQEmIBA/okAOqOKukPXpEd7mdckPVW7AP4R3Cx5tJiGA0PxonvpES7oyIU
SNFx+SvO13u7I7iv13WHUrCs25Amycgmv92yhvhNV5HFwGwaqnL+el6l/35tFzds
uUKIGXu/6dfAzx9qxgLIQb2Gy8LFbwNhpKfwFeDj+TpCXRQ1c9W96ar72CQSiuK6
qVKXdtlXWLr3DqSqv2Wz2t2xLKHwZTfyHIA7naBdLkIG3dQG1QyN5763uR7e0nRp
ObAnl0Wi9Bp6Kn4nTdIn9vkbgeUoqgbNJLIuZ2iB/YqtznUyhXP21A7z9EzdA9OT
eT+XRI1BOg01G15UJa7tUMeK9I/ABiu2+usBGj+XUKfVQdDFNAYEU28u2dfzfR8O
UmhbihjJS6GDqXIYUVNItaCIRGwyL4mkXc/t8AlsJw8DU0XIpCzHPHC65xU5WHZ1
pq5twjvwZOW1gVs5cPyO9alFZmssWI9HzYUNS+/qpMiGoOVUhmdjhLebyK0WeNdV
GsIHqATdS/Z1xIAMtd0kkQWNiJ9b7T7EE58urNtksgLUwBDXru0yPk5mb5YlRdAh
Eo1JcUjm25gHd8h88Bkc5vAR5qT8aN/NHuYxZMDrfqgj8SGIWD/x2Xc0vEXGRMTL
SXULRVDzpAcH0nMvzmkLz5LaS5vXdUtqIEVkieN2d0giXTQPFp1kKerDeFArsiHu
GugE/7RgifJOmwpaMcyXWxvjZ+Xx0TPIwk7XdVLdNS1+EZeiJ7IrT5WVkSOMgLAK
5M4HaoRqMp5GpsjQfxFQZGMsrKcqJ36hW4eptuCtrzYA8fqervvLnqGk4iV/OS91
B4/QMFGLVMZDuPNaYUs88Apn0NgpRRTQHKoQfrKeP4K5gRbOWt8yD/cxNed62Bfy
45SXgwImyV1yUazJDq3cWebfEh5c2bWv+ohn8cY2fgpYSFRu8yRLNGdm6qgWdcb7
eEqDgdIyaCHdu/Gi2UkMCG/MwxC6O2ic4L1mqFjdSzGib0EVW7cJk30XblSrjW+J
y6ctEviSwEoqNXI4eUMtl5/Y6JZBXUI8XDW7iQ/Oa52cha4X3TyDobP7Sg1+CvKP
Ma9EsnwgyUvHQo5ZdzVP0RaTXIY8E13RRi5jtyr74qidK8Bk3ybEk/6LKSy1OPD1
/rjMDAI652BGNJShh/Qxc3VMtFyBnqtONxotEiMtKeqBjqYcYQVOvpXLfj+0FAO2
ot/PCj43x/5mCtHat+6pvFx4PeY2OiZgQkC2r2NEMoW5Oee9yGJoJ6R8HJ2gTGsH
tCozxulE+jF/fJ4lLDK35VZepSut09Hid/R56wJTUOVi1DdTj8SdiGPUobQXukk1
b5kluwpEyME/hH1phi33Ax4nIKfdOjSKNBQpj6/cJLyVU2jxw5yBXvNXUBYMB/wA
A7DCXKSFqSMM/YHuURY4ZyWbC/0VPl+D/Lx79XAgUSwVi4NdEZSqBGNy3wotWnUk
cD8jTtGtww2bSemTZ5sdp3bDP1G76MGpwUPDeqMhCbyDaSb/1IaY2sLX9Hb8xoHh
RHKi1PoXqdMUuSxlNnsVNkPZK1JNXkbZCFWo7X5+RpwREmXnQQpZbpZbs2kqpGHf
dYYi2LJ6Q1+3+78NziLxCqbfwMC11zEU1GA5GFtp/lS/dUS+2/m+hrxvmi8Qp3Mb
3A8YITwrEtS2rqsQWITlpJnf9jiXmcmrC1NQ72rauvL7jERx8nhbNpVxs/l/mCv5
zLemBwm4VO5tsNSr8EFqXJ0jMWVeS87I84uviIjrav4PxryFT5kXg3+X0BTFvuG8
jv8tqb+I7ObTdjDOTaDOkH/RtaweQSGDy3xEpHDhw1YvptG7Z9FEk7Pkg6Ln3Qe0
gidEDdn6kVfgBdAi5Hr4DsyZTc9ok1relhLhvsBuQvnXWU0NkzYm41nBCMm/gh5p
Npu4OrUYQczZakFFFBiJTOJiLFeQTgKCE24p2nEiOR0F4Phsz5aP4+ncW+zo37mE
g2ktbmlYsZXNQ9Npzr1ffasiZhP2o8dHjITvxK1mMAxnJlH5D17dV3NZ6fMG17I2
Du0C+nRhTRZPaa1B4hy5MMkvdyGEa6rCdh6B33yzsCYm7hqsn29FECloM3mnMt0F
ClozBMaiE+lxOpEDJPPXhByS022dkH1woQeWPIHhazc4KgnmosP36hJ39iPKiizA
GMWY0fRxJJlbyxpHob1PrlQcl1osLFFFfRW2TSfTIbw5bd4NxlTmp3c+nxV6TIDV
TCYtuw87mEuWXmxh0k7b0J2kcgtsf8tOXM/A3qjLvNZy31dUkQaXOLfNn5Eiflj+
Nb7yd6DnZKeRFhCYZxyI57HXE4Heo3OMQmK7wXlr8iNbOl/+Bbj3NoxP6oAgOllQ
ztUV67ysSNEQIDtHwq+NG8PP6J+85VsgbLorXXb216LLdxycIaqbPWF1kTpfT9qH
OQYztg9LAK9Bwbqp8u9dPBXYRE6/g5U9lg8o7AFeQswuFBV4fJQjjRwVqKikeppJ
iklXLn5FWTz60bwug9+EIlWGH0+I+lO9DF65T+GukVQ8ejYk2c5IpgoQjmK0EpV2
ZoloVfIahFtfZh5msD9Q5ity51QH34z/Cnq20n0u3OEp6o3ER6hX+HxYc/32c+Kc
QcEm/JASENNqFXAYtGOo8FJv/gyke7RwaDO2vSJge6Y15ZAdkMyuLKpFAh9PXSqD
ImGl85HOr5wVOOw6Axm4KmfZmiJpJMhUNzFqrg+SboketC5dHR/X9SM4aE5II+/9
SsIqRGUDK2r2VZrbHU0989zz5fUPyT3swNkZJWLetm4tla2M4PH7o25V1wRQ/eKy
w2r0bBgdpVTHv72GFghg3Y6d6YJ8D2b00A2NAYrNOmr9iT54VC6KbBcaYaMXkC+K
DSQDmOCN0eEOjpbh5Rs3OE7GwMPjj2NRGEa08MRhzPkMIyV0xPFdEAUgb9HY9Vqy
ZFcVSFB3isNp5n3IzhAp/CE++WZ65XFEGlcZyqh0TtZtbycpzK2veTtL6wX2ALX0
x5C57kOUIZ4hvudaQUrvpAdlqLkHhHWHFQmDVYiiy1CGkCpdM0PaImRLnx2t9+z4
4/rbRRTr/st0cBve2Ivx/QZXQYZA+s8LOhuuqZFKeoY96Mogj+Kqs4llpCkTmE8b
b17U9noD3rjPuyI3zJzTJqJv2TYAspI3qy1d0+KtQupUPRxjiCymnE9v8QCWbHwm
sSeKg05h/QJ0u20TqtFA6mBEvlLqgmrhFITSO+L4FxGEuMZCig/tkqsPGhO8gkzM
8TIsjMRjp0ZCPid/tSFQ5BDLn0l0SZmL0j0F8j96YSqpsCIhqQHeGobzV868rTkx
pIwmAi64EDKW+0y885NF/ZWO5wZbXDc9eQiHUZQyhVkldcOqgpfpMo9aub+QQM2H
6QgZiFYA1p3lpIEoGJQ8ln+vnv4JeRjeBY5ITxFG+v4wMu08Peo4Vx8yWj8HEn0a
9To0kuiS2DsBR7Xkl1Bkl9wdL88CSIGuB0RoQPKEBreZysrqyzVtWrDwqazjLB0B
WIydg8uKshRp2Jm8/RSIQjeqOqmDZuUujbI8J1f1kxBxd4udTtvU9V2W0YqJj3qX
+JZWIPvraqCJ3ZnapNtn6VwwHLeT44+LreXkC/Q62qTvF/QYk9SslocIaxRKJ5+Y
QpVM0yiO/gtT58hzse8BqU5HHN3j0pnwy4gMvMBQlk+sI5PfYjTPOCv/4bevAo8M
JzNoSFf2bVYrR7Xf/vGCbixWDGeNEFb0FugGNxKh7pw0xsyXqsfAxFd7/liMCbtq
IfuIdAleNl0Z9cG91nxKrdst2LWYf6TWnbZ3xMUiKG9N2ROWqcd89fIG83GS0xZs
9MigUpodOYbppS7tLLywFNtjYqIu6zVzUUjqf1W2JJQ2oIBmp891ILIoNND6d1wc
qquMk7oxN+7fkn80JhEdXu1goRV0yo0iW9yEEtn0IUPl+QtgEaNulSH5WeKLIGMn
VYlQ5xmRnoCXTww33ZFAT5VJJwacjkR7SnRzEziwfthU2QTRyR4bomciJ2PMmjPe
7Dm7kJUoifAIfU1nDteiiARiBHmW9Ki5G6vbeJ9KXHQbCw08up4Ow3aEAa22MY6S
FfSGhhdkqqYqoAbI+0gidnusIAaQeMSnGb+JoZ38AC8ihF8Wm6oQnzZx+GTcvd2f
TJqZyhwFGRFtUoSIFwVxSuAV7AKEOCO4ADHUCXbfh+1ZpKK/oQgk4h8oY24ooRLJ
ePzno4UdBwJtEoyzKFo3n1yfWRZthBrZb8PhwglIu28ViCzwuFqlG5GbVT/AGh+j
kVwozAjS/fyp5Z9Y6B7fGIjInzznxAm5kjEbzMPlSEpUFmzIkei9gUANM0EUsHvq
BN00MGZ/HHZtXrhw+l3XONby1EQwTrF/C9COSuwA7JPTF5sBM24CLU+nsbfXT8YN
AHsCGru7MBj328OSeEcchLlXemZZ1sEsmJ67lQJcgK7Y7IPzlolLHM1IFK7ihoTo
IwwhHsFq6RfhDMjqL3jz7hr6p6jvwyzoQ028txnzyZPjD+NLv/rtWQQHePUbcBPJ
DrDySpb783oxattp+/caI/YFwT6jEWFjiA+5rMVuyWNFgitSApDvqS29JXbIWmsW
j7GhJlTVd0N8p09sh93YSa5jaQO+v3raI9Yau119etzbLK3h3ZLnStvMjaFGHwwH
dgb8/BUZBC51qBLmemTLBIjyxobkaB7VXIfmfPkKMmqWvlkRolo85rf7NrOA7mVT
m1qUr1hMHbNyYL7L8vLcIR0rkZWPLiDmnsjoh3lWD4W3WZUtdo2TJh07mf3fXrej
mtLIUFIoxJ1yIdDNoCjKi+vZBRhPotfrphGagx3s+VYuK5BBcIZ08z33+d8M3k4E
Zwp5fYgtAoy+iuhtPWwEzXiR46iMrtKn/QHRdLUxsyhl3yVTWUto2fEJSwxQH1rq
64clh3c2fLMNmEY/AakomC929OujuZpv/0S7efDENB9fml1gJz0VDtvVDXsbTLI/
THq84hHSXWCUA3qcjOoaczUFWni1sPCXXXK1toA4zFa3stl5/o2x0kHzinc4lzWM
Uhd51mv7owfg82UNcDa8dTZzVzxaDcWFH8NYJ2kPDIbkAQWqWitOwgcur0J4pdHL
7KdNjJSPhX69F6OJ+UGHeixghlOp4bCoJ2kv2LUeDk8QwaV2J+iSREu0IToAbYhg
C+hSqujEkxaszfu8CAxd594oZJS87aOmg9Sev47JqY6w/n+hVXsh5rLlCzreEUOC
84EoxKyeqLgyMbaD4unKqZ0lKaCKdIZBnYu3fkGww00cVtAIR9j5tG6gPJUUAcsk
dCz2fMlDZRcoIivGMpvVAMBEOjZR6o7wfmifwPfw0w7jfinhs43HXafVVCPjTuV3
L1jbJKyYW8GwrjehezzQl5HtcAU69vDVGOBMQ1hfQyAo7sDkoCDJ4FPxZOJzZ0sm
TJ++M/TAcB7+QbLZ0SXAnNA0BCL4cYBB083YYWC4/IGma51N3DvgaptupEhBvA1D
8xpNbKEjsarFMNgVCFI9NvMOV/AMnxoZHf599IynzCjF2iV877O70Fe7k1Ats3hj
kSnTDLSrYB+l6uuhLYaCC0wqPiAxXo6i0r8nxexZVptlASa8pgifn1umJRHipzSn
2BUO3cciHY1MXHuPwJ6nSf/QQLqV2wmvEEUnmeQZN87eC7kw5VRw0Dsug1TimlsI
X33Yxaevlk7j/6s+w0b+4DLe08+s5Hs/6bV36+UuaR9EAFuQ9xtPMewy0n2iXsp+
+d+hsUPD2YqIiuwNH4L/wtxQVUA+pyI1QgXOM/w3Iu1nHW2+Swoa32c3gOtbM4X8
utSO5e26/d+50g22zve1EXv5YZ2IIakLLQtWpbgi1aBL7Erb355dPEuqoYn8gGy9
O7FYYxMHj3rZ3MJWfTXXPts8STRT3O5pzuSaGpnu6X62kG25mJ4MqSWBmIC4wzKb
CNXQC3TAGKltf4gZmpigevd0K/l38WX5zalVK+SmMtfuuv3Kc5d6egUACooTCcHx
ouObicfS89NG0MjeESKeuvtxQBWkijb+rpHTRKezCcw+vWGfmM4zNKmvicimolXk
gn4d5mCU2UNUjFZsvbjQlzgzLCfR3DXl9bigdsgc2umzwND72stp7K02JMBa7suZ
LWnHs7cuB0AZfu5RXaYFVUtLk4TnZIUa95/b3zF29DosWQQ+p8eM87jUBZuMobCj
2sd46hj+Seys/w24fW5QG9VCxbQHn7dGPf5DZgEALZ4OWsgLm7RoRuwAjDqK42Ro
CQpMuLsTxSFOwGGVjybQmFrtN+qEQXjzxTwHIeGeGM4/7DCvXemSHvMGdBRw+SLU
ISxUWn+eodS2Egp3FxMUjQiG8aewimROBrmdPIJmG4nptXaoykAYs5JMUg+MtCwU
lO7KOUT7RNQ3JkcIoq2+jPfa2EXXwXgdt7E1PZxtfJZrfLYiSVCKnKD3UohXJt7H
J9G9PHGBSv9FabfUwLDsNCf5zjn/XMqgNRHNJrIMyC4hJgaFNTZfSrvU0PJcfwVH
/U3VWJCbjiMoQaIWftMw/2jFCNYxpNHTUt6XhR2b032ruWBrZWJrRcMTBma9Kd1G
gsNxPJjWB6m/VtvvdciMyrkiMGdPvQR3S+4SWPALrkb73eH4nRN325KzTWA6m5u3
BynIB+pRflEXQM9UkvYRWLbFa2Bbbk0bnhute4RwjKAZTYJ+mRi93oCKSbItfRzR
hvPAFqkMnii/0sg4/GTIEFQH24f7ga3vjbcDIt5JYQNvU5NNyfZdCAlG6zEFom4p
3gxQIt3QSDvgXWPsw9B3cTVCd4GRW6mbAO282AwpEN3hckkLcQT21Is+1cgqDK5p
eLvysgVnIIYFMePikOyhwW6B5NV/OGBKbMvpxsx0qq9m2lSeUgjGI7jljcJ7iR7d
StU3JPuzRjkkRtK+HjRVBeLvpvTN9gyu/dPJyVW+Nd8240sdaAS6s0IvBm6D6EPN
rj8va93rA6GHpA8KOsWE2lWy+lAhm7jT0uVUsSs5pwEUVh9sVWLIIAWJCl8FfevB
3GYl07EqJsFMFEN0U0SjvTIiPUgh+FWcBDz4p18sSjKPFy/rog9iHoFfERqxBISE
rv1XvM++Nt1Zif0i2deYwNRGZNLLtDwv6U2I7YNNEjQZdBFqsJ8OpvhoUFm39FiL
e6Q3WKV3qc3A3aAJx1tup7EZxngIpdyNOEchwRcEOdPX0zmtC4Eym/M9FK9jU+A2
Fnp/KkFsXZ3tsX9FqlF5aJcfrLtJuFTByGyfVXokRHcxR+SfbDwV4vooBBH7Q34y
RKRgySkKedb3KsW1WE8w38lgkBdwibT7XYArfm5dRPdB4bUBY+CwMh1LHwMwYjPU
/hFWzjorYJMtK9QKYejmLoS+1EyxNY/9bUX8QemTbjKrczA7R63YQQQZQZ3Geb1m
Tar0u2ASraK2WKEepR4SXQUULsYBkCes1XpJ0J4KH9TQTVZtw8vN8LsbRt7nJXvO
RbjaC+yH1UpI/guGZx5PHc0jOUffU/7gk9X0WGBfaRc2kvNi7St76zMs4je0sDJ/
M/NiIeRPNTSvLtAKxa4zFKZy8QKyYRrhSppxtXnacqEVgKGL7+bho/mVNvDKVTA/
ZA4nWEBKt+B8tp8YKPi3XzG5xWraA/XcugV3Tiay2YYzxHvSbe5UcVkqz/rrWVjY
YfpvoVNCYwF5+LLxKE0NXZRKPfvZ+dOI3YDaun2P2WdFTvOBZq3/3u7HqZ+4vHTv
kCXiOM6nphMqzYS9txVBeoqPRwW3yP4CIQ8SyY4XzdOZRNK03X5I4q2wzMVdiqvO
1S31z5gvMDyls4SNNAYxYCrBsUbn8fTkdPb8+E43BKV1rOCC6h7lFjmXIZq93CwG
PwjnYo4h83oy3bLwrUdWi/I1xSzjMzGGEJyv6lnj0qKNIgBPkKXrNk9dErXgYYaZ
GuFxmDBU/Mf4D2v9ChCQ5Qg+90lmV2R8ApTqv2pEEyf9Hprd/LL+FuyXfa+No3K/
bmuY9Xh4VMQpTMyxFRFcTM9I6VaPilbOKaVK8Xj3WOhPoh5fT2FgGz7Bx7UDxoRR
kZR95Bmv9S9fsvNxI4ukPKT7oH5V96hsMXHKAxoBn8jalX+nysCM5Im1Yyzv3lbu
qFjCktA1qbSruySQz+pTWFHvMZMMncMEk5c86QNGhe9/5PEhoRzPOV9UfQ/Dsgd+
KCItpM9QB8BaHlsZYayy8Oy2baKDJCEtvEad15tk92kEiW8cKWh/GjG1Ea8iFvwb
G7vvYDSGWmLkyad+JXg9YeKLLcnCHQzSZvsTXYXKAZZFLkD/NvcDEqEXEZrFD2dd
9c3A11bOtlQRLCVqX55xv8CebVQXuv3t4TE5wSGPYW/+4YQQ8ptu6WXKK5z0HfNT
KFzSLKX3Gil6Knk3gE3/sr+NWUdkKl/FoFkUciSsYk9rkibqDELpIlL6ZgD1Gbuq
G7K+rCy4FR3ESHXSd4aw0HvU/GlVb6Lm/Np1SpEF6yv2SZcPBT3/0dJed+PC6RzK
L0MPGFBxIm7Tg6NKmtm8+docChvfx0cCLi/74n4l9+OITniLfms+bZ8BKRNxysK7
StJ5pv6TXbbEBvu/VXplzdpgChW2e+P1cXncFmKtCJ6n9Jf55SvtMa8qFhkIS4ZC
NmglnsZhplF/i54hZ4TLXqEgvbPV8/Uf6NVysOMwYSuACFhVnTXYj5DkjFSYNld2
VtS+Ipgj6Z56wfPNBVCQGeDyrLz5r4dpDa3JIvkAqT22U3fjr62IOCq7HMZ6Vatu
F+ddT2mheoxll4NfZSqu4byja7a15o9Ak7XKyCfGiEnz+kkEYaJbz9iK6NIgQ0fA
gJ/r7KU2bul9+xR7iM+GD5PcqwCWU2I4wJenuhk6byCekpYMTZlI3xLtdmlYnGpj
rP5AdDkjhyCHhoI8RHA4sEUGFxfoLJZyqgm6+CUoP7MyuxzgPPNqoaELkhg6eDlC
Y5l11QoxvEqgpGFEn/qy/uKJwUSS2IkJSsVzzoBWYt1oA3NZYmaPbVy2U8AQLPZH
aY5SSI+Xv/7EZ5mmzQr+gptDxOyIJFRMbUFowmPQri7Tia1FMjGJbvixU4utEKDG
8SHXlhPf61peH1HDdG+YvKK8cCpIOhHpNueTY3qKdK3kXcAeyX1M4nBUKa46NVJf
8p05pTZf8GK0RqYBJkUZUwmNNXE3BsUZ5+TbNrCyMCULYz7Y2BmEofd2/pFFpz/Q
XYtsMbtIyJnCTsCwI1QviAU/syTl5IMMyFcGQOp5SuuDJs2xH6IrJ3CYyWpmTKUP
cc+sbZBwLiWXeFeQROW0awF3kE1trMHUvCKweChAA7Exl1hgwiZ1La+5jSFH9CVx
SxQrra9TFf/cD65KLWBvnCnRTGqd5Th4taQvDCXdpaFnMSrq7EdY6jQYu/oA20EN
smi93sgp9iANQA66CEBS1NmZJbSWlPck2rG271SEWNd+8lgi/H+arSvfymppcd88
4YSQ9ybuqd8e/lvnRtxTpmdPqWPezKoYOM+4GVrV/R+0U9u7pzpoS23jhhJpSrQP
9BdmbDNfjsJBuNnQM9+R2sxv2Zognb4+v6P7Jjc/JU/ZybsyY1alCCmyI2aaLsZq
GqLItWHGuIvjTKTxP5M6rYar7H6QR+cRGzcWVXGdJKhZrV15K1E/gQ50mts9U00Y
4EG5X25HR7t7fGf0HNTb7nzUvppbq/6G2qYwxUzUvlzAA5rvQAnPI9MEkKyyujx1
tthvbAaxvk5D8ZkZ+s9M2tq54JbNOqFKjuWqJt83ckRKjFEL4r7nCz83kEF3I3JZ
SQRVKWzZ5E8HM6YAccAw05tQQEoqwwkVZyU0fNkDfbNGhF9mx5znW4ZO4OryjGC6
hn8z2dHVcl/UTZ3ZeNEj1/Zelr5hBj+zPazADISNtgjUlCId+SlnPjCWwaxKPdVJ
CPnm07FQUxRmMakPtqnRDvf/HLgRwp2zckoi7D9qnWPJyR/ZbLzJP3mCudXUy/BT
STVmevxPVQH1/BYcKwZXkWnb68AB1cOIy7nvUVDYrWA999mwzGmPqIft1gIUi8QV
qHCYojo5HDVd4mtha/fswURNF5hRPhQtv2i3v6Y2QW4j+21DmjrHQ5BwPt2v5dDW
rtzciJROIHGZwyb4b+tjQmWMgPRAVNuFaAHjeZp5fkYsCGY35jUPHEB578wQ475o
rc1nKKFRvHGjTf0wFhyxdq7K2FB+Utn0f/MWL0mZpNcqYD2LFib5JbUS7u4AnGav
2gfs3O6dZ4TSrzQiSYzSZNZOpv01D7JSS+qf6A1vcBTB/sB8yO9ituAq/ZcNNUNS
1KA9qqOPU6AjiV2citcNHAlnWvZw3G4LR/u4NltomcUAg/22mtfVeU1MifeJgWG5
fFqQziMwps3YTL6bTcr4winw4wksYb4tvuTY3xNq+PzTPHvw/7jkgle9s59c89Bo
Mlg7urRr/RuAT92KbTC6MbkEAWByFy37UkGzt934utGx9iGQWpiaOu2EXrvDX+cG
yA81Z8LS+2Q/eBa0ct06UORkAHxYvke26SepLMW9Jiu+x5i5qTfpMtfRRwAx6fGk
6Xq1QQVZQ6iRXkYmU/86MSmHgEhJyGRodCnG3LynHZWV5mDABMA9fSeb3UQRjemL
UNUppQWoJxls0+rYSNT6zuHL4gvajuiHKOvjiSqOMRrDgfyEqHNNhFNCSLqI1f0N
DKVkzVhiBU+8tI6ThoXw0aQHpUrnY69w+uqRTJAvka04viLE13pG4hNDBWvu37Ek
bXrPD46BjGKmUMEllC3T7E2CPdbzbY4LEDnc+47YSwso2XsNBhFPWiJk0z58/4En
ucsDy44xzhB0KaJUtf4KDigHr3sqBZt3b+rzaJ1SFHb1EVJctNsHArcCkbkspL0Y
x5OMdC/T/bTXI/htStLzxuGYFAn+EunxQmA8wuS9AZlkp36xpIVgycQb4ZrZ7YFU
+vX0Wa0yMb98O/PBKI/AR2oyYChE7d9imvHSAUk6QjL5TLZOxHBFqsyMlkO0Rij3
yNwzzDKH3xD/fA4bcKVDocE25Z1/VqXlyJ+yBWEGlwWTbHMa323k2ehhkLTZVgXU
5uOuH97cwhxVCN1i2wYNI0DzC/BFZXF/ztd1+gM/yNNsTzT9QRN2HYzERp6DJTdm
cl4dON/aYqSKLU0HRZ2Qytql6ATke0pcWLH1xLkE86T1w1CAGrghYxtHDhvsx8oY
7Cdnd5Cmz2xz1q4idcbRH9dm1Ci3I1Bx+MtT0Rdhps4RJ0RCEags/H1OYJE31SBx
YEpDYbXTI8zllRF3PaIFyIw7huKdTCx9xgakhYbKbtAQVRQ1uVGxrFHEkSjgpIAt
aDNnkoUJPy+YLWOilO68EEMYChDfUtGssc3eSlupUuse328MFYC5sgK7L24QmBJo
/NN1YZpZC0bHaaqj3QAo8tFT6/auaGIV0sURXAHCZgxgzg6h2sPJaafjIhGMdzUA
e/hYOxf30V+02oLf3yGjLP0jBx39dZgbpQ8DIG8JKpOsBKZO0f62DOXEMq2+Wg6+
qPse54KYP3xRFBE2YikI710R/PwzufCLb2Fj/ezbO+/2e1+tPxCrHgI/6WxFibCX
HWctfoWpaAVOyBtZPez81zN8v29coNhxBwIOyN59BUgtxzBioGywvBSKkRaL6SJp
aQATtLGNjyG+FRcM936WchyQ0nm8quWjZFJU5yLFIGMwwxjEb5B/ynySDIaTq7Da
8vQAzpsv8svesCQIqYfckzzonIKMn6wF8RfvBQL08u3B55KJhXcW/tl4nbYOgUWQ
aH/Ua8yH0tANxhK9MjQPiRFDlPNFzGTD+Roarqjs1UuJ+N2GmtnTkDZ9I4qn9gv2
Yr2v5bADxpz4KZT2wta5mT2NULUJoGRMLGAB0NGb14TG8buFFGRxNNQCHhP4AW/g
HCFjHEhc1ynCWz9nrMdubdCVzOmDNQKbbXhH2kK4soKlS7Ur8MIGT+GexeTbK0Ag
DJssZ6euzoRH1id40elvg2S6pm39ZzluTqg87wmZv/7KWtIc1dTBHs0cqStojIs7
mUDjT32bxYibVwfc9pDV6Br68nkYi+KFqDqve4gv20IrTO6RfQJM2N+yupxvIhY1
FdT37SuP0IbJa6XrYHGG9GBdhSJJK89lYDXQpd7uNvZwnSc41b1JdxYJS/7pRG+F
kuIyezRJXMfIUwFUaS1AS/QXenfsVpEAAb59IiEG6i7VnEu1Fb/dDEoHpzdyzLH6
u+4Wu7DabY9ASf7T7oJLRLX8iuPFLqmymN+iw5dRILpzQzUAwPcGz/v4K+A2Q3Pe
u8LyzKe2u8Kh81o4pWf1R2X8E03U7QYEhiIAR7CLHiU7kquvCJG9Wg6AP7um0+UR
Rb7tydb31IAACagjCO2Hj45LFI+LuguYVcPVRiE1rIPcAfIhViRsLX7PumgSPv0x
cdQQAqgamK+NAwURezJ2P0hJNuVkqtzz0km0zi2UW2oMyFRaGcuh19HnrqOIvxqt
pDmAw7DllvfNIENcDMtYQBWjDtkR1m0JCr5tUyIrbs7IjXa9Z9mZ2ZOZrCl/PwbL
SRffCCcmHi9H/+OWruYfctpoXeCwnqP9bV4ljK1rtn4jiJSAK7FfYjuAqHmEB+Pq
/9Prsu9WF0vBMRHtoI2f2xBScpfCgZ6QTSFRFAJoDrnpCDBVBpqrIVwZWPYXgWhS
aO/P43wXGYYhjKF2C0AzO3UjT6U3MzXZoJ169cWjXO/3+w+Plx/in9Vj/lxT+MfU
mb/SgheMwYFXHe0varxwBTypjyIyoI93N9kQvbNpudv2ulpbYGoapeOs+Ju1kou9
InBDmj7Gug3Xjx6tjJTcWk+eJzuwhhHljPJZy2beuNfSpMhtSD/xk1OhtlYOEwRp
+1Q8okJKwreiC6lbGqhigvPuvUNeo/z17ouhyKwBh7pD2itKPuXu0+y8lV8zuWNI
288Ndf8fZq5uJwZA7Aoeuk+x2j/+kje4XIyqApwx54Fo9iRGY2HjWUC6RL/jF2ZL
KWfvO/HXGqLq/c/nfgyoqshvOZigz8z3p+M++KdRJFxsj7+KYYzctbR+s+uOrAxB
1pTeyYnI4wroF9bf1yf3pR8Obj1IUNCxcX7aX7LrbknnbRx5fGDTBWsxJGzcy9B6
nSpeJxA5UQI9gPrZAk/F22uRcVvrpa2CtBon5Ra5QrzfqZ7JtEsur6qe4+91w6gr
evm4QGlQSn52AWgqAbri6IOUnpbi6yPijrUYzc4xdD+0YVgmj7lgWqGc1my+CFQY
AguP7RA4MxRnQYV74fxbrXj+VBrhUwizBIOKRgBwqAUjzACV6c/dOTyxEJE+9E+t
/u2eVzknnSN+9YABPwFIQ3aY5+2i96YV/NVJFza0LjBN4bnR0+UqS94UBO3e/yeQ
LAi9JaHz8IHQ5OXLSJUBX1DPxhbpM8/weApooYiFDawiia+6oTi7I982ma6kYQ89
obav/vJKl3pzDrNwKE76Y9Igp8UUB38PJnRwcZs+/ucgs11QnqNwbrBExlU9mrUF
hkah6iidZlaa3FGwOdc1tHCT8nSkYbGTksBKwC+h+WF4WemkWJCRyZZOHCel2Tsi
FSd58KAQrCTAwYkEhEMHmt20+88JEf+zPWl9mYIt+Tn1D3NNnoSmGsr4SaEGQBEa
xRT4O5F7ldsFFTu12WX2NJ2oqTpyPFH5DEsrjF0CrcmfykpO5eBwhXqbpS1mxVX8
FMVKJYOlFJ8E+ZsaMENwt+MxzH7wWbpwJdvu/L9loJKl0u/YCfPSXH2GoLlX8mmN
dNLKaYCmwkwJ7EYwggRvu7cK2ubymZuwltvHvHQoFPKTf6xFAiAxPmTjyEztf5ci
sW1io+uLwfbgcKzeSjVoF23cfq4XMFPrqoJbglCLpe33iyDYte7xVAHZIq0nTxVO
QwxS6nlEY/lFn/OpMUQWN4BTdJCB7WrgaRM8da34Pv96xDhBkL69unEBUGOqerS2
pZ48FSCZpzCbEkquWm9kK5SaSES3cuvffOLDMVTqSl+pDYGPWYd6QtoP+H1TyDkD
0Brh0ocEMX4oLvmAptQzRYW7tQeh1rwGQFliSKl3FtJEK+XT89l2Er1mCTdinaxc
gHAkSIXKQT1zGHcdzaLoOd2exgKUhmVRtyO0Ri16OoEnA+EeX0/oZqrNaa9N2BQC
OsFGsmt6Ixk8BRUILBxAasY5KuYjmnRKT7jiz9xNhQ5o2/UylgM0SBmawTc6aBvV
LsU6RbdMidbNuNnS0SSwnwWwZyXtBOIYYC5w5UI7jZtNccB0vGUAVyelkIUiReFn
eeHy4deKuf9BVV9/x1/hvfTHlc9eTyiXaBVx4hB/VuFRR6PbutVsoMFjGYBjfj9d
1sKe6DPGNBezR5ysLAi3AOia2Ek/NWMWan04B4w1H34pYE1fKS6IJD6mcEOikg9G
fq0/UqsddEvs7CghtRQlES0NSOOGY5dxZ1yToEERAK8smyABPpiZ+huamB/zd7y9
PSx/S4gJEP74ArUhS0RFGQHoxgYTqte8phY/JlA+ol2bnz7oWVHMRjBgRCGWNdML
dOUZyzY8FZBJh93Kt+Ykci82dJGP/AKgXuZctqh6uFYPdqzhjdzB2hUNs366r628
WHprSgxlTTzmieyO0B3EHzQoT8zwcivkC5YlSU2RxKhA3kfTFF2EKn77RuULU72a
m7F+MlBKqEfa9G4dOf4LTncGATLTrWegrlpIyAhUegzHwdiEeL28eQ1IfmNEbORn
nFjDzOE93URgrmrsiPSR81aAQx97NYOfbM19PJzUDJfg7p7JUkuVX6JT5F7xWFcH
CUTmStEUIlNbKlA/Xb97j7PPOWmHbEK8e+tODpaIQB2dElyTjhtVaNQ3LFiTQe5o
Ji8cLLniRpDjDigMEmqbbx0IwSk1kaAU8EZBrN1pp5K7fYmxB6NQfn5qzF8rpfpy
G6ouskQnPiFfGb5I4ZQQCyPUx+lFkui+stZbAvoEDYm00YvZLhPZUQzLxZcRvdkf
/X8OCR1WouTQQN5n2cj+G7q6x56v7+yZfM93LV9ps6cfAfLYrbCjCbJ2cuHzP6nO
UOV+0x43YPMbZCLhqXfkUZ6HA96ppv3iDVDLR2dNF/YoFKt5WOyew2wsekQRZ6aw
EGxZMY+bF7a03P8hVdF2SST8xDMuJaYkSAycU7xZ4mDaY+zywx9/1IvSMR5o0COy
1tzUHQOafE3Vci2Txfi9Qn9dnCfTgxVz+5vfysbeOO255t3sYjcCQFJUQtbFJzEb
XRJyvlr8dk7On8mKxq75m+OP2C6L9TMiYvPpeS0OP4+Gi05NnQ4rY7ewFKQrmePj
NErXbqL+/Ua6OI4z5nGhIawEU2josqu4iL2/aFoHuBUk5MCXJcNH4sqHsmZNNb0N
X/MyznYnrZqQpOE6+Wt+xvjTNdrHK03Lr25QPyNP8fPVm3xN0NJqsL0yFAplxfGM
7lS4XljY0W73zVLA/8cf/wa30OT7T4YqHBLKY9GjD4mYJAKy+JJrl+zb3PANL+ue
umEJRSSeVED/7com6MIQn4RnrPjNWQlVsXFYk+cLK7rkH7GFdXFfVJe1/snawYDk
ug4ALQE5Ifcsrs8+3uKeivfw70PqpzODdNtEM1v0XKoVhpjWql+cmxjOnRDskEpA
xmfssiACnQXKapgkdm3aXaOGxjc4WUbl4ObUwZ21O3JaNBpmCtjXIbPp5GhQglsI
Olcgg71hDiFVazGoKXRy+nzL4mzTfD813AW7vw3o7YXbM7t1Q1XdJde4d5kl3vcz
71KqMKdoThT2l+YBz+rtMrHgkFtzbSzKc5T7zGp5XbR25poWY38j9Mj66JONLOlR
qmeFhH8gcZadn93vad6LWyhfHDtD538yMDBIxCAUVp78d1Q80U4RgPJzPHFb5oqp
qvVvghlO07rMR8807rSPB0ruE3SJo6H8djtAgblQRZAkySHAhjKPJIgf6g95AyTM
Cl/JDeHjOZkRCRPJs4OpM3NhZ1U2DaeNmTHhUoECLrGgv7n4oM8ZLXY8CEaBni8H
GVj5+sfe7qDCxhfsv5ggvFMimPEL/gr6j9ZmAXG2TTRDpVbYxexzjYU+C+RaWsLV
F0oUz1wvWQIqDVfS4sKWVcmyZSo6poz9F4tK+FRNpD0DhvcPt4GPMd96NDT3DFM9
PTRbiroI2urbQ9cpKdhTsDnqiNe1CTpxeAuX/ARM3gCqsVD3p6eqCzE5saYcA7E1
9Py6JkU+FEE/S9eJQdU8bCaosNfbDiBLKNl/foXuxYonkAbraj+o7A8YfkUlYS78
YmmjHm3+UsrjXCHRt6xavtJPLR1binDeA/f5M6aEL54APBc91+FsuqBq4S62aoXJ
XajAGVav1SnohKy73mugPmM4W1yDE5IWKprhjiryXraHNJs0aMPPVNXk0ffRCmwH
aAtYVGO8SO7lmhSBFRqxWzjx+T3uYVEjTzto3yo6P+8SA1zVN5k08yJzbIn/Rg7z
aMqge7/11M4ngJIMGlteollIwB5B2ScyhoNyBL7903W1hZZGiyOKGX+V7z2sQmre
9xtQDqBSK+aJG4m/2TPLge7qQVLuB8gSX4Z9/3dTsKXZBz1PjQo02gXvVD8hPWLP
4xHZzfj/0Hishl8IPy7XvrIdXkH0NzoDq8dbekhDXCLfzB3ZvuNWrYQW+ZvTxFxf
kXEUNmuWh9T80aUKe8T9FPa2d4xmTRg3f/OgPkKujRuuu76+pd9Bhf2ka7oCP4jN
RQTDjpPcnnUFGEgE3x4h14xb/gQXzEo4suDCJ8wmuP34/gPTWKRhDLkbYn0HcH5V
uddr5H4Zgi8mNfNZRtb8E78cyjU+7Z3inlN3pByYxvnu4oPpQZn6PqR6bhlmKLpl
khHDtWjUDgjszMZkJrE9pj4GHFIIT6tFdHRMJHDIDApiJZ/GNTJagQBaIhZJ1w5y
KXGGVdQzb4bX1DoFk63D+6Yvo6JLzn8hNOTpWVVMx5uo1CH4H+cJ+8oVg3hQFd7V
jxQlXiW1U7idJEUFStt1LPfUJoCPtPa2TiWJ8GDgP4gJ0E1gugHyA6jlKWKXtSmX
6kKrRkpTQ8YPDiQS9cdaARZNFaAjj5q+nAjWntNvIsuV93gxFscxgnmZ0tZsL9bN
4IXrtzaYS6NJ75XHUwoCRkZ68emP6dJfi1sGJV1kXWE7mgIg64NU29pVGCFnYLfb
SjfPcblbYUEIIFZtm+ldBzK8g5VPLXMX5F+Yb+XcwTIN9OzPnFG52JTw4q8wzZC1
mz1aJzzDjoOsC0uFEoUtuBLNdQyMLJDyrbBHw7AWngEKQR2Zha5JZxgha/qmBAvd
Vbu5ODOXgLEeMC7RvQSOXN2w3SuWVvZCb1dXz/3FEYt3MT3A86IsX3BZLtlkBW5L
NktcrgKp2tL3Ftl9mYRA9NKdu9RwnlJRAYtbWtI8VTQT1pepw0M+d1pnLucYYlug
rSspeTq0N8zWWvW5XS6vhKJiTYTzddsgnnnVRZtTIGTN5FT003uJEK/hv5CQknJ6
M2tHqXyphjA4tCqRZU0pn9o0Kl/sB8P222Mm+wO993Jv24HmTtTaDBvm8VHMC0ac
jXfUtZO27PrhVoSSE4YPbiLK5zfXLnAzPJQrbxsJRHo3b1sFVb71FBj9Bv2lGRqd
lzkCu98rQQyx405AvbZCbEaP+6pseTaBdvKqTy1A+16t5jxf1V3aCT/KR7+yKF5T
Fm0gcsuozifEIhyeSx5vrofAuXzTg7K1CTKlxfCZLjHLg2CDReuwo2P7+dZO+zhJ
hqvnKqK1GU7THArzREtnSe33kRvtVsSRYsrcfu2hZU25VJ42RLFLaUsvEPbSrUJU
DVy0oElCbIzGyYJ4yj7Ut8PooSg7bY7qD+AFLVzejWGHeYuyad2RbLYeBtuXzbvi
qZ3wIJyPqi6OBfcKCVTJXKe5DXPQ1C4BcWRSqBM93Xfr3iBJfTS131CzJ6zyD7XY
VClMXoRdsTA0a9vBqvjnKaUOdNM4gOd0LfJi3AXU5mVVZT/asA38cmDhd3a22Yi5
UkRxlpBraHbpPBAS+6IiXqpixPdvZ3Qgyxaj2SFF525+ERyNy9+2gv4z/XGh7csn
E8W8gVjM9Ic8Jk9HVOIykg05QotpHwssuPiJPcUEbulS8gZuKBtcYCdhlph+QCC5
PG2OYbZDM6gtPu0rGbFk+UJExnRZlh+YGzBMIRtcz8xS4bfxiMj3JPVia5VGcjQR
evg+AdmYem4jFIbjDpzNUhZMEc/l22lAgseHiM0Rk8m2WmYPJ/rc6MV15Ynw6Uic
9tzfYO5IxPuvVwajf70a7WIzbX0633u+auC5CN/JmsbjEmBQu/vhCAdeXE7W3M8s
fhRgs9Y/Q1MQiuXbeMsOwmkaol7rpyFuZimx/qHcZKm2HUKJCwbSPI0I25rtm+OW
YCK6dOjLYnUpKOHZu2ZzXt/A3pcFrGfyuVBE2l72QRSCUe0bPLWyImbDDmgKM/y6
kSdJvPbKZHRC+oPd1g6XGYUaAm7lrynuyWO3cegjwm1GiHHT5+9wY8ecFJl+I42o
3TqwmT+1uEsQI5TQoVffxg0e2wfqtcvN+AlC02uLKWprNgcHh/0YGxZn+qK72A9e
HGhR2Q9tKdZLvFRpFQRfjQsCkVqjZTl465M2Riw5ZX9PVxzEt3Mu5OP8IA1k+i2+
byTdVw3/PM3TdQyXVUkVL8XccYivM5fjoov9GyRHsODC6dBjDqJad9iYlXYOzv1E
DE+Qz5LaR6+1QH4kdYYnWILh07kr3fAo789BcPP9bIUeW04bgbkqRGXcBPJS80mf
vta1Ef5MxQuPc3zVRRk/9/Nnxzw5zSbUI4EmOGBaaH4iDlDMP3r6CMn6HePpDrtK
M8ISiyPpal3yQjGaEY4YZ4bQPw6M1oMBE/9iwU1kV8Qgfd+ThP9WTaa3tAIMDk3f
I+4S8FsUg/09UFLtqwvjT6mi/tM6OcoC/QjPGchzOST3Mg1UxTThbTHvRpQJOo40
7d/QMKF+PTRYmCU8xi/XEdchFtE/BfIprJUFtGQTMvMJw1Mt3QrqYZ4VR9r00XRV
nVMMMWK0KYYLl2Z3/X5rYJ9v18GLz237Jp68tLOeXX2LlW6u53ABKaWmp6AO/e8r
MIXj2EP7q2DKH/1y0eX7pJwRDrnQAi47bAqCeg8uV+a8FxWMmn8In/r7xd9nwc3g
6rn6TIAJukK+tNINBP5XHMFsy9gdBj0OK7+sl4E4eIMuIJD6og1Og3RNG+ZhHkZ5
HdQMpCCi6lY7CDLG9LAKCljIe01OLjRoO3AkQNiuXh0tTmI2MgQIj2h/ja4hQiLC
cyCZjZvbP1mO+cq3GVofWsEo1U+5vzKH4qCzEHlcpcAL7lHt5P6QIRDAfTPP+BxI
Qu4JDNn48ay1AytxK2gPeaC+ux3QScoL+5RmA1KPyo+BoHjQykImwNXB5UPfjUnS
oxcVpkoEBHN9BMplj0Pa+vRN9vcGQo8LyHjfkQAZ4GmC3fs/NKV6M9cd0xhWQGj1
yhva+EBezzjD/acl/kqzsCulnQzt64LY3HJsQDolsAGFB2GXnadNf9jeVMquWif1
Q2tmSBi8EXM2my2ilDQK0/hysNk0+ofIRgKek1cpMYNGiyNmHJMNw6gEPLOn3H7A
gwIWbUyoTEVAtibBC+86F55XKLVLvaISg2MsVbej10HzbCLcLgTWSdn1lzdF1Ljp
dBx/O4Nn1MEynNszVrSTTNNwcb5lK6jyYzdzDYlPtAc1qN4RTXHaY6RBOcR7J7/S
gpnmatnLo1NF0qbSdCU+ZT6V7o0M4tfErkxCc9EWbFw9X9FFd2Bk8PLEMNFnVENY
AkTvLbGNaqiGo1YE+qXxe2nFSd/GvNUKzQHxqBNHuvlg+/Af6E4fqbffpN2txCPL
9JfN9AdpoQjhN1dr+0DreZpApYYR13GgdxUOGLilfpVPzkNa+xQei8HVblZ01SPr
TsFQerTbDGS9Vpr7sgHkKlRjOb9IgciHgGqlFpGWvk7rJAJQTWHLJbjYtKdIdW/N
X14H6POI4dp5Rskxp2cVOjkxn23tSl4O2yZtr/OAK0uefu6RPz+5aHS1VKuBgbjT
kbSqEqxyLti/SdfDzSF5BwVHRDaoKaO0TckhhKnKSyfZaB6k1q3gZIRbRguyAITG
MHKumYejB9v5DhUYlXywLBz/EtG0sAYUpB86NQi1221u3Ux6vp0tRfZSVpdaCpRY
+wIi0Q3QsyJOvmFPpOun1aRyL/7xyQrfhXXqiOAePJTqax+3paFriBlHEF1AAZp1
MOobzff3MjePQOtFhDo1jgsl6fZLVCLWH0JCzfexQJtVLMfLPgibARTC/7TYPeEY
xPhmvMo80W7HxZKjjYyaPIdthBMgt+FKqBnMnNG498xoxPQsRFNzI+Nfe92WP2Dw
ZPZtc1z5+Sk+PGPtay7Tm7VQLrhNAse8CDdMtaLjaaEVsTGIWoRx7zJMZ5n09hkQ
4AVDVcyrcjRFxat2f13jE+dI+DTPwPOCiwxBrBwE3vq+mXJnbs6xJEMQ4ys6KxiV
gsTchwQlPJsksA3VOvam9rfiw0O8vP/S6Lc/N8+2SI1MWU4fu5RQ5W9EqjZ0RpyI
tGBS1uISeT2Z2QZqiwFekwJH3ftdYFOJN2+ioQ4qV1Vte+cTgtjvOWZXsEdiemSa
KOSbM7+ezpxEILcIqiL4NbxuV2rgeZC3+pvsVjdQY5dU73EzaFUNPMRUw7iFSOgt
CnNyjq75aVoV3NoKV4QJtIsuNXGaPadeoDYzuMi40wisFQuek7u8ONGiTH79s8Mh
BYF/ezVLl1ZsdnrajKlRz8wuxDiT/BhtUH0BsHaY9yTtR/QXZMkvT6ZYLGP5Z5UZ
lXQqsnHyrHDupClbknuP74HPLctKGb8vEsLMwXWXoDl8LEYQ3QHgTrQvxDqv3uMV
THzgeDJVe0gAdp05EQjLnonhEZbYYMXFNBVjU+ZpmC2ra+ruAuztS7bMqdLsVP35
RpOXogeqUhu6eVacm3ZxOb2cc5NT7Q9upOwlhN3eR2v57q4CbJ8xmGfgo/Fa82u/
5rmtHu5J25TrcD7suNDP1derxnYAiY1msIyydFAIE4pNeJWYGYCHz/M/ojc7Kmry
bKdew6jUPoiKuwOTqsgHJEg3oVA3IIIaG/GcGm9lu0z6SWuoUZC56nnr0DijHk+k
/w2kmf6Dwd0BlYuveSD+/icBPPUiHQprc645Oxl2qurNt9Ny/wYJ/ZRmt35amfKb
lqt9hAvkI35tUth95zCdBycI6f0JgnT2elSfJcRr97cPc+oeW0igWKlb4Cev4gns
ZAJ9vDdUteNaF3qKcGHsWQdUVdOr1jgHIZcgCHzFd1zdEhfCXMGWTn3oQiEX4DHK
x8WsM4VmgTB1c6fOEVR9+Homm+RHc3tx7VPSwCjQdR6hvovgiybZcR1cdqww4xwH
C6P85OXcstieUZqa5Y+A0MKaP93xZtoLSDgcaUA5GXBlxfck+GU/CxM14/1p0giT
DjwgPZvYK+Re28JwP7qm5fUCA7QqCYLHFY85R1lxDTW2ExTihHm2rcywXRf0D7NX
o1kcFocUnVdoe/kqzN+cgywEp24lqnLoemPg4g+boIyvMz1ymQb6uqHoxE6mehV/
5Ptpkqkv974ARrRuVesEQ9IMA70Y1QsyNA8oSILFFU1ELK0XzyvfXOU2qMSS8bw0
miH1T5Za6/8zk0IRws5bGl9MTYLI0ZuYwbWfsWVV2yNVDP+1mMQ9z6llWsOy94l3
QDg2oINqi470yUqOep97vKQsK1QJnbcqaDA/G8DvzIzp1z2EoYAG1c7QKPSflSzA
JoR5vQkxJOxwcaqkz487wNAFZkh3EL8/CLAuL2FrSHo3H5TD58/bVOVgjZYp7SyN
V4QIjF9D+TnLejgXbwto9LvE2+smWpKnmZBBnGfSI0FGEp4pwXdltkCZJmtrId2l
PJBIRWq3RAOZH+yrbYtit9LUXO4wSmr2BUFleQjaYwvNJBXg7a7OqNT9f+t1vGDr
/4HMW8b6KNQgECFyu6NnBpItCIY2XqUfSBI69geP/rdWB2REhcfDx4BUKS3zF9a4
3t8tUXHLYeMSB0d6d34hk6BxCQUnqGQRgkdRcFXEsEfHE3dnw3f/QmSNgzUbmyJQ
4y4c/Xn5FRu+8k2iZLOVPhlOP+9EEUPqjEPwv7/WoVRO3iWPdlyGQAld6Jddx5XN
wz1aioPBMloR4sf2HIDiV7h6KaiF2QtiUCzqucrY180FhEekvRhGL+e1giYPhHL+
WCSJR1wFkZSEA3vxJOIDRsZxqONXoBeLQCGqrX+FXn9grlR0thTIl+jBAcwjiGJS
pA+35/HHcDO+z1pbeIRWnyYc0Hi5+1nlLGN/HnO87KasUItk1V/XXQB55dfmGApd
wH+eOsMqpeUiMxOya0XSUkIxvMqibp5Rwlq18CvFMyAazs1Brpp2q6ZMG2UmuuEE
CSlTKDkFHQ2/6ulZO0bDyH/bgUloUm3WF2uAluCgVvmCymbWcFjsnCLtoNLqvTmg
GbFDHvVcC3IOATOnJdkip4mTbRjHmTlTY9irdJcTbYhF/5uLtrTupC8GHS1KVjHS
cOTMytvWcMg6QsRVXLwplIHWWI/nPpsdSfSM1BZ4s6jq1O6dz3DCnSvrUjzDp7Wu
AcJHjDPjHnuC0A9Z7+mOjAFhf7K/Qw2bAdsaROdwuxcAI632qVm07fN4tHNynJFd
K/ltmGVt8C1P5Tppq05L1zbswVsO+YOOPbrDaf8MBI+Y5GUg04OPBOmL74SpXdE4
vhtfFeO6Sy5rYNlGdvn40+0dvAQ3Dlt7/zf5njrYvAwnXErVokEFrXEp1faKBHKi
KDO1+L83JPDGnHoxebHqLM+CvZ0WvUuBJK7n4SYCSo8Q8wcSHAQKJCdi0xFopPJJ
syql5lyRtrAtZ6LDMXtS+7YZaw1jdjK8VHMgOFO6btWnKz6DvsTqZbL3ZP2XblfA
b/vpVcXPbvmkMWseugcO8Z+SO80Yqq5hhiohZK/1PP1RSgRsX/38L4zrRfZpi9R5
72ABZBF7QxBu6VDZzFxJKwLRCXIdypBHFu146TVDw5F2v2imCjHcBPTpDC5ZhvB4
cajmiExoUpjC2dKqJDP7UotmSj2p0c2WGOyAKIrfhwfJmFc3tIIWG6o0ril1cga4
r4oEpUFS2Io7Yii1vIOlsBfhbh0CWPWydbi1hfxbj3KI1+x0zyCErV9eahqQPpmB
sbDSeam7r2MpJqaGt63FxnAGf/y4BZ0iCQzEfu10Z5kPv+4ks9CpLwC2O3Y5S4Qt
5iVxPInqw5Gh5vU5A+o5PGDJ+K63bqoPnbIHc4K886RTYb2iF4AMe2senzOSy5GG
V0/cYM1xuxYFKAljd938+eppJ8yPlQWmhEwxOxlTuanzfHU4aamqn3jNDYyDLGNI
d58JPOfG/msl3hIxFBvsy27pfsKiVjXt1oV/+gIk0SQZsBBjPc9NXP5ZfygVwvDG
rWqwPGH2YgmPZlSEDSh1r02xv41NuslWPuSpNFeSo3Iqb+LZx3rE00qeAXGgl0gk
5+VAdrtgRFpXo7420YInhwM9JBtYHvrlaRJorhrfeELdtkm15wAE7vqkvoSZ/wOB
0EOeWNpaf5BjfcXgVjKVr3pyREIkfRKXJ8VeYXXscn/1PzUKprDRDae4rQvHQeHU
bF+4y7RVNP2y5r22uTtjEUpUc9wFAcfwq2R28ooLXbvJYBnv9HGX63YJahTK7q6w
v2/fPLz1Q65k039kjQliv4shxastRyokOXsnez/CvLHOeIVQun/mf5y1blTFzoqZ
vLqvo06UdmZ5HvUOU53XYB5b7NZyc9vWn2A1eRo2rYzOal/sgM7BhJve3Gj8vFyd
7YmYIFg4qJQ7w81EhHt53kLp9vbOZ9Ld0drxYr5LG0q4S+yXGE0XGg0MPpqWVWHQ
0Ude3Vdd0LjC5KbJs7s5pykGgmM5gOPeMx9VhIW/N4PsWY2ql+y05zPDauY+oB/q
l1avhjU8/QnWEfSjOhs7rum7hD1++qnR4fSbeOcH9DWf5GGCuk/XWMhTRAgMIJ4S
KdOWDYXtByXrGjvkht1ozIzwm96mQYrZG2amvNu7YmdeixkCvhxemnz2qqzpd0YO
BIhKXo8rz+gvwxBVD58QmVDW179EEWLDUtOIwjHhJDD+ZJ0tq+reIeDVlcWSkGHB
U5+go/75mG72o19Co8OTINvibbvZECHG4XwuElf0yV2cYAOqhY39+HHoYcjzenjA
HnbRjRotQmR+bKts01wL1+Xwney21gr2KDM7ylKiTQ83xCcu5NBeTwpF7dwKle3J
5yy5StUJEFgqep8ksI8Kcyz072BN8/j1tavejk6tr2eQijg+QNriEGooP5ulM0bQ
fNywyKalks6XA/sRd8dHC4Ymu5Wu6miXeZ41+CoHbT1owVLDCp5wss5Jqa5QSWhC
2VSRDJu+21epuL/nYVDf2uo/q3/lzsmlWDSIBo9K4cmiqPasjsHbcD3YfclFCdiD
C98inqcyQ8fegZFeE4AF+p+GJUZWeu38d9TmalFf9y30LAkB9CSQacdW3qmpvcUa
veZlvqjXWKVgvN0J4WpfzbOpZiCAIfviG6VdjN+Zk/lN+ab6rBI1Sb+CjYonExri
dgneD3z11TxvvJoISyQvg1ztvuI2EjUfVEi5Fugq+mCr9rXJRcWoG5XGt9C4lMMJ
BrDQ8YpyQSLkIVAesVnzYbI/uiryVhR1sMYqdMFq/kFm7cNqTbgkzASBCb6LEMjR
WKu8lRG4NHy7r8WSD1mTfkhz0sWV/mzELcEHxfFAvU6dlHWlqY5r6N6Kd61s2BrL
xydgh6+sO1jzZaYpsyGy9trMbSNKLnM/tTD4hbwY+wxm33JJJecwYcaZGPW8S79i
5Rt7A+dvYHn48QzQSWGFFvqQDTv/pn5W1zGRQ4VNf1r5oZHT19qmZ7rwaiT8q6Kd
yFkUZABPhQUTBqXF9nfCjdDkAVxR0tak82piIllIpSos0tCzcbq3TX8+MfiOU7WR
9RrRw0AkHkBurd7KeCuUvYMgN2R80bMKQzsGNihN/ahOHpxeCyrfnRfKp/NXjHik
5WAmLybCl+ckdvRAcwYUTvnC7QaPxXZUbVE5kdwGbIbDO9mt2lLlaNJkh3Pk5aNa
wLl0j9gg7Ukbdenr6WazJQh1Tkig2NSWYYOc1K/FSLbAcfTscrcEz2ZKcJJLy7UQ
m7nLQl6+Dqo/bjreKKXbHsIpGQSpphiy0zfKJYu5n8HC6FmnqxzLrJYBWk6iEgag
9pbjNfAXfxyXscUMpJ4Hst7wqsonKlXux7IAnTWjpX2vfKEcFXhobbFf8gsexOg1
dzwxC7005Ow1KtgsdTUGyDuNAB07/V54lL0YBwKzOhGKJsHX9T6men25HBHRljAg
QkjTrfgQRw4ofmxPeidFl/CDfHXGWuK7kx8J9tOlczwHff8BWjGN560S7pY44EFe
nsiWTz5FXXHFt4WRrSqRlUDZ/v9TdqbeYHTxbUs8MzVC1KmB4aymvRsVPz9OalPw
vMZg4uZq2Btw589gW4HeAPuMhGzNP48vDXA/R4q6Y18/L9oXFM0wAA2+n9rfLBE+
v0sWiGVzB8mJj6SpUFTk5/Yj9iPPMS5SkLScQlavfl2CtYR8rMRK2Wa8IyxEM7v5
dDLzyjCqSAbbe0ACc4YGJYe+EZ3U5G/0j2J3gZgsbVtUtPhOmjEJTbQoj73+C0Ks
xth+xxNSj2fh6Uq29YG4wH7dFBipHIgwbwIXKHuac2i4LRwpSoNp9PMmOwwFUMwP
d5j06mLEmwuv8qJ2x6h752E5z+EXQGC9nm5EmPs16FklXFel7lyqax3XhX9Py9qq
Tx40AzXNFzyXgX2BGP8PoOL2hkXW9QBi3zmAHXYOgFSJn1lbzxIvfV1e88uqu3+2
ubtVO7SJtsn4Fs+5nqa7aSLQKU+aPpY9mEj+EwX/A1q9ZY00pNpiIMuKbRXSagvs
KC8d3gdBpipz8z6lykAshGgYpnzeF3khvXMOhhlo9BMCTXqPqbi0mrSQcVe7Rqyu
v0HrLkS/UgakU8m4J+Z5s2rd84RqjxowZHFU2WAVr9vE9GAId54nDtyoANhI4kKy
NHiVofbZHLHf1wynszZR3t5tVoG3CoZMyg7o9Co/YOrD7sgHXeogOqNXlkMUkeiL
oJLAiTE/9bvXu8bW+7PJkSiPcPYZUyGrew9i7tKdtavF10mcpDk9L+4EWvcqQA7z
IGx38hv1rq1sKWK7gUPe7UTiImSNaipG462yvELCoiQ3Ort1ntMeJgCthToPGlIX
N3D6l5WGYvPE0UwrRjrc4hrAyA2kMQYKCjBghQJqpaqC1V0gAcF0P7RDyd7Xjluq
uDpklFu2ogQilQr6QsL/zcIl62R5uvI27mHRE2ucqmDghtPwTO7i2Fc3ER75picC
gry5gjswL9/XQEAbpHMbLu6HCJZxoJgp6vRqL+A2dk3uJ/tXuzi9fwTdoR+8dBxM
01gPmCPNG/8hvY5X2U+JuUOUFM7DTscTraKJ+4qBHWgQb766DrF+zylswSK1SInI
zJr1/nhDR3Cr+YJw/xt2/gITF0d3LxXRcul2Aj59ExmMdODmg4thpP+6kMmvnEfX
ULnPV+Y/3xvVr1zMlh6mZE6HSU/q3UHrbBHIljQu2yGZLTjXMjxRXrGC+WqzR2Qr
GZl7hFMco1gdeAbQFl3YP9VlGjE1KjI5GlSsYSfpMULvqwPtbSRQQKlTvHb4WHna
TowOnpo8yIvsK7SLuRkVNoIlyNYbTaNDdit9KZEZSNYs3nmecdxAPJ3+ekX7bCIe
1gGsyHlzOBdJnR24CULMvbj/GDr7xefGmIzOF6VPjcAmoVEezz3B82vMatM8rED7
h3C7ZdHhc33jcO4SfBYunCcBlB3uDkWxHm9l3GdmsMIBYKAfIxJLayCpxRDd3Dra
n1RCxW3E3zLBsQOOifJYt40KBxOYKlJvVldYyiBAIDmamXphGsT92HQCutcdaAr4
X83N9qIDpBMkmSxk3Q0TTnx5M/wQ7sJzxBBlG5czWi4qfGdxJJB8cB5HSD+Z/mja
nmRnYzGDvbL4MxJNXbEB7XRuRj5dZBRI1cDwb5T4Ee9PEAYZ4XRaUpFYk0qDAH0n
DquD8RZc3x16bwxGgRa/RwbwWov/PeEgxAgtGowViBknD0R2XqnxN7N/Aj/vz5NT
3ynUoo/0lyKtVr+2d5SDjwxhnG15nSa6CtCmxNZXHx2qiDaihu+Gr2mQqYu2D/yl
YjZTZAotAGTe0KnEqFVSmT8Fu3wP2S1O+m62h6gHV/ZjUWkKnd0KXwm56sF1oxoh
gd4tRrrygn6kSU2/qoo1dFczYPltRqRRJci2iHduwE7PQVY4j3uhhbYhwzC62cgT
Lj0GbGUobAN/Q5ix5W1d3uPExlNFVSMOyzADzngAz9ERVPEZXFEXjIgqGFsbIEH2
ki4wjoFg1pyX06+vkDtOVsVIwTnAiKX4TISCh4Ir607i+Nh7MVSb3jRHQanx7Iyf
7ejPj40EGhH60TZKMMBA26rZVTS+MoFkxPLRdrqD+O8aQJ251FkqSGk2+hzjLsHO
nNj0IJmbR/AgZjHaPtyi0V66Cau4XNlJKfNC2c/kMQpGC+s65xbBl6sBhHdjBFZw
uZevIG9qdQlpuXXj/jVQfXtkd3UYhTsbvU/9C+TiTbvJu4KMu2tLa/8sEacYgwfY
tcGrehvR+ns2rhqhUwMAu0Gq/tSvYgB0+Zbb5KVZJdCHDy0DgETeiLmSzEpwCtsS
IJHBtnBqYLzpga/3d3g8kPzgYWUrIsFB9Kci1EHSRzhXYjFLCwGxuJd6Yl0/jFFL
NFDoE7XF+cN55kLjouV1pKJc+MLY6pBUm57LGN1I6Xh2g7DrSgU6LIh9uC0Khx9w
obXXVEMi0exWseYJSowMLg8YgCb2nr0uD5CPy/Oxin4MTGFDJlj/WYKp5HhzaD4T
7Pc2eg6pEaOEZkNvAR1wJy9tO9PGuVSTdDIoLOo7EqT8nyAMXNRl5yq+VMBAlLfg
ZOBnI0/C3kkSEVgWQTegw6ujshEa4f4eT5NXvnWk3QN3Nib8s9MeBVrW02W8UnEa
5vtYrE36vupDDhGgu03rJM/6HdS3qe/KGn7i0m0jdQihBfAKKCruS+L4emhmOFfv
aP4vee1Xh1v/qIsT8EgQovDn0aKJ4xgvg22Fs/KwHUp3U6LQPBtkrjW6JYEtQkT1
RXmGH24EQTe4+jRdQ8HNcsyDAVUcfu8/LDADUv3agyGSBNiDwcsjP9FH0q0eqeUM
ainydqEsS+ngtfbqCWqtuL18GNpB2vsrznREQotpxFAOO2THLZ6G2g7U06mTAObG
EllQQZmeBneHgsdQUjPpkM/9A17JvD1nUNJ2lK3lPEa6YGNMBvHNenJY4V0JI4xo
SjzBXAW4bK93HsH0droCHqBpqlNuIsrs4kUrxETJVhdmexwK1Pgnw+HKDxZqN5Er
t5MCVPHMHJuiYX4LRO4zLpktlQknPkrDhX+KUgjry/17LXAzm1GZjVLc1wcm5tD5
qvhc/GI86OO2hq510afRaxIOzOXPlM6G/Ru71XIwBJir8hNiNpPQQMCToOrL46Fo
xgBgw0eDmFoqNBB/5OpZFKgygvAXOH+R+LBSpglzmqQ3eWsrVyh8SVCm9Mb/Eshv
IOguKkEcWine95e+zzra+OZzIJt6Dur8f5h0Um4GsqyF/GoTSHOche4YjaPP43Oi
dRdlSlbGpKxoqHllvIVyYoD74fCQCQ5jlqbitC5AmO2RT99/6MMyDsf2a/p+kcP4
BkhGVXXI/0pUgdrVfhzvs4enqPajb/vTU4aveCDc025YcApTwcRXAczC4Zx5aBg+
I5KnO6mJ3M9Ye8c6iRyyv2enFOPS3NGdBMd4LxNmXqwQ+YI+/x2Q1xHrUUusoLH7
RKOIk6G9y1c1c8K3LwFg6Hdqtq4eM3ffaaWV1YdV8pmF2AuUPnufGUgzAnHRomIg
VLTYrmb/Ci+GdsvTuURSGc+qg0beTqgcAmKTt+tN5UTP+NPECZJSgqDfRXhn0O9s
CqnMEsHVCh/lxxUmts2BUHujCVu212TRQkFxqJalLdDanMExWUTbmkVHflqPyspz
Kpo3LdUR2V0ZGfut8/GtuyWDz5FZ9smqfFvP7y1ArPNCOHtb4ILBZhq6ufPtg78E
p8MdmHdd6e/Fp5YJ+G5ZaXpjjwFU52V/hK7/nZRrTzdtlCtBm8KJ5esQmAL94vKo
EjtXcXCAZXb9HgsgE+yeIVYpvSWgwVgGKDcZESIo5UA73kCcPyfDLQE1P4WPD7QV
ez3uSg0i9Qlo/DVmVIXLMxnceL+T/4kdkcJf/YVdrzN6tA7Qu8m4Tq7FuQXmmCNr
u68migzcWOxvfMP9bFwjFPK6d7FfxuCxEhniQf2VB2xkc5C5mYHOZn6ephfLOrmB
TAFHFcq8VwDquatyD5dxWCdO/OGS55kZma678TLGJGLVygqDaV1cp6NpgwL7e3LJ
kgSWwGOnfl2tLMdNm/OhHna+lvqYq87qeyU5yeDUSJys79JqSYfOK9v/N9eVWs53
DfrNVsWRXGjQIlRKKnpDd75RIlOsSPEPuTK5oDfdaziLIOLRe05RduvThNozFYnJ
V3VqwHWNM5Fc9szWMGGqPe970+/Cy1CeQkSv/G3kihi3t0MGnGtYvvVyH8tROLET
45dconJaY9yPdugkPsEuNIMv2TlVZ9MfOoMjGtAAHKPPMOvmlbTeHm/AEeuCQcfx
B3ASU4o+Cpu7Mn60ngLOST3+5TFmECscFb43pvdO2F1XHpwz72i7N8B3S8qgLnxj
r2593FoieR+9LxYzlTYoezUlhD/2803BaYhay8ZUwusLE+HWDcQIBP0OO8cNun2K
iW5IxTB7ucgustTNEdVbarlVAszIEzEQwg/nnOdrPFnWmCk1UuDvNCHkozm+SWqj
ON70SY5oduim33W6VwW+NazP7kjYktnNgvormZ26bRdDo1uqezH30EyNmxvNNEJ5
N0u/ZoAzQiSkhyHUMezFwLVyZ+BMhFnFl3BUtRDy6rtFmWcgMaWUyVDtzZq//hqe
TWMHbO8e45iYH+jOn9CkEW66xFzKMMnC2foSyoMmQWbNm2C3cLQAmgBYJZfr5om5
3K0bd1Rl+JvAawCVR12nu/F4lzzANKPVkvJvGA6y+9POhvDv0W+fE0kUz6LG0xpU
nLp96ghRqGdqpdO2Z+aLrI9DkiwnV1C53Pc7S6sVjZy1Q69JGAQsd9soArLv/79X
6mzDqXJXiQEUgcJbaQq9Y0x3ex6UNQ9mmJ8xuD1GwJtjM9zlJAUQDcyFsGGTt+o+
guFqKkAH2jHQOfBsKnjf9aum1mK3uPMwjUIyPR6cYbebeh4bcqJyv9eQWi/QVz8U
c/JOBowTLQJqVb11z18V3cjCz/8A3zOQ2X+87AlxFnKXEp8O3oRk71K0rS0l2pet
DmiTndT3O0FqtP9nUk0Bn82KnsurgAUFUKU2kSHtn9J66DkRW6J76Nrn2zJsQMoe
MUgk4gILZrV3xX7zg5vyNTeZO2GMvlntuO4TcRRNw0XApKX9/Ar06E9wecZU+i0G
+ffznmYsBXtwMboidlKsIZow32Ipr2AtpKTazJ6dYdbrFND9KjVORZ081+BGEnw/
cabFRiJ6g1dVozXIlu7wKyDqH/ZpkDHLotKahig8Z/oAW6LFDZnb9Jih90ji+k9L
mxsJOiSCUXImr6baXzKd/oX8EDiRZT/F5i+rafMHjrEPiDNBlS+0vLTO2CceRxDT
n4DhTq4X7jCfMFghq70gqzAkWpIDYGNldVQjCsrmmAJ40lrlcx8Vf5A6nDbwZj4z
NRo/WzPEyiwrykDuj1PZfujFKwkgWkqp35/LkfX2HXUF8rwnvZuafjwcvyqXVdSu
UQLQOxGhWqUpn5kCo4oPa8XZNHD2ichZxY3XmvZSA3WtkeFFPonPRyBspeVBP8F9
nR/jI9aQ8vv/CjGwkDcjH4v18p9xGg2/nFrxWNdrC7Il58WfXCI0kkBbDIxtq0OL
Q7DYpoAHRar6GUHc1vysF5xaDOSwuPI8mhfJGkScdedF+tVlx51x0QJsOgUBBzbY
5p6mGgFcS+Lsf8uqkb/vB6i5tUa09Ryu3avO3RmwLJjjKyJu1KO8ve98gMtxC5vB
BvqtvsRMRLVRhQEsq+9ad0NNjbA8e2XrHkJR99od2wqHPxCLfO3p5hy8yKjphUmi
nsUN4DE6KXefC4TmwF+Ujujg2wvYiI1wGfhvhtSDo+Fay9HCptNYNORq3LI9YBax
mFuFaW/txnD6vFCLuGm3Mkjgenzeb7/y6S5Ti1/tspEddG4TckyMAxxVsmacfKvh
SdrEvHV4ySVCbXcPN1fp6tdP72JoqzZLS6JN5hGsa6HDwctOScCRYeSG837NxkN1
p9uw9b/VaJFuu2pbOMFI2s0lmpP1k+SlMnIJw/OatcTFDw2r0wzpiost8teIs96e
4Exl8HLBJbaB0AyeurPdxNlPKu3uxUYjIo+0aoieqFiJer4OaDTfKEB5muLNt237
2AIcZngo203m7mVUX2c7yfVraXqYhC6z01PzZPmc4jqKrLq/YoThbIRLzi3r9SC9
YmA0sAMYXhxf/g6KGEFQLMfu+ZM+fa8fPcJ9YZLI6eYvXkx2bTwVPREyJyDj7Gdu
NhhvccPfVl9xVF6ChVhK5x2WP1/HYaj4eZOYmu5Q9SseEb1/bVDOA7VLpgXKBwL1
JmjCnDfa0karisRfYxhIEARr7cvU3ShcSbXO+5YS96Q6nPqTeFevveOvqAHkR0nm
XvFjAyqt0zLnoas+YY3tyae46fa44h7WsF0ukdq30XYZ3009mXhdGVyO6F0gPuER
t5O2mlm5mSen1Ad9MiyLTg6FqZqpV01dSPF1dC59rKmMcojy0gsUZbqr+hYl/GvA
Lmd/zGvAh0JcxaEsmtWb9TqUm+rKacFL7k9dFi/PWzQGc9bJdcevw+EjP3617Aab
mVeuNoFThbQZjVWdZ+rW6UdoSKaAWGuzvq5ckcvNFK3IlhESmH0z5b1iJYTrGRMZ
Z2PIHGX6Ln3TkQO9317dQ2FZ01zpBALXS2QY7NPipzL2ZZ86O2VI/H9x2vKj/p5+
AN6jtuv4i39qddSPwH0SHkEzl763oUC1CZivuvz0nTXnDyv8sgMWaxCKAhD3sivB
jaCEYbQ/GhdMKoGlxhI1SQ1vlfc2olFmjG+6IIUKLuVGsXpb2JxeQrBpQ9edXjrP
5bMuSSs3L0I6dIMyIVfCxHjEYNpjNz8V786h1AH4pOUFdwGdcgYhShkgeAsk2lt9
ZIRT07Z0D1mGIlzT7uBFVoVlFEmXSKA2lVKB/QEwnP5GTpAm4Cqvu9IN9XbumBZX
+GmVO3gLhGEQgsVdic/fNOeJ44mI5NiJuvihkOgSkPpzx4yHYME6pGrk5qXhifxz
yBTPnBsjqUOyHWjeGaCvtrV4BnUG1JpOTFOVxs1Opff4KTR6JevydPTYm9IuuBiz
QYu6htGZxCAmTaFSvLseDdq5SHX36CPVds1A8cqbmIj7QMCIEjfmeb1twy9F5WyJ
tTLWKxswI2MwicE3FAP3PvxDuTt2LI7g4m6YCWgH9XZWhrLWpK5KnUT4pkhY+eP1
iP4Iv9RHuCqZ5Pa4kfs3sy1OiLZMlt/9PtFGsiaMA3hKVlD16LWML46Ou43G/SOu
W9khdy7nxVaxos2HqQ5YbLyWISCpDHLFBTYKUkJ+tUlX6PuThgAa9Ho2r3wE9M2J
XGjCErl+1zWZTugzM8o0OoNbNc+E/bRo2exZU4Oj9bCL4rlkpeUfGD+s3+KA+qV/
c3GeEp6ocUsc0BXfv5ksZSDgYH6jbyqKrFQZB12vQEvhhDjV+h8eGnLFIPaxDomd
vOuzp82bmpbIOtVjYmWxTaO/FbBzMCoOK2KRD0gpWw1qkxJVa5k8BWQb6FhmjzmI
pebxnSIsichCmAKG1FYeWA0XBfcLzDT7VaWnjoOCsG7IRZNjez7XVVoBoGx+gk9K
j6ZQ3xUPBFcUOVsIUsQ+4Ze0lKAF59zSOAl1cBupV54yjToNkGrwdUEyFauqj8FN
HPaQdG4XuhlUydfcJO3BYbEqz5KdlYgTfSJudeIT+Vv2Yc2632v12cSxBDuqTzrT
RBSI0jxwBKC3VhCtRTK+C4KuIR6wwf/KmPjUKjITktBJlXomYftnb7Dv2Ie+HrVi
4ybdm8XwuQVya6wf+uTb+o4IKScN2s0ou0OfJqWtsbslO0Ye+C6Oa0VEI5ahDLuL
AmI/CpVckIFBYSx+A8aMOtzbD1LyOz1nQlR5+EdaPwmVrv03NvQVTyyUHYlm+Jv/
mPoQkhi/KMaxAGweosaXOObf9iEOBgg1ATKzrm+K++xA6glhtAlIVQf2Rz8KBTDk
6kXiUojlQ0WDaVx1TPRRZNWKJlJWuQNMzQUzQsDuCrwQ+t9qMDRl2dZ+hpRcdoWN
mfneCtnraiTBetnnX3TM6ihJX1cb9e/Z/bCWZqg6RbGNBJ6kZIld89+4jNswofgX
pFmbqorwqq5PWbEcvdJ2xFKx8s11oT2gFjAwwqNqPxnJixZe3dpdoQG86jpPKZCW
Ya25jKydRYlgrXAXuYX5VHX3eQF0Yr8rdAdEdIujufhNWq4P5crCiAFO6t5ZEt7B
f2SlraYJfoE+LK4eIT8zPpCR8xI5Qom/tXg51/HL5rr/jADnoA5if8zMG2T1wNwz
bmW5dR8ttSxulzSSQtRm7NUYJVsAlVlgP0I3L4Ft0DFDPqxXpHSv7Gypf9IaAthD
qObFgTIrh55XLlX/azXXlmvbW8T/hounKP+pn76zF7MH8gye0eleGeQxRB1b/2Tf
MhmvQETon97dWdKByJtKPID0dFJ6OEoYkjnMudZOL+eEOAUjnV+4CETxmKkfRTHW
1DazvhNXtjAr5OwTdgsYICFI4RIcNS45xhd3Ft9ipmSPvHyd8nxv1rGGSd8GVooN
OCjed2l+DNsZTaT6yqn4AxCmhdU6zHbEVbgo7fS97XKwzO/yFCDILBdnmWJAPfI0
xzMic09cuD1pQEHlG0Mr3bCh8sY6vhenyuhWzPA8ESuqlU9I3aKm45iKfOcjHm+z
/POCP6ISW38igf5QgXFXUhUEXAqRNznUxA5ii6parXw+2KRqoZ+w0U/e5Az5bWAf
GozwItzEPV6T7gdKVBc7Ha7CqaFIqg8CRELutVigGYYvTxTv70II+/+RlUOo95h9
y1xS8s9LAQQ6F13O6IZ4rBKUD+8zzSet9fZnsfBpCYJrdjhCVQ0RXqRnq8l46rHA
B+jwXWcXiAwUIDCWfUndakHi5AumGHcmRxLgd9NryEuRN2EoPTCqHVpL0p25zKJV
ob9aivTjqnNycZmf8SuB52HTFhaXvEL/vIetKu3EreHZWCwExNwetD79+Gmh43+B
UO2AeNbKOFPiguZw/6Av5Kq6ujeI1GraSCkTdcE0K/StpcOzqTFiw8Q1ZwnldwDM
JmJzYk8J9uCz3g9CWoqTtZ6eeOqWYqxy00Ar2mqwpyfwxreWxDDHJuOmiOIieNM8
2g/2/kKUpZCB4VtnQFC/8MQNrafbPzg24WtbUAxy4pbvEhQe/4nxxmPqVN+hTIsB
4ZuY5mtKif+zXASzjo2sfQdErWt0Pq46i2ORTGOqr+YlMbi6HHiiAj0uWDXUo7tl
NM5NfV++KCk/TWbGAb2vwPe470yQYMH6UPhiSXPhx3BpEurCXFqKDulf2B1wRSmA
90c9qBxje+7Yvb5u/KjSzhARYvQLHDGcWG4YNQxp/kOzlc+7QZuAqxCMggDr7CkL
c53q3BtQHBo/3mNEWHvrHHmcUj0k6toe/CB4Z/cZ6Jn4XSimmVC/hrT56fUKWOqJ
MNCGK4D/W5jbA/+9PMUiiIUnb+g9rZQsjwAvE1fChgOiudnA+87G5etbx8VJmMh9
m6rIAvnfwdEbx6XwVafm2C+p5VLzKEVEqi4sxI/QwSiFqIy4Qgrc8470u2jtFnZu
uiRfG9IkflXeyYCxglhfoga3errqbA454orvm2OaGLW5rM2JjVBe0JNFxskmjGZj
tf3bhYYKslkOtk7lq9Ie+ksnafXkSencTI6/gbyNXD5oC60PA6JyyN0w0pAbcn/D
o94Qm9/zLzmFwQoUCNoqjBAl8fZh9U8tF+T8VqnBUcNfHjZHTxhBltPWUuQhRYKu
JsYPjHf6DycC2w7l8njgA4psxdImbw6mendeUPFTCifX+uEaMhO894gF2c2Fue06
p0dfljoJzUrcVEsdd2oLFQMNgGKyftN8X0ExyLXC2mzwlunL2//uVnUsb5VhAlh5
mGj7EvRvVRUizcUwU9rWiR/N+fsTm4l70qOMhGbWjjrzASX8qGvzIl4ej88zAgvA
MFfTsA+yntPU9sTe/iAtxYutClTicvTi9L2xy2DCdCR2GnQyyMtHbffTx+UfCfI+
UHuT5q3GxmBBU7lm5L+Yuo5wYpFY+HEmL959PPLlwE1Znxy6h/CC2Q0eF017DoCt
oH1J5LdYUgJVxWxSqHOAUuOQNZ5xEmNQCWXXH1N1uEnQ0dP2SZOWsuiClZqtVUAp
e8vjt9D4XoCz2znVHYYTQ94T9/CbWQbADSlbHCtiTAhf3kYTk1POP3IaEcLyjyre
AXbiGz21DwY+I7JTrhugyjeK6JhHbci2DfFzWZ+p69PkNrocm43bk2wDskBB4wS5
H1TK3VBYjDtwWBjGUJUfR4cSWCoS6Ci8UoQyslUMYbOgb50FQZSeNA93vL12MTlH
VtXm/Opba3BspXv2l4Y3qZ4xaiIzDqMUUI8qefXARDf4G8Y8m9AxxbYuffWqKNl8
nkT0AUVhTCtbKV/2E6FHHnsMMUksXRXvqKbgZ8PcHvWEycVycKw31+dbNLp49MZx
f7uVVHkCUv14Xl3HG5VwzAn9DVOxgd/O5E9FYAqYi8rKm+wrLBOnhiG0KRZTm3BN
Aq1UO1siNWNx/0rgp6sOvvexG8PtiENV3YyBykfPiqhviSCMj8pZcFf8jm9WWUvC
UJA14Pg7jYflyfbOL/+gij3zs+0c/toXSlRHfTipfugkq+ujWgbITSCMnQFHkRp8
62gHU7Ajs2ApMXCEskBcu8DMpVyUrMUo1CakT+hUbLGQ4mFnaiS4BnkhSyD4TZw7
IYm4Bp4Xx5s3hT/GK6hBmzXbT2PgBx+2+ryPpSN93Shs5IHftmlCH55O7EiEPkkP
LT/SSwsm/T69Ex5o6+7hud4LMnvSMSQsTmuqHTATJ/Z1m8K4KxVEx1hyRTqnfXhm
9JME8lZLc+Zd7HUzEk1gJwO0QLbK7eQfjp+icOYY8uiyrOEtfsaaMRaizvFGpYuo
ETBJD80P1dXoSzHQQ9CI7ykMx5So9GnGjlSmPUIMcnOgeUvhzXwUKzftva0uBNml
5LPUG+Q68nSPqxXOScbuL5GerZl9F81uAb3CXJA2aK9FYLFlUAygmSiHM50JUSuK
ReUdCLzx17dNO6FG5BV5FkMZSJ8JS8TDoqxYFY/fOU8WNTDQO792hCnO23d1cHdF
OvwbZ1U9GWhB3ZXIPCrfyg45JXz+zKDSayAgDfIQay1w2VxNg3g0j+vIqCCLQVXX
nw7D3LqJD3KjU5/vBjVO44kVUzjYQhgiiRcuDVmvVfOiAOrpqkdW6sYq0k8cy0wO
D9iwPHwTn/F+4LeAedHhn1mrazDlXwyt1ZDHcrvjuIiWWkZWUE3UCAjkZnQD5gKi
RQj8oEB0YVdqaEFYQ1DtJdVCZDdlGT36BpkNhhBzWDef6xykNMah0NZz8EpFdJFm
VTsxQuB7B1uqdfZgZpyHvvUl+clm1Wv6150L1Gk7lbAbr4OJk5M/RmWLt0RFoXlV
7b6NIIQxyIbOLEh62kSupzToa9HENfwkIPs02GpdWt8+ah+RS/7bnua244qU7iwU
G73pPjTzqHYYtiszNGqWcIfH8uT5tTa86tTCqTaYHpT466eesLBjx6glCv8xc1Rn
QzpkngoQ9imI2lg3887KIUc0sAAkUGYP5KrHQMP1eEEzTY8XfkndG5e2RwOF9d8j
ACdkVddx3l3TPo9npUR7TFpdZz2xKnSveQB/iWsB83tpAaMOFpaV83gA2I4kqB6F
iRqIuo91XwW9dVX4WI0y3/OnF96BjNO7Sdd4TQ4LKJ+eSMte9s0YmEsX1ux0ilM/
vfHGIHKmIDHy9cmRFhoUNwAO4rwb+0q6eiVYDeYA9196iaX16MlUIpl7khdR5mq3
Qf7c5luTclkFaYda7UYfpDX5RMdCt0L0z6VCEWQxDTUbjjNJfbOn8i9wbgYvZVpQ
Grf0TaRW1JwTqzbRgFctmQPi4Wdv+untkL6pJJ8/u+e56WEorGrjhys8L14X+AdT
/qLRSMNzgI76jCHyEOQ46NwbseUH/j+H+qlavVKnw1MVrAbL820Bw5MtL0codttf
cSeKYAY+Mf/QHBgxJRo+d13tZRm8RO71VDSJZVc0HAGHsVlTsr49WFA62eyh4VzA
Rhn66Qnc85Sn4oeiDvYpFZW9i8SH/xxmat8s5KOPKkGU+92va1Ts+EMiwoY+C8ob
zrLJyu4/PYGg21L1wheKXPAXrNhBkm2c40emxMlBEwSsKj2pCd5phPgHtL2y/nz/
+SGuGxshRTPyVnJCz2peq0zYKtIFKmMxetMjTDzq6fFq1V8kUDEiuOnvO3y3VnP2
MnYu1pO8d9bQm2gDds2MZ4weunUOYdclo6/1maHgjgtZ7qKiqrb80HlcGoY4CcSK
QizabaGI+rd7RAzSCipVwIAVRCsRGwJdqJa1ADpUgjy5x/Gb9lMS68U2nXAq95so
FVHR59EO8Hv11+gRzZ3VEVzGzYzgTORe9fGJ7gsVEWTq2/QbtlVLf5i8+wBBIjbv
4U07r60qqqLHVkwtgIAQ77UuTguMML3o5xJqpebLvzy0DVRUquComwIKcfszTT3c
i+s6tuHv5jirqNKQ1lj33w0PgUTNipKyw3Z0i1bD7B3UrqGoToGXDUOa0Mmmwy0o
VNVpV3uWdF2FrzuadgTOjuCDLc/fkQSMNsfMvdBVcmqtVtQJXgG8nHDG2V/YUjQj
xNWVO/HYNt9MtnDQSbEDDRBmMgFEJSfIsB55XFGDCNCa5BlZm90N9NmkQoHpWASs
A3q2EgcdOmY5LxxGsFGRKyOZIPQeMQ4XBFf88mgvjtqOJLQHAY4Bq2MoJAZbKI40
DK1Fo2cDCJQQ/B9c376J+pVnOMEsC7YNsaja6TeInghrjODJYsfk2a2pza5DYAek
S6o7cJt/175BQZ71xOIAdg0tWwuCwtml1tlD2naOSfcvmTEWEp541q+RbkkqBtPN
Qo6Blb9L+O1R//JWiPD+g3OQpHyx1dx3GL62peM5WF/S77tzYLy2cAk5vU1QWdJ3
B9iaipaJOqAtDn5cluEWzWE9TEG81UJQrdQOSGQBhNWpgngZX4EFtOhD4ZIvBjNf
W5ODvXxMpR8DK65u3z/H4eQ2uRi+0BhPAsYEfMODHZ8BPbj4PrhSBm35L9VqrlTS
ahItcX+8jzjpDg9VSQQh8VG8bqGAmkmkkC4u5eOdKoyyUSihQV9Z9a9gMUiBs0s3
ZlAcLwi9NTsdJ6TfbU7EB/VmXp8CbPiNcCmI4F9stzLocLdkY2laWeqgnOu5vM/A
tTQ5yWlRoxHPQlX64fFqSM6qeQ6V4N7i/2PDvSpDxcjZpCJbfJ651P9UU2OtfOw2
pHi2MN6pcVvTlxTcuuMTHr/5CNdbuX1+QIQCEayp9+kyeDyRqgXKm9V2m5lkmKx5
dl1JqJKSgV4KIRtqGO9q6uWLVAPYewGwCBxNb6GTgtdhdaicHl3nU/AAidncrTaL
nWzIPZ9ylekj+CqYLJWkeVUisJfaHMk4pR8VgINJlLLdWH9Hx9Gat5E+jFyKXBwe
74hHyylTcFqJz5dtQf11ihoAgP9skyNUZeudxqpTzCMz+Mpc9f11OiJOiLpoMaVE
fXoqa9j82QbYGQ5j2vi53bCgMSXTSvHNLXGPChx4zq7SfnGormro/zYqjBDIl1T8
VQDiNyb2htjvRHEZalTHtUekJJ3c4V3MayZ93uUA5rbKAaDfn9YIQ9/y3pHj2M8t
3VlT6GAYeDgw8tyPanzddlsAgs2N1O+4ZnLa24USyoXPzxHdXw6OBC/7jhOpELZl
dXlLFv+Ka7dpp4kkKQUPcS3yoCtwBbc5saa/tqsd6DE+nAYGsSQkvnKlpnOJVBgc
+rJYz0SR2pTh0J7qMyRh2tEOmtJ4U95WOGBv19BJnHMzpIgmh7HBQV2vl/NuTtYQ
h0p5pvtuCcXtOlOVnyycJlOmcKLtajtaD0+CHcwqJ8Iz2FhfhTNCX0RhBG6u6PYW
KIeE1der2/++0QTjpFK6DCUqJj1XnpXetN+3k3MT/3X7q8V5firpkdYu6GOmqw1f
I3DJTGeJ9WHXxqw5XF4CTm9DQ1RqL6bljZBaH+NDlDshm66eAXydLRhwNRKOpnfh
Igm3RTYER0XF5EWUW5EUJ1RszV3mHRDAzUqhgcH3xgtxoQQT1IDX9y+ivHGczry3
ZRkjT54+iKlYU9ZGx+E2Zx9JB7ZMbLiojpzfcH0KrvvOnloha/t83WcWBVv5oD/M
jfBmzG+B7tcBLVjf0yaOLlZn3CKGuI1rLFRKZQfTtJWpWwZ7e5SF30DKvGwdMDIV
QKysXXBadHdmO0A6c/v7QIHdRCs99UhpRNurxXpLJPgi0g1JGI78FJJNc7+wmZu/
Z3qy0LgBuG8ElJifwFfvNELdVCv8kqS3UHGX8pEbCRD0DTYRiVWIHygdZ5/INIQm
3eaKIAnJIFZDwFVEFNNawoqlwe76g2awxN8Ym0Cvd0BGklphYCcObZZvZ2lPL/Du
z5sTdPz0GNX8SCzCyd81lQHdqoc+VfgM82PMiHw683Ruj9FENH1FE9r0QV68K8Pd
iemRSvYRj0aVo8SUxvjvVcn67nwgJAQ4y+bm8daFhsoXdlFKtmRrLv4QqWG9eWX4
AKwT6kp6fCgSjXQANuSJU4O2wTR2lgvc5OQzslBZC2/3nZNiNqicGwowlMrQtrJF
MP4U0VIEqxzTGfBolnXalAiw6R1NaG4yXxa8PAJ3cBVCfMphHiwPQ8kvnw3mLMSN
RUqG4i8JqHcsZS25ZC9itsslBH133n34LQQkZb6P087IFLsS9eTMuXRDNEdZzJEc
9yXFJSeRqCkJrCv8tbnCeVcgkpis3Wn2zSwCjoX2+yCDDc4MCV60JJ8UhYwugrpG
z6kjiZvvGIgVoI5n+kta13Qp3DBGYWF/aVJI6j4E54uLo2fCLvPdjAEJj9sx2ic1
T/BwbKaBeGZQqkCks3k6rqimo9gawD6vr5IWYCykmS0ezjsw0ZHG27hPMN9TN6gM
zZlN/W72DtpqcnZ5fhDlJrRhzXnx0yG7bIngYpqwEPVaAeaxKJ9a6HQRpE6d2UsD
W58RN2BKmhJNGvI2+boXC0nYAIqdCsIUU5WIRD3cg4HsYVxm077nJzWKRv6w44zf
5e6LE1xmZAKgt7e1JTT/MpGqyjHevYmTSIaSy4ko5tO5SPi115gj2nHxKBWw2lYU
eBTRBNhH6qc9JPvEg+9v6TXw/X5NNGCvBoQX9V6/fSJ2Jv5W+tG5e/BbuVPFlZxM
m6M9YzbDXDALGPZXLHrlUAF2y5a/ttLXetnt5N2Zd1cAzrko59glGuE4XGzS66uA
yGpaMY9u6TqVQX56CHTTqaBsAKGwn1nJh9k0HLQWqPb5mqppJASxfKBZ5fCt3Buk
3zWK6hw9snTsYbsi/nfDasUGq4j0RSQ6taVvp25uu8PVY9XWwemwdZYPt1bODulG
MwjgdPnvEJ2FYilBtkCUa7zSVX+1nmhXit1bw/NGm5dj9KNqPyWQzgcNUqMK9EWM
96yquhe9T8Wj6pH6kt2O1PoWc1J33KKAzNducG7zR6phIeVRY/91d22RCkl8DCBy
xzYfpe0WmnPhUof4YBsiOzI3PfX8Sj0VA96Yk1K3ZwCjoi6OYKjAxwJTePVBa0ts
AitxJG18IB8MH5oGZ9kz5zMRlXAc/48AtKO8s2M7PmaIL4OImlKuST9D3scJtOri
nDOnaCF2gfP72G5asS01gUEkRY13Sj4sU3FLTiXJWh8aTxvkBzVt3AwesdtUcCpX
1xOu9yCe8CZZ59oqAxkbpwjZaT3xXwQ4w+MMlcHaKBRQd1ENIaTw7+FoFfwKWOFX
rfsYSdYacFz96ezSfB1kfFBulBTuEBCAOFdei42rTD5KFpOfCDH7BHzLfVmX6ALC
iFa8n8VlQ2MedfZhKVlEYMyeDCpDMK+MCcp0qNoEPqodHoV5dmC4eqPV+8Vsr6RE
sVeQ4JV/W09Ubw0GX5w5ttdnihv30otnfOxbSN40QfghU4Ij65osfh/8MezVXJWM
z2MhwOlie702SOYxf0hyvbVHIDoZCb0AO5kX16gpOEaJuC3U9wevCUcoQ+8FGoEf
7h1ssMoDCuoNN5M7grhtoIZCr7APkwoc5xqUQVcf6IShul8dDIhWQzzJlQG+WUoG
+bcIiL/XSxTfAHw5BWfD96+ReOELI/+dgRGXJk4NKtxQ88pDICJpMp2oioNntDxf
CqCagBb8eVOSILUgRs/+hhzCPLWqYqM/ZuasOEtAupSH8gv8iK2f6M26IpqVMrow
GqLtNVvaubt2Nu2Of91UXnd/81i1FHPqGyqBpDH980AzHNDAB0Xa/sF845MKLd7s
9ur9DJ1aJvdHjGETtPU5vmEqMrbCjrvD0INGgWUzgroNrr9Gk0j0h3pvq7vgLMhp
t+RacTqJV3Wo8ASLEhj7fYlwn2z70SU7jF3goquNBJZv3a1xQc5yACTEu39oU6JP
xUHRwDjafUnJG9CbSKWTQPn6YChI48WQF3tpsZy6Jv/R2ZfAbTLfCRHoPwMkfkEy
cEcryrCG1fBCVEvRPiftXyxG4F8K/TDi7H34xoD96D+rqvzxH0u45Lxihh3qtQNw
xdkA4mLNU8zGoqM01WKHtA5Bf5OWVxMZN5ecUihPYYPpJdZU/QGHLggVMijnO0tT
GuqhhNiNW/Kv+IyiwzTNk0yNF64k3zT7497Hv4fA/qwUKwLpxA9XD2yfn2vOtpEp
qdpPtYVpzsrrL9VfojI5joAR8IPjgUoGFjcwIXSKcZ91NgiE9fIVKwhtU6d7NfV3
OWC8mBqJ9MkynOd4wYEBvFKZvayG+r+T2RVBKqozUnH4DjQUUiyFAorC+lx0SUAj
PxcX89diYXTqmxvlsG+jscC4LQnuLjGewJe1s4tJYxfCkqKm7o0mu1GZIfktrBE4
FmJct9AcDgV+QOd0NhlteEsk9xBGpXYeOO6EaRfyxeE58oJ//jH5MupoZEM1vDn8
x/V9lH0HCvJLjwK4nz7egQG/2SoyQBUEtW3MvaddKWEsjwUC+YvuKpZHSSESYxqP
Bz6srwGAERvbR+F3i9pWkACPvPPo3Np4fuDTQSCbFg6YeyxFXP0zfCNrqyvbzfnb
o5hzYobAmGMlREd555uF1CMHvQHxfZBV7Q41ad87Z64Psox2eDYYxVP3d6JFmOnP
YUGJl+8CQFKMIPxWwlHoLgbVNC3lIVP05vut2KAyqgePB0vrghvBXNAhz4tFJKxa
R4wi+frOtst44gV3flnv/3bIOK///3cdE4+ztXcQoNnmbXiJXdkllJzbecAMIGcQ
XkVH4KfUj6wozUmpr7CBlZ4ghzPudffihiwKXh93mPwdtKfz0a5ctZxcZeC4ZPex
f4Iomdw8i6CQ+t5XV5ywknJWqq/BwyO9K5Ugu2L/KZse+G9k0z+VvPdDKJxAh5kA
7XPWnxEWtIModfzd/9rCLHAJcZYYYE7CVS6fiLAZ/HiV72G4eiTWAOBh8O61NBat
9tEEhW24JALvhV5ZV3B9xoJb9ldQEIqXRcC5n/KDa7YFnwOt/KfO1J/RXQu9F2pV
1TcAX5oKeMxHfN4tFeNj/NMv7mszTUOZU7AHz+ASP5jsH7qJHVj2OiY3LHHHsXZ7
Fioz5G6RvdkYruG7CubDRSxqcMXH9MHJaM25FyGxBYcGDLQqQHdhQHfmpS3PSdQ6
ZQfcLvRmT6PxxYcRdPOae5o639ZFAAGP24+GJi2WO+wzMu1/3L2o4gBqK/AhG/ZT
41N1C/ZNwy+9gW1EWpk3YvsWy44FE294OggoHDJeiMMAJ2Z5MFVbT9+WyX8SVPXc
XoZ8jFYIYvAbDRrGv75Z2MXNj0Aiec82fEEhewsKArf+WiA4WvZ3wv+MskuASHNA
tHuBN9l2PCF6dYntNYxqs+42Rrh13cEoOTEIrW6zwWukp0CgnWXjQC6ChpW36uGu
UAatpnLCIGg3TH3kNtraAxQnr9y81wvkxQ3dzEq+SsPtf7qRxIq5Q0GE15ZztK9J
eZqafnN9mMHhmTRBAO8+SacW42dX8RT1KhVVBVVReTzJKGThdvVtxjGSpFaF6y88
WWy+YtUJgDGj/ngzfReZKYwm9f/q+rTNWzxBO29ClCMeBHm3QlmyA6w1N3XNzeiW
fQFwLy19IZlSUlUzb60CjpIp6xtx3oYsVhQjljDi6f2kdLvrzmU8LNv0DOZxku6K
Tnkvbpi+RfKzinMNr4Rvq4OmGp9A6nFA3MkKu0NTf5pN8l3GPZnc1Z4lxpmW8NPq
h8Zmno5U/6NxhUpn6sToQsQeChRYK0GrIuq8wAO1QgmiSM1sDtBljPzFkNReQ32F
0J7YfRN82T4MLyUM+J2kX+a2w5Y3i1OaKHyXWK7mMrSEzA4CRARVxuLmF4KHw8FF
ZhwszhJIZlUYLBXM2/sTvRZgnirP9sOpaHCptA9e+4pv5umm5a2b/dygv1ASCyck
pYpNMnXV+dxyFr3mOjmtnF9NSEqGWIR3K9OvuYmpCHJITPS5eBSdW8yAdES2OCLk
LUnHnATRK7MrUF/xN9nBQxlFV6VPon4zmt2MPrvOF30mN0LxXzxVvQ72ygzlwI3f
n62ejufdssE6lj82MzysPnJhMeJnwFzyTQArHHsXqs9JxHp6tdrK+V/6VpQo+V4u
56Q2d6EUwTS/l3uxX3s9loLjcHbde0g3qH3TJEiCWyj5pg3CmwdhXgL8+o8KgQKf
9zTRFwLCNhFCWLHSy9y1qFz1lwplHzcR6DioEUw/faKL65QDL3C/W6v+01lHtdCV
/61ZB1VAurP2gGksuhw/48HfgWkp2OXA/ebSm3oihzwO9crXt+kTnPcLNF8rga7j
PZ43nJaLZxebCSB/bWFuArMoG1ZZ8DKhX9FbzwIZlu2cI+8vTRfbCIGd4JwKoRuj
cMZEiqth68Z4e7oDy+WVKkjqqRd/3e2YqG5mUUmHWrAmwmUdgyJ/3nWRvK3CRIcT
5uO49egcHg3sXSLh5jpWp62vINEYpx2h4JwivlQb/R+MOjWXPbzSvoZVETBCvM3s
O+uWAcOqAeEiZM4wDSwdCCo7vDR9fULggkBQoz1BbjY4mPIb5dECzymiMNDLV+IB
tfnYz8skLYgyyhHmVYs/aUWr/nvYPxM+5rs9+rLV3io2kVwI7iUKhMnshzOYrjJ5
ru/D8s5bgJ7WrKNTRzUkOaP70VsKHigtYVsu9kEdZx6WYwI7tPK+3YUEa/fK5itJ
Ylf0VAonzx+y2EQk87fvoOwBo4fnJ0NFvOLSMlTGZkwDC5E2AcLnmoaFFS1PFzTx
UEZPqooLBJy3ibfFPX2af3i1mEvcakKHqqDtUlHjWa0XvOwGToDTYLwFfhb8eiMi
in/JSMy120V7ArJwFbiKW9V4Ar88P0yGZrYzJDHop9mlNFs7wVnb+sS0qQnOfAyM
NusrZW0FAssnB9bZ0IFoe8slhu9voN+cyTmDEvOsS1n/Sq6e16r/8s0nPgLMIGPC
tUajJPjLNR4baC/Y36FN2f6UO4bAiq1TwmrBQjaYlW/8WURFUEOrMnxvEq7ryl4P
0QsGGCh2IujKlZeeozrYk6JTzjVBprV09y+ojse6RW7JCLsZ2KCUuRbnkwoEldTc
VdCzm03wPzgwuek+9Oocxpgs98GCSKadMPPB19WJ1va2vV2VMbKsW/Bu60g/ayRa
RWA7rEUjrSdqw4Enx0ijnwogDRbkK02dwt9lWHw5HEJtesw7FWte3tUYvq4ELoED
uRlQgk9OjPk6+exbycLkjGMbUWG3CYE4oKjFJEiIYTeZIODAky5C+2QAoFGm1vmK
Dnk5fSvIeVg5vj+TC3LdH9u9E/uUr0uZOlZTk2tp0XwQ9iGxHKCDJEhSw87Be9Wq
vLIe3yotp9IZXfkHOVQMJWRaoN9C6TFWCBaPAujXPbWre7XxdQQsRUA/WGFAUjhF
uze1JODZtd0ok9XWm9z9ygZFxojvmKbZ4UdWDK6oR0lZnGG+REmwvyvCgCxN5xJw
CKXcfgiPlbbao0M64YCWSh/y1anrZjrK/00TBzhFAlQqMPSt1tB6yBZVZLiJsTg+
1x8b9c3xbRmyJ/19qoxr9arR+tdlxluQQVItImT6i61NQkN/xDZSo+DyEQh9SlJm
H89vf91cs9BFNz98yCNIXCouHieExbtgP469Q7+odi6f9YtNXomuX27c8fMdAfuT
3iKDLGZEksADysOcUFyK2zuFZMZZCc3JYC4V4KcT/nMbtiSxT/sFE/5PwBwnP+oV
wV92wS2x5QFBTzyySAw6htURrGdjCRzu7aCCuUkX7r2gcnb6HlXLO/XURoFQewvj
Ir2ouw/Ryf9NiU+frzZGtSdQY9vTP5WQ/MDPt5LSZ0eEUdpZlFfbWxstUb3Wre+9
zCpB1re6NwMoi36htveRNIF1UP7+9y90ANqghSwSA1HPuq9AhwW5zFRiKq/UTGFV
fcoFXxALmhnwDTppQPDJwIthxzfEDfGkxq7GwdUkTAMaTgjy2J/HXZjTKhfsEKis
eoMB2x2zmZRJI9goO8FdawjIcbBXtqqkZNqzsxUHV5L4W5UvM8Ja45XXbtZOgwUl
BzSbUv2mUXn5bX8NnyYAv4IQei+xpFiGxpYGGxA7j773daZaLTYDo90O2SEBEJD4
PqeTIEsfz0KulIrQXmB+wwvHi86ADCtJ8lDxhV+Vte5G8uYPFK8kAwRKYjC2sWJ4
6McEEBxRtpkaacg4yMjYxbTPb7S8ahIA8lpcz7qqeZ0ruBTMp/iPzB1q3DY61+QS
T4wFiM6zCcDgKmYxAQ0CXxCUCMsRXh8A1pJIFO7kNEwaiVl7zCa0A01aez62/AnH
KDzztEevA+1o+QzIq6sW/8w8mS4jxBCxh8QbASXC48HP4Pb9900c3+0CuJUA7jbi
E+bunLtNCGXINIo/uddnsC+Cjg2vpbtbvi+flPUlyDI52yoscdY+46pR1IcMW8JM
sV4jkdxakrb8POOgLKMqVwWKCchQmTp74K4QBYAsoi4YwZxqdMwgUJ/c6+0yNqA4
WYHaT8KoeTacSL5f8RsZ6Minxio2ZnD+B25Tq4kqhFvKPQI2C/+6mi9LQLnzLMDW
5vyK6TIwBV27WkLnYUqs8pVD7Do1Nc/j7VWBTnw2CnIYU4NBPp0azClhRIykgonm
OW/2RnTnAspW/qNlt7P0WUh8P1nNVSYKKv3FxMQn77M/CkQMhpBKZsJRi5n1KjeY
IdhYaVBrOVBBfiH5fiqgMrKau3XN2CeSZKUsnMIvQ7AOSiTwf7NvRnlv7N3nd1Oy
Pyw5KfbrH7RLiui+w/pdCl3msCF6aBKMSt5JqOZ64JVka6yjpCMccHriDrBFh8+e
T1Z/WbmoJ5Iyg2s/LSCnrISS//L17y0ESpYV3wW2UqP4m+cY1Zpc97+l9M6QPNU5
MDPTG213fPA1Lmpe4V44XcBOWkllJkBF1Qp8acv/TdbQ27qdEE/sSzpLIbkcu29Z
TEi2989wJEgiaZC+c3AffLyhFfx37EwNvByetR29qktBHEx/+MHP5rttjf8wvfba
yabtXBTumtQqAB+NC9pCxSUWmX17uEGamjA2p0MwD4zoYP4rvNAVsSvgmT2HruE0
9K7LGCKUk0S57J8T0bdUFGGQ8SQlEPWixtJrJ9KhPxqYwKZ4ZG0mHY+Ti5KTMXJy
RD16dZH4B2F5eS5AxnGSE8GPGABIazRI7A8JoDuI2WQ8lzxo44o8b/sy8CTvyyf0
/0AcRHNgkZy3KnDtc5Ra989TN/GB0gIffmHdvKH7721WW7Cm5liVEodsI0oyidQu
x32OpHs+w0BJq8rBH8tmMe64Fy5CI0GTt8NVqR/TZVZYOUEDA5HxC+fda7cMkjh8
AUrdIwQ8ZiSAilI+lT6i5vUCLwdSDf1eAxYuK1v/bXkomrKC6H7rChdOgMt96B2H
dtoB6thZISLR6x+T0HBXjS5C7XtCW0l6fgP0Tp6F0RDDq0VHd3dw3GJuz7bXpJyz
Bs1SPtcymBJOYXCwIn+M9XyZ7weXbewpaBrMtJ/ZXmgtJHA8RbNNl9mkixXCEu6a
g1xKNF6/NtujtK/AC7QHojMF1+FscGRyXl3XBRrWJqFqLY2NA0Zrap595xa8L5Uw
0S1xNBOMm4kgKcG0Xh07Jx1VQCjPx0dJeq4Yi2z5XmxzTg18iy1kMZajG4dtZIxb
Grk41HGpL8F+vgoTkLpXvt8VzQK+3zfHJq8aq90VpveBPvXcx4DUvFrGgGRYIi8t
4O1ZQ27ZT5ES+emAnS2FZbUBDEN5dZ4xU+ACQwT3VkOxUzkSB9vxg4SiLb2Yo4D0
5mbDU6/aItOs6YAWxaSAYtNt6PkMNg2lERu+vUN/GABQkylfVO9wNXPWzcDExh5/
9d6pRxgHR8THCPzT8pIs5Kfd27IaAHQppD2pjiCWBfYglDS17OTX7zUaIsnxA35X
zg8iM6O3Gukl2lAUptlqSGkjlvD8+KjShL6kC34dYPdRiwFbmAjEWrlIG39b5xe9
5cf+KmrlJvqd3Qu3umXUEwajYCXkQQYosiJTwF8E98zs2wH5JuPq+RwcIfbdHOYD
QhhZqSVL6NibN8dT/RKv8A5LHy9PkVoCdpkAbwxF9uxgxQwp3kgW+KGRMNxIMQcO
Wbt/UU00O2qg0T6hD7rOGE/03mKECYXx1wVCHGSCeP+fa1+Rkeexu1Yiq50XyLtg
XuPQrCZivp7m+mPhOH+S0fZoQugHE0PgYeE8s9OH/nssIF+1pSUmkln/dNbvMUaB
pEwDj0kDNjNGnVMt7s4e+5G0R6+WsofBorOJKx7U23PQ+0lG2dQh8dq0V8uyTUxO
abNl+sEMzN+34b5od5lAZa9OySGF/nEqC1k8PK9fwBzwu/Evo1SSTwzQEzin8BTx
y0lO/t9Tc/l9ZGKFk+AyzEsnKuz5Wboiumbx0LUJX4RiNCYO3GYCeIwdDzmeJMmG
nUiBZcm7ff9UpBjfsQFjFUjx9rwK+hfKQ9kw9h3CcSNT7Ul0FH5GtuZrdW72txeu
y9R/233dNoFQWkpp8VbdjFNv2IYloECAongZwns0ibbaElMq4R40aUp/fquoTcsS
LbhHeqs+6pKQRG6c/0/U/ugw6WDan+GwqZIwAE+4KWiRJVwCF9xp/Y5NkcnW63xz
WtqDmfjLLhW/G2kt18N5BI7LCxw3hbk/xE31DTR3c66gF7j3C/mXUMiKq5JRw21/
M/Ui0HjmOx7Zg12ylFg+QVV6SAFHbwfNyT6008lsSdCeNUrdNNp8sGIk2WNriqo7
gFo7QVVw0/ywTi93oJgqKASH8f0zhMBpvV86ifMaW0A/jZFR8LfZOMvhh1LbSG/b
yXDuJdWstDaeNafqoobP5v6MeKjef7pbYn6w4eEmuerBD/KdXYyIAk3vd1HtD2KR
fD7MXqTArFKDE2neB0rEdTU2BF8HLp3+iYGdKj9PvAnL59OVPIwA5QCK6OeGzIE3
yldsp5fey0v0MraBpUcMgXhxxs1OWgane4fvw6Mlf2cIHuFKjGlv2ZFL+2zilxO2
NmjFvoOKAzaB6jG2tsF/1CSd7qXVLYwLPEHOgM813MNJug2QcMCYEZ+MaOAyakTi
/1z97K2duzI+GzzFVCxBuUNFPNc6nbl8NSgFT1nVDNSR/IIGmDnDG3K04Tn9qaDJ
tzomaWCOYGjkJg8fddJBdvpObISiFjuvSVrFp3lfNjgDLBuUAXlls8FzO9Nc5kH0
Nk3BxZD9zlHKMFui0X9NPMdt0G/S09ggkO7jiVJIeyyMDRiezcAkp7GA3nMDErxK
eMeealqq6zjPOj9z8GkduklQx14Rgyt9eMH+Dkfjs2/4qKdKZPzFmmvcA0eQiNmI
ZbhjHLSHWZqxcajHIb2HD6p80jkUFK58tI6AmdngU6QE0o9Ljy5NiAplhycfgtwO
zdluCTndB7xydQRR6wUpUQWj33xdtZVEzyPJqQ+26KfEmMr/dBhcpZQFuFiyND2N
ZacTkqCJXB5eyMzrDZMSzI7kSIKFpkWLoyeCdixa0R2WvX2kBWcnTKuO3UYqLIf3
FslIK25fGP7+OFaTWNspKFrOu4YDZHGTzqHwnNdH3njcM5FIy1gCZyyMhwSNj6Dk
fII/PP1Bu0JK7d1FAS8kvP+FQSp+XNHkO4u9fjEJMYVSOX8W6ib+dnGN7Wr4MAxQ
lWvZOW+5hGCORlOuRrMCKleYo3siZ7ER2ooIE5sTqAdy6+1RDrKnFrasLPFt4wiT
ORwxm0BbpHv3UwRv8n5Wr/Ov2ivVbOv/kKOHBMqaUUE+L3Nl0E71ci7sg3MvjdaO
Tor32xqf+PLFyAlm5hUagxsgibc2krZu42D04iRVU0gzSQy2XFUxDq8ypxDRWVKa
ImSj8Kmv4wavcJmyDaFK09mw0aU6pS1j+qK1w73MEn5dfX5Gp5zRvwI6zXlMRarh
dbw/jWPmjyBpyDD/SpTTsNuD0gHabp0n0xFoV/xg2rOXSBHvDIWia1TDom2zom82
F5Rl0HmxMMtLZV+uBJJwYwyCxfQujLyiwFgF6ShVajftunwEc+X1iqIuTn6nI+8+
tuAjXvuLtq26ltOXrJuhPrbLM2SaSrwDdV/mhsRirDi8MVyh/ZcJnLBBtYMICfVZ
83EX6rX4QKFYy4WE70iRqW6LQcfrbRtZgh4q+woUlE1Vda/jmd+DgdTjI3YTD063
Y+o4F34C1WSpBws9eor5ALj+WpnVqE9cdbfYzGKUT/TGZMHYWaY8JMq+5cXeIhge
XZixTgX14VVfjK69lHluFoNlrEFoGpJnWrlZNs0gmutr2lvN87FABqNdmR5udDJL
j5aWaC0JrutH1KfvYV+kjwc872ZGPd4AH197ZBhMDYNU22ysYnlm6YvsEnodK8L6
T5M2yQtTYHAd48pThIGMCV8w9kvIlvoDi9GzAuPZGQe2Fk5cI59aTURFPxRzPEre
T1fNSsMef8mEkP4/xGTDbHkDl7wAzwCqCZx53abITwt5mDC1QxTkzR0CXMu97lmS
wXViSGY/KkrbThMKQl1snnRxuIZRhru8vOqVXyWsxxyTtzaKWzRbGMFT7ueJHKbw
ebc9i+o5Uy5+udaI1Tq6TsFqFpPhc4JrmnVvuM9M68Jn7aueNzgC5HYEQdXmFjI2
8YGl0g+8BGtkh3wbrHXfxRC/5WbVkiJ02HiG7JazGiYqEITa5Sq8HMtojPul6NhS
LZgB18h9Og3EHFG65+kCg5qB+Fuw170XGM2dHnLalwdylxYV30AXn4i9Xpj8QQbf
1Lg+pqPPn18HvQFB+VGROWBLGkDE1NEa+uoFwMpUGe5uLt8j0DGFAGB6FgvzsQzO
pgOn8wpTBjVrXOPZBlhrfNbVoQAiiyeZegUbFZoiLn70xoq/wpbGCjfnKG+kQPJo
x2GxnfYIkyXK7+gg3A6od3LwwAPXPWdNegdJxLVxP/YwYBLo5tBggSV7jD71oNRI
VqsIuVYIRDXITaFIOpZRBG8k20M8/7d/pQEcFIzhVRH7yBavds4sa6vVBsZiqnBo
dHWHShKL1X7H2w+l0u76To6n0JjEGCxQcuv3Q75gZhkAOgVXu/0Ojg+3Rn+0Tq2b
Z0uBDAoM9N1OKw9+boYLOaqBuuB5kXBQC7NZnwlIdAwn8GeucIBbcoOpcnkUr64w
6YYnKejuzAlZ1Bf8RM7/zOXZxgFK/X+c66AP43irNCRD+3FyWFscWMdkeG9cWvsv
cyCZuf4NHP6jQbI9FRdip+A5T+vXFC92QtJUpyHwaoFrzxexWd4OeKuV9nim9sJ6
Z5uI9tM6o3FW7+1wJarIKYBNOrMpZ6ihy/waGWjwVp1hTNod/HyR6rQ+WoYMEkIu
LL5sCJRfVIkvD5+fNkixdoQ7RBZonmHna/lO7OxZu9w+kmE+y6M968y+bRjVYnXw
EJciPpJqlhpgXul4PSf9YGtT+00fqfqN7szu/FajFNzNNW9HDgtAAHWvyEgn7ueV
QK7Suly4bSaASyb4VZSp9ZWbkYai1SowAnK/6ok86l0e5vZz3KOAXmrOmfqtSD3H
Jlvipbf1K52qcAV5uM6UpGNPHvUaUqGGfMxbVxeMMeb8eLd4bM7yfmuOud/N1NZg
W43bQ1PBZm3XkFqu3Ys3eomyjptM78byNF4fHoVbZsfpT59m71XSbxzsHN5xYdJy
UPH8WCsZ+DzVPgrYrnKkat0n7Y0BI674oS5U4bVFQ7tqsPORfBNAO/b0/14b1ohE
izF9RhaPE1OJwNWnmECTuLxT+nIgjKwU9mZdOq2jOl6nMwWGSQD6VwHSy2cJ762t
ptSA8ME3PaK6N2d0TNkrEqsYnXe0wT7iqMXOVwrQ9o5Xez9H2jObiRa8+qKS7eSF
t+EXbVLndrYWdhS1leCEhjMuXPa0r135p6A5rs/EEg0GIboE1cF1v4yREOyb0+7e
blCKhh+JnsQLHG+cQ+rlgsnxMdRFs1x7nvtmJlFk7uIjdFTgN0oaZ1pccfsBd/gV
lplbdkGrjmKPICjNWlGcWZ3QyY356YvrauTDsCzcLTNBICVt0vRhn/zoCDK1iB6N
CXjaXnHNHi+6Mu+epuABkcnxu+pNz/r2L1zn8OyIN+tqNtH+q3EE02ikWD1MrqgF
7lHJDE6DOsf9hxWsVRu3Jaiqf7lGuqzEwpdGqjvrevaYvItcYoWQXa5+I7gaAF0r
i3jyeZxlLloSMRDkaJkRH36KhHI0sYKJux9f6Nw0e7cyt0YXW3SY8OFMjuzdEnUi
GoWY5sLzVm7Sq9hD7bzb8gp8FaVKO58giiw7IL/IqNcGFS9GwfgJ8Y5MtA+tQNMa
gC4L2422iEZ8sNzWfQTd/1MK50tb29cXjkZBPL577F1FY2MqgNLGm+qZuOjbmMup
AGZNo3pBpCuqFT6quQE7SjtbIfZxJsEE0tpA64SOc+fw7J0fCzimU10HZrl2tQQY
8w2i92LHZPwZPdWu6hye/I1l0PSDGO93g08RvUjn9I1jflZDROZuG6D0qRa2xaBB
gxJ6ElZ52cSGY49wrApHpVy2QBcPmmLkwiCo9u0MkWCEAUWNk4rEYf/iQ9dg2pH/
CIpZYTFOy5XC3yd5vBFC8PlRwwdHp7Av7e2RessdFn79PYawvXnqIiSOKzhfW9xY
ofU04ys8RgYdFZWm9jVnhh3zfzi2auETnF/SwwsMQ6MHOavmk97a6NxhVowKhL68
bnRLX04kvhGYTk6fpUhCwFvQxXhShm3COQOtpdWg3jxf9XPDEwYDaSC7G59wMgQb
tT9afNflr6HMX8NKK8VumfDrFyX3YU6SR3+uuu4jnqSFtgL/jhDil7udvB1H6o5D
1tN+hw2RBl/NtRsNSgfZY+3YAziM7c41y5N1QK57COymcswqWTerLSLuSnrxYpee
zSy6e8/J2GfJCa1re8fcoENnRdJFwIUKlDMjgVgIp3DTcajj08H+9Cvtygf0zB56
DLX5p8TxJPozYtL5l4IrI2vQWfZLw3jDaigXt17JNHg9GvoC42psH+VRxESiNz/8
gUrjZRaMWNEewhX5iSNcRtSKHKgh+51ORGGA4noCASmE2PimyGWIPfhDqQvaFCPI
WobBgqis4+ABDcAaq0UXoPSh5jUDekKox14U4ARgcUSV3hAEBHf846xmZo5aSx4p
OdRvstH3Ih8qRGjSHrr9p4FsDBa6NP7v2pa8FQ07uCho5JRzxMiU7tmsYnaTzWg+
ggDnw128SrALTDbXahP2Mjb2E67RPp25s/UDJm7p/KjespoPkrxw6n3w98J+UoPJ
hSssMwLIQfnIoeD4Ger9XS2d6ds4Y5qTJBi5yhbfsnLtVhng9xdEpfkI5opk6ce8
Uz+drZuzJGJjh7Ff2QAvmsr558DPnmwB93kwcBt1PJ1+ezyPs42J2ufPBS/XgSfY
UJwGmkkzDxHa294GLMt/cUlglHNqBxrzFkwmhzL412jqxqkJjb1RCoZ2NCXnJDp1
xARIr/GRdt35w+U3pM/CUxVOqmlWh0fxYSCEdOLiOKgIskDzxw9IQo7XiCTD8VQM
Z042INQoFjw//bb3ywvxL+YPAFXzijeD2wc2yU9rYwV/IlqjWIZY7QsnzLFoRBZ8
CJnV6zPfQIfkFIO4jDiBpskRBw7Yl0/VxTCkIpJZhdqXsLqdjhWIaB13TNlp2827
kI055lvlPjh+7ZzR/rSS+cu27g59daqC7X6PITBw2uHyuukVfAlREDalsI/6FjxN
iwBWE1vm4G/Y+egkc5iqeaYLaHujSwfoH0pUTuiDBIAYQeBSTQXY5snRzHuy2hIJ
jeNN8+9h4XkPWsyWLEZFdey+xOsuzP0msqkycOtOpH74Fs1wfb/AHcPzakzhAWv7
YgcRIzFeeqQpfec4VP2DtH67Pa3NeSThqbxPaMOtvEPg5Y6Mu7jTMKj0Rl0ykwk2
edNrGMFcsrxF6xWBJDssIHh6mvr5rP+m2kff7iYLDn3Ad0JUWu5VaIqs0Ldv3nZx
ceHs1aOmeLMgHVJYH/+tACg7YGxEDGXRzi6LyFyt6Zsjj7AgxGDMD+3LUsCz7AKJ
L+ltVGT6uT1dKO0zSHsRSiYykcjOKWAvQvflGOgclpXUsNciNsxROfBqBjaC4pff
6dWI5YAM2fEVL8GYc3xYCqJc9hg/RpQag32QOjfRaqEWdCchm23KUJQ2rokmUKzZ
+EcWySMmGooRWJuRIg+1DklXG7OBWmpP6NBLwNKh80EpDM8D8BaXCijRorQWbLn+
tr+vTvlbT9Fg0vxE8gZVT2fRFL1l3xAbj2263NISjxyO1W1ihAY8fURzJwDxofBC
qrsXEKYdvEtJ52oIGZpSHK15XCBdSe8dctPzSGQ9Ium4OfDZ/sWPtS/w+ULeDWqB
J4Y2/UHWiS+FGq5AWt0CpT4uoew6iPm9FatF2rMaMzShZQzMbb8eyPokC2nJlZFj
TClf0fgKGCqDzxtaDi3k2XldyvJvcUFytj7m7AgTmfzLLLEKnFgVfs89lMR/hE6v
CtHPrggImZESpniampdeL61mzgYvpmbKTKgd3J+htk/vxjAJLkXB5Ze/iD8o4r9l
Yq9s+hoGolEcK9CM7gcZqzhqVEnJLTG6EBJQjG7eQq/JK5LNB7Rb/AOH08XvNLJ7
LV2HVTPp6EBpDkwQbM+GsNIpvUefYNlAua0NuZb6ncWePCcTl7ImY+AC/pgukVcA
Nl/wqcJQttffs9JXVnLNMupFoWQJlOapUmVAx6Rcv5zxdtGpFfz3Gmz7UWw9k79g
VG+A22eFYZ/MLDwLxgQCaeZdlTwkyiJk2Y2f/jSjDIWcsDx60L+o2Ro/jz4I90I4
RWDgUdYGQzd+GGPKoTphktet3ck5QWzfqpOAFvn6TktcOvesf8e7mj3ACnVtd2Bb
Uvi5Hn2sBbHM1zeMm9BNulrWX3JME0i0wwRhfSI9MPwapV51CPy9o79QCKc0c1r5
9UqOcx5TrzBOu3Scl0phWq9787KxrUnwwhR68RXh6n9XwEAKPUmkvkwDwZyYvCjJ
kbkMnWEepLgd1lzW8jl/pNvRZSJ1eyZRdtSowAQ6RsTCEl2u5GOk1UwA4506Lktr
gVNNMAv1bioPMkwwJEjQBTyNlbHo28Z8lcczx3KTV7vcPDUSRuiOC287tUHhZTTa
6K9BZIHAmYDZNlId/+rxOJVrg8TfTfj07GtpWOBi4OBvZROmMuZnhr43thHsGgLz
Jl7h9f5/JTukdYPYpvDexKdSVgw0mXlQwCNzufe4p1I3Oudad5AQAaIDUvA8h5XO
dHJmCgv2nEOGevv3GSpzLnWc1r/CK3f4QhvPkT1Pwg6QblQSMOWI/n+geRhfrs3t
UgZncH8aaU9mPosmmR7I4kzQOYJEmLAkdCF9bgZFQBgCm9FiANh791ZU3cQiz8IK
KK96AQUzfpOz11C5XSe/ok+5KnRRXeEYbi80mFQvrPIjEGX+cu2k+n1pJo4eQkl9
CWmRF07u4LASC4eal9Qt3euTOn22bg5dDo+MmrqLpgSKaodeM2o2G0b1cC1/OymI
/M/bcdEJBOIXqyh6mRzfOnaZ/iaslJB5o3ZDsLhxw1EnQ5pdeEzYLJ6CHWE5wCr4
rjlUbMxdee/NY2Pls1a1zIa0yybqanB8H/OvnMgGguMljUxRrdbdHZAVB1HLu2tt
Bk2PlEORmxS2uoS9Gjoq5OIq6SY9D5l0ycpOjyyDUwO9xVkGC05xeSZTo/7PyD/1
wx+narbWRBjE0j3JIO2XzZsyucrXVfVBrJ7mUQXIO7Wz7H2ccSf8P3+PeY/jlXUr
SCvuWKUBbmZA+UfIZDUmkh3Nxr9+oMECawZAGF+Uk0AgtgSgXI2Wh7uoACvWMY6I
jXHnuzsdqxblMbJ0Aasm0ItSjWWcCgujGlZg/W0L0JZp+cXsLnizLRnYLo4byoEa
7gSiuO+Y8KJf9jtKFFiw9YCXGIUVot3dl6mwCWtpfTjbLUwgPD0cgtjUBAHa/0tU
lPy8EWt6qACq0pAb7UG8hiVKbq5y/7gAkCgfyb0Wyuglya0apNv+qZPYTrrsWtl5
nHQzD7h5KILmwcTL0Uotxy+cLIb+00g+L6EHr9JcBDElVxwrNhoecQiqrw4inrsO
9pZyKQ3rd1P4qqiXp5Aye0KKs2C7QrznToiBaPdP+bKjSSVIiqWLm0bBctZdsOIF
uCGd8+qjgivFJSB3wzT2zI82HgeACjfJTAxpsnpkOsfV2G9gc+V922YBRkgQzGtt
x2lj+5uFNBTwi0JBFEzHGhP57ipcLUn+DyMbHzQJirZfgGNeCuqd3AEB/ix7H6nh
pQYhNm8GrJxiGjrDMjDZWBS/eQfXOM36u6Vq7LX+lGLpb/gjRs4E2+vkCtEruQID
j9M+GPr9gktmC5tWxoLaEp0ItonuEea5Z1Fap9RaQSLtBWigU5liePl+kU3GO/oc
sRNt21v4XlidT9hlfNROnfnldX2X8khWQIT5XRK+oV2hEIEjkhxqyS0IItHL4Ses
XYr3SuN0MGpnGLCSdCzSp2tYoCXjJwq1WasdFBW7Ho6uys7fwHmYRIW0FNnT2MXM
uQPz6oVW2FeT2NL6D2IR+YvY9u7EcTBfuLGil7uRhxmRVfJWZDNgioD77peHCm35
Q05OK03rnlbXdZatVInstbQPYMEnvXGJ+0MNnbVP5e+dqfYT3CpiZHsqYIohwYhD
EyZJDYavtRjxFKGHhG/DLAPvvXjUx1d/bU04VNjjHowcWNAAXaO+RZq+YsPgDfng
Kgr9rS49vnvODvQ6sCMLK2TJmwZU4/nsaDns349hIby8FNB8h4eCpt6plx8W5z7K
jdzyYPyTNOS5AIRvruowAjP+cJ+jE7SMa9p+qIcY1h44QeyNm/3knbUmNbuXLTDG
B38HHE2Mw07yBeSX/F/93vJ5G5w56BwqwKQn6pGW9hYu/YMTBk19RXzpa1uR3xDU
9akNHeNDYPJnzKRB8yS+SdyVeIOdZ+H438k54ECy71M642h+DxIU8RJLi+rzVWa4
OMChQzRS/ZO8mwWMhNOcGvyTKtBNydB1teUluFG/FPvWXo8ZnPRf2ahAoksrLF9m
25VtaXpjYV7zshOkAKjIHrlcUOsOySR6mE3rlH0Xu5QQDtOlHkOvuThkgZzEN+6W
sMeQL8V8yrglJ+lnNjdyG0MJ1sIIjbsiTZLvvUbxIymi3a6DkDssojU1ItDapf1Z
9GM/qeSz7Puy5bJJPc5WPmbvGwVNIHILleB00jQeM/Iy/Z7vmJplqU8SxlgTYOHP
SzgVDO09k0AvzmUrOu3fQZ/m1LGnj3I5IhzI7CHTbemS8wik7GLAJU90Dkrg1xsf
qLdasbjJmYmTunoHAQV/5g4qsLN7oioe0UxpY2a5rC1Gj/iZPpD5661CkbjRIu7w
nA7hH55Nt8Oc+EJvv8WT13vPl4xMcR01jfpoiZYT6zXS1j1DzsoQ3K0iHrJlpsGi
lQxu709PqIYdrCaGlZ5U5xeR3xC9mAMT9USn1SZ4Gvab7val7nLfkm8/0JFW7TIm
pjWimax93aKtSfHhFrgKO2v2iVA+8HWbD/+j0eJj6RCZkFKzI79HKYyx6IqWd884
nOLogIwrDmz9lc9LRYixIBEpxR1o1NTrb+CvAMA+JOzzkPBPsaK+JfXRrdVHdwgx
eSzDHy0xDZvP7CzFVbD/TaBWyiWaN5hJ+w3qE1q+VB3LNq/R1kW9UP/gVTuJb3bh
yJC3ZJfeBXqoS13mvla0VOwvyZ6mv3qieF6/QY3toJ4AMbenzPR+4hC36ktTUQHT
rqTaGYL/HqxFG63cu/xFhLPubRWrJUusUQwe99WJptjQIwllYtRsoTrPye84f6bQ
FZc63NMlpIFV6janj0RRO6dEnkOzjn+QKE+Hs9zJsWWg20uLTy049OV0mZGWwKDm
HjJUrPCT3DtvtrnQ4eXEipzKj8Bul3VcvLq5OkVqLBdxdO2kQYqXr4nknPlWr2Tg
S2ZlW08d3IxaBjOlsMFrhJ4NUYqUJKBVl+jOBXs9Rvksodb5tcuIXkQpuJSd7vJE
h24fkCMis8viaxft174RmGVTL56g4Y8IUJkAudi+7GMxGovNVb/NZss2CBL/ACPI
onm7EwXKhBAugeDAbKe96zSAmpU9Jgx/PEFqHKIvpRTLMF+/y5o2nWf5b8MpzRdC
Uxthck0shMgLQlcLCezfN4c12sOSCAmMk/d0bEOZlTgS8EpJwzW/gk1koUcg1z5O
yOUGuGOT7DG95dhpIZuz4ZQVkGB/rq/h3zAQ9lFpi1I/L6548XztKb/Ji6Ps8x50
XttH5cPhHfIdzOtzPNR9xiaPCDSvs/xrVyN/0TKvRC92IFlL/U1gu2ITpS+t57qg
bHNryq6EftKl2wXwZ1Cb+8Qk7zUR+3Flom8fLuNYYAUvR0rCDXHzrpbraRIREzlL
cbQWY3Z+/dLufIs+kUmbRFNqeBPOF7Awoiiqjh6fSJKhjMbO4doWacGmIy6L0VUt
uh54CzffuJTw588PYfhEu6Ai+FXFD5JSp+NVQnhCH9TnQpE/guMyFqc0vBsilyFB
Pi795lcdlrPeO90sLTxBs46X+s7ZrpsfZ/VXMuBNNObTdL8/tC7wYrv1pYVSFqDd
/7fTa6c5gHzxtfdiGKC0b2FxMVbYCnVt1gVufWDI80jPYyNZMOzirjoG0CsvQc0n
sRDT5/KtEtTnarfm8zDUWrhdLBbDSHN1PLDqBcsPhljVOjcd9f90KCelnfYIyo1l
kkUbNhb7SlKn2Mu/oHU1HkqMwm7AkYn6rm+wrWlCk11ZHeJZV7pZfLSXTvTmIoqF
fcmNvt/my+i/A9/NsfntH2UXyS8bRccLAZ3+kR0jE8Ug9nQcrIDadG0/8Ef7qEgw
OzapgwaeShR+JqhcR2OfpvuDCtdTNuzCVtXFH4jm+5CWr/4yQE2GOz9ePjfQNIvU
y0TyLl8j2aa3m1aAGkxoqoYwtc0hLfIoRnnLezCFQOs5vHPRYyb25JX1WI6JDkCy
sm9N9jaD59Fdsyl9Znc2qahifLEJv+oGJBAxBB1BsyO+c+EvNSiYiVTO34Wk5x1C
QL1hFZRiwTUkaDXMRIVFq3EPeDnxBZD4XrnMhtdwcp3Xt8gxHdLOnn5InvcVyhb+
kQokvPvAeuuiCHbgUn7XUQZotLiq9t6iyjignxPGv1NMSUiO7BITUUCLkSxCnWMw
pajZlDlPf+uWIMEWTDeSN+Z3UVwQEbq7HD8wGyoppmTe7wg7M2jGkBLoT4ef5I1k
9SOQNbLnZamqXFGnV1ontrk1J0/Vs2yfD6d97avWGSjX94qnDCwdo6y2eWj27/H6
UeJDngHe0a/tk0bi4abc9IRaZMlbA0AfUUUEonXUmXkUzJHJQZjzrnT0tkiWNo5y
q9Nn485znd86827HzDjZQvNVyUr8wHfBcsoiw89OEPk/eaZL24k7UMzC5UMwnpcp
5YGi3BClZbknv/BHGDiTyWdeSY5/x4HYywbwovmrc0uI1ctf5UTd6xA9INHujHiv
efNa2fBqwv6raBdurrLMTcvzeymy8m2lwKtEoDAh7PGzCKBDUWoKKDLv9u3Bat7q
/7i6vQK/riSuz/pJ6gsTqfSLNDERqypBBbfFK5VY/tr4pfRpoifRRcjmNDtkbmKA
zlT2HDmksIZSzcztHczBksh0c9NV2aJ3xCV8hv5wj9kb5O2jzILg2UyDUWykpBca
2jpNUjcnoKV2FKgY2NDCLNLbhcw8j/xKMbY4Ab/EdDOCXDViNsasj3XRXNHqu75A
6fSA+2hJ+OfoK3eaXLYPL7tn3obIvMPRIPKJafLPtV2rAkEdAFlPlsB4FUHV0HEU
tkGuSnqWLaynn4uBccKqcj6506AUcRNKBuz7BHxy13ENm0LGI6GeGLDR7bzHYfX6
IcP2AlT2AAYEfrUWycmfQONZMV42OI0v4gKZ4fqrjhCcw5gs/hJtuBzNTbJ7f4hr
1yrXALHDtBjF0u9BG4P4JzLtkD+22LGcnmtOWGyb7Lv4K70QgrBL72lNMDpsRX0t
Oar3oJQ2LohKtO0//PzzWVZe8is23Jj8O2J/PLEI3x5s6e3XidTrSXqCTWYFImVO
7tuAjbDzXvy5z34q2Rum3rTPtsIKr1JNwH4JSvCivxG4BT9I9aTOOH73SQhGPoJE
8CLfWedCI3jfpvw/RYb/3c2mwUPdf/rEmtWl5YAP2HOzx8Z+pqtm4xo1kZVg2jGw
BCyc2dYKjua9JOC8e/LkehERgSQdGo7O07T/nQA24WSxua/80gT/r16JOE+qwFt7
PaiqPLHpxh4bVmfoyGXidb+2Rv3qsYy3xvVCz2nQGUu7ZP2IO4BHFvIlSu2HqHpH
ZxGsedtgrmMYcfuWBpUXiawjBBy0QqmBFIg0HqRiVZqG8IrHSfJT7WUkTHjkgsU0
Vqzro7R/rBZjKd46R7Ph/oU4mBPQ/dx6g1o6VqNmcLgR5UZHzJjzN4A2QLQltppU
dQW+LtFKo79p5eHCGdWEvn1fqEC95Dt9tzljp1/SuasJQrpvbuMFFxrLkANPh5dH
X2p8qaFNQ/3tYhtCMULdDAYNeZYwh44heARbkGSwE4L9hUhDG6HWXcXbfkIUEk0n
t6uB4IiB6WGvX6H6SpaGDOSYI4S18baI3CMKFM++yYoT7qOCYR0rg3vMPQbV0oSO
QwS7rW66XvYTct+nXtoNvbZ5PHLZKNaLtFpRA+hJu639OWxMN3LboxFxX9ik0z+R
1nWOEQ9BsjHWEQmKZQ9sRaY90y/SQPuq6KHO/cuSCkVcI/BtBgtspnjepUHM6v4d
Q+kWg5szkPqAphqMSk9R4bWQ1Up7il47loaD7LEJXavpAbHCFb084d5D81IsR7jG
rNSUMpOpEvW2iYDL0rVZJbhxXxzY9pz47xN08o8Qj8f4woi6MKDHfdvxCLwmQUYH
xNkmKxTds/paelRkx61MCOcsrN7S2iaITpyxrswdOuRgTnRrypUnPwRNS9syb8X/
koR2MgKU9p9Lg1U7CVn6X551n1w6U3RLdiRhqqcH011iBZzolVHDJxtez6jKq2HC
W1J56cnml+gI6AeHbCjdMiPUP78MHV1w3ylnibXNl9JE7YBV+t0129FN6/jsDQG+
Ynic3SrkeuYSX38iMrgjkblVG0OFtJVQ0hPr3FRUyI7qdCyEEV7UOn9rZwX9KGR5
J81EbzwmZhnQYMcp+Qdq5Z3xGjelT/iszQM2WEjr4G5uxq9ixg9Vxoe4qVxuPx4k
w47thoeCPG/vBH5aDM+n05W3vQokl6UrX9VBoufFXpwr+SPMED/QPuYaYxDqStwP
KLMAoTZQGoVuorcGW0YeI4uwOcNXb7UBxZ8lMVvaKZpBtUHG9cq8gnXBvmgDgSBE
2/PjxNQHaMmkXySzpsUTytYCzf2Cxwq3+GZwPgrqWrAhMxg19qKK/mrVOm/5ApEQ
lBMG2XJ/613YKhoZMBkKzmJBXc7NE1DqtZR/UPq0Wyn/0TsMgxfRU/3HgCB2RJu3
TE4sbf5ZOKFUtYgWFYdU7UtlGm/0evSmaf6VIKlYAPu37Zy91DkHyKI0zYBG41+/
PR119PpUBpSZQ6VsG1P2fH+KqnR+y+uPao8x1S7b1qCTF5AigO+L7O8SRjLgqNCa
W0/pvqHkWXevJ+7Vy4ymvt1URYxtlcmb11geKihNvEhKR8eNxj8VyECwdvy44cz8
UbHEdgUHkr2LqZDAlc1jXgQ59paPaeT1w2kLSJ3XYp88EGYTsYW3mTCYn9X09T/H
zTPEWikiYrQSfFUjaQOYnSkCmskCoxSZmpfox0yD6/DXVRHQou/WCbKKt3XWdeHL
LBgQ+c6pef1SeAQ0ngTZG3v3hKn5S0FvNZNzfWgjbFcnttOxndEN22XpCWrORuXk
QfWfq3xcuSK4AeOINsFDdhDFLHHkGFsEzrIZ/eKNydSzlNhcNnL7BicPTlNl8hQL
Dv4Pw/Ik2ej65aLAgbsb3HJiViQuywk1WZ1YraQi4iC2smw5nyp+LYvSpiFuiY1n
pFE/zBFhYiujXL6v+yKSrQsHkhSwC+R7vaQsTIr9PVkN5RRYC/CZo6pU5Ho73mvE
ioHJM66E2fTRhkCVyNhmJdFGDxBf4S6QQ0ig7FsDcnK+ppyaTV/qWtumrzaWM+A/
oWTFFLg3++W+Vnni3+/4ACxeHMrvO8fmTN/pmJbklVqhB9qgrzWphKzQUf284CaC
TJuBZUjdVWkz2YWln3dFF/fFuRmV0k6gSCTRUSALobDYWHuczJz0QkY43mybZgK/
f4o1POy8ccOf4qcsggjxaZZQcqFgF2LrsMKukwp2mEE1cyYL5Z+QYVNpyL86QkLt
RD6N8vvk/sRtajOKpt/fIFD9mpsCXogPIqAyNsrAHRHyEjBIKMh4e3VzKXKJdP5k
OgOtf1yUcgeltTXeGxrvPKc9GoJr6IZtt8EH+DmaaPQ3jlUES0zu6z3mJ3y6LJD8
VtLy1Jv0BmE+isjsn58GDrvJuXm3VEM9CGKq1tzMM76pFz4ZLRlRiTRpRH+0GRfQ
6bmoA0h933Eob9FKatt3T0bIqL0Y8wHwV1HjcCQ3ELTQ9EPAuint2XMYguuds97y
SpU5uTn5LhUnhMCa7FuU9wKvjfuHzQsjaAkYZ65TIJHKCULWSmWan1gY/eAoj+DT
P3tHiOhnN80mPprL0/MEhANII15xGoQCFN3ObqK30Jc+vmZZ8vDIvygjXbsv4YB/
WRraHoKmRkugDMjFfdWmwM78LTkmumQIbej63iURvqn7TLwidP/8gN+8lOBGk/Ro
L2lr6+Cs9ZeasmivYgQqjozriS4pTW13jIWu/WdCBQGeWDNy+k0eK8tHXdqN2RSB
ib08Rugj6t/HGKVFfUMBzsfLSrO8X/Ak5ptFosOBKKvwsAne3DQ12LaxVs0r9Hd7
zvIiSPa+V0gLx/HHmYVW5J2AK4cO+kes7Ee4MUVv0mwA7kwffWBep03bgn84RHBF
YrebI2rk0WBB3YVKNfY2Ew6tKKWprnwZTrszJELcfnm9ZtdM1XeZwU/omCIpQaoP
J2F3vXHIb0ZZZ0oJw9LbjeOCgUo8KLceNG/Y2ybSTgXj4+5UPA6fW970nnGEvLex
J6vPQyK2C+DrSp6138TUd+70VDfkbh7nz6n5IO6AAvEplTbj07eIhdDjtWYQbHwR
SVSj60ntkueU1Pcez+OrhTo6DdkJX79GLhaPE2pK2T6l+7Pc6TDdYQ1y+8jJpTMg
nlLJt2mKnyntUGWWPY/amxZo0JulH/sGQEbczw95CJjPsUPm5CFrnH6tz2QqAqsX
Trfz2tK6w+XXG3Nx1kvj15idLxf4yvu1aHbPDi04j37Jk5q3nCoNRG2hH/oXD28K
uFfFDRF1HtzJN0WUbO1k1eK5VepS+oCqD5osgQs+lzoPxKvqvD0ZCUtLnvceUTp7
a+yZgUeihKlNbgMM2JoPJX7eCQNouCYmQE4WECiDI8nnPHpwkl1LeQ9jpkOai4b3
We4PZRUNKBuZmKdrSwYP1ztxWGRjjLTldt8SDoc/Y+uSiaav9DDDgiVfO5vzwzw8
CYf57FWJThKmFOycmG5GtBOTR6X+c431jc2LMYIlnNtCzoqMqbcddoTWRA3RGvvz
YdsL3peOj9uOpIZnMympayz47h+D3EptX9n0X4Yl9nDqHXjeUIjYlbNyL6YTdxUy
jyzMn3n/qwYbZBQVTpHOqXH3rNgtuBqzg9CCltAtgltIbd4YGQytWTM/sTPJMRum
eiB9EZDOgWnMhj1WmEtyn05BRTuSNFak8et6QGNzuM/6jbF6SKnWvHneGjR3COop
UtjLHEari0d01uO6yqeECBVBQ6TRLM5DfLZN1Jq0pC0UKnNRbABCCxM1DcZu0M8I
MDpV9c+IVP4w8BsIzulUs40S7kBvUCAaQCD4QN0jdvQwWDcwFR7PlWyphnFcqc7Q
PIjH/IaLjr4crxVazoXVzz1iJgGxsKwCtVtfVqW3J6trv08AZIaeV4o4Kla3mXre
fQVaNCxcEGmNrPJkv5rgTtZd7kQdxJgQLeXox+Jb+Y3eej4ngBBYcmJZK9t5VVjt
NU96fUZbe3Wl+DxBZcoO0vErQFBOUrtY+iSuJVnwdqsx6+slkWibsfwYUt7nQAmu
GG4aalhGuozxOnnwAraKlLd05m/mBjtzgGHMS9AN9R5N/AFPW4rObuVq3Au2Ybkw
zzZj3dEBWonDJeThReDwVkDIGl6YehJc1jO/fbSUm2QfOz2d3/9Xkp4STi0ilPDN
Pkeb0I5iw2YIbubFBC4ufLhXNdVW2Gkzc1IdY2cSPMq9BT07iFFs4HV4cRl5gDWF
imiAdApuSGUbR93i3SkSckwNeuRTgFbPW4PQqnKbznO1Xi6w3HLBupJVlFAi+z2I
kJJP/7fmAAVCvDHaKBRCUkMcD8jxsIv6Zq51Or9Y7UOysdaXBGgpHmpmGTgWjzZq
mu+wgHmaBAM6veFABUXjQbgEyuV8cTfYmBp7OvqCDpsSizDLAnOlHyOuKlTotJAW
KmKoodq7Bmm2jte+yPgZqY6rnXY+tIQZ4Uz/F3pRQhHeFckP30H0vopuNkrDevQx
wIG9AZTIVEnp6DhqHyVCELXWd/2ZvZ2ZkoZabCmrSiqJQUiN0ERI9Jz7Ckviawyr
oelGR7nGIA9Z96g/2XoI0P0PqNGHrvu3TiZSwtMUJnQi57n4MVFmSOpohGHYCbN1
hFMufNeYqV7XNWzRXrcdjFvRBx6N/FIsDtgs4knk4wmg/rx3HcssYl/sMyiPvSeo
8T1JfA1o3ra9pZMQx4DopKH2n3aZ33F0L+J81kZTQQvfEBIeeZDF7dyzyXl7jvRj
2WIHM1QdU8AaxBiTMbdkbSI4utd4TYL/6JCl0a5MF2G9Af/9sKknFVCm3KE/0Eb0
shb253rlSt+BTajqOvj+KK9a+GrJz35dN+XsojguHAqyMMGNvIXpVop4DxaJrI9k
QDWsjdvzQuFeONp8w6ipNaK7m+zsZrAy4Idnfr+DGliXPkkbe462aiQvQxrQRIUI
uHljTnQnRM/EyQb/jc/Iss/ypCPfIWzSsH5+zXVpcx2ZdV+70yGlRCpS03zWx6r9
q62tBKxD/wmK/g1AcVPhV65KFecp4/neMuTKbZ6GYySLKsIachvDPiDV3pilARUo
btlaCLcG4YhR1pneqicA19QyCwDhev/ohuFcBcEqTuFvA5Zq4alSVKkMODh+clh9
LTPNw0LJCl5v4vhZ/hNHrNvIIqsJbYzv7tOSCv2XpkwiNSRpYko1o5LI8Lyk2r5a
k1K/w7kyfgShxRkbpYmTWhFN0eg2CvVFvcp5kYqvkIYhADmRteIxSA6a+Cr/Lg+u
JqeF+wBclnjGdrddO+Qw6AZhOVGzs5R6rJSha9myRhtmE8RdnOG1mdG98uNGKhTf
gFPdf3QPNc8W0fQxi0uhA2Ha3ApAcEfWVZC96Bp7uyBm2g6ejzPtO4QNWaDnVjFF
Urr3iPnx3znP/1gUA5FpKe7dQy9vLT4uUNzJj/OD9UcMbV27X01UouwwUpAY3s8S
RlQkOBRi5QQbvf/phm1P6nd8QP3iif4NLsOpo1d4IIYGn3BzLtsMiz/mDA3BZU4c
pgl2isrnUAVMAfbH6csbrpYg4pDsi+o9XEMbvgOY3M8irDADkOgLFBdBt1WEh8hb
OH2MQ/EvyFd7syiwDYUgIiJVFTxS4MclFjKX9MDG0isDejxha2NjT5yu5LukPLtm
OwjjfEULqnNZY/u9mwuwnO/ILvpES50a+GxGzAMEVulfiTvme/vrOfD17iyzbyYf
3WqAPQSO9fg0/7ijsD4e/APULEdtVQnjMI/wwDK5uD6VELzyJMqIEx/iMcBUGKes
FrtebnSBrePAxL82jWF5XbUeVXoMlXoXyacqNBNv9yoFSbQj0Doev1Pjqc81Bc3R
e0v5e1ZNUMGe9KGS+UhZ5mPH8CLE40PpBA0CduOEyR6q3RY6x8zcKMSNswbUvmiE
QGaucMz525XkqrgyRzrnkcVmFJ4KCY/1FvpDUI5PVKEEqhqfqmqcn3vyOazJp/0I
avVcvU56yXZE8yjhu2/qAlCus1SB9Fj9Aan2s5Wg3lsSjyMwfiSLm1R+C8SmneAM
5y+clEu1++/2WJhHjkUIWhF5gy0ECqJpCokmqDIeMKZcqn9dWNEGXoi93t24aUmN
ldqQ4U1fYw9m5R+xG0WEivf0Wtv547JeIXnGp/XbGpm2f7S5f29AJQ2OPcwCeTuq
1/dFHNziECOMUWeUsoh9+QXZGtI2TwMmGEOeQxnxEK+4XHruY2m/33kzHbmyH1tF
5IdQqjRbHMney8/fHYmJUhBC14aDmFGdBiso+mos7bt6c89HyEN9aGcd7sC9D5fA
zHIX4l7Df8fPeAgN7kDO5yD/6x4KNRlOjGhk3wNATE92ekpCNG1Fv+g7g2FPuz8Q
AynNQgQQF2hZuuLjs5rQ6qVAeHsLnMewfsmOAs+XCTZ97y3PLa5Ad8TJmd9oN+FY
8Pr9KuLtHSuNWjdrgCtpDp1k3SHVm0FJaW8lb4zPEthqaj8qVWskkotQ19HhiJcp
qCw8B02UZoDskhXXKa+AEW6r8WIw1DxbOgFs/Ar/7uzumext03aTkikRKO3/U38x
WjBMkevF9DZ3mXkGQOQgxBGh46ks92eLMRYoSJeXi/dzDcAmtbmwJLJD0UpbaHpE
WgTWpVcGw5SBQLuN31GdZPOj6xaN9pc9lYPjKJ6l+pRFv7V99llWKMKLBYXVzFJR
HkTAubAf90FHN4GH9TJIKilQQaKVUYo+Z+mP/ssBh+x3LwMeg32jes6+VkzNYIjE
KUTPrGxH2B+lG6qECJh2fKrKaVKmogcn0d4A60FrmeSnxUmonr+P+H3uLiBsmTH5
6JQLj8581P3LzT8Z7FuZSZKZtSUV85qasU1yZ/asAc7ax9uWCAVdPZB4S1UDbgxN
sAu5/udZljyrizvQvq2hRytGO4HYBtdHiY4NXuz1L4fD7AfPXrAJIxgWN7nb5p9A
uFV4NSvMXJD1FHAIXW3YsMqjVg0kEtggSFEguF3y37M26FRCJWMp66bSOcBVLy0j
bMnZ6j4chT2PvQTmmMlYksmKrAy0bJ7glhaN+eHW2ZMS6YJc0d4xYilcRDLgUPE5
6PyYltgnaTsynuOg/Fq0FIE7KsR+/yPkDkY1MFB4uPru/fyre0nrVxs046Xgv+BE
q+GIwgOXiaLsOGYd3DM5OjfjnZrjynSQETugI7v95MD+yXIfoRDT3p9euSI0Nd7y
okBCMM2FGtCgIDc/M9v5kyt3pbcR4Jv8gMQsTEML0EdWkwSKeI0SLHg7dMkL34uB
zMul20p6AquL3kSyRpgDrsS4I6MHbbAwLyBeOmIHEC54itaQAvd0ANoCiOKAN+GB
SUL2yGbye+8XnItUS/Y64rPDlN8LWH6SPxOIvooO3MpK4py2HHLWTc4cKDf2cD1k
eik18O9wC3iMO0OYE0o6C2oSE2E+1mpGSVsouombv4dHcqjwVlWhQtK2BITw0S/l
8jzTETKoKLzeAXNaUvU6SgwvsrKdxVgjKfhOWCKc919PTGxeKQce+yXN0TdkAMrq
heBCpAUQNMA1f+k3qQWWDjCkfamqAAZUirdWviCknwXQiUXW25N0x+S7FV8UJC6G
p7/LFhEMM/LrY+488PXZZO5vsaKOktfVYtzlRF7gr/CkCQsVPyigdIofU2tGdi5A
oBLpkf5BpDKIjUDUc+2JoRMwZt6zzhFuJlSG8l7mVA5I41mxu17rCNiTEaNJxls9
KCCfSbSWbYVQoKmtyp558VbMmGxDUL4W/1/Zt8ddZL52h4F+DfX5eBMxb2HFqXRl
AYFUFEApgYb7XjOqcT9x9rqx7ulD66WAKhI5cRpiNeFlxk5f65+W4DgIvJ42nr1T
ysVTHzgGfimBRpmV46SkvUPs/2HH+T5lRyTdKVqltHTkUVYEFTBrN5+X3bveFQrY
bWcHGMfXpflfMnCvy1c3yyuKQTnRlICdUTsOdDxQttVVw/KW05mta1KS6DKrz1qi
9OkIu/PDxPH2he2r24hXgD05UG/WHubTefqO6hvN3tKVwyUtOh2oU+i/kfYEuhEy
v1IID/iMsU/+G3wRpp73Z5//kcCUET+bjqLeHKsK9gjB2NOCy+QZ9hLUiV0AAxTO
iHvzvwkGOXG57Ga6nRYq0iq+0OiIrJgzKRDl70Yfv1tSYMoAMaff4wRRNRJHIFeW
8fFD5XdRtoGPCl10diPI7qrJoYMU6gTkAxzOYJwEtSZ7p+kVGUzq0XqmZNhuCkBu
7fA4BiKGtj1zoPumO7zRqR4ak9XS1ZIHatHCbG3XVoS8+Ic+BFZursWVSCru8l+P
COwBQaalroqcoZmDCgfXATCvKkqGPb/q+YqzJEotteprJSbe2SU6DocciYpnFeo+
a7Xc9XulLpsuvdfqLfOzby0996Z9lMpS7INHFbDdju0/ParkbxlR2fK+CaBihoh0
285ZPSUxezfOiuKJLlt+70hFAXrwLJtQXQmOJg08XRVX714CIVkrn/P9Ie4QEEew
C7EG+grhMgaRa+PMGzxdzQpX2Y8m4W748C/tK3PtLiAk5+lxAzvC6opfipvYICDL
X5MAX0petm43ffnd1R8P3Z3JCf86myaRYbChsvEtlH/1FsrH2OnUEJIxUcxy2RcV
uGVRtH2NKmfB8ZunHgxPRfUCCr+KhdNqytRyp5+IPYMZUgs00p6W974PZOcXyOjd
s90gs8AkoftXVjFKUI7ztHMpmd9ALv35tzyhckK2aRRE9VuiKynpriJp0iWpEoW4
N+zE1qPdFDWybzZDulbd5g0i1HtSGUAMxJ2NFH65idgutM/4wcXFm1FIDbu7nEt7
f1X9zSYDxwQV2QXiAS3/42tIxiuYmQyqMXoVGgej37K/W822qyLxhgV5d0PS4nAW
GtfpWFeFLs7YO2a3j7ogSok926FDHdM5ZjnXIsIqyDnjW0zbtgphSnLUyDAgKbq4
RuIdc8XgG/wbzWKTuc7CnYlTNw+x204hzwU+RFM47Mct8qd58LiG4t9Ey9e/qVjQ
qW+DusCFHEiKEQtatoW/SfN7xmf4eSsau7B5OVgLnDwUw7Yzmyg3ca69d5Y7gUW7
Aq8cjX0RVyNErE7wSy6gtxqXHHp+kIM3QegV9+Pk0HagFLJfdKb1B5jMpL9Po9SP
RxMgBeQZHuuRaMXce6rPXMaT0lMROCH2onEZPue3SqeeoHOGMXTjF9ms95mrOTGX
BIodWNAo3A28KjnwieSsxXB6sLjfIvnjeQr1NUTlS68ODI0hZp+dz7ejEO1U8yqz
yVxQtKQb1aDJBvtlgOWpbvZjV3WGljTdYCXL2rRWsLZF6qxDd7QRFZUWH85RE2oV
QN1WfbvHv/KN0OLcAqTefxzp3TTpHxypsL48AtMPJOHiizKwbSKjI9QF1ARbVjbf
qD+1sKu4903ZBwXz8tLj9BlTxXWvQQf98hOyvX0wF5XD7Gpa8X23MIwh7hJME6gX
WfHF2goNHlGsHUcAvkO2U1kfvbAkEm+jBc6l/+pj2eNAJG8ICMAUwPFK5w9so3HI
upom3+oo0RPoD8nRMaqZdS3q7oyRm2S5bqd92ktR6qo1UY1RXw8gP39o5GTQPP8o
wrslLX0AH1Y7p83lgYzLxap1r2I3Be+Y4JpIOm5vFVNlEM1bVn+YOhAgIn1Ws6cf
S6pjFd5K4dKazXiVPhX6gLboDPZemdnmB8qoF7bJL1Ln/DJdNeheWPiId9VdLmg0
w3KuSijN7BvhzzxdCN+EpK4LYBJgi7ojJtBPbW/Q0Pu7adDYmxQxjTPOm0NiJB8r
3qpbT0WaGwee//LeMnOtrTAqRSopHO8fvCVqIWYq1LkW/0NHEIFyf6h6k4ooHarM
NCxqdIWJc0NFt7d1nbz4CCPPBrJVjZllrOSOEH0WmoJoDDQZS83uN0aJagRuPBHb
E95wLY10gy8C2KnxPBzPRJr0y2tl9lv3wmSQ1Ky+mXPgV+MXDGObiPNQEcPKME2Y
uQ8T9Y/5k5CuE0KAxkJewxlFvaGfg9r0gQ8nshiYNBHOcpnCgEjXTAOoSFKWUGik
LAnuXQvOYzv8nMNLVqTHlz1UToV7HH4uLx4lq/3UPLMAy+k8KRs8i4rMiAdUZilY
9IUy5cMxPsxQFj59uQbRY0F17QFxDipxtPNCOyNC8mMYZD3rO2FNCHaSAHxsYVZ2
pV/2gabSPkcx23QA/seA8Xbt/vLkqe5x4H3PiNywmmwi3LorN7rbUgwDtiIcJdYi
RgrMMuClMHmwthq9knV4/RLeCQv58pfrEzz0qP2ntT4CUWbvjagewyT0NtGSqEum
JNz34D8iAjMSDM+WFM15GaSUH9j6rvAcOyNuT0z3yAj2Vp6jy46Btk7P1u7ShHPJ
unV6J0uL/hUEJlKRU19M4PQsfCFKaCaz8342awY1TuCk78fDzks+w11AnrywtTF1
Djh3tBvoFBcxC8Z/qVW4Qw196KeGR8YwoRhfpu0GBbxdx1U6+aPB+HVQlvRN+s3o
gEws2czW5yoYlAFUF+Y5xygLgxU+jAdMrDl9OS07MeXF+hGpe1szHRlDBs2LURuv
QiS4BvZ98SS23fb2U1S/OXyYNCwSf1T7NoHAGEMbtfJCe2pDwwmg8Uot4PzRQwkM
oHLWOEIIBx5UkLB+Xk9chU5a3g8FUSIWhF+K/XbOpqNGo9rWu3dLKmIMfJwHeQMd
TZAVXFqsKisnYMefFRINqYJ2uRy19NOOHbDpc6Aq3ofphbNvx8UoKVdAgl2BXra7
a1FB3Qj3qaIw1UX99Fc7NjnkKQZl1Hyl24gBvt1KQv2Qq4JqHr3VKvUKiZLll2Wc
s28FrT1NPX2Gg3UQj4zSttN3u5wp4Q5MKNw3kJ7suibhmdJ/dwSTXEXaLW0tnWKV
sXaQd0/m3SoHKG3l/mh61DdC7gp1vPLpTfiJRMvi1v5fg9tAPkt6/yQUTHq7Sf3U
5Qdh3ufB8k0Q+hNsxZnTpgkjxk4/Bb+qkkSNQNlEt9+cX8tAh2U1tCr8E+Kny98h
azetzUZ5WdFcIwHGeBGTBoR9s1WeS7zaq6ZefRN5Ff9P73aamRo7rq179tVyK0k1
qtH2uL+NGojWU7quzj2u2e6SnaEL0RxF7BMBC2TMKJBHbEeXKejIwZ3BIJKFhccT
d/wt7cSai33smFuR4s86CY4awua1dlVg2z0L57VOkyELYgYid45uNyNDVP63DBQE
0v5xLD9qy7+wZh5e3k13pXFu5pR6jdFhADY3qzYtdxC6io5GPpvGF3JhgH35/CUv
YuxaP6LjMrZ4775kXKE9/NJJlMmPoZiINfB6zqu3AAWkNb2AaeGs291yteQRlt1D
YRLVupVf7KXhZcNYVwTfKiOByI5z/oc6ut3vJuUxCI0/WXbKBF4JpyRiKr9Fql7X
hbrYtBsfJfOhByMJW98qIpEZDX/ecY8k3OQoYXsG+YuSbN7YykvoMsfXj4Ki4VSZ
KDmGAt6w80PZjoLBQimLI+XEmLwKCr5ZQ9Av1SLsVwRC8wOikWPJNZgfGn+RlyzU
ifHUn/6b2CwgjqjnLqhCIEhYjGlzY9upiZa4Fu63Ies2kDdcsuGV4rxkcuQlntoI
2vMSChpbXKdT2ibhEBsui3UiqclUXvhiU7cDAMQSPBPuFwLbckR/2fqILG+HqKaN
L4PF9xyxR04ZQmNVNgi4WE7zC3JHOJiMOJcH2ZuOKbnQQ3TQlMMbUnRsg5i5+7ub
tZpb+Ghpk58zzuRpztxdiAvTGPjdnktxuzf1sis1kmGOKKr47OYz1hp2/bC1U+mx
bSDSkTxRqUN7XmOZyJ+2wWs1lbbcLlKx4LS/9Cd8a7bHGy+i3MduRLDge2DGYb/2
ugRbwupWpuab6g3IUp0EqCeR55BxuUqCF8XBD2Hrll8NwxHcnEPCDPgz8X46IOfB
hXVouYinF28tDsLaH3Q13IxF8f7gbk8Sh4IOouvfdPBmvqWSthcBz29J7Wxr4ih1
8KQiWgIZm1KzhbKtmLb/9tQ7W1Dd7bnw70ivR1/EckOhakppuKC/DWZu/yU13jS4
+LU+YkZk+KiRuZ9ptis68xpTx8MU2Yv1av499WFIUx1cPYwZFEHy8ayPxPQ/AK7N
oc9XS1xK3kVN1t4zdhTJVKiY7R9NtS1++MuYl/nHvZo+bs9QW4X2Trfa0pl/bkki
77t6NLQaPsxaq3a83ZVQGg+oeV4iL8qjg/ojmsH04evc+p6RsPregZWAnRmrrA8I
VWrer/1f3VEIbfmjONc64rCubiESS0mxTOkVItG99tLmT41vOZxCsg/5pQcyeTSn
vxcp0rECjrkVQ6IEWa/wbBNXRuhY8vWueOYpoIrj51FGEczJdSZH7w87EC6vQWK0
C+aJcIrpp6VAlJ01VKCKYSLegiulm/zUxQyl91l0Tvny8FQXEe2EiU9XVXHU4Lwt
kCLklxoZEoO5EVQz3zThtBePUZ9wGpFZrOGSIHWUOAPioGvE9giTjZ4VOAN1NgTJ
TPka3djp/YJeArqyA9/4udcaBDHkvk8+t+gk9zQk44esc61oDBrq8yQexQAgyOM6
lugHwI+BCjUyh6/hazMbx+3gDewEnjoI4MKUMNRxTU1HjrqIf+VeBdIseoiu5/ZP
vHozhmfCEufuA8Z9gBSRVHhPF912lRKLQtmQ5uVtG7T9xz16irdFurDUs47JwBDw
fxXOtmgNciKoVIhEEO9nHGCzmaQoLYv6fSkZK7p7ZqC7+5Fr6/JrViX8rMdJq0AS
oO7F4ZCkzvX9S4fafj3PT85XOWkKrefOf6p1g9hXmXakuhkTaZqwq9ffOdqKbE82
8dNbSdy06/6smOXHoLGONCNSXHiQxLefmBVMqljJyBANfRdEK00sr5ouQo5y2gYj
m45GxV6qNXzfFKMU/fFmOkC71nUbZv2ZvcAwNnOhuqoqa7bL8wl3Sw587loYPtaN
NdoYu74daznqPmaiN5oG9KsLZh4PcHFTAanPktwEaFixpmhg5nQopXU/PW8f5tej
NEbWpBBl63CTwGC1oXE/4gAe4RU6ebvUEUPx8r2tg+u/bACfSZBakGI89+uDHBpQ
GBDW4JKbFvVnj7pn9Jog1s5YCPK6QhxjAcPyXjNjMnLg4h1x3276MlMR0xN1ZZGP
2RmyN3t5/F+EbEyF1yWWIxcFvFS/JSkfhLrxqIiwan+nWHKjKEmxXFZzYCXsiWjL
vvAdBE37oWRR8e9H0dj+Q75sXqxcYrJU6Nt4/HC/T3PC2y4OSIDmIcxDA1d+InSo
VK6Lavr/kWU17k990JtWagl3T275wetAnxA8xb9fvGtKPO+xVUODERY8kiufGori
jLUL8Y7yFZI99P1TNveucAUCSAec+IfP8sg1MhsJgsIYgEhFV7qlcmJWRIrudacg
UzxfG0d7n2fjHblyFj55HBF6G8jByCOIM0+S2fhDrOeJ9Ov1ZDUqgBpjjsbQkwFK
TU0aIwaEfsfPX+xuDwuRurY+pitmvMLqux7MFvSozN0gIq8jZmz4FM2a76v37LYW
LbgSNJBaf1E9N+KAr442H4lFyf+jIvXkhPZR5bXeWtJQfiD6u7uKcAq1oxkxpK/v
GRDBoAZQmpfmiMKh0YaHwl0ns4uE/o+TPHhvBVb/uJiuV2ON2V/HHG9bCmhFZPJv
IKqpzZug9n5hplE3SvwcGQvimqGpS1nn9c96MFDLL4HpMIW664xWk3DmlrCYvD8r
j7MeXax4UCufCdXUJJRD7acDPhc60M2HvvQVdNIZ4B0KYBVNpRKGQ7hlAabybYAX
gIJZCvzKvK6gyzPii/60Zq6x9HnmOmMdsMNSagyHV4vvYtfg2CuSGDzYYBO2xKzb
jWR2JHM7I+Cccw6J6WyI3Uy9foLTA5uFCsRUwGBrb+S59p3x61QjGo6GIHlBCxpG
syMejaUO+SN34Qg0RZ0OwMXLVQnynGwbbL22VInynucQfuSh68nhBUIvXRqeERNE
ueG2y9p3zeQGNaEzzQW3eTSQmd5UWEDGJUxTTcH7UoFJIqu3rw4fMeUWE0Zin/Cr
UZxLggouKBN/IGYVbPXJOfwDqW3bsM8VBkzcRhLMZqo6NMPCmh4T4RQzb5oLikrc
vdSK3FwRtrzIGUSAbFLd9fbeDwOc346yjR39G6uCIP9bcjd++R2jG932p/Jxh8Fe
QeGuaGT3Fbgb3cscARI//znMPp2bNAmbdv33x7fnOEsft+gu7y04M/lBVHxQ1oXr
gloDsmfWRxFH0EotwnJW1SzlSxSUdYdeW2am4cAH91f01wMDgphhC5YgSJTOlgK+
xWItYELWZXSL0buPiVfj3HXyDry6qDIBPa/pla+5gocAyMzWPOOSNwmN6GdNBFaz
Bbt1Q0tvIx7Bw9honcN4QSLxYMBRRp+J6TeH9peL+Gp4jY3CvOjiXaDpWQzxUR2J
D7wlxLP5GwmikFbm73dlJD739Tr0Z2viAHSCjTQM0ldPQ/vlNqVyV8/YFoVXypIU
slIqHkMaPF01fjE0gdZCnjHqMrChh94qLMheozYeMvwWclZ+iXHzPUKGfpK6TiCf
++bowyKsgyj1C0JYbgF2sy2lvpmeo5uLz6a+IPl4OJR1QOnMxdSz8ICyIV2zipKz
UNLe3GNxJNNhi0GHJyjmkEeUFamZHOXn4fDW2XcMWLlL1rSrlAPQCVVXiVPK29Ol
ogZOlOErgYDgVLcKTop/uFiIKuSFGxy8HfLM9TxHMiMUPfUepcGMzgzp8G4U94x5
o/b88R+wCk4w+LzY3PDVv1tVT5YyRtOjsFJvCZ2WJWaTXFHshAfBnLcmCOC5+eg3
U0yornYjYscvJVz5mmKA5GOaqoq33xXsZ4V2m7M9fMY3aa6VVuEtu+jHRqFU4XNj
EIXAYE7BjpIgfsOt4tEB7i3w7uT3xmzbd7PJksGaGgnqyDT6Fa6khXmplfi0Rhua
1Ndsk3lzcpnJVfOn9RMorcVP9geEbAH1aNtf5baC0eLIAcL5NAKuksZNXc3jOT98
TBxj7QyQsledeq4BiuFhOcx9FmNq1ohahwukgcVLptBaAFgYKgxbx+eVONFokraj
6UqGxBO72CrHPb+Gs4VymbV9hQvBc/Brq5K+hkil1gyI8gHshmQAhJHb4+izIqly
dh5hpHyUY8pR7irTP1Ykcdx0LdxHVcAqK0Xu9+uekmWlZhRgTzGOVS2ctxTq9duc
TGn9YZfIgHhUj27krskDeJFV6F4JXVTHdTYYg+auaNBzEWR0A9NrZI15UqhsepW1
mSgm1BSJV9ByFZ/U//9mcJSMVdSR43b4E2qYsXm5h1U7V2K0Hc/hcLcb4Tr1TfOp
Wfy8391GP5C5iuiDr7sOF/iq5+GGyzluudtQQxeu/VmhdnLrPT00j0QGungvibn4
lb0mo+BIzBdjKyV7V35IKMeqc7qGOjQ+zI0VDz0a7j+LrUXCvDMUu2YwLmneG6+6
fsEyZoG+53qXbnUyrLrPmkHVPMeajoV3OJBB0M+NubNU46VjKbg/uCfYjfmB486y
GLMn7Us4liDcCyjD6KHXrjB4+IcJnTs0kMsNusWN3QrMsMgwk0dV89g38GlRUg+e
PN0UrW3bIfugcYrSJ1E1/5gbu4sUm8F5Y8Pn//uTKXFNeMdhkyidHPLQUSH9382C
UJvit66x5TBF303OBgqWeQAmGXAC1/QUDWBM9l4RfR+1u63HB8oF4mQSdn9Hwltv
8Xzl9Ykv9apQbfaiMGU5Gm8ABjIXQB2jXFFZO0ICKnUUEObXAsl+5tqhT6urSTm5
kOzij9fcVCYdeC6mWvWw2hSi0q5J8ftlvFT9BkoSufNtNYL6NFvSsqwf8JzriUmP
FMajjY5RlH//lON0w2Efd+jC/N7vy0SeEUnlU6GJxP5Xi4Neg1KeMWt6FJdkRdce
YkW/RAz4F5CtvS5vJFXyrAU2L01uaEw6tbKm5d8AMazWDX6AvEi6x+KR/OqoMDeJ
fg99S1Nui+DvGY0oFEqLMGhFhSPQwIux7DLWGjmR2EfCU8V1HVTHHJ5CvAJZOsbY
xi3BNNXgoxwSIlZwGFflh+cTpaHmuLl7L3Kqn6pwMK4BzzQgG15AoMDZCDRgXNsw
Zwoj8DXZ+2kxRVoVsNcdiGGOjzdWkK4ytEt/fDSyXdVaJNO8DTaNlQDis9D6qnn0
jQw3ZHAyH6iP8/MQv8ouNpni1pUBfRcAmMG1V2H8uJRkEldSQYSYWlIKCbCsuNj1
5ZGCQEiCghcuOzdBzHVWF3Tq4+e/+kVaq4dPGNiib45YzNjkoTNiP0Kzu3QuJjUV
/TrkkJ+wy8Ge525+LOqQlLGGc/JfkPovRoUyxB0pfkRQs/qgUO0+tPEMWiGEAsWK
gbDpdwyHAIVWbR3m7ozUPLS0UuGct0kxg3/YZfmb8wbb8tFEhuwk1/iSSxh7t3Av
K3gGHs7uvFw/QszincR5LaBrA0yt7yiHrLOuWZTDHBfVsla6+es6nSw2iiUSrCEk
fxGUkkvOhWjVww03Za5Zd8arlRYBqFF5Q6uF3lZwVNzPTnMMqQO1tRaZC+/qwwcH
uJK+8skDaKoH1qt8kTh2chMPmiuXP1zfIkB8UqFWM3RDIn7l+Nsf72eKo2fawpTE
4eIVMtAExv6yK4yPDBmNVd1djY0dvwajYayCf/U2g9HqnKvlgAk8azz7v/lmwHoN
3eV1iKf6FzAIc/dHqPczY+FiE1h5MwdCMPn3GuFRCD0N/DD183Qmef+j0pBP7KOc
rzMmfh68L/tXoRLCV8WaJx1HenbJreK3wMPp3XltOcHELQbh86/70FBjPz3HosOj
ev0lky6tuuPFd+NYeO8bNAZ2e2KRXu4/w5/MLEmUl7RZEV26SaGAjNGGPg8I/fEi
V/SZLeTNfXN3jE8AMJJQ+nJJnpyoE9PW/VpAFTlRokzalttI/pp7EYyTmJGNpz5u
IxEMIF1rBiHGoOUfnFGz3GZmhrZ44/WYWUQu0msWeGdFZpKQA9jtLZ0CXbA676dC
HKjfXqT53hC8OrGDw2MM81r+cLbAVUN1O9fnA0YBD/SW/7Sx9bqkq+qSETzzQfOS
gCDunE+DLRLj4gRFZwV8x5JzOhdSAqwtH1M1knt7SNS+vknN7+faXCHRJU/wJvrA
U6QgAuab/okpSLgA6ss/lcOpzp1z8EfYeVj1QlDF6U/gNuw6snYXWIgnXEGu4xoD
UjmEQ8yLI31pEKu3x5k8FMhaD6sG4eNdDj9RLjdvCVPFeI5dzzeFXpPXwsiNl+Rl
0hKjELhoPvtJ2lD61b3xBz+4RC474qisHs1EWGlsPJkDlq7e1egi4MU1kIS0gP7R
VhXhSdtKMjiWvGoVGp9lr7lvXYCmqBhGijxwkx4fXfNHefZMqNrv62vAfJpZMMj8
UgMbUHcVNkG9fMh+qRd7/6FO53WoO98wBafZtoFaIrfuNoOeDOfYfA41v5ohQXCI
GvfKmDOpDTKeLc8xemr7/FE1BKf/wsd/zSXtAAReB5+eKIZtl0H/aQ7JUdjk44bd
VNyhdRDBiSNajQE3U9Q98TBhyjcsFxGvBbY9ZPPt3tweTtYxjD/M0wlrvpeJ+P8b
YQgO5HHU8LXbp0jjuf+qNfD7ymgSJ4h4s0qdF91EOFIlRjoa5n+oylEJn+BczOcH
6zzeAKU2UHg+gDA0sk3O93GgEfyjXKU04u/bw+UUrpxhCM1MQsYLt+eJMDRPLpfy
bsOettqjN1eye+NGxkqTOkbkOLqSoPJS2POwzHuLVkk9q5bJHsk8HgUJahz/hGzL
0deoqOPGXvJcaTIqVWRRbblI502cFxoWHOTzEh+e4YADbS5lrX/wzN4QVdNT3c9p
Yf0sQQVGK2yyKhe/eo9rcr9C72cIOjOtQqebfhGj9KkO2tvv+nau+0AObEwBAd5j
CW1Vq2rsIK4muxueop7pCYX6u+PA53YPRjt4fAjMXQbY68OVybbZukaShDBEzZvy
6A7HwYdphA/zC6fX5lN1n7fdgdhaLae8yXVGIIDPCKWvylzJvCdV1377Kk2mcBFQ
pTNNFuToKIkuT47C6x4OBa4bmEMXNrdyILktOBZG+pRWL+SRws35kJhkdV62WBme
kjv/RymAbfkGVQqruTTbciUVG0jeTF+kmhNvAsO0zGiscpgHgS9Hh1FkmwDxLMz7
8Ey6Sa3i9onfZyWOQL5R5j7wBJE4REl5gEFYLSirqKbXgD5ApT/9bINl+tP7LW0F
jPv8PmzKOXQ85ExKaAWD9iM//qaQvy+EPD+uEFeQVS3c4VV65z//IfSn0VGba4Ss
vHXydAq3UYSQBvf8GdHNM5/fxPAm3KKdwtnwOqm6kZPfOW2CzZRw8VAJlF4SHfNO
mmIrHsJMrYHI1gRWG8GBOvIb3r24YJaJ6YXfb3LaznHONYmbAZv+0O7hXC/xiIUj
aP7MGO+0wtURGPNOqMp++3ek76WDtgZ0gzgMWY+WQiTlLwZHdIqG3jJqhJdr/Ta1
wcMiTygEW4l6RRCYkzKlkgTtICQ4zgu9nx1Blo+Jj0w0ldGOltJL2dpdxAKj5N1g
4joWAKXl26+Qu4Kpop/jpptljHaV0HI1RgJxWuS/xZqhZ2jUekMy4LsfBd2GKJf9
NSD7p6sjEfeZ8iSrQcF//3m47jA1PBblyBmdh5mVvNdIE6NZ9VWQW9OjmksywYKK
QxiFEv/Y0X828L09yRCwCry8gBBOBY+P+SxBBmGj+dzlEyleE1INY4iEs06CwFOT
La16AYkLteMhhdDEb+2qaztMlKtFJbB9PoI0ufkFrTIpIA37rCWDIB+IYhnjVvDW
mXsFmCP4MnDYt7hwBQb/mVW5JMGTUvqM2A/TVbTG8WZ0q7l/6PG30ihE+G06v78T
4NIuYZyWuTRKfQElNHWXM2+8Dd8w9KcaAwaskWK0ZCpzqv7tB/sr02aHR0H9QyCe
1Oa4OcJOHuuCVjr/CE0AxquZgYaffv23hBoIgX2Rm4LVdRyHfgMEWujp4ffiO9O4
l4coD6EXB29HK8NaFybMAA6h1yegmBooDpyjKrP5VnI6R6PDDzW+lBQdFkeHCnXS
yFz0RDQBibmOltGdZsPFvVSVVf3Az5g/6bcwsbTegEiq5tjXBhioScqrWU3tOlD5
iYOonv/5MwhGZ7Wn/pAtOEZmlA2859YWstlUJFGV1h4IDbFV91pk5jLNd3xYftqq
2+nWWbQz4heK34muSV97zPptf+ELk9tAylTZTgSDtdpEeChgO+4W9HvJzGioqPzM
DdH7uPkIv4vHQGW7dsTfGIDZSiJA2BS8AR1NVjcrUCtv16YsfZWYCpPw519/NKO+
fs2BvZGGC3sxsBUqii5W5S9+n/crwbnvhiInSor7vIkOTSDsK7KTMg7SpOOc7+Mp
spkKxQ+knhhmMZh/Emg1EYqUSdzC6ndR84e2yzp5Jcoyt0xZlxCbIfYdCRhDC2Bs
J/hnBeC8aT/L0bzWil3q2ArgSW3EdQJAI58Q7Bx9tElfqvRu77OqUyQtDuWaOZz4
p5dkvIab2RncjeXHZgkTZQsgbF8ZKVq45APF2nJ2Bwf6EcuLCeATb0mOXK2chpei
t4L1CsnlaDCuR4pHXMiPQxs+kinI7bxLqxJg/FpOo9Nhhrd9RIY2UhECQu9+TZlH
dBibuIN5ZOxHwSl/JQYsNLaIVD+gbI0i5TTaxl4aiP8CVECz2Gxxu4ODlUaiMnEx
GCzZDl9q2EYpQbOrZrL5dDBlyMFA6W8qeeYI9X8gDNE+7ffq3EFbFpckHwXHuWbX
7Dv4NSTlyYDgxv1c9CgoKVhgSFsrrM1HR/I9wLIa31Byf1eC90seoVbu5kgiZFIb
TA7TBs3/X1QfNWZ7K5S9OgkQMG9bQIBPDOxC1rIvj+uuSPVN0in/ReKZSgCHH36A
MTOMygYLyMqWMVy1u/MQEUVaOVUUT18K5bfrvQtmJF9h+x32hJl7QMvyzON+B9B3
Fil1Y57cbvENFnjFc0RAR8CSZhYVMUSX7kGK2xCmX1XUVbg5H4i1wf4lw1MgYMf5
LLyLgRqWCD7tYMia9mkeb/1ojcoWizzUtBor3cLNTdNJ9VBKYDvSscRIIoUGP0BD
P98W5ZF2R3sxPBTWJnwdlUHb7hKYtmc3mLThQKMXcbX9eovys8Lky+7LYjTjxcJq
Zy1FbCn3k3YVQCr3BiCxN91ofMtMn8htj2RFLUJicPPMWcLoKzEWylz6Rgkqdy2r
qnn/pmPJQoBBThtnYB8jy57x6BJgJPTmueSv99xpCunvQqave9nIN/NmZ0hPd0nT
WSmpsLP8JfKbdjwiNBg+2iPrbYS5cEaJ17GsONvlG7jPWXkrWuEJdaMCRSdt7Bzt
Hp+CpvIl00VM4UrkRJoYyQXA2g0ICyWHmqudTYFt4fIfTFeDfiqjbTA8jWbK4DrY
BTuniLXpVxx5bm7By9MJiD3j4i8wEEVAUriDRbee66XshA+t05k2qxyq9WJ43hw0
MPpyuvdv1Ee6YTsU4p0aWHR7hpcVTF6sRhsSLgmpfgvwO6Nn97tGu2jmJ0PqnKuR
PppaqXz6y+vHGCt+rL+sdP1JfdQczQjH6urc+oI58Bb/vH0xMWkM4a4vJB2kf9R7
e+x8j9Zgk29eN+pIZJiGeKIE2/5hJR9oYv77XJjV8fvMIOHE57V+UtbRfEzkAzQd
BetXDV13r/FSVDJNKfwwCj7nj00zQe7hdLRAv84Thv/+E4GjspRjW1uNFHwv2Jew
g/uwpNyO+4cf8Y8cjwAxyO13TFp7U0xJNBlMV4KSRJV0XUP3vl5yJcDnYEKJetMU
MxyQfiRLFntV8OKRuGCkk0aFt8wKsUC8S/i9BjNEgMi5g1j89j/meIUNORhmEPqm
90uHh068pySZZ2oJa9vqJS6GoB4PFPmTWuQt3mtGomGiT4LAv8U8x+6MR9T3d32S
uVaP6jA4O3wPmfaTO4cfxXYMBjso/OmKBTY2mulfSoRqP7Wy5EeZbSJvEZV4d57V
DAXRy3Si9UmziIN5TgfXlBrUDF6iruimQmMkNXIAlXn8iTvkYEK2OVdSDsIx2q0U
hXd0F9eW/jYXNYpJFAkC18iYHTGK3Tm1TYsh9lWF1FJA1D3HlaOKwooyorxTRJvb
xPfe0ukAHMF8QbOwen2BWWnYiKe8626HHY8mnsb4oHQzmTtjxnFNaOO5AVR3mM4M
OWOGpUiA9qFg6jUVgpRB4roRNAgr0a0WvZvwa3yruykWBeJG0IqwrWvhVf+7RkQ8
ULWUGJLPOapRfUb3xGDV8hkwuOLOL/ptn9qa4e8WodgZlP+w/pMbC784APHZE20R
h8Y4eFBHk8yDt52kG5QmUcgCPOXfknzgLx0mUILl0ke/COrJevN7iD3yGqZ7YfwL
fafDSNCrNLzZs2szzIrDJz3XdvvrFsrOS71SFDnnrjuTHCNyjkeUbg+8UHZG9dNt
uRFRgQ/KDnlB4tA6bt3eqLBicAAscY97946HLf3e3Ggmv+Nts+OUgrG/I5aFlmDG
7pU4w7HcYot06b7//UaVjSBN7dUR15GxnSicXXEnf5XEH9qmmcrMl7ZGD1OopOkB
p96S2OoqrcKB16lrSFHn0EgIwJTQ9Z7cySpN0n7pO9nqG5sJLOQJPDQ/PlmfkSa+
EJirOj5aNuNpb33hjNAB+PPq/ixTCpnfc9Lwz5R4/zxOuzk1r5lD8gSD9SUUTNTl
H590n8B57pK1yaCGJfmdAUCcN9rVEGgHQbJYg+Xn3X3sdkmwTlnVy5eF3puc6Tun
ygs2zGmTY5VyUKYaIHEnBXNIDajAMkJHSZfD7znqyGfz9ITbVCRlv0RbQwD98tQs
cVx2YM2PhRFAbcSl7kFtckruJmR9dRh/K5UyBiduMVDRSNceIGzic3hMhE5e+gIh
RnWqQvfPMfURidDOloJvyLUy5OWuw5VUMD5oWLA7QelQtUHJ2Qch9AT5olkfEAT/
qtbpyrgBRqKDVZ1LHOjf1sL7fSctm7pzbISynaCQ5UwFDDy4zFgHVIiI4scqpLTv
rVF84H/te4oKKlEHvpiwjcVQq2APkVlftmQuNzGC+AhPImfVYQZSUVxR8QrnPeNh
NwivDmVD2rsRCXjxpgdyH2JlJqopTpK9fRmSg7CujL9ZuNNTgOd8GxyeMZqQOIjx
KAiHCoOsW+z/DAlbWImEJnS3IxkrEOeFDhkkqL6nJo5TD/E6lw31OcuNEAZh2AFx
2HFHSE33xtTZHxKHuc5OhTVhKAR2OnmIZCz/OAyq7sCo8cEa/gKnRaMhmlbf56ZC
h+T6zcD/zOm4CYNHxk509URsykZhBPUHIN979t3rcMVVM94RrsF0srcz5JQJO6D/
Wq/uIDgo2Zus0iT1b84jIOizS3qcIKsZgrNcdVox4FE4XcKbHhXrT6dZm7xu+tF1
CZpRuAL/d9XmsMYRfXduIpUfZ/7sUfT6gQdUgh6ysTSTgI5W+RpfiuNoybAFO69j
lTM8Iov7PVXwM75yPZY8eMz+oO0TsfWJmZ/Us/rV8SxOFrsLcU2avdrbl8BJFTVG
68ptkCW3G3rtODt/dFs5hiey5rTYf7cOwYNftWO6pgmu6qxbgOctSv7VmgKRrqKZ
mOCcubIS73xelG3pEuW8fqaUXKeM60TyzVoO/BU7j8VrXkNKiruj0wpPoLxHUHiz
C7qbecDZShw5CrjRXU/LdWdVJTXTdFClFeqwoxMpxWSOj4XSfEFvOtokxgBNq4yC
wYIQZSWis6jG4Wj0IZgg9Ka+nYZL1RefTVlkpl+NhKDFTjZGl0KSIiqG/B/NWTwq
699/1BpOCw3kfk21jYoEX3S3qNe49R24oufMnqF0gnAYM91g4g2yhVO77Ff1b+BE
zkKMxdm3GUFsTzkn5w+cjJ1Rgx4WcLdkIU1PKMrOaAIyLhEfzQ06Ks25PcrI+hZY
KkHHUujpTuXEVOEHFn3W4oIdicT0Jtce29t3MaPzpbBT09I15caVGAAtYAtCCuCP
+52nrDvWSYEStKLw9GYA01NS/LHaD9IQXOsJGef1PlYVFRWwoAvhDMZD3HLmz6ap
fhqVc2EGQEvsRn1vWV36WUOAKDykAxVKsDLQZUobB7uuvXUs5Yb1zsI4oA8ottXr
zhZodM45bFeMO6ndYOEg4OdW6+Jgxo4PaMp0UddNmjK67Nk7BFU4Mn0Fe/JDXmDx
8w+kKhE+T0lHh/4ZKkI+vMkqM/7K4Xic3R+vEVXTlOYV+ZKRx8mZUSmirYlR2hxM
FKNuGZA1+yKFbCyaisl/dWde0XJ9FX6M5qah7CtrtHj/M7AdoTnpHLTjkwBobbTx
GLyZxV5uugwIYWxP7jWMXDpC9eyDuM5yS2zc3fSCVRc1DYE4xfUdydioL/JQLDGO
Q6G8WXKEf9CsSEuvzHFPjLjcBE6dkeXd+DqNr1Nuv4wJ0i/8eQruq3U+IGyAoA4D
jZwI7s9uu1kVCLzFcFNpwxmp/BcjthX65afdjh9P2ZxHE8cZ4XnwATr24S4+FNSw
VdLHPjA6A//J6YAKEWnxFUvKtn/2TzDmhfuUoUA+qsoae9sH10uE5uj6u6/wT0c5
fNDL8E/ggJ3k7i5ksd16nXzUUMh97NRzYWRg4FFrMwdanlRp7O7n/ODVOu6zMfdZ
hwyGU3wVZ0bTmswBgql0M6qczRt16KHrArUy9FX3ZtpoKensiabV/3lsrHckcAuI
AXB/3/ayUbGMm0tTWuVGgmcA7beeweFywSVxREKfUCaVffNref/Nc6OB6W/NRcPJ
9Cl5IwTIws7T7oZnSx71pNT+XFbK2AJ6Vt5xz3CuRcMnZ9gFFvFtiwvYq40gBW2l
0l6nWZdQrVD2ReD2mS7LqtRo91IyugrAJLYJU0G6NJnu/3vS9V58U7DHaO7zSAzi
rvxy2JPXQJa76Q8U21NQgSiWAnta/vsB0nNemHEmSjHZBri4RFb/L9tXZOjksjvH
+Yv1iXofvIggvF70iYS3GfaBn88juDNB3ZQjcvDp4gB7CNAMxKIA/Uy12ys+2Q2F
jkjynFCa3SXm3D/KeSFDIIcPBVtgieb5FLd79yDn/Wg5PnuBu4kbq5RCqfFpUTz9
Ljl3cmK1Xpxkf0pOt2CBg5ntrPqq0K168qdeDUNlxWabSqyVp85K0ORBNCd8WoxH
t107jVUJ5vZJyWogBxlLYY7lTSxRH2TKUwCR2CrP3LdH08Lto3olXotxxS4MEEOc
9ZOf0hkX4JBzjtPQCvANqjKEXSYykp/3gGJAEgtLyW1kQk3Wq840VABlx6hkBhLC
s/mSl0D295sMjx5WcYR0ApILHGVyI0YHpWbBJh9I9t2W+192B/v3ZgujXYdCxOMI
v129M1kE3Iv00+iVXT6FJ+uJjy8BiwhnGT17GD1PosPswsBOaoi7OjdpXCgt/fYe
MYssX0ByZ3ZYBGBbvpMwUH3p7GShVs1oRhnRCBeZNmhPSYqBnpOtKFwmbCZ88C60
+YMdXTWCMhvRAevYFSqAvGTDfCutpyQZmPwHiaE2ddiXLUx7AIZwwmqFTrttuMN6
fPIy40Zg9zvVDUlsUG3QEEIL4i1emkZKeV3gjZWlNZtk9p7lRQgy87t8uhCryp8h
d5NFeIB5nK56jodLywuSq6/60MFzCXvhRu7Px3Wx2+jrQa77sfNi5pWYg4u0Ktk6
LhT+bIflJLOKOI3X3z7UgOD4+Apeqt3Axs/aC3wCIfWj+SPyGOZoYPRg3JMJ52Bw
XKcsRMvoty9EOz43QQAqpxsuHInnngxKmxaBgtvox2BMiGr0al3IaWeUmKDsMkqZ
psOrgegJGzH3lekfIPmHjwuKT31zFpiaHE+Mi3RPi5jht+8sN86ZhjrMTuUw8E2a
KaHHqKkL04PK8p10cM4IZw4qmftuM6o00axjCnH5o8rF44T1LK+ylQYrvNqPm0In
kHImN5jEnvlS38/BB8CnQ1ae27cYqsUNcYR9WR6XAkoZzYXXMWFDU2R8DVbN2lG0
6lfbUIpahZOcf3bRleQYM+U/D3tFWvZ8NCuFcZSDBWsBBhDjL0O4LbBGwtuqGfpM
+w2+BXsCIjIjpF9cU7rQmpRRtkawCbqtUP/HtzLuwAClXYNymjLM8ZlkDP6jYQdY
Ga8W5VGuEru+0frIoHt0LFQox6r2eTXP/XKt4R5BeBQt1Jz5f9j6ceQZlHHyyNUg
5cENYw3D7Kkj5a3W7VTAF1Lzvmw/6mIltOBgIxm1yfSo2joUFUZ1kLjZFNSzgAol
MMqaDgBzJ5mFbmxYQAMQhnkSez6fms2/Z8vah0zQuMXIY8i5conJMuLJV5OxqNQc
yCkFD3WPKc9KUjeCzYtMs3oOz0ZwlhZxA7pBl2pvTodKHlvtuSlOer3TWRRbQOFF
qxik+VJv/G7FWdQZ6XsMhQIbeAPE0DVHgNhdshz6T79ZS6JQBf3TLq/dQ4VgqXW3
1pTi9j+06YXdMOCxqDbSdzc1ZBj3/ay6CvoIHGj/hBwh5RTAHINwyzCwzRwkmigA
JjGWC1CH17zwTwHXf9HVJeJLr5l1/XW9CYx4bmQTeNukULatahYRYA/ZvpN/11jy
9kJQ6dKfA/CCkcwL4CIdh9+VnpS/ASYMDf9m7TIDcpPb+eYAEw7O9bhY1u+kc9WP
AoaQ6qMaITGOjagUKrlxQSbQAJ/cW0NSMBqmqLbVRV7nHtnyLUAxZ4UvoaTS/ayJ
EDtaq/ihpx2v6aKj8yiaaqOVHSfi44cu7Cv5c26V4A+9uR4rXg0vp/d+uJvA7g2V
n+KE8rNyXhNBoZrG+h9GPdGS4AgkLs45f7T9VIVAFFS6hCVhZUpv8klthVKDRjxW
TlZftjAMfXC86L2qsMAWtUPMEfoXKherBhKvDumISKcfy5DeDVNnQh7WRia8/YFD
iLS8Y0mDxahEjqK4/E3LKvXuqaQGC+NKGmYazNgl6+AC7fzlyTX7jl9TlYdDbtZD
YCnHLsdaqeyb36Wchwkatrzbq09V2oNEos68t50B9CepAfXOWr+mbrFf0tg0CYel
I8JXPIBFHpceSOpoYia9NURlvNOP2HogEftWDpwjDcLz+25G4z7d5Gopb7E7hkXD
IR2O71MOHZRxttNEAZ46j0N/geB76CQNT18U+KuH0u1BkqV7LbhhATjndeFQt03W
1EBubcgVUnAGI2d4M9OxJPrDabEpK8GnN3VLZ3cJcCyBNL1ulcBt0j/KvS+0yapk
bSvkW1KslbCAzc6EyGmPX0+d09+RhWtp14EfhoClhimerMywtHDxgCJjVAuUrNlE
dN5XBXXNTkwwh8Y7ApI6bcjpOAX+9aC2bxo5hyvXNFWuSY2oLxcY3IYr/ReXsdd7
bZ6f4vYebgLIJEwddqXWcuXa3rMg1oJEeTtEBVESGII51sDCV1Rn85gfT4U0MsSY
XWNRefW8mN9IqIjPY8DC5N3PwHIBf6xwAUIwEsDJjYO7ygx9V5oOG+tnEyluG56G
OMEruk9ihbfWpFiDclnFTdICi6pGRhv+5lMcwk9rFvCWHTYU3uetOZD4Pr3UG+ks
yfNz/z1CUI2vucNQNxrTwCbNb2FJ3lwbkfYoFmw9ae6UiLIEs1nGxaC3Pj8LFWY1
3uYWso8gwGuNEw9IMgQvAuf6XfZFBhL8dLCbGU2xd7BF/My0aLx1bCZg3RhmvReq
Bbyf1hde4yj03fNN79TIN4/tz6gVfBGNldTlJKf9qmpJ1EtzfyBaV2pNenCF7q71
icpw3nptxF/1y+vs4SLJQUB4smhdrzuQ0fcFzFU7GWsgDe7WL6SG6dfHHFRhaLT5
3h6MKf6CG+dpXSabGv1r7WFoyZb26CV8pCBNzxWg4u3zoBf2I97VOYdtsmZObNF9
xy3TF10uYpptHCc080WefR/3ozMNJDUT/axsmh04P6RQ6hh2PLBh6rZOY1OhQb91
4w8CMJlHgb4v8yGLaR/c+h8G2Gj8XbaWWM6/RxFb+KKUoUxfGNtta0NJqMyu7Odn
waNKeiTAuNGmBhoSoJCzcMA+jtr1ApI/DAMH4Kc6a19J0cAEthQxrhU85HSy2mQK
COT6lohzhR0KbLuGBjrHmGnRtjDbdZDTAaKXMR9XKoDYiKr8c92KrffovCB26nGp
XeMKXJ0W4oMiqSSKi4zVXd4ZPv4ZfBcIu978Z6a+nOYJ5fQwRTQB61GBpYBuoe8d
Oa1w8/fOsQ5yr9IrGxqxF2hbYDM3lzLfcp5GkUtKV29b6b10GBGGtEA+3dkWYLIb
3em3rz0cQprhjhyZ7xQHN+30CKl57eA2iPAwBOdj25h9rww09YMrvvtAYfXEAaox
XTwiSf8xHwjMrkAjFXKZNhSRK7B/seBOHRRyDmXgHOb2F70YfG+waH3UYGSNLicj
0yYBRlEPmggW1BoQC0itvzPbM+9lGMCsPfKkLlSFBpkm8i3sXuPVQlbDI1m4o5ye
+VDHW1033DyafIHAtP70Jz1DJuMF3Wp3XFzAQtN7JpvZQBbs7i9xIicmZfGjqFxJ
4uP5BCMXNK58iWRkGDac31wm6ptLSfxxkrAA/vLr473csPvoAZsVkg1CkTG9gaUF
2ALuIz3JIHpNnjsH3W64wrsU7LCTDd3HG6gA4P5wNiGRxBKDfPd7MGdB/lyLq7JF
0kgQtnYf+IpnmRQk4//6kJVUMSVuxpmr9N/dCAP+/p/hepD4jF8uPpipVmIAjcOZ
9kddHKO9Wh7qz1BynUovQFksWAg++63OdtByxR5/co+KJIB31x+Si1xQHAp9pjhH
S3/cf676jsyGQIOnq5chR3hqqPjzYVI+dJ5kzjcI4ZslaHiem9wF3k57uCAkQo6L
9ghQ0W79ZnGuWb6oWM6ycx+1pS/um3yT7Mne2z2RZPIpstb85M+N27BqHPpeqPdQ
/aclTXqYbOb6ReWDvN+4q8UfQIWbCmVqOya6zOKyUr3laM9UZFYmdWkis69wX7b9
uCaA5IqYw3eb+EEwZUJWQoaaol2W7bBVUF8mAne91CfFcTF9lqEJjDflwEK8chAC
q5Phlvd7/m4+j86e4qSv3THAWQwhiTUtvdo41cF4Mep5Gy085FA8JT1oKOBR2EkS
1bDTF1R3aMuUkxPxQNonOLYbUcuuwCGRMXJ7WPaNR6e60tsKzeXq8c/kBfA7OUe7
/cN5tjM7W9q9sDLGwELmZdePV9+RcDC3GUjrgol8mAjHpiqQwrYaKTRW6PaCpuJx
TT6+qKcMT6tvjtT40cyUg2nahTKeZMj1Wuai/3nwjf/vf0wTVdGgeJhEpxxiICay
DzTiP22GlciE9U4mxCsLvyy/EB4BrZ+ji5de20cy0r63U92rgf/No1FSbvtU5R5O
p+2Cdz9sp1TTd3GByl+HRfZmzM6Gr/ZRUgBMaOddCoXqNB4rva3eh3UgssFPtY1N
dmF3chxU6blDLnyPy8bFFNwCyvK4XU0hamPgWDBHEtHMF6NBY62c+CoGBSci6pU5
ohpyvXCwVaV2kcYhlban0M1Rk2GJezex6+zx6ji5ncYXq2rdbW67fb3DbOhIzUDv
06DWdq6lBcYx9FcKpN25lr8VVQbePBd5W16arCvYPEqGZaNyveHvmf12zqxWm1G7
aZnwKz8nmvNY4r32f1wM2aoDfDaC0r/scbpD4DPkaTHFgVROc92W7wNgaJd53a+e
D6RTu4DVwo6FS+3MnKuZ2Fy39GUGaTZ+zpqnjuLMmi58x+Y7zAzuMNOr3GvVzjue
87AZ/8BEFB+sPPsZV2zvv7/Pw/VkCIgkNmEbWSCxlCgereVHI2pi3l0q6NdsR3cA
afLNAAW6Iofrbli4x6cXHueE4ALz+JxC2rnwO9/nTHXYOQlFUmq6SBhuROOir/6L
tpwNgkN+cRxXPj/n4wi5/BsYbAb9iyXRflEzApCFv2SXWRKBbAdc6rNYCqU3r1z6
rsyNAlV+Ma96DyoRfPHrTW7G6FLfeXWOlU+8XleuDhSRf39oi7ybC4DrNk/US8Pe
uaz/Hs4c9anWZV8g7Upmh5Cc5ZsuNLqkMiBdNZ3g1Hl09xAp2Ta270Gs1iGWL08Y
lqcXIKB7Phk/F0jVjJWu3ZdQf0HXqop7kcQu4YZabb1hoN7xa2KyDw92zhKn/Erg
9mKw9ashshU0kK7kyaK1O+RFhzH0E80XQYIFNk5ENeC2Ap94qnOXJcLP7UHWvfrd
xS8B01GcvhhSgtcVyKsTojRSvvhekgamT2a1eAxSP3dHSeyz7Pf+lvrFu4LJ2sFL
HpClXPTf2bCt3b7RVDLQxsryDPA98lfQNDPFSZtd67c5SuNMNGT4Y5vNCFXrqtBG
XqVMxVwiiVWtC2b/IInLik9LMUyoHRJcmzDUkG3jIfgIW5PtHnCBPwFeMK/Bp8Xh
sEMMHf3vdySlp9HufhSJifH0r6dbO4bLhZG/Cegni7VNlQYiQE1VlR6/hmUoXo5d
mPjtmJuXwRj8AokSGaDt3kvBtP0zN3ABuSdEWm8fnOdv3vBsU+KgCrL5TVq7G7SQ
Upf0gNosLgEuJlXFt26szPo3Q6bcUCZEKIIyNDDntB+B9A174NlWy8a8OL2Iqc8y
2WkiGCK1g+eFgLVck58oGdoDLOM2JtzFlL504DYsCUYI2ITJn2ReqoZ5ZMErPUVQ
G8hFanlrlU0BzOcKRr7M/BKS8XT459hFyutoUhfDNQjvhtKOdlUhiXx5lAllKkNo
iHLUdHjBVwX+REubJG6NOHdVlhFgCnL84pQxjXdkpAbMalN5AWCO/LbK8AJt3nKN
Fi/yBQnridj4EGOS5tsvHpYwQwdmse/Q74BrUSaY5IIOCg9pHEj4PVok4dmrqM3V
fCehHs943llhjScRt7RRByYvZcUL0rsMpzbf7PDCG/NVc3UNcmivK0JasmfANC6u
aj3Q28/LfQ3AVm8v5xk3MrR46URPTSsLTV+jmIqaR9EH8VsxGCfv7waHL3eDAqMi
u0yZSuMZxIrswkObVjcMI5rY/uRJcqxMpEOGa7Z8OoShD1+ICzJi9f0xR/hseQxG
l1oylVSqV7cAjGx5ooHRFxFxKFR5goDYy7LV/CjnFflBMGtZmRMPMw1CBJlHHsMP
tG6g/vD5GVrWNJ/Ve5ZLvRv8k1xPrTj0L1WF3mqpksNjJaBap9nFiI0HcOJpuBFv
WQSgyVgUJwAf97I+LZ0RGi0qOGapWTn+mbAyFYCeCfL0HsGPCMKQdlUF3E96OUL/
z7PkL41+NI7wFrlOMUL52LGKW7zIWuuTikNTxmSicmXmO8z9MABI6P0cyWcAawVY
N8zVo0qQ2zkiQFebuJXcfHThtHMckjPErm3+AHqxkBqWBxE72I3Y+iJg7f0zL3Wa
s63p2OLp4a2sWTX+8X1eSu4yc1qA36aacRSSDnf15WkeUMvsdzAdh8q0v5lcAFU6
ri1ORjK+Taekyf8KSrS8FfDzuBtNAZdyNSQhE8lLoFBIvldhe+kNdLa7rhGCeVts
nFnxAVZrMfnMDGgfHjXLBhRFjI5/0f6Vymq96DnAT/my5xPTtt0diiI4qna4Ap8I
9JP7JN7mtDVqXQYjN5mlGVuDoUecBuOr/afim1qfN6piOl3C56ZQmQxKUHd6+CXd
Gthy4GmE4qWAOqY88+Q9iHe7hf9wgu9MGL4ufcuZLbu8IC6NOqix9H577dVTVZIi
ja32JJSHQ0gOhneZgEoegJY7//cBYZycLzCHvzQUQy7qYQ3i6WIC/iLZf0/pvxCN
Z7KUJbAijmfcJG166MUrjcpa4BZbfmQBOgKN5GJHSIftxEYIKnI/5NDizdG3ZI8U
L/eRcfWd5cymGpVo+lcMeHzdhE/lLtL0GS0UMuvzCy4gvWZ6sMu6P3bq4Z95ThWI
NmG92PXm44JykhdheM+lENR5k5qEvkIj6XNrMEiIkCadIQWvtDdiPQTqeJY4yq0J
KWcICeI+agiJ2za3ggwagaYa13dNNt8MkFG9pbeT9phZvy4OabXibENVbhLD6lRr
a6rDDqmNreLWsi+FEC7lixMZyfl0kYyMr/X2f+JWlPHTCyk+swloc0UJ0x9N7kpy
291Wd0wCMRXyZTXFX5wVK4vFb0760iSBGlGOYL6JUs98jUUn3h2m0xPrvqjKz79Z
12FW/sexfOnDd0LUILZSMgUatWujedwF86ykOaapbroQjnd46fPPxn1Iv5FhEqva
w7FopZgr4PqlffW7LVQDLgnnYPpvqvpFXu7cI/g7RqfD2J/f/kLlmIZQ58ufpVOO
Z2uth9gMBDsJ+v5WFa7MipdU8luTu4sXFr08dmc+BTrigdfvOD4LBsHneMZQNHzf
FFfvceeUu45y1EQ8Sefpbc2rp2eJkYc+Ftk4lUqT/WG6i9Ku4mkRXZfq+Q7AMzL0
NE+9ePtlUJSI1unaUnjLuCaaBpqk5toaCMkd9xEQSnzwyJ5HW/8uVPgkwOtp94Ym
m3SSc8NcevQJHve8Xf2IsIwMxx3QxrrG2GqPE6ZIaIipnAk5c7TxhEWgC+U807Fw
sPSsi3xK683kZbxJsM4AIzZvuMyMiqRCEm0PPaIKS4Bzutyim4BxKpiuTSPGUksH
LVEhwd1gGCCmVMDpHDSx5cYFtMcnT7wzbdrKghluAohodYoNBQEPoFRQ4/LeXDkE
Oa4IVqSnsqhMQyumAm/rOl7/nZ2cu4kNiAsA+3cNxMlKxJ55IeMTdP27yu19HKlv
kyPQL/Qzlhd9VJCUoaIO/EJtRN+VRUpZ7XvcHkADrqCOdDYgPko08etv0p+NCuBI
5FEirtm13IuDhmOhjvOwVzzg0eNZOCAVz2dktxKkuXT8OD+A6th6RWlzk7im952+
W4cp8EY+/tLY8SDhlT9XRLY59ou4+gjXlrGqtwRW9gdgyyzuJH7+V4AeGdQMwrQe
C7GMFIaphZv4ozcKuZM7FP7QJ4sP/LLUbDXpjuvnNyggSxduHsB8EDJgmtd7jSRV
grr8KrymNAIeyJqtMjt8DOpRPrdovPHchfQWkKFQnHylhqZwP9UaC9xCtcEAlNMv
WaIxrJLdOmuuWXpNO//1mbwLQyIxnhy7QxnvE2DnWX3upsBTfoo30TQCaD8loVB3
BfOMuESvb4UwiScu3053BN4Z9Jq7KzJK+dU2HOiyYYPJbg+Cvby7FtZo3i/HgmCT
CZlBx4+D2P5XoNu5+TIjcdIDKuxENmNEDzNyaLQNfyKhk5YTG0g9vo/c/ZrkvORi
NScVjfSbmRWmRGLOhzraq7e0SalTMoLl8/ieYhGGs1AKERUuXCrBOH02NZ9gwBM3
vHQT3DcoQ2GWVE4Nc3a7fOmGlMlXKDCxIU8Ok3jTYGM7jYPje+ralJHowir39hJP
k2N+UNmOjMFH+QxIvcxysRTtd45s+sPbPpBwWLp19pmisi04PJzWDF/CGnALF/Pn
mtJteFwzKfJqouz7m3zvZUj4iWFizDrWQ/zoxkQf4dPI+ec8fqh0Ti8CiIaP15EZ
xfbNlTtZVi+ls29KeBUWa2NQCRJ1NnlqtYLQisvlar3VMcJnal39MYlpJH1qdapj
dn4vt8gLpKRdqu1eEdHed0pEC3JZNzts7C9ggCRaUM2UYOu0zZRTq+5iBj7/pb1w
BIJvlZfZHWZ5JaFi9GOKa08JwkExpRbKB699EODloltg/PpmoVtsblqo124oRoCf
kv5kunKFoAw3nkwKBF5tVDuQo26fKzAegCcuuslVUDUfLvnFDJnGxFGqpBesfof0
oNIHhswGbnMBVEz5bz2XiGarCDFf1jmrXnqz7srNqhOU8o73xM39rqeEwiZsFgBa
+1L5g3MEh1xfGDQcM1K6lvWf0BjGzjNmGaSirWzP2G5GErfrJyrhymodj2JlQ+fU
MxAwE+V4gJ55+XZZ7dsdyyNo4wF8X3hFmMUJ7Y7v7wmd/oDGjax3281SVyc8orqm
5Yvej6poM9nFT8JWBjC5fE2cCbH4vmoFhXVJLlAOklUpXUIVRgvzry3w23jaAEyj
vO25Y5eIYl4fBYBwYmBHN/6y2HJHxBh6uVehqthys3Fxrag7a9bhgRxcyDBPdEJb
oC1KG9lzlBRaAVdjuXQyFZcxy6LvcvPN2ZcUDa2da5auNz2RuavyZgITzE8yg/qW
x4vO31YZJ+vmPfJIToPZxm2NTD9WM2O2bfBqrljMEqJ5q80QvkmVepwvMWmYSyGS
D+/RScGh0gid7W/7uv3DRHMw/KkeVd4s31dxLm8hpBxG5CHyEtOD86Z8B5WIkchy
eDtUjrUTA/16l3FUJlPV/KPaCbk9YiwGbMcDyYs/Hxcd7D8AQa9c8LxD/TLEQy9N
m/BNsp/wSPY7Ka38ANgHN1+VhCS73Ikyc/3N+fyHHtWCKG/jHLWUOrxfPIKlb3Gg
Kxck1XzMB1ZBL2GED7yjt/Nj6SWnH+Qg7GbdQ5NcxXNvRDO9OELX+H2C+0UO3yBw
DsiUr89CAo90pkz3rgLwUvewoA+zxPXi0rLO9mr1w6p8s7ew411EKKIaTkRa+rEm
55B9VNZ20mI2/Ubg15eI9lk8NxTjGPxW55iReIWHkFTh5g1grkrNwCe29D/cXHL5
lZKrgFtcHM9efXbu7CsMbs1OTBKPwqZWTp61uL0CsBmdeyv+WBjsgp2igjje1XEQ
l/qUQ86jwOpDBmfOFc0DlxbPFcwuCuAyEjW0ta0+K3J8XsEgq8rZsPIafdtOlfHs
dOrk4KjH/5iEQOYSZ0WBX9V54oG5aJcHGh5mIAeLxsW9FiZiBsPH3v4gc+n2ZNA1
hk2LF3v72WdFSRbpEM0ZcIPtAk59O6ySrMbZWtZqJXQGhhHpO/4OyvLD+aqZOO/2
aeOqcBfG5czD8YDGFOhPTvzS1Dfu0482utVqhjQJEd/4z4UdjEhY5X6CBzzCTxX5
VG14YSldQn+Ch3fsLTT9GtgYV/gXlrrIFo07Ypj1ylzRW9k8eVfurbnox9crVmPa
pXIHrlhHLPzkxB3Q3+pqXpgFQ3MYKutaurncCu/FibUAzpKEa/mBdf0owSmAHbdH
tImHIrnPEmYJpL87sl+Z1TlLhaS78Gw/AAv337aUo13VagY6NIjhNfZJhVFK88rr
JtZEk9LGhx6VnFz8qCfviVNBoEXBulve4eHjZwIi+6mclHZH3UNp22Y0Un+Dh0UU
bwA5P+JbxgktCYIhl5Sffzi6FO3oIhrty6NRvJjs2UP7ifPq0znaMf26ddnKXego
KhbFuvVIhcuaTr3kNoWpLbNoyag+NG6rsMWMkEkDK+73WyB0BoA4tgOo97Ze53A+
vDS21AlX7OHbaaGBFrnFzbYLzmiUxN/Ij2+anck4uOFiW2yNej4p2u47s2dWCvsi
2zhKyQ1R1iYdg5QAO3F5kCesUJC2YGT7ZAY8MYNp4xILrirroMAfw4s6VTMAIHzS
SprI3Fb02C019ZNldcSzz/2gC9tRWw54WF2MDQdiE1FeWDc/UAfEMVj/ROvhXGxw
29dKWYY8cLppOs635sy2YYGBv7oESVYVq98/csdUXOjscUzEoRr1VRmlSyjx7i8E
Ek00jOVoTBWxHZIN3qxk0m9oW+1qvOnu1E02IHFFsU/4b8ZG76KG6i6EpDQFf5E2
5j52v8infFHlcv8nvZPwNceCOsXF6doZTcEJ9v+LEaqW+YfXF9fAZPscb7gqUWoB
LD72eUaUIpvhBW/HY8cUo7T7C+6sYSzHSYcgbxLaboe6StBKAE7va8x1BQ9yF1tU
Fcibc9kLFj2ptp1yaun4V/m26rCSMFlmlUVQii5zZJA6UMqMpy5ye3pCudhv8KWz
v9N55ldZir73V4KP4tnnyMqtHzlDhcnC0viUoBw/BfW4Z0++m8Wv/pWRvm0pybDh
uOaO+BPMxZEwIvf7LjdPoi8Kn8Ns1JkJgrHNV7zvgdYabGXPKSyBE2PG1wbBacBi
5lxN97kKdyLc3e7jn9cgKkwG2zTI3kCWXi7HoR64op3SLnlGoQAXJoUYgopi/ZPv
CMtcakSZ1/ilWuJ81SxZ6iT7TpFdpPCF1zO8f8lb98QFF9Utw16ojaZJ3eU5zXuO
xt1rGdL7VFmGzPsEoRSz2/6Gra0t6Ijx+5n6q05mu2Eu5+AMDDmEJ0RPRqDiK14F
zgCV3x7znoQJ17auwHJPMBZgODuXho1vkmbyHYCX1yWAZ4LDXZhYg3YDiqYBOLaM
t7WI5+J/DlGygfGOuyee00d69OFCA6W+ZmldXlnQiEA5cCwsHUPHDL+N0hwsoc9I
44O0vwi5UXWJTSoJWm0sYnk+85XKQEypW0UbkPjsHIBjLKRVDKMr8aWRIryA0PBe
v+HCWXoc02GNMt5CtYiGpbuO7ZXrwPWukdLuaPYAElciByiBJEOlmbdDJlC5/K/D
eO3VhQw3yKQh8RVEmnFhl+nsKFi6i08HB8rsq6ty2zQZrA6INsTzm/qHWf2oJnRI
Ez6qOEfgqTUqEUV18JjimZrNXfh4l54t+qoCbIDNuFYy4ZJ/t7xisL6ldWyOsIhz
jQ4NUU7tMFxrFgbt9V5xj6Kk/VTOs8yCwjiVdmXHDt4yg2VkNGMWjSNWhnyWKC3Z
DiJSlrR/D7eeBEfonrRvHRLvFrQBuPGvbNfiBukeTBYtyEufzAh8gVFEY4cq2kta
it7V3iccPpC7J0LUZOx/Vg+Njp5gZ0yuex/Ei0BKSdD0nb8GkmRfGdYHNStuuoAp
yVqZU7Zv8rQb0VO6f5k+/fZ9G0aTNFauNpepxziRt738J8WMlEsVj4EHax+aOJXs
KjmcIebQPHXYidbs+j1fgq2mxqW14u98oiLNSlT4M3dpg40oaC51L009iYDTHum+
7UCRDRQEX4v19Jxd+LV1nr+KYHPe6HN5O2hgkoC6vva6rYUs4La5J0LSsgbB0cE5
rG/nhO2tL04Hr48fQRLXiPBdZ8Og/wL9+RVTztW2xkY2cRA+skpxATUmkV7zJMu3
I8HdzkjLQqLgJKCV1yDJyNHxFuSx8wTqviYKcrdh6iiikn9mu0N/Gumj25P9wN6i
WMlBbkZ+y9/Fm27sWfGsETDrDP90v/Lskw/SH6CwLvnQp+pidrc3H1sCit+YYgSR
GwagwOtf8BYf+0KSwQAg88sVUHyhus0sJ6/ZwvnV42c9XtcSz0hzgXdkRWxah6MF
V9Bn4Z7dAIn8XLXWw1bEIm/BzNYQDzP/KYOIKDC1OUtKy7M8qevJEtQcTAoxJ+qy
5gicNeVaEUqM2ddhaw3tH4H7t0m6zxfNt+2LoUgAoTscUenQKXRdEki4ux0xcHjA
0bZl3iWYjSwzetzFSbP54AQTGosJinKkzN0uNRaeFgv3uzd8pLxAizQyG/JFrDMg
pQN9YwXqF+FhL9iAhdGf/afFDyOYvfa1RnKc4/z8fO8BNd9eAYoc7kj0ZquggXQb
3k4yclG1axJP7ryDRqKS/fDB+v0sFkpwT5y5DcTrbMo2tgdyNLfUQHsKSsIwbvwe
u4GsnPJ+WaJOsjOho6LJIAwwBVL+AkkC/HrdQtmubVLcpZg6MRzMNLL6+VGrzmUz
2yoDp43IoZyr+Nqh5efdVA5aqAhgTj77l0idQ4ERg27/uBY0XpVfMmZbcP9Eaxr/
BuUxSJVPEK5yGn7YmL/Kag+ymOwMajWo0IQuO3eOrGw9IPF5sqaNGBRORBH1+AAy
6ekcZh714Arox4+nRKB554cAc1dfmwJVkNS81H+8dUdbAlcfSac7D5KiABpR2S3k
b5/YFhhxbUsimyaHPhfHGM9Da1sCo+QG/Bp6jWhY72wSm5kuWWY3FD2krAkYCNby
e9jPGXEY9tukuKqc+6DYdE3cE8h7yArhDP+r62mp13b2UkadbRQgQW4EwkhoIUoM
j0fs3IxQYwrI8V9nIPp3LUCPcXaeVFoDpgU4JZxdlxlyJTyZYhh3dTegU5SpTPif
w5lL2gjhs+aGUkqRWdcHARl0KZ1cBAoArJ9f/RkL/+J+ZE1Vno2prtD2kWZYRNDa
IXGeIqYWKXhm8ZVM3nE/XM8wXH5cxQ5zQj6Q2mWgIh2doqRP9ezxmKppVgYvZ4AG
hqRzths/bi0u5fkAqiuAwZs65oJDnycGf3Zzdh/fojJ4Y7uc2HgkWFR8efhgq28n
sNYH+LreAEnKx04CCns5kn/SmO+3X8Z3h61lZy0XGTnihrL+Dl/DPiIvlp0yTsA1
P9VJMnrAn04lliKfDAtu7teqhdZZOld2BlGgGhYDabrF4sVT3VgOK4bTi4LO2LEq
mOU5xrXVlNruxDAyoiC5phDs1OwKghQIV3wETLQ7ouGymDxIEFTabNF5mM17KfUa
b1oJdqFe6P8hBVCcwFuFYjqD7Yw25DHfe4qncaj5n5bzep+pHkNt+3JGOlilWU0p
aFH0n28r7EUvnYiBZe6DPBhezZzKnMYdUF5yYymR+5nAH5EbyAYnOLanAtLSECRK
qk1lG/qBpUWYiHFS/lXQnM+tPOHS6kNwKLLCP8tkOq98w6NETntdal9zA1q7mafw
axpR3E3T9BCPP/D8UJBAgVcKwGiS/ohrtR0JeNzPYhOuBAAM8aOGGxPLtFvw0GPO
dly/C/qFKxYhEgopldAt3IA2gEWmZypT4OOGdj4QNFHWxJoP5gSSW7Ja3DbBlBnL
T1bNsbf6ga9kWZWocu1ZwBJf2Ge3lyvOgypWHuVK5LvPYJIlxz3nmuyX5AR04/uO
g+s4Er3+xlnaI7yWft3W8dhPHlLXQpIg5Z/C+Vv1Z5zAtFfT9lMSVGS/rtqqqykU
mVkw0FkqLSVCPLRPMzmqXgRJqsz9WEyrHS1yxwwxuIAM+YxzIk/yX8Ry4yU0Gt/5
By/ui1Pi38q4eKiDXSIe6ggw39eMNGHtzSyo2hE4lZGKlhwTLE//J8i17UNyowIh
FHHuVWpCIZB/SRNMl3SWv0f30ubJqJdV+T1IHvt9Z5kgifWwDpaR/ap5WzKc92R3
vMgslX7HCLFtZsw1AEyrqGjxdnALdhxM+yw4xzZNP7LKOvjIvojCbMbjC4iR6Cly
Zq0WubahasIsznpt/GXcgFOdflJ9t62rKe+3ednrWEljXvAMRoS5nmJqbuX8omXp
WP9Qd43XU6Byy39enEVsB3QeVpQIEQ5mcWZTr4nlxTTSJRmio8aAt8LsqAZOtI+E
b5JRXUBoXMRUd41lfOd9UYh9bMmaDBQylPbsa0jTRvSc/EE1tEy5eepa8aCwyiSE
nUliUPRcJy9Pys3sM/6xlAcy7iZUapq/udJyv6+0xrj3OEoa37eH/Zyu0SjJ6Vu7
Cu/YN8fulUjpym793d02D25Z8hJFZJqfbgtGEOIEPX5nLFXYT/tNi7W6AUcRvsBG
KdBCmGordMBch+yoe24fDmFmG32yW/LOhF1+Wk3EJYfcC0v+r0f/KeJfGy0nkYfR
to1r/I7Ipw2Qinut5avfv74eXtFSzI4BG2424bko+kkw2w+q6jLMNsxaBUiKIg8G
60xZVUhR/OD7oo4K1ryyqX2DhnE50ySWko95LUe3BZ4zgq+MwiKyA1VhzawKLRT3
g3E8lUG504u1YDWn3geahYMnW7cxkTbpLLoFMDVRVV19O6mIx139Yzz/mIA3rTqF
Qv7xxVCzQyJmMDx/W1Zb553R9+PgOPH6r0tMGbydYZKuFWXqBH4CiXLwbc5B9yIS
x4d9zL8rOxdVYlVUOqJoDlEiYDf+anQWN3habT0BlNUlry2CBcneLlnxkcmYJbaC
sGv7zeeVdbSLSJ4GYwsV7idzBC1ruOpAOOxJHFUiU5ypi/lktGyFuhRMI5zWb8od
kdIW0kYcnJrNQo5N4SE+/2GiwTemWWoaz42TZsVH7GxVs9mXDAgZEEUHKesOPG/7
a+1Y8AEcFiILEea6CBFKY15lUSUeSf2oGxb1WVl37wUEfzoQXPBLUjX4Bfc1A96u
ODH0h/cpamSXxh3Q3TWFqwG9fqOBqsiCTeT1wMhnpVQ81SvcxHNcKJ1deC1ZtVhX
MWhg39zNgreLV4gISWwRCv+l8vyB4NIJQoo7zcgnTo8RNu8euxuNAiFjFIy0CSxy
h+bVdQ6Cjjsc0+TLMcXi68pFbN8PNXhgl4Yk9RvKcIZ2Q9G1Mj+Z01b4f2EZ+5Yu
XaH6Iccj9s1SqjxOmsrC+3H/lQmgygP+wcpYHSpF5i02mUJY4OYskFhGZ+53ryH/
Vm1SCoUAjvr6Fwfo3f4naP5K6EdgVp56A5eOT4iJvyFjuPKsTe/Gazddf4cY2erZ
Ppz2kffF3Tv6xPDU/g+Ds6nedw3RniVMUFV+fb3rxkmO/3wrgj6o/1q0lFFHgjlx
u6Cil4fvW5+aaHCZufn1hleQfD1uWrNoPGwiofrFTTX+5L/Ii2AXUGfi2v4f/KVT
aY3qHg9gPzSmEXx9uVTlS4AVLd7TXo8KZ980p/lSfxSiNiRbnN5jugqwRNht5TR6
+lLjQe1DHi02WBPmIAZmdyvq6f5GlLmaZk+P2V+0s+uKnsLebBaHBDKWqEFhW1O9
nmEckPjHHvOu/cVtVjDkDkDKmf5KlHdNDe2hO+Op7fFKDrgCwJ+iisO9jeHNyRO/
Xc8AR/aUZMYZAIe5GteZGC067pGLoayStYQQ3sWyJ4FGQZ6UETvzxIdiJUGS2LTn
Sd2zn0EFoBuR9vB90VPpr1Q0AqiT0O5CA3+/iZGk2Wxc+BhHBuNAih1H4ZsYo9t8
h2agoWcfyUafoh+t2yQ19sD+jTNEOEtHkIJ/wOUr8FuGVhfNgUItICXQmVehPfER
jZemWmYWya3WyyJcIfi8blLi3z6V+w2lSlMT38Z6eRKXHYtni83Hb5QV5LpPK1pY
UTRyRQLxWh2Hbvb9Bz1KAlo5GRzjh5HGF9pM2RNJjH5ugDzjhPTlwqjaTrB80kQS
yYSLDdBaIRWdnB8s/bki3Wd0zyS3A2gVsKLK7oC3ZryoxIAtblz4c1Sa7XYgV2tB
b5GOamFMk9voIfTkhB4MXv45ZMr/f6mKS+dsGVkVeL9COpX6uDEvPha6V0R1pews
tRk4B7x1kfxaew50QyfqHe/6wQgWJsRC239LnoefPdVs0jJW+wLa+Qx6KVIFkW0E
fEMy3Gxq0ftTEkR9tXE17PgeChNGY1zuXLF0qH4iF2PdZPU8QdP8ln0+mbyRDznc
EDOxOu+4nwf1Hv8iJRu1RNEwaWPYQF5dRzqi8L3oWbkpwgkuchre3EBViPIh/2MQ
aOgFnV7xY1E9qM4egP/F5x5vfvAA1MDJRw+fesSdt0yqkT7wukAza8fFs42YsVQy
UmOusEtSL7e2mTYFmAacX+FAO2j6bv8WTNTBw7obgUtejJ8CuOe9FNygZj7549aj
ODU0RTBQ7ooy300zOAYs5hrDrkfv94DmlFO6irq+t1/OA2FOSyhlB94OM7wfU9eR
zw7f9Y7+AeyD2rBCYHd1K0FZOOpbKDy9PiHxlLDqq+hzXqtjCtFH8HYfv4HD9JLh
eG1rUo6YzQf6jB3AcRLTDSeW1jucl6FU8FaD9k43avWC0ad6paUhuJwxGWo3f9Nv
9gLSN8PfNOABMGcFOR1W7DOBqDyjGqXWVHHTJeYSz+ZkpYbldXrL4DWZbBAqmbqh
nvu9K1r6aYKnHBvvIjFSpc05fR54oz71eRYmyuwzALtr7a/6jDR3hClzY7/T/rTa
heNsExNEyL0uErGb86cn1jQBDu1KglApyZlCp2Mt4zHKgLKr6S3h9yg5dOrm0Xfv
/66gtg6gTtGOy9eoJE/ZLilf9Zi3wMOxnKOvCdcGyqhql9CygM7oSFprOycUXvOJ
qCgmZCw539y9YdMgOxSjclFleI/cHGO3p65FNSefs5NIFypB+OGGt5or4aG6WEwX
VywhPUHbZg2SyWEngGqiS7qXDHhoF5PuoqMInANIgtMEG8GiXmrQ1xf6YnHRNf9O
cWFdVGV+kEfyIZKBNY1QEWYchmoyEAz+f+7sEPFVvUkvNiestLhgpe0tWAQU2Tjm
k+IuAtFFZwQbXp/E9y5wAJeVLlyKOPv9jDkc4FTmrvhYZNtnSDgCB1IkTihUx6zn
v+mEQujnKfdiIJpRNOtvDsyPzfJQAivcC6rDWT5sbHD8QqCRZ/UhPsGJb2heqlrk
jQfgDPeluMX9bEm9CVn2uokDTF4DyCvCUUtL9SFLXTaAcZNZ9dRHHDIrSxCjGsTI
wA0pvoPrktQg83pt4mnThPO4ri7JhOJC1nQCW+CCKQJ/WQJWTN811xsKoPQ/oETg
UgL9+glZIaEAXqrbEiJ7lxiXN6Nmp78WypkVnnpDipLT0i+DifBJZrwbGmtVCD7Z
D16XAF63B68CKopBMsI8IgGI7BFHLyhxHn321pOtMWmuW048xj72+5IGkHvc0aEJ
+EFUO5dL7lDCK6qMclFZPcEra6kD9PCq314Bs77EEaUeYncCgFy0RXnU1vFinUmt
xSHGiB9YJZoR4cuK9uMtWimOvbkbV4RHKWzMQsGU27Ixq+hCn1LLPZHkLr+QQjC5
PIs1/Fp51ylqu7ZwdX51YJO/TNlMJVBiNJ4xGcsybx+IMg5X06S7cu8bXUcCMftG
DGhm+6GEgwKTrKuI0YXiPWVhoQK+XFSgGy0/AlGQ0SX4QFLWVm95Fq7coSgYh3FD
yh/FuBIBFtdEtBuZxyLF0GHXRIVu88tLK6hZ7RtZAqx0KdP2ZGUKJEMfBAa4mVwK
+GxZf4iR6E7A1oDzrP8AVg8PQ5SM3GoP1ORmmQXgvJ2SzztjcjGTNfKizZeLYkYT
OLHZk4/WDjA4mTG84rIbv9kM1X89Z9fw5D+emvH6CRL3++1PLo8/dH2hvKUFI+ps
YxBhqofKBz3FAaalRTM4eqan0vwpGs8heYhyAvw8MJGRsngTWinl+ofdaAehuRwF
1HGc/OxWwsLippYeJPPrar8MMcBRCK8PajKs5IZL2IOtb4q8gJAHoyKhpmV5haiz
IY+m83zCDOzsKDvPe9UDL0/QZMXwpvJJHVWk28/h+y8fsKvVJ738byDRFVScsmsS
NyYORQNSNXyse01N+/wDsN+I9dzI+Ns/wUoRT8zcAytziH2gsoR4zDPuaMJgSqBw
tznsSJI0i6I/cz/MKJ+IJC6l6Xs0nsa36VTzE0Td61ym2kn0b6ac28Ef+dpyKRm7
ln+8/gDJsfVIR4qqQStzxUrIycKleCBnXhbPN6yOnEb6z3gJP10R1krRuREGZYyH
J2lbLko7QL178vhgFtxBdyeKSILTBd1jYT+X1erCXvI1FRVIUrOvSyWi1fHxSh/R
i/Kzq1MTXQP4oSPPVK39g7a+viVr+QRLZXTPP6o4AypU1XikvktTCNrENa1SkySF
WCxmaayWcv2ft7mq6cJRB4B4qy5ddlU8YkPouQ8CCpd3nCuyRyDc73xRNVrnqCSV
PBkrDjCsSwG9kXRr6lWZQtgVdbO5odsK4S4HCCAR1WrFkxBPlGOGKdQxKgElab+I
w/P9ApXD28w1yg0pQyy6zbRiTH1mz1BnxUwZPJ8g+QWQw5clfxv7fdSaiigxojWE
WKvFgW2e0B55W/YuzCLcEjdyPNT22984l8lGs30PtIKJYLXcyqbHRkhJcTetyvk7
RM9bzJx7JHEh4ve4RUJvZ3YkUcxaYkLIxzmJR4y9upg4e8JToFjKfOUn6tqqQ4D6
aE0tceYfdf5PXtX/ICkSzG/0NkDcXaZS2XyxfZWbG25kaQ6x6Lc7lVi0tSbrV9BB
kPUKCWm+aGHdVzcAENyVOu3/vRif/7OObh3FuPYGmboNpte1sZVp7vjGyFFS/2dt
Ty40XmOkMuul1kMuh3/itDWYipWbjw7/Pur61OQNSRPMfoRb4tzaHpaScYmBb3Bi
JsBH5UMR8hyOjoQ0o1uDtgxMCZcs8+KHv6oW/eDe94uAF5x866K94a26WWM2Pd42
1YzZf9RxNA7glMzKF7H0/nWRKaULFYwUUQgRuJU6lRO2HSOP8ai0vqm6VBUya2Qt
rzzEUJ2IS0XFw+74PRHRxAt4xRoQq0NPTGAfJI6Pk9yJKD7arGLGF1fzckzg3005
hyJQMjF9fGTpM+2A8S7hyGxPr1MvJboto7dzo8lIWxyRegwITyuLuopWyydq219B
Z97N0ToD38rtc/xeW0SkVLlKuFaN1K3i3KsBr9LPd+On0ya1ThNBb3ALYYGDKOyl
G2dn/phwtVY3bIoss1eDyKhK1ti5ORybwyNo83y43uRs7Jsn0kOuwLLjQl6r84vi
BoAmiY3JKnc3uOv0K1ZCTlfX+0cjh/pQfcR5dXRBob+XLEzp+nEBO8uoD4p1DvXM
RcCz1S6v0AwlhRh8paoqzwrkXnHtKRZSzU8uPUz7lDPstIrnwPzCYcRf7JZaVBFF
IPJ+6WXzLttsCEVSzlBuv8WMHApGQlMh3iv8eFPWHFPbpUR9ve+dxiMV5eQn+8pr
vMymXBlYNBSzJ40B/UzW/kXThtLvKIJ2xfKcHxsCu/qQdp2YChEIs0xAa9EyDJZH
L81BvBNIMkuy3xK/+7H+fhunwG5BqepgJOVKTZdE/ONIHnjQ5KzB2o1IMsaGw1BX
xAzbCxHjvN3jmzP3yrsmU5Xp+ZklE3kxnw5OVp/2/q//7vG9c7Oy6KAbiId/mep5
tSEmcZnfoJbJa7mjIm03u7DNDoCE486k4KnxKb37rLJ9UQQO8GWnlGkcdOae2B9e
2CpexRHfVUjw2l3YA7sYtEganX2AyIwTpOTUuAb/a7nFNzPpYeUR+B/6jOpHPcbk
arHf3cNLm/DSb6raSnikIU5DpBPLCjFtgxQWHWB0tYM6SWSrttIFLTqe/oL6596k
dCQQoYrsq45XQ/LQ6WnFLmcwKzrb6gJNbbkRxexXTtfH+HsMOS0BVJTPWixm8KBK
Mcnl7vAWi4FJaNoXpebHiEZN5MCjm4nPujCgcOY2qXINb57J8b2LJSHzB/Dj6kpN
Tvekf7QDO9ct54DJyURM6W8EnrrFlRc6PNVqXSGtWyxtJWkeIcb2/EGoEAR2BBkx
Za7p9Rtjqba3upGn6plhB5ZPX1Gp9nGdN6uzwggMeqBvfFRW5RbuQoPDCIdYgsiE
iTbtfbkafWxB6yzAIK+qeyELNtD9FjeD4qCga98Dq2u4O/xma/+7cNC/6wLdcBrv
zxu5TNYvsAEvEje9Qr50l54mDswIvLXYxg5Ag0R5wjivxS8HkF2fg2w/I/1soOX9
6/b5AQ+YhfhJCn6LO6MBMfUq2G9GERZBcTIDYwa4nZt3Nf4Sv/GKunIFOCzHPfvE
bKpx/pPkCfKJSkHWHn/Eybm9bNvCdLTIRrbJ84qJDCz7nX1fWLDNbnR52HBoZNhQ
1HdczVl4lvrTjyfdnISdaj6efZllM03MuJQ2CO1PzdleRILSPw0bl2T6/rrsNar8
HG+18voqUyeNcfrEk+t6/LzK6UzhdI+XiMjfuxXh6hHR0bHGOqttW8K0KR7Aqdbu
Aciog5KqgGWeZb6XL7S07S/vMUPDTG/Cg8gN2xEWeF/9bfUlD1Eyi20pa4gpvhNU
yu5mOj00hu2B9AV+UzTG7xd42w09R8F7Nv+zW/dbR2MAfOX+v4W7rf8HKEFLs4Vm
EvEtLlwwgB99QOKLjnPKqzbdwtNHhjM+PZtkLSAhGF2ypQxay9CVxPV+Qm+p9u/u
20oOLF9XhWt1WXnTvsRq6jeVmzu3oASoMm6vt491gZIhjyzhntT8ssUX4XHTe3Ex
ogWYIaZwySpkXTd91MqeCK/uMT9eZwt8d8COgHXVA1rcy9ILeONtuRAowHkKiN8s
KGX68cQ+tvJrqvxxqZge7/UlYGnli1o/TjVrk4jZDhUotcaUm4iHI3JQiP3WpucC
IRaH5XpiXuYRG1KVihf29CYHLxB7EDMS/VNLKgSAx045sjcrV4g3GMjP36bTswYb
1WC2KPHurOcQy+bkZMEB2/jVn7r6PYoYMTaLezrXvfEYI+jr6NUzaziCZeK3197L
KdqCLDaiMrdSp62KTGKPge9OgaX2rV3nWWiwLgkA4uuwtUPqAY+Kze0FC/OeCNzh
cbUkRpbarDEkeIGafLOrZtSWulZEiyfw29idB/7KK8nLc4u3/5WlSRy1HPJ257tP
59P3zJZpm4NnS5TPa/Ux4n/GNgUcWb84RLBqJkiaKtH4R9Ae/GbhbcK0itK/AhKh
zq11+FvcWGxN7++anuqnhbTimyR7duPgp9mPBcRAs4a+2yT1QafyvdW24iDMKjmb
AkHyQLlvA3jnhIIRmQl5VAw3ebNQ+PBPnU6ue5ys9lDbwnuUfF9hsDHFFvUjIT24
fh1OyqIAoFBgMaGeUMs/pzcqdbJD2nivlsd+9iWb2om32BMJBwORaaExGf0svGj5
MMesMJsmxqoCrzEbPAkP9cfjbLmB/EhJWUPh1moPq3FewKow3kmCSz7beXGd2ntJ
WL0TRXY2T/wqWCdGPl7F7+amXHKjKZ0fdYS0ksG8hrXIYNPqVk+JK93S+2MhGmSy
em9uTu13EW8JePjpS5F8c3ndPNIf4+6cTKdv1mA7KoFh4nAI833I1b7dO9DBMmME
ay598jEcTmI0A1d6mrKy+nHpuMfj7CHg5sV/vBFbAzCJjVqclnUyoOBAf5lRr7NP
EF0HSY9ttz7YLzwAZsZX1Chk67CWqAk0R+JVY9AqYcEH5iEAFAUHAQpJnJuTcR+0
d9aXBzxj1lwyiJ2EDczIiY6kbyka3qYvWd4wCVcWJiIUAfLGE7mzBw664paqDVbi
rD4a6KAHdDLQ1E++KdnT5VCazk00s1tmrnAUnQQQ5q0FrJadgL5zTYjs3YRGbMZj
XZzyvpyGW1QceYJgQrZAJs3hM/gn5iOXKVAQ2S8ml72t38Abr/WmNeWtu2mhRIxM
jUsJMV6qL3Kg6fIV3xa6Hk0+aZ2EM2BfBzMLlLuJ1JAGQjY9h37ELHD9ICw7Oph8
Lno7R6bH3/echuN2S0gJWRDu2t6l0Z078awx6y27z0ZeOq/pJBxbF2wMoPpUVm/o
MAbl0nkJTq8u3fi5GVceJVDK+wHfO7E70FWX35HIR0RH6heNyBgF0JUEp84KgrkZ
df3heoIwmVwCyZiFZ5dGpqzFj/TZkOcaG0D41THviCXQli7WvhrEZJJ78fsKeJpu
/CTRUxJ0yU8qBYwg4cQduQ8HkjEF++uLm1TQgc0yoNhdhmxx/SZpOV4j5ZDtwvUD
l+GUyaMf0+r6z374T/eKkA+HgO2zd4GrKJnopybTLd6r9EdhyHbfZtQz/IgOJuvO
1UpgYqkVQdm0pDRjjBF9nyrCWwfIihc25gm2aQkjYhJESnIrTpxXnZkIUqeNeUKW
76Q/Sa0SgGsgpbOev7FjAPG6pWVxakyysxXVieIGAX5z/ReZYWqfm85Xt54qPkjT
9wWIgefDqYDprkfOc+aNMSxHZfdXIPSFygp4W01lQBeXUjPVEOc5/AI9wfqfi6+e
4oe6vHFKLbRG/aEsGviVHse3qREJiQqMZYaEmbwgnhkqJ0jhLySzFMm9Qgh/CTkl
Tf+h4cYhnlOSAmGlHgtLoJNdIqGToO0LQjOsezIeILZY1R9MiqyfF+Qd7kD8n9nr
C1V8WJws0c44QMZ5G2baekdISPuzL3/qcfNeu9Opcy1NtQ9Z28thSwI4OZ+elQ6P
mmkSTTsbW4GRDKoGS18JyDIs4V/ZTaeaTL6/Ln0/lSagsBnQAiW08Sas5Ba/Wfvh
jEStSx5cLFVNKu2GSJyLdpmgDG5v5bNQ6Szw+UTA2jx25IMHZwrigGzz3gw1+1N/
JWW4MG3mTxj1o+Mg2ecqwbt1/yfi17tgBg13jz+VkUy9XQYTsLXTvaMpAUblCVFN
blVkX9dByp6g+IFVLaoOUDYi1StBcOKc3HjBcAXV+DCZiEg/vAAwSpCkoeYbjoo8
NCQlVkRTko/E7PaPV+2r31pBYy+1MkagG98FKUyyyIcS/jt/ii3AkwT+FEwX5BTG
fgp+K5DJ8AKx9CloweU51I46GGSmDQb4tIg5gzEqAD0C+oqrPFP0AjxMuujDYvce
aRHWa5B55ubdYuo9vLvtdEYTsLVbcEXTi83fkSAvdSz2ttfwyAIhkAXKZ74YkI2k
HcxyS7yqo/0MJGkxEl2bdvMRnKfeALFDbCuegvJ7u1SySFle0gMUe4zcB1Tn3etk
XctB6FOLWVhTy0k9kbak0vk36f1yHm+GkFDD38H6ZtToUbfF/IasY9gph6dC/c8F
Lpi7KcAUyVfvq6hYucTTIGFkKpNL+YqNygiHa4ZXz2hn714N0nH9B/aOFUEPZGBv
FfvbLFDj9TtbHlS44R4XzParWf+TV4FoxbYHt/b8AMXZYjBGcjYmotxPLg8Upchk
cczjPR3FR2cDeIpPcx8E+J382AbaY/U8IcNd0dvejmSbbIsqSfV5SNgN9EN7lclZ
rKL6CbhYNzWj/VmHo92c5W+uP+m4oZx4MgOAbLGCkQct1JUDmnZ4dkWoDTAmdHi0
gG63vyy5KhCIA64IAKxcUNg066CyhaZr8YGR6WFaB/a2bYdzI63btuoaci06b5mr
8ts+Pses5e5yMAALsDHbcyd91dsNpO3BEY+yRswkxmxxatLlP+lwR7tsj9Wbk75J
ilqJueId3KDY+PJFnTxpRHXHLyBYh26SLDezXeYSgegHo+gyMcwPu+mmJneyvVDi
RiabcwJqD0zYY9Kjdb1c4W45xa+FXFe/g7vglF5Ja+9Dadv1TMbzMW8ayTFByYuy
FcGF2vcyuIbgPE9jjAs1VvfvwoaqOdysxJqho067yLigHVAH0efGbUMqS/2X9End
+QC+F4+/5SBhoM8Aj8j4/g1+0YW1k/1YjlVhxKGOd5nd9y8Jenv7uQyO9/lQi9FI
qU+B2PsiE1s5suAEzK2bktVLMuMAkrS41+V8S1g2LoF2UHtLSZpRP+jDKQHhRs03
XeZJVVU/Hd8hfw/ymNqJ/SlfBZc7XpK3/NGAMaoZY+UOV5ltQyZOoTghAcxzRuKh
kcrBDhiekN3rnv6GzK3ZjQWuCWb1bSv/vfbhFG++2aaiEJ+sIS7xTluZ5Hx+ghyF
vyLw8Gb4IoGJcsU4taJX2H+eiYze9IkhPhv5Wn5kKy1HUmnA5uX5BjKvI5TTaknz
YpAhmeBjbu7WmYRRHpNmO65IHTv2pnuJB0qvbgvfwx20zUbJlBBvMrBuewhOsLxb
dD7cNaaVfU3lvImmd2NAbkoxQN15v9vB26S3yWcnP84cPysxIBu7X8zym1UfHkDc
4gEeCB2bFnj2bHiZOVGcdEL8ihpOn4wo3zu9hRIb45g5suwKpz3z9Q9ZCInwg+EW
ChrnqY4tNAQqtHKVUgMMAXOtMpWMvt9CAmQOvPyS1W5aEeYzrpuoZnWNrHV6j8DE
RgGFqkn+N7huY9ycrSIB2Hh42B+ALocq982sP56JAAGTulqHlUaEqoI5gwTi9rcX
SnChxlJgnGoQl84kvFCsfgjEc6+zkuCU3Ayq4tjsxCDs5fv75jX8ZLPLSpaU97+N
k1OMHIgTdUzqagvLEtfU7iNqRTpcYLrrScJV5uAsPJV3JZwdbKH0L+wMDHcRgOSf
+OgX4YWj6c3znSs1y2wl03kj0LQm32KCMk9CRTxklcUPaBFUiX4QmkWJIvxpLm6W
QO4Mx0XqOdJ53yuDv8QEj8i22kBTkzni/HswCYNb8V/g3ZMLFQVhq+QL12fzlYjs
1OCJXOpG+KtBtJ4kF9ZoI91JIuEtwSFwCPGpmjpiBvytCVW9Zq0NK0fFPACHi1uv
sgGsVPJsD7u3+xvvIVjQViaMiAl0HDMiQmZZMWA86xwIjhHKwr3a/8eb7Et3BCrR
vMghPJE4L2IZxYMROEYYhCZhO1ql1q6IJ1/XB3wgveR6yMV9bdRN/EekJPBPujhZ
QOVfgkm1WkNXWSLbD4LQ9laEntFoWLi5MTIVRjLqMSXYPAn6+bgNRYtq7RZ0QAjF
uScCF4kdSyZl0GIUWfmnyceXvucMtHMlIgCUtoB6AIyYxFvfQJXWfVdlE03iMn4O
SnPHUcfoSfKdQm+ag8lgQur0n2zUSuls4CRm0FZmKg5nAcKml81bylpoFRCfQAKG
cBcz3Zxr3I4nBFZq0d+as0eFVNfd3BAe2CM/GjwSENtEec/fIHAU7MUSzdlejg+l
ExllWz+708EPtNENzccfvJm2rtgU9qIeW2JVS17F9kakI1BzGiGsmkGBWrWX046B
E1EdvNxitEF2UMJmphGSTeYKmhLOg+WuL1dRTBoIPjfT6UqdeKDNNXNZtbj0x0H/
8+sPDPFzOyDU1aKvfdvxSgBsGS9c84Wh5tWNZnf4j5ySiw5FCX5aoWabCyUcdro8
INH1amcY9RjZayjpEgf8FQGIap4kE7+vCTzUYuz0pjBypCBeX0WOaa4n8s40/i+I
iR7l5OQYMFW0fnqyHQZx/yXQ3Zk+AOb1jzhupxA2wdMMBZadPGBnslDfjDfphKhS
lB/Lr1zH035J6fTFx5MWBLNtHw/f7VcQlO+sVAd/ixEfVXK4qadOliwlOkPRV/Ln
icW5bkxAsVxIAZcXCYntA5SKEts/8+9jbiHkQDw5nEvIct56glK2NcOVkCpV5tDj
jnG95zC5VYxm5TXJ34CUobP9Lel0RLUTD3jKaNsuvnivC9BwPRlTDH+J/PmR4Lny
UA2TxvhUZMHa4AmD2IfyaCXB2fxDVjhW6jm0ghsIE/co/GeNCN81ujy7pePUzpbX
YcxOx/V707bF9BD2yEC+FYtJNlBtGR4twImnPsSijgGZrz5lGZnSyeW/zUzvhXvH
TrC6+F2aQJPuSURkfSa3NU32+FjstzvDDOdslERez794/8OFKXJOMGHSyZy/B4TE
hHV6bllGh0HeR1Dpmgo3H01Snnre5T7HnkCWYCqqon96P/78wQ+jQT4/AJNcnLyF
v92Ro7IzdFTxtgdznSojKOpw4g19nBLp/27KTeFr0hdqvQBVeJqb0sirg9y9MZ0q
g8DNMGDgIsK6n26cS7aFex4dKpNPB/VAVJLxfqS2UqTExyItc81TshP30BBNAf8v
AY4VaWxiMEsCWNh5/B2cAyb7Y4B2b2JXh1T2WqWdvuBraUnkczpmY4Vztw4Xy5Ab
1pSt1t16D0KKEVeViHWJZKy/XKA1AF5nq94RTGgYEoR/E7aR7H85JlKMgbNYPXkH
NZiz9zaK1zV1sY6uAPHsH7GBM3vmCbIxGM2t2n6eTyQqZD4ZvrZzwB4CpbnOTuqL
t7ey1UszfEweJ375trf3HRQzqHulfZaIy7Fc++m+MTww3VQWPf3b1wMm+1wI0nZO
ON3mD30Ao6Dfxe8uF16rO80gEvoGWbV68wo7DFyaevLQTNBvnYoxqBxMeNanqNDi
UJibxi4pMSI31kx6q/rTXQXHYx1Vo90XSEbLzq52kNM2axD7K+LdYZJMtj3vLFTO
3lBbBk3A0o1LrPIqhWOE73DifZs9se4YL0Jfsqnbff1+zW75rtsKATP1ZAdA81Qg
dgNVhTY/rXHO/Q/qKwq0iuR78X1d9Pruyx21QoJC/iNatOI7zizvnghyNKQx8oi3
Pllhq0YE87tyNQfSIw1yAP4+hvB+fmRxnOr6/5C4kgmbaHb7JTuVEXpVgdw1qYsk
OuHk26sGecX1EnjGlSJiMxj79cg3O81kYC/f1+Zp8DOFL4U5itQcHYmZXGd/u6NX
E20K6HQznXRQwSi6tIGGT+DGtLtFbUUGnhPX36JMza6Ww6B+SE1ykhNYNImTu/om
1TH3ohnU753zaAw1JYb9olFKDpEvnRvCc78EKeQKzOzwgdiPByRAt5Xf6ROrEM6d
yzei7t7LME1n1OrQ3BQuLE/GsfO3EtIVbx1JHPMIotW1Bq1HeSFO3aUzv+P7y51P
IPzbFQLD3E/NSV83FvA8WuKrWfJ9XZdrP5r9PrEy1CRtoB5mXYqjASGDlkibsxVa
aMI8asnrAWUv8Y2ZbAlLLSbHZAzNMHtemtN08VCMTIIIHyoPjUZA3Mvg2uT0Je2Z
gOXIDisukG1Z0HXrmSZKqVGcf+eUi3cNzhG8qzUCCq2tY+1LiZAH2xKk0cDcHL1C
RDJmj9W1kVsXgQ4IDKD93OBJuf/NRQC70DrOaEvZXnMJMxXxqEGBHgRUZ0HAqX+n
aVT8NLH8Y1GyeaT3v/MpSWxGDzj2rORKz8jeUFzw6uGM3BcZKB1ZjcFqzk9EY4GB
b1AfhQLgg/KVmc4KGj8saXe1gx3FIdET57UtCortNJiRFJnkCZMx8dAUp68mCqbE
c1++vLw8QX1V0eDwrAIPaRVcj10BJYEckBOKiAwAaV2QvA2k+auZAH9vZ1EVITRM
FOBjg0mRWX7pEkQdXeslK2kc4p4iTJK/OEmaxeCM+kFh1jWrzYvxqQR527m7x8Iv
sz5bY0+HK0Qq9R/vKabFAvTBGw05WXZxGo3/oHD4vUyoxCIZSKt8zGjxFmv3DlBO
q7NZKcUW9/9PO1K6lAk1XoA1FV3kx7YHGW/mxViDoSVWw56Y2ew41+7mLvUEGXS8
Ck2ruH09zbv9rPfd+Z9RfkMRaz18VBjSZsIlV9pCRaxxdv1KFEITC+8XRhhis17D
lBrn4mTkCJWx1Kdg8t190dJyA+Qlq6BYRT6OSgY/ok6D9l06fy+h0/2ik/S3xwEx
dDzVjdGu2OWJdwqPUigE5nIpRI9YwCXXfK1SpTJ/nlk7gSartnwuaLOTuujTYUx+
7AplXWHMEf1h4TuGwNbNMFndHntVGRVIYkTDwjKMS7u7zk3n1GzTuKcBhPDA4wQt
D4PeXt6llfRhIIuj4f2H9BYQdriJGcgmbQLGA6a7kZYPJwAEq1sXtiNLLi953QXS
5Jmb5TGtqFiYc03Zpos73jDq03z6pHBipmNYYZcM2bu6Qx/pRwGjOQC39/LGgN2J
pHWG7gm/NByicZ3pJHJrQhsricE+T5GCa+vyi8x2LQ7oU0EKrY1/dD7vM0p9L25Y
hopXzAuugcgvzJqurmD+/ZFX49xwslWgbqyofgVeh/K3044Ma7OIfzgyMYMEfBQo
uXGkNE0HX6OEmM/qoBqh81kD+zylUU5pCMkk/I5WzocPdpHiV2glsm2d1wbXxNOA
on/sRlgRoVD5aJk64WnPFyJG4oehZIDE6m3/SiLW5uTDct4v59lmm8Hh0z1wSOa1
GDzL2gsgVE/N6QFVDN/g/3acKi2sQVN6qbaMpTnK+/G/VLHbwcGgVSFDG5eU2UyD
coZiW2PPO+khUrXkey10q+z131sSO7vQIsYEE0lA0qZpE+5N8K6aobHemKMvjCUy
owdA3tFunEy/tEM2VMEDQgnCrCLJJtVc5OJzWHjWgzaTWeLZklmMjFWOw5vmjwf/
3AQdkKspmhtrh4TLf3P5EdEvYdvLu5hMkltC+GxiYeGzQwNwoGI6fMONNxm0yMF/
eCg/W+9J60b8ghnVGxVMXu8WDUXozf4mIyPjf696sYshJhEfWy+94+tJqqe4hjOu
4Yy55aOfN7xo0mV2ZFyaiCP3RHwXKevZUQJdlU5IDrD1EXgZ+xpce0darlc3q2Ka
HJJr2ypD50ZdynE9c6aB9CDMey4r8aVdS8VF2MjkjEAQknnDz0bt87PT6gl5Kqe9
cDxB+/eWpxjr/6n6OCOcVuKfqboZ4At6wYM7QN8N1N8dexbi3r3zuTRA/sXohn8u
ZXBl2yoZIybm3iXKC3tHhfRhhPCWn5uo1whzsdl7MIpBW8oRtm7wgdGsF4QtCY2X
zG9ZrqwifQM/umIqms14cUtk8UCLaHelCy4HJwCvMFzVVHoT+/CVEyp24/YeUIOl
asNXUcNdn1hylpRKXcQ34xw3kxsCSf/TeuP4djrw+G611C4+pIAw6JwSVhQ9q2Mn
lcWbm5m4KuXZfbIwjt5vAreXCTQbi/XSkUqiwXXXl8geU8qnL+FeBD4XvFfvFJFL
w7JaqVNVBEKnQSQhWSYUc0WdLex8vejhWhpG9+ZHDI+s+ODIp3LS4cmPBohLnVhN
CIMe34Lsdt9AQgXwhT1cXiYf2JClSfN/bx7fkLcqa1OAuJIGhVEPBggx3Fu6x9Ep
1rxZFgFkEd8rrFD4johOIcQx1OPYP+gReSlAjbhNx3nSkHNLcEY62VT3hEyWr7b/
TdPmMQNh7SvqerAFKlydXegI+wgvl/fng2pqBsN4E1nc75cabv/72al+1gAQWzpa
iFHShuclRRLI8zOlwfPIR3Awgr5nWEHVuLMYQYProKiroMbcnrSKkZr1x/JsiCLJ
DqKqraVgKztfwUtaXXFcS7fVfjh8sK1BBvkfO36AqP1z+9/mrwoREszHVrS6KcP0
cqo+zyf7I7WIAaFRs63p+WD7PuMarVUzjw9BCy9RiS9AtWeLWml2QMjD9U89acvE
ZPtsmIXIGihDhiDnlmSMdogEFds+YSkZvKd+P9GQn/ANY0fjUKLwXYUJDR7s/NVI
hpAuXUIYRStalBApmA3s2wKGmNSvL7oMvKhVLU7UDC6pklr6NYGSk+Nlh482VrI+
eRDraJ+zMln/JKlAW+ZcTlmH7xa03KPaEyTl5Ky1lEB2sFRf850zUNDa+/HxAt0d
wsX0XELh/hhGDfi0e9Ruy7kzePlE0iK8/Y8EQMakvzlPqveeIa1p/M7nzwXORQSZ
FW9PvGCbEn/SEImms1oYJUol6AW329kZ8wYHvwe7q/xk1uF4DCYGvcVZPDab6aFR
MEDaj6O5J5dKX1KkBtzlkFGHCAGAUftugOFFo1FS5em18htiAGmunSEcGSMb6E7Y
dvOlDqOpHacpVYfXs+f68FR8Fosh8cy0I4EO4mUIN84lJaV9rxK5bCc6CA7t3lVF
36U6AKvSrvNZUy7qsVXlQlbZkcvyCQ0Nmf7+LHWC09wSuPumcLQVc/Wip+TBV+Il
TEbIGE3i24B3c2m6WNDePR1MN09I9BEpgB33dYbc6op4ys0Ow+85dkJ9eHXMhKnZ
OpnAPOcdj8yPFepI78io2NjsSIsM8r7Xctx9wCoOKHIX63qFRSQaLRAc5Ut5iPYi
1s9p59UEkniOU+WfRaCTCiTks8V0uwuSSouuNTvUa0ml1H9mr9FP+MxKIlkB+dyb
GANokIBHWDDaZQgAJ+3IqONBYcl7qiliq9vD6ngHxmqqN0V/tKEiCK1qrwXRTplg
TZ5vXtFeZ4ZvZe9UcwLD8b9FlQL23qG1J8OcJHs6EEGbfhQxAt4axgkqCJ+58eJi
jevNm+G+ValtaFCsq8IyVRq4ADNYCyV/O9ffInNygDABSZ8HozWuNjtvGao1FTnU
ikoUxRQ5mvslbbqW7sM8KApDxHv0DnDPZrRHEuU+t+/Ryyxc5TstS+HxD8tn4IDt
4U847ukQAZJPBV4JggD/+yDmA55ihpD+P4AotBpOtEdE+Bwdeh5ltiDWGoT5TTeo
OPie1CicjfbpbaTmwc4GZLvdGwgaSoU1LDyBUnxvZpRgJ5Y9liPNhilMNByq1RZN
J1gT39nz+gEAAo5uOk7NQyWjDSUg8Lm37yCangULx7qiRTay0SZh1mc7C2RaJiAh
bfdkLCZkMNet9vpdqy2+AAHmNuJFFRWgvI5pPphZnEFgtL+lV/ZWPkaQJKv1Zxv3
dqLqs22bg6yAGz8s3auUDj7JnwWDzE4TQf0SyYL/sbdoOJjqmbEhV+j26WPntH4N
91ehBHCgWp3gjXLDyOQr/VY6ewgzaD5OkFmNhs4F3s/v1stRXaHQP0vKyZmU7Kb5
yZPPS4++0sYSGJntqcsrGiSyifeKkJcBHNjtZBEQbeaxaign1BWWftYcY/OqDnrs
JtyEZZjpY8ABkMBhfHB8Rv+R7ioxamNEvQaV8Ih3uZA6gjO5mf5I3DH5VFSw1cUG
Uxs6adHQDkRYuNwm3MuG1rvefEk9drV6e3jS6hAjjWwdEPPNxCuqXFkliljvsi4V
15PgTUO4sWn8Gq7NdoW+LXhullGIgivuc8oGBsXcjeZH5mQyxVY9xdLFt2716QDr
GMF146yVPo+8LbtpTO3awPEVqRZ2M83YJPE/vsiOo3u7nZds7X6MSTBAA2/wDL2G
6aNgiGWGGSRnVRyOAerijHlJzAFnjzWYf7FcAgOWu08l52T/+vBP7WCnzD21Jntt
wq5iFNL2jLh0MyM62Q9gYpbTcPOfKG1M+aaqspFYwQazowqFLiR+VY8APMgIDNel
8gm6aGz6h0b4yXaKqzxNxBBG11ktNITRT18taehephBpco5FekPIuu0GCQ4FQFM9
rEh7Lq0Xpl9nGM3FMq0AjTx311FmGIp6A00fXG0GcIrEWYix+2UVQWs5PHLCMY+C
9jV+D4noDDz/303agsRqUMnyfcQb8lewZdV1KL2AeG4krh3ss4boYyTbKWomveEG
zInOK0nPPgJwWVU9Wkf9mBACJaRbk/D1LqxPmmwZg7tevmTO3NwzcvrGQpgpwWGi
WjfbnS8HEj6ZTSkZBbh/rIYA/L68hk//EOSn/7pKirZ17gjnQKdJ4kDTJJGrAQqk
9JCEaQqFynWHwn8KxJRom+PGMpHWkhkrRtLf6svsHFmsa+vv9ICKnxyKYBmLwIiU
c0yme7ljo/YKdijjUXkN7sKHvvHi26/Mp+inxa0AGrLXNKn0QJODTelr+NuGFslV
n15R3lYLPvODPSWmgS9pzJs3csfqY6T4eGCY57XXdkjoV4cDyJscilqkfCygzLNk
93qCLswvs7nhLgpt/cdHZPlpsrWeQDXSunQIK+YyObolfNSDmRdL2kK5/hl8E0wv
xaOJNAnFaoCiU3+dOoWeEeRkBdjr3ZMcAj/qQBs4CT95kgmnc8F+T4rfjQYYryUB
e3+EMVWPtXS3tBDljlQt3pE8urr+xmXBMJoO/Na7kV6gMLBS13af05nS97SjFHKi
stMCA9WQF6NaT9KA+iZ633jt7TwPMZaj6KE8cM+CTgSUhn5D+XxrytAW1BdgYfM0
NGmOvG+PpkFtxx0cYFMu8wv3PVguLyKR7QN5JEm0yXE9Ydw3mYpXUGpDom1qgfN2
8zAeizJ9vVvyk0/njf++ZM4gT7OM/Hkr9ncXgL8modcsTE8msgjWHrLszXNZpRDo
1DLrBjtXw1axowYEQy3UBZyJABe0AfF0n0s8YKH6NENZfeImN0gh/mWnXrgdlBFM
pQteNGlEcF8rBoAUM1tGzXfRg88A3DX0Vm6y2DBpVAH2o74q1O/sSYORQYwVmg9O
E9+YfEQ8pmx/J2QzG2mnZnVCge0Vcj7PU85OAJzZv51p8rh8600uBwBvCKBi7pgZ
tdRCbqMw0Qw3AfEN5LqFlATehV36x7WMZnTnkuDjQECzF+o+GsI9tmoi3SgsH87h
uUhbXX1pWdl0LTsNyWAcCFMaalIIlJpZgS8YCjdpu+a4xs4a9bH+0iAxuZa6FUoO
f96+chpr0zkvvN+McES0whGxenL1uPrd5CchAsU2w3axlw99HeEKZyUUcM4Uecn+
ZgRi/2poTU+wntfJBJ66b27Rriy/guWGgzYS81c40Se86rp8GlBmFl3hcvNno3fh
D89mHNwxbWNXZP9sCb6A8/6ygpc4W1OC81j1Ch6IT+ZsRxHrWVTJP3nDcHdRVfnm
dZ6aiV9dYFh/GZTJGtcyQWiSCza82++dodcC983RqOepw8bAEff5fn38EohavJqC
6BJDold12sYTvjaj1ceteZGxOGELsdMVh/R1oaeJTko/VYFtDbq93DnjxqQ2pKmS
3Xz5KW4wrWduR+YqhZc6NoOX6fsRAOlWkzGbmEaY3FTQvkYm8hyS2Ivu7elzQEub
gdn19QXeU1eOkcZHNA46FMOOpEwrMYtHFjt6kJPXvu8otc31PM0DhVl+kVb6xU59
I5Hm6Cnlp0GpVxUQs0P2JTggjL1qj/bca0seZEIg6jPECslO/19Kbg5GhPf2nWjj
i9dpSnBHDlCM8qF+ZtE0b66Zj/w85KKZDxKvLKTss4igXM7PsoCckUBhh1guFFsg
2rfPl8eKHfMZkrUVZOgbkj32CgPtFS62dNw3AHYAPxN/BxGAopJ/oK+s3F0KMcxU
Eyx2WHfUqUTwNOstsV0JxQ+pUfQpovIhfoEET95UErNRq64u2bsQSpH4EzAJqM+M
l998TbRWU/9k9kjPEj1N588HlfLzbojOSeD8d+N5kdpZgkAswuCxRw0e2QDUP4SK
lJguOUMDmXiHBqAXpUBXc0R5jTKbs7DDYwCbOwb6J4Xmb0GawaZasVOQmGgNVasH
yRcYnywQASHO89BCGlmV27bbiKz85BcQ5ifoDRUZ4b6QsGjYa1Pf5MB8i+IuYdoQ
dn7lCSo1N4Fcsoic/jLu2qKlAxM61FeOlvN7BRLtbFu7Z5REYDsNtOK1yIQ254Vp
8AnQJYkvA030qpXJybAtAuBQQrzr/xs1QokRzRoTPKQlDD9kroyBeGTuSD/RX3tu
daX5YMjWObTkUNGaG0hLeCubD36uKH1Zi+N2Aa7itScN0NG2CamK/DI1feqwHf7t
P90bQfkRQxOMpRD1xzhmsN8Ez/D3mrUdMPa34NjQALg7aOc9FGn9Eyat2pb9FJhc
HMkH9aUoblrlgxiFAFtsyawwCT2Cw3sIfqj9poz+Qg7bzhbu0oYm2Z0JIparXiV1
GCDvyRwVM07RM1EO0K7KQm8b4aRu2p3LUxOnwNbPFoTv2+SKIrmm8A7T82yWPeRr
CnBCxfxh9DBxEhXr/UHiponxYC8ZW04hVsh/3t44QEb5Fvw1Lv4CA4B4vdJQRFLM
Get3KlEbO7nZnWlNey2AqyoVvTPrzVLcChogFDwkWLZ6UZAfSl+GTYm2exxmqoom
hsPnwX7o5X2JRhF3ANZiST4QK7X20+oJRNvhHEkVw1nnwMTCSH3nYWI29uY4oBSo
LElWq5SB926CxJh9h73px2d2WUVREgJSRipvanm3W8TE+lB9jHXJmxsS5o2fQGoh
gYgMD4ZfbNQXTEFKerkU6xjzVT38Zlq6kewXaOtXkvkkNbigaYSN8d8+bdT4sE9X
/rLAF1x/U3Qx79K0KKahxT4incjUJNU7JkwvrmX4cNoD0J1Zh1ac4Qt7IgLcJRl+
c6kSkuyKlxWxwYZRsKLHh8gjZG3QZNWKiOlUf/nW7xDqAnvjvv4j1GBw1XsYH1gd
8OHE1KyyHIi9Y8xDmwzHb42HLdNpf0WXhNs49f758pFrycrhkhanJtpcwpaf7mAH
B1T1qzq0DutaErw10PzTtpE8Lha4uGwRmpxjrAZ40IKGrtOI9JMpND38LFdhX+wG
eWh11OVhchwevWY1P/jlBnwNDNVxWT6qP9rUcBlfmelsoPI1/P4FLnMuWSQgXNVA
Od647SFKYX5sU8cN3U/Uq4djm4A7iCZd6BnSUKttox086HXD5k9vFi9iShp8gatX
st6GI+tK/RE/FtQosWpXrbwwDfRdfZ/Fs+UzVf95y8j8KDb1sZ/I7GYWKHWuqfeq
YktTF4kDWngTkbQDZzTDkBpz72LXexTZdplgTqolAHhcxNYlW9sAQnCwpctu8xja
5ObuGBRyJG2hxLYVFlwp/N6EFH/ojWJPZC9zz+0fDDRhfAGvcCFEQJWTRXDbc+8g
UOY0sgJJ6fgTfiUpyRBDIZ1QJB+CC4oag5mJE2cV/QCedu8qD4ayNYEk2DZ88FGV
Dq14ewtVTdIFlq3T/To3lXbNL+4H0gPYZcuEbcI6kQnGfKx9E3FKQKs2YNRdNavJ
axEhl9nAeo/6aPCF5domj3kFv1DygCVQoD1aLJ+VTW1OQrGqeZzgR+0bitEH4Mkx
+fSogtat2khe0BIAFq+lNiKPf09HUlldvciUfIdCKcTsUiafN393sxo7slTILeCA
DoB7CFea1lgmHmOkm6WjURaLA/sjgkBdm+tkDXwy+wpUfOcvYJsDZKYY+TOhYMmt
j8oJDWpuFzCOL1PRRyoVT7Y1rJlh85TlpESGArMECOBaQgRrENN8jIg6r2XgmkRD
YE35q5V+Fu2/r4d63+GkJQ5Gg1CBn1JyouMJOFiFFtPRs8L9M257DrIp+mKwiNAE
HAVw8+gLT6wKFNMLnj7BAJ/2lCnd6FjKLWy1VjK9kLDSvowc0movzjUPeS1BcF3q
3UBn2yg/b29CHyS7hshUAGB2CDe6N4STPqfElYh8Kb/iyvZxTTnJB02FcbtdC2EP
PIWhLZYc+rkamufNJLJJivwJD6FJyCyF7DrBQoX4+W0dWK1x9DvoqaeHpEhd4pMZ
N4guHLhDmtZFQY5YoaMDXYaMNLyov9TqsJasMjWjc6LfZwdmrNAbpJbYFcr8kcqn
CgR0Do1lZJI3JUIjn8TK/UAzobKXb8AebkeWhN+7/+W9cHSUErskGNpy1qIKIGpt
XnHbY5nnbEO/HQ8XvBhl9kZFVosbmq3tXbV5KaN5IrVBBzAp+npK9ClvGUK3zJw1
1oS+04xWaLWtTGnCTybV6umnS3hH0knOrwbJUtOnTRLLYREeC7Y4Ed02XEaVjTav
ZOw1NWijBQarNYqu9+kmrJyVqOUDR8cxEQVfbLcDZUV/NeeD5ev4MwSdx6MysLmQ
gNCN7fWBYQmiY4qg+N2gL1lS4oP0aSkDULGcHChHYzlepFNmMYW5WAwXMJKloruK
oyXJP+VTVmvsI9SwJAqQ6to/IR2R2axQW199YPbTP7wpF9Cluvq6j1Gs7UOMSXCj
cSySN9qhk9iX78weMi01rblkdm3pHPed3kS7tanQIipKJlRlieRWFCDX5T2zxpgp
r5reny3LmrG8XEsO+utABVoEZXtEXTEop8GgG0FTNV6yh5mEvnxZuUJbCHXhGLtO
osZesVIGnGxcQ1KwvuneFnWUnuWUwewH115sHj0bYez7DF3zzhXOZWnLpjr3mZXq
0CW8iPoSHCncYY/ZbB26ym/XrV03W6eXvNETFSNS5zdnaa0xM0nUlBmspyk47y1r
7dCi582bTLr4/UUKciWlXKWNykB9Fa5QoFzDPjStRgtS0NDj6v8KhBNUAokFRcJo
qkWGJdaH3KfT3cxvdsLm1dWfe0siACk7xL3oIrlPqs8fO0XsvaRY1lGlALlSS25r
rOF5Y3/qhUkdAu3T2KoZRXhgVj+J8rprwjWbc/+0Z35JRh1GMjZQZyXcYSDSMu+W
cVBgWrXJSutaja0sH2MRIBjFpAILq/2/C341AOFk6toqid/GjhbTf3wOOYnaf78q
3z2ayN6bIzIbO0FEFoPiPPGHV3ofByfgEMnB5HGtaKtwAfstNIQwA7e5pxS4b2xa
nYnIzs13U1RhxzQKZWkb536mmxfW8b+vlaXEsdq3zD79WQXlZRzWT1/gjevUNh3c
wmYKfEIfa8QMuHkvFfh11C5vTPdaWNlaIj/1QFoopO1rvuxrfGXBYmXh6cISOhZe
wk5tuU9bb25zyNtMUTyjIV2stwKPCC+i49gJ6x+keOZH29IaMAsa1iVtZnW2JR0W
FTgfkJV2cf9a5cRECxN9BshlcRpDF8rEpnq0UHKJX82ViE8Jpi6i4+dd74i4tAjd
0M52BF2W5hXEN2wE3ztIiA8QJVMYi9dQRVQ/0tRyf/FXBykRZm3kkHrNi1pFki9W
MjUwI+/hQ1ZUM5WlsoYvcrQbnawD0zlh9s3FLnbywkf9mdxJnxz1QGxuQeuBT/Bf
fLG34uYF1ms9nwDJPxk704gxJd+op/IdtPN9U3uzQrzvvLd9cX+z3wTfwM9ZC2lZ
v8AQtGjbN6cPvHhUc5SwYwasKRXWDUAtfXLH9wufm3CutnsfAd9AsedKNsQKeh0T
za8II3b/VRQ6Vm4vhQGzCyg/iQviVb9OepkwrIh0AZyhRpBffZ7q47tYm0ksOAEV
CxMraBaBpVF3LDn2fA8Ujx3KQCcg0JKJWzG042m+0+ealwPtnR9wvJyulz4sJWVf
ckXpVneW4BcrMndv/fCjjInWn608YgIFYKqbmEBMMMQSYVCDfqeu7c7blkacq+d1
E94xaaVVEgyPFXt0UWJYbQZ/E+YS8tfRG+pyEdsaMdcI0yx67E/ZWJU6B5vhdbNF
Wgch/zC6ArjqUdthtY89yM2wYer/CZwzgcS5gFzXVNTj8GNyikNUykWWJU5Besdh
SxrdGtvXUJAZTogVHSvpAm0gfHHmoNMcq2P7QNHudh+6lTYff7ecRNb6QlVTNiFD
TuNqiMJgYM53XuiNPSyxDSxkgzRBt8+UCNjYBkW3JgMtUcQGZSVSYHsto5x4soDb
RyqcJ5uN+jXBdDlLP9kpnixMEa0KVLb6uMVOdGdaATBnJBCN+gdzwX1l+XsOHUNV
PgOnqMPKuXyUxoUGD85uDp2K5HZicDJeqDZk+FN2UPWn+RqMuu37HHicxOc3OSR8
TB4avINZbFiVerKBPUVBRHlWN9Y5CYESJaMhswNkdTjIIjadVIPqZO4ISPMldV9p
CnqW/QVj6mV27FS7KOxnJ9WMGw5xXmWDAWHy0Ip+g4YDAEp705UEAEZEkl9/BcH7
jpWQQ0aa+pp6inDWoqr5PfTnOWBsWF4Ym8hStjQSPVyFiCcH++RJON43+Dm77Zc0
zzRGuN4a7B6qqXqLzu6THtraYt2hMMFPfV+gTTBpdARwFUf0jfnvVPzpen+bwLUg
OSz1OFHIYqUCZtGpu6xkWNf7YXE5opXMbPuQioM715g+8RWwLk++0qODr1VqM9Ll
ErUojT/EA4g/cDXrwto+FrdDlJZYT3xG72Jee7gHb6vNuHohqoykFW4TePh21FrW
XGGmrAyJZiihh5Sc2twVFWJQICupp+bOs0tDXmjY+13eb+diARwVgUzAZm/Bfb2h
ksxiPwSfvvbwmnkVjhcjasJhxixjbKM7xUHRLgUou9RXfX+paYmaf3m+PrktOkPT
MEg3jH6vuVUAh3sbXb7BK4Lo4vNNrB+2MtN5gLfbB6Uw9l1J1wOCsf6PNsb4fHsH
bC3WaHmzvcXvUEiSWxX/o+ZJ3C409eYqQzNquo0Xm00hDiWFUcfBkt6auZeAYlrY
OHJuTq3v8+nGWInS0QTZouT73TK3ZSdpTpI3FWwm0ZYL+g4dUv8KTb62yeGrunTP
vj1sqpOj6DEAm7BysKcgQS9IPI1j5YARKrU0z4JpQ5msVUuHfrgsuFTj+796NeVx
wY0HhygWbKpksRRk2KyShPSD1j9YrINS1gWsUqVKnuWFgOT6LWNiWk1RX7q6qr34
mXhrLuTsX5x2c0ojopy2zvL5qCNoUT0Luwp0ttHmaTKqYEbIStaPHym7CVZ7qoKf
5LVjZUTv6v087wjZkyqKJMq9ffFbgkZ9wbHB9t0SYXV8zCnn/XQxg0NgqnWVwEu0
XLwigNoiyxECOcD0zWGH5bbffdXc7hCjNbsHjPF3Jh8Yo0WCtd4knr+BJfspTB2V
kEcfCH+jX43g7F4XlvE+KkMMr2QHw0aLF5i48CaIFrgZkjoGu2IQyLjJepOj0C4a
567uVCQ1c6WnTZLn2Tc4JI4MGBcAuJVr1YOcM3aixpZ9MthT9xGOVUog6C9jYTs0
FYAfYADsqh6Fh7R9U83Ed+wAFPoDSJUz3lIz9SaFezaUQXNZ09ywCtSfoFI1il96
O/Mf9m2y3x5iSc+NFTQKpgEkUmyzzLlDZdsgsp/iTe1Kt2Z5v68DuGFbsF9woRco
W4Zds0woHugj1GBb5mhW6DkNIwNeSBM9Dv+1MNNxK4NdmWXend3Xs7+dGkteQ5nd
N7K7sM2XhPGnjm/sGuiWx2Czk7SlAUz0L5NLOLhsIZNOENVHx3hzWQnVhxb2IkSo
MbnXzRrXSy3+fx7MFATgYdZwg9A0+2Rc/QRT7IWmYZAvswkNkLVjF7qRznl11/iX
DtBWXD/DvP0K1HSCaJCneWiJuzyh4R0HG2aagPqoWe9zQ+Ke3RcpP14u963I4t3r
bAH9ofVcFhcjCW318pt7YpLmzUWRF4IlxNfYMxn+vouTOIGHORjGjKx2FsLSFkQi
9JyxvAfPHvxK7CslQqggv+wUWlO/dVdABvTjtYACWPSaYtTNJX1ik6fLG9lg4UcJ
LZop8nYjybUSHjJQHpS2N5isE9AuJkkNQRrJu2m7NylaWuyIUF4IkJWZJX71Yjah
JH+3L2GOkKBccyl82e+CoxvdbxhIl81c8jMTbZwgwQJTu1ihviZB1ZJWd4FlR0ra
GGHR6QvmuuXaT1ipChk9wjqrTefyY1oXJPY12gwLNpIbX58/TeoqzAWvralEpZTV
FbUGYaMRBFi4s5ci7T2/vjpfmiEVMCSuyTItAIaqyY4xQ5SQ1kqzu8i0vM5OBrF5
4LnwZgBsm/PXcDcnlXSVB5iYtWdVDEznjmI1U2JKuJGXlKKEU/YF7t96qUIY5WMK
2pjLYpPwigvN9FAc0EocpkXySYWq2JgnLNwNPmmTAFJ8SK5pZaa7f1Jkmp/LRG2S
wW0qOzf7JlCRKPbBy2NVcnFiX7L2XW/X9qqU186bSjmK2uztY7Sl6TJYicNX8KtB
knaKXCl7mbhGEL/W1VGGnzuWOa5LTTa4qhCr4gL2y0Fq/zH7f9VgfhZ9XUYD4YCq
VwNOQXcn9BbTOrU3ybH1Xs0+IfKOJDB7tkuJhT+tBhQRSNnu21NYf8eo2MBun5+4
aDIzKwmvFBVjcEnrihIWddqvvsUvg5ijCNyaamt7XJ0SqttTh3hTuDEfqFlIJF1c
Gf1NmbfnDioKYfwAi4HEGxF+RObER3E1oyz/PLVmd9ohU6R+9kUq8Umw9/Hx7kYi
0yZOE4YY3cCNmNrApIg35kBUeE/q5PPIFgi3YVRhcnlw+ZF2i1SMXrePjVz1mbV8
7dARqC/wKa4mxdXlgf2gsi7Bc7ypvb7hX4q3l2xCb2zrY9zxwwyrUe+m0AN7ZDQh
mShWPkccbhG0pJtsr/TL4pSD28heCbzvsISJ3Bp7MjdlVHvIjFoZ3G4nec+pT5j5
aJGgBRo2fza1rms2DsJQid4fFDB97abfmBGAQMVL83kY5oDh11WM6UG5KLef8IFu
HsRHDzeUsynEIOxiwwtxR/z6D3Jc7pDmTy/FKVCnblvpjpyo/1W6zVA8LGk1BcJN
2tT6ciPz1ze49awLZ/wV8v0YPj3Uj/HjlIQSWxpll8Ej3CJrzHaV/DHWS7kI9DAY
3PEmtIW4VN8nQViRYjTnxu3+0vJ77Yvh4vPhaLxzRk/b+a1EbNy8NOI9U6lf5myA
08jroa9AVF8JgXEqrt26O3sgkvQfJjRC4rhsvZVhd1aoI8RuWwR5pVYwEVdjwQXP
LNEx9iF95DKknUQplBNLgWEKkDDNaWZaU1s2pmpMUsuN0osgyiKt7h/JeQe7zlO6
RgopNZMXxyxct8r/Kzv1xJdi2C5jKXudY8CgM4MQLAHrVcijZ1v4Y2lbVyLRUCae
hzGC9KrKkoynAIuoxLkBUie0EM+B4ZsUP4ciIUZmu2EfcWieuCSdg49wFip7IMJo
MQrJnM3sPnPu39Mm6KMCH2bHBkDs+2RIXTRhxa0e7tV/9F+lMkVUaeknCW+U3emg
3tLgKOKz9AWTiPtHf3sgRByxpO6+ZKLDy399rYh3aXuCIM2MEpRBiiTHl073P5QT
B/Rr+lIb3LVIlrj/hk1QiAJqDvkzRG8fddOUyNzP+AoEE85zvXbUX6N8iOk6jJ73
y0ZBmtdBXzCDjsLZv5nNrOtdBmwJV41ERfX22rwesZKW0Zrb2xnoI2zZ1Jsmgyo4
m0n1XcXXW4uIVZARPnahBNxbHuuaWC3JJ9YKzFfMaZHfs9e+vfQootDy8KECnCSD
nM4wO3V2j/67mAJcz0r0PFvQBnHrIFJMUxCDzeTV1cTKIpaTilPajmCoWRwIHtBc
fFt+OptBNtpfSpbqE+bv6mOoEXzm/V6GbMpiJEiVMkcW7Htsp293H9BkUvkgF1MW
qmPVNfbVpPpywCQtX774j3sjGx6hwJVJBQKoNZ3+D5b3ro8yjwtobnfc8M/NyOLP
UXbRj3pbg2fIc5R2TkykM1IOYCu8+ATEnTF6i52XPUsz6AKH1hZj0wuDTlpA57hl
HIS6OWpxCV49KzOs/jbRpvHAkgYtffkc9L4zBvahsQFl1Dv8xm1W/qdGGqtgU7LF
B4YXRRrDrXDthYdA6cball+2TXNIU+SJw+G3i/mpjynDwCHkJB30blQ7hB6jvMgt
Ahihk8GaaVPd15LlUFPfFurE8/q2k3fjJx5Y4okXDVYaFAwhAW5ImWIgNp92loFr
vEVkn1oL+E+8Dy3qYJ9tDHo+4cKLW2TxbCn5RLKKgWUL4zURceN9wAc3LDdX+qfF
uG2mcylIhazHLxdwIhZisGSf421I0FmdXl7Ryd7O3HQhryZe0DAwrBFlGkZXuXAa
BnNoFVQsfzlOI2KAMzXsLoTucw0dpzLKc5mMvF2X4fxnZCYHUvqNwhJ94IrqBuUX
XHeLBFPdn/8Ta360tWNKZDL2XjEE3RAf0qV/jRzYoT0VmTiqgmPkbyeC8AIaAq2s
ETKwmuMDfNj4bdr7lTLwhHdlIPMKpRttaOCZJFfm5nPsW71qErR1Ni73ttgaovmm
WKO/JK5je3yS/b6n9BdHJ2nuBbRPaNV9enR8aqO/9WKhdcIQ6qBtShu31+iCgW7V
YGVUWhpfBfygjRNav1FuOeiqWNuVUugvFQJPZ7eoLtr4P6/Ascfij7X0V1Bp4rlP
QkHZn4eBzxkZcsU0Tvrhx8B9FxGfdcnF3EbGue6NDkXlB389CEQYTwUgiUVb3aOt
5sIGzSWJw57q5R3ynplbtBZwiD5NAiCTlijbxgq/OiMhpdIMMZGD1caAqKfzTPKP
9UqAmFhGtkmgHJivyMr2xV9F74bJjSpwVW8AqF1i/BixZvzVKDW1n7vKkvEv4Cj5
YspibfDD+pe4Lt6rfYw8NxgZ/haVamfaVE0+KaICKBzjjwE+nNpjKUAo1qHlwQu0
v77yxI3Xd8eMJnQXXg59MJLxgZTfDwze9i5P3PpAylBmtUBsIbLcbyHCGurfezhY
/iuzKKkPYSlJRjn5pNqI46B6ap8zaLRW7ss1nUic14iVplz/W7WnDNtwA9Mc/c0t
GVwXgHbFE4/eGu2aUdpKjsr7uwczapSnjT8AJVE04K+gJhPvCQ7CI1epqE1BCuaa
s0V919t8hWPuSCKEMOf0fDKtuJo83+UrQlB00cwpaB3fpgKErwaaBAaePqI2OI9N
JITu2joLuwAzuL/GGyxIabQSaBaEBQjNUwIPPYHD+a8c8vd+n9nb45l3DW/OdEB1
hs/MmtT73gMbcI/yKS6xqOZDuuNDDANYYLo81gtweCLxQuIkNclYZc0PE1n/esK6
A0kl5CcSdpRy/6Gc6ySxWi8OAl1gDKyUpRnnTtMg1egU25M+VNm8cc4/5gXTA5TH
PN25yMmwaDRvCTpDDgYjllN+6RxQZH+mLGl804SmUNCaJtgndWV6+Fof8snY2lRh
AKATcErAd+IhjxPoy5DH8BaRQMzuw9wUBMtCLQXUQzlJbO0s3jdcCJfo6yMG1+GR
uJgFTrR4dsD9DqkncljcDpsdApCZO+8gsbNnh2FU2czg+fYM9lAUxEDK9wk3nItT
AisQX1h7ioeSPYxsdERQvQPWjmo+xOpJTYZ+8enxo0ga1idmwCf54+ULQ7N8AA6e
GkK9S2ea/3HBT8vxJ8nqxGJHZWVEGRQ41z9OEsQWQN81WIQmM/dDFJzoUeS9WzNg
PXlHbA00LbLbcf8qgk6TpHq/TXVxMdJ0kPhoVifOAnmlujNW85yhhRRSlUfwQJm1
W55Dpx7s/0Df1rTrOwQxvqlH168MyYQxQhAkiTCZMDRw5JmYf0yJUXaThkCs6Nyk
fOOSoKAWxixEBDyDqiYnHyh/B9yxnL6WGUV1Xq7SQmGCZpuQCb9CCF/fqlFqNSU3
vmOxR7fWHCjI0wug58GuhkYus6t24sEFXqO08xBCD8BkMIKJeDCzqVbfsQ49HaWg
qPDvIg6UkNphlTW4TZYWgi+5kCWf+/TzO2NDZHUcxlJ1Hbt0F07HmTO/WZ5c0ttZ
kuinWMs3VnwKIG4FQJ/ttd1ekBb1h4FutxdhLsCSjEZWe5AfL0OZtVnFqQYnJy5H
Qplzw5BA7BUcQnvFFJ6N6S/nkUPy91OxMJeu/Qq+TdEvaJjhfWG8PHo/6QjT/MjQ
bhxlcqlP4waVsTLrZQsJxrQhwBcHTchpRcRZ4MiijrNYrM8dp9izzVBwT+DZhHi1
gsIiSuizU0WYDAM8A3QNHdOGL8o7Vg7U6cf/ZchfPXaDUxKzGs+44jMOcN+QiF84
hUmwCEeLI2DkyzGXVQ0FEmIBYe8wXtBF/RVPRyxpsql3wpmnrvQG76P7ARXuEBjW
RtfKC43hQKfPr9dYQUtU4KzcFLy4sIJoOtdlOjRTUWAUMZbFZjpp/xFIKtcNJUyA
rbWeF0/5fNMASgcIFNyxduEIYvBK/mtpHMmFuX3dqU2lHODr2TS7OylBfIbj3y+j
KnNRX2iQT0giQywtR4le6oDmnIUOdT43sHWJe5BjfXOzJZFABUKfupv1y0mOTNLK
gNcyIcfzwt6oVUo0MNgfpd5lW3vxypETiEM09CJOTWwbXeR8Y2Fas8MMqw3uE/KV
1PCyJkb47UScVmrp/IOf0wqDdp0rAfe7XtROCGFFa6uJf1TGwr4sIYiLlwaHEERZ
hJkYZy3UFUEI3R7hciefQy8kODZurmef+Ip9hgy6gzvepsaLrK3FicZalUCnfmrM
I6+KesRFKRBiIDLzwTyHvLBU1SmtW4YF84hvBbVhWNa/4jZMW+/q/PKoGsyl36WX
VoRYu7hqfPZhmxO4YeHn3Z5RVV0V+Aoqof7oOObfJO/mf8ci4baKO89wlOoHkRHO
lPzPBoF8gqBuEWu/8ruWfBDgCQjxjE1vJQDupyY08BSRWWVE+Z66HfE4QXkSezVQ
kvk2tzPtlUsk4LNgSYGVS5Lpltyjo5XnMac+26e1AwFOXaD86kp8TcezUDLwfAQh
XcgbchUwHqmAOic0XQ8wqo2Rloi/zXf9kFlTcVrex5R7dZmeHaiGwAMkPo0GKTcB
BS6PF2b/R2paLvsFZh7tGl7teViP0Vee29GjxmWcs/PVzw//jrDtkBmrJAbMXP+k
HFE5cdyvfq5Hsx/MKiZGke7dmNcDvnsaI1HMMgLjmntVEM/gNqxiwA0hUv1GDCZV
dse5TtP0HXiYIYtUS2pwITUd6tNhsDRkHb4Ewi9J+mvx3t/bHAwS+KpuN4LhLvtf
ZMJ9y9HsjtLLTWljaTVOQ+fuR/HXX2Tl6GrPf5XC/fEwnzyOtAA/E6wMMuohfxl5
1Thn/jA5R020T1aKOiymOt+WggEes2ffXKeKGYDRBo2KnHgLHOujXQhH4nMWfmRI
LmFw84xd8wKkHwpWejVNl2LykqpGPT8tU6r85sW/JqGXOwBqJVsa71dTgyHnEgd2
SJ5453QIgrl2UFkRbLJQyc77MC4j/OVY/1cH6QK1kmulgFhWziGBNebF+9H2u5a1
qezy+/XYe4ycHw15jC5/8kqyNsgjmoTIhrdoH518gtFk8il/zZEotpIrxOr1cBJO
VDhTz123G+gyQbOSuQXiqn3w/kEndxV/1roiMOtGuEeHHCFSNTj11adDsD9UEgkP
XFGggGiJPYpx4gQFl2WnacEFq8B7U/b5wvn9hoOiOMVFixGKu3c6qK85MPK0zSvO
ByrTgNdzV8L3bXnKlFxjn+jC1mYcISQBlHdD4aJ7x1otDSd9S4A31DuiNW5+bR9/
1ejONrye9LORGZ21ygcP0GrmtiCcG7T/dA907uetIUGgCAMpv0juTnD9Arfk5ZV3
uN8R+9O6bBmw8VzA5UhV1nTjo254lk8k7NIqjRaxG7brM1FRIKMP9JBvADNvwZXA
WbYu6c6Fk6ZdMSa1AzFK09WYziGgFH5atKFrtFP0OBu6RbAzJULLj7x21VxK6ik1
rCqnlzyMMunxRJpSMQ0HzO+jMsQ5OlVRgbnlJZlni4i2JuCQ46v1zVfJtXVK6yKE
s7TEupt9vSSn1RcIsl/oYbPcdARP0YQBuCmGu41amlzDKAwH+pcrfyoPumGNM9rG
jzf7UoR9H+NK8gQ/DHk9iY34knt6aeV3dbFVQCiA45m0jrHtdZh6Puoz7cBX/5sA
kcqYkMeKCnn7GUL2lvxXFI/xO5Aa6PZIcJnV58KWZiozvHsTuv9pXK2vfaqQP7S6
LdOZ8m4poqh4gsip58he3aYVZQtHQuDn7U93X4+yxcOxjCpDx6IPWPnDiA4o/LtJ
8h2WOFeYZfp9TWdhA2aSsgcjnaq/BBAYiZZUOAePav/+0Rwl7DcSCoFU/UNYCwXi
2Sva1Av81VOZNe41+q3ZwIbQaGFEdyeRyebDxb7b28i2igG93254jHTCeJcSVBiy
2UREz+h+jZG1zDmhawNkT8KDSSZ/uIOoqq11LX+6Y+mrPtCHHGuKpRDdzKYuANZz
rxS82/lPVNQM/D4FJWKv3b7xImSpKg7Rg1Cmz+dHehJYkbsx0ItB/l+GaWAAWrMN
UzT/YYxW+aXE5aF02ViKtrx9Lf1fNq0g1folrIEKIusxWzZgrA2OE26pgKPbbLi4
QYFx1hK+jRyxBtXsh9Su7t+Sqe+J141g5sBFnfQ7oeZu8Bx4PYwQ51wXezjfBFqe
XJCH4l1pwhY9C1/0y+1eJu9cEyizRYRonfcgBKytIB9s+pxfuLYCycEwr9A/GtiA
3wk1ZdDZSYgGgARWMuq68idSgrT57/KAdtv/CYt1AkoElsFPN8hC1j9q6SbrEOPF
IG0t/VZULJQQm20DilvZ0++gA0LuvF2eIXzOqJgrMs0tY5xi6VvdDEs1DYZEwgLW
CAOBVwkdPTY77Zrzmfus3mixjGZO7+CNOcmTKnsUx5aiIXR/skehlHPPy/uV4F3i
exuwLtcOktdz/omad8xKcPLjCkUJ2kcENIfCtyTXvVSECJe45sSHhCYH2uBKt6d2
Qf9c8HRsONEgrlID3CY0z4RDPUeVFJRzBCyvkd2hSqPCiTXqe/tWBpYrTw2YWhrh
StBVXN9g8Sw3pRyUMfzBhMCxR9jZ7blL1J6Xpto1pAfnkxTez6YJhCaw8kRSWSH2
i6xEOohnjYibe4q4H9d6oVt/Bi/BAofMrNYJsN9Xum6DFnGTJxjTVMqZZviiEP77
07adVzMJebvhNJvyWmY99YuC+DRM3h4+nk6r9GfUdnrztUZwyxKVsZ2iBX74ZCcN
7gpU4Tin6iH/YhMkMZQN38XzFcY9scuAo4xrXiVm6wFRg18lcs8m6tSaZzrx36RK
FyYB5eDQ6/wxlpfG7X9q82YzC94d+cQD52YtDLCiN22MwKN3mqDWTCc9uEhX568i
30/jZkVCKYP9d5Y3WHMJf1d6om+7oyoe17KwZr/MInGjGeKIaBRTcScnw28Zutp3
4/WDdK31oFOLQhrncBYl621pFT3qzPRYFET/kZsgsRBKVLztQ+8oqLyQ1FOQZEVl
Ny7PpntvLzOZ3p2xj0Bbnv3v5TrK3PWYeYLG0P0u163n2+NmDSxA7xFvCPoOdHl+
SUnchTlc32FH5qUM8A3e+TOFMGLAVg+snidHERnaJXP+xD+5dzsh/O7bZtdjnBt7
CNHkTqrfQWa3qKMx2sgNc8dLDVNSXZzDz67jvvJyNB07PhyThA5lbTtovhkZGvTT
Z/7ODLX/fH0VRT/60shc3KZshlL6HNuZpU03U84lYg4YBF9iAScwsuElZCHygstZ
3U4hUWm5hGpxPEAbhzs/4Bmy8lcUc2QVOBD5Mj+nfEFWlO0+ktXDljsx6EYrQYy7
vupFQ06LSQwOdFPfmhpbopQAZhVxVIjX71JtCDPfwM1E7uy3hc0AycDryqdQR+yT
fB2PTSELreLtSLYXY1pgCLF/Z/ja/vIolOJn2iY7uJO6E86K/oD92naRQEJgqZJt
qmo0aRJrI5cV+ma8jZq4sgmJPemUJNj3+n+ZatRCHZzXiSTvGbgVOm/i/fOE0UkI
41H/1Qo0Jb/z6CbMHMBGfXWYC6CHd8u2HmoLlBbTu47Dhx1tCxCbIy0DOgesl0aU
5EuPnUZ4z1xVVpgmNpXwBzd/UI5jsvcniMpimO8ZoULqbwwECiXR8r7O1L1n3MUK
Y+jqd+O1puOBSTYD+1eCOgPNixQE7zvfIhFj4Z/jhbwmmB0e+wMKqiniGL8P1TDc
Q6J9kPumbukkQOV73dUDOu+a7VDT48uTJQDnlGSktmC+dmJu1Um/iMBgLgS8kUj1
TmFf3HqnObJPDhQSJSHvAmy0fGFcPX7H3iOm4B+N5J34kBTR2+DRQKb0fyVgdPse
x9MpW7Mtu5rYYGhyB/3I+igAdQPPIsDfaTFM5HTl/sTcaxygXYS2ihdtnKa8XwhU
aVuST69rWsQKUEbhkTYpUS2DRiQIU9dMFqvJgWBp4RD2G7W+PAkid1sbg8LIFfKX
xSNzinzXletubekTDai0XeW/y5dJ4vTolR1D0tdkfckrq0TtOyXoRKITZQTDVMSt
68POeIpRKnp4yFU5KmCwzf64rwtwJBikGx6rVK0EKYZoO34MtF8ObzQryQ3ByGla
fCA5ZRcv49PKmqHWWghOLLdMqovR+7y66RVGTQTTqu+11CzuYALLPBhQXy7oIL3l
SUk/3RV+Al/ycYvBPLiJitRMt5z2AR8xw3wpfidqI+tJWfGB21x27MoKC6zZFsCg
YrhcfHZbryKnJDYzx9fl7IXdPH/wSTBLkj1Wz3uOLnUPYFu2tfH62VCaxGZpJjGN
li0PWVRA/2gVdB0lUNlrOvzHxw0f6hL/i1y1jEsdVRpPNS9bZN9A98qsHpocXdvS
uz4s9OPtaSLBDa6HMMibfZzKXLGYVBqxpLXpH8/WEtuZAgo3frjciWUdUBMFvScb
tH1/z4LxP2oFuWaSc/0geLahATkybe2ePtzlGz+oPPZiwvWJrQoT5lQ+unTqAHo3
SccSIMcitcxSTqVzhW9B5ueVdFAWRWig29bBCDuPftr/GYMGlZNnb16mwt8iWD73
jCLd4EUFW7Ikl7615pnHY+SrI2QHTXCP0xhB9SzV0dRoYC2AL2G0i57AZnK7HX/R
JLrYP3mGjAimTFWSJs4qbMJsRLTvY9PCA9sPuYnmvLejDeJECM26WYgUbbXWtReo
L11yfnnTdkdxwEkQBrUJmg55WDhIj07mSrSiTC037WfbThZu0t+ocZGJht9ms7IA
UYyN+vtbyOgXeDw/SVTvqCL4ZQ569fQNzcwqjPCJcLkZGgXVZojSK6lCEyhwRD1N
QXd1W5NC3pP/eACBGFZiyvPI1OdnKAEcHj0Ub8mP2g1N18EMu+B/Jjsnqd6DA04G
6xegztxrGjCqcewQLFbBVwCOpnVcYUGqOIs+9b1W+Pec5fNv1tqEwhI7K7w8ejRD
1mHh/lSZOjcWrhcfGWl0e+YHvuvzewhiDF/dZo/dBgJQ3cZPaaPNBqcHACcQsmnR
yqahAjZ120xUTyIPjNCF+stC80tamfOM62d0qEvEM4AVwz81GGd+LxtKl5obN4Id
txEn7BTIn5UdiQZPEfx28dC22/xwvx5W1ACg61Fz000LDVRhs+uE1tLEwTY4lprV
uVxKdDwBwyo0977o2vdfJGW8tAuggraPiGwUW1auX9OvNaHh+Ryp34ydWFH9EzBv
wZr7/3ZETI46tSMRUuPHVQDQrF0WfM54WDIRX91/hDLcG/4hazm3e7mLh4YHN8nx
9qfRSDGeAp7I/mVynAo1/M90LNO8gfzgJn3mX/1YHUIeZg9uA1YuMFwzJXbabD4P
GtcFQaF2zxWBk2KFwjKrf8bgPEpb/nP9KdUIhZWuEoEZuMoSeghBArgXWlLqy4ly
bw3O9H3D2Jl83kvuYjNeKaVmtitc/up3mo43tn7j6BWjqUgvwAK51dF2nLm2xh+x
m1Cq/dP192z+r4+hdL+A0t1dqAKIaxsR/hawpTUYF56+N40f1NlIiQUSdHloeD88
Kc6k7wE3TNN3KSUaEfm54oHUHZVsTUBMPAZhsf+P+jY2oHTN7HvjnQS7R5viqVIb
NU9CZTEYKZySxFxiyZPxLVo02HUdbqAmCVzysDOzTHAdBAH//2T02gSaalmonqDg
Wn8NFDa9DXPz9MSvvjNxmj/INPQMKJzhVd/FPp8xIpe3TZtYGweuQH3PMcswkPbV
KcZuDM3zHhLSiomS3B7x7jEBEKkDBcGYbdumXdWt3DDFCNI29Pj3tw4Obfvqv+6A
W/gtueXf3jON0Jd9VzBPoUzmtxiw1cw43pPuIusX8tSn5qUGMP9RtL9J6L0Ea+Cj
uKPphL6VEfX6n8AqiEYA5DLee6ua5zEuM9DCck/e1t0I5VqtrShh2gkBVGxkWMx1
kGycQYPKllPGLURqLHneNayXmQAQOL5TzE8zbTy0x7IWlh+T7QpyvzCBWva2UiBE
7VXneLttdNnC4mruk+a03ydJuVA+zWbv+Q675ICldSIGH47ge75R/oM1KNswZk+b
YXGtTnH8yto+ngYQvTZUxv7YgRYOSNDzeUh/lt3XreIrkNqrFjOhcekC/8H/+sgB
fUd60MGzj+AkUtoNTYuzioHGODypugW9yqcp7G9Pluj+iKDZldLefnfOdWxeG/9y
My0ErWBYXVP3RuWbewIIf2Rmg2hpdqJOfYM5ys4y7bBl0DZ+4woUxUD6OLmgfqUC
WtXacB+/ZwxkLA36V7bkc8jTb9TeG7F7+eFw5G6BSRrOHMyDOe57+xjga2Yl2ndZ
tcY1Vb4pT3UAG+2zXyrvC+cvhTQIxJ+OPPhaFbRWV/v3N9RdOCeOyNlsT9XcbfYn
DngLTIPv8n9jluv9BelEJLB29EzDG04So3qckEZFGBlUd3cHSTxhVbsPi+NhsyVH
TaW1vPipvPAntH51jkiwVzbJGZkHXPrfCD20hKsudfDtFzQVzrRZA5h5VasbJWXm
w+R2+PTv03ejIzAUmiig2VN2+mAopWdyU120i1J8z6LmYAjP6vh6u5bHXbXgt3Mb
jHLLZ7AoH8WmafZUBC7QlIs2gQWPw3B3bihgAP4ye7pUnA+GNMTVWhF2L+x6bXav
MELLlmEzoxHSt9oqrDvoJCGE52P68IlLmuH9MD1U5SxrWcyrgD1BbTJxzl8vDtfH
Gz/Z3c9xSfFyXa0ckhUkau7ktjqz6nNQP9KKj7Dv9zNH8uTPLVaFCL0wMs0BQaAQ
mOHXKHQr/3uaBp3pyjURBkSp4DkQVfBXahWzOqL6o6hfAHrFxyFqmVmkT8wNocMy
3cGCExvW8S2mQmcKu/gnmNmwJ3lE4upFm2aGMYMidbpgwu3Wfa9DI62cCLIVzx+F
9GcohLW7ZdMOsulS2UKHhn+eZ6x9s0+cmk811K1K+LGSzF+iV4pIeyr7zxNY+os8
jQLs0zw4pZKhFN7wUgdrWvgYq5jRoZ2X7HtVejBAkZWyDSmuUJmZ1y9+0Xhyd9g8
FZDNYMUlHpBs5Py2EzlNrjqIZpm8sTpio2EsR5+ldn61iQhQwbiAkka0XSJgyR94
urANUcygTlj58/b5prNc3L2cLCAGt3VGRZ95mWogxQCmRVl4Cb+B7REQaPGijdwK
bBP20dCDQXGOELfGi1FR6QQN9ecHCTvN/Ngs5pnlURPQugAF8PA6ixm4a9pqEsKQ
77R/QTpah7378zYxsi/X5Pah2fDfHtqGC/0AqWFv6uyPvfxvrPaxQhAwvEVIpA6L
wlKWfwPSbDGv5ziqdDrjhEh4pDLVNkV6U8YeWkwyupeFGuFSfrYQaIu996FNdpBp
uwSAXsJn/3djrVKyPB25wJQ8rBilUDLVhpwitCvFQfPBES0ZtsdaTA33xngIqjCL
bna9Fgmay7O2LqCiOKSff2Gs1TefUe558ULSNBHurjjdz9cuOeWDVUi17uWiTw4o
x/SpUwMbkMd5lR26Tw+L4BM6CBNuVqdHtVoqMp6BzOlfG+NuQSAOnnK6IjSfiwk6
KXmr5gNtNnB8zgaDDtuuZLtYbKMarm6fNIzywiRZYKHYIdlGoovCpF18jbTjS1Bv
jgrT0+2CbXUJ47RHJb5lCRZOc3DPwYLbtdv7Ab1E1KSOET598yN9pRK+c+CQb2cA
rVDgf/IMUfqCKhM/iZ/N4enFQoSsN1YDweccg4BJ8Efg85ApLZtpSMnJohuhacWk
iwZD9GQ3m2WTX0g79zAL2wm9wXFHgp/p4GYqoQJn2XYju2Pnv5HF2+aZ9p1P8vXj
f9JnKkLzJxIcxKo+RnvStUX/HgHXWyJIH4+RbKOuIU1flHnNKyEPEinEL7WeCG7q
j/vE7LMDar5WBSAwbPQMK6SipBoNneRKH6TqGl7dN8PdDEwLFC3vl6M0KN5pCRDx
H1UAb3jpCZiGGH/+eQEAyhp7cvt+XBEjX8buygpwZfV0wXA/jrneNUhHcy5eeo10
ntlMH42ywnPb670EjZVJq/uqLmN+SifXdUBATZu9ZkkLHxa6sm2efZR5nZGzsa6E
L9oVXi/0GyaZDWI+aPLrCboO8yDdvIUw5k7sBiD8kWkhRs7UXvIcOlbsjFJqD/SA
7ObkL5yLG2XASX4CFj3M79wZL7D2aN4pqIy39opwdEcsko3OFdkJaQt2BjJXLACN
g6APrX+HbenXebcVWo8Pa4qrDWGLa7wwNgmCmLqCLjP4re1Rz1DlxPL8fB7LgXqQ
FdDa00nyD8kt8pW8vQa/9xNYIgYTt7oxcizV3z5pPcnVwiX4DRmIr7y0aZafxtK+
F3ZBFzqjl9iEoq5OEPgvT+goYIGgHmYCNV5GwS8NJKWvhkeBL8Aoo5islYkzrtVV
lvj1bwPuL8ofHfkBpMes3iQXkedikw3ynSsvyzA7Gzi/JiZZEYsNFeUMCQm++IN6
Lxc0TmiEH5uWxHvW7Dythbo/zVVG2F5x35K12LXwHCUZ6MT/jOkDRW9IKdIgz1On
r77iQv5bXHJqeHs25bUaaHYT1bzAv/ttZSfGn54qbA6PSnLB6utImfIeqozRHNlx
vUjddc107su+8NpT0RM8qEBjbA00x/GK6yxMwHXuQgIjr7XvXYgKJOptk+ivADs+
dcvis7N9JPJTJQJNtvUSM+/HtxwwFyihrQfkQ2V6yS5YyEQodkhoV/SUBikr06OP
1OZTuStqF1yfaFuTa8HrIRWlT2a0xg11cqgySuDqasBKnyi+vVOU5zvs2ee7IZIf
0dWRgfCoGE7Y1GJPDhqR4UdAQ4FsrgJfKzfEbjyItZof5qfQYXcsMXZ2kALKrkfY
BvxiTe6a3tMRFhnXZ0+3/7LytiuJsAmlJc1pHq5RLVNRDzYARxpHqwTrPSV/u5cG
97DvhbkczK5GD1m0Re/z5mSUoVUwekmyW28F+ipDmnyO+scsluVgPeOhgzFZcGJu
OnORSL1Q7DG2beOG76rI0ixGTA4oaXGzJ/jZaQPBGC215Bh9fop1vvTLAtlOelcj
Ly18TES95xk9pUB5ozD0HFBOt+oN8fQ2yBdS+tMW+1JUi2BZA1DyB2KfhqTu6reS
NaSSBYtdU0yQTg8DXgYNk9n7Okk4SJ3Vhj9QsRGAm3os+fOykit+YKcAKGfDnjWP
xeM7hieeJC4A8Ot5F4kFsrexHhU5dNg0S4Oir6mmJMfSu4JnCTbX8cGnay3X/uR2
wBe/Ve8BUJowixuJ8DkpaAl0rQ1V3uXj09Vpowtyg0flb8zhl4qfMAHCA1dkh+Yz
gSuiZdVBAveZxOCcN4wuSgYg4KRR8bIKDCgSAAlrwnS/BvD8xwP6FGzbGwvxXV/i
uzu6Y6PiHOpwhJdrOcQEqA/0KpddKbe3mFobqczj0SZAQb2xmb6vVuvdBx8UQIt5
fFoAMKTwtIkdBlQy3klIXhy3TWU8rwJTcvAio8in4zmtD+uL/Ic+dVGKCqT9HDSM
mODq2pzw8nCkIYh4K25NzDFqfET/efFMOS6J5jGh5Z6FgiQZvHffSazsVc2lBEvf
cyM3bPXKG32m0pjpF4TQolBgc8M8jErgeBz+bVXUkSVrMeUnTRteBLzZkfPx9NBy
t+LsFhYcRPzS77qtJdRVAOIPZh/7eApwrn7pPRVoCzHFI50oCYe9IMVAPL3gMMR/
RDasRlV6CjwYgDM8JfFFUKUol/Yt1r+pJTtN6BSg9aNoqMuAkeMwZn3ZbWiqdy+S
QannTdHjCArlJ6YV2xB6Qd21Tyl1UfnopD85psvVXgkWr1rZfDvPRcDAb5sLFMjo
9Q4LemohvCEdyb6PN5J+U2FlVF+0BfFlgHOI7JhlM0IhwyMAxlb0APU17UbFuJHf
+6iTJBBwaY19G2yL8qaOhh5H/Q6UjJ1zyGSDvcDR6LIn9qmkTcitx+n5+QWYfxnI
I6EPsDxxR7NyGyAA1QLlWgaMG8gSl2HOdyCbwg68KB9u4VamhwGKYVfyQccRB3Yb
7eAKZZn9iH38QlcsgsXnoeQ6Na5n+iK8rrCAXgypSY5UG7aBpFbJN+vSfqdzBKAx
iXwLg7i36L50CE3Vgpq/njoOGkUsgGcJf1JbG230+HPXHTi39fBA1O/VwgQTOR7R
h7+BC+dYCvIC1Tx6wKMOAAY6PTD6JMzy8LZQeMu5zi+G7BAfPWOhFQ1UHoK/4EzB
t0mjyZ9BXLH98Fnzu9oH9/61yiwbsLe6lYlZTkWdHbJbNTzK1L6diJV77DPD+9fy
4TEWWYmFuFZcebFwEJvZw+epOnHwjxIjcM2pT453VPcdP7CuJHL2WJQoXj+l+Ni0
G6xS0NPgYsdQoOe8HvpN84Q8nhjqSrQFW+Ng9gAewLrAYaKIZo1LDHcY427vtk3O
xi9AiSOv7ySOfQaDuQq3ZA+Fas1JaQH0mkTXFYdzUH57TwosmwxZni+FUJB2ObZP
fzHOa4SXhCitP2c4/cU1T01+gINigN5+NzxjrD+fsH6Haj3iNdZCjJvxL8fOm/0k
ADvAPQlt0DZAHK606mHQlDw5X/16/cPEo5GLei13IqYbZZ4pS/2rBEv5tgclHCNq
JkXECGoX0/+bQbbZ1na2dxTnlMQZIKj1MBuh9MIedzF1bxTASe+DW0Gb5S267ZdA
BhQwOAnEmxAAmHXM2TK+p9Y9hFqwWX4j1wimYTy7+MPtShjleQlF+j9x9M6pesbA
HuoSw2xMrHP9G/sjYC+sZE7py3xWtCvfoYZ2uy+AE2QEVuk2q7SQlFPKGH74zefE
eD/PXJifY9qXlHgL7rOZH0HJc8gHSSzYmjqDeEjDfeR+mi7E8n0WXBtNiHC3melQ
Sg/7Z8O63iTuyKMqbCZqVbjT0A3KYgDhIgYnAcmqZlXXpnreFgesvaQd+GtIrJGu
Ejl1VAJzqxg+m39RhFfl1sajpZpZHbA5U2jRCDv/qumsTx30BLN4PnBEYK46H4Zl
sXHS0SrLifjNCzOFUmVLNcehfXvooTEDQhJeltJZTAGFQVre68PbCRCitZj5PmL4
UPbzmrf5BzN8bhQO+cLx/zHaxeYiEHD3eEmebsnxFMt70OIcdHKAb3jHndhyexZm
1iFVGMNzObYF8VMdxO2xfagRh8koVFaquiCpLnYPboOAO+gGrF4HORptMqWcnBfV
ni9VNv+ZO/oXAEXBWpmNAHF08CGHJFJSLolwwNAq9lLMRWANAfSv7OxDjv8qcqHs
ZZwMViBXnZ6tD6VgTdH3rQ0TQVN9zY4gTt24swDMRmX60087bot1KD2kp0kUiEle
lgMo2lOfm09gTeYRWmDKj0wk891iljQdpuxQPDd7IUYA/q+1wQBCiu84utAGiSPo
vf07S+aRQSKlYjVG9WvLxUYgTILQATiM+jj3ZnqGekMsD/WkQ7iKX44UbhfmCbEf
Lotptxy8ij/aC3/UKcFQ/06GlEWp6mq84m82QK+SVriDnpPlcJ09E8vxd/GjlUGl
oZnh1x31afs6TCi02UKzy/9aOiOQolhr4C2FPb0mHQHE2FJJU5sZoMVqtIVwpxHK
faCcJZ4V/AmhFqpEMcLR4bQCoXrx2pGTaZ2mhQybS2fwa4L8caaJelsQ0aWOkhI8
VcDOHfS0EotQC8OIuxQ1zvNLxXrNZ5BTBTgmQT2JWFybbFtYMu2VhPR57mXVSagw
2YRtlHirhs5HnCEgDDq1p/JJnZixTOeP/xvWEaHmg8a1JbJ1mp+kVhank987U1rg
L0wuARLFjqoKOM7MZe2BTRjfeCJcQtTR2MBtEUtbP0/iSUm3KTQgCeE1bVlYEwUK
Y4CIC2wWsdpjbKui+b9Dg7G3uHGfZIAZlPAtSuzh96kS9adncpfJSG3e7kmrwrOk
ScVg5lBeQrx9ppDs2M1x5sk1oCIllfYp0sRTNEeRnFxFvYo1q4YhbonQCdx94C0P
NxBxY1Nr5eVHsTBwixkGVEQjlhqS5hH+SFE38/TsMTVtLEtZt5pt8TOCu0YgPtUC
eRdLo1iZLM60EHR1Z3LHtHLnwu7Cuk6LzdLd4sIX8OA3YQ0e4fRqqH6H2BRJA85i
XWp1OTUYg1uDOsq6ZVFtvTjqXY4CiFNqpse+kFeGAR6SPkgXz+JhOSPzg7GlDJMe
Re1YkwLq4CXCX92tiSeQszrOR0k03V/n1owEZpYtW/CWjopwRhqY+buiN/6GYzlz
MYywAp1iVZUH8CxICguxb+eey67moT7EypOrbbUFeO0C/p3e7fM0j/pY4CJ8gsux
VpfdlptAsFrEq1DzM0LyMsWATB2lWey5LwB8IWynGRYBnV+4wNLNedc8XOTqEA1H
zXwmIzcU1rmRaEycgKfKP1asNaLvErqYJCgJhHQf3cos5oR1qDJYedU0wvKzNlTW
62IE0GXcsBXXE5TXGQnZWCqbK/hjbqK92ZGB9TBY3V61HtERyHWssb8R7MlonaES
ccsBbhNtuzxyDI5hzQEL8Md5CRyk7BNkUigU8mawsbVQySKwrQxdwj505bDEGIEf
+9+kyIJ+CMtGT2OHgchECKwoSG7e7dVrSo5rbtYsDtIYH/J45KJ28NGZ4SonLE9u
Vgj6gchlw8bg0Dn9mD2hxO+IEJODeAAN2PGR6HkE8vu1CzE/naiC219rRBqS+7gt
BjQ1BnWz3jUhFhP8zS/2FtbHLVr/gcIniLs13vuA761PPehu2mTC96lrzylSSc1g
znFE5eMXZs9eUrv8OnRRjqR6R7AsjubDbonpX+jv9hnyUVLqdeFaeeBrv+tCfjG0
ysK0BqIEZYlMrb4BK+2UylRWpK9P96BFiffc5VtvyHu0e4pNFEf14zjOY46kVY2B
u9tvT3ZZtKekQaKcN9YVYTb7gv+1QSgf7my3hVVRiD750znI6b0/A0pzXvY53eTN
WslWgZHz0TBgCTka0is+d54rFaVxeRmoGX0cZNkIffB0uW/9T09JL0eTxho46guK
M8FjrUdJFrgRaHQJgyZcGEHguCEesyMIZABSJktXmuwYo8SV0RUPkcLtNwvhn9ux
gkQbsY9hX6xOEcShoI9vxiW+/3sK2SNRCfhiTHZRNYPhNgg8CMn6vBwrTD6YQ+mv
z1M3S38dox+e2cX5+Y3d9pf+oDXD9Atpl4K8mll09d8RSCDOUAwP9lxpyPr6DIb8
7+gQolP07qTtWzI0kCIB2rV9BY6mrNs7WwbJf6FKzBUCH2n9zZHTfeX0kaiY/rmb
j2cDEAvxE0xY0BRGDzcKGpYCc0/RDzRcrY7Du9qo1PQ7+oNTnGG7hC5wHWIIwmZs
N1VuJKTqpE201QjvoCUdpFQpy5u+WRuK8VtnVMgzSCRo1iuiNvE4zmDvSSkhoyJs
EZlKDd7inzVe0+9OcrZgK/XYQuooFr007jWYVpHWaNzyTjF5JSRznx/bT7I0f12T
VA/9tlJ2mRXCFOKv04+opi9t+c0NUQW4Nq+WLDgOgVirAvDFDoyPruaE8fzVQ5AB
vORl+cHBQgAkTZLWxd0fNUm6fGiho3WwVBtyAYu1qgbIkrXOVWuQ/ojaVorIZt0h
afBFZTNm94KaM+1XYpo9eca0yArNfCHFvGdc3dNYahOhsrMeF8FoBVildEl9vrG2
EEufM1a+HubJ+1qCELyHHO3kRMF4gfb0fRXnKj5F0JxRI66NeBG1wUp9sfRvhoDw
8TdGrVoZ8Ox8mDtexDf6mn9pSaGZcSugTrWp84w7t+BjRkaMbM2Xg1womTuWT+hs
VI2U4UKR0w+C4XmTvDl2/oEwhhyjNMcauN3QHG9Zc35AzFzZ2VQNQz/4UeuhYgrI
1eljLW7HiR8doaw7UXMSvIVVsZTuuviJBoZGMhCY5FOL10LN+hQB1O/FnfIr5ALk
fmrVbt834l3QyWhHmhc+YqS15rKnPX47AHpLYBjhL2rPqw3KNRHMNdShnqoIZMP+
D98izWLLupF/ocT2D49OweXb9xIUVjB8jhgjcaip/QL4pwSl5bv05pZsMcc5eEsk
Q1iHUdiHrOoUSgUUNyl5bSB3eJ5qecMdY9fySqC1RUa44BDsRZAFVxj4+YehWsmL
K7767aUlgBHXZ9CRFGSlOaII/otDQptz69mFmplDVOp7YInxP+uiSxnxpMOUhFUP
MZQ3IHCKAQBY7vJUdd6KqXb87Qo2K+yis6QTkW9HLlFX1vpl3wFOjPjRYoQoH9HH
0l5+NDUobgw4ZyTkGGsz6ZNRE+wG6Y6UbdwrVikrU6AxOuFihc2Z3Ge61keAWP33
tE6rCdgohK7B0BZO3Qt54DoWSqz/UPuOI6vySx3YgaC/GNjn72Uzq/ROoHpUUBsy
arSKBD9Vpq3khyEGrqXHrmdVVm5pIba98WradfE+wo4G5t8D3ggxuu5sw2KjF9u7
LhVF377zFogoP8/WMf6ovcxo3LWnwH8xpUNDokwOFzvnAvU2ut9r/pWShyqCjYAa
PvhVASBsrmQU8gNUufoP//0TVdDNhEkpR26Er1u80AaC/LREpQhfzpQbsIG1f8Il
/983p3Pq6MqagNMmKODGnD8Gtv8HuUc8hHg6NF1OvUL+7AAdhUSbXtBsJL24Fv5o
jMmXkZE/DdJRmGhcTjTQ80e8dnu7/B5/pPPPOzb+xUaPswUlBnutVfi7WgRrnm8j
9xzRMOCTftq1VQiyMQaM3F8AtUaNfewEG1itTD1yu9qdJTLfZAJK70X9nj8GS3zv
Dti7r7IOETwh0pe4uPpZBXGZdWY4e6c9WZMkASjYYYskN8emvS5p7jTMvRbNis2r
lMWyXqKkIOmbsLDqBWPnl1CboT8oHTaZoL+SScOTCx3mA4UbS+pqu4+HrClDBjFA
prCLqTOfEa0/DLwuPTW/fob9R6MkAsoBsKq+mjOwocjSMBhlEMQFKLhCS7NhjLVU
XI/zB7k3Sa9DhlrCgijbCWGll2ayMiRZJ0PhUMfVmmRqezp+6zB7eh2JOsvdVzij
UO3HjGZ9IyfE6eqicuSCTuit2reVQ525B+aDbzqPKZya+b7U01jkrV0tPxSNY2Lr
mR4KDkHA4Z/DF50FC0PPlvZAzByIeUeAQ4s7cVYoDa0JzPurfW+O8b1cFDyk8Ovx
L4szCU03n/q1Jk/pknY6+AiGun++xU+AI03J400/telZf61kdJEytl25mv/elcG+
622Jhl4wApd53oO8WZVn0SNwSuN5aEj4NUYLnqWcSNR1aYvidcpPNwbFe/12jpsR
dUnN7uc6BJhyfsVeS2PKUS03e/Ibf26gmQBQVHzIoRVAOXpWZB6pOeZJgEvx+RQU
kipwstTVOTFETc62W8ET8gZkysUWYplp+nTKfRUEuogr/Vg2W4a8u2qx6+wJ+Nvw
aXcSWsz6TCSnWamFRroKIUvwEbiqsPVia+EZZKKylLmfTxx7Yn96VXQWqmQusJkR
GYG+kZe9ysBHIzpReaQ7WWTNvjgC4200rRaZ1F3U326ag/tutocpwCLLKYA+PGKI
xl6OloMujBOTW+gDlgd5NCe10BXkhS/TiyKjABAkX9CAY13gnThAdd3wC7JCUvAy
GeF9eXk4L1PvuMqtVZ6cjSvhtGRxvg30+Iu8+oblYC33WgvC7VD5fe8UMn2FufDr
l5Va/gT6qfqibSkxRojPlhpEm9ONR9ZkCFV4E717rHiznM3EJOBjjKvZQRq8h1/b
xxxkfJe5UDhqd6clWvDUaTgut8vtPSAZjJH/9tru3FFk/aQvfslMtbTXsuF4HabT
ZaEq/P6QoQlriK+9mIBoyUi0sJnN0ukeYxy5dTQc1vEqYBj9kLnMjGyiRwq5sBJQ
uYtoFFJ3gKpIwosjbF+sXZZwSrRSVp2+GDSOzHFkEMJrsn7edZNNqw6GCOaXvV5I
AuZF9iVmmSVi0oWcYQlYs3txiqPdd4VP1KB/ASilQi7rX0mJrQv1D8ZUHBfpAC14
kUWWiRJOc261S5GewYiK5yqKADMZDq/nq5kub0XD6L5YFFIvAaXRyLzmEtjJs9Sy
3QiFikzCn0QPLBOrm7lbO2uB8kMejHPPVR1lLglUHgDMn4KIQNSbIR8Wdv3hBXRU
hHoL9miDOW3aofymEAcLUwRtiQZLO9FF/VKYPbiRkzy/yft+p+9DICbcfABSw4OC
0ljMIu0peVmpJp3iYWxCBXqZfVuVlhJmXHqATubB7AYsYB6dsjdh/sLYnVNd4Kpm
ro5KbPtbAs0gtSocyI+4xsJF9kSjChNbQAow5V1mnkvGglvXUAwcoqCKIkZHtAjE
yI85xPMzNO6dZagE/DSYwAvM+5oyvaJtHJ3yEwooxWW0uhw+Wf7Z8QYjVqnVZkxO
sIu2TPmpIoIY3JSCL6HhIokEY+fCBk1cWVfSAi1SL+tzurXygdQLRGPhOtuvIGGp
F8zUtNdZFe6mQa7HW1/R+LkKv/YN9rhbGHNymg88vRNh+gAGiwFrc7mDhvSZd+GO
Nf9lnhvrBbMf4OUf7oWrJ9ZOBk1gqtl0175LvJmX6MAVdEngKqm094B4g9AvwFBe
NCuA+uNIRddZFiG8EQgJWmLQ1WduFDP4frnp9o7hb+xtiks02/sQMYbCdaL3VHtJ
5gT7d7+OU1pxOPzg3owLk9Nu0jkD31u6920PobkTk4vFHGIXMweWBIuo9+1rASJY
6/eStHjri3wYYohQZZfmaIr7bgwF1VdLvlXYRYxLOXD5CBHsbf+jJkJYyPQxZr//
r/SzXCViF2JE2Gn8wvCfjnnVPNCEwyebtDqxwmeXCmeLrZ81+sQrJJmO2C4fepIj
HeT4HI5Ljr1YLrHetqSLrNTnkKNDQICXmBTiWIkY/WtYaHbWJoFS/qyMn4Te0c2y
Jb22Sc1mCRWFGUScB5elIUCsLJDy5HyT9Hl7Q4YsbXJkK7zqlnCgIDw5sL6GYcT6
rweCMN3J4yueBZTxK2NMkeGoAUEbCxAn3NYI4gFkZZDlNuHh5yIddIXLsmxgEhVb
9DfmDkWpZSOwraCod2A/C2Jqgkzp+DBJVOBHiVd0FGBoIFH5w5oo8ajb0EnjSRUJ
95Y2HI4oHDltA9OkdzBViQn7qq54KVZMYhlgFEDZZXI1OdtSHLCPcJXA0fe2s0Bm
XFS6hztn9oZdundd3Ho9wrPC6IAsxgAdDJ6VVXfNVGMsIKjRcL1fnF/dkQO6Mbat
+7nm5hv5N8otCsfNchp1FWyGWZs5go2xoO3QYiCtAsJXDQewSEkSLUxdcCfbyDfc
3knyyx0vVYhxXM/k+5Rbkahwm/Og2HHEOM0BrXlMKrcphGr6sdvWh02IhkPDCm4a
vOf9nJcCkBJLBmVgtlTbLJBd0qKa1Yyu91PDXzrew7TKIcqUelurJfCVEgmzBKDo
0Mo4OFS3P3lmI1CF/sZ27ON3tn1X5NhnO12HBqUaIp6cQy/dztSZfC3TjvmxBNYj
6pWCLykvD8U2p4/9hvErvhGKhtA6IzbD2DWWjfKOkcrLfDZeOnY8AIP7wH3z95ur
3RdRtlmzR23ekvlcwcBHxc/t/fDxSCaWTytCEXnh/JsZPGSKWcPcxX9yYxPV08/H
w/YPTOvGOWW2zagz0Gdc5/qbWS0p1i1rV3ZfliCMNX/kIP25dIFXpL9IDAS6Tmwn
5Yx3/rYDv+NKTIygsLCqpXqDBuSIKXAcQOwjFtNu3UBpUCE2kywKJ9AsxSIMc/Vl
vu1kl46/yHk/XOivnXjiRYHVaZ4UT/jlpPNXy98YudGEeZ5KolgGQSYOY9nrbgAL
s6xwxJ9h6qOKMPHbFYbaXsl6zbufK73QPGEVCNX1z0cbfxKwbe39i+/5KlwR92SA
NsjYCTX3tILkJN9ftH9byN3KMz/W9lUvdh0q7JaqxWnKdtYPc82BLL1eTDz45EeP
arJyQzjsWBEPcx2CbSJjEFKFrttV7qzsrUy+2nuRXaHuycma1ZFq9ZJQM4xIZes5
VThPGg527ae33LUJ+tsfxR5hgpM0qQ25M7x9PudwWS6KrT53NsCmErPhOpycDqIO
OJcwDuhHbCemuK7uSkKzjNflgd8xVWGmuWqINco9GBh166PFoLe1FiW6wz67J+C/
cVK0OmIvTL832QprG66aFE8vdpGInbCT58LhYiP3muzfvLDEx1zOwitKoM5zAKy2
hxNePwVBp2YQH5/Ykz+Vw/mP0jYdp4ljxikX6UVtlIf/TXUdOgQQeSh9RCcHNnaL
M9rsJf3Qsb0OvgGvJGKw7Hm5mh0x5ao22d31hkUgY60wVK8WeLWC6cPgiuQz23o5
aGcKBu/3oUYy8tuxfxAOh1jr5ANwhVwsVV6HOZJG/fmNlaa+JW3hDU8U0ydF/lDx
Z5US1J/4ad3kJeXLjAXmo1YjxQfF1ASWDDo5W5S6MjdEOhjsryxKH6SWKcSjou8H
tfBgE0OpQL0F7Bj2yMw4F18IMu3FhOlrMGt8U980x/pe9GdVfXct2I2qSdd+SmeC
YWjwEe+1qZFSGQERrbSrESIcqN9TrOFwayPN6Ju3G39wwsvQ+/fbbnMAxZ82Q2p8
f0Q+NRdRl7mTsGXSb8fhMRYdR4Z5I9O08lBn07T/UAO9itidQTkz/MYZCn9AUyyt
U7kVv+eVr2doTEa8Cs3rATHG5DuwoqrG/i4kIvI8OCSrI5HmyOEPX1HJJLzSSvGR
t3Wvq1zqeh9V6V8tiLutkbruVVqd2LFegmt+3x+eRFB3by3wpJzPi9O271b9odAL
adWgTbhiZhqApmnNbYt8SGbvoGxcd8ftxLL0IEWgrSyaDhDC5WZ+tlffOG35fyK+
uvunZMr3qgSbPvV3egqfaxdR10FVBrlCUfnWVtKz0TZIyL9q4nVFzv8J/7a3CxTG
dOGOMv3c9Y4fhGGbhiOVrManOfHTabuJUdh3InHOnkPYf0lPaRrNYQV6c+y/ZaRI
MHYjFSoQ+1HTlE0OBv2Tdsa9kKaSp/zpnfABd/q1U5Vk2d51WansLBFQtTK/6WKr
RSkxgIfA22nDmR+BiNeqRFjpPq0pY39COYOJ8MxQtN403PGIGFsqnIJc2BoibCpU
67Sgqmrt4DySBiBwSqy96t7hUqvRHRx1kZivEtJKvprusJY1yVvc/pIiyX2JIb3W
oQ+zGXtMJ50jcd/JrPS/oBGymsBCUypt74oGUufbPuHXAgnuDXVRbU7kdfyLpXjo
rKmbRIMOyTZrtU4UGfFFSUhr9E5b5qTAl0VpfB3M29TKwT2MpMscMk3Bcfo5m9So
6ALVX7JfkBFbMSgCCVxFeAQ+Qacw3YPMJAZ0ltS/sgYXNlJOu2O3NWiZOiuGke9l
uMTM92Ggms6DgbaxdotUCPMlswDVSbKuCRS81/dfMVDo8HIDqZwVyyZ/9o6VXIa2
dP0X+ID8/gEUHRr4U5HpgysxlKpAKCz/9rPB7AlEkioTMt402SKomN27kkwrHPkD
3EstLiFJWH1SY0Bu04XgnNls4qIATxbAl/ueIVbfWPLKQT/x4aj05mfnYppgHbOa
T0UuVZQjspzmjisUTa8b6WAR2DGamF8yJA2ll24ey6uifG+WBN447XblM/XiQEDx
lHizzUGiV6/36xhk79nBA5QGGlRP99+irpexjTgdkGGuR0Y+D6wi6lqykZsly1oU
Qho1mLMSv/irR+Rt0OP5k7QxsoChDXpfM+Gryz7V9VcNndEwEH4+6/afK1/+RKrc
HPDXn+f6L42rUa5wXcrPQoni4wnK1UCasbdY4RKrB0sZz7KlSGKSovGCePRlO0py
/xZ3aLSPYvltjQ5DswXgarntDHyw3CQZ9MLTtGUV7eafUQ/ZUuEsxK4t9fd39O5w
csvw8MWRAF/qY5B2+Yv1P2dmlGTM9F5BNyOXmlzSL5KliebH0RgOY6HEgq+ou7Mf
QnyISFRGdrzT7GZpXf6RgDouHLf6kzleRmCslvrOyWAByCGGwRgS5e+I/renhFDM
V6Fxpw2fAW3rIgHx00x7SSq5xVSDSyQX9imfum9NAhNNwHYnyG0ALlyIojbllbK8
YPaBCUrbxDowKR2LL9zLYnbYZII+j6GTfpj+wGBYPDq9YLvXroLNc0loH5vj5/iw
+LJGVzxuHHEu6mzKXbpgcs/GT4gUU9+lqpbpYMWst2g1ADXc37+Wb8jLyTvjGBx+
L2dXyXVQTNXaP/d45EedZirMhpKj9tI3KD1rwj7r78Z3bNdSAPlkCth2ZSBHebLZ
NICvMsXeCn71CIf5F/LQMWczFiAst12yDJBLgpiGmAnUAHAacgJrmCV3glxq4+5o
ypM0A6x1DG6TgR12aaYLy6ZKvTDP8k2kUVge5jPWHPu5Kl+LSs1z7ThgrUcHQ72G
xSpAt8A4ZeDVsNaBCCPxPaMX2Wj7jnM/gnfbi6dQv0+vGFluUUi8izyPBfH4zXOZ
C+i+6ZCCUvBVM06Y0P7YIbDktP64EIP8ows4ojF9lbUl5tAC64gZlqMg/JFVw6+X
xruQAa/3yzVnpM/mDk8RAibxOzTuyfTHDxXuh1GMIN9IGUOXJBTdgZAI0VQrkBxl
tjEwZXXvm0OLdiIRdNJ2x44AJpEkGvfiBupGuo/J2VQMud2rV0szEdq7RgA3oW6L
YW3mOD6udssuMYMR32vnCH5XbB6Wb8aqeO6dthVuAb1xddv4m/WClR+srz5gax7g
CvSj61Ag9X/EjEkc3YzPawOCX0qTOgRpLPFm6bz8cOEFCyBR7IixhCb92mpvnSHq
UJo7lhFnMIP9NTnz2lYEJ+qMQluRBqWkytpE4/eKjVxir0oiGzBD8GxrsyElCwr1
zBPG3kLUDqKY4vp4+cc9d/HY3SAPlo+MrFkaI82JUloJv60r7YVg6J5ktIeOtFX3
SW5M0OmnlpGJm5HHgf2JEHSGvEKC9Cr+xn6xz+NZmixdpA4mKmTA/BH1JK3SmCeb
O6GpGNj6ACr5HvSTHcink5TR2O5V78JEWVuuvRq7HB6ZeAwCbOdKGD2SabvY4HCN
vx/Lm2FU/br+aL30wAlUUBvyX8L8yAbvUGp+H2txVLjKcwdA1czwiqwZtQ8QKnRd
dAyFypQfygjnWV6fpzTWdDJMzfyntqwudc3DwX2JZGl3ps87UL8+91LukO8DcFNL
r0Wgt9/DnmxTlqGnIs7nkZAsRaR7eOPJE/TMBfuv+vU9AeKf4utR67gA4SEKBHt2
fUYmiP91XuBK0n1wjlVeCrIWLZcTInnvdYGzXrxMIbvX3o3ivpLGamdPuSrJXuSo
IL9dkX0rFca/kMf80TWPTdGAMsN8R/ovTBaaxP+mi2ZQftPmpPJvJ41NmA166i51
Nm36Z0oAj0rwOfkj+4BLSojgltQhbjr4yfLZXy/FL3l5CZkw7XlRn393p0N5OA7P
kMyNc4PvaOacPWQxDazOIHo3EEZQGUbclt5K69orvnTnu58rRU1MDwWxLejQIYrX
6qfUm1NCyv59QNOc7T0uMY53W/GrDZpQRYtWGMZBtuVfgyOuDZGmVMdOVNjCGZ7Y
UATE1+EFTvg+7794kJZsWZaLVul1+uAgZm2yp2/csdJnpWK/7ahJ/Zzz+svphDTT
a01u1mdnNTggtIYeJgjMxxL2YgDXbKAUXZJsDcGsVhmJ5knx/OENAU6PSVy5xAtF
RGFct2t54Qt8gkZ+bCy6I7oyynPFhjvR00lb+UP8CNmxC7sk3l1pa83BDxQe4KhH
mAIEH6zpMl3PM37XgtxjOip6iEGQiKlE+dPcKSvddtVHuIk2ls8V8Oo9XeXqhTVz
1VpBqOhOJStl9LiZ1HhwEsKbN2PwA/qWwahs1c+n5RBSezqEngRKeWUoZiOM8mXd
R2cKqNCnk3Q/7x2V1zk0D9fOhu7Uf4GT32HmoVCbuJZAAtC76ALq3bcnssMy8KCO
m5bC3z4ie/7+dxsA0oamqi97kgMLbCHcnyTzU5m5fjAqPLNyKrdaLQa5FXlemXOe
1IXU3erOtlpKCML9mk1/b5KOfX2k2PWbfCjJxSCQXxDg1ua2SqBJ10/j3CLSMuqp
YktIRitXMMKzESEmpZ6AnkWpe3o8bSPLVfMjyR0CSyZr49sbXR5zwvrLKWoxynIM
eUrpRx6hFQys3ZurjZIYUQTaT8hrZ7TfbsaZyP9ggpgCzMAGYx8mvicz/VMzbg4K
pBJTXlLSrH2h3BpBq9z04yzu9ExYhjZj6Dcxpy/x0J5nghE8p2sQIQCWS+BADOZF
uBbXNJplfOQsBqs5vOJN01YBWJoiOtEvcAIzoXqoVDlLTvGq+ndT2X7UCUuxUdkp
u63hbPGVfW3sgXT+Kh7UL+DZUmrw5R5bSZOQpPHO8DpRAg3IilwE+TUhiLzGFmh0
ee0rnCBdC7HlOosTTdLLtXgNOgHbLA8ZG5VCwB6Ij/U8R/SJwP8PN3MoQTsAQ9bi
n6dvm6+MVJOVXeOxqBFBpNr8fplyU1fm8XkhpHSh7P/peEM/K3vbCxq1RY3UK1iu
NU9eXvqDvTt+vb3UVHnwKjw1ilaM5JzKmilrJFIDYunfbPvCTBZgAZlpWnnu0Icx
K5ThMPeABIDeRUkg8T+4K6FyidmdXV3BQ4fBxkCQKSaulwmCTE/PdnX/ktvcph23
5khz9r6rbGPdiza37f8PnhS0V13dwOop4dGf0DlJtDR3kudavj6i+Inr0T2W5vPB
WMDIQ8CJc33nzgAyxH7WZ+N54sId02UDuuCu91zekVPKLGtB73oxr3vtXI6+d13W
ZSiWuKEgfSLBtxQg1B+zzV/pJ5OwgfkKPA05/XwKi470XStmKyqjUGxKy63yfzL+
W+CXYqYkWJSvlu0RYEgtxZcYaDnQToydNYljNznFfjmLYDpvt53jJS3BYHKQNQgo
blr5A99jJuDytb0LD6/6L9tN1R/w86OjCq+aT/HUlzR5kOX1DfgyZSuQReWysuiO
JH8lRdLFsibtYpmZI8cNFq1bPG2wCLrHDxOpbovc6MYW+gQECsiwh1OWd+UpPHh5
vysFiHo6ouBwsJHOCxytOrqqiO+WYAxDanPIS5ov9v/99DuOhnJMNiMKKvOWyVyk
uC0232xYQXlWNxW9Ajz/1uHqCeoo00NwgvZPVvA0/2bEH0WVChUnXW+EF3XxHfjT
yNxc74QdJWLKhGF64w6k1dqKObtmOVSZ1LZcaT6spy4LAX3NRrbn1cMwxVYc0iPv
pcZVQfEqFMrHU2Isg3xFNVcYGzKezsrDF0BXsCNoCn/g8vGzZSCSYyFg4RvX5rSB
P9WTQG/Kk6YM8VDGJqh6NoarA2Ormhsq73AJ+cHsI8pMgtAs8A0rTQzrMkk0ooyO
xYQs+9fc6m5HXf3tjKAHzTr4A38pzbf/vJ8+q2dWcJGAA51fusrD0O4G3GAvfOr9
WbDqA2rTprmkUzESivz96iaPIYWU1YPidWs0gHjLc3uvS/4kUi0BlqrgB3m5mlZn
iPpQU3Ih/987QD0KQaM9I5JmxCbqWjurMuKi8X669pJnvpFqqjBW5yz4SYsrVY9h
MqOyqzd/L4gUK/xx1/2Xbv40j762mxAhGiH1XiF1BRDtxEGlMWLM5k9jSugYzoBK
EFsxkjUO7rhtd3Jls1WAGTKOYWh2jthdsA7FQ+UFLfHk2Q778tLLI+IYEcHahemX
WgV7ZyQYSIOK74W7pcaUxkng/9aXd6u9wq5CGjlRiHeB7LGOge+ShP3JtynV+iw5
wG/1FBsXyS/IKvWhD5Zsk5ihUvh/TGZeNxFmSuDJxU+V89Dr2/LHh5Zs3d2EIVnl
x9u/ReVtYV5W1FRNA5jB/QDdKrsveSUQdq0HAWxM/uXtPWEUlyfsqNPDsLhSyk8U
XT8rTaF/YWJeOU8KuAph0iRdFrooso96nyrqpM3CYbTlzSU/5aqZEXjQqrFZzlQE
a7GFqo2s39Qp6mXNJDDYFoJksoU42W10PB+IyRITs8MWiqEEv4agM7ZQpR4UEIBA
PJq9t56cxGKjNVD4oMscvTjw9Pg8gV3Svb7JYr0SkenTrdle3AigBjnvW7oy0K3i
u4f8YnrZQHtKHlU3Hm+sRvsAek5sTYFv47jmYG7rNWEOIDhrJaJOtkSGEXeTNVRT
Ek7pf6RBxG14iVYML3vyhMSgWR8ZW7lT9/uob4Z1/EJJYLPrARFGPl6oRr6v/Usw
xQ2Wdz0LR8lUhu0/QFxkZI7UH8YILFQt09+MZnekjOZEJYUogM0l/NgVxjYpaMM+
eRJ0j1/M3UnIQVo0UeyeRrzBOcEWBFE4vGs86D57fV/fIzn7hRk3YMvqgWMVzajo
ZmBNJcevG4D+1sw58xDrrrMLiJpIp1N+ekDkNattSLUXYrsPMRVlRaULFOJjzBZb
T74Tiv2EphOAFl7vSaf2TgfKYQWVJJOYAI5FCzFxhEbm3vMTBSJWR4l3dX9ioRO7
ih1OZYModqV4pF8pCP+S+m6OQ5uAXS8a9eYTEj4ANIGKw3pGXUBovFBKFfCCFD45
AlAKyjbi20n3uPza8scD/b7noxOSvPHjbaTGOTCWQS0h/LAVSLJd2h0ut9ZTRShO
aqmYK6zXoQwzBjkEqqkuhHOtrFjoZ4POxzrl/lDi22EcdxpCFNOXaeg8ixjFUHoT
fIiYxB/1VgzLrEud9ugTpP0EBCVCUuqAiSqOqV6arSi5SKPCkPuPTCJ7OmpH1YR2
EacmKHGQIZFc+xx58MP4AkZbyxIAgpn2H69ZH6xzocQFNV1B/sFMfq/VtYBRXHul
igdGIU+GxE0AGU4HQ6OdzSHWhYN2Lc37yKjyX7Jd77NWUFbaSP6yEznHDO6KtcFv
pZG97QrS0e5yhnSDeNb4AdFqcyh8Ko3zPrkOWPAoUK3c30JRmE98+mtDNZUpG4Ji
CEYg4eyPZ0t+0ZeiImwwjWthXIBr/CCkWDlxsClvA0/HWmIfw81N4OwtschID4hq
bzb1iCliYdijYeu2IS+4i3IwMLSBLDQZaZ2EPFH8v9gZERdlnWBYHtjLud7to871
EqFX7vKJE9eLBnsiq2tNWpmsA6erBbCwXdwYVqsaA5BZ3qC5ezF5LfC536u3Beq4
yFFrenCZNgL7k4g14qU8GZIdmIhoBQ4XmFoOdNisImIdisiKKiaoKluN0kNg/0dF
yYgW1Mm/gg210FPwlYrfzJdHGDl61b9RNCSGbIcvZt4F4zRDPkDYQPoRmmtrFUN4
/FOL6F566R1lTiHTff4a/J4xhLnunQFY5f5Vu4cfNylRz0Ks1PTqn+3T60dgAcw4
eXvGoW4MZFn1WTBXJ6o6/KSFYZty8LlagylVuldhC4ViW+B7FDkwsXI2GCf4rrNy
OsW4fTFqMOSm0ETZlP4mFHqd547rvLWlpvFcl1QBeSm607ttUJ7rYv+/TslLfiJY
YVO9aXSRzOUO1k0DLSoFrXWxAsAmWyCX4r3edrsXJ5E71CFe8fIIbK8cTNUM/c3q
5xoWkubJWUGIwdT5SDRwjUcn9qGN4CfC06U+NlQW90r7p3RIlvJNsfwgwXq0imlP
dskjb2m2dqfupworBceg5H+6ORGeYMELrI0IKrF0PJoLwCi/rRG6EXa7R0HowLg6
a13431/iaiqVbBFmD3CqmlFRAIjuDESfgoT6IBe23EzKXECSdtO/Pfymjw9pIrZA
e6zVnCc7jDEtg3BYazaCgLlAH4VsA1e4Z6VPZbU1MDG6f4oL3sm3Mn+O1xM8+s8Z
RTs7Rt0nn2CNwO9WG83YklbM26Vuj3zPr2/IwhvnmipXFBWa6qErlxi6TNWWc+E4
0CnRHbweaX33qCYAwuZXLPFHxX51ovF0MvxQVs7EN3ptk7NuL93wzkaJxOaPJo02
dY/Zk5MPVNh7KUnPL+hdTw5lzW8xMRxiTJmKQ/4llIZPpmTk6d8BZ1PVhY2F59fl
BpDArkjC/AV+/ITYXPXu+CcNJMBJxOgR6QzcIcBU7XP+evL+s4iVLv56aQwqK0sK
YGgNvP1B9M/Msrwx6lclNMTe8ylriQHg1u68rIz+pmiziYMIITOCcuyXQdLyjyZm
nT/l6vjK1FkpsL0CEgWSLPBSjSZnCL1nwwTujGvZznKxbXDRs55KCs00uFq/6T+t
MV8B5rccxthbDaNgQAw5SUV+Rzy7ZsA2dbmx+0z5NQZAF/NIiDoYxN/BKAl/pquR
CkvefZINUDruCQPWEZh+S0VWQOIvCOB3bDNg8FZ/n6yOien3XLLikdtnDm3etCbn
OD/+tEVMoSU1mCofgoCO8AXHOppBS8hKnJ5pt1LwVCkc3u2mRlDDkl+7a5EIhFm9
2j7DtYDCMQ0UTL8HabSJJtyFBnbJVoo9TsO9JTEXOaJAxmkBBG13QWRUSJMqhDZ5
tfZE1L6exgqEh1PSUf4icjnuIJlYzJTxh13UEcFrA9cBn7HLrVuS/Oq2AyKcSAhP
fZMA5LLtMjunfTCzRPT44ol6SvY2O1MmxawawKmXdQcGuSM1sdaaNvKpCLHWzdaC
0ndIJfJbp3rTT0OJu8jL70E8gP3bio0ADXddEXWpPXwlPpf4/0VohbCosmY37nYF
KyffeAeL6E+jCImM/5VnD+alStJFndtQQHV9xo7tP7ClOLsKPcvQOp+F9K0Yt9Ih
Xm9QY2P2+p97GXPQ+DlyiVST/gbg+RRjJY9iyYbo7x9cR0YOvV/I7pM5+oM0HW3O
XRaq9XPvRQeh3WIUsBV/mDEiUgw025csxI1rdXNm4pad8ExxbhjrEWOaIM2TJEEL
6Fi2n+t77uI08yHRaKaLlGiXuCDSdA1zS/LTcBadA+rHgkEXkD5r5elgTwZoq1sb
/pLmae9bb6h/H+lAJoO0/CcUQV0cAWEMS+cE30ILV8B0VNa8vsBYEwBWkQZfCGXw
jEfOj33BE4yfBPqOsrT0RXXclw+6Ot9Ck0gXdVJsT26rDVbsR39a95DF6iDifDj6
2rlCDK+xAq9wodDaxZeFYUVkvdSv1fOPIqFgyQA8A6rvYnNoI1m0aQIBT8e7hlIa
U49rXpClUPA/YdU0n3KdWA6c+VMRXx4t9TIWheThNrbhSTq46kwGc8rQXuoKVhVO
hIvI+5cnBC6NxNTVFt2z2PIapKoN2mSThKV7475F4DHOtfycR7xT6PTdLYQde6+V
irkmIei+TZDHHQs9bj84Cdq/G0MMGc/hM9a1hT2lXvo1seDi/lqAsjyacVzzYvBE
HwArgaQgXWbjcPgqZgB1CjfUdYvhvmT7pEMve4jkIxzVJh6sJQOHkOhoYP8mvhXt
CgxN9ZRy4Lu1ki6uOI5uz7KCxNAR0dDGSID7FbQYOTAl9LSLuZG/vifqoSw42WnS
PS9rlVFph3+AVUThcM7LJnNQj1vKuFjZgkcgvu9E+RO35f0FJPiGjFiZ07IZiOmm
rDLpy4jkJmfpBcCwOyn3eviKV9V9MHQoY0Vr6w/CqUuVWOpyvWHG2RHd7fXBVeXd
py+AteHHb4KM27Zp3r/RwFCB8WRWg372WNa2zeLDflStLNyMN0Hf30QGljCzJi8C
fDDmwCtTUbJw16ZcTgigaLawerwCHVN3M9ptqTYVOAoG35NYtesJuwDE1BNR0fFn
RPuj1jj4trLhojlC7Wigv2rGqUoF0xeo461TENTb7dF/yFLPaVQtuauMC/zHc7cd
aR1sLvr5gyXzOXc6Ye+fEjUulzKWxkfHNkymsb+ybmIXX5YtBi+M76vO3yXVXB4K
qmqJZAl37ow0RtKpKqiU6/EvNkM2Eno6iVhW80YIjuvPwAhVvR+k/zXur4ueTtLV
0YqcV8p2T5aynfBTWaCFJ1jE86vhIDMzhT9BDphNHFOqmR6y9nQ6VSUj2f/Bxsav
k8B/9UUU5hBo79YHtLTem2SdEiHxJqwE/DUEJmjtrxEWHTKzYoai1eI9OczN+Y/H
eoo+fCd8EJ9BRojSC59zUM+9I+lrL6WAyltbpHroFBNeF/+LeOYhi/nzySYPeKnX
dIt/R9j5tfGhp+k419nRUwsxdxrt/Rb2IiHUiKgsmJZBDhOiUSK6nTczlLrwHOEa
fOkVKGGNev5b6MQxCVUwJzxydC4ub7Pd6JKbAW0HYD6v8hUiLvVBzjoKh+Fq6aF4
B8Pzs8CV/tPdIcms9UtmEziUhxDqzmrDThsSWso141XIBekPnXuRr8LLeJvJQrq/
wXvSQT3PuTjkuC1eeF5+pHS/pUjRGckuiFO9hLYUek3gmMmzEEBdfzcxWVEn9Kmo
Kdni3HyJNn440xDRxv8PN6B9AR75AEbi4IZxwUVo1eDddDvxEfJ3v2x50Iu23Zii
pfy9yHOWqLA/f1itSzmqqm+/0PuwtuLKk3IvZqUJ/OjwskxO/oSSSYu8gIDBTKBD
djhamj0Aka5X4qTArEdzJmleMjeT2dHk2Gv5Qpe0h+3EhI8eav+V+MihdTS5/l2x
ORHGAsn7kvMFTG0AHhPiSfz7KLSaZJXWcpKtREHH8nOKI8f0Pd1RhNwAz4x4Gv/Z
4dO/oiUCdR0RxxSoskJxI3j/pE2i/+LdbF51E8bxl1o4hbR8XA2XPZFtNCUGF5tx
ey2aaeT3IUNreNE7vsqoKUJlHpBp1bcvEnlh4w0oIsomjVIaD5fqFvlkXQfz3wxl
15bs++vbpHriXTLVh8HDeDmn+1jo9u8v/vRVzKZ5QHscSCuyxAjFzue3UuBt5EsX
wNoR+vKyoOqaYMviNVYCiod8vq15guB5r6HpS06922ElSRTxF0IDfgAh3qtIj+VG
qsBbG3E9dP1GW7oa2g64+9upAJ/LQevN8MokIT+MRAvDh1l+pe7prW7kSPcqSqNo
gz4dmfL+DaQHNNe9XWAuytkYbqf4tqaOAM2fYBaxSg6fuzq5WPiRtENRcwsYyLrF
kebtTsq28m1wD7agNBoXonShncu9GEBhdanxyOltADWjhLirMsnDhmvHhNEQZsI+
oBR+OT1YZkPMxlZKppeM8GRjm4bDliuUftY/MvkY7zi3Uihd2lXEJd5oKbxg7jzl
I11zkM895kyVkvmYhE/UZob/wA3xFBx5MaF06dg4uzG+EZHaK9fvonOK3qUsnwR4
+EVypnjhh8TRPPXqHfPR7HAaUdC7O6BCyz0Ao6KRBAXovXbLJ1gIwCnlYs3Kkp5D
jbNCKfgzWc0DYRq1wCkoYafrKuzsE2uWskK4YDr8s4hGDvHM0RlCeTPaObxFN2BH
RYeOVQSCVMUmS+QXbSAiJz6a+XrusTyjL+N9Mm9tmEqAli9EzpohkA/+vIhmwhsj
vuxQ3HqYU3DJLS/0scVRIDeNbcl6KNjKYNbVc47tXJ4I8nblxullYAD2IAhI4FUW
qLzKyQZOi6degUwFR+APo25wY5hvLKXdHeTtNFqBqAQUOzykOnrWKpT39taDQJ9G
rOZK1PgAcnNJEISDS0Y8KNEmc5TQD8LG0idh/shwpK4T/MzlHcIIzfa8LiPUVdcn
qWtRCfP/VAzp65TQ7CDSN8YC1SzzQXq0nQCoUv8Nf+qCSpQMbInF7nUpCoQdJTwn
nXXVpStxM/0ZomGArFErgtcshPiYUg5L/kQbeZe8+kQtRqO8GvNkz6JUcj/1zZRf
8m1graHmw5WLJSF3kRVe2iV1xGRuEE43mWRcY5I4msNzrjSfpMGBHNGCygeqlxCr
fhuNOFa5Win4mZA8F7H9cnH7zhgIg7UY6+Gqo3siPQALaqdGwEjfXCFkdKCL1OTm
M+s8wfiml2G7SRwNyE/+bJI4L0fP345A+xvuIsb7DSO7+9LD8D8Ok2PeaNN8lb1O
Yju2AGj4IVVz/vlNMFYjL8qtkhEmXhL5A0vU9HP0lVknke/DqUHf2TPvRvbzO63T
XXJzxBxF1OSU8CVbRCKDj6G98Um/ZQpWjZsUJXG00BIYCo8M294Wnr35clD6NP2D
oWMpuZK1hgcJ6m1+xd29lV0XcsSeK4XHNwZynW3/bUyhWEx3qp4baUopQSokogKw
hIAc3tLoOg3iyGmubCUwe2NVGXPQDz4alV3i/f0viHni95eOo5697x7NMdUeDWPO
8A7VDdZbdMHVewSGWSeN9CUEMEXGY39D2NInwZ5Rv4x1a19xXBgB1qBLhPe7yS5k
nYozQ20z2t8WEayUP0kbw5nVXFc7mrlJfmEOTCEwZRW/xZ3TvkIMD7yGK2ISS77P
YyAnm4g3/bLrhFdZR6nj+q6nZh0sCZval6lBdi7diI26TYiIQJGZP2FVCXkB8Ndb
fmsT9vacotJ+rdvTSZsbvkRVmrCeEfoeCUUT6Ze8oxA0l3FyWBKC795rsVBfrG+5
3CMbF4oUxq2vv78R4cepkxNmLrU4vgYkye8gGvrl4vEQW2tkS9sPq2Eepr6H7b9n
LpkoY3krjMFRiZeYOcruot2rANPGsPTBqgSQZMbC6uWG+qBpRH9AUnEcQ/1zgv6K
hqAO63pkAQJFPTmp+QbJAiOqhoABiN6ZkhXrGRy5l7dbBpYh0fomxzL2GcvRO/ZM
P8Vxh09v6jY764sqHoThS5h41sYL8ajfnmmleRFUn4j9i86lbK3J31GNPorB5Kl8
+6Po/cetFMfHG+I/sj5W5Pdj+KKcHuLSQqjgVBgBtytYqCh9y+GB2Fkor7Lfj+Yu
EHOR3EJBc5BKu/fxlpG0EbEdSSUXX0EIfT8r+Fe3vDFWNtAPCkzP1nKCVjT+sT6c
IgO5p17k3eRo2jmJfn0VN0O86i1yx4q3BaySQWYQfkITbWTKwUMMaRKDZCqsJ2Iq
Pbfz8uGLRHirc1R/uN3CNdsgsAIDmSsW87z552PHQJu4gFZDDNn/w+3ieaAWuW39
uEjtb2jIRP2nfLenLkc+Mqr5vJWmxiXWi3lm6OSDYF/DTKiOlgT4DSTtuDzFmpZi
Y46WFjLnJA8HFtzpTyyOn4z9/d+CbaIQM/WM1cf9dnAuTnDF878G+TJUJrGgmTVZ
GAEe3/+1BhxhwoL+r2SKkOv0FETrfkbN6++cLP52mRNT5Uh/imQ40Hej9nKVLo/p
D+GmScGYPY7eBKhavpfVfHmugigNdC5Upaj8HSiEaI8DbZKi0KD3J+Bm04TVuoI+
j9KAUJIOLIrOsurPZ1LK9Zyn++jQuobF29WZq9OP7WfuuXrD+TKZ9THoClM/LxUf
pSphk7jw3rOBI4V+7VhCjEguYNJvs91FqANmStJZuuBuMUlJdOiHrPtSTqBfOsbO
Exa9zap8A+oYFFDqab7JZVFF6EsgVk1EL8axeXUTRgxXyJmEF2KDRgRSWCxvtWNC
RWLuBJWZnNXHt4dU2PYdrDoK+b64GwhkHIaBPa6egk0bF72+9Sh6lht65kCB1HDj
QN/tZUAwImTcrp+pHp+QpPFoBE3PGDywkc/Ib94Kkd5iPskAEX8kKtom5TGWtRww
h8okzXF33z/P8aLE1+IvPaziEUZiYtFUGiaN6kC7jzwyYkpGA0Xa2NV/RSKBRJcZ
ldQhMYdtXQzneb9SQQkVWKl660to8pfV5oADpgXQAa0RiMkF6FNbvBCxy1UIOdJI
S6unKZj18PNDDAkdJr8rHq1+EbxzMCJu0VqqFi6BlWVRiCESXXFeEn9hHyBSW30R
8S+1QL7KBdyb2nk9tAI/RIM2XlEfHqUGVW/XJJ/GcdDZQuaZmyWvIAk7TUp8Gczf
3azNi/EAfUi28ozJK8PoVnkK3uGvTcFqVUNbPWx5Io6D66+Sm3clsKqNkLBr2qrz
4+cifMU/RFxP/6ieIrRI8X1F9ivh7JEAYDWZl0UkHJaERrZ1qIu02AXtAmUBwDa4
+3X89DKKTfyHYXwGyN88LbaDFn63QLNdMmw3grhGbNoWsrO0FJSHA90GOafZhL0z
T/q1ZMIf9ByKj8ZPJCEyufMZjd39W2XP8gvZEhsVxnH3JC9Neqn34TXrKcymOzir
xaQj+bYW6OLhLB1d+GTq3lk58Ogh7D+2qYK8PhnmkNRa62EfWX5dRJ9vmixcaqFs
8Uo1BJWVGhyy0RIMsDKlTVpy1ORfM8M/+L/ZNXkqJpMRYPKlvFBP/qSKWjk84DDE
RpUZF78Tz7t2FEZ9GZma8OUkoVivbsKcRHV3Ev8AcQagrhKNn1InhGk0tIY8NZzV
IXCSH1ElbpiADpIgnXwiRyh2Yrz6t+3OgAKG60WRZE/J+Go2Uj00Q6nzu1mM3bfa
R6y4GkMVWHWVze08qKKrYotuwvxjjXBU1bpSu19dYgx2eA71k41JdaT+UQw4DfhB
b+HZN2+9F013K4/m5b9sVtTISIcHbugEfUoNg6GfjFz8AMp9ABzbyeOKrJQJbbVF
ImqXu/4Ru78UGkH+EYVnzIE816lMtJoztBQNNd01kvKGj24DaJZ6jPz/DcwARniz
YlNoUsNPB8l4OO9QRMJAPOPhpLZOXRj/Zi0ZG5vgAHeHWNNlWbEcZfEszPfAyct3
9CWPxjCLE6Ck0wx/aQ9YKMzwVhP+jEHq58VsioqVCcPvOB4hLiRpTTHbe4UUBPbI
EgjuTQ02PIJqPhMWe1+8ZvD01/cRv6kR3Tkm1W0W39O+fLZOUJK7Awx6Adq8N0xW
IUdyY5rEHJKLKZrFehFgru26aiQ2iQfKtYvcQdcOeIM7bwTZYeMCxY2EahWAOOZh
8SrB/U9q6oJKEqyEPEghIucKclkxSIaUjfSukb/Q9sUcKabbHqkqkGEggObdttwu
zZT+QXdRbTuJcxgaSXkjwC6d71VMgZ4cluFFOXB7xA4glhuYOzsyjYdHRhYiIXfP
gE3eVD5DUyhRdrpE3pJ2VZ3815xoXgWJ4I9h1dI9Ej1GElig9FwhuScuOn9Z8qtK
rs6Egom/x6vobTTAEjW1R2lCDu5qBRuOMxBa0G1oOGBEA/cV+YQmSJ7qGhC1e+AF
RGSWKGz6PCijVjZMWbKLUq6ofxEMBTCuX6BIORHoPM38XSJo++2Jy2jJw8Qv2X7C
xz8DGh5l2l3IzhOZNl1SbHjmBHWmg6bnWsyPEXATNQmsfWr8oidQITyWjRLO2VjP
Y8f8xJ4YtRbDuWTOpEKNG6dismKw7Wjb6VSPXPp8BzZWmDjxsnqJptJEOPSlC9VA
KLF50fAmxmebDkMF9KpHXYKA57PWz9b6q0jN01kHlXCwPQBrtPIYyUykkKDbz7BS
DKqK7pgi0TcX8OeriN9w+ZcCyAOpZ4ebzJTBiN5LcKlWtRiFWWCVOuH/lIKWzSSz
IuIdICTNm9UQFgoNH3N0szVe65UQYO/Ck+dcxaX05mDriD7bRpnoduQEHWZiHoCS
hNON3Nv3mCfeepNAsTPdxq7lAcHu4sLCbrBVQR+s010DNQi6ei+L1LGQEwCKSLBR
0LZRwzX/SBjPGZGwa2eKIqwDtBRGg9c9rSA/IhfC00Fdk0rMlcf4djQbwFjgGJRZ
0hLBvxPtPdqztNrcB1w+FVo2Od24Z8tN4erC7I2ZWKrX3rkgcOWFEla5RGkB3B+U
HPl/yKc00Y0NQhUVsQHAF3ErXqHy3wFHH3o6Nzg0ege1qlXOmy/RClXQWJZMl/3o
QpmtFfgosUIhmHp+7Em1Vd+BY0zbVz+FeREW4e+lDVw0OA8VtWpubja/lgsMDQVu
7ZqFNMQpe2bu1fRB9i4afi+z9UUgO1I1GZvZsgzfunaKkquWiT3k8AILCG2d6Y0m
En47NlpWtyUeOzldB14YxsT9eGblW3IIZL+wxYT+bN+XI+msZd5BAU8cugbW67TC
8V4DTiLI5amvcBuWR/h8q+UvSF8THsBkPg6ddLs8WiHzzifLQQMlltXlfNWeO4Ow
UkI+4RYZswTqkxz+6OoZvQ2aJLfRFBkydHkcnyGgCbw1llAUxm/Aqsx3zn+ZQeaI
DgWncQ6hmBfT08xa47RHp+kkfsVZ+/IALpMuLtQhc2ylHXF9vbHoV3TiGHDPAuMx
oRJtDOpUhqdCbnM7BxMZ+4wpqU/ShzzQ5V0FJOgrZEXULdreElpv62bLozB37jau
BrFkdUqd0Ts2dXgm8W2uX15gGbLk1ax0ZeSIU5helmyaECDTrmRcxEv9E2eR6wJ8
3FVkH9b7xYT+T4g00jqdoz+jw02LnvbNqUEsr9OktJyN7WNu2vwXg/giNYcFYwkI
teyYv9E4QSn6DQBOfuro7wkh4bDfBummtis5+ZrOSBhnTpzzYIqvPI7AMv9SR/sD
08SPTqKv/L6JAmSo5cQJoCuPRSLIsKWWE5vmU/bpbQxhssS4267GDur1/sNTUEZ9
5TUXXSMfvs2j1owWy7KdjOQDkeTewqyO6tmbTIFLaPZSJPz0otsaxmDB9aHNCyld
MMTFbDt6psoWHGo+NG62aOkVcm28hMasKk2EwGqh8YRQQF8m76y8vio5o9dIeRB7
OTEiPI1GmTvk7OKEnIkiKgkjHfXDR77rC5tIBvD4OBVm3Mrmnlyghb1uFvWc9ae5
b3GbUuDn+MQFo4FpbeFMgM6A9ksT6/rGrBER5M3y4O7x8WQEyrj1b6nbV2LzE2V9
8Tl9Fr0MtZQ96UzWdVdpGnA6Vi6Wc6WTpDq/2gobCa57N3xnC8NxZ240YqUXOgvw
f80EdBG+TMM+iJmfZScYf338pfYWkF9GtKWyzbG6oUUdS+mURH4KKdaBD/I71UGz
jQokYSo2pv0qysRIBB8d22JCjcMUOSlHj8II0HN0ijnlFUbjLpm5YOmUzY5b4kaz
dy4BAtLJ59CU+W2hX6I/8cjBnPDII/g9ExOMvwDImoOv6zQHMPdVBtZi0N0Fdc25
LkuUdigqMjiHb8/3rQwGvm7udogfoKSFl4ofhE+feXWVCtDGo24wHNmILw0ZkTS5
S4AVAkNFmTJQSYuR7sNbU0qcYu4RwE8kI8cI1t+S4GyZJ4Z7+c/YWS+ZJJMQEp2n
6E3Y0IgV/4dXpo39FPNtfYWs07cTo9UKFKorYQ2QB8sF5V/EVVw/SYXRiY1OTLJm
QDqSkf5kyPXeCi2yGyvyM5m3Kj6P900NkWlxDJWmPBp+74mjvxUOLSkriYYzma6F
o3rJPP6FTveyjeB+LWz9LZykmfXzJaXV+mhMYTVcbPZqGkh97aM8weIwckQCP0Jl
bjDD4t1p7/cAeF3aBVtCZTcnENpUFohPHFS//c2/uWl6rsoExeeLTxC2caylIqeS
rfhPw2rOPzoPx2lVtw+9MeNdVsbUsys1J8KDQS6VR2WqJlDYOzS9Y80JbKBVDpQy
IcokOfjRvD2z+ijOu42Y9E8JrDUaVJOysKuNEUsaD5/rJ8jVHi2XO6g+tLd+ouIw
ivsOlq/GJlH+BfNN6fve5co5guhEI9IMjJtOSOY9yseRbwkImCPRLziNnVslTzCu
ErB5qYn/HiaUJNj/cryjKNMLbMvRVHZvjBDrDqVxRh2GxkXpaHCt0SnNsgvW1wxL
Vetlx3KmE3W5hTwRleE3szp90hgR26GjytTmym3kh6LHmhTgNz4ri5GcSRnOiIp4
KtfLOKCj6nS+GLsekPcXzTpLBG51Y7EHTYRse7IbikFQm2RSNXt/l7NrrskGSh9a
k3OtUSQWExaiAboH0txY+aRiZ3T0bTMXrS9gb1Ys+q1uBGGMkJHMj6w5Yx/iT40U
aCU+M9CtMYO1THzJQbcwbPR5xwlGG9fyYZb4o69pCXrNLhWz5zLOxtcXhLjiilu/
uNjEEtpBl2nkOhJx6UeuxRhj12Ii8y8cdw9zNWp8Jn3m/7oEWXd/EifLGVrCsYWc
/41V4b6N9p2rLDlgRqfYX2v6/g+nC9TBPK1v3oYMFjV1J6O3wepvnI9/hp7HeYvj
MXWpqgreblnXXTa1mCQIYVmMfiyNFygKph0tPcosY2fQdWHM2jyfNHjZ/Zyzlpo4
LjcWuDqgoNRiCYqZR9JUJQk3qcQ7799rWK8PBazYTvu8hmF0L9zxaRyeI/K+HhiD
89KUx+uGlR+MTtkPS9kgbLNexI1W6fE9vEZySydBfLP6S/4TWbvwDsI94PDTnT7i
wnz/c2pXjNDvoO5DbtGF+ItePaYHPsmkzSacYuEo1uu1158Qz567fxO4ADPCx+6e
fSalyuzQZ1aol/ZdBPcnHARqhinQdlkAVqbSjlzDuAPlRYCp1n8AhVPv3OeoM8fV
LG4vDsxcDHt/He0+S3gt8MLV/ZSPnFxVv18vkt1lXpzmwbQtsj4d1qkD/rHfTgCN
t+n0O9I1Nk9An1rHCuGGPM3kWXHpMz9hzlsqEr1nsTKZxq7CoaJAflerOq8wfiOP
8AIqBhdcnNCmADs4ykdJXmmbhDXrbTXp7XGn80/cnKv1U+z+hFi62SkgVNq8TGW5
5flw3YbxGvezHvLix9KvZXRapbJuBlxCByjX4r24BGlX7m2ot/Llq9N6QXpNzblZ
z8OmRnuNNPbrLeVY+x+hF2HyiVgbral2HI6VThMjU0KE+PjWfmRvElI2fC0Gs4hZ
uMuDngoIgMZ9Iqt1eiuBUJVFRNEZbskbcq8PtvLAvKLfTIiUgG9sShW2TxgCITen
JFMbjHriL77fh6L6iaFQTimd8zOlDr7pCOTPhFSl0M2WBW7VLX3Z+ajhmTc+URBv
jR5GjmLg7+FJEVqZxe3bWGm31xfvtoldTk5jJ/sZ+nhKMauoHevMVAGm8/JOuHYA
CKONqAnrL4sKnO09jvbPnDbRD/kELuqCJnI3IeD+/3G+KEUL+0Xt+mNDp5XbPVdz
2Z8spkkSg0dtD+EcBiAOjFmQOd6x0cjcEOjJOCTrbMiG73RrkG243STbN3o0oGjr
bbUfZfxNVjtRz+ObUb50390OKrEkNCgYtLBmWnVnHif/RnizjCJzCa/FftBt5I/K
hlNADUYAYVlxTEFqbf3wxlAmFYKT+DDUKDCVdc4nK7RkgVZcibFyvoxFvGPrayXm
jPjSZYHNF1UUxHcAZrSq708U17vGbsT65hZGEKuzuTMpF8u8u1oknclmzdAdilzL
4azNQ4/2AEnj/i4w0iyt+R6xwGsdAwXp6gWSJbM02UqfpquXuLyiuonFxQkKzUkK
6nP9HNuHuWZo1GIC7n1LAom50kEyDpQ0711oCswQiHa9bm5jqnLaLmB8tpATQCUy
3Nbvpgmkmt1tNyW5Yx67wNKtc0ktbQNw+v8Vfc/uCpuJi7fagonpR8hiuNxPX7Ye
WXB9H9sYgTmFXga5YLGFASwaWQdV4Yuyit3PX2mh8wkDRSeZoMqAHtOLyZ6W9Vaf
MOY5yx6l+t1+rHVbweIgm3sOgO8805EdANk9ZajIYTG0nNmMmT7Y27lUx8u47w4M
SVPp61uA/AZ44leD8feTQWzGEHZJi4q9KrHHLI+kLIycFoCdTX+Cu0ZGovNQyBZX
SAf0VmTDJKJSGBb11C9h1kn2ZFQ8yH7Nm1aFl+hJKJO6an6ap8Y1HI8HTJVnC0mg
U7MvO63YSp4Li952QsX7rqiLKCOD1Sgd0Rh4o+sMoD7x6ge9KEXCNrjkZVcJr6V1
s1R9LVwG7+Aq8/VAgitLHert8FwwWowyibQMu1mIS5eFje3L6T3dmfKYSJI9VCk7
KWLDbu+JBYYa0tNlDyY7Hl5PTLjbBkhvqH3OYB3Ma2+Y5zsPa+Ve5vUZpySSZbv3
Tn3sky0if7ISy/tl9vqaG+XMVLziRr3KGqgZfMuILqbnrkqCdQmXEw0RPBr1SRV+
fQNlzju8fVqrKZqU+hNUIYYYZDVdKAU/5zrZKBFSgQsT8v3LQ8DoXaw7YhOPeniX
tgV/aBtipgDyRwF0VwBRK0gCEB2vMbxHtXpRJvZ5Mslkk8J7EJJUoVq87LbRYhv8
D9ihy8CWLQIxHDU2ijOhsl5qHPyj/3g1UuqymAhq1HrPHcoNtrEHqJTnsOcGSUfL
eQLL9WQ0lgsvlhh9utDIPOBoYFNB9gR66sYUwQlECzBmJTPajLU7Tkdde2J62Wao
iwlJNMLQKPaRh3HtFB9xToUwQ9s7LJmLMdc6A1m4PFHFjfx93hTkFHFn+iosFxi5
Wtzn+3oUClkE5JhV1nZ/LCoeCDhF8hU4c0dV+A5Co1Spe2vjdFVCyHhvecueQMGe
t84CsKU8LB/j2+V8r5bUAQ1cHRv4xUJHDTdoLGAgD8M1KUNH4d7kMGBBYYBNJ8Nc
Alf7mEt76t5UMf3l8Who9S5h4TvqlJIi66NrWmk/1jIOt9ajK4T3BlXzrbCZw6fQ
eZMFnZtKLSyhhgJBFOziOE4ISEhzK4BDjuaycSfM6VlAFoKU03d6fMDk3cDdn9wU
KnZLytKKu7h0eEz+1JtbFwMrDlZvnsP6VSPlinowWY3TacqxjU12SheniHWXwUWJ
w1qhIdL1FoMY2nAIQB/5HjTifurDnHWqVqZ6whtHM0npQmDChzUGIsSeTe1dZuxY
qe7zaCxF7eHQX7f6ULUyOMsAXEoZO+HrEOo8Ilj60xdPc5KTHEWdIqLGxoPLJGNu
gbbFTsUwdazEo3QDZM7K/AvUSvp3b2HBzOgmpleNzhPn/sgd2VyAYvatP2GkccHW
CS4QmmSxpyR+QR4w+Zrmme7FVv+zhRZeqXVw3xdgU2JKzGVL588UYJGGxGxUq/cG
YZaHi+TwBOz+7GLNF7nIuh0taG+GE1SdY4z4T19bujsdP37p9jjMZ1khYN03ky3h
qh1Bwa6iUvY1sfIPd/mexMDm20iv/cZJpFA5JsHKe/O2TFpGQfN6shQ66H6C7LcR
09yZL4vq8tDGRNelhNx4gs6j19T+YCwOkaqmNBII9aO/qXaoj7SGhAl128lbz+sV
UPKODg2aLYWRpcWeDYqYH0eHdi75VI4l9dVUfszFMlMeblMcSwCnNWqVX5VKPuTc
0geRUW2FJv7JcvkxuGLKplAZk41sx7D6tfcHGoxIeF8YB0VZePWz+l2opvXYuD45
3XNiYF3NbFFNqW2kx77o7qUajfk0f42b/fixsmO+TpofwIiUd4IOb9DP2JUUCsaG
l4peFaw7cdc14Cye5iC9RUKASD817j0YEW4CQ6pZPxSFBYJr6wedxFk7iDouGHF/
jsrYemB64ecrj5VBtMTLmAWrCknmqnwaFxUsi80Iywc1ptl67E2TTmGL6nxrRbp2
2uTyf2xMsLYgzWQacHpJRC5wpiPxtpDvQmT+5DQM5e6yO3RURuKlsWPyMnVPNmFK
Hrq8peF7rFL32r5Pw6/lDPIO/t2pyxA5vngYIV++2uPE7IjclmU7W/6o61OwoSJo
RdBfCVAKTjzJJ1fHCFoHBzq94Vmtxt9AdBTavO0VF0BuXkce3ZcfJQoVQcjUgJmY
wQdeOkzWq+WRrb4FfwXss6XXC/hxLdk8QU4Ah5z4uLV8qtUtHXFCzNqX4i01OFDl
7fkNchoNNHPRX0oJRp9UgGHSGbmS4j2NclTM5s3lyZOWDGcl2yZpWpFesirrhIsG
nP3dgA7oYCjCIuKIPukp/sSKg487dUqUYQJ3cLZX9dFW8oBpDHwIUWG/mtzj73bH
X0y37joUi2gWKjSsPT5EukKi0/mceKV8s/xoXyeuXom72zzL2WrKI0T3a7S7ThJb
m1TuyM15sizs3PihE0RzjlmEU8+ImYyAVbefwKbh8slSSn02aGKOH97MEnyb8P2Z
yoRX3cG9RRWq3KXncvQYlHpgmpm23TLdi/C4yj1pJULlDq0DsBlFMTI75wooopG6
uAtkDPDWFlcQr5CeE/KuhBm+cNuHV5N8ZGLo6XdkwP9gOyjY8efK/IQjlydWf2kO
qP/jSfiO4m6trGabnSQk4VD5B13ckrU17+gLKeYnE04YbN0JyLcCRneZq3CbGaKC
YtFQHJ7Ja8VbA+kDM0BqpXKT9VhCOzUJEPRnNYZFfF4VS4EUckZbpbJwCHFHGyYE
B0UtNXu5ap1oLnVPuvI8Ir4QpS8pyJ/MY4MHISzisyDw6582xL+qgF2wQGTc+Kp6
qLO5RvdxAHbqMNxpxgBk50rFwq7K6131Gbw5WYsp5J9vjJOc7PQ719+u5GJ+3QI7
qHLDyYemA7va7stz+FeFMiSlBv4TtzqAu3bRGvcFd2s7J/SqiywPlEF/VOOxegHZ
eA+kPN73hCFIkhTBxyI2Twrj9tRMgC0SwumKpb6PudjM108F7zL2k0kTxvOQkAZw
X6xPglqJ/1Qn3UgkWUpH7qd6cf1MYR38JNQQwTz4NqJ7qCGjMQpdJGGmQLwGMye6
ZoLIw6KlQx6HQ4OAGioQPRWbzUbiEwkmZNW2J4JbUNyc+B9/RJ7H/oogCP3HXz1Z
lEKv/8vdTV4UktxUCMu9hIHJIQibm2ov1pnPElg7lvHsiM1+6cTqkdXcpaOdvqKW
UyGuloDmT23neDuDzVkIh/U4yKQbyb2pWnfYW922t31IaxQjH25D4p/Lq+Q2IUuR
OQJ0PUuu3VrqJiVnwsfH8MKvLfTVPE7tccl00hO0wDALBeW0sA0Y1IE6E/nqdHwR
U19cF8pHSQlsnpCwyLzZAMi3nTocdRfOMs8bjiawXczQoClEIx3OZk5jWIxbkitm
nP9WNsnBktIEaJVq87sPq2h6Dh26CeN1qL6Le7UkLQy8Zkry5DYMr+DXljjlTbi4
oo8DnhA5XdMacbmcZ8AokWWx8/KXxvnQDYSdG5OtB7IVQuxwhjDxzpg4LaWwzObX
PqJNHG5hPYsR3nKzJTXhVeOYYKJ2N9MOFFwdgvZTh4CXYf9kwYBC8G+GtbDTfkje
9i/cymQzAbaZzx8w7yEC2Gwc1yor78aJ9g3ubPYJ41mcxJOezfO+smNjAjykDC3H
IwR5QFXUNR6AlTot/oaNdwgn0JY0T7Zm6h1MdrLuoFkyVlvPrnWJHcZYPeFZfR4h
nunS8Vl02d3bc0rLqz2BXHKoQelPUhdRZUH7anaqzTQ9X5ACV6F1SZ+FhhSRbTya
x67i2XiJPieYM3K7Opz31MuvuOuPe0BiqcO912ctbu/jM8PmH2LpJ1a6lt65733R
T+v3JYH4KMbl4/1qPl0PO58Qydh0xpOmXzzMxaoViUPPeaWM3Lfbq7oz2y52HlI7
QqzS4i7yM0h1RdhK3BsFvFgC7qhjFkzgDeWhF8XUGwZTVgiUEi5UmJyTSQY+9aqa
sV+wksLq2mDla7GNZGq0Vw0Ygd7EUYGV1YQzQrGjSppNoZP+lizegqfRMCBC0IAb
0kXmMlF8gNCYcV+1KliTeHhoN6Djj7Gg9ICttg5fZNwCSCOTMLQxtlILFpfKR4Fc
y46JPtRDxXPLfMBx4YOuhFbhDHxl2tIk1ZIfgpYE9UQd1F0mV9+nGhBNUBLPSOlH
bfo98mYpVE2dRXu1FR49GAmwUIpjQ75rbp+gfPqBj/nX5SYhGvVnWi/JJrP5OhuP
9ikV4J2E2JxY6sIKQMiGvTYtlb3pPd2xcnaCwAF83XVDLFB3VcC07bAHTbCtDujo
qKx7w5IQPqtFi5iz2Y/I9qF9HK91SehoH6QF1gsvvYcYwntZtOEp6uw1HLNAwE2O
kV3Dq8q9QO/N7fkYRWN0V0XEJfZH87NQo/Qva0i5ge4ywW8W0hWeoaFRwlWSQvyn
u82nx1TGo8vhj3IBLzCCnEE8OA0AJSfNX3j0m9f9lR0EeVhRJl00Te++z1kenxqL
m6ILHrQZ+VUoA+D17yZNuwI8CArqN5yR+9ctZBteXYKsVmdvhSngavlc0JGksohm
5BWhgUkxVGRCipAV546GhLV/JkATN9J4iIQIHcKuA8rpM4C1JLs/FJ0biWEgqrK4
vc3ADcOOiznT0/n73j7JZsFxyE6knimN+BcCYpO0XiodUDO5KtsPPbBcOECoKwGX
c8p1FX7d96msE3TcmvMQzi6q/a4GETF+taqfEBeauTGdCebfiYMEt+YNS4MpgFA9
bBMdxfu5Oa4q4mHQfi6dkoyJ35SfczN/mE7RprEVkDvkdwp1I4ZncEARJ1kQ8PL+
+NnOTiClC4Wn4T3hYoH50dK2LE/wlBrJFTNajUiwDaec2+F73SnWCRcP3rxE0i5w
1+Y8FXIeC/laDaTlsjZpbNzgfXfYUE1WJPAmxk7X4OeX4TFTpT36/ji42Bk4as17
z9GfcH1Q77RYXjI0y7Qdl1M/FqTYw8qi5AYzvc6+uIy+IrLHzgX8l8IkvUKkg7R9
jLkw158NFQ1FfMJ1RoyytpvO0bDp4L2/l+Nvqr+jnbRqC+3XhG1U+xb6R1Yi5FZA
MqTpFnqedI6zUYRzfVO+aneE3+DrOqT+xrSUfqiid+OUa1KFQPgemKIljfpH6IRj
uIsd1avwaEQkw+SwqBNpbz1dgqi2FczPg0Xe17i0PKBTaw//QH+IO2/MH3EqsW4T
n93M1FBwL9LoZ15Alf+/mtgLbVXM8cBB2BAaFenrBOEAyB82okrrk5dQAnPoNTtr
zv63CHFyisQV5PEklG9T+CMqUbgU9sx8TW0KanuUE5i4cQPgqFw9+dMN855WDNP6
4LHU3GaJxWfhv03NI5q5wu5C6Wa/WdTw8q3K1Uto3fGn67C/SI5fy327c2vknxvW
oNp3uYvGfGPzLYjH+2nwMLxms+lncRy7EcdWquYCn9qYk4Ea65SWTju0m/ReRJN6
3WkHJwQlLcra6TAy9eq0xNAORY7MNF/wVjok9mU9dc+G1hthEfrv7Tb5OGU47uJr
dtHKvZVg4nkyO4KBjYIJTMkkE0nQ4chv+blFIhs7rtXyhEndSqotKKYdkzB7QLiv
xI4ofkTOB+RbUmmLRSqhs2l36+qrbAz3Z785isY3sLw2QS4onYY5l2gl/SHaSiea
5fHbwhEtXxs+55GvhxH/qs+co+qXVu1VVS5gPwUrryr80zLTo2fKoXM73ZsXrCPQ
Ozx/r/vQFpCvyTrsSXU0Eklzl+YKeHra3scDSZasWFcM9izxdRKMIa9tF3/ALlCY
YiRAryMC9hswvoxCgZv1Mv+svfNDdWBYsT+KRI42oTB8rl85V8GOYBBpwqo2BBB3
BW2GeCgHHqHF0EANn2sD4SU01YYhUUJfBXC6wfJdKKl8GJaFhAeO+bYyf0EnQo9k
Dg/Ie+/lOaX/DMZVI6QudLMyiDaJB6Xn2l8fgq2cdFvrBhpAfdqfPvN0v826jZ5i
zDbVe2RWDm5bRuXeJy38i71nQrtDUpPILkpnLtkXfMZXlNPxMcQZYrUsZgDtpILu
nVHyVMkeiievgW3w0h9tYJuruYM88wHJLmNlgtFQXCcx1D7AWDsDTD665+vhKXep
ql+fBRTYXz61PWRbpfJwnGqyTMHHk/poAI45Bwxn02VdXZ+SQyA5FSl85FiA3WYE
fAVjZ62mM8Z+RR/AU64MuK8pewHKoNJrw9HD7lat21p9Zya02gLxAFux3lku8yLV
wVIYwOzOPWbQtFGhRAzkBREZTKGzxnmG57dV3ZfX69u6JQGMWYkYsTCzUbW4Qi0i
xBZcbudTnxLdqd1qucZb/qaBYtzkgVgaoUt3XcCDfM2Em9vRaW3NlU1FYr9Q0ymv
9h3FV+8vNGE2ktA1KzpYztwOCQ2+4o3K+6nVqLUbETQhmLLcSWQI1jOfomAZwSwN
ynTdX95vg9XXT/dGZ8mTIAjEeV7t2GkdH47efstkegyIuRIC5QA4nm1vv9E/skIh
8f6Xikwo7ItUmuCIx04j+Wqoei8OzNaLsVnd0W1Xzmpplz2BK7prWg4yoxZFSWXZ
NlaZJKYmhHqXslfSnl5Qq6njzXiAJviEIJ76nqAV9+dxgMre9e7CAZEgkESyUPxL
8VZIXnL8/TGI1yJ9Y2e1YeTTaneTWCNqaNutoHSDUlE2fDReJSy6IGy4c/yoB9sp
kZRlVcr7aNN4L9G8XnFjOoxlTnNpa6SeHCNwr34Phw4rX4Hk7fELubbPH7W1L4xW
uTxg0Ds0ZyFBg+XStD6MD5CEMvOdhbL57DdnEV7oUtp2MLnO22kDfV2pw5iYB6TH
UYk/1oS54WVlZSg4qvaAUaLduVuis77o5zA8Cy/4PhHABTcDtsVP/nCH3/R/NaUO
iWSV8uKW14tltBwQLwFimMA51SoE2seTx3PKkCdVqzme+7z2PLJv2GLO3fYO4D82
3LkRHQKf990gPU/RXDL6OgMg53LkaBU+2hJ1KbzpYSKI+tcgdzNZOHzQtRTMpkvM
upRplsUqnHLjfmBaX2F8ky8PMvGTZZWcw5dgmcs4ztvCxeOSvhhCbdetJibB/SJE
qvw/dLhpCbe0sd56tYVHHfz+KzASlI5haYc4MSW8L4saJWq+PvKCEtAgBXwq/hVa
GFJFx++defK/nmm6h/0nuDF82JIJn2vwtTxnrEkJ5MT2Nt75cAp4xc7Mygl34CkB
mBxkjmxDc6e+fmtdLPtNJCtbDnTxUPP1thUZr/b7aQ7CC9KWmCLGjsZi4YvcvHzf
+30HfQbGPMz+097miIAxrK0n1mNRigm6NZDDdxpaWal1hU9JQ0gtiHbG7Z1Nq5FQ
lWCWrx5Z1pNFjnQH6I+iR+shAN+vOtGywG47QXG46XzKvHLxSTuS3Dr0065UJ39k
M8mH/fyRRD725mpzsYi/QzIo2/GD0jgm5ySvCbAO0wdM7yWpb4UvMD9zXR4dnzAk
NsC/LpIQr3/dXXCvUSLyZkipJeBucL8sUxgKPZGm2G/hx33664Xgm8cWU4LVQPXw
bsG0cVxxNSUO1IIsoGnXNxZpsIXV9hV65gIBZgBcYiFIwDnsIgiFq2JpGTnbDlJy
m78wcheDCdJQnmYd5WJ6NqGsJtWJA/RBAfXHLFuKWlVw1URh7Vsy2IZS9AGABCKp
eEXQ0+typKj6PdvuoWxhC0paTNnniNutsu/y3Cz+o5igJqN0IRZPNiThHpOxiF5+
+u5Fnpy2Vd26u28Nvai4ltrgRcRV3DsXBbuBtFIrsolLJMNZfCYnnFQDm5btCTco
mO3Rsu1BWz6OhjBO41YfcT3AnqpE80kQ8YHX0gL2d6/QdJuhBNEzhXOEBcy7xDSx
GlgAsk0hU1UgYK5/YLMStB4+5q4sHlJNxRqzZ7Ztk3c0H9QvwBG/8zGx7IXcASYT
RiRs9csmbY9qtf2FrrPsuz/F7mVb7i6SjJTJ7lcGb+d98rQE7jSk6ZAhjT51LwBT
LPzR01b0omUD2OFT607s3DzXyDz8iNifshh+DG8XtNnRHKc/jkQ0aFVBArTvwhS2
asc3d0ymf90uL83Ud3G86W+qRSOUoPHQwgrj+aSqQVb22MM7oPrA5aiFVX28SJGV
+X/R92oF3Mo0Y5VZjzTuTpPpqtrrLgrf5mT8HYUNLbkCyFJfEbyxapcOFTdBTZ30
lVmODXIq66qgMnMeknc49rbRZ2k4IV9s6X29kw5wWwpxYyfFIpL3p/eJatNbfhYQ
Xye18ndNr2ZQJKNd73VhcCN4Z7VpCHGUcjrHRWo9cSmwdFlfi0zXccA6N1sYnl/l
2gAvY4R6LGZQZ4bzhDOXEunqoodtr6IgD6SKcZ+TYWbO5rsm/ybADeeg5kflGPiv
1NSm6Oz3Cc7c/M2wAMjUOKLwTRWr1EBTWB9QOnBSQQng6Bn+OCtPM9lmufeU0IpY
+xEyGnBXBLpyY2wEV7+en7o5JlDK6Vwe0aCgsNO4F6HrmpHBkZ1DzC8AnS1qBB2R
GbJneRgaNydFiupXqNJqir2rK/wDQlqfYQm0yNY0NNr5D2Di8fAVWdFsFqyl/fiL
p67WI6mYCbaszUhgq9wCma9NZ3oXTmGh30hb9NELAqsYRuliet2DCN+8/5ok5e3d
xbXtDtzYdbrp/u5lSHzFZEfKy61M24nS94JE/TNjj3uT53/mpxMnOHtVq33pj8W/
7N4V++T9aZ1tasfFp7AAclxixfWULBApjT0fy1i9lrqLxMwLefMm4kkj1WUrmh/4
/u+WPgE2v2W5tnmCyh/+N46RbSaVRNhfumpLVsfiImoS+YC8jBOJqAOEjS+txbgn
htqKnpkuibnacJ47RksF5d30avEoW3V/IXoX3wG20EzQOAyIiIF0ilsMCY8np1KQ
yaJbMFPXVMRu5IJROtK0ILjgswfJNfgl1Der1BYx103cMPw6ymv/Ojq/I3mqcdl/
3PeA2Ksqp9Q9yE+EU2KCwcu6IIIgdDkbPlAZRBH2P1MYh0Tp+QKqIKbBFqnA4IFv
EBHCK0NhGNu7hZsRA2DaLIiCHVg9KUSBWOfMb4yLr0Etidu2mF2bCU+ufiCNCPND
pHjZjMWBOpHs1Dmiq9lJT7YnqiumUESWm2CZp6N/mDEvljgII9ZvX5OAS4ABfZFp
8BGTfoWlydP0V7HxRhCtEj8q8qrV+V/KSnAIyKe8VM1rB1j8C11Ulgrgln7yU8T/
GYEj+cXoyZuDMIzl7iv6W0t/7/5CDjVuEMHKgwhu5XcWmkWOWDDwU5E+LoVd3Waa
ZFf/iFQKB3XoVZgkPUQgOu39lYSIp88/SPukPom8w6kdjRrpIonzErOkJrOsNhan
L5KPOgurvm5/my856kySmfIxPuiKySgs1U38qzqIRdbUe2AxGD2TG9kP01bsrnvX
ZN9ePOYMvEtiZc+DigdEq4kQYxcrqcnaEES6JRxXD10JCD2YJvRiFBuHpz3OQFJH
mpepK/8jCh5g8uCC2M3ThN2O0D+bULip5z0U1nFcmHrasCdfdnm+qDSlp7z3AcV7
Ht0Bi0J1Eon+Z27ep3Bdr35HY92jBwY/77y//PRXyGl4UZQ8536FNQXimQlezI1I
8IDrdh6TxHsCV1uJJnPniEEQIziG48FzDPGpIWWMScjJ6nuyCT0min0rhoX1SCpt
mLrkomqLoIxLITbcdSefXc3id2y+8gR7kSHdp3M9giOkqHhyNHv6t/ph8fN1myed
w7eQdqjbsE8vahlEDJ4S7OCqfFQ9ey1TbWXxZyVhG8y7ceDhCxN/ZlO7NrT1lAC+
RVOCFN1te2eZ+L6TRGEqAge3n9BccNoKHqlJTjsSY4Em2c7EhgWzJ8FyyE4fYQ+6
54cSk4mOKbV7YwnF9dBVOpVcU45csa4jyKFhGny8zOJTp0M0uJPwXYRvcGrgqJ5u
GgTWk/oaEK0NNk0YlcS76X+nLkCiCwRBFQsA87Tbgn0Ae5dwLIEoT5hXzhcutn/8
CiqwUoPwP+14bjhk4sjjsBnPK905DJu5zeMLQWihyE4kJsY9GU6QJRIcUgIGpXQW
Cq28TkzW7Bc1tCw0XnxBwxqF8/QBUUCAPGm9jDxG4em0A8Z1M8PRcgoylUBCdP7d
rc0+gDGN+VAS1V8BBVoIluTsVW6ay1MEam5trzp809cQh27ZkosDt6WSo8u32Re+
2x256cNjCFZOjJVkoBQMrIGe6jZvMEeE8uliNzj88D+zc954q1Xu0866Wa08CBGA
Fb3A8dyvotxdtKYQLTbZ8x/PPx1+VGx5mwB0Jmg9J4PypzGyKDDhaYyk6ujnofue
p1f1tgIgWt/W6iO4eub8iJCmYoaesNqwlJ6IWwfcM2a+1yzJ5X1QKWyEAxLYurv+
d611L6Gp0ROn/M75o+rlRqEwbHg9jsY1sEzQcWdCAqPxAGgX59ISaKPCtkxZU5P/
VTIk7BN5ucAPUMHnmLVO8EJLZyxV0DAEOGplXLR5MpQoCnND8pdTD0mKXXEcz/Vn
NfY7Goyu8OhiYaDhDJSLhODZAvPTwqvgfxZvKgYL1n3LMPF8CVHJoVfPWGBV64qZ
Xmap3zMiiJXc39J7JQwD+Y5ybx1BUQXOO/LAXgaDrM5mON/CByl0FVnlBZtIDOCU
eWVS0OC3GTt0dt7xK1ewSrunkE7sAffMoj8Pplgeee4gFRtKhMk4rnTv21UKhO5a
p9cOARlqIHK8nLoEfIZbTmFTA+KzSZgDpD5z9NXezEeCdDtzzB7BaglYqygIY4D6
TaIR6k04BgKtyzIvLvRetBJcFUgLM6D3gnsN0G4GMXJKsWrGV0xsjI0yTY7O30IE
BVHKLbIZzZu0I25pj94YKQI7er4UXBhjLlLpAvNpIHdcO8JNs3FMuIMAfRP3H7QY
SJcIE537PkW4tv7xCAit3wxgaJr4BmJQYPyyd9JAkg6UiXaw+pakX9P2QM/EooIK
r+g3bopSAyWkWoDiS8EfkghxmeEdb4doE9scRi0DFU9u8gmTclsIKhVsocIhD/zq
57sGIpHS04t5WOHnG4+fRLrTrHL47MJ+XRqHbXSdKgLHMqTBpO6lLPO01I59djYJ
by5Qt1KnFUuTsQcAKck3oY0wbToCWR3qIsSK/nFzC1sMSaeLCAXWWL9M/kYcvOT6
eLkbi63n6U+Omj0JcJL3opF/dsvfZLuiKoTcft4DUSxkHnK09eahJGqBo2wgBOaO
7WMPqmWQGWAL4JR7Ld3XrmSRmlzZbtxpX44yJ1aGz9634BIPlR/3Xwfw2kZQWFJR
w6XNx9/Qy+RVQ3JjjzmKz5g5sQMxz6CUYwTUd3dYc3X77pex2ga4NVDemyBoUlXA
b/CNdxIEPthXxkKUq7ys6C7d7/zvi1dJPnPZkskHWBvKt4dWiB5OqsFd3COU66qk
q1LMx/cLWN/KFECMum5I3jDDb6Kk/c/lDTJTGjtRCY6ruOmgJScY0CD8cqdIhwDA
II89llkUPE5hzAH1t9L/ghOplJfJ4DDAHRRbAp2R5FjKl2Hv5aSiujrtbBd27xmm
/zJY7h8Tf54Vrk0DxWWsd+4bUp1/z2h+Qspdldmd67apaOegQs4Fv6uPL9edDAp+
nMCeoPzOthIa5hkqsYW3tsjv3w+M+YkLDnVQiM4YvRXTVzw/+oVXekPYxt22leHJ
blntg4D1Yzwu0604e5uZ48r6LJhjFmQMBe3dUdpNQvPetFjHYnQjcs9fdZshvziH
3hwOfrIOeZYJZMvF4Yv2xdOJiEvH8WzH280+bcNiIqLJHKV5cTcTKMObwVoasAYG
wRQ7YJI3OpIiesACH6uIlm5M7WiolCT0TdyQXD8f8QSOlD+8vTJixQrJAJmeXSOu
KJOe6B/MBTt0Nwt8WmjxhSPHNnKTKXxMn55fCwUn+SQ0EJ48r0rMAP528V/WgLCv
EDjd6hWMHZ9vcUgzwZ7WiCg9C2qMiHRN4B8tt+hHOB2G5TOKMlDRwh6oyZOSxl0Y
cvuB/vuivDHuX2MrMQlHeMMcUnsL8OBnpLI7Dh/sa9LbA8lCbU8Fr8T4NS5gxkFr
evLTsVwvW+e8a0yfiDMI5XN/70hz6TrSu6c9VniA1vE/jr6ceoL0UIYcA0tiFF/z
VClYvurqqiGXWkSU8bE+ZJN+YklyX/WgBTDnZyZ8bxlwxbK4TItvIxkLprpXImkq
6K2l2FcbJg9dua9znLVivqgJpORDKAtcI7E+y5cBzvTMGcz21YFGhuiwji9/M/3U
TMbosNUsUPGRVCd7Hqy/RNG+ydLyu4rhTHSW6MTchxBsfL6Ngm5QdVAE7Rfrp3UV
3EVPcDEU3ExjT8bpbSxzZsbijlcFjoBiP043TmDJkp+868QsTryfc43buff5BHV3
46Do22B2r7r2xUyw+0XbiAnOmr0WZ1eWzgSPvZX585pDHidR2cs6RyEYbDXoibAU
Ud8O2wBDPDikiH7OReBnqVB53KFGGXPUp1HOrqsdQLgStvnFSUxK3884QGvv3UUJ
uuk2BMOMWFn7rwv1p8sF81SqXuR8je5LlZMyiKn2O+W6b75JxpGeAKRp2ytHqKcg
5M8xsIVHsGwVE7xx+W196+X1hF1ozOEZ7y4sINHk6diHxVgdgOkrFKhuWWxpRKxm
xcCKqVF9fiTsGneHE1knSBIIZHDLsAaCL6GHfp/blc1urqwhUBRRMSDuztD3+vX4
ICTWWkHvWveKdKuBxwVwestVpY5pCaN0CZ9/bOvxtX3FbK98f4FlrNE/wt3foxfq
1T234xyDOElc1BL/WpWr3bywVjIRdFnwTUUQF9B3YMN7P/GT7M+nfTsHn9pGOn7j
3PK706x+aOzMTLoilCmcVYoZbXQwkhlhCkhaZOdvy7NeawzFRwmZqPfnwl1Q8MPo
ia7OSS24kdik9FNnuvUw/uIi8IIQDoXAxiMeFDCM/2ps7DvO0mmlVBYkgHayqQ62
PVJGUSQIICZU+/PGVkIqQWRToimYPZkHTOFBJ364LkuPrd3W+9Kedx/OhQ6paYHw
z5X30FpJ3dcw9e6bZbUenqbwUjPcoxw2jKbkT+OPyq+9FpORlXV/Rn8TMHe2sKbn
rc/+rCmtMUcCsrXHqZsXkPXa5Ex8O0YX5za0RUz5tSut004zT0FuJDKQ0X9lVMTr
Zc9bN7cFKLNyPvSBM6SU/03/vhTTMxpusbnVyCquu/D97DLk2cRxwoKKIjW/04Y5
1fazV/BkXWX57Z28XJGOeeHxhQvag3n3oYiW5FvMx2ZP984QsnTfTPvqh8FWOl+8
pcCOaHX+UWsmzCV1Zytyh/3vf7GrQXCvpyyw9MF5/QLJmDoHGX/2P5hW7HDNevqO
f0PYqyY5Oxzy3Pg5ta1eFQAG8qOyZm3iIBT/qKv/WJKsd9fd4OMldr5E17IDN3ld
QCsDxseOOpSzM1ohsT/yp6kKbzaI7rD5CqBARQVvoUPfKQ5Q6JCvgCQHYM6goR2n
1LxiBhqFtETn/zkCgoatJeau0gaLPHeGzbVW0ydXHo0Xr+ph2BFOOLiMBwK8Bu/D
JT9uY+8PhWDdXvvb35I7Heoiez7yExz59HP8rXP1TSHTt4kWM4WJX98O1IWpj+bl
fymQL9rANXJt92GLTZMoJ03CwCal6IH2La1qGPuF/6ygF/SGbqXKWswNgGvpcnpW
P7bce630BTfEZUCbKposyNaUFJjd2WOwdQjABetT5cIB1eSbvS/MWY3MUBqXcJZY
wO0/+8MdUkZKLJlMnUgLuGSjyhXi3qnohTLTCsSI3WUOBtFUjf3cl3Txi4gfM5lq
QSwzond8uiEXe608+bjuzcF6jZ/lrcFRJtJowR1+HPxL2Qe1D2UlVkXXvhNvFEuM
P6Es4TxtZ2cX3/QyIhTpItgwpijWfzEWvfUCCLX82qXElQ0waB2TUT0yKp6gOwsN
YNMHn4SHL6+yPWMcefJR6ZVYCqSPMO6gY4/N1fGFSFypsU259S/el8ja9qCyLm5Y
PAl75xDfV3+NL2O8qJEJz/dSQqanGWOhyOyGXAjKwxCa3VSBd7lU1vJwo7mzcx7a
MEpzkIjIfv6vg3Y0Qjuq4Y2j6TeflsuICUHCME+J3cfShvUmIsrCOYVjZl7XTU/b
34B5UMSj/FQhnBoarAqvDsJi2tEOpX+FRpt6ZJSMlbggrX2SejtMfMXw1TSPCkj2
QE5rYNCLGgLw6RMbiAIp5vMD52iANF0q1QK471gTmue79TN8p0cgsKLLYuaUI581
RP+hTXNlF3DpM13b/ekUtDn5ge8gCfeR1SpDehqgUhXtc3kKZc2bTrzMeQYMNduK
Q3dCwVy1fXCL5Xf6LcS3dfKv+3VxQm9t0XW7f16/8UwbacyfOQketz9Nnl7NJyXw
z20FbjfgFbXIIUaM/Bvzv0234NAvLSMmAihBKSqibhkqoMlBS3r6hX+8raW9lyge
raHtQc5UhryVFL1KiyXyMnk2Zat/xvzZZ9gCj+pCYYA7EkaVA8xS5VoLZIo9KZNJ
Edi0SCAMZbVYBM5cCOfILvWUX8/iemjS7lFrxC10VIt6eW/z24duUf1kG/EPlItW
9tfUhp09/bUR+fJVgG/CtqQTaa+6z7AduS8VHY2wpCYdScOziXezqXCRHAu2iZqy
Ixxkb6lRojckMXjTHxgj9jifQlt0ND0CZ5GVSXsEl2NhK3dCyPQsfDHkw2gaU1Cu
X0gVtzVOo+RhPQkhs20rouWoGFcJXxqSkUnf/27tcBLKZRuKp1S0F26+c2MgPgvi
+R8qMrxksb6W6cPAg0Syj0Wv0cMfPq+9WWEp4ohh9sGeqa9UTjhiCNiWeCYjQVqb
mS/dfYB09Oq3ZLPXMtkG14HwBe1lsT1zLf23rdlgbvuNjE9AAWVCkivKatHLT+MH
ZqyWMCmSLA/MII57Y93q+yGZF1DRGrwo62TtLg2PZ4G+ecaiMVIs1HsIcdh+Ijm3
Qyc7qYjgwZ+x8WLo821vTSBIe5YSCsp140shC0WM/zVEeG6j3lWX9xNTguevgWd5
KaVwCppPfPGLpBr+VuUSUeCT0oPWzczJD3fRsEPWpIQFEfQMMrYRWLvLiGzRUpGf
L7XKhZ7KOsj0Sm+zM2wmpermCxJJf6H4Ar9V4I/6DbTUV9+YZ2xzuk2vaJ1Uf+Y+
/b2+E+WqZdpO06+nyy4tVGZ0+K4L2ZftiRf1w5mZBifgQItX4fjU0cOU1KVmsfmz
uqhs6nwakXI/VuUsLEbTVV38MgMjlWFAamMwAur2T2k5ZYqLL6UlTXS2SX1XWgCA
SXqY2RwB8438M96obBSpXyh5jAYDQIQcAyS+4ReaXTJu/sA2/5CHXoXW9vHYTvU5
+3xm/I/Lrd7CQelvt/Zr+XqhWTepx8tRzdeG3CjMazlBSAH3Au52LVpNOnPuj2L3
xlGptnZgHKZCMoOhVI3nJSK2Q7G4NUd2+YeeYOr11UOhw9suGM6evCE4QhCZxWmD
MeMIVPeEe1Gd1F5m0otfMjbXdZ1LzmBIlDNGOryTcgGz1eyQbMs8rGwNSJcBjCIg
n6Xmcsc818Y7B/nGRGoNp2AM/eHuQ2O8gzJ2q4EyDLduBO5ar6kuN6ZkJpMYY/IL
PZ4RXHFSUbZ4sEv4CB69v5UNtrYmznc0XN6xK63eg4gZ8JS2vzwivppl3u97Oqyj
13VtO7xZ+/hkagYIqd8SKzcQpo3oPsm28ex+Roaxn5zxyXJlpOA6jNhCHli4H778
rTcj5SG4gebyzbIubtb381c4dghcgTgus4rZ0qSw06Tqrqc/oR8tR57dh6ttFZJ+
GWg79h6flP/ES/iQgNtN/GdUY55YhmdOtJINI6z7Y7A9UZnPNS/rd1IjI+rcOx35
kgOR1qgfq9/l7J6L2f9d6MPyzwwrIVlgEVC0caIYs0qebKvuA00Bqi4syZ61tYxC
ru+w5nZglvZc5DpUDa4AY3lDJBOnWmsKNQb5GWJv/HupZRDUtdNR1ju4YOxEOf3o
F3iYezotLmL+CyLmDLnX5xsHt7sYFWnqUnR/M0zZRw+roKBB2y/2RSNuXl22UWZ3
QarFA8JjqJEG3byurVHAVQo64A/7+tqGoFjooQWgkDe+4meYtW6sVRcmH34d9sM6
vbXHQu3jHpHmqmVzolWXJr/m9fVrYgHsRs6awOOcf6kY2d5gzZ7jbHF/+EwZjN+X
4B69cy/UfQvCM1KI9AsOmRWR6urcg1AkcEgoh3xFT3rHDfPMMhvrnuzBua3kpABn
YeE8WYF4/bG+pMuouV4dkuibMjOY5Xwmgne3EoR96jHmlhislPwW8kmVypV98XE5
m4MSaiV55jdatPzuCM+cBDchKOS0txqjosH++qpFj9M0sC4HbC9r7/jsTOFmZBgf
pYfUJqkfiHWpc3l8rM99j70NWVF9Zq3W/t45Pqr5JmO8nOhfUUKwF9EwKqlplPN/
zgmw0RkUyectbhpG8V0uBFTni6rLfct4UYaNVkncXB1+cI+LkME41CYy6fCE4v4G
ZpMk+Br24Qg3iOvO3vkh8AtLcT4RKMpOMAwjxxfTnglwIsVsrqFuQ+bvRtADrsDz
w7ci/byuvRb6YLhGG5Arpsf7a1KWpwq7mFY8s+T9phPQHQhh2l751EqS0Mx10ssK
hqQUsMuebbvwdt05ACDBa7VKbZzfylFN1GZt8YsVUeDQWVK8CQRY55aDIxblp516
4BS9o+T61QOIYdtqEYtgUreaQCWpQ+7T0zWUJyFA5uyks2iwh2/FCYDu1fHzdEtS
PKt5plTmOZHw9ZCa8N1fpXxfYOa9iupLQ6MAeeamOokABcjJSlqVyXNx2Lewjolt
zb96cuzJ65vJprA368TO6Ff8Y78jH3ZGgCFU86CqyVNCXSF7kSQO/9Faq7K2sAr0
CAZqhHKYz3I5ySThnHTDZXjuUEDiTwrZ79KVGBU2UaGppS7HgpmTMdo2Mx3XOeEf
m+DkGwVrfWYYzlfjv+EiwbITQDAF07e7SLoqiJ0/YBZGibuVMDSIra8/zwyGgQ+Y
JI5bD5FzsiMfYqWAqCMpxP3rXhIrUJkfTLglJ+cw+7/VBC7QEPtWiceEtMJOivn6
wv0ZAJE62K32xWWv7x3EIEGvsr3mHse40CmJuV5sQuK/A3XsvCNOQ3k5h1LEXRk1
mgku21qKKLtMfBfCYYlqT3cYYTtE0S7Nv/sUu0fGy4HEQQdU6bM8K/8azoYgZlnV
S6FL9zDPud+MU4/j9Xab7wTClchD/7XfQaQgnbYRelOCmXpdPeBDfrmknryw+z3x
Vj2KcyTAf/ud7Eq+MetHVLHOEPDyfmVQHNS4nneVLqTWySsoqz6BPZywPdKC3aT1
XyaLsX8gnZwIwKK7V8EF+cfR8c2FUXEmURsnOJvVmCuGTyJMeYthlWEV0BrnECaG
D6+OgD2r1LTeoQsseCIkcxs2j7ZlsO0Rty6vEROGuhAg6MKMsOkEEbTL10OJ39iV
NvwAQIFaYIVhnJyV3GvTo6Jk/JreCk8e5fj45Yj2/m3xNXI6i/nhkWcD3xFiIqU3
fJ6Vq7YhKGYQNDY0nTpyks099c8ecJ/TEGNfatpACSHF1Atre2SdR8V/S1C31shr
fY29/KuRbAbHv1stMvK9o8aKuTke2VhmAC4fX55nhxVCWdhaA25birdAJSk5C4Cb
rnUQjxZvKc8Gm6Y5C5ykO47MlwSSrGOVqnoS+SkRrtM0F3ahuGEet0qGX1gGuVsc
n6C/Cy6xTRppG7ET5dmlxWL/KugFHJQ7r3DGnh6cse4dGt7cI7cXBp840jgZXP2G
E16kUjzCJKwiAaM4RcIobxg4imdLj/Xa3eGndnBUYeMD5y/N3JFVlk+OAal/9i/r
rb6zl3gwoYDh0VHEa4ChqISauEc7GiX4MNNL5UQlu1gG0byWvE3af4c7+4NUq4dC
vma/m3adYSlw40hFN1lQrER3QBuBfK2rTeUg3HEqs756rHlg3dyuyma6rEduj8qs
F4UE0EGpY7S2MEFiOatJqFSFwSRXL2QFNsL8o/VB+GA5+RnsVeJwvWA3emUscyT3
5DqqmQlsHb9meMySl3cwZDRJSVVrWrbS0TK47FysbFow9bm80nrNAmGkFAv+RY03
2Hw8IzURj9iwmB665I9f20sxMNCtiavoQZrg/6+Qduw7uXQk37YjCuIQ+dstT590
Bck0K/o6fnprPDl8HnFXHZOBZ7QiTd+scwEc/XZBVnXgP+JEYKzSk0LfnUCddoEf
aKSv4zYprZvxBx+bKBfJp7gJoGNvTgDFp+yNk6m78453Q6XlaHiUDaFs55pkfmvn
Zq30A7f24IR9f1uKBMRgqwQRQjPluJekev8X5SKLDqZj3GRZY7IifBax5jRXM15C
PMCF5y8CoQX1US+KyOpTv+bevqLBYeQX8x4cD0rkV7U4z096KNZBWW+h028OoetM
j/5QEwIdjMewPjq1NrpdVeeKurv9t0vLm8ixumyXubxlrllxmcls2Ucw6W4CBi6C
rtqrzhVdMk/jhshajm7k7WPADxOTGpSqR8ge2W2XOTebD8l9j3Pbxy+cMcP2+lv4
NppNN5R/eyBZysv3XMY2NP4lXi2mEYgEhufPxzZT50OmnJvDqK3ntCCOH1hzhMVB
4ofVddPzBbX/KywFqwfkbrWyk1k9f+qY4Um1vtY/VKj5EA1fcElrC8eEHrJmG6/k
9mJeGV0C+G9T73Cbs3HyvIsjGSWBwlCPWpBSLZdApjZ1d9jBUluIL8I757HauWNL
z0WOi/+a9ScSs2oqbInPn1k9KdYeZnrdlLtUSCcyA0CPFoBU433FwVIMpcmHywgt
KiBGbpifLYTtGInlFUTiZHuenwuzupMlpVkdUuUxvrimIqI6UkqcXiGzVegDP0HM
XfZ95DdC3Q6wCRqxSQEiC8hpumrPW6NhdkTeOcMlIaisxhIulLZ6BmED8hFRxIk3
LEPMjR676pyYBSbQ5GRDjn7JNO38FbL7KebP5aQdlvJtDoLZwTzjS8LsbN5WTG2m
Fjso7CFidThXqW9gKhXuzIt+3rM2NR93iAenpU1foPeQs0P3vcDNW6ezsmwmZUrj
3XozUiKABhS8QHO8zBqMHZFHlHMRR0QGmGduV6x8XAREGj9rhNJsvRRdw1DNF+B3
6hGoa7oVKL1YV9+MKnoqUVeFZGmT6/PIXmeG4fUKsg/cOlibL06Ca1GimqWKXMf7
lTP9QB00YWwno6c6T/Spo9PzX6K381lkWYhdbsYsbbjgjamq/LsaDxkBlXjZMwq9
sf0RfxXAQceqesES35xfjRvHfzP+X/KnXfKpIjAgiS/+xSDBKIXaPcSlxC+FdWrZ
kRPE2KrUREduwIK4bJcfebKP6YVqUdPilWCigFtKrcMV9jTOsT6UrQ6kQoo0nN/x
obSGfExibs/HVpoq/83u5R6jenc6+1KylAywbdCccceRJOWz5Sn1L+TAi4C7hCJQ
+lDapaSTqYlvnvlbEM3UhuCC7PPcMk6AXbTIASqC+kGQVUis3+lpC5zIcMOd1qcB
CGD3r0MPQyXUCND+eWxILIYVhlUAVLr+7ieSG+gcwBv25f61Ae6Q0hT99AewY24x
Ge7rk0uICmNwXm1GG85c/4q4kLXUDoj7atsYuD/b9F1Z0dPRUeCOhTw4Je8ZSKaz
ApAsdey9pC4EPETf+SCvEIcibQuff9VWxBou5OlRobu7LkRmRx/jarmk2IRzTUfx
Qqq3WU62uDNdXRHnUDZI5qnEBDwA+at0uaBL1LOUBDyKcZa95hj5nmnEWV9dw1na
CnAJOtHMpCLHY85mcSjo7MuljfzUwpTgzPdhMCG1pZcrmEvFNV8zjcrrSMjELbcR
x/F9TzAGV1FQHoAzo/z0BxSjfNTr349R6ytVfS5fqUWXIN6rgtd72nf2eTHMOEm0
2DoXTCHKhAvyXpRCaXW4zvQ1NjsiKISz1vwSqBWIGetQ2g5tk2HXve0QuVJqocqN
2sBMMvHxqvCWNV5aO4+sClVmsWyqb09nf6+Hz4gomar4DDZpSXP8SeDCa0N3bkmx
kZlg15Lm0DTzCcOIXOxC8iqfglNB5d/m0Ob/5YZfbKzrpakreyUGcI1QZIzoRIJR
FiS0gsemCYIXRNMoMeLbzoaJV44oZFS1V8e/+/S1y/nttha7QcrODFotQuxFiLdw
TdILJ51yBDF0ckWBx8/EBGLSwqaNeY+gkvHbmDDHqpOW9d98gWdSICpYrQc4uwXe
aXrCnecH+N7md2XoA+Ni6fCts+4p7/C4okTkXO6W911q3FzkCVi08jRKq66lof89
gXC8ldTaVIQ1Vz4F/iXdcu+Fh6dIAaMYLM+N8GELeix0+X7xCygGXRfpcCPvFWf9
UKKUAYxX9CRfnZVQQJVGdWI7aQqGqWremrQBcKhMf4Thj2qE5H/R2Un4Oawx2A5I
2z187KSbF9k69TgTQ6+4c1L4CCu2Azaacy257pekAXMAylg66gINu11x+4bjW3M9
3wiLyYWAA4Iojq3yfJ+KzcYBLPlDzR3vbn9j3nc6NEh729E3i3SBSYHWOndX8fTH
9ovnQxi9JzYQt29CWf4kVLguuWlFvWpr7Sw5G4dhOwlEHl8/3B7CQjrtMSAzlJQd
Nf/MVeeyK692BJX5XmV5f28uP1vbayoQQa9uOgbpssVKEpSpb6ccquDPJ0M3QYFz
aeusfWr1mNizfRcIIrVZWLrQBBGi9jTQ/SwK9rKqJ7/g2x2KQ/GrFiwFEUpyRw8M
EA8Iq80arv092APVd5RHGPnCy5Q5xcMETM98c9QCjSWAX93cryTv+guGssGPuqq8
WIn2olfK0iaZN4HdQJ2aY+JdHeA8UMyfRUl3k0J5fXNfnAKYJbp8taEUVSofmAPz
zNrVpUr9fBBQhi66SdDUuWZYGO7oJCp7lQlAuvnVTTzZjcez5SgeVUjQMa+oDFtU
qTgMa5JosZKEpOc0pClTW02/KHv0Kny3uwnVUIvlUA/1vCkrjyZbajmHOUO4szVY
21Y9dRxeFpKq4S/6+X3wV/8hB7pAjXbk2KACWPOzw3lMguL29zHvvGsGTOMKPQ26
WR+KF9rI+5zrV0MQnDjDAy/DUp/sys19DZTaI+aezyieuCTLYAUw+Ke2j/TbOlY+
gAUB7P8+IJIqXNIGVEH+hykwLf9vLXpbSkhlG+3k1JtTgloSCAyoQosjUCbNg/9G
aYdmZW3xNeMA6FHL68cA1510n5L623+VhjrWBWEAczSt81ATOtKCF01tJxjYoRFU
uMyjSyF0Xar5hc3AITnrI5hpmScxqY0wdDNbP2ILIVRBbBb9TBqwKzjzbkk57sAZ
LJPlkztv9dZMM/1Z5bFxSnkwNRIe+bOi9g21RIiIFnefV1JmDO/TtZQTbtDmhZzF
TuJRAWzpyQGE+0gPTVmBbkX8QmmEpyHlocRvEC6OBis61A8+flFLBWricz2RdV5K
dytMOaNPTiElTSBqXk2mGBjDNevuRbI6sEJ34fSK9tWWfaIp9tAKP3gT8OH82l1B
uR4UeQ+cYldsty4EHg5s/ZZkJuNHs27gugc5jEPArKPe1XZUrC/dGSVNHgS1tpEC
eaqprk7QLS/MWoCgnScfQEmb5XE55V4KwxrUDJY3FYpamfPhrQow17f+WFcPTYQh
bWeOsl/7RQb9SjsSP6g9kN+SknqoAcV1H4i2Xr7IGavg9I6sANQp2GQm03XlIZl7
NVFkSJJ6UBLDRDn1GrQTfpXWl/crw/spG0/gJT97THQFzjjHUxxWLgsuo83MsRU6
HZsEf9aWQ6D85vRfH0s1NLF9PvuWux3CJxcina5XVPlrXqlb9Jdg/PL50hAzLTm4
j5QmyDVcNoif9oXU4R+7V3kC7O1fpTXtSlRweRIIjUqbfhAlxuA057wrh6mI8DFF
/UjbfMy6WQUrjz288CQLJ7BGZkecU48hHPDvzPFTLJN8Lhnxbu7FpuI3HGBl3XZN
P/7v5NQY+/zd4j1ShWvuGhI/9WSElleGv9ezwOquY49qdFmiJGAJkFQ01nsfPpx+
iSoy5WL6unGaHGoU5HCaj1YZtRO7EEavSRf4BDYEXYE8oWB0bgPcT+ZAgGPQsrIB
CNKqzQsRnMJtDt9Dk1q+zAJnEKxByXxnPDKlaIKk5QwYOAIRABmatUgHDBLwoyET
8OdrBnpoc4IxoTPUSgKyhB81BkrowQk28BxSORVqDws9NlufntNhwAPKr7Hi63oy
mNCImNn89lDK9Z9ISPOSE8ZUa7NEzJbw24VhdnVjDXgwbpiznPm8DgdcqOdkCbZt
fR/gJTCTBz5m2dL568XioZMJuy480RjU8lyTlWLMdACvQiy+HKoqxT6s0E01QShF
48YkwWqcDtwjQrRSLjxDSyLJVaF9sfReROTY+/XPCik/0YDLI1Wv9HP1Ld9KFJTq
xpB/RwTfxPnG4Uxwl9qVeB7l9s4U77UwMyzIZeq0D13ONIO3DIxre/HBRO/NPiWo
GY2OAZbP3a1+ELLFzddyXIOzhm1w8qyVGuDDO4f0zyfseBjIWXnFxob+T/cuW78t
HBJyDs/RrE7ErQ6R60s7gCsYj503uonF2dC2BRGISY9J0D+HFBezB1NUcFwrkgQc
ZxdB77yUAAo2YuH+V6M+nj9ZIbU6J48NmI4C4M1s/w1ivgEv8GDQx+SxZu6g1GJy
6/cKZMNBlcMqJnf6Dzo9y9LbL6NUi3y+gmoGQG1Cvi7jcMQph66JPwTtCeIuz1DC
U4fCeCj5jafaboMt91990JEzqw2nRssFLbpThPVNEPzAlQN9fF6ZYKcd7NMqPLs4
lADEtUbtASizJdtTNbLp6BvS3vw/gE30ZWf+0bJDDkePZL4MQ+rQluidy2nO8jLZ
xWII1lYGyBB7zZsrTcIDvJJvR/+MSVbho/AZaZeTKp1KguCtlN6ZQE+sVHSl+T6A
9F0QXB4DUjiBiwa23ASoCtKuDmg+kCOv+hpeltIq+/V2DF3yzOXdf7jgG0kdpXcJ
81Y0ENs6lES91M3cwwpSEL/Voiscx6bvyLQfhJ9dkrZXB4ZghN03JTrf1ROpEHgr
MJqoH8PKSOtxgvyxmsasd6doxLKz0s8qaIZHHmnCjfuMds/BX4V+bgSOsRq849yi
wA2RYE3OlMFmQ3rMYEuQSyWxeJcmkR1P1q+rgaZyrcGuidFuf5S+Z2rnHXdykRKj
tYKgUyIXocntX457jp5ce/YlFFQB8Jri13dqsXjQLIsU4tRVHTz/XbGEKQHpujXD
i01kI98hV6AB0neHYWqZ1jVHxg/Cuu/TDDXQohCYSH1lk2ouEgAWRoPhade4ArlD
LsNNNbtpBvPyMp8T7M6AJG1P1nB/OTfaW+p0p1jKMBdV6k3w5B8feKum8194JnRX
+nbdzUEfZ6uXuDiGSyt58qqDgxcIzrjCtFfB0UAOKquE+GMAgje4DLigXuGAy2Bn
xxg5Z+Zh53/iLkWbLCioGXhWt+GUJ7js+pS0eqrgoNNF+wh+wMVrw0yCFFI6CwwQ
pGdSf7Ikb//Rvnq6MQHvtogxzhXbBXdWnXq0VtJuN9kQAqaIRXNMB/bSKRcqrZJ7
ZI2lTXfiydXNZEjA1ImxEGyTMoReVdnZbW7YVoMySi1X7Rn2+8UnC3gCU3qXLPFS
aPU3nU1juuEUSyTZydU6JBoRjmiIM+XA3HHXuWrn8oT4OLTdJuyP2S/Tv72nzgof
uxcOnwepa/1rZ1p1/sxbBOsg9JOeyb+aTcq9XlOrhIb3aEYdMQq7s4K7m0p91VEY
NJqDKX3iLzJvrI4NraAm/MdUqmNLwKxy8KrkuxzNI/QtP3f2xmE3V0OWKR0f7kmS
tdRYZ6Ymc3pBB1dEo3WiGxP4ImhNjQG21M3fw9TKza5v+PYbKTRSxkoK5nXtwVSF
mLkndHUlal9XD1xTwxqp4eY/rcibrB81f6bNd53FVx3cs2wByny6hHWcHqvsJZw4
zCps3nqJ7fn0vaUqO1k4R+nh/AJoWumV/9SDUMcyLWyNlBdZlrylTK/dOmtOG41x
RCtiuimF08LZWmjLjGrEs05r0/DextTQSgtrGY5M/F+KLICsZsX0WRni7VSIHrJs
08/ocSbt7yhNb/ZTmZHyS3NF/0eJZEyHvnKeF9VcQ8c+fhZ6NPE92AiotKSt+4Qy
GdXzCWickKfPtvOrwGfmgZtTMTcJY6ic7BB0gDhmJ8oFJb449jXbRuSNFUMlzWgI
QLcu8mnGxDRAENbfV42MZ2wpXXXIkg3xv0S7to8tQuksJncKlSKWpRyNtqcPqRkA
4OpxryQj2Ls8CPGGTaT3mZwiTN/6KWsP6WEOl8+boQVKl4Br8cWGTvY8r5lVYZOT
KIGUM7YaYLlK7Em95+0ZKIf8V4JY5UsrUCPmsa9G2YXqB/oWVyJ2Ny95k9uem4sN
hZQxt6HVypH9/4TWu4/ijMD0x1yLo/sUcYqm/n7whxSvT4VFwri75brFeXjXN66L
5NVmkkpkLa7sT6CPWdTmbrIcImN9wvbiCVoA32DUur/VyKiQjSqXGs/Ibsjcyb52
Z8BeVNd24ezqhzA9FHXk/DWNi0xdR2m5HQk/X4oQ36rxMs58AGdTU9rSnVDY7GWP
W9quEFWpoaEwFuMXniCgCYdkxvp65uUlHlV8SSV27owEdzI5BGoZe8xTIr96g8gE
+qeJU5SsUKUy5eRjzsDrM3cn7TuaaFSYxowyd41INFCT0qN7TIV92I3oIrUy9N7N
/eg2uQlO0RDGOezdWUfTKZv76WRGOsFD0oPjOsKcIDh8GshoAoIuE0y5dOWGyV9i
YIGIBFxu3nxTWENGGFzuTWuhkUIZYSmVxxcORPSpIxxa8BW/IEutF0WlYbcNBegu
kOcifaNp9bz4cbF9LQmd6emmqM0BWpUveNFfwZ6jZPHjZYPIGZwIWqyCu6lVfqlp
QwoSPQzvEgx7Nn3tgLZOMiogbfDiLCwYNkd4Q5LmBXDMEGVvUAUGtN8SyjSnTo/I
8QkKtm9ky3/GgxfLtOkLlt1ShhjjHUyyj00CYzx39nNz3pZlVV2c7CsUunfeErkq
FD/+yt1OVEluCUt6wjDcPp89drB0yqFqTMLX8npVa+tx5VSb1xk9pZ4jCkdRAlbB
dAvLwvnHaTAb1Z8bIEKVu3qJWG/OOIYGPa4eVXThRHuzLOi68jW5W1+keGKEW8nu
BL1eSBO28hZ5+73QmG8Hc/1JAl4qgZPf+0++kSBQIr5F06odI12j/JIEdy96uwd2
MGp9iGf/yKpDPuxo3id92wBLzlaApp2kWOkaoKuit64UIt2kpsYxxNnDlPjq60Yy
NXRd+gauth8GvRb7/UHonCChgcVH6SZci7FQUFjHC+1tJGXkvhGys/be8ZguTmOB
ifNN7MBU8jG7aCQbT75ulpnhqIlRgGe2Y8J7Fv7Y4ISudwaBXKyeDqUa5Vd0EENe
Bvlmy3Q2OC4kHw02tA00H/8P8znhbLUtodWRpNM840Vhvgub6OnmBf7COJZfaS4j
XmHo+vJ3fZ3EM03RtbGurprVxXtw6WsGmNyGruja7y9C34/XSLZPrlJmmJUKDC0y
vpy+i/yl4K38x2uTsrQFpOA4Y/QoKky1hBjUVS2q4YPhLgOqK0gTAcDAXXSyVpUQ
pASxnfFSMRgh4XueL2r6LDMg3RnnCwoXAVFFXXoAXqVrXW1iCcjptJjjM4oR74mh
Iz7N+mhUwsn26hsVNoKNT4pUOuIAr887v3LoiskoYct4FQyEFoWjTKjCpzTwvEJh
Gc2ZH1MioKCNh+lG4MMCPkvWw6m2PHAjszXC6U0scj5A6b6v+JDdNhxad5W4pFTn
X15Kov+HiajDFgOoskPS+WPZ8OJm5Nwx+6VpW6fp7ANNYAaPQPmgfKjJLmcr78JJ
QGO2Ewd21R0LCxybaA1/4AgAU2UHm5u6uKRRXPVcN1zhhdHYywAlwIeEkm7sgnoL
cgXKrPF/KEQBzwzjTxrgYynK1da4cvrcqDHXRSMyneEMRCGLSyS6+oWUoNIem7ZP
M3/T4sLCV576G9cBN0utq2E5/ds5EtxRHKr1qFLLlIFSnMQsmxW2wwBSgtseW8bh
tSlapSvGh4WILS4jG3POmOKlrKwm1dnAS+N0cFeJiff0FLg1x0VeP6HQ04oNzW1S
L16jwB6hhnaWrawmtPvuCHBjLE3WpWbcb5G3iiIll9Tsii7ikopJ5r6/V6UjcalH
gTYAqCAlWho2/WW6x9wNlZrxoG3BXmevlOLOEeUXOdGRR2/zmf7mMOpBfSupwahs
YSTu3kkpurX53iOXltfhTu/ip3l9Ar9MOtWUji64VnUQSmEq3baxXPrOs8dmeiU9
0/CLFYCtvdrr5Oa7jLdWWF6bbXttC0rUUpMmzevo32HNfFSU3NUTHATobZhBGQgZ
PixkskCEIBPNjZzQg8IYvu2FyjFzM6dczmBJRUJvqXMQXT7iOcVrghf5zPvXgyLA
htZfNS5wyfnyMFA8WM89aIi3nH7LtmjKaRMtzWwjZbx4u2iSRZWHfhO1MNrRl09f
Ap6y/2QG2eNV8KpwtV85DoRx5+oqWIa6wcMtDTSNFRSoBFgXPd2ROHjTml30I4cH
A+MLnMeG7TRVS0+WuWlqiMK2gosOkjhTWpS+xVriG7+4w5ZTkEGIhMpmKEVXLP5d
5WNGyEy7spNZ2EVEW3eQXWJgt1rWCb+GztyRqz3pkBi4Cgp9ZAmgVyAn+I4yHRFI
s21uGYUGs0+jkTKjiP9LIi8RIuUIUM3qh2Tayjppfb4WxUFGF+efoxfK0pKpRPnJ
ApML8O+uI7rc5+vUQWG/5Pez9yiGDgxI3ml7bWyu67dGXH82HY0xqET/EnxqPdXV
/asvV/Tdn5+2S/6WCqPtfxJt6grwI60QAvxB5ifj99vrUoWiu79mxkh3+TNX2g7M
MVDZZB2c8nQjhkyyi0+AgqO0R6vcs1W7kSaPj8JyYM3wIg9nFbOG5ZXhalFGaMYZ
x/K9MY2luPh1plYVFiPPCrR2A8Sie44d3mhUOC9QUtXgHK67Vl92Jid7/all62Tf
vQTNP+8SCiYa/z/yld5wFc1qKjCHA7doeiGXa06AFzC/Mc/cseyL9c/3tiqYlw4w
Zh7FDqb5hJ0BXBRIKFUKwyepme28L4al5LaporKAzCmuphPOf8XaUEtnO+Iv7TOe
ENJFIuqBJyNhZtzlCUhaKDso85tcXBQfqsfKI5eBVs4FrxTgPKHIRp/zv5XnRowy
zBoPSTfvdpUq1su0pcwMVY3oTPdwIA9Hs/Zs4wMgiA/wK/vs4xcPyPI4TFxtzZCz
3ogZtDy4GXAhWtW9AnJVIgFuxy1GiPWVB2neUw5kL34xgt6h9cLhmC+dr+f40Gx8
0+D5Mw0HYlENy31lq5rWEWwykNUoCjgGfmp1VjtywV0QQT8s+FTrt0333nY9kEh6
V6oBqDXEGr/ufJIBT14CfAhlnDSBIjuoOtQC8GPzrP3gWX3VJU6PBDuOGq38Rae5
Mc1+8mTZ3QM4UdDwiNjcxvXtd0WYxg8py56zcpEcavt3ZJvjRcFCBHkoB2FvzuZI
ikeud4PZ1lN6Z0ZfGtRJgv7vlcVezgNzj6RBUgv7E7MPz1vr5HldYcUX3TxHKqhN
ym4aruNnXiGldvMiNU5c0Emv2i38ARJ6wrsZOlMYckEgWGPFCyBxLz8I7xHrjZf5
8ijDtxYxG6CVroJqkWKpBEgLM1k5eMSSy/+mOn4szwrJB20sj3HHK25+JfNgwSTr
gZNRKRfR7DqmMZlJ9LlHJltXwBgKIOOdeuiKTY2mQB1zzN03aiQRyzT1bB6vNaYC
Eo/khhIGRMOtcyr0jZemd4tSen7f9zMBphag4+Hn7V0ZQXYK+UBZIR7l8d9EpT1S
vABQeXQIqfs28/T52fd8SJUdEvHqoUISP2nAmoLNLipuQLfIOOFS0Cm++24ybzSF
ZVeqDoxANlWjRvergDBIUly5/IWWS7wBYhbCAY2DTXs6IIsseealfryEF2l19DXa
RQi8X/nVqEgOF0kwHoDcwSv7D9cGRpktoRWU+Mc1rgODL8ERuYwTpglhisoDNRWI
RlqkImYt0HtCNKV9S1Vq4ektNEMbS5574ZzGCj51MrEiYnswVilrUaV3JPQpPlWG
idZb1/8/9+4q5gmYoyBuZw8cql95pJ8gp+uJ2gg375QMUP8dA90IbplgdR3HDtnr
EjQFC3acHfPIOjWwxb5KtIxpRACYOyBiaJ+c637jTn7U3fc/VRC4f3MibTaZh/8g
0An1cOAD+lg40RcLH34m7PG1v71viHBYI505bdjcnTpHxDKQpMCLmjNlB1XwktUq
aX69Hepuh6QXnEKOXns5goMjdytR4hEIl/wm9E1z6M5jvCF3cTlVf/PuGlvENNnD
QCHIrRxpHmIo1z8Ms2YHTYoS9fYx6jDGd5oXtp1FxAUFik51m3DuiXjbegq8QGYe
lyhrGdmnMGTVmt77l2JvVHZSjDQsrote6LrV5wHp+PZc4RoppYUaI7QqXwRv0I/1
GqHn9Zb6bdl+g3f0C22epKYHQVSXIAsJd+oRZpMoIYczW0sJo8MrHXkjEiGZMtwa
NKkPPmwT6D5NPQLJmgPuJZt5AS8lhmxNpXjo+tWsxEgQ9FvmLXP9stOrSz+GVhbn
CUeJpHENqkls85TASOpliiAyVoS/4AkS3BukKoe1qwG9+jenCw2lCme2phojjm8e
IXX/eC8/Qv552N998RaUp8WJ+77fysegM8kvg8MmNZooA6mr+tDTVXeYJ7hGIUg4
7IoXTVktixmvqe9+us7F+B5Lm916Mdjl25YIgPedMYPhaymCa/0aigf4n+mZv5+b
MV0gL+lVsVdGLs/vBjArQoEzXA7xjY9/518KsSwIQNbCqOPVzqhIO6xX6pIFSGsV
LN4ykRlmzspuDXdyEzboIt6IkWvkpQH9EQMezEmq6T8TLoOXlzDlzYCtCeihWJJd
MkDU15UjH5kqLwruA/pCXjHE80adcRXf9Vi6Sb09OdL9ua6Lt0Cu3NkBDj5pu7Xn
w9uAj53tdVcuArLfsBrNgqJd5cMfL+4xPAVNyTOKuwBfIomNo8GKHdLlFakG3I8N
P5B+PkWmOKqMaIJwoSM1E4YRgcvTe7UvVU6bjPhZxGLXsCHbETE03QfE785n5fdO
GHQlTx7Xbh01llCQDbhnSimt3H4ixNJh+83SXRIWlQily2UhK8g2mjX1kQIBKroz
/nzO6kYhF8R9RD16+SAMiGAI0yEw+B9r7NDWkIC6G3VLIfkOVUNFfZ7KTnB1ZXEZ
bk7Rj32Zd1xazEQZiHu5mVaURzp+9vWsqY9c9HvM+PmSjOcrol2KuUNDG0tbbvbX
Xm8IxTnW+rTbJBjnXlpJdMKQ/sLbiegYmWiBRqGpjI3QeRJR0DEMca07zEHgqQVj
h7w6a6Ds+G8RgHvuhQe1+DOJD3w8XMhGDBQq4oLBwGHttVD29p6xsDTMhZh879OU
lPAifNGRrBQSlxfQUUFIo8to/awMXn+dKgZGCVKHskvZR4NMnZ6VVRfFElU3upI9
U57LzxZyvgt1UfrayO/1scgQzgLLLjxCaUXlDkO1TWHUHCeKJf6IsB3FSWwF6Jgq
XgFGy8FanvST7PKMMce6BdIKIrooKH7ZmdmSPn7cL7njwOXZO6feiUh/Qfw4SoqQ
V+uhvA+UbF6Qcbk4LBFeoiJsiRsoZeqUykqq6NznDAKPq0c2j9syqiHiQyX73SKB
X/KNP6wbTwlGwfXmyx3kaUlpuEFFlDgf8pV+1kvPfJwroSigwJsdcKvpSLWq9oaI
rkwrboSHk+HfktWCdru7eOy3t6AZmNaiMvo8PlwHLYZriy9naTtzkj8ayjWkAkc6
6/03muMABvlXSVpAyK8eE+/0LK42vcFDUekbjigN1/sybVy3aQuvXdndSoegljR+
PWh2e7XUczx0wTysoDHX+txIvd3dVje60Jft5CwVQWYcBM0BjarOxfaXZ9TMer2G
DcgsjTvEDtOXOGcVOMCVhyl/cHt/BSytOWP5o+SlzmjCnCblRVoieItdDVPjLg/q
AmQjKOjFvgjGaa0yzPNJiqgGPMUXbBbATtrc04d1fzIqW9L7zLCAwzwQNebMufs0
UNOfiB2anXhOyrf4Kf1qtxStAUHKCO/dhf/lq+XefLzL6wQkspcW+LfzOKVzUUpZ
D+B5NQla08BKjt2pjOzOcddTCmZWHuK2QDSzs5QRY/2uQ1nT+LH0LdFLI3M7kaEZ
82RhvNb6zaRG2kDQ55REIsr3Lbtp3zLUodmbZDl/ZuRIoooiJEo4b92osdUuTuhT
bHa0anftzP/JHQNxbIz/TftjjDe9jbBr8LU01KpXEcBlP5tgUor2Mtp9LcuoblEi
UUzG+2aJ252/vxPmGDsUVu9bYke4iDqcOldLzokDjtsI3W6eIciGiKSzPyC02eBj
dRiDbvEnuJoqEomzH54/0jsJBTGKDT28c2Za1x/7fFAmZv5SSuWolZEJgaQHjluF
RevRHBelfOFKv6zr3+4svWtYv757l25+7GThkABnZIvkv1zjnjrrPSBVXoi7WmGI
89yl8PggnW+9GcA9uEJfiArCs0/dipKmTom51qUCzWPHHWzecXztcY2MKeva72Ra
Lakq5R6ckp7GJ40XCZg0W67U+OAeuYNWOiafi0noL9EZs1U5cuyQuf2Qp5pMO7lX
tdTaAxgTy2WoLVV4kETXzg5y6h41kRrVjeNeuFI+3vfbGEZT/flL/YOF4l+KC19C
NAQoFHbc+NBTjRxOPaCSyh6qGC/HYsBilPSmTDyBiK/KhIzjVdubEevJLCFMP64p
OcP7LgraxmeBAtAyuJ2XfMY0gnD+Ga8UHM6iFSD6eN5jIo/KotoZXssdt4erCMbm
IenfG7ue4pQzxujwWpxcQgLFAHqUUiD9xNs0+CtLDPOQ1iMREahZat51jyh8QVo3
/E8CzmOeJ+5f7SeiGJOZHBx3wewymSOzxFlcUxeM3TVgD5jKHdsGphTdAbeoJrxH
CNc/CcHtDxvx1u/umBe0Tk7Myj7J/nfllBKZdq0rl2nudqJXXlv3uncDbnMS2wrg
81Bt/tq97abdkoKrbfkm6usm7KjnNtfzs2v9/lXAk5NBjzCZVjKL5aB29aXwi+iu
6/Pdz6A8wpUY1xFw6UxKhSaCSv3l8bBKl901Oa7zc60SS75AwxfForF4nRgAoFdk
efv+XkG4fXGgDOf+45Op8R8ob5MNf8oN/xHr6NywbFH6NbxT8U/84CTAQa7ry/Yv
x1CBJ4O4+2NFQPi0NQgkvd1vE8Gj2vXimiOv1FkRwNIEHaQbbaR0fqP9KgC9RIFL
HLloOJgvH81gA49a55kA6a3rqND9x2nXFY87W6BB/99ROqUHOe7QRrcV8Th+ogPF
3GP+NlVmjnWqH4uq1s4JbeIWRJRvSp+/yOsL12PYCtJTgSj1BeLNVGwsxZO04ezj
81+gNwD6aeEF3kWc6yJvei1U2FE5fYnHIKCIzvklisque9N5D+ouCnR/hb2Ohs4N
jsMYpXWZtQIeSo2qDV3cKacdekFZkd9NpefDieY3j6YIGboWvdFr3Zb0HfUpwWH9
3Mh2/q+DPNXOnxNJphYHU633Ie2LmOd8N1Jn+4beSm47mcC9Q8bQVHrLG3b2PNku
1J3w0cvmhEyEsH0rvoMEG0Mv6sela01UGKqTVwIM6aIfx5Ps1PKeweoenev2YLWh
5xGTgYE46epz4Fc1L0PzFTB9KxId1G+46dOWReo+cHaR6bZNptTVYJLNKM2ed60O
iyR/8CvP1RhwLpj/79TUCfZ8vs8XXQeMvAqvealRTUfHl6lXZGJxYRoIeVQWW3MK
LxU4tXqrZSBp+WYI6jEfOYgImiUIOlWpnvyZ2eRyYCM5+0fM5Kj3DAavfSJQtsu2
YRNzJrxLqkzzzWTld6rlaafDUb1e5FLVSnHHvJDWSK4oRgHRF3Y4mrKJYGRjNNa2
zWsnc6dpOZ1ByWqU2WiCtt8rkPbrVN7OEd0Qz8WxNGyPD79qVXTDe2Se152+I1hu
PkBTdQaH0DMcj6zFI8TVZW4/wBnfd/ki4SluYYGm0pf658dszesuw8f6fPY7loe5
l5o/v+H0t7FtgqCWLNeroy4f/tzT0d0qdjlgiRKPF+i72Gzr3hQAFerzWePtVXGe
66ftivtGn9HrsG8xy2FMUzT9MOEkLt5JaQiyVv1BH/+i+fwCmiCXDHw2DcqMAURF
CMyueck7n6xdpXf6ylpd9azlGtaHtay+SPvU09U3dehX19ERN/B2BFgS28HHCj1Z
I+8J/KcMai9R46yBQWSomrwSPykkPu94u+IvJTU4A/+pkAJPGR7H1TkAKpVKnmx3
GbMjvgXZn+vGH9OCk3YP3HFayHUSx8wd3yVNECky+KXZ1LqR9OBZdyqLsuJwuj44
p9ie9gujlyfFi5K42Cxp5vPKP6VzreqYdYwcsc3mSDplpGxyVUnVpzvq/pvfuirW
zqDiVu1BPB6TqAs9+SsoO2pNnivhQ2FNq/r7QuOXDo+nRxP819oa7DjnEmMtAO7w
X/t7ODy2iyzN5Du6t95TjHGcpxoXRqSfd2p+69sQsyWhNBhhTnB9yi9vmJ4hS2eK
PtzC69vXC3YDRfVXI3ut3J3K7kYlCCWIFZ7Scj/xRWhD0YcgOb7+JWaZIq85XgLT
pWetSqA4H1hpNu9A08laD5d1gOQSA0JNsf8Qlri/J2bYp38H2j8ywgrzUmIpAg9G
w4Dz+Iv60iOlEX0kShuQZ/buAC3zHRM1uqwoKfJnCoib8MGXvHGE7uFkZFbLL0ak
W9gvFlTk3BSvuny623GIJxTEFa9K4jFplUlEUbEgEtsbycMEV/j0KEXReQpgP0uh
wgBlxt0o+yH1DdqERrMIzaxES4ilKeYsplDelIOgaW15fkcw1kDnq0Dq+zZ92usE
2Nc2QBwcnUUXyYg10a1Cmv+T5RWALojs8MNt5g4XgdIloWaSogtRgTFxplykJsrJ
QtqgykcaX9T7rWJ2kKx6A9f+9BYQ+kIJsVp7XCXrbyJnq+Kd5k0oiS/lUGrlgtSZ
puGCzVnIoce7aDvN5ujaGh6VL225wiRhGwvwxNIfhO2aJvOHguxxnqc1eNSm/t1B
hbZn/J+idDDuGYIymbpW/9Ka2xPOxO9Z5eWZB7qBrI04Iub1VernFdeO6K6+Myr+
bU70OZgAg1WI782PFkuJuNolRpc9NpEFc925VFLg+mqMsMcCqlWSkjupLC49NoNo
XaFOAZ5aKDgC3bR+OC59FFEuQowrRHg+5zrWHZX0FWRqXfoehRpXVCZUB6iV8Dj0
YfglQM1AUL0WJ/0U+ywMx0RLcd/0fvWEmC7crVIrMmIvD+14aHc/uNrfdYN6brjq
6MvmU4Gz7nCb1Absxf0RWLQWElNi2jTVbGED+277hZReQ1XuBtnOHpnW5uoHt7AA
CbjbTguYO2MCQY9XzbCBiqT5VT0Iylkty2CDPLIeILRp2uzNGlSI0/FjOGpbhcad
YlUn+hTjt0WQkAiGP1xJZEgLYKbj0FyP6Fbbe6zqvs+UFCa/hZIRIsVtP9YhR8Cg
gCVkz4cv8h7RYIfpQJMVnfo5kYwvgZdOupeEXGcbhI1M0kBH8AqY+rOiCCq5K4hZ
ZXmjdNamO/T5IiMBScFdMdnnXgZb8gB47KcPv1JdRTG/mD7TOnvCOD27HNrE5FV6
qENc0ZTRzhDq7JEIkodUt/RKxCVq7DXzJ3MnJTtnwhP4UqjdyvP/QikWO9/k1qsy
iaZFd5JobjSgJau+WhduF0NWBxAwatMc/OIwLhsYd6Bc8VqYTCHea8yGC58QCcOR
/VIFdZE6/fsldoMUVQVNE1SG/27w093RKK4wFdgz3EMKjB1bqB2x4tfCwakVA1Kn
+eW4l56c8l6V4bwmWBpnqTxhd+K6fcPcBnAxEgsNkQDH4fCZCCuR7K76Ad7/aXFP
LLSKMq/5RHc+Mcb0Cg2jldDuSIBOhrTv9RCwg8cJmj1cVfXex0LA1RSed5W+0fTf
ZRVMBp2CsCQ6UCvsneKxPDmlRZXMJSPqok3+MmXo7mhgwLq4D2ypSJJJ7AZlKT6k
nsGXSoi77eqKi47YWh23/rCyGWSPDQBlCB6Mkh3TwRgJM0OUSxvhoccwboDKQlpy
UqWIj6rRIgZ32CVNrKs8RvVN2D45aCHxKxuCNKShMPLL3deg2YfrNjalg/tAHGDF
GIfzw0VMk1OEbPj7AhpqdreM2U/u3UmXvAEBShiQETaF437WDBx+mjxjHURcwLBO
VD7xWQTjwe7SijaI7/a5XIgt/PRP9zBVbeQvk1cRrBP0BKTUxgnJNPtsP0Yj8gon
4bdcHynOCm+eZR+5FgHZbiGuPuIxFsSe743cfh8rGpTSSqeFmdl6pDvh8a+ujMH/
edacKTQG1JJ3MFiquvaEuSiWaSI17jxEKbNmFAroaluXlf6ZlBVaGkLRbZmSAzWX
+H2VAreiZay6cxgILaW5J4VDRU8TPudTAnP5IwYb6tFG0HI5kGU1CT3BsEwu//5R
lpYmz88M1aI2gMmJn8NJMRvHVLkAgyUY9rD4aQ+Jb6e9xqbA1ebJ1uu86qiPpBJy
zw454tQq5eW5ckXyY/sLwTx8j2mJ8Z6kPrN3tSBbZUaIVot/FcSV9Bn33BW3hXib
Lkt/R41BmnzP8ECgkjfLbHX02muarX4SPdVjDRF+gSbdWLtMsV8n9SCl95Wz9WBZ
OAZNm65+O/YhXY6BTDWJ5IJyY6rDU+36Ae5i27INgnJckfB/F1GFO4iDZwwZFEmE
N92O2P8/LCztJQb/BBouKMWZlagezbuEJILXBLp3VsX/2fvPZweIddYUrnsGhPcj
HcpMqWhcDvzCpPIwNvGKz+zh9n8WNeYs98KdZUMwLGZAAMLnJtEOQfSpPCD52G36
eyiCQdYR/uKSlvXjfAM8EmiITKYKhABtMa+Xot5c1fZWU8beHWdJi/rSsTMQ2Ixr
BtBo3OivNDeIWJdVzHdJcQFefJ8kcngtHYuXCH0np3BTeZjmqWVtPQGI44IPrMic
ZLjBTGSQAn5Y+v9YCYWBjT10rImuoMFDRvpuEEC1+OENBg/uryCSQvnTKu4xTXNY
3vMqZIq463rj+8tNP5Z6zw+9jHxsgC/omtiy74YQbX9IBOVQZXxnj2w5wXC6gB9W
iRrZODo7a2L+AkeBMbWpbvfbhRccWH23rXAEfO6fKT/QLE5xKHo628cDprWvo25k
ck1MISW7zTT/w4x82NtJvW3WQR8/JOWjP7o+mRcSM535JX3QqNW6ubOabv5j2yCK
H9EXbk2iic97ekh/gF+cbS7o/rKIIuv8k8fxz1exeM05vl+hMfiMwH2Z9YJFqgNc
9ZfcXXi43V+Z8XLBUL5VWDDwoucz0WMYV5WvfmHgc1IkOg9T/TznZstpQuV3qMN0
RdLS/PNwRo+gaTXvCa+GcinyTCs9kq1pvB7K4+wDiOpEmCFiJykxiPxk1x74WZCL
ptvKzRnSSUwZQ+721oUJ9ZLgjaGb6/tL9wGOmo76owXCq3M9O+9o93qkmWwI8xR5
jwh2is09j/4OyxSLMNgrvVzBctWvXZzyo1JVlCROqDO8vN3rZ33m5pVGo6OtBVt8
BpJtiSks0ctjIeADcsB+dHSkiosYQQ9EPdp1o0CXa7NGIiQrxx91OFvjFBIG2xd1
PVFaij6Xmul8KHhhdqyNnQJ8ckrvgJC2tz/5aoOzWyC+s4aU85vgYaMIp2OE384Y
u0WbsQw4Ed65zCki83lRWSdqfRndmcuxcUlV8ChxKispiOxoCoMJlMbd3/QiF8EN
FdvqjZbTUOoxqZ54o2x2E1PQC8Dk9KTDkVrRGfKgtvoU1YKGrCsBYkyIKrKqo3nn
IPysgmlPUJbKqx6XYZSUbMiHuB3jSnQXliYYsjOZQbIVMaABXLUfj8FJW0VaiM3+
WhhHphG4aJNJ/h2fv0zE0sXHoUf/dt0Z4aRXEE73KYkRsY224X5KbRGTCAu5s/AP
0RXbPj3WMdpv321qL5nQFucNv5hFWlllF6DFaOM2FxErD5Dc8GzAbHtD3fz/u/AC
lFXSvOlI3wrf0ITY+8QykWdYLfgkTybYS3sMza2OnZFwmu81SjlHNNBJBjGenWku
LSb3W6eJhXqW2w349ID/ARCe9FJyf8g7eFH7H8cwrBbbNXVRIMKrnWWEYhJTXK0C
RRedqiPAzeaBK+8iBO1S9hLtQR+z+hMH5ZvmqVFvXZ5GTxZroD+/DymbpRbh0mj+
1pvqOgNjYEnIcs2ZMnI+PtJHkS4lu8JVs7a/WNpoNwYwBeGwt6EZbzmlPHmjRSr3
iwDdnZtn4qUA+ocGB1TAO3ACmOMSoYifHyQN76LoEJg6VkTUsfmshpuq79OqEGew
2BC6S+FXlHqaKeec/rAg9xuWYKPF1JaMful7gedJG7L3Grhn84YGdeYQK+HIs4FN
CzfbBi4TD+47cvmsbutOxDA8MfXp4i48gLtxjfHcOsDl4DserzhRl05uuPaYsbMG
YZ2FgXWjTRt3SXY93qgbHhcr+ouxGIUP6ujEyY29y0csUgH2HFrzWc5mXz5s8TCM
GxtoVx6gQB483aP97CssLcscv8JvVqc/ehozGm/CX28Kw8hzoAuPRmnojy0NJpwG
9G1Ux+BPv1WVcGrczFQ4CKydwokegn/W+4WyNT+ejCrmtAbhjjshV4Gc/KbJgF4V
tV2nz5EhYguwmXM4Fv26AGHIgTcmAQebrRZBwqSMIpqreoMFs0ZC0AT/smfKrhGZ
rglLht0RHeqzr0QSfHssvegnpiG0+LL8T9SJSuY7RHE8K/CZ5Ob5S9TxJT5Ar+KR
ceBapfld4LIbx6iFo64gq2mwRop6J2vuNi/XfY/j3UC0H1RdoZMvvyXxM1a9Dty/
fvWQQV0vsQwTE/WcjGBEcNRLZ+3RGKUCL0WHNAikigRhsk2Nx5dAnL1xwx8GKyvN
7G57WNMPOxkPJdVRq6aJM1DlKIBIsE0yzr6WgFV++WwSmNtxmZ5q78OrWhCSrWmC
/zTAWdTOqiqSdmkTixwAUDRbBhlcZ+sOobi3mTzq1LRqHp0vKVN+/wSxFUaB4wpJ
DCr5YA4UCAg1t7AF86qv26239sJlpGrP/RfgN5t9mbh19QsPb5GEQsA5CB7ZSm4Q
iXYY4J/gAfZxsn5GMnvZafAa2hJcrsW2askfjRPwOskmqIVjiJR/Cut/3ySPMhy7
Jx68v10XjpalkujNPyIambImz3bi3stYI95ngQzZjx0WicJzzx84U24Y+mET1vJC
4DP09SBP6QOPX1utfEPlHqB204xw4pycuVxpn3KDLzbIAXfYQq7A3bMPDHew4WfT
uAbaSZfGwpvF4LDrgCVUoUFwI4KfHsgL8dyWLacebonGHqj5N3qj1Jz1dGd2ZXIb
wlIrPtmQMkHHq+lxisEsIXR0Tv1bPP6RCf4o6ezgBKQCZzZ51owMxS5zMKWkZ7N1
MFEVLoWgAIjvIr8txaa7fSXoJ3ByR+TsXLbXFBXV+GIpm7aVpcwUmmLhj0zvAYfs
Ub5Zfmvd/qnQ6gXk82xthEq6h5wuimu8nGAYiSSKk3KzrDS1Sh18lP+voZr6ODV4
A6+B7ZHHTWHVPixYNIumFkLdwzcauoxmsZurn40Fo60soNoGj0eQJZIOtUUsTYL9
kqCxDPAC3jmXAejTRVw2KSdYPUDK/QAeAbAZn+F3uWfUaEPqH0HBOrdf/jvMeTPy
X0h5oALznMBnTyay0DoUQw+hemhtMn6Qrqd1MI1txTi/eYATxPmbHJuVcoNLNRKe
OEdlCJdm1xUuyXWxba+PHdRQFNr9aouGSaqfxL95ssRFgdvVod0QQlhUre/X14Zs
sVjMQwxL2CAU8yJ/kAMOEc/l/pZBzLRkAa7m7eC369ojomsVEz4LiWHZG7j/yPvT
MPpqMm2T5z3DFX17c5X8X/VXHZ0H0gkNpYAexZIZviEu7CfMRA3ahW2AHPakRqZZ
Z76SrYdd7f2QZgMzfrtr8RyoijRrhvpzmUdUafmeptaKEGxzgLpIEcr8TXcAC+At
WDDO/owgl5kmCMxR9CrEyyqBV7ib3YfEM+S4p/oC7b8qoGjlwT8FjF8VqYGj2xWX
UC5IZuA9bk47l3WZSUDitGcK8DRhIlTIDvvkILYifOox+selqkQ1XJ5UQs8rivgs
C1EneEfOne2ljr1tcqA9TPYELGLpBdG1xcCHwe/CfoQhZD4CbFwdg7rArhC5vWXl
3SapM+SaPBVD1WXJjp3DkzkmHyO8DablLiJyyjXHWXeOrVCkUc6F8+QXaiXYSXjz
8QtDrAJ68t0Zo47eeMUYxyIgeagW1QIduu2iQjnv8UCYyFW6mu4/NoSTbX2/IKdI
rTvD3yKEtgna6G+Xt4FILxH6gkpKRljYI2BfHjwLEWvxOHmZGwsNyQ7/0hDpWNMa
vCaKa/o1AgyegbeTe3JncumrNq1vtTYNz6blrugDknpDUVlnjC1prYC/+taGwDLm
kwFDaEJrl8YDQQBGqk603B8LGzFWFqJ1tw12uLJbtqIVoBHF7ulnX3rMKxhTdGon
GuwkFtLiwwyWHB6yN3qd2h8yBSTWolwEEV8AS0LJ21yeaOhEDap4vlImBV8BzPj2
HZUdJmiZSWagqKHR9gYOIGn9qT8hNXMwO+UJHdhv1LKMgYRIuQfwBQ1EIJP/NftL
/NCc7gw9G7N2d7cS64RhhtXi7xloH95dvzwqJBJzoA2mQejaeS3F2YjJdoIJIZBU
82Q1aCsS6zouEHYCeGcD/6Co6u6brJB0JQ1OWAwcm+J47a/vnWgmGndiXGZbpAmo
k2RafoFgNKkBGDsupHEQQE4EAfD1Dt31VqQ/qdR62rdNTgUS9sEP2Uc62qm/5lzi
y/DHzaeAEkyBFB2ZHx4hnMCgi1aL+CCPnbPB9uLWsLL0IO1VOcozwzJia0DvsqPu
lGVSqLTQW217UNeM+TzxhwFoMyleHg3Dlz7tcRq9H8Zt9tZS3uVb+vu8feHbjR28
Zpbj/yE30pLstsMkV3N11hdmzgl6h0/KE54i+aw+N874QfZLrBPDgskV1kIum6ds
hnLNob9c/IiZJcmVA1c3i4+NP/61egRrW0ie+zW9Jy5oDO3y58oXCHas+PgYlgGB
j593LzwCx8FT18GkqPpch4WMyTXu93BVwdEus0BEpmBCTHYe82Q5qFcpn/ZY3Fzq
kNHcoTW2dPpCDuJNGXmta4jGmvHHzaF6TtbebvWdVg8v+gC5gaYI/Ma12EJ0TGnA
rpUrjpPMDFncFUT0cicVrnXktfQsG6/JRjlB1pdtrlouHIdeSBOY/8bfeJh5fqYc
GpZPr4/tNqdUf9RCxu1ww6YcVm3H8tVKfwV0r8ThYARArEKbKt3LY59NDXg8+6yM
Veh28MO3eBIR9amseRn4pEr/5GCQXmbDtwK2yyZCIAwB50SVIE4wBL3STS18eTD5
UlbG3lCwr3O697EHUPpDs13OeUkS0gKtedO7F24XJttmbvVu5ZxvkinkOtTigNbZ
OdvQpYf7WbvresprecalgjbGLNHWHLsjy4M9UlqGT4Gid8pyu0RMSnraIokNs0nd
H+iTTYQ4osIxEdC0n8bSJQm6utYUzPL5LABGfQf13jB7eFQCvwkEvrWXYBcy7TQ6
Y+9OqnrytVtVJtpaNH9BqLyetjY5GfKg7zqGUW3YZYEBT295Lpg9vYpY/B/pCGJV
L9G2AlT9WQczeCSNnCXrz8yNAQcI4bbo9TNeYWpTlV2KGycxMlXWGigQoGGLZj2a
L0MMceaAaWIklhEjI2e+EF3+cFdLq+P9V/+K34frc4mA1Jga6l5I74xMdD63p/J2
RNKCl3EUWgp959InaB6aQ0I2IJihdNFHcbUrICFUtraP93lIXS0toeCcOHH9Mk9g
D6Z2Wy/5vWPOb3yHRluztnLRxWWYd5N/cp2cRKYwnn0f9805F1c+e3Imvti8MqGs
NtAYBtBWY61h8bt+dahptita28uXiDVltGCh0wfK5lcgEIRCooA70TmG63lYucLq
YluPfw/LTaHRvfw3yI8TNdNsTnGRxDgX9Fr1Yvp7Pa7Y5mpCowwBx86yEW52driX
uN1otWE37ZW99+DgZrJcOF1srmwY6yVwcmyXJtCBhBQQbdCdwcHMUTHWnyU7MXj1
/8Sls+BVedumpySN0I3HGeU9982YLpJ09SBI1fCPTG/afKBj9mM8Rjsc5GjW/z0z
bbHstHU+kDx80VRtnHUq2XEl7lHYSLGnbyCvsNH3MAwk7xop56vi0TukS/ATHVDl
4kaov7t7HNh7SzlBIY5N2y622ZE2rDkSKhyxl7kQPcliCBpZDf5+oIcIOCh4wYV/
yaMkcRPg9w0dNdmG8HTvefTmAFzuIIDJkjEv7+/pcruaiuuEOCzhT+24xo61m5vH
kE4SPEk1tI4gN4RYZh8qmpPPuoX/RGtL+aD88LxnUcwYG8VN+i7rU2tk06yLr+zo
1QXhZDxw+mMJM3xnxaFZvbX2GVW9OoETLZsWO9yKFj3RfgLYf1zdu63f3aiyySWu
n1+rpcEIa1LTtk7towOt36tYP5ySAq7JkTtnfxhY05ZFH71XXHG7EMfs23n5CMh6
UA7qAJCrVQJNuQNlT0KsrfVsdOjId9dK7N+0E0ZAk0pP/a8SMeOnOaURjSZZqya6
3Ce9y/CcCq02lYeWk6c638ZYdLKdZNaYb7E9JDJuMjIYaQ1fGUAkffapAZIXPVl4
sOG9KYFtEBBJ0mzPzo0QI+y6M6Tb6ppIggNJb3pjg8+nvPEeGJsCodmEX9BnfKpx
pQm4543StDuuFq77iLo9tooh5zWYNfPmOIr/7uoFV6kkgg7zF0KEEX8OOKvLx1D6
gQIp8nnxXUmRFTzViYDgB5calYzIIzfphUjwVAQI/wyVKmQnNpSeQPJEPYTgGK0a
R2ZOEALN/4g3tS1YJ3340IGie/BXR/J5NmTyfLCJHEmwwfMpu1OJqXoCgIaZqoNQ
G5widV/wuoy1pwVbpyHRxHDb7rcihLxya9mQarj3voapNw4s9gZlUZn4/EA4eT/C
+92Kdg19R3Z2CETeLmKD4YtHgXrNKpJcBtfeLOFrBlPLdSbT61kuU37YWvToweRf
2q1eKY8y9ojgn2Yelw/lVXdqFmpwDa5+GD9SZRLKieMs4y8ZGhT8KsHJTJ0TMBhc
7Y/8zWzT4pu45ssbCIds/gsfF7jWeGfwGHwLd88B6noYSjroRAnHmnxaqgWBjroE
c+NgaGmrBQHX6bjsaGod7qm5D9K49cdknibIYEvt5/0+HvVqva3WPbSvcV5LHTsg
EMaOhA4TQX6kNvxyg6X71Kv54rAAU8MWmzNkm2EXyY4ACkDT45bQNPx/UfrHC50Q
2jqsvvS8bGzgn2fiqp5qC/obimVwFn0coe6ZVg6PXxF+NGWf3ZuJ7oHYdCHRnDFm
/Nt1ZL+goKYWQ1vZUI7o5aZ0nGYTYgBgG8UsaWKR9ZZRaZ+gGEm9/vm0f8mwp9vl
2geq/EXtmK+btzliE1aEAjnz6a/LFkrSLOnmYem0fr89hbC2Z065uBWcgdm8AEmW
H5wHZN5YNLtY+urqB0btVD6OFA2m7LU5ngshULOnWjsElazhNNGXYdb1cmvnjAyt
r51/zxmUtg+3Zy5iU8xdeZqUq5opjGKPRnklnJBsB1mXLuqYo9916f2Qi2GTuZMk
tfZy3psFAjizBD62ogm5COqO85Ep+9pdXk4ihIB8O/kCd1lPc2scx0a1aC2xOyM1
+QHt021iXccLDvV9a559ITvilj09L/mqy2lUIC9WH+jdBVDe70Yb77bkdAjuS3BM
PzjUTfFitMO/LlYp270zmqpG9j0BRrVCHllWpeZ9B/bjry774/C5oHCBWtRXZiGb
hWXMFzM32vg6hiKBHvMkpCDhAXzaaWAXoVEx1rFoopIb+y8pt9V3WNqS4pt1RYTd
HcJXi2R4OPfSbw/meCDMhZKxwSjpiO3s1+RgQRlYVhGudrwk2k2wVgN+TH/AuBls
4AjS9KaTWlSrQ5OLW2vYM+jz8FtoekGcSz0mC5/ks7G4o0EOalX51e4iPlN6aSIP
zZdIHdFDG6VSY8SB4eiFsW/uQWrPtZ+ZWpprs8evpHzboOlSrM53t6S9q0FfUnO8
5O1HEelG5c3u46sMVAnsNk1Xf6p/un4oGmM/v5DAkZ8fhcVIAehLFcbeBpsVWilz
iQU43gmgTI+AljuDHtBIPjbi57NKRzxFnVcx7SamEL0Y8KVzFqtiGqNzoLUifW4y
iOUyq4rJVVzY6xvKH5S0bpPzouVJw5P/3t6lAwpukxcTtIfVtmTYxUeGQX9YiQKt
cVqZ9HgWFCI2bTDliThA9WumG8B4tRM4x2hy/VyN6oUJcpJJic25ozDwTNQOo4TD
VUHAW7el42S5KYpeJ4OTY6aHyUlvE7XB8VVRxziWLlA4bjtL1AnymPorMSdvkTax
ve2w8guL76gR1zaouhgRca+aO/InJiRRaEz4+Z1XzaQ4mDknY3a3dPZ2BTvEm/Zm
24nydB/d2S3vmg92M8y6hLtHitALfkBYT/oKVpHRw1oX40E1RNbYlOeaAASzhRwK
F1yoZlCVV5UZXMM0FlDrmZb7arFfNcwpJJzOX5bwT6yR2B9lvCkfAYjxNRvMoJVD
+MhIzF5UAIsjqW0mWaGMEMfswfRSWGpVaW/F6CAz9KkoLzn3T+ROSGSxgVw2+kiA
rcE0FwxKliABOfCmWyQYXl5nF7GLVEn+h8u5RjDZbhMDyScvizufS1CEo9kQmdUx
VS3XPBxMmMUCm9XSQr4nS8Ne/Nw9M99e/UyO2RqLlN+cNSEpkbu1I9jP3ik9sfHy
rpr9I797JjVp5jGHQuqjAoKcHxJTtKrN++CpCIuVJCLMrsovqu++xBg2bgjiFL/n
oj4ZcJVUCZt5fZZtb88QSogbDi1CMQYhRkyWvLeZjAkAlVDxor+bDwpScNhDDGaz
ZA71d+Rgi2pV6Bzwws5KBl8Nt7seK43Ev4NEtyFNib5eMFL5R/XkWWOz3DP/yLbf
se9l7Nuv5AnLzpbUkl+pjd62PwMvqgZEpSnpMDlYfvG0+o5KZ48HBEy9DOWKLXQL
Io1/gjwIWPALQgDB/NSGwjxb646CzmlZgtZhZ6NEuqgIWJE+ATDK3NJetZqV4umt
BUrZrdl51qIrw/r1owydBdV+xIJHShuttrXRQVIakO5+1fBh+fw6cZe6YJo2yFLe
t5uZFkQPkx+gh/vncGcn4oqcecsZrZ9cKdMez+WULLsSXe2p2NZtXSCMbSwgh44N
X4RsqxS7xgLcC3HAcXy1MwnX5xU46N5JekM11a5XcZngDsby8gT5G+npx9BRBUh9
38/7lI/+fAY6HBVqu0zjIXYPKxYsKu5wMhvEXUoI6HZuT5Q7FrnAPY52bGFBZEcn
QCvu/iSIKiYZktjrQoCNWVoMjHk0wzvSBJSumJC/J8N5p02/ivVJhhgTl63bQ1rQ
spoN5CWaB8Rbg3WI/pgBfx3IH1NrvlfQflD2PfTn8DEJrFVYS2EYggcyQ/LIFnv2
ckqjjokGgfSDFxjqPtGYjDVj1M2GIzs/MhaltadJk9UJaMxfrL5TJ7Egi1Sa62D6
ypnTg1T3GIC7xd/hUK503Csu6zWCQ97ZmQ68/A+SFZ4z8QJMeqhl1k6MKNk1bZJ6
DCbKGylRuc3GbBK3/VCdQWJ18lx4O9QdQ4vp45Pkzf6bxkMK4azk/KiXKFOv83LX
RK8OFH+jaY1QKnntPBFLIOC7gRPMi+UTPhAkYduQO/tDj0frQcBxVLID1QWyFzs6
wB2dBCy/ejpVLGPcUctEt2qgi3zb8dnanWAKmdkjCIiAheB08pqEoUqmvi1zG4uE
LIKiFUvHN/2Y9Bm8g6bei1ImeRnPxgc0bRQROWzqJFnESTqgwwNyW7ZuIPGlET3f
znpBm+UI7B5Ky8rO7hkQQhSnLK7nygt2EwJZHzqMU9XOOnC/xLlXupjDNZXFss/I
1oLe6IZkDOkOYs42yGxqArggA2ejckzwD9rvbC58hZrnTcfUBRDhlKKE6sBUYuYI
CrM8yvnVqepLhmdB0HkvMv161+OC+81DaGlhCGAIyYvgem3NIZCKDrCi6r4B3zdU
d8JYU2H39jvXu2nrxftQ0UG51WCWqZHjomQv0qUql+Q6VzHOSbkEmukrTACrg/OW
PN9QuvRgLT4KkdEY6VCtdhmQJhuhvpcHIGLhDLGCjuVIgQUqOfQQ+Yf4X/80Xoje
fwYaagaO1o8fCUe2pS5QMdVKNxz+8YljGcsrZxUg60+4RdC8flZj2GJwUAEkQzJm
kDxFaXet8bK2RxKuv6rLT47XSirnda80s+K8bgZNUeEB1ssSJxU1fexiBpsNzH5i
ZZ1WuQKf2d2f9yG3Y0+jqOxfbOWNwZU+8ewUROy2R+z/o0TSc1Jh9DHK9ZamRkXe
hmq+TuVYkoYWBUrHfuBtVvMSwSOc5yjbIdNOJONPvGkPm9CtAPo5A8gu6hrGsIdR
jZ7emZ/7jDo6/V5eY5rUcNMYJ7br0LBztrUq/6Jsmmd0UT7wlkggf/Y9VAKoct2Q
oA3VRfQaTaEFMuhixD9TyJKzXUUThfN33qGU+Wz7qcdeQj5ISC5pAlKbwMaE0505
GwJ/2mzXdOX5JuGHfGGNF0CShIs0SxZwea/6wBRXpAVNaN9BGmJ9v/d1hElY4YRU
5ngGu7KONwd0bI1iafDp+U4ny37RrqDjc5BNovxrOl0Zx+CrhRPK/JxhDGpLtj1b
w87DNNSmijH0Vlzfs7DUDHx3b/ybhYv37CbKGm0ZKp0DoYLmeUKuc5fCQPjF7PB6
Ow6QYnu95nNJLGdYPOodhrnZCYeRnlnaExuaCWbwRfHqq2mtVT0jkPa/RzzIksSu
ObJ79iR9Ld32LOTZhnsrF4GyUSpTHmoY/NolxUjWAVlVxkqzqbfNbwUjk4WB/a7I
lehMFhCgdg3cyK2cGyNRZHmQxnGlu2JbT4r5epx311dY4XUSXe11KIskPGXTGypX
XEBdKJQj7tUj2u2KumRahIrkTsDxoL21ujjG0913UTP44LNlcv+fqB1t1CG6m+Df
Z2lIB9289LDA8ztQvF3MiBTs+aOsJeigd5ARK36eeGm/kMf7J+Ud14iFPHEDFkN0
g31rLu/PV0fJjXVqk6ppAppbNqANQKcXFJtmN3o6c6LOFzt3vjYtiNganaMdDERU
YFfRLpGsr+/TUQG9qauLaDEv0IereY2f4iaf3AWzofqwx34k4OZavCYLtS6H43GF
igXhPhmP/RuSfy6SiRbNNVssmXExxjwyGb/b2bV5o++7XQQIOqn572OoQv45A7bh
vV4CZHhGNtXoH/F3O9GoTz/RzSO3TFNIGsIrP4e7G1a3p8tM8HudPWxDJh2AuUx6
95TPacspNaIVaW6flloO6yXPsKhrvAtODEX4pTknyizPJY1MnE39CAN+bsZ2WuV1
0VUN7Y48qTWAAL9G3lEBM0fJfimoX2BFgfxAKkuKhmWkmL8NoYkGGw+uAyOcmQup
twhnYZWgEzRNl7tjBRIusrmmjGs/ieXGSY8SI8tMoo+W3fu4tGUClh3E245feKgn
5BRoYMtAPr3OEKBj5Ntwkq0VcdDpM3JTmPnMfaz6bxsT3yRlbmX3l0k2lBu6p+/W
roKr1PA+aDYLPcz/3HrP28vnjC2WVnz5GXFt4mw2OlWo0PwORt2mKD15IXKJNvzA
93WSCJvarcyMgTqFIQH2c9ogak1ZFyNk/cYJrUZA+12pGLqI+aDLMdYeM5Gr+8Hm
6LGrNpV8rQNrCTgQ3E/7uj8jcRANuuqL15GHiFWieRFp8B/J5nL7T1Ll+dABgtOl
CYVMD/5l8raV5Agx0icy7HqqHb+wQOrEPFAD+1UlXrfWyjmd2P51UKcgLu91ziYT
8mL6MkqkDerZuaCk02RSASYv/4DgZ1OKW/yV9WK/XepBTMRVAa2lQTgWEADdDzCZ
3lGVragOwmCfmBYZLyERC/4WeY9vNJUokNbbjwUSqJGngAObWUHLzkImxFiNCue7
WhUneegSQD2fa9lBOpELY3lecUDzHTWsEkQn3Cb9J5W4qFjnCncC0UGJACSN1nAu
+x7oJObJApStZMh/wo89GO9BPA2nxBqvExRfTPEybDW4qvilolfJ7oRtEsP7OvXo
Ptncq8NTxfJFnF+IU8VTBlh1v8fb4zBvtA3PntCEQxSoMEEk7oACHzz6xvrhm5sD
nV05lwwrbCuOhtexfyEB7aXV1V0y8/tBOb/JcpymV9vZyXFz8GEaGAW9gvO2Q/NL
6jKWs99ZdTgRi02JOxNjHiUSXlgkpymFq8NiYLxLVbjnMjhjjMnkotAXG04E1qOc
7WaC4xyaDYW9hmV5+p9JKHa3Ptd6o++QyvVq7Y47R9UKYJ51DD1F4YDP1oJRNrTR
mHP07HJopxgdqOBxV50s828+5PAmQpp5U5EttOHLOKbKvJfScjlacs8s1rngpTFx
wQGJoZp6ousPMuw4rd3nkgCWA0dazhiOAAndwEwFAk1s157eOHUrOEHKrsdQGP22
+Zrx2dW4gsC4GcTVj4O7M+g4J/FikmQhhqgsdq+lErWor6Gd6w3cGs3prdZIzyRO
6cNGWo/MXywRxNPl08VZINCX1VYT056VkKvfsEBrk2Dho3j4dFPCBn5rz1yEVbOG
9mN2ka7YO73RIlfO9+B0Gv9TveQ1i9pdDnQDdG9pje76VghNabysVSXut1xg91lZ
k7603ADhKalLekLnnfM/3S3HFNL3f/XbdKIZGYP2BlFSSkoGe/pFC2qPWgffXyP2
cH88EeNe5xi3lkvMBkpyE1Q+pwvbe9qlqec6eDnaBVi2CGoG5Z0kXSQc9eG/ItEf
eOxFxKgdKYsIqY/zeZlgxlMT9NXEb9q+RDmJ5mZ9W0sdamj8Bccf7nZ16s10vNz+
rNmN7ZCtDaZB5T9XTmQwjF44VjpfNqh0+yZoY+xHod5joaNA2CHWgO0Mw8BQvQbv
wirW+OQM9hOWek8C7wvNpETm6M70PgrwzV/wXoVDgTiiQlnX18paR6synWInJlyX
AIrEY3XLaDE7yO1Uh/TYmnflV4ZgHLieK7T2FHR6POgNiZT4Iwdk3J1y1igEs4FQ
TvW9jC2ZEBNWzuENgMWTHT6vlgMqQDjaEeVoNu0+ZPME6dyhq682PkEytzpNYaaM
6bViV+PI7mQqClaE0pLj1KkJ4WgPksuhgxG5fXirg3z34BvrX2GJqpmwroQgsFUL
7OongN23BOF9XncdAqlzmbx9+5qSYlRXs3L1KALuZwczcyGhC2h+qTiyWAA/55AB
Nz5CHXz0+N2EdTdTCs69927rdFUPjb1r8BhUX4dPA2lNpDvQ09F5LIUmf1nVl1Jn
PQRX8rMWK+4+Mq9Y2R52xjcNE5wRyZwnjxgqi3lylhTXgCVlES/5mQsiKsxcmQXi
H22I3BHkal2mwikoj7OfA0JNHwdZ5oPNazU4ffOWbSnzYsiUXg2J5Du/NAdHRCR2
nZz/bOpOQJpWdD5xrpqLX6q6ATbbj1TWFQnIhZsVsEKqfQkcKk9rlcAS7om0u3gu
kqLe6Kpxr0JRg8nXnBZ+GfK70CR46yiW9RLNZ24LvFnjm+SgIMJv/5xjMpfB3vLN
ivAhgvLWNRsjoLkWNBwPfPKtXyAF4HHUM8W1rcKbl6QTEum8hgXixUfbApRlnbbF
l0U+/zUA34av06EclCG4C44qJPRoFuypM3ldXiNiWf0OGWKCcLjMZ6PwXZLzGGm2
5svbRnCwU3hodBXm6wyN6hpC/I6hrcx09c0FWkIRVXViB9Yo8XbYtsPap0bf3Il1
R2/gfzavX8HtuWD/ZLcq6aIwbmfZB1duW7a9oPQUJPZw9yBU/qDwwPtc7dV4Txx3
6TUgwS5esAH0L2W9Q+h411Y03fZinpQzYOClQJbT3ALU5Y+gyN4MuzS3Z7nBHDyC
uTZMXc23buxhjXxW/hKmyVRsLCSKW8wxifFv81YiXma5Ppu28sz8IUAC0RKMu8Qv
rRjbtxjBQl1iT56ERdmD3chRKC78MJf2BJMJVU8YC8xsOSc31yAP9FMPu4DTmH+u
LLoVeakBU29mNW6jju22iq2ibgT5WI5xqG+dWWe1u6cc3DOo4HA4l1jYANCI5dfP
QFvscFpuUl8oY77vlGww/aInZud/XdahKak61gCwewzKk1o8kdsNjOah2l+PF6ZP
S+cVlnFtjnqagsjBj1cBXFCLswZKUMdMucjtvfrcjzpfjTXZeOoO0mZmhDQovz+M
AhPGQ/G+uYalOX4jmFIh50g7tq2U1USNJ0ijtH+5b1LV3JhhejWXXX2QA6ULTVyF
p1U9UQzKvhJJzO0OH3LCi1ywDqTaopoTtlb/GxNbRGGiKoM44MaDrO4gzf4UZpK9
+y74MvX4R4K5Iiqhi0ZATezUaWXiytpald79RP4rdCyuStiqMu82IlRjbz35XSgc
8GF8RGW+3TxxSeBjYfpRIOCgvuS+CS8tgCVaAv6S4Uyc1kx1PCf99wlXi7hbNspW
+Ccdt/k2ljqts9UMRq+8csiJK4s/h/5iudilBwFV75ZsfRLKiEtxOsopqIxz7u1P
PQlfN/Bh8LMPRVP4bkDOMe1C7yuQYNwM2N6Y0sNqDpTe/k1+ZnFBPCMbXNLKy1ke
/zyHhTDdwkdB3nwhv+cMIEuh9OhWZ73vau6zMv6hqgfBuAqRB5iHQch0QpfjBdeb
4t558fCmdTpWAFzcsX+lSkysB4MS45X3i2ydwlyS8XmE+r2/auSg+ih9b3+BZOm5
Whaawl33wykM5K6Vik2KFxkL1HzSlx3py3gTGkoHMcCmttnR6mcgUgk2l3YMmTkE
13/HcCWieNCVO3U8DrGio1jePirnUUkh9KUNY2keDqgdsc/wkxXj4Fh96JjVNvn4
GjHX+u7Gs515rWYsDUvZPA1GcTpcx7Nj/rNqakEOD2gZC7o4aJtSodAGpIPAkxZq
leDw9xnqjlMiRBQvFzET67oG87YUtDRxhVMNjZZovi4vXBnnsKJFg9726FNtAvig
1ZjcBUMD4w5a/eRapHaaQxMjaJXX4BHMnpX8Q2Pzys9vvBNnJfehUsTYnr3KQ2hE
q3GyGUsYzOuDErGKi4PDRXgZkYIWYXK9r4GxpyLCyyufhh8uPtgEM1YBA+GS4K6g
35kU/mOnnK1erErwXzV+iUZOmRTQnKmFequiWkVmkt9YZaK1GbuAy21upuqYQvN1
e+a3/hdfTorf/SuXQQjkjvBy0bVK2HVwwwXxj+qN4epCzEfS8ATByjp6AoQ3yDPI
3+YydK7BDnd2AC/oxbJIpNjBhlkCiccviJYw/6Der/rTn4MU4XPFsnHZmVaZ+voN
V9GKtHBhzZoeewKn/NEgzO/yPuASJ1oTzO0+vmCKG7UGTOSNHV6qqnjgYAM+92yw
rsBda7Y5Xt9Z01p35gqhDFOdnP616M0eObceGNLsMTvAGAAkxZ5n311QWqmTtVLp
TyTLRYjF8mgxMBK6sTO03918xXVW85JEKWgXvelaKgfwXiy8CBwNnFh2e8xQlItV
yS7kCkv+tGB8fx0SkRG/sgJo5PspCUZ56frZeeooX2G0MuPuxLJ93eBy4obM2Ptv
IRHNcs6c/u/KXbdAgJl06+OQJE9BDr5QhFTfFAWPXJdaRzfyarXasVWuvfn9kQj+
mYKmPNHybgw7mo/6zSJYDZfNQGlY9V6bfZXdF4/eMB+QH/Gcuq2F47I4DKW8uClR
esG6RdW5ZW4ivBDPr0P/fJ7Fr3RTwfRrx1jYW4xWQ8mAg2lJdub7xOGS4uKf995t
inLcW5bsNf86wIaimdEm1wC5AQHY4p+i/9adnmkua22UBDb1h72iJDOxzMTdQrBE
smIvyValLgaAnbqZ35XD1kB50ua+P6yM0w2LMM1k12A+RFAvl3a3oHBngRTi0trG
yh+PP9TrBLkq5ktI9ocT03JPagZDn56T/Zm9C37xj3faWoHb2XSStf89KWvCtBaJ
DG01jSY0wPBFhh2+FtcqtR87yD3sXznuokYFMGytaOW6Eoc1UK5PisPAtsllL7NH
2UVW34mHEz6lhQhJfHT63kWM0DWbkNyp56J6AN8y66Ec+L4T3YbudNowCfppVWJB
mdtpPqqDJoqPIIF8yHjDMtJj+9OgZ1A6HxCS/RCDxrmRZtdHKPpRAvsDB35iEWW8
ozKvIk25dTnzo46w6tNd+MmX0R1oX1WcJU7Uztc75rdSWk6+UL8o6ILrwtdBkqq1
k+hAn+6X0gELQs8OhZbL05pg0PvT++V65r4ydkzw199erOXqeupBzELldrU1M7iA
IRsmmt42ZsT3/k1GZiibzc/RvSsM/Yz+q0OoAQl5JMIYV0rOnCkJJcq8AxaUASgw
3RrQ8Drtju4PrYF2Z/hLJLGJbEGfegPjdHLR4up8ydSJFTct6eHKeJo6O69apYHZ
cJTgqCHpC2o+OjnPIxN7w41pJzqN7Y51Re/YuCg29VwDubw608JejD91qD2x9SWv
KOr5hZve0PZpezEHFHDmIrAkMR0O3twCrHnfNXYBhwLU8ojKIBpy1DaCzHm6bb9n
cdLuasiqxM2RW3/HTOhyCRwTHVu78gXgMw4ikr7rF6v66nhyTyZvjstvwtO/GO7f
vcAVA9Yc7BIJ7Iz7+VW4ntGyS/C5bw+/krALkPMKrjd6NYAhvG41OmDexXtg1TSs
XXIeEtTgD5Z+YChEu2FmXH5NTsjP25/JieLQ6VpsvNiYICJ8Gu0X5BwDp3U3IMpg
HIhpWHizago3EbXZC5kPqQJQTJKJUcNVnU5McXuQ7ZEbe8n1ACgt/KkgE5RNehQk
In/JCgcTc2KMVlF+VyJ9B5he2eX+Onuhfa3Q93SM8NtTRNQWD97yqpBatubKP0o5
cBcE9Lnh9ZMbONjBnT2bhngw64Quo6yCqi05+RJVAm39y1RdT/xsF5GP0o7j42AO
zh/fdG9/hm0AlM7G+V9YooKprSShTah0j3iOkWPMrHaKrb27J2a+rJVYRcD1crNm
LIKa+ttEAPN++7HymaR07LesW/0pe/kp4Hnlg1wvqDlhEfzpYX0TyO4Qiu7Wblmp
QwM7OP8LBnCmzgTEn4kCUPWnscd8ViCA9pPHk6EDj1nYCSSj+mOasju0kaBklYPU
hU7k3ROUy18+G7QnlpdaKkMqjohBgHIgxDFxLkX+JlEmU/kV3DN1cMNxWGpfMOHj
ogvpKn81m90Ky62anp9y5MFDKHRDU1IsLK8ovLHB/Ij4ibuJNFwUKEnHAsE1h82l
SxHiX69acvbxeK4OmBmhDyaeyMW75+kiMqQflPY9mBeBv29R4bLnJj6nsiVxGXFU
UoC1LZaAShcnjCXFnd/QZx/MoKdWK59tigrt2p+tvUKsBo9cMo0/saMaKokcMj2B
rb/dh6gDjcHlY7AZax60Ze9em65r6BVsLv7l4NBhlt48vbLkN2iV7ePwzaSyJYmP
ox3ce1xfLsRxzNlb+hYJ0QuPakFMXgTFNov4JGbdUlx1v/SW8fGqacC8gKI+UuUQ
Pt0Jcj5sTMdNLtn1s+hnPgP7et2DJ9zZTfmdLJq+ovreNanHGGXyEdeHzRS2L3Rv
Qdo5zBq3hfkE4jSd8ya9s+MKfs+hrlmukVSmKNaC0U12nQjzMvyKK8f55oUGwAiY
ci5aC5Gff4kzf4yua8fYp5tDqMWHQCoKvSM1rtZzUjrUkK96HhNYbmHdIkFYi7YO
vv+HFT3D9suXSMTOaxgUiR6zOTTWr0LOw4EAlB3dPrVbLd1spnmBrjxQuXCQVFjQ
DKp6yLfCyUJx5noMAgJVY5tbwL7jFkR3giz2siBXYw3EGovuOEJtbgA+adrWa5LR
oCGYosHQC9gop3MATKCuYWqWB6keAcmp8udzvtrDz3waCwukZ465ZbIIljaM3N1i
p/uZNNT6J3KcBxpw7NrLngnuye+7HYu1T3wIqnNZGF8Xmm3Ay9YuExfjWDKAmq1p
PrbutviLa54cVaBgMvT2ihKb/6w0t2REEP/Dt/9O2HATctGPfVPTgdrLzepc975D
YMF64+1v6sEvKsr3ZbRLzEJeO5Pc2bFDtJTa2uQOSsaME149nK99dVNJ7kHCp48x
JDAjmj6ATqfL6Xf9Wn1j3wysPJkgyHAOJxwBJ5OdC+3x4q7NT1a7gvnQCNO8uBb/
7tEffJMl61UW8uWHKpz9DiHEHOt3AL8MlpcANgBucpIAsKCwRkma/T1z9+Q6dfVL
yB4FniR66EU9IbhCqmseT8ABTDgHGdzsvrr8hClighZ3BxCGUF4U9zJMWIOcu0My
I4YnopEFd3iTp3oIcjDXyMS0kx+2OQdMj+m8AnDFx8CGrWvY6tCsZC8V8mRtgPR6
49JSvUt60cUufCYoXUjMlzGH2Fes58JOQ/fbMAPwPTli4+7hxOIRIKtkmEmpQ5QT
UfyxhyExZ6kXGy3KuQYFPUfKqn78fKC5oo9OPUtboAAZk7TYUsKuehjOGrybjPKS
m/2PW//Tryjpu7k5yOECm//RCdo+ov8GeeLJMzprPg5t7cAbQSJa7WwFThauBKr7
comE4lAwxd/2DI6vAqkAx5IV/Ee7mSGlXRHZoIr7IFdLZQhjn1F5Q4iVxS555p0A
lHAW3KjCW3E+JGSNoqGwJ4o0JQrwQN5za+6hspBxyhcZGsKAT1y+vlgYqXX5uzkH
EICB/RQqIkBo0cu6tjKmpZhyQQF9+KBXQi+xsKYd7CSHD0GLbIemlnJUXrIkGBX/
CIlpYJZhDDt3MNN7/LbiyB3sLlji+hM6k3s5o8gktG68msCclqGIaEHATI713zJQ
q9WHXm6vFWNL/x/TA+Sv33ChzryUEczHfE+tESUxDisK00NhN1IPDnZTSli0ujAv
bfR5MBJ56ZmqM4UfBU9hm5mUvYxFtcB/fllvs2i3Ww8GhlvoGyB6R2U6nOz9/xLF
h/6l9rYeRzBCanYQqC2Vt2kaKA87pgt0HjM+tZK+yGbCNGnwjiBIf7VNyMjHZnve
1Bk1rlxo6c1RyXngG3s/qwv4x6dE/FC9AazN6GhANW3TkTEgjYiLYYmBzSoMG+gM
caq2h0BlLGkTTet0UibnHODtXnbhjMZjOCgY5h8mhQh2OJKuM5JlhGixxaV4Y+Hz
s7u0CNHH/CU9VVtgN4/HW+xaBR5gIP1T5F5WRfw00aeuEBCU2PiNs4cBcul1jyf1
0hJboOAjv6Fw4dsPfm2WarsDyEye1IJU4Q7u5TRnMKNisNnzITjE2i3kDrDkm8Dd
m8rTtXoOuyRtxR+nm6qNisbrFob+1H26sRHWJeqwIISSfW9ZrGN/ZqziOFGZqpf2
FxGSnIVQ+Mv25LkZ64++7TbIMFW3u8hgrcu2U96NnlO7DDYfykonMnIlVHg2r+3g
oMmQdGTvtuw0tugfdtmSOnaaR9AZRZ7CfQAEx9ehIK+g0uVvc+f6JAN0NsMhlnv9
h4lI6OiLKyfVIK5rS0mnKR/uOx+cdxIQS4H6K4UOPbmCDjSHd1zWkLnKSt7PFg79
or2oZyHGiJgbXSroKWCaqgp/dTi7pmYcY1CeqiWnTXb7p5/p8XGW6GdPQYoQnHBC
lSZ+WBYzXjCrCDk1fxwBGYfI3aULa+9O95pFxRKO3hDvpGPUziI5MirhzXCHAuJS
edGHHm4r2uuFFeb6dBafA2+6+V4RpuOjXaws2EJ1Gr+XJx9RHlJLjLMmjId8oUNo
dTiJYmqPvCEYCd8Bap51KdaPkJXCTD8Bjsi7nS2V/oJicuO4CkbtuAMeN8tN8dIy
7zSxSKudQ5qRjFq6VHjFkkfeGuueMpn7S8X79Be00mZoM/NmzVEPeslTbXTLwCQu
8tdqC6VTqDT03+n8Fhi2Xf1z6VFdhcglRkG6VxIoP1i95AJATpHPNird9Pwk2QBD
vzcu6QRokJZZAV3NR9SdQQcgb30uFxS32EhVmJZYLZzktTCXdH4l+hispJaa+CwA
2IziOt8WV0MXgyOg6fWB/uQWexAIad8y73Aj+0TF71j7JKMjpHkPc8XU+575C2ix
cE5byUWksFROuoJyI9cN2BpabxBeCIV5VJe6jYw0gSBHa+Hy9E7J+eH3ynXluvz2
v45ZM0+U7WBreoKrxzY9ZthNQXBw4Z4vBFbGEtMpzhVxQRNdRXsY29Uzb27RAtIl
3dsuFKh0Rfdde32PuvuyNzGmwifr/9M/dBM72lzLCOuOCQXoQN5izPWeg1TX784Q
j8gDnikq6L5P44VNg4byDItVke+NYjmc/dVHW/kDScP488DK98RlePiLl1SsEhI5
7s3s7s82MqhSJW2jhg/J7H+kCa9NiH1Og5riy3oHcehdQ/+RDCp7f82Un0jhtahf
liLqRAaxq9vSfCIzkjyNLobimiSJfr7+/TPXSHJE8D4qHKnPiPrd4bR6HRfoMc6V
4Q7IAozLnmLwfpgIQ7XNLvKJ+WHtpDZzDTI4SSU+lXsBVVSjmSpILoFBO+slTW63
Uc0JKP9vNgQnLBuksvEPQeSHaUCRD1NbQmh7A6x0RCMe3l24xL3ObaQO6Uio/VxQ
z5XZLEszSiABrGVa6qpzbpOA1FnPiJHrHXpWQsgW9KCSmepbA17w/UTS4ntDPxUS
f4pREjc8K3ODPN54Rk4jn+IvQ+scbxTBkcwApo9ASovy3oeNUoSY4Pd6FDe7aHVd
EFnzEte7acF5GlknIGFeU0uUq6UrAayb1q56C+2rN+BTvrK5jOPHadTWp+1kQyV/
yytzZszKFsBjXz9poNo8mlMoneDMdFzRi+diqF0uUaVEUoF1KRgJAIs79QIsa45d
7N8QKeT0oSpaKLVzeZ5gQxDAeCZbSY9tb258QACgs1Yxi35mVTcR/tsLyTIper2s
A7z6o4UF/391YZfvOKNkXlbaLmpSYMDBuFwA5usfwtYzjAv3NNwNKth6kjn0XYJR
Cp1t8bwmslpxNVwLAekhbDCUH7eQ8ecJxMY4GeJrUqO2zJq4RdQuAzU+AgsftsUo
E2LfIU89ALx2g1mIeQVLEnob6Mbwz/c3oTsbxvxbhUHy+ir++hHgWB5UWF2PW67U
FMWTdssu5bXFEvT05TjlCD2ixi5/RW4+Zc8yNZs0OOwMVkKyf3rVTqPf+qW386jG
jlvugLbvClde3dWTB2gxcPUXY8ZHYp7ivBFjwuU0c5kaVoU4HJ0ZO1S73O3CA6pu
9T+btNMdmxuMXqb3g1K+kWz1B1R936UCS37vcK0/BNgH6+FU5WtAQ11lyVtBeOsc
9Xk5+MKaVuIhZT0XhFtdqKxRD3SPErGbLx4ljaCkkNHZDVZlmqcK1s8bO2meezQ+
D7yVzmZAnjViQbn3ZAC2XyabchTs6vD6fE/AOIuE3ct/rKgIaIT8QgcQsjGHbbyv
z0vUIkSAdHrAO1/0nHAywrc78xUOVy41/kUxyEKBep42EqM1eJHkFlrWgudfpxM3
28l2gCeIgImlR7QEv5UzIuQWyXt2kBX+whW3JZ+djgNJSy3L/j6D2hdiiViCL/DT
3k1xJsfPfV2DFtibfL1OMBk+aGhlcjRT8oM7NtnDkB4y1MSTCW4Ym5+WiuUUEH8E
gIl/enFWDDSvI41xIaa3F0Xw4lWWfYkk1BRAZB8ebRLlDKnuKVlEwirprx5w9IIF
fQWgzLbXwqjRs+Fm0TcHw49qt/sY+UB3FINgLxO4nci5aCNXZIRQCY5vU4MJXGMa
LLQkfKj88F6LWGh1g6aNeDrZs74qhXDFRf8hpODTN1T/T6pZgN6A717ruXuyHvyf
sGyp/DSjcpFZiddDBFWJtQKig1C76gxXXqt+x08Xtxsak1UAJ5QR1urg3RiKlqQ/
q6/Gx/dnfYaPdCOBi+ajAP3B5FN2WEdBT4y/t//DB7eKhCZcE4cE1C0mYZAu+Xe2
lPJe7neMEtY9HyRJfBcSNVnGcrbYPz+nCksZKWql2fojJrtpzvQRSFfcQdIfrxiB
HX/4EJPlmkgWx6FFEXrta6HoQlNmxDuJIJC6t/Kb6EkJ0oj+/Eia8PSA7loassuK
aVKBaqd1nMpYbI6j2Iake07zS8T30YEG14eT9nQ9f3ly1AhEysEih46Rb7t5zFZr
rgw9qdFiDX/R162bO7I58ZDQH0ADA0W6KDgR+FlKeQo5feillTpfSFWBmSC8weCj
ohZuoTzyLIiA4mp/z6/R3V5uNXtg7GmMT4XxtC5x4ThI6nxcQLntsr28zyz0rDlm
IJnz9d7lmJZK+jCYbfxPGJqyPGHL/ieVGkZOCcN+dyGsfa9CAH6PNZCRMZwnow6h
IeGavctOei6vDpsn8U49khHQ67l1MgEfu00nff7oR/QDCRbYHSDeQULoWXP94Ma2
RWQOKTW2Hfg+ykS3wylV44ZT08SZh12MC9XKFagyXzL1N0eLZscpnszKuAOhbT6n
YKJDwznQpL0OlSANEGZB57HuVRUAuwRAv+dzF3YEuCNQiAu7GtiSQPrPa+6QNvZa
blFVuqsVp7SH/o5oyifRYof4U5UJUw0RGB9PiBkrrWuCrN+aqhD+f2xEqUCljdN/
atjcsd6TPzP3gPWkf7TExVwAbi0X9l71JDbEkQjWvIFbIgbq9KE/+34KXGxzPM5Y
pwNW7j2rOJfaJYjlaOlwhn3/QGSUU7wHHKRhVl2crQMhJeaL2XmIm2YTvv+uMxrD
F74g8yHsQeTN34eVS7RHv4p0OQL8HfinfW8BZcmbdnfyGDpAvnNirOjIhdyl/Pp0
hinsHa+hvEaUUmXVsJn2Yt9Ydc89wg6kmlCdWxtcM2vAwRMS03UuS6fvez0MCNuu
6cJDAk8Fbsm6Ei0trvFAnl9lCBVIAbHWHsMCcsJ66vHyJyePhmGg/iCD6UD1oLQs
A53m+eSsgKIytSfKu3kl/OJYj+IEs0gUL70ftGfsVxPr93W8F5kEui0FGDhhIplk
cr0Vu/ksnWqclAcT6dua4gebTGHKkQ9nM1taaDt9CVvTWNQUlZmC3QIdXo/2uaj/
1Llh9spYVW9/RT0qOV9B1zeLyNz16CfEF4Abq9t1Ra9IAFw09hO6bG5e7w9YBYxW
WckBW/Rb+vJvghCAFUf8kyBn8BxJCsthRW+8dml2gUgDo7OGNPW/ioeJAy0V3zzP
PB3amVlp297IubrO/UF9CczVhVSClnMuSkvxv4ygrciQnk/HPiexZW5BXw1ra6aF
pMwPX63hs3FkE1oAsQjgmp5hRF18pLu3f9tR+w9woWxF/wwdxbZEj83HhmBTqUUh
OXk8uVctBynUOylwGH9kl0J3spDcPCTX7ODUo+qD+OhW+pjp6mMo3XTfhG8yKtx3
1z5OI9lNsjAnQF/HPRB96kWfEBnEdjVPicJVXN2h6B5zA/aeAsZ+2iYk+In0WtWf
5WyLlSJ7Y+EuRb8bUJZalYc1qgTB2SKEkJB0/zZng4jVMGCBLGci56cctNu5fmOp
Hr7iV5ntT/mSpRXYtLKa1kO4iqP6lNYhgjsrWeYeolloHMNp9MPdG1Xw7cTjTiMy
5/CdnFKq2bwu+ZbyY7I50HfeEvB/eNMwU2LDzrlohWbnwUsYFzZzuQR7MRR1QAfS
yq8Bb/XWdkKkAftFRvuGMtVWJQfTVlGhXswK68FYgTUiNbCxhz6oFYAgchndBChw
gyusZ4VwTie0D5VnWGF6JsbWVABV+zxH/d04YogGMlnp4IMkmM/qfkeXt9xyCkoz
Y4EoYAPCcZkslMpE/scXZNzN3Dwu6TtM5J7I1uY+fEXxkh9QvrmxMI3vid7tbGJI
PL9yx/V5v7280Ej5llnD+xhHrSSpQOx6E0xqjNAdx62T+w9CBJOsDgd31bXvrH/N
5KBMGeiVTAOXNfvndxKZ5F78L1gTEnA+MsyC9cgJi3vH8m0S/o3BLeFhL1Wf/kOj
/dlrO8uMxlfgUlIieWAwE6Vx7Uq8+JFj6jenYD0ryTkItQ4gnqmuabsN/c+JJY4d
Z0C8DHqbWVvfJM+dJT9yDSKPKjUlTiGIiXEV6M0nEwox2exEtEpyaeqyOZk2OMCT
rjG7NZ6YjTlRsM/J8t9HO2GWfFxCbp5tBcIvasPUucH2L22BB8m6JPCJXX2L7k5e
u4+fAea9iPtv/Bpiz5vtGWbmlq45JFMYiOe/fbB+q4ojfTLysqnXA+SAN+sdpWxa
Tc3phLOvhh6/bQH1moMsbtQsAT6nQD/IvxrxXEA/5VF4KJCzusLp02wea73h3JmF
9dxIj4m97FFORzzyAELAlkj0lg/HjYCUqmGPiysbCit9CDDKSLos6KkhM1EbT1w/
EdzRzsXQJWwD2mfT1J3S9FDr/si3WSylXhvQ1WDRjXBprEWhre7YifLXy5+5CDYb
80mG6nMoRUw8jiH4o4pN7zveqG4zH/ia8QyBomanIXvm17QgAEHGoTy/2PqLqn21
INf/Kwv3K5smzEagWHHIERG5OiC7tSHA36StLXs1pCklOLhFw8kLITc0N1jS7yQQ
nDMspzSjzf1Z3I/iEV3CfJ8VdQjQEBacExVSlwW1pBvrl/+DjTUCFrlhjhehLN+c
JlgD6V7jFATs5e0PYLGOQBU+JOg8gEirmcOZnWMxvXv/MZ9R9pwSRnedPb/O8Ve2
6vdwWcWH1DBKlJ7dAtKR2VnxuDSUxFHXSwCTpdAwNl8yxkLWPSszIG9AgOEzlGmM
y3iKL+6+I8erAlW73wDaMmS7eGhJiiqcB0Y1ywFaJJ3Dv36r8VEZFLge7JsMlzLZ
+4G2DolrMHuiXagmyIjQdFx7LzDc/nvjv5fARyp6pISCGtiT56302xn+WyQQByz9
n6DgrY9l0yFZPCQpPtZWkalLq85zbIO6Mgvq7m/46EFJDWIPpeWkNhGO2CA7VUuQ
RzmA+jqhYghgXSEUk1L9KOwJ0AW4DiSg5AS2FarfMJP0NZ4eTyOnXKZ8fG7n3Kkv
aUHy7oyx/K9OsciRdR9MxP2wI2blwUUh+AR1vp42UmEH863duMLXNrKHCshcNwG4
JSkG3mpPyUo5zL54wh5aI9UHjN7QZBt9PVS2zQKdKSWyVipDUMeA459Ve0JkbHZr
sFY9L04RilV/wpFLAunjBF7JBShfQD/jJoXWG8GddzQS7+YMks6tdQuMvjPZ9wSf
6echkneg46geVneGlL8gSJTfFggxzGeqM/yj4d66mqUqrvbBj04cVV1XEsL6U36w
zcvS8zmPkKW4bC2GgvMLC6K7esQc0cH06rFN7mErIlt7F/SfFPCfjg/ajECzLKCz
zeRmrEUZGTvw7or/+adfc9XuU/llRIk3DGhmxVJvATYNrkF9o6ECSPUAKrZFD0fe
n3zbnKDZUlcSBuJfaalL6/dYu5bNW/wft/wafOKFXzKpIuNmhfPywc8e2uc7lL+g
Q0+bd+kECKV3WENiHtU4kb0wOdZjTKI7hX6blooUOqorxBwfRGQvqX1EVl3hROMS
jFhIQofToB34PXuXQltULnn5EVLVsEmfEZgvFD2qsN8y5KqLM6rmN7SvcdXymN1b
UHD3R/U6iJlBRMzU/rCnSJkCetilp3nroQ8zrgPsbmpLw6JPQZb7sRKlxjpYxhdK
04hnsZPydpgwGjUoGoJ2daAdDBTJbMKFEDQL/ZMXJLafiNjK+AE3x8t7Gw2Z8clF
G021CzMsmopM7FxSj1rK3rVedIulyI/iU/JmEh5w/sgLobAWJCo2bU8hFK5sP6l3
Bnb+2UUH/DTamepNAY1Pep4LivLG0P05vTtlyPGNjLcUDS2Y2dzaOF+Bmlo0HKhM
yg+mr8epYPYOLJTFWJRzL4B+DxncVe+n4seu9a9jG70SVI+hBRZkF+sjTZZJDlit
TifdHAoqPpyJUkTECSLn81v1WlorOBD+bUgzkt7RGGFBGF6HQvXq9hvbbO4/mw7C
KPs4xqVATW5i1UmdOq4z2r9YmzRC1JclvCygcATWVzls38Q+cUxvlYAkTR+Yug9g
iY5ZVYxkBeWpFvn4PuNsJ9XSd5ol7j+4eE4ofmh7VxN9JQV6ZR5h0JZR+CBwWVyy
s0n8aapfC0lmKUMVJAiF+y6VsOzh/5MtHtD7+9HdPWwhH0rrv5wHcRH6+jV6hga9
zi2T77ILQLDSXnc5Q22Pw22lLHuJ8xUFJVCAdXNx5S+eU/oXionQjkjN3Slbk2jw
cRWilwWP+ZbYe4KlR1hJfwxxDlvsJJJtQ91Kp6K9HBqeavcW0lLTM5EsdV9IGBGn
BjsxfhOcKXTKbettJfzz5aM9fRBppazC7RS4W469s0fx8NtqnhObvk5o8TUY2NMu
If0eqv+wpZm3uzycN58ki5Br/ZS5HBEu9KHj2khP7B1N3285PjGERqpCzfCL9qXO
P7d3AkXd+T6CxtkDULSZ9ZCkmlz8p+R3O7+dU+uze/IWzHoOzIm2Q/MXQPwg2amb
QDrfEr0tESk7Vp9THEvrbRzuGyeiDSSh2vgSE129wkl/dj1bh+WgtRL6eULTst2T
BkfWB4WI7cxKXdOJTPjSS1lPtOzV6sRB6pyb3Lk8dKk9GEWOsaTw1NGim7pellGO
4kEXgAAXtNX2P4w9fQkGX6gvHWwSWuiFKYSJwI1lLcdz+e9Qm6B3yA/L3dm6ytH7
aIoi3w1gjpGwLs5yOD4d2gydzo8Lys5pqPQFEYkSjR/x2cIokao3oLvCD91baeV+
ovRzf3cQkw5E0AbR9RLwtIszn3Awc+z3WTfGW1NQnLOxHb4HldlMGOWzlyixpd0c
xq7MNsC0OnFmTprB2FbpOin5jbQhAFhxPNm8VqOf//M6z4vDuI+hMnOcZ5fPCbDZ
HtCI4YjJecVOtdxDrer18HGol3rG1QxJhEnWULV3qAXf5o53rKqRfpY+z89wjcUO
IJQeRuzjinLd+Ux8c2irOwydRakHhySytSxxaaLaZzniq45Klwsqg8sdbM+t5IlS
74wi6uryLk2ohqV9df07RSHyXxsaP1B2pOU0e8QWWxTeAPKimitN0aUi8JnBcpcZ
F9g4cfH6FTwsGTnpF5F14mgw9rbjEidJQQBktjF3uUMq6zjTdtU5XhXidSrMHofC
O0AX6c3btrNKPcqQ4OiJxtEaK3pYAM0QWiFdXq8f6s2QgqzUVUPjOWhO+41VS+HH
HQWmr2/399W0AfhSN3e1/JpCXiqAVqWpj1TcJ2avuOSGRpK+TkP9SVzJwoVGL6Jc
SD/CLtB3osxM8BOh91A1rZ0+seWxAI5aw5vTv4X4wDI0HVH0+WEyvoaIexluwrMB
2ol/X5exd7MJdNEXP6UI/GKiF5kYSeek/ftjT4+bYhARE2Kb2F7RmPirjOiIuBS5
KbNpuqFnRHz/xNJQScEBcCgnCVFJLBDUJiCfgt5gEFp7BISV7kVy/2wsyjZDRnzr
cN2jnR+jgp2/KqZmOiZDcsORmCaa25fPf/FHSt29MMDrfmn/5rFxcXaOVnpKTYQG
HShva1rmkFPvSpoju16G/NorZ8l9I7MPLFe589X4CyY2X5bUvlDqWY6hoAPUFTR3
q2Gg9uRViDJg2s11vXQz9Qk/P0kg15CJiF8VVqjLOXG/MJlxtk0PGsC20DdEttpt
QpiygfM6o1EwZ0ym4IY4w5Akz4kBVzFtf5fqJg6Hhi6/JAvWekj5VJcK6kAJKB0x
xolRavM2O2R6BRIfS4DanaPY2txO8oRANdgk3E1HQ1AGvQMkPPHh69JNGf7JOZo+
TEy1uyog3JtT1NFn/+Rxa7W9Sr+hMkDlKhCXsvEECIyJInJkFUGkrRTYFhnkQkv7
qPQe6ORlSOZ5Uk0MAycVON7b+4S9PcBcDfZDr26QYnxlwAONNG8kRN2QoEIGfrOE
vy+cZL5HcBdg5dY+1I5sULFjxF//OkXr1PLVG4YaaNbffPp7kE3zKAgA2XDv/wwc
klgFfEKjZiM3LI/xL345HU5MqghPsUeGZny2JVqM1FMJfIy+ZpTmp9PkT1OhjuD8
/P0zxj0tqmla53pAJlw7CANHFqZLVRWs+1rftHy8jLSydqKMqi1VDRZsWw3bBVje
e3/50yC23paHgXSyI26NX7s62GZUD/dkrS2I21cTKAZ32TRJo5WUPtaBTTdjQOH6
leQuNujBi5s6Bm2SPrnkl4s+hMPJO/O/MabeJJErLUgHSfh05YQJW/zq1oVBObDU
nOEzH8xpwRLrH5EMdIBoYx1Hi8mNXCNn4bVdRygpE93LsMhhkFcNVqeH7EpdSEnQ
TaMXuaZF+40bCgsvVOrzA0Bm/XV3mhhd6VQq+28bHh+eWuSsU5AR6EQ5JcaX8yGS
puqYIAFo9Ry0XA37D5kCc6uEHcsiNLSrwwVw/5loEKxjSRHd4z5klStQnACNkgNx
SkZLU78C0xgatfi+ibNcUuTTPTS6Z55iDuYUmzIe8UwX+1S2FMTgofX32CbOTDSa
E/7da0I8CabpGbs9DDoZepWfnQnOD0vPIWbKaaElXMIPDO64942w+SPkVoWH2beE
/r1qOE7LWifL+2+TOIxYlIoVVEdskvhN3SAGttiUWX+hK50m5UynYNZm695zbhK4
3+Kfw+gzOUCkeByAAla6QZ0TDFAI7O3xk05ed02PwHfWCm9nrmyhMNxrS6moC7md
iYEkqiT4qYqEqmoBqBQzLjA5h7WlaCNAty7Lrdb7a2/I9HFbF3UgYhLzvdEJaxQr
sx12+tOpC6LFOv+FUb30xIcblTDJr3rDDJNk4OIrUwxgnJ77mlwxQjBVmEo3/Z40
gKGTo3ZkVZZWyw+bQOzPX5tPfTVFaX4f9GaxHAlp3hup6elN/FBAGvQrynnHccku
rzUT6v3JNmRWRE/N4rM1FOrUh5yi3Wp5PJkAykFF+0Ftb+/dLBO609SXO/hEA9Pl
AUSjInvwFXquXboeXUZLLitYy8UDL40VBrvm1qDLwZx+5J8e0+ZEsJPcizyzVJiV
nd9KF0y7TS8l7U3E6xJLpSFORl2lZzrFr71X243DKyEnJvZm0wy5H/MW8ozfnUM6
PozI4GxzRsK0VvKnbg+Olp8KBU4m1h7VL9Y0gaoRxu41KWxHC+CD7awm+7/Qb4u7
++sgHixSWRfQqhZ4joWcMA1D3ZbEudjEEsU8jFi+XfUCi0xENKNUGfjt1joA/5ZA
9MDGHit0mZ8WG3aFEIyxTQREv50INXNHG7aT5OpK4yBCB5g182nYVo+QqILK3z0N
NeyTUQ1BG6ChrenLZk6KAZo+Y7n6LqXGlX6f9QJ4GwrxwKh+4tGRwVIAk7almphf
RGZeaSzCGFAWEAvNL3KRydXFMXDu53/BV0Z1FjEfKVp3qwVL0py4jvEFohuxmC+7
1LZKwpPZnpxa5ITDnpgyt2vN4stZBpPD3jDWJzOpFjPxMumwvi2Inp9jY6fYUm7H
5p9wFntfCBPCs4lgiJAoZjp7mbb9XQs+Pomv9R6Sr1cZjz4xbqF19xBzfolEmfd9
SUaoCkXif4wp/BqKOnsxnQBJxfioINv/sNF6NAUPLDGqfFHim8SVUdr8yx3TBZ7r
T7nV5fA8sRtqeojT3GqR/hjifZG3P81xIIdckD2HwrEOb+OzKFtWUB8iC2LdIfL7
wup3uYQIQ9U+D0gL56O43fBHNuxnmLXYhT83wAJEIl8ZCRKCyN7+wV6b/8tOe35B
AEqSRSM3RbvUExFueb2z863JTieNimEFKHFidY/r3AIJ0X7mUn85XtTOZJRzPnjE
LvmDzt5ceGwrjAnrouV8WlphuCn6RiFCMAgbPLlOo4daCehOl69Y4EkNfHvcxZ2W
ndhyjTnsP3U0nThrzfgk9yryRRSusbgjfJVA4hJsGCADiyxqkggsmPYYio5NjLnL
e2Es0aqxh8Yh+0WPYTRfkSYEg8/5vvWCimBk6qMB7bqCk9VFXndlnlf8tY+e7CIU
pYr0nHbUTX9DANBfB0OCTaW/+2lmu26ttIaGdTghQ11rB9ak7T5PryKmaI9xzveD
mlH5kFzcIZO+Y3hkPMw6n572rqpSfD/bBwFlr+I7ICVsWyrdqYzimYKULBhB39Dd
Afv1zUqXerhRFckWMoDyA+fw4RlRiFbCi7sG2MKbtrgCYf+KNMmK76bbMqzXMiW5
FQ4lq9j9lC02HKAklMuBMArXvYd3fHRL2kjwZ4/pVqi6xC5fGPw/F83RV7Btys+O
e9YUR3Vf7XMxjdM/JmSPMb0+oHjE+1aQkRs1cylH2FhonTqbwBUvL9OqswERxQZ0
S+hlRaB/zqipJ0h3bxu3Cf7DRyIFbX442Y8mhNh1hCNokNCB4MzwybEJzNSOKJgR
dnzEaC9kbtKcHJqPfbxKQXEFHDAeeBPrLg8hDsFq0Z8KcPclm4+lXJbZIsVOJYeW
hsFCfgVWBI5HfKGCj+drpjwFpDz9tLURTWGQZkSga76Pz6wbMCeYTbwoqTlzAt6h
+unK6LfLIW6sc0HbekoZXX1VH36HUKPUb0rTV5uaanioq7xLcHiOl/S8g4s/HBCF
Vd8w80KCqdllH9N4cKrh7OyggS/HsLV2NYnD+3ugEGyPrZxVJ5iiUtKkGGZ7hfbK
OTGo1lTyv0oAXYkbsThhxglyw5bdsdGu3SWy/GHC7RG08l1pApqogfVoQPhhYGHS
qQkwNmE7QzdVzNOh/2hqcy/hq7cpBa9OtNxyAYNfa+MnPsMiTK89dJFZM8UtHaSR
5EmCQA02xDZp6uOc1yla3xaqse49HUC/V+NS3G90ei8Z9xqapN5sEtvXR1kCSvSt
DFh3665ZWKftYLLrVQH90ztqCMZTLjBdpmtyt0Sv9/pSNcfn1adO2pUZpVSwZP1w
Ozgh1W+MMJDefFGZFoqDfgV0yLMYLhg6/9zDet4rwp7JIyFNG1TqLWGSH3GbfoC7
3Rxxd19Si112GFfhFHA+hcNT+hUGHVY/mT7MhacNMkryy1L0N6kXmqyNLp1mMg/3
RY2qQ1WB4LnOBJplhnucDAiYkdNY609XsyF/XuKJnM8O4ZtVKO8cu7euBH810oRD
47ZpZWDAxrlx4sR4iWDwuq6fcTGMqksiPB3BtdC3lA9ocPIhE2ron/sxyBze04vs
VZhdSMzJADFjpuoJL0wpMkxTP1+z39X4UpjIZd/k6jmwaiamZKXMrsGaEMxuf7ld
uLI1jbHxUyt4U+Fqcsr3+qE/JfuRBJz0VHR8HrbU0iXEmQV96kvFs6BAQ2JkD/F8
m9G6v9r94QvjU561+PtSzpoaU810n/5q3Kfv2D+dCyo98ZHLRVYbt2xZd+0ETRX9
DYsRdCk+R+5K2Q4+3xW4RusNE7pSs92z2BtkKQQ5jpzz0pxcqrHl8VojcOsHMWiy
VkP50gwFFbkrOLVRZXqiN8OqkLRZHYQP2NOjhcDy3ops1chVUdLz9hkFue7yt92O
viWJiYSt2OBV8v8DQG4QJ89VrkTYNOmJPvNpHAHq9Cuz+8cPaWdMZSBOR5rk5Ww0
ZO0/yRhHWAsx8U/B6QOjSIYl70HnUKcdHfOkTBIloOcuGVnxZQ4IJw8/6iGuelIH
a1Wnokd76cVaIawqvTWAItc3d4sm88t6xLmyqqiEj+xafNzgy5DyeNgMHEOw6jYP
bNFRlZrKOVE3yMTNiE1XTwao53ItACwl9HOXJT84vYphnIiwtTD0vOmz4H6x/gZO
WezvWPaoAdGHqOWAmFUIqyaC99L0T5xsy1WWTOvQjKedP80Dw2ZCmJdxx3BT93bV
R5PGSBYIkpgmCxrbhu4An8GD8hDGa57HFJErhGEQFt5fJjrBHKi22p+QBZ2GSOIe
sKNHZNNmtay4isgz1Vi8k89mH6R5hzPOULIPQtyuk4GMDavSyktWbtj9ECsKiaDu
/19hLU1HXWhRAZANZ1OuRwFj+yI96IkXcZT2Ew1/snbPTxJ21fx7j+kKzIPZyUCC
7xCtO94L4H7miYFubnhMKcXggFR3nN8HrJNtKNvkATMq+JC1kHUVBa3A6biifnbG
Jc/dJMbl1lyXdOzY/XOqlSs886GUSZDE2SA3mpeOgrwjRONR9BAg5v1jSXkFg1g6
xhSPJwRv+LX/ZFnY5MG0jEHpMWCOb6J9u0NR/sSMzwVeQVJbl2PxwLafrx+I6/bb
sBNgVIhj1gpW+dWwNCRfMss72DPZtW8vLFJA+lANIS2F5LVMJA4FlTl7rOj5d73d
5PH0cfQt35Yigk2ZdjkSvGjIQeC1+sGAPKVfkJ/xrk3gbSffrd9GDQRKIoYGgN19
l5JJOkP7I1RA2WkvKc4L3cn7RLG2juqB6SqwSZ9/kaNgOkb31fC2e052mhFyIn3I
+YDJYwKIiujJnN4/rTRRPGTbMEDi9uCBwHvIuU852e2RW7dc1y2xT1/gDLdx2t1N
y0hU0pKDO04BxPzwNwiCvQ3k3fI5zO7WOF5jP/X4rf4hb2zmHDulQ5jie7/3NxcS
KeuVF+mEoVPJ+3u5d+Y0g6+Y7Vhufj+uyW/O4YOSdEEhrqa+jC0qqNeCGwYKgH6v
H2iCFjru2zFozLp4d9V4zuIyNQU7iq+rQFlhUkBNweP5WFZom0UVja0iOKDuK3R2
/5djCleSZPE1tpT2UmE6gx+PRc533ms6jI2e3OyFTiQ803VTMZycUDGzo59Quf9C
K6V2SzE9UdjFixVogD08U3aJ3+7CjP+9429ANRTDoO5w/VicAz86u/7fAFdPrLTw
w+qITtaTu7KyM+q1dgFJ9GhYqdxeC8oh9Nh5/oxE3zymP9000UoO2WB7FZHnvL2O
vT5yyZ+5MLa9FiTfcM4RGOdaYaCiGYtsQe953jnbveNCJHdM5tF070eUFCI3IBnA
aLCRbW/dsGbvyRWCIiIazo2XtOgAdpYNWQNWUG9ORsThiJUunp1xD7TK+YQovAwu
CrM0ZU6Tv9nWFkr0CnpjQZGAr5Msw71b3vbHqzX6kEyD/6aTvL6DyY5T6SvPtX1/
yzvz2q24O9gqqdY5GPmBoK30jW4CnAI53kljMvF6QfLyOxB7+rkVZgoFlDvuTrGG
6YRsvhpRPfS0MMitwlLf8jn2VNplJZWo6ZlLBsMEu/TouAEPpA2hQLmRBL2arF/5
IkJHU6lFHlVSWGULzR0fYNBSrYwEYLdFIV4l7A9kLq0ZxNChZ8t3mJuwBLrz73yr
sTlYKKfS4PFg8teE5VlWh4f7MhzMqWyuWEcvS2/m4YO6Z4RIImoAACnVw/lEKLt+
s/o6oPfcf7Nm29VFNwxZtx8XTBvgSLUmt9BINPCb69KokPPixyRcH+yT6voPnbLk
N5jHNaJUOP165z/F7RY0vPh0X3uN8LgO+e6hnsPIb3+S5hZGnLqUpnuv3joap2xn
aCA12Vtqmffrpdoqw5mJARZifEUR8uAwQfVjzRZHCuqU4pVmYldqiAp19zSZY608
gBTjZFzVVP4qweJcOoDCDgAZE9W/14GuPO8EIteV/kd32XN2/6VcmJ4nY13Fc4gm
CusfdmGvnJzd9lQGoFU+ykarfrwXVxlroIsjHnsA5sU26iGMqrt5TYQEyu3kBTwo
5WZHrNfe+47yj0XJBzWyiPSoaYFXAmIFWspXeeGuD/tUJdBror5EYsilAdcaS80C
CiiLEBsMu1bqlOf8/u/rgsENZhVO63lse5dnRJ1EmlpwMh+1kRXePTD3xo2n7zCe
2jaJam0sTFiQrZLp9LeFaR4ZDD7tsqjEJPOB+GQ6iLdlFkirNt9hHDd0r2GKDoUw
P0HdsPQlVOE6KiR+iFkdApoIfZcQMnM1iSRRnT/ndDBEc/b1KFCWKd9wZctA6jj/
7VoF14ijknoBX2bMMfw4NFXr/v5QUBzZCXF/pnZD9o/mEfAD1RdBZRKW7+arVzoD
uVa6Zpcb7wEOO0ET7ZSrB6Yt2EgBQvluOQk6uXwVza4lq6qNiPmCJ1ub9jrFWad/
uWSmWCQLg0Mk5Qa53UMqhO2XwSHeoqvL8D6IJbvPz3kDfbhRPr8Hygy3qmnZRusB
gW34+N6pOeLbiRNg9tZO0wCCaT+ImNGP52qXhlw/P7SP8NTS2e/oQTMvcIQLMuhN
fPmuv64NJe11BKE2fg5Bs9a7FcL+3punCOPHMWzLmjgEr+zSU8yCSJTX3p0m1ZOG
Lmf8vwkfc8GBxVIbAUNOlWg+wqfijmRZoS2h+AhoiltfQdkog5Qvf5uZzRRujvIr
F5UVZPW54OMYIxlMEllzbS6mhr+xDwK2MN2LulYfR+22V6NU151HiOWBqRl3PKSE
JTQy+1IG52G2A0gjQqBObwWIv11BusPy7ZkN0Bibm/VJgPoNS4K9fkZv08Wpzfei
KPSjN4TZOI9bas1bF2i0s3fdAw9186V8/ITUQRB/fUsTRwOm2V2Pd0r0yv2xk46G
siEJt62ehYU/0MTvUGm/Zfx60bC3DYuXrbQOPuhViMAUEdx5k48sOllIHFKkOiID
2d7KSySkXxwpIoZcAhyEYRLKebwWHYpQIE/a7ZgUnxNLo1EjcPJELhmmyovcTAt2
vZInVIb5+sCZSSOfZPJTPxTIN8TSSyqM0V64976Dck+6Q7QrPDYWF/3rnwKUWjXY
wwZo5Yd6wUPML0sqlAPFJUtfilWrIv6kqmTll7i4qXQR+1q0/6Q3m1XgfP6nDa7r
Tz5/SzUEBxM+/T3uTHRqsCuffEjr6TAwdsGSlYnDHJhzVr9XqNR3VcSGbxJPKVW8
jqX+cOokrGtoomBKw4xL5xSMnDuGQjoaEvRuS+5EE4GEfbyo0RsImR0mFilSQd1L
UvzMSlec32sas1xjnCpFRJpUG4IhjiJBWikBjAJqq69GMGygefgTCRdrgVNB/PZu
9JTsP3D8jQoz4EltGX9CbAGBBps+lGKmjkG0muSHnW50zy7fPPG/sMJNpUhFHzyd
OAxbmd56Z5oFPc3l8yW5jWCnfHf5fx4zUDMjT/6YoT/LHxnEwg5sf38fmo+jvnL2
Mbnp97y71WmHQ3JdIY/jpaOVqKFH/gU4ixexj+ymDHa/VNWRJL6r66iqyE6a8nhA
yKJm2OOkXAAST9kAn3jcUKdq55ohX3YSPVuNapinRWA98x9OT7ERt5/8eWFGcDuN
UKa6g0a3CiXmyTeli5N6joguxGd6cfSHkziX5tW5TwlwDNUsRsoHpvs84lQZD9hF
7zzaDRqUoapnjHQAI6fuw7bBpeeoIkjQdBr2m+CBQrWr65H/irrHG4TfcnhQZ8DF
nv8QgLPWId8E8h4YcyEt3xeB88P2f2opH2Gh3q+CxKfxjvg/40smkmpbXneYnPPY
3G34u20mfrD1QX5euvgP1o7fBeYHgPJ4NtDr1shEliZ5L3VoCgXb69eaN1ik5onp
6cUTRgCR1BhMhDQnjdDgnzYAMLarZlLAOk7OzfZVjUGQIo7WIqgAlroD0ggzfJYk
gO9iZUkTAf1rdczL6+D9uIpaulZpSVS4A6ldn3ixKNQkdwX0E5hlm/KYHF35mX4w
W3oTXbxi88623+tG2Dkz4MkPQHsXFz7eccyZXAzYVOnwRLffv4oYtV2ISc7HpzYL
OF52w60MrFqRQvivzLUfyLcjgsfOpYdqUV44c4Ep334oCWGnepjUFQWNz1qHFr8R
cnbYnlBUkNVXdrR12tRpz5K5pg73g8gl6XPrmwoHvR1M7dqsFB4Vo9JiPja7toYy
VUFeIN5Jwls5fddUKw2+atX6uvVMmzAp8bQOj0x2M5sRFfUM+iu4GLRKukVWtFFv
g4qVwzTLS2Ht4GxL+7VjHM0dX9JKyHJ9mhYT6CIv4TS6Aw6vAXXi/khX3rlJsue6
5P3Th80LWvhZ9URW/RU9JJI/8kuNNjzawHwFjET68zxgagZfMA3wy8sTWxC3mkuy
guH/V9RqyNzK42vpiEJ+plctoe/l7QUZ+ZHziwx59SiVoF5K790+JhCjHek3bzSs
5fNw30I5nm3fVcQ+sUfFbaG/H5iuGs4a7o1qmhZhS5U/FTCeRVOMC32UhVV8al1b
K8lcaJGOGgZuGQYq5YQz/xa7q0+9ltVUtlbcFkiwUDM/S1+DWgZz7kcOY+yeCUBU
/d6orhu3Q2+pCxp0ulAiR/g8Nkd6YEi/ExF5T4RWPDuLqXkKmZZudSaLqbnu2w2H
YM1Y798XlVbtY4iAeQKpJcdf+G+C+vOLDpW7wkUqqaTBgS+4f7xnjiZlGmwJRmP7
KMj1FoycrubOB2c/MAsyIlNjJSf8/eFWzVcNrJMZTcSuA5mOKqvokQL0l1X1MaEj
rJAjTEzk4GLk+4TgBhcnkneLJZJ8OAQY4kvpeWsbwzHhWhwQ/79b+5Nm7vLM4HKK
LAKOeXvFq6F5IZNo6d7G0M0beno+2cdy0YZeJjpTcZsVXnivHlAZ8JqaHxC22Atu
/E21wqPn8fGs50BlV094XymO3SMGb3hiUWul4iMeBxgpsPvim2HVhgluOvTu641b
haSBcPPp0asQAwJYhGc6xkWnglB0a+jGBl7Q18OOv32JAt2zieKQa5zKpIysuITW
n7cwlgPPhkTHkFTVAJe3fVTnCbluuOI/YUBOv3bzAqdPmLJlPuWqosRKTSTwd9Wy
Zst0TEQgtYBUYyg+J8xerrvOyb7i6ll2rR06WpmZB1vJLOffbeFqeZq8qEIw8JAy
clYezsUzspFIdtezmvjCcc9P9hHbH1zQ4e6otRRqAELiDSAPDmAnY5nqc/mZL68O
dCrVzaU++6wDYQ29nOh1cLUBEsUxJl+W/H9hT8JYvhVMF8rNYVerEMaGFKGdfT0W
Dhecn0BC2/tvIRjuyUym4lgAHUzROoVQG0wTVHj8J4X74kxzZY7tbTk2MbG1z2Va
Azdq3H3xjo20L2pzmHA0LGtOkzFMq3IlP/2tmc5aa7i9JYhJ/LYUQv7D2SfmM5/0
+12ZB2HwE0atxmXDpeblPC01e36wsmRG3ixbCRs2L9Xp0Y85pi+6Vyhq7B8Kj0ai
Wo6/e1ZgWz/ZEP/TFtBUlmvv1L+aJWQNLR0CyIQ34ppI23eC0p2tVOxZU2VRcA3c
kv/5roTFhLwKPxu+zcd1mPCO7u3cCzJvkh+E3FKcmI4533uakfrsqwRimGqSKVQH
0Sm//NvN5hXU7VY2qmIZ/ah/G6Tqj1Pux1WR7LVe2QQoKQI3KC6r/ftMCJS9hQPI
/8E+Z/cZY3yDY56prYJdGDJEsAmhhkZARueU2Z7XNQOKU2DVfIhpKik4yuZGEGIk
ezvNAG20Z5hTOW6CyzCIkxF3ia9rCoyRk+iD7jqRpOjSeAkSEq2WrfoW4SJ1asN1
FipnZYyjEJvTUV6jZ7UlbSHUhJYzyxqgwHtnnPW/gfBUtxd3MWzEOV6CTwE7ZYk7
jiW1lM2KnYbdgZX0qPBMx5kieozMEYrZnz5mb+90Pd5xKvZmmrJhfqNBwLECsYUd
7f0fRggoaRKs5lt46QLIXIo+zj82CezN2ZQh0cVHpttpB0rLaVIrWaFKcxQwfCj7
hRcOciYXUQHEamhJubWuQqVXMQ9YsUTD4WQB29BNs4OMP1f5//iiVZpQhWj4te3g
nMImnIA8HWX1wCB2xVfbHvmoVenga5sE0VyzS8UtPXW/4wrp+RL+FIPKPzfvEuFO
pJbcx/+K9x3GTuIWYP7YAGdNupcbPoShKr/MFvUwaSOfvVjJVj5gOs7jfeGktGIR
TvKm8Ur+B1Bb5HkSsi8mwsJMaBIF2w07gAS73yhqRIPUPFUD58gK30XL4jafwJf0
KG46Gi2BHiBrXpiYLjlqhlx30sRsjAZMvDgbhHrjdzJhrEyPTrm1J0Mb/8ZdiDEn
gTtg1TV9XwscmhlRCnxIC61rCnOXV0KG/oRyBfK2IqD3rS7NfvZMr3bp7314YPG4
l9ga6TdfhLn1+nxG8RHFjYZae1OaFf/z249fZLZcWo2apCoS2JZebcRpSC41gaLZ
14v6LUAsflfEfi0KNJtihtbiCtZwSNYHPMk1GTjYd8g4jZrY4XLH8Iy/GHXn1rNz
mFG18yLdqKdd645gQXAOcQyl0GamsKrgrhN07HFdeeMnix6tl71bRWy5Bsf5O8jb
Z+aGI1cEq+17sDGPPqKJtkbef2ydZTmmMT1pu4FRKV+jLMLqHSRJ/JP+VNEVNF/v
WjzBz1wZuR1yl9/50eBREtChDQGAVn3C1nuwy8RW2IrMP7procZQQPJ8v3dt7ipi
Su54EqmmE1IBFNOhj8OwG9Xz9VYYHqkA/X8oDmK4ET7Bq5x3zpxb/WRuECVyGyz7
73Mio1nuAVyGOG+q5KPTIwPJHn9Hz/4qqri4EoTwqZIEb4gWNOULKKvSqX74MqTA
bTkPVkj3VjiZm03WTeSkreY37IcPu2kRlghZgh94dhYQJKIacA59NV7bpsu/8D3t
kSDR9u8ufrubUq97IG+Ty0Ewrd6bRkEhoip0bBT/jAbiCZJR0v247L67zASVm8K7
+SBiaDGa0OFHsLyq8DaGdq2fxgv0Z43tYyGMjHHYJVk2s6Wt8OiPjyuA7e/Uxktw
ihHBgSGILz+7D8nhj27O1tBQn1aJcp3s5XdyJ/WJOSOcbZnD0IrdWHNPRDNURoQK
rLGb6VYdsV+D0N0wAIHyTaK8bVevZprC5yUDnPmMItjWYMEamHVF5SoYO44CRyBk
50/X7Fwh9IhgsoGH4mllJPyuxSNXtE1IiqY5N/BELl8uCbapem103PPaFMcvHimi
sj+Rdfpw64ar9sFknDDVLnAdi4AsV14GpDhm4ihqz/3qdvrwFBEL7RyVk1iMaF3L
pTN6hSANqcpma3ffULcuIUsByCon9oDZykj+jhCSOqUvkS2IXdiKeZllPLaw7PsM
kW6OWyCLayB8EXUm/5sWDNuwdokOBIrmEDJu6qO7poSNKajqQ0RFfnX5WKMEGMQZ
RtjVjshDE64Q07BrzTuIXzmYhSRwFTovnJTUsrhhL9GaBb49zLTEgxsXCEXk0d4r
ibbpRN7PA9WHaygIU+IRkh2DcXVjMUZ6MgRd8kXmTQTSO7KWR2jQDLEofXlIOXQd
tL2FbN/8cyJz+qZORx9pkQEP+pEgYYLuleNs/3izPQdP72Fk8odwAmL95ZgwEkAp
ldW6sSZyyuvDNVo9FN7Tyhe7kODd5G5JROoBOjA6BmSXe7LAz6zXLhvBUsZRukUb
O/KDLnKT3m1UcSunzhN8qSdimMTq4ulas4DzT7yOnf0CEGWTloUWYheUZUn+0a/w
uDQE4y8HnKAMKhlF93n4Klzdz/5JBTuuS11B0pX/OMmAwIyX7YfkE1lFzo4xr2Dn
l3XOfcaf5Eo0S0mfWAlVWRTgp8YdsOIhgC/kJtz3P1OGTSepI0Ir9/wHyw9mIXUK
Uolc6ydrFKn4xJ+/FwSYAmHe3VN7IkCz3HpJpxNfQRlN2rE5YzvsHcyKQHaelqPZ
OErK5SaznOHpx9PfRuqlGi0mtMVQjCnSbZMzaJ21wKVkkfFlthSxhGE0ab2mliEk
LV208ymztCSYQ/nIU/gtm5wAaRcJ6UgFQ0BnB7yhvQQhLu8j6SJO6AjWOwHu1zEu
jFvs17MYvwG+zharWvAybGHfKU1ePtuppbxJ/5LA0aU4M1JeP3gOeVETHwlTo/yX
sB5dMVoHPyaFKVs9Sn2hsx16z2Wk0SyBIcmuUOlDwGgzQF4h8xZvJVMcJQlktsQe
ybrx9jK+iaA/7JEXJQ5PkTRPXYoYczTPYEPuiTkkYUHiMXVXuBLsUG06ajd2XD0x
/Do7X+GIqdFlaQMKI/yGU4AM82n5wgGoPFzi6F1LX5RZHp9nmqKvgK0oogcO03Yd
2tkj19B3ib0Qhp9M1JHeHXbS6ni7PLMrjnL0Pq7YTWBS6T4tFegbdhUj8Dho+ZY4
pQjdbQcq0VGOAzvL+IRc5Qxzd86OsHabBPbJLwe0Hcqf1mYfJcfOXfCeS7cjovFv
7HMwd8uobAFZLN5DQUxE8RZd1838zQ5lz8EJKpulfWuoEbTVdzirQXuD6UYFOedP
SHXBJ3cEjxebzxqFEoj7pdp93R49DwPwWEvMk3DKdvrTqQ2Ou5j29TmTyUiM8V6k
b/OH0HKUhLEB9tdZHt8861B4OpwGKGKVkhQLFQle4p8rKJq/gUcLwHfPNSM1W9eN
Y7vDxMtVMPDuVV2qLgKPY6eVexqrgx3t5F5wKWgbZmP5XmWUCRh6cOPCEzV7hNP5
AVwFhtkONJb/e/3y9CYk+isZTB8v3B5hEvEzLcsWjptsfKR1iFlZ/IbuWGPmnef4
3PcW8TftJx+5eCaCkWF/AYoiSoferpEncz60Zpp3lwHmNlMFCmV9Gahq32EsxXsb
Mb2yhhdA8zHeRx2Gxi9s8df7Hcl7XzC8J2vXCWdHjYxsEqgOyJgHmlgxFbm4yD7v
aQ6dtjEis8zSkDPCPLi/JYHIJK1kx1+YSZ97pnQhdGFLilF4LrqF+g97GqIr72Be
seaM7pSVLi0DnWdDc3rK+QV7uSMXScykLgsXrQRwDpSnUa0KGilQLvq/2R1H4Kv7
+c50u/Gt0bb/ayVPjgqmDU878LcLVg+iXvfjElj5EE3DqqmSqQiWQP3B0CdQctz+
cLMd1Lvrf/VBIoyWuT2sFDTaBB157ZHl4kosw+A7WtJvxpxKTD0HYulGPrEBqt3z
dpWe2XWtpn+kZ7I1xs1pCt0yNou0479GYfr6mEbnSEUeG7eQs2aYZl7AmnAJxnIN
htRDpDXjtkZo9ITj3j39o2IE+SPNDa/Hd23MqaiNTfTjaJRE7Hj3N0InvaOY7QTy
hLxe0KfMdhe6mcKFR4szv1tRwpUbt0g1+R3L773rfs+D/1iSDu2fJbxuTJ9gTSJl
CECv82b//g9mQ4B5+M3XSu8M1B6zgjKKObpJIN/YfMS/WC+uDy1AeZxCj6rzJVBB
AEh7+k8b4U2nkqKLd8G4l4OZqmibvWI5bwjknq6mfFj7r6tYadRe9qzjaKI6eJw7
b5TGSkmulRCn0kPWD4b1ZV3eo0t5OUY9p3Gb7YRuS6Rt160HMHkUSFfZyHwWb01E
BCmeoqrncosO6gyh/RPUZetg/dbjGCGrV+kMCOUFqmz6nfWfd+sqQyVghRoQfX/Y
mbKsUIBbnoqHtlsgpKqw99xEzaDqoIGV9XqSW8o9x9zn8RYe29Y921kpK4jAOfvE
76l4cQmKG3+caVe8O/BP++3PDnBigIMS4qA1B/y9Wt/JtroPsaJs/z3PI4aCNPai
IqGDPGqpwy2U5cffyLv+4h2DNfS4plOiW1C/L2W8H6BDSrqQyVCVo8CW5umakMAf
33hz+wP+BKDKGOYbMaj9PERCMLGP2Schlysb5ABHT0vcYY0oOdqx5YvOEbng8fVr
GNRUwQZYJ955l1FDnoga4/9rOXo51fVNrwjUm4I6Gt8YyrAlLBeU+D6AUUze1Y98
bY7xCb2XTJWcE96ZcIuXpPZ6hF6w1H7I6ZPEpwIxbLAfsodDw8PEc4nMWPAkQjDm
YbBFxM/fg2SgRQ5Eh+tKkG/RNXrnl0LbQiJpDOm5Q7UegXCshMW1qY/emhujmjbF
uBSSG3OuyG1igY4Yis8zc/0wJnVJNWg3/ruCqjbJisi9BjJZ0UN4UVIgLneR5r0Z
v7BPL4xjAQyqGV/ajdLtk4uXfv2j2LlsYDCdBrRqtyqHZPng8YydVQ7z9EMO6C6P
q4KN3iUcz7L9wM+0o1Kx48KmuckCteyJTofsGPfQI5FY06CX8CgEXh+LDDM1lxG6
/CVQCIExNHe1CP+OGqstzYLddkpFonm9gz++SVFlqpTAHSxhM6v05To9IcDS4USM
Dqr4ThMr8gkQPilxfo5SaJcvXignGj0WfA47vwJntddANqltt64SafO9al38WLwn
pFMkOtttMnNXQZBelShGOOhfdbRrEXLM5FdMEMEOSMPxoeLYX9D9SY+jYU0btYGA
R6NQbnL3rzpihIoRlX2W2vs6cX6t7KqM8kQIYDigAb9oetKlaFLfSIeegwQ56ODb
sTjgvVetifrg0Zbdd/q8RHHj6QpNRo2nMGtgLXn/5aB25LNDi/pg9NvaeZlmiVvN
ggSKzRJCqPsdBtIVuUra310CSuyb/22Whmq5Mt6Hny87iSrI0B6OEESweldoqRX+
F7vu9n0sHPHX5g4Td0DYBvl+PtgqIQZ3k3xF8/xcQdklK6jdy4Uh5YLGGW5GkO8G
2YbwMkNL5ld+q+GD5VtU8YLOFP7cwHJancuhIX4Uxus1zsUn1XnE1dVVql8aCJvP
Ozj52bX2+QismFShtttwXw3OthKmBNfSo6e0uqA0EWnYcn6JmQKCNV5KPA0bTy/b
ba2GgiJH5sh9beZJWlSTgxleoZUDX0p5pq9xNLGGdk5KCOWt8HiCIZp4kvQ81Q/d
sECfCEDyL0n/BgtpvrqSQKJRxEaRTdBUx94EVo8njhAoW09R7km5nKGGXSgPB9ro
o5roqOm71deOwMgf1cRP62NOCJmEjZUmFZ6OJS2wSpfPTeW8E69XcqGe+BgC80aT
4ubwThVDK+AujKS+JiEaGeFXiix9tyksmyz5ATZC/DBuvL0xY9iP7fwkuFxNb6sR
VeiVRD4tEaKv2X2qyCRa8RnM05UW9jx1f9lPljOtFppYDlbwEMyKsHgA7r4I8HFB
aAItG1nr5KRG1BzUzSJu4oCJzdMTOTcbMrGrqmoTJ3Zc3PeaHTSgJaegOiozUnmZ
0l7h9zijloRfKKeMDeeQP+NCjik+8EpHV/VIJ6pw3lK/M1hPKZav6dmbYejHV35w
jhXIW5QGrCoVYCD159R7PNT5iB32o0ja/9zVupPk4AB6GTV5FKRzXHn3Faj8pnPB
qPImxitmP2mFawV8LOTqKmBWbbnG7jXxtUQX5nV2orzIZ84IQcJ0PIrpIJ3kJO1u
8cuILFRjR3YAae3o9sLsMS0LXNC19Aj3Ouq9O1kadZTfhASwsE4rlNsWEbROYuwB
nvIdj+jLau8sdkwkF9nqQnAMgFj6XTsYkLORzbuIhQIfbsLLjUHPsUGvQJFz9+iL
hFHxceIZwE5WQyVnVnTiAoAy6Ydnv2hDjkWLWDea5Vx+R4MaVnkut/jqN/8iDMrx
y99QwQhwUwChCiA+/CZF2I+5Qw8W49Cah9EHJIvjIx1esi6ZyakEiyntO1yU/+3W
ORZAM3TB/IX0OCwT7tKZesMW7rvMvQXHnwkNAQFN5RWH88y6KnqE9mj11ozxTmgE
++4CHl07yeAbSgs4rxscrzIu6AuoFFopNQ0QM43Gwg4Vxt6cxVtuANFr7zJVH+ZE
pytRZtanW7DbWu7OOORGft4R5poA+ha5GWaqwasMWX0hVbVm93JRCExYYXRGaWQ0
+t37l+Oz5b+TsFBSx26IJZTQTvyPXF/ohvj6KMR2WtMmMLkEeuXpJsqn9sAxvygY
nlCJ76+0wVzliHfQapWk25jm7YsBMt+Ga5WBLeIJMs8l0WrdrTc6qdfUiACi/fg3
An4mkwrqG1JWuCLz820S+TbTyIYet3YD1QeDeHeMua1pECmJSYXowcSixIPvf6SU
Dc7iz8bbIOR+v+Vlno4oOoHeTft0059gZFfZukx2meGWMMcDfTiYfcLbworTAVmI
gir5PGe6EeUeZVW/HCojF5uxs9Xk2cwebUlOEL1VsKIPnqKD3HhdEIUvG1J5OwgF
xyTme5BmzjTISMk7eWmyO08KSs5tsC0W2s4cRLzlZGROGV9XIfBLTJ55x0wpmRAO
XQma7C6ktCaAZX36da0hlXsxif/yewA36wUKKz/E2Fp8pElaKdOBjRWK0BGT/FUr
CbgUmPb6SimpKJbQF2D189IJRHNyaTE0W2gLBhj8E3p0VgL1ao5/Vc/6gjbFTo5o
oB5jrKkry8O0YC5hZgrv++/QJkNUxQt4FaAMlJ8pSYqCfX/P/XroF/71rKTKC5zg
p1jHDcLG+ht7Wh1FN+xYcmBqWZoh/a6zpHGraTAHzhjitjE+40ND8JELAv1slODU
zKy1UJ8xN2+l9Mt7GT4K/NRef+mpGGJx4kCKsafsyro6GrCqS1GZMagzAFw94ihH
1T5q83jERmcGOOaamamG1aXXLPRXPFdy0xYRtdPA6yVtOV62yEK30OBTngj6gBqm
xznPTx4I+8igG3aObcKhG6rnKrYqmabVI6vfeLThQqYQWB1sgdDnARI9W09HO29i
ILeKkVw82hzAEQKdpL/6wH17VUD9dpCQK+jNnhJIHFnJO82MgLg16aU/4peexy51
92/srV0tWm3Nvsh7dCnMIlHCXP8lE6PUFCHqrJQFXRpDe0Kk3Kcw3R1DHn40C+MR
/IccAVbw1alEdGOvMiBnZKlYE339AGxX1mpv/ghYyrFalLBp+c6XoRJltbrD5KRX
MGRwsrq3hVsKQiQeL27fVqBnWYOOvBV4w3mg0GAGGYxNmzQ1OR10Z+CvWao8luXf
TeRFZu3vPckEbcOF84jz35BGoFJ6ihbngykAxvfyyDUC5QgQDuN99s0EDV8q5run
UmtyJjo5TstzK8589kypHl1jAgxHMmZpkJD7o2YerWPMUO/WXKUN5kk3jlxyafjK
ux7lcNp5yBA4+9qNoyJFkDS4VeNE6gN/GXTy1sqCJClXx2GKfAhGqiIvu3EcQfwg
KGTaktthtwVwllkxubvYARpeXvvVFT5yacANApJFnvs6fNjXsC0azKba6WHnf25a
Gj1Khszx9naxJM/FBL5vZsguAaVaDAl/qpOPoAfunfhKlJrnJ55Ljdce8U+HS/tG
P8iCpjmU26Q85yzY6HfQ8rBL/f+JgMSFPqWvtfAE/l/i+zaM7nlYSj/0KeoHRwYZ
o0LSnBC8A0lKX/5yDFmsvUneyF5B5f4Y3Z3iwfWUOxR0wtmj33Av3dr3pPZ+PZWL
FBVP0cs6yB0lIDzr6VD2bQkFFepFEganX5kHxhjROd7RZtpXmGSCQ83jCFZQZ6fp
2rZk3UNNqKhAWz6VvzQl/PYpLCILpAqgxOh7F/m+fP9/WrjYMR8UsjBEofFSKgjd
dYlIQ8nun8A1jx5AYeyf6npVZvg/kfRCwXrT5cBkCMss+LKg7oMTLXgeMYGvvyp9
UGPg1d/Fs/yaEhCE/JaM0hwcjTSv2llofRnr0piYCk/ZYiiVrF8FAu3Gr03h8ls4
gKmZgzzq/+p5wduJK6Jj6blbLNMC30Lf0ihyHX5+lgy+w87PNRrJyNLGPZIOW2y9
2i186GA4EH+04R1j3EasmO41X+5+JGeDTMd2aRLmEKRQtNKHdHAsMJvTIMrHXN/P
vCBMA1LxZsoNYvz3gxu+3x+2LE8t6CgEVG8raGTznVtT3kpqdmBYxPRFgibvM1Jy
js4q4WM+JhK+Je6DvmPK/JLEUkx/mVtLTVy39wKJyNGQhN1Rj/p5rmQNuCXajaah
fA1wAcj8ksoOaTzZIDkrKOinJR/mMV81xKtoBbg574xcVI//tYOwjlzPVDfiXHy4
1pqhC/CGhBQAs385j+5hvU61KiK3hXbpQNuwL9RC0Ma9cFLFBUNjfmwp6LAvmuNM
UAqgQYh5IaVsgID0og/qAYyjVMFISfzVh/D7XyaOBc/tykrcUDF/7E4NUhKJSIeq
YpKyUQ0abwSWost3DN9GjHCy/Wd6kh1/GYQig9zI+ZuhsJUJQAqbOPRr8vbMaQcX
er9jightVOOLDtd6wOMxfUhUomMW68B1IqByZvQmWAOd1SjiLWEW9FLD5B6eIbZp
mLxe1QEWjrwJVPT4jwZVBOiTqlOCaiJXFWKbgtf1QB6EgiOdbWY7dcKewVOFbjpo
EaPI10/Bn+pqEURsnmWs3qJxJ9GezFsT+BaT81ALvtvKJdTRHy/lMPOFPBJ/cHT3
evhnkfkPLIi9honY9zv7r94B30KyFv2YYpnSM9iGQUOQE0Wlf+24sd78N3fNdg/L
GBnS5ENGcqW+Wsy1eBU+L5Dc8ZPNqg6ivrYZ6TjgCPjOYMYmFvpb66Nktxb50Rq1
ot4XBSqqhuIRDMYm52uA7iuxaBp6zhdU9T4nFy9Dcx/c1EedMmT4aH66WqmTKEAG
Sci4XrHzZ+6CzCIiSqR1zlQfWz7B24YfAea3wLPglQWPsBUtuI7OeE4kbkyLwQ0/
qDfpVFiNsJKHeTwHWaES5LdBkf83IPjJ3s+8hA1K8X5e/Dlfu2fhsOgyNPh9+dQ6
fh4dRMLk1g5beBz9q0+HL4dDL7TtspDoTLM33WnIwocoru0Beye3lBPTTktvzRY0
rEZaZeD0zVNerBYOWZr0OdL+JSxI5rW2UCGeVbLyUGg0Vmlc8eP2ztXwfghweGsV
qM8NFcYbiF5O/blOfj4o/4ha6KkrcpRoikU0pEwbB5h8tN0oVoIpuDVSGS8TqzXi
xtQWoK8l9LKnAMz4TIXJeHOZX+L1nlgCx9D179qYHgMTbQqL5U7He+wfhxbCk7lq
s4s+kEoJ5KokJv9QIOmEeXR6gQe3uS3QrCALJzxTMBIh3xDNo7QAGJqo03IkOGOx
VdkaoIQ+R2ZSv3a1jFTSGRKL22Wd7nObBVilRJ7QI/j5kmV80gZIPg+e7uzWwdnU
6AEaVMnWImPuentVFL0OfOe1gyOH9MMDEkfoECTPHTWcnMQahd+u2hhOyOwmgK8c
tmm4Vm0QFK6pJL0bnsJnVyw+1hP4ktOkRZBktH9Slsnd7L0DMDqvCQpUiXEb2DTM
aPhac0oMzH6qbinS6W+pliIIdNOpFjnXcP+XpAzxoGG4V9lJrtlDyYH+OCG+gJrO
15kFI8VRoz1wprJzLwToa1HN2eBiPxnYkdefy3DIK6hfqsqorgRbtDhvyrCeEie/
eU30RDooZLxkWTwaZowNFLh2DWvw0acf+dTULrw+/Jei06QpqbKIPHJorsC74Zeg
L6F9m5OYphXLrhJecXHaPePW4KsJx6gxsNuVlwgaFMAOo25pHQoIJzBVBHjeiCaX
AFRC2/cAFl/SIRmTYmH9jKLJwFUHsVw+rg+6W3r+5HOoiKWZT3loKMox8NVKEPif
XizXUnoUyc5uEoKTY0NqyZNY6e+gZ6VTL8R6UxVFtFU9BcL7QjcZFhFu8/P4GTL5
WC7pL8+KBKoq1Ayd2LNgYUYdH1JqlTkzvb/nPiU9cJcbGVPinOQzLuVakOjYh/Wo
1mHRjJbS9HTsycJ0G+oNgXYd2gjra5Tb8FOhevXqGFxzfmPeNSQzzW7RlpDddQzj
wGO2YCuuZei5N9yXfB9lIIuI/rETPlCGCvnjevUC+oOnccAX7OMq4BbD+JvNtJFc
YsLWucB/jC0NbZLd8uslxbNSW+jw0nhcaaNeb/L7n4zQ1jCTTKzBJpEPgPiVdLcS
fnp9GuatOE49JthoWzzc5WZ0TmJw8sUxFCdHok99gT4iChCkxGI2WBIrhshvZmdR
UckQUUgLTtY+jFD55Mh/L2j6CbErddC9jeAOcLZI6gDFWAHo84YdUQLaLZm8Ofk1
pfCGVYGd2Yngp9OsAd/k1c0bgSIpwRmzV6YstGh0tt1ZSmjzqgoakSZy1q3a6XY2
y2dx2uPXsCkk7CnJJSzfzB6ubd4dvarQDZpZAQ2IadbxVcIlHxJjWYhriVf6W3r+
y/6H5rWjrS/q4BshO84Rc8fDvloV6sn+y2ZGO9e2ONWEgSWnnTzsZ+cMRzHm9kgo
4x2sOdt3dgka93Y/45FxNcDu4+PEwiMIXMk9yHhTl/7qLcodQoQeCHHgq6Tc7VWD
gk5Ysy22KTBf1Zsd+gSbcLlK6rR481VT63Si51Tf7u8dBSFozrjjYGbudIayaqRJ
ZPchKO4pyrR+lWPeRLfYBZ+zT9hSERMkvYdduNsspJOhF1PPMicdxlJqjJlKGFuA
xjnMxCD1I1KO+IJ0mVsiU7tXn/BOlm7VG4FUxPf1Tx3jPk8FcEO832YfTt5LgEeQ
4JaUnrJd03Ysr3t8XP36eSFz76wNzarTKT6EnBbnsKuUpDo1w5KyTsr/xypyClr8
PS4Ki+3z4WaxfrKpjquFR+Ny0vYIgUtUpOCyDerFiD/+uFWSuEgs1LKVgKP+jyLK
EEmungxHQ2/UOjsw5FkjXLm1+6s7tKl0E15qwE/yjZWixyJbTkXdEL0fvDg/PFp5
JGANwJEg2WLysfoWS7giq6BVEbmrOjcfyoYEyUDGXmKCuhAbU/t+psMZ2g1xP7Z/
xIHgrKRjzOTKFu0FAjOvfL7KvFz4vX0YnKgsDNvvwX29SimZg8Di+RITkNyjqhrd
r4KYMQPq2jW8v6aAHS96Mt/sd3oLAkuyi2YE1/Qoo3Efu83hSSyVcuET5acJkmIc
DSrHx+ovSfqjmjeAKQHwhCLATV7s1Uq7ixW4aZIO8tkEwWM0Q5ZrHuvHhwaslaAj
0e/VEDvCylDxZA5HU59gsTq6uysWN/f9c5RAui/1+RFUbcKvF26b9wUtKVXdmIZs
5RcHX020ktWU8WFp5ZDD3FoSWraGVzsElOJ13wf8tCTgfsLsf29QQPZLPjnOTlmu
qXajZw8XIF5gg+aGm08inrod+TTXYhKXqsabWp4rf/6Po0Gq/tZs81fHdEGvbFhF
wlYZgzeE4BXEh7ZA3P8VDsSpFoMauX0tRnexY8a0VtzwGg8/9S6Eg273tZnCHFGz
BNdigi5mTu2VcsrXjaremBcvVqel7d0gQqBd8tUsD+RNEdbq8B4rgtMY8QaNpAIU
Dol9WvpgMHo4fHmmnDG6VjTUcGBtuzOy5qWHRlnmmoVBfpXH95UfKfMdcT0s9JE6
gMaRXSIgvo/4w9Ma6/KW5UZyH6BOwMKQS6YpVWq1gr17WjFgmGrvfXeuIRU5DA6i
W254GcuBrtlE8Pta1iEUUquTWXAtoYWc7dFEe23+BLCUb3o5ntMLQ1MJ49JS5/ky
qryfKszJTAUnG8GpjIW3yJFR7mfVbBAiqWsFMZRC5+P3G0ri/ZgfniPDqnyD4rS+
el/Cw9oYeLLm/rXzqv+byobeGUeW6+/46EiOIfE/K6R6qxYZI+GTFh+OzJTqwgey
pVSogfUXy9LO+yY30HX5krGf+6i8Lc2qV873W13wYuIhq54kr7GBS8dFjeSIB7Yc
mAc78rUl/qxCSrLbJgR7Zh+TX6rzdlDrGS3CxDlWyJu5cZGrz2SaEEqo7J0m6AJR
DyJFCtHv1E0TYLqXZPWkChvWagB60d6M1A7QrfQgq2x8kjUtSHjlqrMGfcm8po+S
8DrrIyluHBx4lvy/KCeGIekTtimBU5ZNBu/EW6sTtNc/28jeh2hNv59ssO7mbFzg
vkjj7E1f/kFkqKy5h4W32b/+pjjwoB7yNUdo5yAvG+9q/95ms4lkHf0w6pM9HVHW
6CZQnXCV2aK7jXnwgxWG1wmmA+3CzpO6VpFCmZanwdTI7VWRmm4uTiMRyuGSXYTr
iPUWwwqfRJDfFqrZcCwo9jsiQcOe1VeKnjEvB3o0vF/p9MmAKTvFTz4uRjE1SLd/
o2ZYkNk/5KAjZ7+t0qSfG90e+OX8zEjEuhZThiD1lgxd6j64YHh6vIBBzL3Rd3IN
RsTem6IC09CO1eO0i1UUiMt4mIcq+mnPXETZd7+HwzIHFv8vVFBWe6Xx8wPx5Q2u
pXUs8mXgslgvVMWC5UzDpXgOmB6ErmMCOp83dIVrVJ+riQl+zy2sGaSrb07WCkJG
ZVG1vRCBxHmkCG5wmWx9VEGbVTK1PR2i4W+pYIf8THHLolkuyfOoWT2HsYABr0Rt
k5YLii/P1jOhLnawCdqc0xCTXRgmFaSRqPtjX51tY71IQKAmLVw2BQ0BzWfq2Rf2
HsYuQ8XQqgpEJA4qRQ1+ZSoYGdFDH8ecMHEE4JcGypw63eSCGelrCQX8VVDGtPW9
9nFHIuZZY6jgNl1mhYl9L4hlFCxZCgAElQOQX2QTio3yPx6h0lkmr3Hfhdjr+3tQ
5gq/9jvLoId4V7JdgwtJfUcBc2GnKmvgJXw32uVXsD3DRahFpl/almKbA7AqIJtI
/Y7WzOwcEFHm0GgmdcRk/WIYSWs6hbi9whETgJ5XeoJZCMsgGSiVEDHsgj5/9sbK
WU0PBeKqdJhLLFwsvcXJV3Dlg9xPypuwbOhoDMIizgBKBQ60AoVoznHcqAjxvyHh
kPbBqH6jDVCpNaOok2JsmzERad4Lc7TJTCq2hW2U/lRgux+5c1CN1yUvfx/v/1rm
nDlIorjaA7pG5PvfdiKy08Owlstrq4C6BiBTJFjS7dZilvHGmazoJmKWCW4OaMnD
GwNS3Uubd8V7VJN5Od6NWRrGu6qFB02p3PmjitPtpRQwSpf5uinD2MFfHj+p0JPF
it/Pd+57slbAukG47/a0tml7mCYawaCMk5WowBM0edEmkUnrrCHWOmfVXu3OmDde
8rN/jlSjLRwjt9riJTlVbBLKVDJHnowKCLu0CFmjrAspe1LSUIuzwa16AnhPinoU
B9AlS1lF2kwclBKzUKA7AdXT5eHlJkxhLBWsNPivmz3qfl54d5xRmI5U9F3bZXb/
j6l302imUCWUBOWfuYsqAjyuNapfsIoAY07ritKelLoR15dAPG19SVS6scTRZzwH
2mZc3s0Igy6IT5Kl7dxiW/xXKKZ2dcxCoINyoioYO2bqADRf2U+jpGz4NPAWAzKq
19N/U2r8Glm2+Wj9j9kE301ZQIFhLUJfUliDYN74JxGHnVqayXnrZzLNwuNAwZ/r
Ku0QxJqwqDlndMFhx8pRGi6YdzalylkwIjvqitlNFfa1STTfqBV14yi528m9HrEo
IF8etAHVWpCNXCAwEMi2KWNbCQhkdMIXnMvBYfG1iD167U755XtaowzRp/G1jQIW
kqnaNLz6V3c3u34b+KEb4/6f6JWF5Y2q8jvToHgPzK0S+5J8tRh5+YJhL8nAEhmn
T8sdeZS302X2L6auCuo8IeiAme8VzNRrzfe0YsQ2NL/VjI5zFh0q67OZG6Vs3uHJ
DNbeN0A5u95YRLAtd4Z9f4I1klSj9vpU2BGS73/u+TMrJvqsC6CiDVB0+PEYIimg
Pd4lK8Go8Iq9IPWGMSW2IpCHR+/X2DoysCL/L3mprCsH9zU5eG8Ij1QWEo8Okp6c
CNOOLJ9xmgeVRDWCj59WOQRW1NAsDGnG0A9tvTbCj1UzEj2hpCTWg7+33MjL83xj
jVA33poRXM2q/6y6pEAWdoS/5dVDuC7vnldiQDRJXIlMQ3QtkUUy5L9vfImj3AVA
1Sb5pm1ssufAMtpEzVd48khHe5oWpiJpaxrqOr0N7TUHzmk9eRe7jfTCG+w7TDDL
qu2r9gKYn0cHSlgqbVOdT2PdGlW04QU2hT3gRoQFGJSb4q9QEISXHqMmlLSYTw3w
J7fAnZGENE+N6KOEnS1RymToMXnOJirC+22U2FAAfurnrqIkEcTN57jMHmTVlfEd
5ot803ETukLk4fi/6wu5V0Gh3ZDm43MAXjC/zkN4C8DHu600v6ecJhtxwDbxcabY
nv7W4BzOTp/Uv7dE4C+qDSfh0RzrmooTTRog3x94vj9fi7l+N20PrHGn/YrQwtf2
eHYZX6gxLYNQOs5rO+JRVpD3XmqQytNJQF2FDrMSZLnIJKR3Z/7v3jc6gEuQWO2y
ROX9Fyk3yHztFrw18DooPuNMyKk3MKJMrIz2IibWf234orYOf34aZ0G3HhItML9p
u3LlWBvGY4tjwgi0nahrzhJcYkWww1rPTGwrbppZE8Ohx4cGb+xkdzXYhIvLLu5l
AoroVLxvYNIKU75JUr25OY1CmAwHSRIBh17M5TD3CXnMneW87TqJlqFNsG40hOn5
lYru3e6tRfMIa+0gJmEdrMMQ9MPQOpzs3C6006aNjVzCaz4bEwY6UkwYyWdag5Hg
fCjxWaGsWVPvxHEpf8IALb+TepsiVAlHbV49wMxqSRPvyOJAag+iOQu5DtWe5ZJz
BTmK4zIWbYCqirG44Ad20BA/iMoLUnMivqkP498KcBQFj/150kjJyp/VSJwGJqi7
WR/paSZmRJGRx8eKGprfeyYn0BLqmGm3hlf31s695lQkoWWntu6C+5qTOYiTtzWC
BufFNgy0ngC7bqA+G49bYhwJlD48Ctc8gD4zHlb1tr7rsmukwf+9Rnnte/rBYira
zSVMNpbW+zusPnRvTG5YglaCrQFoCgcLqqsHe5wPTOSisaSPqQoadiQxGUipdp3s
QhlpjMgZJOlVpco+W9iG1kBssQhfVlxJu1cgtZt+ArbDrME3p3Te00bcdfG+uPs6
iShEfYKWNviKuChCuq8vzgeNm2VkiCFOiM9bPaV7adP0zTrvbJWZjU/eptx0iI6d
QNC1IRUgRz0AN/ZB36me22+MSF8B5Vtlg0xYW4CbuEjzGujfzIy3YY+Ui8RVkhom
8ZzX6Je2XAUKFf5LqRkroH/+BvPMf6iYHXGUB8VSd5jtmsk+r1sGTg5b8a+S0dHD
3uxOCfiqH7qNjVHIPN9JqWCMpWUT42zXyGZiCTTCuiPnMHa3LCukNavJFQ8jWBmW
NFVRYEbu8zQh4N8T7bx4BxSAm75WI6FbXefSO8Yj0sSakQtnELCBgBbMyxAEKIig
DCeofWmlxXpYorsOcoAdoYuSLt4W+ezBRjFEW5ytMJg0Va2+Rp3QvpV18TJbMiwD
8OFFOd04e+VYwXXTxZWSb6Loi4U6wguyAo6XCI8sI5jjFstmck0KpC85++Bahduy
9CNFhk+UbLF+Ye4Xp/O5blKKRr/365YaVA2yIh28c5Xm/Dk1PjsAekzoBJIlHoLY
AG/U3fHs5N42gYISkHGERK3dUNZlytdSXv7IRXyh1NVuDpcfq2y+oCBEjkj5gI7l
neeQ72pElGJU6EQGb8cESsDEojfU2vj/e7zQKjkPFwUzLw6TcvXtWT3DDEMpiJX0
kDTEkUatZFChAT1jb5N0avhSnkppvdJe1A+MEkkL/OQiR/64FI1MVJg6cH/3qzPL
4yRL+CgeNcQD0rAg3eeEG48V3OBxogoEF8cht70nCUOnUyCrvyaKuAMQ1rpbtTuy
KaLCBqnR6zIat4hDFXVDfhjHR82SiNpwMNCQ/37TZj2rE0/XZ/wxLLdLvnN5P4I7
TgWtZHo5eGQzClKui2lLNAXOSO+3d8NKTrvaE1/r54u5Rh4BgF8+b8tkiYw2MO0w
duuPcgJ62iuxjvGKLdbkBoJs777+KAgZCMb/v+EQ7zhmu8M/kc1bQQ2sVwCGGwxz
Sr5sXXgaKKTxm4/7qFwGH2KnRPqKvleT5cRfX6uvMKbsI/EPFtRWSOwNvWBcFX3V
jSbUeObKVOdcYlUN6oqrVXv0Vdttb9sNJHymm/YQ8j8taO54jCO5Bu8XFb/dP0oT
3dmxM6Ic1qFHhdY1cir38It8NFU16pSbCJLHXRoyihanviOF6olXuw+TX5gNwq1o
VCrJn32KgAP7aTfzEqqGbLADcnuXXfUI2wnzoDe/ekd+aeQ1bHCOcxDKQOh9PF0U
veCPnh0ejlWNzfnlToQTNdx8+4h0XVHGb4GwmmHfUS4cvubIDUFCyiphATRBCLfS
Mk3xAmfRBR3CtTfUzew99he8oRdS5A3v4E7j11S4ZQ7gey7CBieYZ9XfRJ6pZ+bY
N31OYG0E5W2tMsn8/syyMVTYWixipy17pPSFEMoQZztPMCgmTSF17py0FukkdyRH
MW6v+4OMH1iC7d5zYVLeGkgGwM1wjZbYZCTnVO27IQMfVqke1jDGmdP2hKvRaRTA
NLJNZKbWV4jRQ2PnVIvF7+Rc8T0wCPkQYyr4nyc4LjfsyYv8XbcrU1JFOzDv819o
76i7NpOGuKitJ2crccP0r/rWvYbgZGzGV2B1f7r2rs23nWgLuO6SgCJy3PL80mfR
iMyg3fely/SEMMz+GiMC6AdkwrZyP1Xf3hOe9yFj3ywZP4IU3++GOfk981YhbaM3
LsBpthG5IDPoe1DpUO/pFwl8XnYj21ZYc2tGdAEtS3rQdNI2Zxl/ia2g2z9sXnew
TvkbkoDS5oheLk5lRMwB5XT9GC8h69/JfcczR3jxBIQf5SUFscsDPw/n+X1vYa+c
r8qfQsyJja4Iefhdt5naV8UYmNKuGo+9QPu5BIZVc1Z/eKbXyHXifcTCasBToP+q
s8lX9k8NlyLwFWrlbHfJzVPpRt070gVSk6dWkxtIYKXjQGA7DCN640sYs6FZN0PF
qHfOBpN2ZmN7iiHWvmiqaYm7XDs0D/0OXITu1KNfPS2RXEXleujfSJA9RA7mhdHM
I/vfls7RNL5QMIuVyCepq/JW4CtVUjW+CjpTV2Sj/vbX2K4SFzRkxIWRgkAvM5L5
rODB/jNH5nRT9gBhET8fCQKq3GtPXGj+hMV1kxeg2zg1G1ccawXBGm/5IGm2S7I9
EC9i5YwLWNfr7iDZL0akqWPqi++NpT98XTGuHYw1VVgpkvVCEPxOil4napGxM8PO
v7MuLO1PtE1OIUQ+JiI8J+xNlSxNd9udpHtqlg8lvJS1TMwtQxQBS2dzX7IehsTC
KP17X5E5I4ZrBRrq/LJ0Jj1T8g7MVEY8QmAFKmNFfbXie+s4A4Tcy7GmkNxmnToI
MGdJoWAkeV4b0w91h8FCnSY4d4wyoG2waNIERZLUH5YszTS6YnPB2y3Oph3OinlA
20RanQp6ZS5j/PDyJ+p1YhDkGf0XBAD/Q1wP1O1JWm6uALmcLtiOuvCCrW8vsIdr
mdlmV+rE7kKvKxZA8s9aWs8dIT0HcsjqE3fKoqXUz7OkuHUwdtJVGuqVZtOXNalQ
cGbt/x2qOxKxT2395gga+lXzDXi47X3M9ufTyRE6WKiaSpB9VJxEcQMO+gYShHf7
zAtigEAw+EDzdPYQ0UP/57JDjsiPk59Oy1pcIr/0Naks9wgYyRIiKzLJRDHdyA+0
RjC2cYNZ9PDziDNA5QayEaereJnmnbd0HtvWMDnpFY/HTephkP+LJH+6s34I+zPX
Mzg52xZvSDDOqbQoVGXH/HmLx60HKyPZz4BzsxO443qToh2w8kq00XXk5+8bvBg/
GE0CmoKTaguozbjFAyTZIMLUwgFhDiA8rVhZaNzoOo7ZVCj/77t5agSYYO+wn+HC
CDvdgIU+rUDRRdC2NGdCKo9iPlBf0AJnSQzsAE2p2P6noMPSIxcl6I2QRQXuO6Dx
QOR3lx89Rp9JY3wF+W38EGfvCbOBARc+Qlj7NIjO7xvPQ+RphYAwoo54Dpw3iSag
kZo/RUFudDWxM9/pHWUtPHYYTtfphevBiWxtm13ROzYJSpk9BniOboPBy5xwXPJy
xONF/3tz8lCuJnnaz/sEw6l2Lk7tDNYWkzE4ORs/mYlJ/CYp49YzVjTIMN26jgUq
euvHRDDRozJUqeErRlQeGwJIv+2o2MpdyRVsocBSjtwmny80h1IrMaLXZtnhY+5D
48c5X0TGqR2S017qXWQ6KkQS3rul0859/7zMO567Y/SV5EklVkxYaC0edfZojVAD
zS6j8NhovGtMPZ+1GtTNDMCd4HFt2YhzM4iCrpBey8LdKq9LX4gETdhQpkfNtYvX
Wr5zRHcbcd084yLPDTEsXqdotV+fnsx1cpt8IL9ixg8BOpDdfN11XSBxt8HLl8Yw
BiJv3oDxu6+J5OSWglu/9vPY7xDSu2PSvYsoQUdG4bP0Cf/NdQlPydvoLSDuaWBk
/Ngc8DQq1suIO9ynLkLyU/Ffi/D2t7y6PTZAfKGx4FWL7wAq/lmrxNSAi/puxqE/
3KuY8rU1kwpQQ36IEU1d7duBIq1hH1Ooo3yMfu0f8weZrLcUgnivL7U7j2BlXCUf
F53z0a5zoT21dgVHzpO7fOV8xDv2+VQXMs3c9pb+i5xhY/duNdCGAAqhjt+cSHss
rpTOVioHyfcoqXcz3cZcxh/sEE4gcycLMusHaQG5WvwRrmSTF4RZeN8FW25RLqt3
0ZjhY8vVYVBhTE3MXp+LoSHDHHgsDgCMP7NdYtzunfZpVtNbac5ihIstcEVpLeTr
6mWPHDffy5h83A/QoRfKO0n+WoN2gjqRFwvGHhn9FvWDXuREUJszCRMeN0e6Os68
ESYDTkZ7JQRUEfnVnasDWeoauGVeF5MS49BvAt5fGuYzt89optggSYIHk+YuvbPj
/Oe8bNFFmkZE6yzLHxfnTtAg+6Uunlr748Yvlxd0hF4VGkNsqhvG8T7fUcrkdmvy
yz4embCATd2BpTfAURlFQNkOA9suAL1E0IoMAhVsCSOOl5+i1EtTvUbfQilrylTc
Gk+ptLzcmUS2AMrtDL5ZORVs4hgh69HKtfEucwGopzqRQ7M5FOnbobBbgp00yZIE
dZIKOhP7Mkfbyp0F+PmlVYL+Q+Yh9sEqlE88kMGxU3M6HM1JT8V1LbPBQa1729Uj
61Q9hiG1zfy4bEJllIPmfaUBdEXUKNG0xncYhQ95gdtt3/uRHyl4/56npXJw1Sxl
X32RDH9qFhFj56VB2HA9SoTjejiMEdObY9GefVqc/sCVeliTkC7PAovK67Cy5UME
gkKYEpCW3yzRzLBVVNH4YvmsBLppwmKWs0D/zUCF75lxFlCXW30PoIz5WhYtDV74
5RhKFUa5bmZ8Q4fj1vGwDCOI67BZFh8YuK7RslDDOCvUWFhp51OBJwyJqJ5QVees
rTGjL3D0UsNyQ/5jhf51hqaICleIdQQDUD1R0yh0aJV8kU1p1/ajkbz+cBYK7D8Q
a1zWbQ9xkYA6q46TdI62R82/3CfXauuDC+p4lIz6POfJcKbYze9zr1Aewk4oxCTu
GYxC+3PFGqbz1MwMaghmcg/BLiBRoqYNwmPQju/YlvuQmT0Bg1TCw+3zCJ1hImw6
0/AfGngBkJFEgeGM9U7jEYQ85gpgMrbzSbkM+DZB9JqK8CvEk3L/9C0cZJge2UFS
pqd5tdG1mwGUq1pQI/+sd3dClh0XrXGQTn6S/M3RRvJnDDrBmn4+dlFgFfiH65Vy
qVXyuYMKPf3KGgg6sIZcqW/0eNrcbBp72UzpZaJOpjs7XlQwyox2/i5BkXXSWdxM
3pCD1eTu3YPkyFGaVgosZXRbXYek/8Xpu/kWzvvM0G93+wTQiXt1h0tpOnGYX4tz
UGe+ajHGmZKQY4U9RikwgwuGfR8CrKW9gpuxMjza9TwlH+Q1NUsmTzDx49R5EPMP
muOL8LXf+LuulmhIfXAOGkVnGCECfEY9b8bWGYZ+Xqsk8+l2NOXCVYisBRMcac2o
Z3yL3N8HlKm6YaqfjDreEPz/mL9iYdrZ68SAlRkTaZ1rllmAUjV4QdJTJKPf98Yl
1a764g6aWDM5v99Mazy+Gc2yTiEe07tfgQXtQGylvImtWQWixS03AS4m+Tu8RpZY
/oejZABlx8HZ/vGW7Y8dy5/4SQXTnOfoqd0YThS9PBQ3E9ta0XyXB/D9gftFqxro
TVAI8Yv2UJ0s2lnwCBdTK+XdMZ7QrjoH8s7gHoEXMkH1rDaU/mguZ25rwzB8v5RE
qy/Bm9/LsE+NiUjCaEC+PvwFayLn7bk7tU/wbO86MZcZ+8F/dfiZFcHsTGY7Txq2
2aXYfVQFpWY6Xb8ebMMeWf2/44rS+3ke8pIUTIr5HBDP/8mNh7gOJdAsG4kbWo70
Pok5aiBQsqUHsQHSBmvaPhRwt/0tgn+xoSgSgFrMX9aL2zq6X/w9pyDua8CroBlk
Du3EtgbBN5dgrTC/MHvJRBswI2gYWsv8qMLzpirm0KuVCzBFQ4Gil/EjDQ3M8pyG
TQcKjna5HOBOSWSF+nwUKQ0JVWOX0+RxQeyS960+o7c+iO8lB6O4MntkjM0nfSl5
wn3zdrKmp2rP1K6JSGO7qG+F1pE+8lcnHO9nen2MV2ln+AoH51N3zHp9y93yl/WQ
k0ygvkkDP3Fd0Ka9bQJ0fov1QFdpV5lfqo+w/hFqsRRvMtx4Mob3bcsSr5QTJVp/
PSek1PmuuWUuXq5rbPtZUopYvjRUzKgz+N5VDDvTv5ZBXYsoZ/SEgixxabPIsNvL
sdZ5XzqHy6K3Kkjz8cAqPiKQjAu52L00mp70OcoTKEUga8JrBkkUTeraoAIUWEkQ
qxHk+NKdI6KB1pf5e3WG4V0SSKGcF1Q6DPFQGKwP6QNGvcvavegIcigt8zwmv5kE
gVtqJQtzAo+3lzIkkPXxRpzFTYM6PkP1o3w0r/Qxm6J+DF+3RlsLZ82gCd3zR2kg
EFyAp8m8DvLv9EKw6vxWQQP4Tov0QIN2arT+ZlFjIBXHJfwszeDiogXET5OZEEZB
ZpmWyIwXNSaSR3X+GHvQ6kvjt2+It67WxTvxSlqBjky+otYxaKUGcVJQuA92i6A4
c+2nZVsK2n5lEr1fwtnveCe1obYiDIzNfgSAlMcOc57xxJKqJY5Nxgfat8kUj0kf
/aKGmIFGZc0meaDvIP9ZlQQxeLgBaeYfIC1ktw6vuaKaRMQxWGVaENql9rQQWbio
eNyJ8o7Y3jqY+F9tWSpebzvBaqCb5UAoU3/dlmq5eAVyt61CmUmTUsOH1UyrBsYu
tS9It29B/SVP3fedzdEBhzGWEReyOSqpV0mfMU9ljypNfKXLz8iXxXxcXxOguKUr
hAS/FUTbOlC+rep985X33gqEWwmEr3PDGdw4OeyS5SOBJZ+EGnlJrOw34w+Pwib5
Jc6H+5LZcD506O2rLs5in5fhG6J3A5WrzUj+fKJRvnCSSvaw5PeojjCS0TeDvJ59
rfYPp5o8QGNxkbLWgrATblbM5vFPe0WTVFQTGqEJIcPWgKXk+r+erdFWt9n2m0/N
1p7Yc+Unq8BAYBSYeoF7b5LobymSQ7Fuijok0QsEdmzZIfOZQnu8xXwfOZ7ryM/l
JU9csyXOkcHJ33UEJz2axov/NETAOSpKW8HY5RGcywby30hdUy7fkpRKBuOTgoz0
q7lHK+SeuD4XjjHlBderM9N3FUV3WtNExxC/0ExArk4rjzJazgk0+xyf988tAH9D
ffiGdUHjoTe3bZnHaVOqSdynGGZyF6lIKk18yNdLCZqqe11tBFnw78FDcDQnwdnQ
fb/Ntdn0JZx0/4zL/iTSK68Gh3q4JIrHVDWcoWmYkTwuS3rUoRojBNRii85yETHi
Hxq7qwZ82X/CbxHosdW2clQVGNLjhHKXwLgXgzgqUMe2k89kQECEdIeT9NwwOnKv
HXpNMzHSldojwg2EDbAbo8/Po5Pv4yGmp48rCvh+eNxOilbhguiECKpDu9euSCIn
1lt5bYbfYlHvKA3PZRn/Setgy/8Sx2Z6xxX6bxc00MZ5F+co+oFcyjZwV4xLLQeP
TwbRvHz4hTb3HXwy99xZ/rgk/HrFLFdIBLs+rXPD0ODE1McBUX7Ra4WVSsRjLQRQ
6JLN7p+Ew+UTwGqZOjkEf8x6+5G9CTGN86EaoPAA5GPDn6zQi9Vl940OaoFv8shd
7Mv4dzt21fvI/eWqH4FdVf6V2Wb2UgyEk3lyw6GeSVVNC3xY2iTCFTuZUv9dTIuq
sxEprhIgEkklT7oT4GSC3unpHuFYBxMMe+PqyKeXJPdONWdNhE4KMAJMJh82wZth
qgPV2jylwG2M7DusOEtXyexyV/X1vQiDrX36LsLT8HbmFySEY9A2Vy/3vU5nIYfJ
MpKRe62ybhahkVMHFOofGDskLKByCW2ieP50xBSxK6b4vUFBNB62oTmmmxM1wErG
kDJne2Wn7YWFR3sks92nFiPwUokZT9Uu4vVYzZeCAquICVq7aB31GWGPHdJQEeCv
lJU4y5nt4HqZ8p+I5DqzC6RvcK3iucS15xAQ41zFbxpaR4p/Gm1Nc1+US6c3B4yg
V7zbhdCbRS1MSdnhdVP1lGNiKGya7VKPw5iQwRTcNtJOI95FFAIpu40m6HKtaynT
sM2xofoXNikO3tc5KyiZ0cPdZxsjsj/MwnSWtWOOdnHv0fBeChUZslvjv631On/A
UyGGBbwqxnUCx6xcz1rb8+1ZlyBblLWzvrsS/BOVTqt+jfBApFEeDG4xJtvwEenx
0wvNr1TE/XVBROCtL+HchRph9YiS87oGOZ6J836HEElmhrqJPHo+MMkPxBKf2rPH
TtAjXLLYZoFACIt4q5ciOe5dBJsieg87775dtV9iLQznN4qmExFN7qaGkSQJ180Z
ehHQbxcMT7FojSFCkh9qKtig2b5wonkEfQGlFH0bsEtJYWTE4Sgqgp9nbILPemqU
Ns9igd3iwiYgSSvGLTueMFIOlzLHuUhuFEeiu/g8kGJNinQd56iw8BYqHas9zwih
TqpM2kpK8wBf1flZJpGum2rOPnJOX7BaNmGbkneuY+iM3wMpS4CFHVjd/hXeFUbD
VdjoOgESUf01FjxLZYyr2k/kEYy9+8C9fZjnhXKfwTw/xLQt7TZ3Aos+mHf7Niy1
fQMWKsSfWMgl1eFGNs2bPd/YPYV3lJCTVxJ2rexIKWBSRHOKU6SFDHkG+RDHCa1Z
kuByTs9Rd5iYTfcms+s/gCBKTX381i6TC9glgxcMJpTnvLft8AfV2OpRr7eseqMG
VmLtfHbQh7n6dPHPJEpy4bx2BFNO4lb35SjY1J1N9Z1vsKWzeMqeoRd4oScH5TJ5
iSxJVfzAwbkroedyZN8yNlrguyy/Q8/DUV7p7ootJdKx9x/R6WzEeVbDwghaPQj4
r2geu/GCEGoG5pwg4MwoqDpPv5ZlvJWmUZKZ6J5QwLyyFnFapAQ9Sjw5s3Bwp8F+
tcSsXh0ClsdAJhdH4Ky3hxctLWimd0Y9x2C0qJraJvVhhMi9m84Ly7DluXRBsE4y
lycFKgU3ZH4LyFo10FIc9EmQAibOGm8f4wrJuGYjoAcHc6OxLz7HZlhFNnftmSx2
MTMd7SM4h+1uc7kQVcUgP/YSreQbx21aLj3qy0e2w05Szlij/jv5o+ib0YzIizTc
M4xhI+jIlDJzq7F7kk3DtOBS/wJHKHh/RpDSZmxAVMGMO4CvvFAfUOdRwdLo8jFF
gpBAsJeu17uiH4jeJiMc2F25j9LpXSBWA2N18Rjg88oEP7BVSaXwPEnjrgxAtTm4
SQEm6smxmG7HwQ7QFl0ngfyOKVp2PbVe08ogLSOnBgeLF9Ai8ik1V5/r8RLISeyL
3bPFpoiK1b15fPasoHlLx9q9+LTrW27yJxqkxp69b7aZg2B7boNdq9ZjhgJIbP74
XBD997AsuvZ6h6sJZwV6vC3dVELRhURuceZqbXzQbV/qtRNJNQfMzI9OjXzthciH
qQYpyaP3JbeuZ8BVcQTsAXeYNHM6wrl4dgi2+I7DeA+td/kqKMVHJ5HNRyb+hhY+
oIUfTgyTfI+w+6y7HNSAuUhgZ1Q50gOekgDCKmHGxXgzumSjO6b/nbDbhebaKoqZ
QCjmN5puDvxtgnjdZhlhXclzAKR6makPs4H2rW+xG7/+Wy+9vuuP7cEJXmv3CeXz
7JiwC8ykc57kPURM6zNZDSTUQ9m+uoSzuF2zXFNq2S/lrXRqBSUo8dDeB38DrdNC
/FzBlEX+UU6ChDDeqhDZtQ9RFHZr+3IbIKDqXNwXiaAp0bKlmUhlL95+JPwOIutM
1BA0EPuqzeN6HkOX3/KXLjBaEUgDI1Ad4ZDP3hSs1GsRD7W0okcvcM1a5gv3G4zb
gJwUosQu+TJBC+qwxa/zqIC/uTu6as5UEO/ob2XbAfUiNDrikSN+ynJhQwF5JVuI
zCLeNgvk+0nX81ZuSuV4OvML/ND0X4U9+15KGhSeJmgmXnYzvp6tA6iVNeJu9Hgw
39E+fJXuranNWGVUC1cZk0eaK8uKo/H5DLZpH5D/jVzuImIx5OcFn9SiOhR2NTx8
2228M8Adi3+DH7k6OzDdKbCOM6yUPUsTxX0kPbJDhy5LngBUX6aYzWJbyoNu5sz0
1SHGy/H6qAgFA8Zu8Oh1rxeSD+DhZegGCvTOajHw4+HmCO1s6Irh8Cs0W9+vX9MC
WhtktFqpTscPNSrCbUT5yRgNh/hzHfsYMKE+RwuxC73o5DlLmTgs5BRBX6hHX5zx
3Ni3Fmoc8OecfJqvhxvWLdIYy4wNxvYRnY23MSSjsvrVCe+KUAQVsKd1ytc2THX1
W2cYv7cGhIQwh1mwBnu/XRnhUQp5EETn+9WIf/iRvK0UetL9B8MXeFMz/3IxVCxv
usU/9in8HKGFbwlASEXCeSYXcfn7WwHcKxHchVe5SbFgp6Roapt4jTNqKrt++Er5
XF0yyKGdCS2lyl5ZjmPZPRYte1pLwO/wQ0u8nJcE57u3l4+qwwEwieB9zDMvuwbd
nK28Zeysj1z2JtMN4AHwGJex2HQwtG4KTlb3YcO8p8F6qJpkcI4cLWKkWNrbUFFI
PssZQMozbPH5ekOStl9hx+fYsq4mexTbILbuZmqtvicgnwPf2BKHdjnC1l2kLO8T
3ZVK1qsHPWFEPhy+VLTXHEzAQ3w/IkeqY5DkmSvtc6Qf2Wha1N4+h8wT4AClP56R
FsVm8pTJzbbrb8JRXk0Kjrkfkt3NZ3BqMiRdEcZxj/eWiOYeEpUREzelA+KFNLqU
N71J9IbUCnZbp9gR7P2omls5TXAPOKWR6EUfZbXveJqqXQUpXcb9hNrgfzlCAmD8
lJLHjphfzVEuNvMXkqyTwFq6+v3nfAFGAkqPVGlTSj/rU7ILNFL0EYP1LfS8MgFk
/m9oBCIhj8Kh6t85OPWyrngJNzX4bLIDDsNzl92CIHjc1BcgYuLf70JUgUJL8jBf
AdUBD16zQlbZH0gOMqT0A+iVCSD0AXt22qkwEyYBXfoGYPQqbr5bkEZMAYx1kyi2
+CsQDC0Om2JRYK/y08uiNeb8d0QPw8/moJKx2Bq3cwLR7QvAoxmLXbwBkIFgivYq
Qy9USIbT7MYShnbuFQB1u5KqYH+py+ut+OaztrswZj4zgImYlYygBSVeDyFZnZ8e
vB80VW/eATnM18M23o4qAhvl4FD5JPAR6BtC/SD7a/bOgKePKoKJBnFzU3VeErb1
B8rgQ3wSVg2GNrR5lciIErt5ESBT/IQfpwJI+mQPvu+pP3UbM1oMUBW1QeBK4WBQ
6MQOM1qSyk80OVzZrrtYhm51ctmi9qPNN5aGN58ptcFyBp15YSPGb4Uabf+1Wrx4
Jwf5lqf3Bq8KCpm1xz926AbBtpAztB+hHE+u+yhwmYF9TA1zAzrAuCyXS/qDnHXq
w6P/LrUnAXmxC3wXrNsrTzXSsNVBRDl2coaqRBJJMFi0JdL/4vcEQ0Tww4HZnbeF
yJ6JZnQRQU9GbrupIlb7TZS0wwAKvCkZ4HWwUlznbals2Bwh6yWWGifttZUTBe7g
iZMx/g4F2/S2VQ41oHJlVi0qDBP93iOhQvld5u1TjBpj3gk8P/VyUumua13wn9bZ
ZqPv/xTLHWY38xECvSN2MSiGWYZ/XEADVAsU2DtPhUB9lVJ9h0CzLGs1dsW+4JL/
ueut9vFs7+BTb+x/zWn9uc7xYVtSX1/Xk+dLEGIMnsrV5g7a3R+A3HGVLME/l1Ny
MwQQHo6wcGzWloR2tOpWw8X8e+UD0OwfYBq6eNeuJpjnGjhYs4NQ8Gol+bpphC9r
zBCOdeVZLnxwPeZ2zhIt4GOkaftXNN5lNmBS6xpHd/vsFN2iaIUclxbapcayFaDj
bZqMhP1ptAXH0mTxYi+4rV7CvXibB1lQjlGreti2vp70lP+8ehO74lF/R1friZfv
UiT46ht0L1BEeY9f+IpUYKO5h+QqbYS3Ca/HO/1a2j98gSeIz6B28V6vXJu/LoJQ
xL1ADQR+tCblUt8pOxgtdFFrqKwgCIfHUc5mTJCQONPbpotaHup2bPO0ArxSKdeG
ShExjo6kWxY9Zd73ylAJTGLVnRlYe5MQII5AF1i3vnjIX9SEDNw/+biso99nCx0B
e5GMygVg8UjogMZtY/fVxvazPSrHoIUua5XEgz/VPyL2ZVAdHFjpvpRrdfBEn5T7
kCJXlBhMKRzT/R9TyQiqxd3zK5HN5J4769680nlOwXIrJ0QdlyPKijU/xB2KkHa/
zAJ9yAi/67T1mKoTvn6E2vLPKhZfH3lbPdVdqu/XIMESO6wQp9BlIOc+ubpA72p6
8EVERXMByEfV/+UKjh28vCcSp4zpvxCvwRxgJoHz4asKAR9cyfh2scoAtet2Ez1Q
lG7SRuHFt1ydwJBiMAQUpGbImoDKde7xpWUDPDA5i2/kHponXnY0lCzv/BHCPGgC
HukxY0oMfZjjh6+KMzae8sQRmjKcmpJ4yoJ7m7xHWsm4XmzM68d1oS88509Zg9+e
pB04HNh3ADT2Z54FC2jJ53H7zIroFDakPKjeTCYw3PWWQ9L5pLplYWQ0c/YG1Jwi
sewqsi5sVORP6wE6TezuTDnQjhyfZ/mCsNezkbL5mnoToHJT1xoPAyOxyQRZogAv
KkTUNMBE6HiiMiqDQ5C5Z6yM9OOFVCIdo5Yq+0C/Z7z3+TiRMQXqYiyFzHlS2ZMO
zDpP7Ds2+HY/BsZnF7cZ2ja0XPowsyyj+vlN829Gfy6fZSXT+7YP5Og3za/HIISH
Pmazn4DkdcRqrQfCoHmVAYyxepAgBEC+GTAz2ZOeIEpQ3idw+F/GNuM868Rfhsc0
3OkrEJdC7FY0lYjCvxGB+ZH6rz+sGPH7RzmoFKiLV0kggLpOJmAWowzPTbwWeVe6
a8treL5OS86a+WzXb/4EA3r5/O5VlOrU8CEzL0S/WleJwJxZXeSgmjiP38r5Utkc
QVlLyu2mrWfne1UI74vvk1l2pDpJxWF+6FAYk5cxLWrbmGCeG+yJlLrgDxQfUy5p
dKbqz5K8JsPqPRopCKuCC+OyNCYbG4LBzGdCr67wSzMJV5E2vMT0I8aLHcuuv55O
Pn9GICVKRdapIF9LE/G1hKnS/CjdFSPAtcfuWQ28AiEhPrOi9vhFZ2d/1U18HcO5
rZxiIQb6r3WIdpMLImUKXpfkNpfnWmBLm5zeE3scynfbHdSh4mDFIyzkevAVTAK0
n8jh0bwF3orMmnNGvgwImFGh9jBljJKovbuIJWr89m7qs8/dJmdhZnK/cHkfTSsk
SbdXRdskeR7qQL+srP4v2xILV1V2E2O/ZKW3ncbOG9RuAt09nu+RKJY9yooyHpYT
6u+QuP4AUXw0lq1ZeoOYA3ohlwavTuFv8wk0cuTuT/orZlXDRu4CjL+Z9eNWy8LR
gCET//pk0F7BLeILpae+g7pxHNRMaDGtU0yM9dPrWUhaat6yFsBUD71xjBHL3Tbk
bTErmzhn94Qo9tLlJk/GgLAw88go8UtoQPFgdtMPGuSZRQ33Doz06CHQx+Hk6f8t
5qIdw+qj8FDs5Xm6kj3m2s+wyjDMilI9utPZznC3vP+ViK8W9GJwkkKUq+g7brnG
iLxBLvrUZa0jltRuepiRv6vVRkt3m6iqDOV+kswFCBaW+HmvhrIhucZsq8M4q8nQ
D5dI9NkFgi9E/NNE/WbFoitQmZc+kvbQc5Qq7TNhP4Yu3uZzRE1YXGohOV56ua5F
Xg4zH2tirGgP9G9NZpnKIf6n4KuFgSpfeIeOPB+BdoF7aNtxG5dt88QEYJQ93XJD
ntqw6wly8P4AZSeVsb6hBt/ZXF0C8E0CPutWQWljPf0UpaRYtZ4+J3HUdp5SXITQ
P4JAIhQPE70Xz2Ht9NncOmpNDWL0eMCe/gnHUetTGgDZFRxT5UX0ddOYumt+dus1
DLOW25jzlPhFDeKqV6qpzG1PPMQpOdR/XpD7gUWqKkNlm1yo/QXCAg77wZAcoUgr
oW3AXSFlwWVIru/XZAN9D95UdJKSk4J6I6/3whqmfrh5sQDHNfBSwz9mo0672Ya5
vSN6wRRbyQtq1ysnc6KfSw9+VSnLeM9L5kC1r2akxXN5t2IYz7g8TvB/y7Knl9xz
IGKjG8nXf1C5+fwJJcAm3Z9ldHJsvnlFs/qVXlPSJIUiKWeQzSfl50c5Hnq/o3D8
c72jbY9HrIObD0qeTqDSAeQoe3ihDS2q1n9q92CJIUgWVAHnsIOWvlxcWnRIpaiD
58p8Cu3vtcQi7YyVmC+W5vLmUIDQeyTJb6Z9PWWojxnGXFUi54C62zOpEsX8q/PW
keI8nuDvOWKM9VXfwcq0PdaO8wwc2SNgb0LIfguG4JeIM/X5BKw51L+YoP9ALI/J
cOufdgQnRYQAUsS/UcPGXbDILeZ0nT8sE7my6OWG+GgAPS7EK2wEku/u1lCoOIdZ
EvJ9CtUfVwgW+/mSOXCSgHqzAQY9dms00TXbT0iApC/CCdYw7QGk+PlQhSU9/m1X
3JbTCLtvMBkBUjYyaYQFO2xtAmxCwUu1xucYnxZhxBOMevYH4viB7KZAg8iKMCNz
rt9EV7ni9fkwszXSJ6NQAmjwCaC3mUfexnZRe4c7a1YwRgyE7GEPNexsrdDCLVIs
znQxduGNu9Sbq0hDQoA+mSXed4a9blyGtSCt8Qbjl6vAw2IdEk34omagMA/bi/oB
QYlYtGApPnqqP38SW9GqE9uLEhhkyCWacnaJ6CqUcfrGRmNX9xQTVwrn3ueu76QA
vmf6uUS66bZ4+kWkOyxheq+we6uRX1uOIYmjLbVHZ0M5DI3lZUUcCxzoOMaFUbar
jxfWkXm3zn8BaRRtmbGIHdgRI2JrQ+DYiZdsh274nV4XH0pZhMwvTUekL0/fsL7H
X9LN9j6NkuaUU4K9THq8RSr9q+WkHwGBVqbufFtxdOri8fOfasrAc3blsK/APGcG
LU4Gw7yVt0pZURU/9J5wDSTvOT4mQ4/BjBgfanHZqySEf5jvxKV/qj/y1/RAWCsu
vPtHVGxfEFvUrUuMlvZfqmAxEY4yhluKRCdI2RkndRS0bbOYdWuV7oqbLsmxgd56
92nh6rhEzsJkGdjHADzy3uDQLLelorE2kb1GYLH/wDXRg28C9jEZuXu0MJyDAWco
UDFJjjHr9khXAhK1o55ma5pMntKwh8iNlNuekXBhNfI8NQIpwIFWlHFmAtyKsHOl
TcXIVkoE1RwaVWmpTzKFZKVpaZbpDRpA5yIfNwUaEGk6TPugAHSBSdMYyjDNWwhd
Fu2DsDp+pHw6vAHydW60/pWAPeLaFUzRJxnYXhLcVOUr1Ak6bIDPKYF763FKt01p
yKlM/CwPB20yVgflHNuB4v8Zu1N84vfbjvO+wihvQSX8DbXSrpxRV492vgo6qDNq
ZeuYDT28FIdVtU0e2WKhOEheSH60apR4sZh5vKDB/npEZ/4XIOUcdyHt8tvgUk/V
1ev3F4GY6aMsNLEUfW7fT9EZWSmOkn1ctWq4so4FQgBo2SOyc3TBrNXLvNswFXoV
VgTLKa6Vx84lFNsQlQ2V3GvLMAq+z7/4aaXrQg+P+aJIxMrFMmSTSuZ4gBvgYZQV
L8o7MG7MFOL9e9BBXMOtO2x+8M0iZxO5kd1/0vLsfI6ZZDNuj1Rr8bKWCEWi/ug+
ROePP9h8HZ5xAd7AHwZ8oIxd3pcwDDAdsfDsu0LtrHEBOtxpxbjjkMWDmRX2UK8F
R8BM2dw4umlNbUAKjJJBuEKWHemBck2DfDGBtOlztiIPJIo2gzcO/TZ7DCBBELPh
i12Ffc3VG4kpJNy39mMZuzUkfGzPltnr0JT4oCeHzJ27o57+y/IRqPDy8Gwf8WUC
Ubr63iSUlP+sYSf8IOHYXo8uyqK0Ll6Om5276Yl+5l9oPvoQ0dseLB0YIaQSH/ib
VRcAOkq5PNP3VpdhsNrdZutKTS5SHW6873J7YY3ZxwXfC8WBzfk6rLnfvN54tfro
0LOCERTr5Njmm7gGaI7W9iN1fFC8tsUNEsziqvozGMv+8ggUwcOYcSlEQxYrxWhr
8SkB+hxJWk/Mf20qPs0uFtdf4pSHLim53yNIbjK9ZqL4ycwnCGvjK6LDs+Jab6o9
5b+3vuZNcampTtg6/qXBywNNcdzy/pt4PEunQCFqkm3G/OyY5ufaLaI8LJzYSrVj
c56cuQKIbXpGnnqXNvVpA0RIbKKrR5I9CZ5/q7RElxWAxg3ptQY1yeZq27rJZ5yV
b4vKl5HfEiJYsPlpWDcwTDWOQdZbq7RVH2NzYNw79bO62GUzxoK5Zud9R4A/4mVQ
aH8I1DtfiNph2wfTAM4pnaQwdA+EvGIu0qxTLQTF2RLzFhchvsOMqPf6oemesg/8
rq2xHbHGPWaaMEs+KED/jPDlG4V55F3J/9stj0oct7SCCSEbfZiT8LUAENJYdCZh
rbDUvpcoQhxaQf6PWf1q2hIrSULPbGOvXXGnCk99x4VMauvFhv9rYmshCQU6kS3I
UYThA9vjmEiH+dfm+vJHxmxeg77kp92qfIgfqKelqYy2cfW1pQ5H/T9hRTf/BtRv
eeAsnu1ikaMKpxyZjcosUB4lfSG7NMrvpK8MyarLQiJ3G189a18iQWfj6yFCs47Y
rllT0PrMp5oqRfJsZHLRZx+vVdUCU8qawwpLUoXdjGnGQb5PsEjdBOTvtCzTQ4j/
3mKkax0Us4LBlrFCgRtoZYRC9G8zBuqKOfPVTBPXR+bnXVsvTe/8705Sg2Kc3LIY
1Y6uvVM/00kSCKPR+g5Z5gGwLsG/3WOBtKaFA+RxkjM5YjB5snbXdwL/+8BYgRzq
qzOMnzHBlmYUZAmGhWa9Sm+sD1S4FXXRQQXAXVmLq0SX78LCNNn88uk+s4KOFhKI
EqKK9iD1is13vnYq0p7Ms/zI6ngkmSH5Hrq9PDIflEDGEf44T8suSmUIHASLBhZi
UF7gn/YoHmLGAZVEhd4G9Ddfyp2LY8WdtIEHit+scdiKp1eA+NfrFuwSiiLjx16v
zY56SCyyv9jUHn61eoO0H1E1ZEL7EXwJ1XcACyt8oylZQHwHjFfYEdj9a34zg6AC
8ggk00OgeKg5PnWIEXG9/sjiQT5FwzxDJDEwmAJQtcmfMYAH7vIq6VqIvjtk/Y/Y
V4LZcgj14XIf5V+RO+Y/t5dA9caWmGjZuolb3lxTPOHwCXhWotQQK7m+McgF7nfc
8N3FUn89KICHi0wxbc98oUAhQa+fj/vrsGbV8l2ndHOvEdVxUBwH8ixAB4ihl7Qr
DyLkIYrK3nJIJI520i8chb9Hpn+CSvIphen+3LwLf9RSf5S/zkdDG3Tc52qr1O9s
4D4K3sg3hO8VfSYhDewRsDjD3vmOvuoxgh8i/VoyTNnirLteRTo8fK70tHAHHjNy
Vd7VCaMNZ9sbRYJpt3oVUr1KI03myJU/Dl/l1Vhx+PGxIK05TLJpvSBdOjoPXu2r
wsl+5vRUE8TiospT7723vfGBvMagS7bQ2tPiq5L5gbClkTEp3nULssZDVm/+YF3F
+ApaRpyFiHCsZbTmvBkMn7GKUE5312jTmI7Q1ft11lbF7yBrLKr2fAFKmtkTwoip
XEzx294ZIcf2wZp/Fw+TII+5i/iLEglIA12adIH4I0bu5JI2fvOmKKH15YO3U6l7
7k0RTcgY36b0FeoqIS8BNyrRN6C2qDNN3c9W0nD4i1tXGw4zpXFOArrNzNFR7bkS
RSbGvTBdJSvqSZctaILHhcEeJvSoxsSAGBKiO+pycj52Zl41nSU9BE/CnJChVbLh
Nq6PUjgjpl41pySR3m8ihVhyjU6lfinD2fs5bp6NrYrV7DcvEJRTCBER/thEVnqW
/KeW1rEtaltNG1AXb+K8wXCPHb7WZCCS9WVWsTBT0JbPrH846nxarWwLcKwYWvbc
fIQ/foDJpie7ODqaKa4eqnUmiZfLkfqu3NqseqmDM0n/r/nC0vxYoMn401VuKqnu
VWHF6gWR1fR8zZJFSy+pY3yssz+5F0DjxbaYiZRX6FYvfB4sc3ddUt1Nev6bSZ3y
Z+LbAwbTJlE8LFDR/jFEWDfeyH4Q3bf6vzZlWx3MNsolopsVvz8Z2j4pbZwEb2ux
Yb3QOhTwHVyugN/5y1KqqtkW9ZietHqKF9CK5WHx3J9idqnMtOUPEgS/LSQRBS6Y
AZsPHN+R622R7aqxR0pmlTsv5sFmqqc5XMUwUkzYlVKhIHf2FpXRWacMt/sqWGyl
GiyWy8iNrs/TKUHYJqvPQorRIjqI04Yzup+mkPEBVj7aZ/jjlOoDYQuq6ewwCuZ7
V3syOwtY9nfVjCmHUkZ/qEY2GeCOXQyCGG3o/KfTvKU9+BsTOzMXd3Xus0Wf5mbQ
ow2m9d1Koo+w4O/d7PNgg0I9ym62xijzhaU3WdVFciDcrWFwJxK846+Fh23xFTRm
Z4DqPl6xEiieyV1vAeZzhpLXHdwKsJ51wM9dFw8VcqFZIfKeXx5dpRhnRS/btKvb
hov40L5o8NT7FKRA9uYAgg8O53Lm7K+vH+HdiBcvcxqhUD7I9ICPr/E3NnUUQsbY
XLsMhQtDmKdl76S9rPZHz88IREBcsRcWRVlBSUpwS5KGNh46atgjAP11R5rYHg/k
mv8V9cN3oS2crD0NCIGny6hXpXbTArL/pDnEm8CUGBFqnlFsxYEGwDnty0xoXyjA
HavFT7Em63chVcgwE0KG9o0HAubDhPCM/chD2TLEPc32lniiXDn0pnuowOcie1AL
G4lknYypDlcaX5KrtX8Q22XFDqhdiXNLFM5AhBP0IJ4mh8ubi7i1szKbKNwaEIhd
B/qEVPGLznZ1CLEHLm62zkk0j+H3RtRilSfIUXasfKVtpMgS9mw8ctFl/K3HXEok
fiGSNJLeT+46jxYLvpfdeWjX9A8CR887uO0eqDUvGvPPANTpcqhWLWmXRKw2/ktH
lRFE8L8NTp1ouE1yAkx72o4TebZMe+r7SpyzmvspamS5oLEtcP/aGiBN3jTMtnim
RYb4c1WGmngjShZuGZACklome7Hs12d0xGLp0WvcBgCM96ohNWJZ444Dc3+ja+JY
sh7VfngZd5beIDqRqvTos7GbfULuRwkL64vJSo+cuiyKk3U0xVDhpHYD+YRfDBcH
oGh5Uz5dkPd7OfeaV//tpcEoENFLJ6AIcW0pWz0Rom4XHtR/hyGhFkKFb0KGe2Ve
frbuwGUHmXoRgvNHFZ0iysTHRtlbTxdeVkLLXUhES3qCkRpJ9lFm5ekSrCpDIrQV
tlZJiH5mNBsQ/zR+VLNtvM+R2JOiDM9O4DisZcKXilVhm2hFj9pYEXz4XGIBUxXg
o0uG4lSAuKhTWFev632uAoeCPPZauVLZqxGH+/CG+KY1vKsh5vTxq+7A4koS7AP+
G4yUDHzYjO3n+VI920n1lM2oJ2IWG4KmnGYxDx1aKTZUOPgGu/QHDQQbssZyLwdy
f9iYxfFGsdDWx9mT7EvRll6ht+EtyKwCn6tYkzxODlTs/+QNFZW5u9X421tDV18R
PKDj+Xcl6njUCgEA4cyqXOW+WSsG6xmeV74c6kT+IBRkfaD3pZLhEe+Xpe0DZH1q
YsTzSweGqAOOkV50/IRf7bPus701powmXtxVdLZLisWqlhaLTvlkBRz47y/g22Gl
4xdVVvTyqe2SYuFEDODkBNFCPfLEJVTEc93cNk2Ff7a8Nk4fadaTrhJTJfmjF0n7
DN5RVlu1Gz5dd7mjuFK0p2RsPndSivJlDbb8kPFOX1nJD3ugEt9lpoUo3jJHXLgP
nCjx1AHP5Jr8GyIc+zTUiVO5awGBEIu57Y9XGdKOdp5VKILZbXyk6XFvRb8ADTCY
cEFW373Wwx46J3nV66Rw9R0VRRHjpsbTkm6ASNxB8+PnHRjAqOxKZNRzBJZMQRd1
vQ3DGD2TJC8M1eBmnxJNIDsqKR3OK4nGKMfNzwf0N52FG8nzNEbErBAhqSCww/HY
Q2JrOtnEctTFPVhB5W7U6SAh43Dfsd6ISNhE2/453BDxBBb9hGiSzAUu99HMvSvy
1YWPXnfNROe5Jv7bbGptGa9oTCGdvRHjdJIADLBDPvc8hiX7fjqgDe2uR8D4HLA6
FsN6pbY+jffNchzSP4+oH1JIev2HJEmYpb7wajaW4VKnW6yIFHwN0zWsqiQ7gaAH
nJkNaQXgpniaK+VqaFZsaJQUc9swrrHslHITLds49E5pWw2fBFRTMbNhtIqgU4C+
mEtKrFLcWTL66JAs6R2hfwWT084XJIzF8F9YLVze3ZS9/+EJx3+sj7T8HZxC5van
fjzBVDZNEz9eY0P6Iat8KJ2jJ6+PJCIASEtgM0tYPBTzjVmZZ+zt4tzba3Q7E8Kn
YywbUIIG3ZQH3cTNAIuxy7LqBioTu+5fMIvDSFO2j1gr6gXxD2hbYpe74Vk4c3om
NKNlWB7NBEwJMtMa1kc+SwWdZtEHIn1KzWpHYuZL6nIJ0PvsM829OgReo4SmCtri
Sj6wZYqsPWHBoTRMAImPEQxg+SDl/rw1Een71wWlUvd6upx4edXu5+3WJyeoGJtr
KBDtrjTm6yku8Z9DidFmIWcGcwcT8ZKJxp70io5y8lUThjIxsDgHBF3Pp/JsLHpv
uW2uHICJ9dxyR+lpHu+n0zyALPd/nrFU5ok35+5vlMd7TZ9Rxo+dd2bsTDh8lES0
n2cVnYQVKwDiQbfn5eziSjNbsH5fVC61KwicV4u23IcCepVFhk6/01jB5fl2u/Kz
lZNqCkhBVZ4uthVL097gdxBJRoSarb+s1KXz+vFN8/kT0axXfiZSyaD+/5BuCeai
2jThv9//YfiQJya6tK20mlQUxKi3ghwVZSMbBIu6NPvEiyHKOeKeXNVk6gkP30xo
8yA6t0b3ncqTvjfUzce2iIZZ1Zgg8Gtljhiy7UIlx2lUmeMl3Qp8EVz48kvCmfIR
koAFYCcefXqVST3nd8vDN9jvJESODiQf05MZtB718YKeqSSiUM/UDD7swUYAaEJj
hUSZv6FgViOD8+w0ybrPcj1tSebGWbGjnZ8RwbmimCDWfe0ntgT7PNYMAxv2iCuR
BU0mraHiyWekKf7VeTdprzgTphLj54tq6I01LcMFkNNkaQaLNbjmyayP7GempZc1
kEw5sTRPf89Dc6C37GFZfaVrJ+UpusgMMd5PGKYLY3gRf7keD6Y36MDn+Cb3ZllS
Vy9LcfVU6iZXYkYSvBXX2f7gbvIY7xWxqvXaj3cbjShC4rIEOnOvY13mtKYRT4xX
gjBMFAYujm+3esonaaQu8Jhnz2jSTt2sRpXP8fd5ggdQJl4m58xe7RSAUI50bZdc
6Gyk9UZqEF7ufP47PhKU5U7+M3cVcQJ/G0GTvBFuvwjUc/aGcEZta3zcYEu4GAU+
xXh5dl+Z98Z8b9oe4dJeiJh2j/D+zid7fvIXukA3z2RugkhuAPW1cuIbNTw3oNI2
rK5Qgham5/BrxjKk0OSNhy23WRjRGyerEcSFx/k+DYpt5YhqnQGBSxpTG8fy8j44
yKSD17Dw43yxhjIEMtirkz/TgXKhkrjn+kt3vRxmsJJqbwseRl+qBAu3tEcDuW/l
K4LKKfwGSPmMsrhp22PPfujXSTeLmn3PjLfpGBkDk9/q4VJDRlma46pryPX6MAgI
teDoRPEoOEZG2MQhq5voMA3I4fHH+KOxVK3AZ6ya9Z8XVsW7zmGvpQgW6RHhuhaD
0XK0ElzIeRPeHi1F0Lt1yNc17nrpwbEn1to85qn4SDWS7nJieM72KKmshRSjs9N6
OO0AFbKB6zSMjomFBYQ08qGM2pkyDEKwo7lm2hffchm/1Vddm2oa7nY/k6x2UcT2
rLFNwvJsaQ+Vr3F98Zy9utMKXxB2RRXdCBzv1EloQ/nmyvzEsO4kY0dM9FDTqIjc
sD1OIa7hxp8rHom+US/MgzmLbYFOn2pXiP8XKTvtv9vJgZCPznlt31XJZftKq8CM
7fULNR3QUVdB1FAgrw7mYTQ791tKBKevRq4Mku3nS8jUxtRj+SUFnd9vW9wHIvDu
UKfj13f3vwIWpRo7FcB/voGS85V1gQj4Yrgu30bvzRGMzxwRWkLjMqBzYnJZ1z8m
9tPyt+JhvbUCcluNj/QM37xvMkuhYv92SNtpmRupWHRyESzJKOsZ/RbQxRic6qu9
TmR+vSOreoMm4elzJriDgmISJHbiJvaGfgNyHbT4vYwQbkQJX7pEiH9PcITm2neG
hNv/3uuiMgtUqqYj/3gOjB7F38fPFWhCA2XZ0IwQjTmF61zENO8A7i74ZXPDQSCV
+a8je0H8DFdRJbXvkkoBCIhEek1538kCNRSLNl8wtX6MRLXOXac5GSiT6lotgKf0
jnEfx8RiG+JB1SgAirUHQb781dXZkfYS+4bsGKCN0P0LL6k7SUQrCPJAgtXcCFs4
MH7N2VUDaopJeVjpN3JU5vnBIPsZrYHGX1khAb/lZTQoSZOdhTe7j8BglNH914ex
ENY4pNFCVYx4npEo9grcYkhC8abMeRQ37FTL4K15uFiVJ2hUerEPDSnPv4eoZqNw
zW7HlCclKTRUOWXOc7m0+HQb+JtA1X23zCo0oz2EQvdWMPIpTBTxeFgMnXgMafTc
GPkmnnUYxMCNTxSzlDmX25cmY7kjfvyzoc0xG8/kuI2z5YhZ9hrJFD/BDAVTL1Wj
Va3kepSzRz/0cKe/jnFZ68F/w1QhKtN04/8u82OmKdr/iWZN3IEqeLgKpnAehlci
txjCelzXvre8xTySXSIUULlIB8HJd7l07dWDptaLlr6vVqD7AURys/Sq1dYQRlbN
PX1BjUU0UGelrHZv2napxgemK0fyazYSB9HoPBcD4gCNuy270IgvNDViq+vcUsMs
MXKSrM6oJVu2z/+LT66qlnmWNqx+s1/k5VdwtG4RyL6/YcydwclAbpidE4QIcjjO
DgYrZaomPFIscRLz1nnVWEeDUoo7fYsPJ2adH6dFYSs224msu0Nyu9bJW9X2FbJ2
qShzlBUa+V3I+poU3bGxnvoyW5XRrw/QBGXWX7Tjquk3kqsZ/pfDNDDyI2FkVAzj
uL9N3v5T+5BtwbY58cm2+NgAG7eJKE9Hy9w3ij1ZQIognd2O8Nl6Ti8EBg7w3RJK
1oXiU0DpLuad/8Nu8kdbdGQJDXemtgjyFpPw/YUNbGsIPSXJVlz4yVGRsUhOY6iA
Zl9gdrlzIf3sLxRJH+dWB6c5qhIWbtTAE8zNkXRtek2JbLWU1BC3Pp/cpHVBUzm7
Az0AZnQjqpXyavu4cLA89x6Itp9ck4NJCZVnsjyGElm439jsQoAb3Gpo8h482TkY
JfxX6rTskIzv8gk1SIl1T/osnD8mNkTHA/K4AoxMrjnUO9rQv90dG1N/EZvyqW0A
1A9ZLD52tmB9YnI1NGMu+/uGwcajohEyphQBAANJ+dGi5yOXeWsdoqtQXrOSFUWi
WgCcs4ziQnlk4oWNVNR0qGZFOpQXt3oJoukWXVxdcmtfIC2TrtEzoejrHxmHfv9l
x93gwGRMmK+xiRMUVtv/ZhtQr4yy6RYSvZ1Z3LvFWV/i1leeLRfp59LULR4WU6f6
EXofj5uBUZYW+cFsy3WqoRoRl+lTxLv96qGr5hDaVJzoO+jEpJBGrNB/dTVKjJU7
dQWVTjEwiLdTnTvqpmRyrn8aBnV/v6cYtGFvWs7l+/VeWQ/TpyQziH0kyAfn5Mla
Om3JX06JKiWWTVOIoYD1EvCKzqDXy3ZIPJDaRpThm73To2c67ANnfkX/VcKND8se
exGrXhC1He0WbID5JkWQvlJZFieeRRr+qWgYDgzL0YzfN782pmpbNsHTJLNnpSMv
hqXgAV5g4zpNr7d1/KuRmNiLvtIQZO4zJOlokWqAOy1grLECO8COagI3veminbMO
HgSbT4VuGwrAmzUdShaiJX8ANgtC7IcCdmbYeRbi/b8N/IUcSBXJR916xzhORaBc
leRltGzfFAt9C6EDQmq+EnnOqCwCBWRzziED0oRYwpFIWlMJii9Tcbql89sxduO1
zjgxglBY5xl5XDKTeup/aLmhl5HyqqrYviGYLMhvraOMgCoipZz2MyumNKRVT+bg
2fvGGRJy906mbyBjRX2Yt3FTNfWvuD3YqgpkBX9wN9lS+wI50ZAFNU/KjM8N32/s
25MmNHv+iIVu05BT4//pawNd6Ozi1JtCMuR7Mg5PiqSjGluCj1gXGawohCDgKayt
XQifWaQ2BxwpNCQE2JCwtoEZ03Z8b+r3hrWXdc8hd5/UKBXObnERbOpn3o/mL1Bd
qAZL63Gq1aQ/d9ksuILSpjyj89E1TvAqUajYvL3QPyvjaJUMkKKbhXE4N2pg3Lfq
dXQ7LBZEeJrvlMkmTLYQtOiFO8TQnfATEfhu0EXOaWAAZTzZTXlDQyV2pmvAguGu
qw3E37vu+SXhouGUOwdE0tRBkaRFEA8La5oQh8F0efKsFFwj+BU6uPUtDnYRzVid
hOVWMvcag5qvSq7jtHWDwGM1Oxq8NsYC6q8u+lKKa3P7+BVMQKPJDxPK+B2G42lx
UMzlm93isLp7vdIj7CqvVABnMtOc4TLkZpZgRUOkBqi44DxPZX/88egjd1S/QKFG
FEdo8qgqMkoBntGoEYiGWChVbJjp/c1jzdTmuGj86Ee2OPlS+/NtbYUBhjAd0REs
dUXJUhpmE8GvhZtSWHhygplcz64JX4uIgPYsFCqzJb6WAfZm7PQyY5IRsR1tkbJf
dWyU4MlG6bfhJYZVZ9MXRWLE5TRVGkI3bro1Qdqp+IRxaIIVske2iejOaOXSraPE
AUtPQQ/UXCAsB2aa2XZUtG9pwho3k1t3o7z5PbQC23BNxR9Ry9fE+wjucRQl4BAi
aqUx+Az5aVqoUH6XJbbkj17sXIGBPvshnUgstOJgsDQ3QYaaewoAcfjiohXk7yns
yG4EQfWVzdd9GwhcJ8pGVPi1Py3vj3yX+rmupCIWMZQ4GGD2L4vz5NcIy1csKKx/
cMzCtVabosjMloUrwI1meGrCZPQafOm2FYsv8yJKg9yigGR5uvb8vrUmT2Usa1vu
3NV5FtZdAGFoc3GG2jfEKD9NItZlvhjrCc2JOjbJwYjmLW+aKjoFNXerEkeEbRQi
vt6ka/YKeacCuowlNukKXFVJHGUPAGicMBy/SDosfTo0d+x2jai2oLc/TfiNiaj+
+7cNazJBEEi7apG88DFHf5dU6OXmb6+RK0iHL/2hhSHXWHwNR0MAoYGV8jcBVbGN
1x3YGpzwlpSK+CoKj38k8wy8JggQ515oGmR95dG5pP1rcC8mgwSeYn0Tsm9yo5SC
rxBSXcQgur1MI9fCnu2cgttCQEUBQw2Ju2g3Fdren0ToAkLnCK0kr77RGtdBa90D
PX7BXTcWbIw4FRphRAr8Ab+5bI1NuhcPT21rsl2FaUnl+FYAdUZOVHQLdcyxMqUY
Qk8oZK0zhDX/XmlEGQfRQ5hWUgVPM/88FDS820Wkzw7waZ6aWwfqQ9SMDsXxsSPP
2Iq0YpPQez+VkCBYHwiS16XjYKe82NQYwr64WcbPkVR+xo1q5RD6iDXrhtn9RYUO
r0UuVnXLugjWgmXFsT84f0dYJ0TKI9w4z+7icBZK0nzbz+06+dO2g1GmDe4siTpU
E5IIh3czXfC+sUs6HUGrwPY83x1BGXYWUgWXMxhd2ZzmzLqJa/kyif2tlpqYSoEl
pX9VG3MRq61/pdHxWpdsTxB2nOnuCRo1SrQi9VQrcdZFWnbu+Un8II0awbwwL+/d
/FCHTOk2Dy74rzVSzeYzOeMZFSkA9oJ5JJJDX9mMGH7Lr3GO2dZuF/Cgdk92N0OL
jO3HBcVjHsfoHf7hGjSNvEdK6nIMlzInBCoxgIKwftjP8TU9ryb+HQEMIDXlDSxU
51lCW+uXpgjXMb3a5oXgwq1cd1ROLaDJRVw6BitqULvGXv4POuzfxZNNzm5l9hC9
ZuYywpW2bwJBepQrZww2CswNuj8j2KIBEsMLfBR4saEv+zIk/jq32Df5xVH3XsR0
qjyxQOMLDVeAJCZZ+121uuNOnDJZiPjWRC9cEzKDSYC/HCJV4JXp/DkzpZYuxyMP
B0T/fz13Tym5Z8ZUl0PCdb3a2Mg+yg0gRgpYiYWQESR6A6qsm0RhpwclVWezvNHv
qqoGLVmAl8eurQjOL5FVi+ts5fWc1Bd/2JaNmA0X2WDdvDcU/3Aj/dvCSLihUYqK
E6vdal4dkboQptZwZCUOczueJQMzbj9DzJWmL44uzHBoUNd0rSzjJE/YnNU7dvNg
oI7LYtMdx3hfpZgY/dgog5B0162MaEygR27JGAU7+/qX6SFwFsBRRCo0mgL6pWZu
5Gqt94ibJXTLU09zN7m8ywct43mSNkf8fCT8NNXua7biYp+hBS8f9w6gpz9AXZH2
HiAcmvp0TZqY64ghF619r/Ck/E0cIpkIxSmKhMDhyyUd4iB7hSScx1u3r9QILNdW
crILiik2JyEXCxiLLfcUMhax4TuOLWSzut/pak5X67330q9cv1OhORbu9OlSh/Bs
Z8LT9KLj1tPaUhmFAhiGIVURTq4BDNtc+LkIQIRvqNUW/s/CpR7G3s+8fv1yikSj
VKy+Ma0k9i27xf2LKvajaEBd5f9f48zkmACoP+qqwk+p7TlWLAOWuusS+L8YDMuo
HRGLzLC3lMqUHsQ6yWaBrIvFRM4iNdvHLVvJE+BfFyk7UG9k4t/k7mcOe6TIAKCi
xbY6laB8sNZHUYPaExJZKpolhi1z26NVthBTOQf8c8Dynw0pE7gDmW4ebLNwWcuV
+gnErHIEEh7yVu/10Tpl8Aj2bve++kJ+FyT3218Fg6ijt5vYXQFrK5L9oqKfP9ze
PAW2Qm+jT432h1tjjILrisQBFi6oHCpq69FSujMW7gwY6zmRRGMlrUNJSoEZCQhQ
fb5SsG6muuLXFm7UFyJwbFy2mdUJoDuS4yqUDr97lhhtwQ03lQJS1CWFUiMJEfqz
rGdxy6H0swQQsBhywPvKo+lX8qUXNG0HhRal4e6RqSzciXW6sWffiFFUUg08Takn
laoyig3FrtalFfbAE9ZgveRmTwLacKCG8HUJX2nHzTMufvX3Cu3IvP7Y7OXCRXrK
iHkYt8n2elpHpdeiGAlSPxSrMjwK4kBLI+J1gx36cBDLe3rxDiSBjCt6KsXx16By
fEBN/BOy7yQw/J/GotUCMVYiPAT1F0aRTG5o1jy5w0OEkcnSskpbQPA1oTO79odx
O4ic/27ZwacSJ58MPe2l8g/QIL/H8dJ/UkTVlN/hSkSLlBX2wKpHJSo6pruCZbRV
mOU4UUxt4O6mRmrSTxh22KqiwcDueE8FXBY5hGBIUr2pKgaJAInj2TchAdIR6nFX
obXCZtAMSgItSitzOufC85pllfpq433cNJFjZ/Y1tCWR9TnXhq2Xek8REU6mzgf7
r1iwno1ovJ0Mm5/niCPn6B2Mr6M2DVLa+7AUbRG/yL27cB37Qt8Ffwa48v7Sw8fz
uL1E3w8L6vdfx6mG5YZ8lBR+hLzpbDE4UxcvBfV+ME2kOz5atp3IR8wbQb5wLWqh
Y3eVzxqAc8fI3u67aaS82s9fORwYNw6j/m2Ab8RDPV2cfUxYU8k7Nvt/dsBDMPnn
qJoZMK6lYKeidE5sLh5Le3kVDpPDVKJ3aoMFCR/RhB5s66FSodfMq9i/kk7CGUwI
kbjzWAA4v5jPwLFw/kkdrRw/W8uVBcSJD1wYrSsd08TX8DESNTouEHjwcrdowA6b
UIFUIDxKx+5kwke3kTlN52c3d6dqDDPJTtjPGjd59JocnsMQQiN1OTJRvrMavq2D
QZbVsAZTjBhMibvMP3ZTsauv7GiuubHuOOZ9TTeWf5knP3XPs0EeTE8+osKQEPv2
UgP+0pLChCN/mN5TNNZhgnILj3xPSdljOk9tENuk/WpYehqkUkk0itY8keSozbOB
w1HPqsz4MUgYmiwe//+B37AC8O0oXvq9y2pyvAlDSiCgBOwKWdymiz6Jlc2JCpgw
kPUk1U/sKG2agFrDv2IWP5PKf1X09c3Z81E8QvRU+xb4rQYF60NneHowEA5q/2K7
rbkWZ1nQpioJa1Dk4Mv+JaFkm3n1LdetANy6qTN44TJw0RUzP8SPKebEIpl+GMpP
x/UQsXz/m75KFFdRR3oq1Oc14706hFYIC7PxOV/DnWoYzKOXK/UK8bFWIxBNvxCH
qFqH1/4fIpAOc0dPGBfhAfZKPLGPZmsndqaAHwgqhdFLKF/+ypAWEQPG41zMtpaw
IJ6qqt1geBgl41aEh4EuKmWXkb7HVxvH4COTg+ReU6A712zDa+mYvsoa3xmyFrmV
0rguV4i514uer8TdaBK+zzpJRhEBgG6dhcUDY7k/AYhKT+eVTxmekiYPkkvXmMao
+P3QY0rvqJ/9h97gQAc/eV3EFJfCb/02JALu4OoyL/hJdefsmbHsQXMSlpOrYV0N
+BA7CvbWD9GVFAvZ2QtFmkvTsrDhIdoEAexuA31UVnBBroCgDZWKN+h+u234EUqI
8MRa3CP/WS6AcMr7Vhkv+0keNvU0fRQtp+84/bJJozbKmqOhB2oR7qc4j7Lk7PRQ
grTBgZyDlfiusi/izAbFG0Rkp6Z1TUTfHiqY+DaqwpC4lNBKUkor+ySLHJpOsuEz
K/mjQ8l+R+Dhp3C3Nz59NKt0SFstBVR7WwSt9byGIlsWWRA67lTVFtPAJPJE2IVK
Mw6aIsASFOL2h1LhVI+EftxBYNLYYY97oY/XtNa2+yWJN+QV86rIlO9esxviZV6O
BFE/6+YlNAx0D+Nqnp4EIR4PtPpoMVqSTJ/GoHUo6UVV+uyg8ru2BFe8Mx5WITcG
1+oZKsgEjivm3EGzfhWg4rzUS0UTyKqGJuSLIeDfA5S1G42kW2crX5yQg6kccec7
XBo5qBGEUVQ9o8oOUR9OFACAzrT5GrPxR1y/ycAhPw+J+X1OiLPxYBxO43qO4LtM
pXrbAi9SfAUL1Rc0f4pbH0BuS54LFaGeXPF03UPgIAjdfsFRxn7gRsshnvwiJUa0
iWMDUTRC4frx/DXyK+/5L486Vtxtb0GOaVbXfkoTbiCRI9/L72XO9Y/tul3V1ri/
Z0MKHbrNa669fJu8npOXAXOrNNiCs234paRFJetMtuPJj3MhU34iA2yaZJWRt7pe
9/cSonFZSSm01GUKhyTOm3LLlRshSiyFlhM7zfb04PMzwgm9cP3CL5ZJpf59Aza0
pXvN9f7G0M5sWEEDHiTw/EUvCl/hNyoMpUzVBms/AuXOzsCUPQkp5X0S6KPlwxPE
+SG+DkcX+F12I2I80bHbgwTQVKvr1kEs4GDQImvCkfWbcae/FITEt4wcUoInKd8F
zrL0V13Nzk8UARAE0qkTDyXv0JgOsNh2EQpafruN0x+B3G5Xewnd1BAZ/2FvSwLe
ZKMd1cH6FBbvmzpFkq0BkdRVHLoA0iEMK70UGIKP1k8Ff/TJhK29N/p/MniBhQmJ
G6Rk8NfZmqgNlsItSK8Yjbt05E9PFgZSEy8tCJ5HstziqYcpFesqseyUv/OJTM9Y
hSCgXGSuZOw7Mo+GFsfq5yqkKr1xy658MILhB2nOFq+2ngTK2XuXv7Zes/+7FzWt
4hxdwDj6X+9OxyHxe7SOs1HyLwWKWkZmHDcJ+YVfpSMhnq9yZiu5bgsQgwhybt3A
McrufgjoigxRFe29cA0EAKhzacFbNAaZRsICedZGHYVe80mWzInCGFZ003mfZkEP
ZNZWgQk4zwi7RVPg81Za9lYdvT3GJzrO9i4vtre4nRaudcNlbKCNMdLDZp1HXLt7
aZwwyRthVhdk+BfeMZpj+ie1YhBCUujMqwN+p0XqV0QLIEAeHt0cUzKMg+WP+LhV
zGflwOSVnc0NAcFOTfamSBzCn2iMrZjPA907ylhi2t2mNPGp3OQYmUt4K6pOGKQA
7ydK8yLinmovCDJFcZgflljzoa6kw8K3szSzSeg2H3LBJWD0FZZ5V2EMf6CvAMMA
YU1lJ+inykD2UBHXb5QAO1zQvf48MWdkv5AWLFC+AEKiTjWTY5aX+s7qk2zLDHrb
diB4ym2dYK+2BpK3mK8/TmnOg1myZhrPd7d6JoS9tS0frshOwH1LYYyn8a78Tz84
ORgZ38Is/zsLdRDsAlqWQmpWtbPdC0tIaDbt8uImZxzWIJFcByMVlzfXLY2hb/7P
CY5ENd6SdsOsCjsgF+qWrQeA/sO1qgt7UUoxGKeagveihAQ3l0776bjWVLVXptnQ
3q90vG+/kOB2wDbADr4hgRcfeH+NgyTOHNHLoYhpFJwAgRAwCQXzsM5fOVjzDwnR
iM1ZUBnXSAi0pzasSFW22YFFFCnc8n8V+fN5ZaI0u+Fg3RxJOKh7DzFKeYqcS0r8
LtbEyXUuw9mw/fPz/AXV0XKh72wuwU3+FRYAxBi9mFnwg4AN5WzXvFxJP7Y+RpCS
u1j4teWl7tnsUHCABYAaAuBiOnpWUCEQs5rb2A5+Vrc/Y9tdeJ/4UAJ3UekVcukB
6yxQvPr2T9PuyTAh4QHdAx0IIOT3GWanQ9VWMbX4oHm9tTSMtFFAxFShosqZQwb/
HbzxNmbMcFxQwJpYPRAObh/4/z44bu+NuEVv7YmmH00Jjd86n3Ad7iHCpFBBVzMn
1biOsbSrZleY1MzAlTHN/8DQX9DoegFGT4ePG1UAI96tZnPHQuPghY3Jd+3c0GUu
Dsj+obDciyU/F7GprTAfP1vO9kIAM2r/Fpfq5ZYg5ey2J8odVoCjNOvOK/MgA5T+
4rb6KZLvGQiMQpEEUsdKmFGMe9u2pqGDdG8nBFSPojCfTTx0mACVh6jTkV6a86ob
yYf7JxfxnM+/pTUHIozYd/mTE/dWZ3+BOztKEgdD752aE2ffe2XW3ImP2oRsul9s
8rXOwRwkLAnjGkkanygRl6KZ/A5oYzXlfoEKIDslH5YCtQvGkkG7kQIHjOaY9DRT
ef+jjzO/q70sCqiXRJZ3DtfQ+30yiMIyFO4/BRmCcrYIR9Uf4yEXqmyQewAwCRIE
w3EGTaUPJbTe9Zn+Me5B5KV0onmYfEXzX1bk9tRINZOyjkf7tS+aRBR3s2mpSlLD
5UQYfCJf2UfixkPnKMzf8qQX/P60dQ9A1nrV6RK45LbPKgrRX66QsZZtwVQHX6u/
XKIu75Eo9Rg0uIHMTaEuwz5+dhUtaXbYWkgPfuDiM4mx/kcuzsVLiyRX1ai4HgSf
wSPfU3DDYh/06Atw0zzz0Wu/V7Gd/D3nfyvXCWM+VJ3qxEo3Vop+TY8ITGDefShB
6b7YsBjlXV+Jln5Ht6LrKrwaz4dhRH9JGsCMVsjAtAV14WaFU4oE/gGNKLbJiyxh
cFT+HPFxRvgjmpcdjSqmu4DB/ghkyVWJbpXefF+a1LGfT5GfPleUVihzXvXrU3aj
Q9xOKv/dZxzBUb3KNo2dFtF/2rqqUC/LIzBHzmtV0dHihwO/8UBcH0xRI90b0v5p
aTSVY0xa1h7emeFtA0kEQSfG02d29Nb0M+Q7k71iQJIReJ2/zOPuZ/U0Geh/2upO
2AxjsGUlroGUnFDNMcgz9ChkGXwTJ8ziLBBlIE0hxetiyVsPGtoVssGbgv0r/Vr6
7HSvRrI7hVbmE2ZAuIQOSEPM6yQXteOEBRtdifzb2xEvPdCzJdDh7xTjBeQCTHV9
UWHLr4J9tw+SjfF+wdhNRRoA71Dc+B8QLJBesqzOXKgyPm/VE6PwJdamanjX5tdc
8zfaEiukEaOg5GSAYxSsiZg7nfmuUbWl0taIcWiMzIPh67crxwK72wriFM/0Z0X7
HpO3Nov6IahFZsT8+iD0L6J+08YFapq0nQSa7MShPDwfhEJjbWyaC09BvqfhUnbi
P0RhVP113mYX1oW0johsmWc+cKAfI4SFColq7NIG/Y54GNjuNtNn32y03xabmpJG
/jiiEVFPcEBR4/jnXvaW0lNxMkDpIx/As2d0e2T9kywRmXC3f0sThnb8HU7Ipk0k
7nzAKfOI1/cVPiPnNhF5Y3kfwdyth+/TTAid4HcvYgLH0NLWnyZOx4qTnoBNO4KK
9l6gCR7xdxdDiU7vk9RYkcjldrCPnzSyOz3yJcftqp9yc3otbIwdW5U8z8gdUQw+
oCNx/FIZWNzjGapvLNz594A0/9ZkpG2ESI/MF8GcIBM/lvjPQtPWo7MXLcG0boLR
coTEt9smQ9y6rOBddODbJm3CR7I+pVmEH1WZmw9f2u5dlSFxDBFFTGO0TpDYig+T
9wejCmuY0SxIHeGkbD4+IFs+fyDuLIyToY5DIYjJ5hs8zi2vvu3pEbAXSXNeLccn
lNDBenDFN3BZmE0pCJ5+e9QIRp54iXT8Ah0fAdc/DcRMzC2HuxNmDd+gKXiKP3+O
/7YwUt+SFwzp+8b+4f9F42My2NZXeIIFHPKIkmn+LbKoteuYDP2rZPoqD9UAgltX
Cp7RtrCX5ojFkunVEap4+TH67XVgO8/lHvxZCs2sj/QoW/1sF5cK/m84MwSK/3E2
PJECn5RAPHvLRdZ8PDmrxWX6i0CaELTcCREcm2bf0T0c1reoZv204W5tHa3o9uU2
MVwfIz5z1/7/3mam+L6fWK1zKue0b5HIk31Gyuw0y02MSsIG6bbjY84qMmlyxMMc
4pvphFL1FOd1BYbFjHApUGAfCTYIeWuXYp4agdoqZqZBy3FyNNHEHUrGPXgUg7az
JAMONkIx571Tuv25CLhM1QfK4qZUKAksHdTF6sOJ/eL1sLMbEYxHiuC/LOn1OJUk
qmDaj2a6vG49do/x2DwGSJB6nJvi9925MnnLx/b0U9VUSeduhTjz6iCcCb/tcA15
qXn2cx0GEPDp63uwPzxYrcEXsnnw88WTtjJ/HL8BDuA5h21nj8TE8sz5Xv4nVp7V
0dwm8RWCPRrwcmq1+h4RZBoHhsKFOPX+EherHqSBOciPBye5U6fC48kBEIPHJheW
D79Re+drNktWESHYB9fRJ2wQr2UhWYRyp1HpkiJFpmIbRHwohegeX+7QBXMfgwn0
TQhLn65lvJyf6TUKWMaEEt39S/1fyAF6gyrUHIklsEAVfCfdP0pQGjbIkdShZXvA
O/Qgzw1HutmG2h5n77WyPohyMtIurFBmklwesFn/TEeN+yxhYT80ZRq3NKzth9qX
ktIrS9lWFwYG5s1lEdZzoQpGEnLi1jSJLC12g03iPbMt3sC6Uqo+zIdifY1QdaaU
eAEwvyiW2ESEqkrsCOvS9M2n/qCqMk19Sp6LI4KwnV5a18CtfqqDsxKt1SiqGwn1
/ZmWhJquLTt4i/OBKtNkwvnRIoapYCsvSQN2TrxHDnXyp0gNdEMlyQC50qvlXqpx
V8aW1lzWu9ZjuO7KWeQzdxxP0pMyt6ZvxKwDA5hUflpU/QhA0mjYG8iSe64lfFRC
kwx0AkWtiNxUoqWOeLyeHNyia/JhekyAW2Z10AyxoTKTqP6nRp9wflbNIfSZdg9T
+35eZKMwYLM5rlv42sptJsnMaOjkdeSvTsDz56W+cxFrgBMq8ejGUyl9lcOm7tUx
L4CPwQPvV/NMDYbLus+GA5+xxnHdt8gulesqe08PCzYQ4YAlRXa1mgAhDI9efJHs
GN94BXYZ8bEDAu/s8CSmm/sNj0Ga3KoNbbd6JKGC5g6zOyOjzM2gzj4GW9qf3wwW
v2VPzIZ+EFil+fJOBIbq8mr6uHIshi5bJYs7DZ7n2fkrYpHFOFSHVuVBn4fAP48v
PtpovJXcqvDqZMdojvaP8c0MlLDOsZd23uS3ejnd604FDWkWXJC1xyCPMsQja6Us
rUaF3ojQV7KIzLoplXC9XrZC5uTG+YaevlYN5Mzv3dmPt/fTyHErjWss47Xt2LDg
aYUH+Pr2EZe+Z+iUmOTHmIPUYaQpZ4ko1/uD63o+1fSfMMvdySeXAERJfXd8gqGl
jYDGkEhjvAc45pkGgeBkJ5L8yNcQAVOb/bVBmxPSnsl5nSSu+BRBGH7e5ns1HjLA
kru4RgC6fhhFQC2u/gN8CSkVZpVH6gdc2qVzKuPYH4dsRS4by2CZ412Rhrw+57Q+
ly9aEhoAp3uvDys1acBj8caaCP4QBp62OrDn5v8LLzWP9znQjv/4D5vUk/CTbHxS
bnEOE+a4IFmaYyw65djb02RKGUqVnoZAmQouxLzuyHL7sNNo/JZXiC/UX5M/hZqe
Z4/sS+Rcbx9YBESm4PnNfM0aEVBccVeCJ/HQtCk5Kmg+0YLjzFEnQO7NXIns3Txr
iOppoeFb59PU1XHMBD79oYI8PKfyOTd6c8jLHNoOmp71oe+GKJkn5Z0fPcqWBy9h
b736EszJE+/JN2BsCvCaUwIFWx+6+OmNJQaMhcWAFMfV7IwI6xCdkqpOwG6j/47t
sisf7ly5D5To2Rv2YxeoXhb+D1x8Om7RZbmaSEP9tzCaKJCxwklk+xHptr1Xy4fm
cOjVAPsXVFLzPNFgoWnxeIAwdbo7e64Jo6XSVHvoSNibSfDqm3366MO+7B9iCZ/X
t7YqWShH0JXxs7onShWOR2QzJyVqZ/Hq2k0cNyR5YVmT3jigXjPqn3blSKNQ7y2U
Ng+jxQ3QXxB8d+RKNXH2Pjra74a2z98KTgkv2dxsAvOnGFEhDEnr9nzbF3JOZPvl
Chrjd4DPhFC6HA49pOdZiyA3qxF7KF6hMI7RgkTw+q2pisGuabD30BjcOxfQ6p8M
o2J5GkLKqmdR3XtaWDnWX6MprqlrwGUw0K8ZdvdrqIMvkk7epSyi8FHy4vjwrEa0
tOFYsXHUtRXBDUS2FuI/50qUKX239MvIWkA1YWO/nMIK16Rdh1fWDjkLMfsAQPPu
+pzVdabzqqHe22wPh/+TwcltnofBRbuclwxGlbYC338oTcHXaEjj5oBOBxVfQII7
6mS32qtl2I6Pm2vasfPjk9H5TMctzFBIkZAtYP1mZ7+6VBGfLik4MjUp8qGWxg3l
y+VzA/YkFRVk3QF8aGqox2aAaJVrdjsBQua+o/5ayVY4Xw61z97lvId8N6k+Foyj
3t7fg0YJFNF0n9wQMiRU/S/sOYg6pf5+4MLj6Ly0hVe6VuwPP6uuNm5fXOWfbXDe
0Yu+oehEBADAJ8rN45/FNmxCHAo83XUWLp/8rFVfOj8VGQ/Ul4NwXJ3KohqnlK0d
uZbG5a6wsid6QZgOhR3ZZB+Xrg3ELON9yqwzSoXzOFL2bCQeCgLxOyov6K/MUE35
hpQL4EZfnsD4HOhpRS6sa3cmJ4beTlqLy70Hj7iBdH4/v74HTQ/GnDN5xmutOrlE
Uo687wUFaVDwuP9FxmJ8cRNDpuzGEevbdGTVvPHvQ7Hwttf3cee/y/xmzLS1zZBE
yfqAw+17qVrtak3KHcXLjNgnKBEOAAMXCri4nhRrl7+OSk3AOatgbbfC+TxLasnd
ukAHd66yj9sewB9ZsEZMEnvkOD0ziawzmbj01mBvRBNOX8KDKdamLpWQ0FXypv6h
DzB6cWLzpifc5wnpJksR+eNWL2IpJCk3Zh4Gef5v0JC0kZRbOop1SqFvDpYGUZuE
GOD6GHeBBOMcqP8M7glBIbzN1LiQJ1JqTaMr1ZJkFVhIleR1cf8SkriW8tPJ3jYz
nrpYe4wbPsCP7uOcnPCd/lQrAzf6Atkwbho44kbgvPTGAtyUzuonre4vqrq9O+fR
HUDdEABek+CcYrnHnUrMU2pwKXSaml0I2qOTjXJpftUHds64BRCYxVjoNRQUn3KC
lAZgxUA3xH5THFPTiv27p9vEDmntnJGf+wmWevkD/9flnNlE60HHrFFSCBSK/5NC
NRsRf0+mGNLF/T9E/O2fIlboF/N+5K8ZIv7+z4/wX/S7j5OFj+VCzl3uNbqlTcJv
8a+GolGAFWzKWstBuMz4KPL6a1bkgRe+3m4GZifkVzfy0S0r15nbJ/hZ8xuN2wqU
AZORnxnMqcobRdyUqmgheB/oTxaPQNcYVvnGCiRg0Of69ndxCwk0U74+ypAwPknW
gb2+WrN23lm0CNt7uTxpeSkYuzHyDlF+LPiBcihatWMJKaakYzODd8+Iw5S022EW
3aNiypUmTLtNDfVWCAZ+U0AJ5vhPsNE9kQymGzKuSh8zmNlIWgnmmUP1mQtI6B6n
cRJNQGu+jLNbizDrc/yBMp/vTy/sU6jYQ59s6m36aU5uF3vbyUDB0g4MYieQeele
iY1m5BSkuIig28+96PL1qjTrGzJZXWFVpBgWPhvRRLXBnkR2sNOGrFxLnery27QP
o/4XeIqSeif827MnIPuqPSyJJ00wYhbPFDHx24re3iZu9/9r9y7Xrm4iALge9puS
VGdp3sWZY82fCc8As+vhb52+H4kdEJl7GM2wXD0lSPoiASCxPdAy1I3/lAQYjekF
zSp4T2cKAzF6LcyBccoMM707cJUF+wCep7wpMBVblSYNw/RF4VHmr60SyuJzGjr2
IoeteXn07Wt8vb73qPpMpmvjHiwBqEpGGCs1oH7A+P8sbpZYO/jL8XxyNxgFs8qX
nHzYSC2HseMffWe1jt1GccDzGBFGzccTvDoapdde8ju9kaHRbzkL0cfGxcNIo0Yt
HBOx6cqRCOGrJ+K6vjUPEbaXMvp/ZnCXCv0wEXFMyy3/WMsAYQ9QFTog2xTQl0GG
CHMf50nRDB2psAIfxvRYVlrWIYs9lrPJybrR02r0fN6ogPwNpgXABKngRt82sNMw
srg8jDbVXJX3/NqQygCz+quV7hfKkokHh/L8uGCynJLRkkrJ5sFZlDkYmLV1Fxs0
SMXlYNOGJt/jtKN03mn8emr6WZtSc9N9iI44nqJLIZ4pYnVyAaofWIxVdzQDuW+8
O8JNR/pVAu3xDbgD69LrYSwqOEMQvvnOwt/JmH61VzCjq0SlaEgcLRrqH66K31JG
5SpRhRBw1FZOlOrvPwPfJXsTWkxTeBkNLIYZNrgNnHyqNbwmqkTuwqUnQ9/AL/P9
sasnitgOr98VvuCfqEyEXOWmZClQa8hXq1ZMv2BrshVQMroI+gPFVceBwV1aqaxl
fVEfNy3iSs9A/18je493TI4ZNGg1eFmz49VEdy/zI3IqYUSN4UWdNCXgyfIjHOFz
isZ9eUR21sBUpnTb+/xmu5y6MWyISkKB2s4QwNKoxyl1+Riqhc3vU2uEf8JozvUB
ebsxkAhJnniGZExtnDfZXQSd5ci92Egz0iiRUbIBzS1AozJfEAM5xqVpSvkYm8Fz
omXluGXAonYtGZuITGaOGOgZpTNLDe49DUDoWTPKbFO9PwCgipOl9l4U7fkHZF6h
Lzytv+MRkgnMNydUDv/N+3mzk/r8Q6wuoiPe4hMguKf7T3GyFNNk+xP3rncWngat
tjOYltp0R4QVoB7pzB4QFndRbp8Y8aOnYeS80nL7C431ElJxkDIM7qR/QOdwGsDV
BVEukn9zPd0S7lGuKAg1hv7TQFyKNEifO6c33JhF3eoOmEvC1MI9fJ5KEuvOtKFQ
N3P8a2xoJerVGHRUustUb5BfMRt/GG5f0/vG7uPEPSa9YepfUSc14Dp6eDaHAfhl
4rTNHnjV2VHByK75gNPEXJu2LCAnSYJkw+khquaFA0++x/VZ2fAey0+LOkruVgQk
gY7UrwTVObXxTBaQLzkpFeZKzp0UUl/fLclkvBpKF/oiJ8HBAhkBeXI6SnAFtpPS
zO+xRne+h7m9Fwr0MUKrsXd52AYgFH5TgmFmLm1eQCiW1UAYcBHF0QYjYWUu33a3
bY4FKc8K+IeoDOIkFcg3E/I0JTwVF9ivHz2Uv0HvF6IcN2Py/LegoScVPeAmk7r0
ZdeEWKKbAVbwwo6lXHcsrQ+KIX7VRGzRUwwWPhEa0CLT6hg3AJJBHAZ/XLnD7nZJ
O8H7HwHgj9bSEJa+DnNLmvijc8K41gqhi+OjoP6dDQ/Y4KilQXS3kFh19/HSkCtV
6+hhQEQZuWXpqnOrJAjMeNz767ENWAtVsEMVVsQSA83f7DCiyo4mm7OCMFhWcRcB
UQCj86IfjL2kg/9FvkWHuvdDtMu4y59FL7KM8DMOZvJg8Ur1iuJ/9xMUYE6B4oWn
AnVPFRh2f96ndaBkBgad136jfBHqvT4ofDhHC23PIClU1J+tFMcuWf60WopdQ6go
9neOLRf9lG3Els+XF0mjoeKaMNB/IkSWgYcNSdDApz6yBMNQ+Zqt7ULwrbeMStBI
bsm50tz82KlQgv9rTPCiAD5m5IH0DLXziRXkAn3KDAtwDO1Zdsrji01GDMltILkE
/ByOmTui7tD8TqoS9+H+Vs4RSdnxSeyjs7aTNypEdH8IVJHZNO7t5ngYYZVmwdoS
y7lzXtRqiSdKq2FDemNCHdLlyow9/BumLmg4S1NTPu/fzxl5MYtBHGfTWk/SuD0A
RBITjFIulC6LTjfW4wvjv8yLJUJq4BYXwfYYnRWrpG+CQi9Sw3+jGIJqGoAiYMRU
jo1M/zAd0TcyT2xiecC7UlfVOvo8EIzTbCLkdzxekG05uqqfS95+Ga2EVmshsKZI
ZGc7D3aKlUhUgRYZ+mZNGD0O6N7uZOBMu6zcWq34lVBNVuTOUoWpnnb0nhJ8O86F
B3fUKjfQxZlS/OcBphO4jO1OT/Tc3G6G5C9VuTE0edw/cgm1jAJUbs5/KApauWIO
C1VRcM4KPEfq0bXXYrwg05oCxVkX85qLMfqUDgpbPzTaNz+Dhx5FNyaQACgYytQg
gQK8WKIcGva3LeSlUrZ6Z0o5DVQY8btZy08BdR0a3ur2B6QU/9oEGmBFMVVXMCbJ
isRaLcuUKzekh4JSwIiz9okMu8jUMacAscde73+5JhWlDmbN9cCQFlGNuZ29NLg5
NU0600PDBkWiwQXvq3zIbxCuOCLIVwx+vY5zEl9qImXa2VBgni+iUY/FQ1Y6H7JP
J+kuRFv5IJORGvcKdOlbRUhOb2SlYv49oVRK02dEBbOLUDBWIal6YbTGaQW7BbxN
miSPFhWcRz6SoDN3cUKAsySVU78o3DDpF/q8gQMMMLWI5MZiZVXac8WIQ+JB3x1f
hcVsReZ/KdGXMI+AF5DNoCu4mS+gDNdIZM2iw9ggKAkUAFXn+GMvpaxOL1JLds5Z
LxcUP5MRz94WNTGul3o5YLbTmNwLDaOW3+frLg8VGvoHKlHXATQaQK9145hCMF9O
Sy53losseMpxQNIlL06UFYHdASTjQNGnOrLrYeDojYCiMb9zjmZZJ3glVxdyY2ya
284dFZ6hWogyb99ldUU9nr1E0E37Q3Dvjv9XNqdf6a6XAfxA+4mCD8QoXYbybNqG
Lrlp8ReI6gpuP/OL4xzbfkZHaQQExgR3U9/KcEQCyr5vgQ8yyOXUivc0RDEJJDZf
CqChFb38qRZ4HF3cnZI/wJdOnyC4s6SYdHjuQ8woi29ootlCKTvSyGz12BnBvbDR
34tyTbJpvACHv0edhESVZjev2oQWl7lLDpFoGolQ1qN0GivOQxhX/9e7V9DeIwic
2Vx6zUI0EG3KtXeoS9XRnf0a0wRNMbPSwRHSyGiWguzW2AsvrTjbpnGSytJnPEeQ
utMCxsj6zr2qzpDow0tR9Z9Uy/WVgKTUIGJXBqNlZmHFl88XDeLi4ON/RkWJxZL+
RS56v7IGduDlq5F70LNsh5jnlugJZZwqZYaqnAUid9q47mMcUW8cl3IV/OkyBN1Y
oPoF1pf58P7kBUwy+ZstAxbm5VqGfhZicRecQYx+FMSzMRakgVjtZcl2B7BtzMVp
jDXcZ5sWf6HVMNVqAJt3slzQwDjWckYkyFBvH0H4PmiibbhISrLUb82wLbf6MQwK
/LMGDYkm6o9TWr9vYR/bYjVCOafCukbbtYApgNt63jiJW4MwD3Xg53v6tgaYtkuh
2ITem06iflA1ywqGWu7IySmvpOqFDlin6AXTHyGxZ4RSiJY6aKQ9FosK66JA3jgy
CaJscYsUV+Gfpo181mDtPLtMiqLsb+orctb2eHHZXnYgV40L/D8YQATiiizRLSs1
kLMDCOvXhF4u8nnt/hucYPWoCV/tyfD1vE8kpLO8o6aeMqeucBJVImWyepi+1DIn
uJHzFR5MUa3PVS9zh2Wc/LZutT96n8sQyq1MxFaf6aRqXm9y5jNvFu5hh+6IpMLC
O6+F0d/ULIBdNcxx8Z6rP9pr9RGe1VRVQ9pxpt3SYvSTUE0/0CmPEIVm0lR8oRfJ
8Ts9kKrgR0c3bFfclMGDI2VkaDaWwgvPqR4J4NCTWGRQe35MdrKGCx5KrFNf/Rl+
LAVZ+3DYSb72t09kZdhkno4m2kydh78EJ18AdYSH3x4qjLCbBlpTkeuDvAufo3rR
DKdS2hU4of4w3ehnRE+FyjyFvKjz0hn1zUueWsZyLYyLK0BJPYSZmPjcBu+4x3Cd
mcZ/rqgjyiAUkVkwPnn9LuBOiEJ7FHwYU4ALWP5f3HVGfoQE1CP822xGsRb9b2VB
WWPF66/H5JcnUfjCiRpucawKGPPDei18AwxO2To1ESRKNIod8DVn1tSUEGuXbh0O
+sjdrxQqy1D0nVorD07rdaTgJsO+9q5NE1NP+ane+YeTxcJbNDu2/v3U274msU5s
FrJxlb/ql6qDqFbetAfsJsinG0JaqsNN0EoaG3/LGn4Yf/k/fp1p3bMCrHxiKmbg
IsHwswsfpn6IuMbFIMbi2PE5eQw5gJDGuQaT58Qvs7hPPxkObzQWm9OoukDTN0AL
n8Tdw7xPEzV7f3pNobPa1YH+FdTBhDST+mgWOREJq8HrTmoe2FQNL/P1IVdnlXh+
xGRO+JRWuHU2bhx3949NMQHUvLRgzFh57eFOgOOlOPcoted1YoV7eOuwgeKcF7ch
uJ4SOzpHDTZIau09sMmghnQlJPAKMX1BuPMjPx3OLeNyvjmLig/24VEWj0cU7Jfm
AdEqAs1BrlqACimYMvfGEAnO85bdWkSbh78kjlMJZWviL5GAxHUDpuse27IeKKbE
PBY1Dau6SyT3rPTBReB+YwM9ePfoZ/sYvxeItjwQHP2u2qYShrabM+rhVZ3+HrKx
3WVRS309rRD8WPhg8ZcNVdaI51Hl11XU96dKBsBLhq1LT6q+rKqIKy/goRLAI+N3
GY3D/bNJiTHOy8NAoG58qrYYKN33bJo3Q8xmudrwsizFOKTniMLCE+sWRn1OjF7+
O2dk80Dw2/hLjddluZkwRYsOBi5/uAKPkwBRQ3KjjmoV1Af5CpbT5ofXnePkddH1
BeSrF8yftn6AZ01d4CRKL05KkSNk9rRdG7ApdH291n8huzQWP0i+MjfgfKhmGvM+
2SczT9PqzMaTRZKBJCCaVsKIzMhRWqiQIpgRSpq7B3hdjZpXzEySxyZC3iWTU5Zl
lUt0032kih8k/lDri56izCx0pIaM8OQnux5RldoiF7w0a1Sp53wLfGJNywrAlt0w
NT12r9zCOnfnmovhRrx0OYR19ibhZfeYrk9Jbf3BtRFvYJcPafDVGtzKNqQpkg/l
iu6qVs2iND43yogI8VSo8jZJDlEQicsCBFpLTijjWbTjZflPG+vrq1OPeYIXc66y
/1apDjazCmJiiCx5ckHHh7K4n6t9nUMjWiUL4Hh0rV3eG0c//B5w6jw+1TXZ3Aqx
bjMzReaCBSPBhl62S79XCJZ4MvmwrPo27YPUPDd07tDHL3FCBgky/BobSj6B9E9k
MSz1920QbtMsg2urPQtv2dAj0+fcmRcSUsR52QGIJeJnzWEy7pEtgmMNKuZ2Yd/C
w8lxfaNl+iqs0ofrP+mvTPQfDgn4xKwOR7qHIaaVXJEI1EgPscOCUmcBDmAuCcdw
Jdq5te/vcvG0F7pJyg+8eRhwZ47lEcpHBns3u6lOaB0vryw3GkvdKwD+7RR6NtBU
zOEtWY6t5lrPyU0mlks+mYfXNHWnS6fUrgWlnVXfpdJJz4LAAcOkztP+3ljYQ1iy
KpmciFVKUTQcyOphnMppfBzWcrG1mBZtkqD72XDmfE9hLkrprjFQYXrpl1ACAe52
9dgiFYC4SKb+XLUxyeIqhZ0hTmjJ2yRMBBKs/ELill5gaXlQ1r2C96VnWMST4R5v
LMjt3/pFNVLuN4E9spxMHc+EYY+s4jsnQdK9OcmM62QYWAc9OKi/A8nq2U+7DkVp
k65w/WvuHmkeQsGnbSeJyBepH6tXVAgJNezaKnVzoF9p65Hrf4CSUcjxqgDHSM/1
YzQMAafAKwiotpRA5FnxeIdMYd2TIvYjTWfvtkVYt08yVTGZuvLGkonlOW1YlafG
VMVAfOeefjCVNzoPLHlOld6zBhguKSLrpMzqYz1Ia1XQ1UujR2TQVrsG1aDoDmM0
aEx9WKNS16iqSf0ZCnllpnoCacuX4taJV36BQUbXrb41YCCapPhECwHuZ4pYP5iZ
VpcCZ66rXYcblbBfmc98LPwpSdjcP1u2j8/HNE9c5zbUKFmMMVv1ZURl06h/Hio0
hnZRoywLvbvk/0n1g0TSzkgIY22krY7IMk7Vc9eyayttChrbV5LLrcM4lpZmu6Hc
p4VknYQgsC0ROEFGbTkMN1se8Xw5iFas93EUUnEIGh7YrZw23jJdnJmVmdMj30KQ
hTjRJrbw8qgIDEW110TvmjGmr69XhBez0UWR8cyJgpv5tWnLl3BcEMcBCe79KXY8
8Hc7TMr2PAXx/breMi2ISiO6/4U+DDh5Gc6TlnQk8K/vnUhkIJIeq7DD4vCLOJ6C
fuTju+tdbuBdt7Yv1d/6Gq1mBXjwJvuRYpALut3pYfeEn8QLRQvuEBU/iAeuxyMP
5VBTcrbTXuGWtOl6F3peRq1AZMz/38WHiAdf3rLeO4SVauTq/qBr/tMe7CieNriy
DpZpUWOUpZsqJa/jlUPwTAfhWEEQq8GnrejIrNr+CvvE/0A92yVVJ4XS8pQduym+
rEsSYgiQl0eGtgrgI27+LJqSQnmiuTHaBMHzvo1ivNPbSeKgbumZEsatlyH6zG7g
K65GPqWqFePapGFH8CpRYt7nk1RQJZP9ckawrDx/4ffTcigym4p0D65yBDxNGXjb
xNN4i9hiYAt9tcA4Q328/SG37usjHe4PMFOzaW7/AANj4s3XLUqcvWgzzzw5srLK
pyFXJ0M1sGZFFv2nUmeBU8hsAae9+98AqF23K6nD6xD02dgDSAv7MRWTaV+oCfHd
Ohq5glg5IvbP4vG04HdoPkwSe+KgHO7AWxOQrh3smHswd3vMjokrPZ8oN7rkKgNO
HcJKl0+i3LkRQYT+uCcthsYJPhGgUDG7+q0oGXM34H9BY7lv5iCSf+SpkMNKLXY7
7NjX4qpLvr6ph67MVShW1AGKwyFJQh/oAzMhDsttA3nt3Ul7fNc6sCw9jjkjKQjh
EMz7EzPOc2IwP1OnJBASRRdQuEuLFL5u9wDZqAL9u80MY38x5QbFKwBSokRLxE22
WDU6I9N2lNHrGQA537rm1OocNIL67ueAc05SD8dSOKItRzc9y8C/YBy/g4S8d0aw
z34DsYXeO0o3u581pY8UZg86LebF4Q4M1aln7kp+CybwkixNiv/nA1KwxKGjRNJB
QdjMR/1rRjzRZTNcYbRTP+T4N7/pTaaeS+uSs18+Tc898H2HvBUsoPfm1NdyCv+/
PPfwzI+LuoAN/uSCy8xXyufGGlevp+kIOQjNuaTZJHzEmeAaLPBV2f3rq/T+JZ9j
oopU+KDqvcUsSdfOUd/PfzpMHMnbWxAU10Ul40VetVGgDeWMCyABaX/Z6ehnG8K3
H0GQdhcJI9oVQM7OrVc8BA5ZwtdNAJnuGVa26JAitwQKX55T+s6mp93HsAMEGjQu
ubrwg3uVNfypXNgT2tZhYagn2u4/sFCoWr20TORkXJbh0Mhqg8k37DHLynjL1tV2
Edy+oVMjeXopXo8y+MMcsMC1LAoH7NESNey915pioJQjQzF9L9ygSjeJbjDyKQlj
pkWq1XgaKhOaES3ieSw5G8QcI0nMQct3/r9Jf/aCc01a8r/T0q7calMpGnXmB834
YaeWz7wOn/wCMCbPqEeXjHMumlvcO/KhkcK7ZD/zLtoilB1v1NdovT85gKhQpoXi
bLeO+Sc/Z5PoTA30A7+huw94z/v9kRWnqzNk3W+rYw1IA2ijdLm34MCP1SQmoRn+
hsOo6FILbhCU/GgtiXI2aiQ6RLwlQtgm2w0h7DKB3x+hWYvBkstSWfV1RS1Z+4kY
WYQ/emonNusms0bb4uqT80IA22uwvbH/Algb0PujkqOF9GEuNusVv8jyO+lyMefP
vgSvzLXLg2jVEgPi6j0EWxHhdV8G6vHOXtEqRh0gDojkJPEqlKcdWML3dTc8aaPs
WH1Js1iMd27dBWiDYi34f/8sRtzclLWuS7hzdd+b7UgAaO2DMf/PYGKu+rmjcuVD
xc2OXFt6DJaW9AbVaLC2DM/qNN3zjUY83kBSC7MCIRvph63QqWZRKfQXywyz5wD8
I1DUhLJjjY03guo3tWry9YaWObxdkHAABz6jblnnNUY6bIOCa5y9JDWPRrtp7rTj
iieyM+SNWVvqS+19ZvGej3sjLPCaV8XoWpalt7OnHCz6xrQEUcTnUXIa+AeYTX19
UZ9PxMJVziH1LHqG3Fs6c1antT4TFS+GzKTc8QhN6uxB5Ag3byHH5LlgIKHOus4A
9txc0QHDzKGaJZWmGvKgBQPwBZ0rIvSt4s6N+rVXLImQ5WIbknIxPTOna4tPiUDg
WBJ+IrxbmY+UU6/jFlbpXwTgtSuu15Z+e2I4C+a/0/dU7wOVKf9iJRqKT8CZ6S/2
gTRcQpKGu28/AsYx6EelQr2N7HOEN7U2y3hFnqfljBVDwfhPZwkwYic+lL2lVkRD
EJXoJ31WXBXTX3DmTSRCr+93nUuJ2yclKk7ttaaVFVHgokO4liIZ4L49uUTtHxZ4
R1KT0X9T9HeYOmumLDJqFr6+cm3NeZ9mcvVcFRt/28dLhUUUsdRA66JPnqiP6HSc
52vD+c/GwnGZTMa42A8hHbmk9LL6pAaiJUCMy8YiX9hq9gw0ZVD1QeZcVtA1uujN
U1b1LGtwQ8dIZ8z0Euvkuz1g0XYgjnUoUdw7P1tU71V10r126vMJRxXA7KpZ5C6L
dsI+JKp0yQaZcxthoZQ9a230J1Px4plsSwkFzRfx6xRajBQXZCoFsFV6Q7BgqLhK
RKeCRmtc9UxTPPuwns7u0jrllCLZ2dbBd8QZMhjm3i/tuCtwki/e2mXjBP7bWlMl
d5ZMtAcHliN6VzKPJ87CUEZ2F/mnm3gQX4TRTTk79o4fPpnHAceGFQ8HITv9gDKx
u4B5R08vlY+IgTljPlZMQIN8mDExEDWacdFlj/zz/Jzfu+Ht5SC/WxPqGuin8TC4
UoacYHreVacVAbIpCg6zs4FlIiGxKE2cTNnww0nkSutniy+cGpRiMes+x0ZyaoZn
/cfMK8XB5EiNyG58vN4rVUQDsuyEFCDpatXyGw3NbolY7AxCNVlWogqLk/MNlnV3
uMWJBtcTUaYOGBZCyFdZzWdd6wRVZi7b8NgDl6HJUlJdu4hm8weeDohKuaPBCbNS
5VMzCG8Q1SnKqlY5rpau1hJ9wHxrP5q/9OIur0UViZFWMNaik0qjQB16S2kNPVvP
SA0IvwmdbTH7UNYWh8LW1NJLy5enC2za4rbZicSyEWFmx7BCtnhgh4WrYDLXpMqy
US8oOy4gIZbZDP2wImT5cMdESLK46fSqXdkisvjY01ttlmVjsgnplZ6bB0iJrpma
hpsUkR6/e/Jx35/zzjixD2IZYA/637RXCvlDhTRmer0cViskQ8UbTFM9vbea3K9e
x9s/J3x1XTWKz87a2Hm8Qcjm30ZQSyTBt7hhsD1vVckNuAWL44A4eHpNwB46rEsI
n2myWj3fjqfOcThR+NOkqBGe5CHgnfTnYpubePy6wEmlM4ywm2drdLD+Lj+2f7o2
GHOvtiGZC5lSIEzTM4n80JvzllVTeXIZLKsNHEJDJXw39CJfl53xZe/BYHpBxr19
XaHAIL3pjZLnmeifOWYLesGov0ButZF3GQoE2HPWd/WZAM31phNzK2gkoJKMkFtY
PvTffeuyEratZxT/Vd/WrUxRCfBxTiqQsbL4G873T7iznOP2zQqTRueOpUbGbGOl
d7ezDlkDicEpgu6HHH4je6FyzF4vlYGBbN4PX4sbACOAUS5havnxHO+ReJzfn+iT
LveFwNTkqM2Aq7X1CNn4gOdhMdOsgXZeuWneJ9nT0apHb7b2ceV7emtVWVLlSh5w
weyt67x36p3+lGlyEedG7An79a0QP+6L3LC/jpvmuQPoQCQFUCX6HRaO78/iWTYP
RC6pPrgZ5H/d+vQ0gnKzE0Emf/uAszGNuQpsyXhfXAnd1k+W+ZQKMOWG919wQcYM
N8XXuyxjvZ1kLeD06tmp8YrNUSyPbpe51vH/XtZObFR1CiRvUBGFQxafGHff0eoE
qB6UiSqk2urIi/WvO3tHIuZfUkRnlBXvc/OgREG7m3UZzAXKE5HgrCE6PJSrYzNC
4ArbdqDcSMOw4Z48JiiNoCd71spF3qrtUuwXkKNbdW7LbBdvxfvYkIJUXti9DJkP
xfvgFbGRv1/kaIlswfpL1OupZE5zTs1N/OdbZuFq71FlcnZyKK0M02alZ2o4OD5P
0Hr2HAPeTzi+oZSvMXUQPagJVwezYm2ja/aMqwD0oosvZEsYjWtHsHNhLOv1i1R6
M5R4KaJkQBUnKTeFqklAcEOl6ougdkAsOXweb85CPXUNcmIDPQTHTmm8lYZ28L1F
7TBwP+kjC+uFAmsuiY944kjiMuP2tdFUAy8VgwQp4aCLx92uGZdcJHOyryKgFyUX
EHzje8tGTsshPl82fYpy7K+kX6dZZce9QQ/TSZ+wY7C9DQn0vS3G2Jb4pAninNbj
lpGvLgHWMyCByWH/Gt8kqx0MChkaDbzRSyEgjfWqUDG5C1vEAf91omyUK4luFruo
891rhuKkEvdyaFcqDIuhZDie4zJK+56MLuShVjVARrR7xbpCaDbqLYXkxF5k/qrr
jvwzhMMsJLfhm93T30fymS+uEM+6NUNMN0MP8gmpKOjYWpOLTxxhsZlacQU7nGfk
j5ycwoZyJMksk1WrTuHw9IE4iwgW6Q7px4Rn27hOmGbwHagbktM4a3E04wqZLgNW
WejD8932UTYgUJIrNA3j00WCiPFS5d6SBtstw2qcJ2gcPCej9Xo32wABLTPbHvYD
VwQv2VuCbwsbBzQDT2r5BHFdRI4fMEN7/elQu0roFHIZlG6Qri4GXD4u3Y3Qk2uB
uA4TbxcL/lW9lFMm3Z8l8uJ0A38J99XZdjKTEyHcEth9SFJ7hZdwbJs0TacA4/nl
vhSsCDC6x88ZiovreIibVtMQthQVlgYeF0ZqECHDDy6bUDA9x5+1g6Uo2Ab7/PF3
8JCQpVcy/fGrVAGYsqM59iX2eJXZU2nUjTIcqeBsCwAd/H7D0KLEPxoAom+oofmx
PiLRWamS6x0mLNzP8adZonfokFoggGu1E2U23SGOHPGTHWZr9zP9kbD19omiM+Y8
ab5RgHm5i66gttFSzDdTCwkmLH84x0WriOxzD3O2VZicDH5gs7JrW5URp3z+qImT
8Zn07md3SWu8v8cvTRG5fhkjKjfHgqcgAx3sJa16xAohwRNF+An6yDcoF30DqBri
OIMJendHw2iSTi9SkIJK9Mz+OfBz3qyj6UTWcNVaHiOXZ3vwgmkM5HK/NNFxr2X8
ZYwfpBecRrYXv4lPDaGmcn9xZ3Nfg3sATvbX2Fu4ulQtQ78G/lep+48vRNXVSYMg
Uko4ECeJlHyWMLR8anTGWrDWSvMpIexlkennU/LRd/HwJOxwsxx5rsNrtCmPpWx2
H3O667MZ/N5uHP0FgYwcED4AOI93/AYaBgkMwEHkd4uc0zE3f0OFlVmOKrMPUook
M5gYnbfKMDAdkYFWRTztmH2kbBcgVLweozAIJqxpXyJSRLijtDjYLqdKenPa1Pjy
vD/cjrPki6NXSUakVEUIynttnYQV5D3LNeKW9c6fwl0ulb3t0jWfVwXEMXpQCUtn
ltXqRrTna903Uy3dRSPQhjAkTL7GENkj0v6vf2kOIzmrNpJbifloYYerby97Pqv9
eTaZwFil/JIs6A9Phvz80tlUAzNqj5wMH8AgLYmZTbEfdgyMiGUDpWv4EZFVpdry
b2yWc1GWySQCARthOhVJGh5/P4defyOAZMi4AFAG1MsV+aEVkidyGW+Cmr2iXOQN
bhuut6Pi7eW1uC1UeXsg+abZPmtpWMRS7QL3EeJHH5d7rvkQ5QlhABU0fOFLRNX/
Ei1mBeVyR1x/Tq8WNOe5zMG8hH1/IQcv1eQfUYt7Li3ywDnEBxwNTy9s6a1xqKGs
UwaHO7VIRLqfoWMpEWe+2YWCUA9hrkFRQsnzrwDHCUM0SQpM2Sl7QBHJWLVcxp4n
YolvQlPKpQHE3hCDGy3WFXcUz5x8nFmFN1MkUACYF9iko/6xJPR9SGO+aVEcKSdo
lqOr7nCWObnjCDJkKX1FlWAwr+lXlkdek9MLCW9LNqEg6rke4L6Lrum2s9u0pMyD
+lp95dfkq3rYVx3TtDCn3ItSTaqbzTRZ1RwvzL9a5j2aXzb8McjvR1gMGTDvnksB
XRfQNAsYi8/QmnjNK/hVNA/EzRmXIjGZHSpUWZsCd1TPB2BF3hYruf1oh4lozkdv
YbPattgrN3+y+N5fdpqd65ak8s5xeiYre+a9EwBfXlExqsi3dA/VHi0L+eoZcwEm
7UujI7UpacClf2mDD2bU+b4OHIIX+7zIdNPTzkIzfEjuGgSUUGOwEMQa/2zoykT5
Cr0JqyxM1nVjak4YzCa0eT/k6HoK4TeaA9qMZ/Po4hZWOvI+ytoKwIGnh3QlWna5
TnKtujAihQ0IWJpYANRek0rOAMZf/gglkT+DkZlBlP4j9IVLLcPdy2YL7/orDFrP
JFZLGcjZlSqR24WVsvcmqm+vWPbdecOIn+pOMS6UsPD5m4s0v3FCHTMpEeRJOU1l
kxlnN6BVPAjVwukVr5z4efRzpOrY+Ep37hoWaQS6L5Rwi1wUY3NQaGYx+HLiqK5t
R8EsNetRYouy7iQ1xwdVdr0rnUP3b8aDj0rIujkPfNI5uWl1sby4ctGmzKNsZtqs
O7ocBNJi6Q1otEhRLkKNZi2lM9dm92hi6OIgVuap+ZgVlLp1du1zVZJ31yLS5waH
+KmS+9xuKyIVkjuNsHyDUqapukGAGLRuOkcX0GQ+ERBx33xSO/jiMwUrD3/ebcjU
+RKaBDp67iS49tCSEecxHdgY/1de7DQ3mZibHPvaRxUHdx/jUyk5UqHKwwNEdXGO
hkPdul/NRwRqcBezRUbSBUqfrMmk6UvsanRg6A7CauFcHisZBA29oGkX/BQkz6YH
suYQfcK81ci4g3ndn82fAX/M5b3ZeXv9mcffMisFlR+vmcTkeoXQAO/6cqkU1KBO
pqYpOIjd2AzVevYdQ/2rwBixV5d42LPJYtXBnI7OhKYMSSE0X12Ebtbo4x2kgpmF
E8+b3SSEHJyL3tRaiAh7lZO9imveUEKvi3ry4+DiKeb15xjp+YpCZuVLGzxBxop0
B3uo7XUwZBwDReU1pg3XnQFmkMREodUP1a1GLGfqCxzwjP9dYQRaq6HC2sRQecLr
Lb8u79eArXHQg4mHRH9lsj62q5nb5Iz2FiXft1CTOLoEaqNcoUvFxy6gilAMPw/p
nARu1CXQlOaFRDzB9mED5bP8mWXuocre3di9pB5hDoqfDDW7AkR+KaXEF93NNQjq
zGDmiMEi+brSb7SV3EaKCd8++iZdC64VaBuf8Qw0GGvZI76dw53fBJ+VaxDBEhuL
FbOu2LPczgmIasg4woRw9lViOwYGSCnTqVrcxB3dXvZw+t7TMYnAYXFdryNZQpMk
WZUleD0iHSTO8jdgq4hrCJ+rY9vJGXbNsymTJWcCW20Q/7HHSqNoMjBi7pzRdT3S
vDBknai62gh3nj8sr1zQo0Lgv0Y2Srtp9dMkgVqW/YthVWnr+MS/6Xt/JkYnvIig
TSwG8BA1qXg18Q4nD4wij67GrJdmi3OmjV9yTndGwGswbQEhF3Ioys8jbd5bHW51
ryjqIEWNO5j/xqvwsv9lzdt41TQ9ACCbC8yUs3l2ksNA7FTWeTtuK4uOgHN7guty
jeRp0aLC2mNmzYpyKYaXL9meNHAM0gbt92K5OW+InOHPF4E9u4PoofwNRJZQPp1r
K/l9O1ZCP0Ocvnt+OPhTJpi54UD9cmZQgKrR3rmd9uFXVHQAS9LOCKDE0+LheJPB
VJ2rVo1n0Mm0HdDU0wUOg07NlTWl9gVRTHRp6FCJRYYEyM7XQeVf/aQR9QZuU1LB
0RQ50tRRJ3GeN3eXDr0SnF76RphCxyuVy5tgwrE2b43sSpl3fZOAVVXBXxaoF/N5
CKU0dE+vV3Cx1eWTvzoa+wJZdiO3zKbrEBRpvVZt9+z8D9hHf7NWHxh2B4GdS2dg
nBN73urHRAzj2m6czSJ92U0pO1vGKF65G/eWbmxChvkGJn+kvjugBMQw96R5hXl+
/nKKeRpFDLOD/oBUUIw1c4sL+IpmVLt8obM4z9QFN4tq1oGeelYPa2IVp8yRXRc1
soOIdXG5+n7mj6+VOMYp7XNO5/iFvVT7Y0NDaaIFJDpElZwfDZ66uVVEEcsWxBva
DgBXlfKwVjTaG3YlAYTqeUu+zIjy0VLNn0CIG0loBF0SrYJg5huVxHXSoRcMEr12
LBJETCNp1gOtEf/bSjz4lCcJiy5MFSbSDog1mLzBaWw1Mq2gurJVjtqa0ai6rZ4a
OnqReqLAPHZ/bcNEUv+teyg6XbSysVPN413tLu7betd+PRI0uj4GKzThvK9y+/fC
m/4inQX0HMGHRzTON3lTIIUOX79+AZDkQiGU5JaDQK4yEXNR/CiQ1M3eznsLinQm
37QkMfk0dUlzDsEkh4kFwyEv1T7wBy4xkGKv5nl3wwn5YmvVdMfw+AEt7nTYLlKN
9RsAP83ooHnF97UMoJHXz7WFcLxqmWcyJT5C9nu0irOAos12AmW+79zmInZ+KyhF
T7fr2/Oph7MNNHBKSmR4iKhzwzmnXCAVMZBZSO2jxzVxfHsot8idTGbjJJd0UWU6
9E2xDumizGqw6cyxg6LhSGp2BN3/vAZOYbRZq7PmxdKMuzbc76STafrljIdMtnzj
sQK8c7tdiyI9NKrE+SHuQp8lS+UGOzM8HI50vkBDX3QhLBKSIvDDRKRDPRneUCgg
s7Vf3CC5CG8lXAC4lMjfyXfk1+A69QzZGBizm+qGIxkk/RXfL3+t76FaKza47EvX
UERGKPp1xebQYqCHqBUuIKJEevjM8eyWtsO4FvTql+E5lkMOVlS/aqESnwt89ceP
GdIwGDG1YACbA0yN5GrBzUr0chA64Vbq3lkwPcYSAmOS9QojhQ4d1t4ik8nMncp8
almdU1newbWL7iL2sL7tPeony5lFm+T/bv7J4CZHNzDaOcMF5Uz6UFx3gGTqjQRk
jXRsd8Q6ZxTJJRGC65lBYjAzo0S7eLk7TUQ+VagzDjOGUoWimnr6Typn/s5Po1kS
Hbz8tJS8yg3GCYz9WMan0IIw01chg7WOXVgLLbBRy4IkLWy8kRqiLqt+B3Z+LPZL
t7dIgOqYSAjDjyuZJihAqX19HJc/2FxMjNz7m3pHbYLKCg+b8L2vUczG+9+Jzj1Y
bUZeRySyA1ZMBi+ji7N4T5hybXhk/VGFDuAxb/eDdOgo2msqm4WO+o+dskp1HU5N
7u7GykbMRbXLwC566xv6zpgbBZ3OpgSfiCAGUVtk+eZU8y8cVQzsliJr0MDHlwiM
iz4HxhD01mn9asURJ6qEmCKL1BV3QwM8MSABMVxZtHa0AuL6i7mbqUhcI9wFsx6B
BzceLKQDiCQ9hqXN3s6P+W/Qd1usmAjltE/MO1QpcDaQenZbKbpB8F1UppDuOqjt
I53nFgUjMHadbL5r+6bjNDdQZqnuvinawB5fBdr9OP6iM4hLPpJ4IyurY8j6Atnk
0NS5r2xzISkvB+Dqj1PnEqdNO6Zl2hFMHJRlQTY3OUnvEZbHTGzOAZ7slbQQsmal
Z50xvW+RCqQ38YORc+gzGb+oLBCFpVLVjqzXLaJRb0NUvPGk2oUGKlHAffPsmHYi
aoGkaS/nqDx8JN09dE1hEk2caL0tcsqqtIlBrJydP9k/w4ta62WUowYmJsuQqH5x
LoJnXvgAE3wNm3sCuZrMx8BZaBHXyl4VHELm0/V18NgsRs1aczdz/LfS7FWPKRFV
XHWvn8v7d8OGRcPZ51Y6iexizYqyrtRKY8ss6LCxCE2m2101nWgtgKKiXP2Ex/8p
Xfl3yxBiAu+p1aJiyjn+ck6y9fzHe+rZfzvROXCj7ubzrxTHLIuKWAgPd2DHSG5j
D3ChKO8p5c3aX18NNp/VJXPHIkRLA9jp2ymBglp36TvNKcs/5Nuh+zFuBKRy7ejn
CxM6XjlxkaphwX90Bf2veivTi9a895H7H1adJO4D468nCwQZl2MYkcYEumPAVHG0
r7yxUbF2UlljKD9OPuO+99UZU257tYaxPXcGDbXpxDhI8garhtLTZ2M9Ir/flNQ1
iGc5TjOnWO66baWxk/+TV1OMhEqVD1kC80MhUaPUONPvHOYrc1KfLuJEm95RvEUg
svP/p+DFVQNMs4TNM1wgTnLQZxV598yrhSQwg/PrEh+W3g52wWmSJQ+zHg8XTbO6
ggnQlgi3diNd3TEdAIo5hQbe23m0OfrhkxWuu2BaM2NKlERxnyZWQR7kub/y5Mzl
vkvRNOoqqFRZFp8vwSsh5ADWv9qW9d9E4+pfsY8LRg+GBS+uaRk3Pylv5eCmKAE4
oeCeIcejtehIKbiAIKr/XVLzm03P4zFeM7HnOOyViT4gSuBubSgDWcs7RwoSvh8A
bLrA7I3HaQLXZFuVb7XcDVS4oNIJv11qll1BvpmUMI0Vanw1f8+phYk+/uwSkidX
Mt0guCvOu/AqwB6AHytY5jZswU8/HnCghcqq0P1ZRRXZ2VQhdJ1TJ2Be/0dMtSkX
m73MWYx/pM2aIeMFmgNdFXU562GL0x8vztg6sssQwWwGRGQeOSrxP3S8K2WzNS4h
2IU5rPU4R85cH8XTGdP5l851iold87Q9NQMBr4/gyrvTDEA6kYYdMSxl10o+TKru
U8P1sN4g6OcPz1RPxWjBY/zWvg0SC/UIbBPqHACYcVRkF9FmVT91wiIMx25aoLfX
Cx9JdQqAiRgdS9ujv3Rzwmnapb5F13egLOqVWv/Tm2xKStxAXUxZKnfLbssNDoJL
xtOlLhKu3bI9s/32Z6ulec5fQD155VcAEhU12uxhjy49kUrhwgtXpy66rI5tn7SS
C0hq+VVZVTYBAmXB8t7dT+u4ncZsrUF/noQU11EA8Cd/C87apCX4Z8wuILKEOXHb
s4AGg3SraCd9ad3CDCPtgLHrW3aNt+0EPvZ/odMj4/ZpLqs5quHJthffZpAU+fjz
ddWipB124cCHBlsqSAMaV9Xrb9VCblM41QeMGMn+ha7NMFfB7COMRfVKL/bmP+0r
TOqKUxqX6cB8+ffDYa3yf07B1fGrsFon9fuWEnHrC3AKbuVa5mJSz7U3Vn0bEly9
yVYhS4jid8HYeUQoJbANFUwS2eIKmIlf3rzOCRQNmUunN2C8nJc7IIzNlVoVPMhM
oK/cZ+uuwd+NgPx3GRdB4fxYbOAKq6umdzntzXBajJpIJkglBs+//EvXTyIYBLVu
lF+tmGks7c8b5tU4hwdeibqQuWwl9GuCkvNcwj7fTBRcMSZKO8sLo/MEq0UB9Xwm
1u2tPAGQBkJCnomp233xIXJLxIYHIrITisIVQRe/dSxq1M3WnIkQtQN6pGtUSpJ3
2v1uYe1MAa3tzmnYwc3J7vxaISRPqzJSrCbeQd/Tkx/KW2dl+O5i9s8uTWUgtCJa
j6ieoI9kuxZ/vutt1Jc+ZpOPWAL4XF+/9l20xuWsjdh2hSSSQlzjf438vxdgBhdc
v0j/GYf8mg2a4hs3mPOAdOLubHXMz+tju+A20ck2VzAXQpyGCch5rStZtV8KxTkT
BcP3Bo5lnHJ36AIZUGTyiyp73nTMFkdHSJeT/cwNZlEsPxP5A5KJeiI6i6xUE9u7
7FabAgNubyPnCvTA6jm8yGynL13YNSkUPoe6BWTEKZlKDLQ0FZoj5jN7u1p7ohX/
swuRRCIUiHtpSvEc1YbTi9FdbRp7MUhfdpeIotVyMQAW3muG7rwxySKMDJnqKxr9
fyHgKaI02j0LOzUwnqyhZ5f3FrDgwouiFvn1bMz5rXkcJhL5ZEz1y/HSOPryn4Z0
iajIDncQQhxPrRNl0Fjvs/cVcHNO4406RF5ON/V98dyL3e3RajQkFityeR1NPCbk
oko2OLC8W0MGB7OIb8y0PMkuKbHwX55XVIl9IPtV6MzFogXJM1VFOLoTBCyxCyEf
CnZ+njk+dTL555hx+jpImeAo4SVD/lropfTivwotN45HssoArklumRiwhaQb/McX
PO2kp+cGavFWFPe74gkfEb6+cA9kSGIN8TYqQ0RAs/ld8+BJGOcv34csmJ6baNEa
pi70VagbafXD+3lBzf8iKnaDEwDQvPzAZFNQL/J+htx/WeKtqDQ+8fNANIHT7INK
AIHKIWVOLNf4/u9McnQ1pBjeDf+dzapLm2sMfydM5V+4ZTqdedrzKZBFeI8laGkc
QJVYujKtd6RVBAOSZgj18ndxK0WmHBCCtJ5uoadwEtacNuGOUJ0gpynGWzVwUFOo
MsBiqgekKiPOvVaJsKuanD7iFfP8ttmJHmqutDvMgT2CHk7QF+k/pQAkrR+rIKwQ
GHfp+WdW6L1zAEyPXVuEFFcaUt0t6fCTuoBcKYIVIa7QLLQ5XyjqhvMQdA2bMat+
KLipCilQNavaFvQ6OKu6rT23fQanu6R5F1oFInvdUVY4Ageasxc+9VZI+OLJJJru
ZtW2x7Ak7TTxo7paS74Ef3cv3FL/24ac9WttDDjByIIVTKal6QlerZa78CppFV9l
jCOiT+aClE06Xm6eM6Bjhq2gL3VsIEoTXdvtQ6gXAXCd3hJwu3pCQPnVY5whMPAe
yDWGSiYcEitrl6mCuoCFcKKbio+GL9GphJNCkmiHyD6oCYlRmKR+wW3bLrMEoeK3
o6f4RSXwEeCS+vwrYLh0fcrxA0vMvBLbpHKmDzYuqpRCA77I2/FGEHlFSM4xuxlG
ToRs1mKCk1SU66aFspElo67dR0wIqpty3ZmTQgvBXadRlv3RfHNy3OVKa0t1RB2d
1Uy7luE4ZGs8WKlREN/2qQ+bYzsI6lrV0qZL6bvIxtWtV4DWrzxgYthL3yoZaU3n
iNmMXzQ/9gikvyPHNlyv6v/rbsqZBq2y0Smihr6iqYo/zO+weMPhhtpfz6SCWqMe
MjTo7lNpCtF2aWjbGuFrg0cjXw1bJDYogqar+UoQtLq3kHIvQWPdybVurhg2Vb2k
CQGlDiWBrIk39To01tC7R9mKwFRrh9di8K/BXAp/2XG5Puaxgj2boPusmH0690cX
oTzLJ7B6i+kUJb9dPuyLAogDuVqZKRKjRj9A2bI8Ht0wDehKgEJ5LZ2cyZAaPAV9
yDzewU+s3jeb194jGjW71jbpNwX0GhqGu1ud3iRPcGJphtSEkFGylD8Wf0hPjNhi
PYyLH0F57/ppoBhWGKhAz0Te6II8ljOwSpJUrcOFkaCLWbz1nlncOs9RO/4tbZwV
XXzvluA1gHcgnxRu+jU1lG1qBmCaYjCcLAT1+cGUSboHVpPu90ObILH5JyXtz/ZT
Pdt7GS3MYvBRH1/cJHVDzMKoK63zQ06uiPWdVSv2n1RiVZL7YE7SiHb9yn0fCvpK
Xji6tJ7Xw1oGEOrZTbmgYtOeleV+iBlgk5JcBVhkbdpk3uHRdmh4zuZo2nwWe0NW
cMvO3kU5OEhh55zkftZ3y+h4hpN93b5I1po2iDuRuKbsG1in7RuDzfIk+JIZajBr
FTE4R2P1nBjeLf6aPfaNxu72414OPr4lqUsZbbltlgHwNTkKgAuGA2AK0So8nH7g
uqA1axPdQEg/2oWDlGIsv48FZee73YxFXX2LXClfP0CyVhw/F5oKcZXexXQ8aZKj
v69il1pmFCaoZyRRKQfjb7B4m48lJB++QDSAVSvepZvwiarXnpFDmq4GE2557KpR
/TSOM/k74eDXlfMbslbRv5mul703SyP20qCP+78/uhrzqr9Qzn5sgs78UTUflfXi
H7FPLtcR9Hq8YrjwPhIQWU6ZNhqX7i606bJERRwYupuw65I5tQDRK1mPt1hy3U2W
jpU2ei6r3Jv3N5wmcrZC9wVNh/yetXFHioRWwnyMEv13/qtf3nbvIDuprBRH/VuM
THo/4L6+mAvUZqvMXwAPQeLLWgawRA8bzd3z+OIRBitLLPaCvuEmTOXiP/JTaJTo
l9R3lJn8Y7uZElFkJuAqYYmO6nP0QjWe8k6Em7qCaYNcx9DBvEjZi3+XuHciIVsF
E5uxABIbq3chJWgO0CTJRSE5GntlgD0Uz8Qrb13aYFF7zzLVFcfb8k16kpw1pgv0
HC2XIXbHenxCJI8Ditlr81RfigIEUl0jZ42wkDdV4kKRLBA09IQPR0yhVU/8bb4p
D3kZu21bD2CNHlxbE/cOehhTouW5Tuvvj3Cpe9qKWqsJuHqGeOfUYGSBgQ/LmgrG
YkUhZrGTixgFmEYm4CUh70503snWvDwVWmGKplOI2d/Atytz+ptmCseH0/Lt7fOA
fFGKINltDvRSKPXnxsNzUhS1dlTE8x8HteyQQt8I/Zwwq749e8pV14VJvv/PbCbV
hUJYoA1OoCYC3wmS4ef5jT5bGN6CwzPicmoRq4XAL2Fj1GsuY4lMRpVmDctnCwie
w4g8+qpxxcSkbzUw/jpwWXxRggJYXVxRdID152CH0tqYbgRvqiWOzEjmQnUBgrLf
U2dRF00oqvsQBlq0HG65qntP9xWuwLNaCm34llw8fg/LcKnxzbtBzdHgvITb6e+C
gcI/4UHM5F7AhZ5Aq7Y/PwHa7Th6Nt8rBkNnlqrV4mdurQT+L3LNAv/puqsnEYXT
ZRpFgZKs9GnB4boCL+AmUKyYg/2xTftLyCLGcH5u7SirR0LSwCN1SKerzGFD9WKP
RpaEoQZ/Tr454693JM/joM0eueUJEa5IrnjGXEDrvCnE0ezfqvGEBkCWuRZ3N51Z
qVN9zP/1domEy1tJKhxm+WjPo3jj020xdctmdMn+AWZKsMr/P5+tbTxE/AuDHrB3
FQdQAHX/sTpT3EfGDFvnYr+VqZMW+EWBwGfzV4B9dx0yBrMIfYpkZ59TONQ7bIs8
tM2m3Q4lPlzAH1xLgRcduMaZRjDBPmhWojh0WT/asW6rQz5nH+IZr6G05fbbxuny
K9rMjpZQWWzQ9nhgKgUDUTmoHQywfC6Y/fKdmgxKYyj1lTWWNIT6pyeJWqgugYDA
5oUFasbkMNZtgZdhBmfZlImj/oojBidJ7K9+hXUiP12Wd84xKPfYMvxcsS+9w2Tq
0/trPXewf6JdWbICOkdSThgycEMyj7o+fNe2HtSWXEXl58dKYFh8wAxVwgWFio7O
CmUN94TJ1ZG7IoJKEnqW6Nkt1M90fdPE+VE3iKWjAPph9+nnt2/TyZOs0H0XW3+6
UMUv3js9WM5R/wd6+++7cezZFxnBIFw7plMlr6J3srAaSz2ToC12jdyOwI9CgkhD
F/b00zSbcmsPE9ij3RiN1JUFe52GTHeodN2ZNAzw3TTVhwEOPKLPwmYpcZXA4+G1
b+3hzUNGH5Zz9IPkNmZRc747V3OBAjbRsSZAJeBOS07Pu3Dz/KzvUNbcaApDD+68
IgckBSOJNRYNgoooNFvaspMl6HY1OT17aW4c++8TDil/DgX8t+wvp9YO+zKszGm4
oC44RdXZ2jfo1sSk6f2IlLZj/adx8N7iGzpyFEkTFltURa75oBcrgYxPATHTq9Eu
4jC56vTYZg9iE1PjBrqgCQzwQ3l+XPo8cdyRPLIuK9sBndo5FHWoviuXE5SwgEKt
g79AMl3ZckcZ/qMHlsoRxVwI0Yrg+baYxqUXtNjsr08a0kXEEaRl+yhm8t7+pHcM
MN8nFOTc4OQfuy54gw9FiaCEuZ5TYopJ4tZiV3raewi3jB0HD2dnI/wdn4AQxxDT
5JG+vuN2KUe4+1+qQCyosxHNclv6Y3f0s+juXdcVwK0fHlLTRiHfDrgKLBhW9Kwa
I9Lv5o5HKxLk24sRwMxztdnyn3Ziy5U8NgoSCVVhJSnq9jBtXeG0UnTeSildiDdu
LLBiULPf4uu/WAUlHVHU6pNLy7S/8MxXC2y2Ilqia+S23Z217ag9pQ0TBPWyvcQT
GNrycGFoLxK13qqPf3fxg3SJo0NK+/fk78OIuhq/650ZLq7Q4tou26WVmFGkf5fo
vBMRQv7cz43K1p59kguFfDcGHtqMMqN9IMF1cDdz6AcMdRWXt4rTOVQUCas2RVHn
CUs18ga4IgTqfBoOn171/IzNhN9DNrr0Ct0LsuiRBGHlDCBuBRMXW1WTp1DIoy/S
vF6bAjjVqy/OTOrfzHgdaq5fgZpm32URxtOh8ep3iUCquA5aMZdUMvHW3Wcf7zpR
ll9QOW/pO+TBD9aIAjuR4lgOIvK+OAGtGqgrC4uD6sLn5s9M+QzcdvuNO48WJdsi
V0tDneG51YtODZWZOhV4ql+0+8TkHFktUFy2TsHt/cVBRt/FSSFRNtpguW48o49y
h1hP5U4EK+PwoWMRzmKv56HGMYvdb7UzeuKAqkaMA03fBdxXxGfCp5/ciPQAU4Fc
0NMPNN7Fvo/ZMqPe09aV/pqxD5eZk4kdOrkAmUgGfmxgRS7sd2EgMloQlCV7XyCv
18wmChchXEbrj2TUwvmdOMDfY8XhPdkoXO1qMgxCKPP9WAghHEl3kdaftypJcugP
mToXfQX8OOsJF/dis2lzcXi8608/JZfC302rw01s1m3IiuWTFth0h2GiuhmKlTI/
+8soJ15N+/WPNuaX2vNRHUnN2CL7yBpboyvm9LWMxvm+E9jfA5L23RIPmprggNti
AVvt6U1aDiJv9wVHIMCeVa9OZF/JFu3ZdT7DRyAFEgCF8/kxfdHIO51nkMtDGXJo
lMjR1ge4qGDdkQmWrSZp7ZVQ9vJkx5a47b+EPloq76KYXd8KYTS8zFR4Jl5YOCea
LLtGgo8sTQ4kbMcn2QAA9GRkwYcIsLmJucABSRifJShl+0kozmqA13l703VSiK1p
p1/VkLNEweREgEvSim9aC4TJsyEAkstXdRGg2YCoEj6k3pmxChkmatdEUJM7gSPA
CJ5kHq6B9ws1YcdI0gPcmI2xpZhYiuNdaocWrUZko7t/QcVAJlMhj3W+bfws1wbj
zXEEYNo2y/lQdDPzpQoWUisbQYP5OfHC/5jFbCWIqzFKK3EuZP5HaXlbhPs7orrA
CRIGaIQ6HKNyN1/yCWesS8XTOngFCzar6V7HtiBRY2mpkZvFvScZxMJnwh8f+050
1C7DbLCsjeyGFmyK0yCeWPyGS6iQobOgwSvl2srmcMz2lAqHqNZ8ew5+1dYsRfJB
d5FEcObuuckRDMcQYMhRtR+jTYS4yUBIOhuxrT2pjwgx8RGvj5Hy48DdF7LPwEkj
OI1PkaoK5hwpqu5Kt5OLW0kexr83UJRCWbAc3zWy686ucyGETRn5wXDhllE3V4SF
uIHcpcOkzRkmkxDpu1UIRfrlNOAtY4nCl+8n7oFZ3telqM60KQffENEAJHCswO0i
tU2L5g+qk+NAejaxSfNUsj7mTm0jFX/xM/017H5TCOOjeCofzg0idfO2A9gyxEbo
ZIRtiF/EE/5AtwLZOmeJ4nvam3+qwr/qpL3ZHHq8es/m+qu1v3l6jJcrcYfUr3BY
DCsQnh5Q7lUt1yYOKAoV6wL+o3EMvGJTk2SaEwvNhxsmmlzGAhR2plRY6pXkEVJc
ZIvQUTONWMkqzG0c11DGVYd99t22D2l0m0gsNFC/BCVV0tjVy2xI5IEMUztrz5CS
voVfHRpbEvuly43ieU3wIeTEFKcRFVOdqppnuwf4Ah/cTi93a2BkX8XmEleMBPpz
cQrLDUaVQNy7gG+bAcg+luI8lWjlMWwAwAkxlu1S33+GqSHDgB/8LT1OMiiJG3LX
1BNaGGp0mE8hGz32DLJtP8FzYi8s4N8jheP1sS0onrEANWls8fOhH4SoK0vb1cId
ikcGfB2kWy+FTdu2xl45QatJKW++HJwDwecvXVLheZI0oxCmYqMl5NK8mKPYrkQ8
zE/Aegbt8XPetYBojo1iJACIWRLQTpaQr4hHTj3xaGZ0uUMINEbQH5m7Xbph7BfC
lVQSOv/INF/Hexof066S/M2jfKaPNIAHQwaYGuKJ06ObMhUQ6+38fWYfoHOPDYOw
rG2xXMPnGhasXs89W6cYDNcE8lf+NBdPtqLlSR54IncAhgF2ZqLqOwBecnecuv9Q
ygIxKieBR2bShLaOLJiCuJF5a/y15f/YPOkNiJGS3rkU2uYnQX2MxMSdMTP/Q/7F
J9fr6gE3K2dvdMZ/ISqOQ/KtcrFxaLdWW2ROrrut5D0l2Amiw7qAl0t9mvOJhcy9
i7nh7GJpboq6imQc3YUjcWKYpxRk8o6WhLtF3eY8RydqzmyiNlSAyw5dmv0GJHL2
zXAECbwPTIGc6Om3xklZMbltn6F5Mr/XHA3NIYUGdKPXHfaF2eUg/ZePZ1JM9dA1
e3rP0uAPzUfnwv1zjKOU9QBk6MD5cvtO0GNWZTnwt/7vVGbaRusOEx56o9NYBI9a
tgRsLJCFzqrN0kzSjXivytIYIw+599NKPpAJBR/4KveFTKGR/7TMHnP/hz60tCan
PkEBkGqPKOeHVyUzUxMFSrkMonQNYxS0SqbD57PC+iZZfqQ5C57FHAFwCsHqRZ7U
Z4UEFhoDz/e0OD5prSbUWRrcmHizg8THHcqswxG5paEm0JdzJXb1ZHXKjW8quLbS
mKItft8D7mLwAAkPuvA8pApESYXRewdXNCO7mN+c6NuiMZwq0+tIc38fNSdYitTY
z1e9el1d4+v3zpKpaJG6j5JtxRqJy8j6eZU5Csk5IEAMBLLNUYf9y8gy+cV19BHn
NmpFK+xfijuLs3DA/t93YD1DDjjuztian+B+QoEvUCMMNXQUcli42Eqb1wwUT8zg
Ya/YiK7Y56SjkD9fU7C5gmz9EQ0zSMNq1hua2/OvRulnePOqB2EV+GG0KxAArr2E
ZR5IsOoPQZ2PwU/39gg6vGfSR6TbMwHiRUo1xNwp8ecwgOp0Ug7oWgzi2vcaDrfB
koJrjAcz5pzUPuyl7Z1+4UuiYOQfgVdJ6MfaOn5N9xg6NBzikIeyQQHU08spN01d
xW2+WEcc/eU5E+Q8JpNtpD9lye0eJF4RCDllgZFiCwGJ6DWqtkMntGrLblncegek
CzeieSclTGQ73nfjCKFCMUGV1qwMjGbxM8HgLS6HLc3YJBB0rdLKzt9qsYu9ILgd
wB0/5kEkICS7jUt1BX+cCRjw9/r3QGOq8OJG8IfyR++M1VMVu7uB1/RbY9NH8Kkp
pMokbTXS9K4cwTI/LQXilv6XKLq1deziOI1MD3+iJ3F1+t5shxG+ReHmndumj/Vy
ji0tuN9kqToZDLdunSd4YE9DWjm6EQdcN76+/gy1M4H8kHIeoVsXyyaMC7qomZWK
dtreJp9ms+dvFnANq8Kl1k3bvu4cKYAondI2OqIp4USjFUM1+LJ3dAOKj9fmiMXc
BSkfMxzIz02UOlZ0WV/JL6KPBa4uEyOceTF7Sven98aIMeWQS8xk05P5Nqu+TXqX
lrN4oEVrPHyHH+6advQASaLJTJLfbePg5Z6WHNijKmREyitZo4/yKJrbEBA65ZNn
Dt8HX2cVhICSY39bgGTMle/fEcQlFYbl4rlCbAI6uyMYYdbXFLc8g3CFQoGEEi7q
IOK+68rR4t0474LiXfgTsAl20+Pk57vhoNhumG4Cm5C0XAASst1btUtsXvxUspk3
9OY4mQcVSNUGCHUGh308TWUW12HheAmqgYH8KF1hBTs3vE5q49anDkBMYHk5ev/f
kfrk3EKPrvsu2b3kTAe6PpO2xzkVVR4HKfkH5HYfe8uqf2v9NalRvpN1Wbk0rPW1
QxoncIar18M13Pz5csfxQwLmHPfjegJeV9GGLbBM5OUFIZ4g9bDL1gNtzh+aT8R8
+3xKwrm4ZvlnMQw4+qQsqPqtl2dS7sFchYtDRl43g5Q0065UTw2CM3d7jCmffyHi
YoG57hL2nG6RPaBN0v1l+W56vlbJjnIUwRSePfP0wwAUVvc3q8/snqNaVgKuLPac
cdSSjZdKQBm/Ni6kutpLQh7Opv/CtGcNuFiTeLXMoaFPVUyIjUTMCgRAMK2LRMzq
sK0Op2lnggLS773CrsZVGO41Tc11oTsUkjUCa+6YW+169mkG9a1mnJzPl7xv+3Am
M22ZtJA4ofHWLvNqKD3H0HyY7NkHiLE6WYmTZoJBkbFjRfI8+CeiL9SBipjsN5G7
woBFI6YQ7kIdZZc/kjSOY5pzVjxrvdDH9M70UrW6/dwrtevA/oKGV9Wu/m6XWiCM
2/Ca+LivbOvkTfM/rnehGZRt3OA1518mOEClxBCkNTAQPC8koLXQr6M1Y8xzpMdE
5KxNJ2xWw8ghK6nxuIKGbXKM6tGviBLQEPVtx5x1pDN9Sg391B/k0/vAg2I9RxBF
g3nqrrS09ZSemV7HcK7wP1zKGFPYkKKDW9D5JSmHKQECFboueTqx7G/gzKotvX9/
hnqBY/vOpYMt+hD8KEeW6ytMhJimBXU6pbRlZfntAkBuaby6Mm33LzDHFJguYQUg
YdaJ/6zFdohlhMkF1dfrwHV0aCDFeq4AXWLeXmD7pKJ/J7WMe2VoLycVo4fCM897
GvGqaOmDeCqYx1ixMwIDtvKACnhnVod3Bty6AWGe0HhuKaJJZkkqr/xoq88MSOCf
UA3vUKNAHkI9wtPZct+pi8POArPNcTW0J1FFRTvZijuk2AxfeqwV7jIE83SK5FxP
2tfBmPqaJB5Lh5mWJtst4pgg53ND65+my+UCiF+o3aNCiXGmouThZNWRYukwm5Zt
FnkIjYrz9Er3iTpq8HaYxqZ7E0T2u+wP4GkB5aWWceMeWNYUde82b5wPVAVWxlrs
y76d/9noVkU/DLma1Svr8pOgy6y4nRa09k1rne1Ji3jmDdRHepl1qYvXR2IW2kgd
0fWmSU8klhOVeQxeY6Kj4lnsnbxWicA2DhZLYGRRrAFmm/7AiXrhxM4Z74Z5onNI
CcrgoNAOdmaodZqOpdcRTlrNPma3jEW5PoZMBPCbV151bsJLHuXXdxf4S5S0vgqI
Zk9PbRaUVWEhWN4WIk/9Xs0xbi1gcmmtCejoT7Qxk0/GQuInQvv8x8VruSq5aAAk
b6zmBSHfTR0ZfDw1zCJG4+LM1CeG0XFELyk+1nUNKhfX+vj6ie8VQ2k2XCa8O8ES
YgI+eD1MdEmxJbUEGTSZ37+haHq3CPzkRFczGCnSeBxOcu3bgb8d0wxKoI7Lf7Ne
dV3hFODxT1FWKX5zOtRvMgozjHXv0sWsZxD/Sf8iPGIuU5bC64Q7Q2HHagNaYJXH
6Yj5POp6KvvJwfcJdJQaQ4kQKqXDgyvQyZ79Q5k5Cmjn0jJblZIfNt6xMJDDHC2S
DZ/4WUMKseJn5iBvQNKxCEq9dJp74NE0Wl7S/kyMEWvyu/dy1Q4zUJFyfXlkTYCv
QDa9EShKqqQtofdplqmNWrWDxp7ltTISIsq++k5cd+fg0SZUIdiqmPv56JOMz+OE
b89eEVN3neBYnB9uOGTeBeVe5WxC7d/vlmJsL2TbbRyF9OEB4g88uop3E40M62oJ
bzx2r1/WhmJRb41tBtt5jL8fw6p/c9rNuZuwGk1fHf1g2l95vejZbOewhSDkMACF
bd8YIlsi5KWsT7BCvchYD4GLFlxnrQDizYltgr8eLR7kfjXc0EmuGAtUUhMsk7iG
zD+sFpdL3e0Shh9MnS9+qYJnXdwEKVTaaHhml01hOmxogf2pCuXDfrWa1SFJYmg0
vlbDW3U1TMgIKWA/vgkWcC8Hqvb/iHghO9pUKDi4rC6pnp24Nc5Dz469Zep4IAKk
4MfIviMaR3oW4O7nlh6RfwTXUOizwQzGTYUFHgxuGzwlOgT3wbI3WoQsVJKM3n7k
XAEMPtzD7TfUVSUx2HI0VumoR3o9UYUv5VmImutnw0Ny3mTwqA8v/A3jGTs89hFe
IbRgQXjkKMSXtE8Vf4UT6EfQNTDt7pz958rOafpIfcTNfLOweebyf/nsOHMbBJvM
LJMQAH090hGvuBpyVGvrlNWztPI2j7JaHKHztiUKJh0DFyRlS5E/1vn7N+Hxubwf
iILAuZIZyRYkYCbXaTRx6GrVeD1e6mNulpWXC8aDF5hW+SH0tNMVrJGp8yNdEoGa
2KiHQQMVTfTW8iXXXhfORh9xx9ixNu3a0Q0I2kZTZ08oSHjg3KuVbToXRYFQH/BK
jZWJkC23yyle3UpGcPAAu/LB+vqExwAG5BfAPV9GiUDLGF7MSn/ZuqiMbeY5akaW
vEF6HYhFWyUU6tye/IxSLSO4J6uzasaNks40uMA/sPcmTQUzMPb0Opz4jnVNyr9Q
5U2ahJop30HGTw68yXpUKHZXzzNFWNb4b2IIfP7CoZw4GS9BQzPcUmHzvLIyiBYC
csLluDAbT9vAmxsPziPQDUq8MCiKhfYbIVJuspJ6HFYKT44xkC4Flo348C/Is0NC
Xyl+UDQZHx4KNOiJu8DfSEDjgBnv3sivBmH3QwZPB8lPGSFckTHeXnMEQNBBOfJJ
4VRym0DyTzNPYAshCCMrt1k3EGue/D+S07bLBQiJbW8e4tGHRB/trAC6GgAcU2GE
daER7foCj2zZ1QT5bitBlUfJfJEAt7U3/HiiJAdK8Nwmu1yPwK7snTRlBo9je4w5
3M9Fsx1Xenjh1Frk88IlfSN+Bv/6Dd3ZDmdfUGfDE547jYe3eUoEek1K0UkKzbJE
CBSP/JM6q2kuyoJFMZ/Y3vl55C2Qz9VG0JTC6TR3HG4lLRtDj5IFQ4PDvCwX4a6F
tgyD4S9543wtYFwbZHOrPRLZGCTkRlUloL4dt0Gq4UQI0+xYcO+ctKr8+LXG6c1z
odlellPadAc0m2ZVp+nbtAz+niu1K3ATA/PEEor8za3PtIm6u6gOvreJmJz5PN7t
iAtU+qUnDHAS2GMcYjmxsgDxgy10a2HTjPrzCbEVT1YfhwPC03KuA6CrjPg0gyky
qS9rLjITefocanpCJV0jxZBmBT/bo/ss0/MUl4gWpu+gJjAxJPbs3KWrjLT5Q+3e
8BOAiqUFh1oXwdGdyEJ1kUhTZMrzcI5NAEH/a/k7HljW1Q99qFw7kHmGmUbyfNS2
WZRr0gjv7xqlWOmzd4MxrhTFlmlD+H1pvi3LF3t7eq1LY9mROLe/c+vnjM+st/Uq
1YYEhyOVrjOGgVjRdWL3XNHD7Cp3V4P4QCbbyXIfDppLqs7rkwMakWfwIAHQ4Y07
W6apDZvfigWnjRK6IUNSBP10Aa3ioZpY8BYoH3ycrVT6RgampeqXiIcTlk7z+7ez
hR0cBzfRnyxt3dOISwKPOOrMbsiM977mgRTB3GqhdSwBSXiIEWucYZIZ8WCb78C9
dRWnMEsPe1Vcxq7tGowCLhmurhp0chqQRAQDU3+eAm4O09wf6eRzeK1sABzxT1dO
+rgbzt5tr4RcEaDWCEgfbfCkRIzZbkZJYtqOOi4y9dsLXB/ZTLKIDPR2PKXN/iuu
AwmrhSWCaS+pqeM2BMzGB8MyR19Ofoxt+WOUSAv13DHzmpBnQBrxT4wntGEfdvvm
rdeZUCK5wf6g3r6NeOK2LQ5PCOD303D7CkCujroepk2k93r0EkpFKeX2kYc0yGav
b2r4VFiElPy47pW+aOKvNxtVMxbcJ3Qm9cd2DOdDg+kroaZQq5USzUJtXtoudUHi
eyoWTOYH24jX9xR5wPNMLmBKYyiGJUZaIJpAktvtXXLv3NS9ftR1fb6ijXdjAMK5
l0ynnEUonZXPEbpgL+KJRP1mpczzl/9Da2A4+6p+b1orvG0NG5fyEla91lPghE/T
BpcNWc8/EEb41zGlqo7JEr3F3kYRx0EAUTJP62uY3e9fWl5vW5oCaoaXDMM1KURb
LnXjJ4xR+Su98FaSB8Te5XZ7z6Q0LHVl2ptZnmYHn0D+ji22mjUGlNxRdG85esiM
ZYCgV1E4gJndlazrF5VSq3hpc5cxloKQ/gpxd8sqHoDMjXrxLWZsGlVE83KphGjG
MGHcZbJcv/2ToiNRv/Owp6w2ffTz30hfd/VVPwIziryqW4PGcRdncrwbQKmjmrVD
sn5KF87JQnUVTU43YaoFO03hQpS90hHGsrmJumwm3h+hCg9umHr3ALQ/YDlitWa7
BjVt80o/JJSzrrmh2hupQUo5WnL+caSAYs6vC404vVP9B6efi62BMtyWBTqb1G39
k1bD/BLue0zNUSo91W/zJ396kRMel5Yo8AoejVvyoQxleoHqXj9lvpJOSiKVW1eD
J5DK2spTH/tRuwUrTAhcFZetOL6rtbVAr9uOTUHUvFFM9tqLKAjY8UC7XhTwvMl0
gTDU7izq/l8YPgZJ9YerKJA5NInLPeDGHRipZHn7dR3oDZoIyF7Nuw10fCD3H6oe
0lSYDqhMAg8cBYa42JCxi6yAHk8SRSeeLdsyn3HbXnU8YbzctY7WD2jevmlKNj13
FiooGvQXylZvCPBd5k7riFtYjuZgEoA6ubhCnzaoUQOfTW5FlS9fVM4CnnwhcL4H
IcflIzYT8XokeO4kIgzK1CECwqHUi/V6qbtCdDRlwrgyVqom9xLRjM07dUsP7sQB
h3TmFaLMtzNj/g3+V+OogGzicpmQ5mO4PK7EYY5xsVZOIGIhTV91xBEdjJDmkRv7
nZj2JUb9w9/6ZudB0BsB5fMjQhvzanYO/d3+u+lcsHuO/SSBioeBoYnIxWqlsfgN
yNj1ynkHrEIPouIOuF1HzuFz0tW3f9oD78v/Qm+4XOfJrsV+1ugf5cB+PTtan+uf
b3htxi1cfVZ9Wz+czMokH+JSjW5JmwmzZb553oQLmTcHc+nwM8fqTs2DZD/3jk7n
hd7jNJm6yRfmsQ4VStWB0nimytqpwUiv5DvjIYpXAQ/3GTMQ16H9TTfV7A9AQOef
nthd6qJ0EW8d18yHWRQ4QNwGV1sSbzn6MJzxkzTpcY6hWc8OtN3GSpc726NQr3nl
Fj3zubJP/eJLaBIqaDk5mZqoxqbVi/r+K/6+NtIsjGEBAnE3+EpKSJ1qG9kLaaat
07vVHr7qOjmRxRjSW8rXMNDr/i1cIrs2K0SDbTrG7VBNLFfuSolO55b3XDePoN6o
07zhSTR7FY6FqpGVrDJ5fIizm3jew4aMcQjbtyNg1vP5vbtFixF6OlvGEzLk2e/P
cEZGVhdapbH6U9JBkPeC2UraPxgWvi2Aqy4LAKZcA4DV/owmjvxSVbb2yJW0Khm9
9jf/PlIIVpBc2vfJOskVtbHPLz5j/BZqiMWPA4Tg5IESXRiM/frukJy9svDb7de9
imBA5cubS4H+eNSzZumIwYwoeOslyYJT3kixv8d8iWj9nlbxV3PDhj2KuVqUq9Ig
LTTwo6A9xBRTstygEYbkZTDB9OAj6993ymW0EQkZA4UJIhGP4n1jepRe3zbNGBi0
dHazmv8jINMav5oshJhqDis1ecF5TSmmu6pnLb+Ok6+XXEveZCPGiNiYaOVtNKWh
+7Pi8dMDAl/YZUC43CrAJEBDVu2kAVUX+77dGAUUy4ihx5FBeIOG5V1ytu04PM2Z
uoMrLTvQV+NDvhBPpVk4bDtJBvZonk62iA/Tq3loQqwKVpDSKFpIwTTKd18FdUXj
dfD07i7+gDpPWnf2qk26pYb6lOduMAZNzvYNsPFCx8lLn7rLHmaq7OK3B5vMLcYK
VfyMww0ihMGZIYH6Epn8e03bSG1nnFkV46lFgw48arX+079AWQaMeZEYZ9WCAphR
K5mvqes5keo5t2jCcR4UxPO2wCdEIZMMbgRd5mk1sFL63wY/buMOzDo5k34WXh48
XOZP1JgLQjmjWtDlilJUJV9HxQfo2lBIhreBHgzSyJv0xGnRMe2Efa+LvfAczPlW
eJP7SSR67iNzk5Z/142U3FBKXEkb5/8Chf9AO6rSxeVu10ABsQf89BVhTywhOf03
Urx60s20OjJG8fHTHYNO2lh16B2C7gR6kiZ3Zh+7440l0GDmzYNHvjdCz2OkDWff
f4Z28tUCQlvZCMHN0VFQpPjGdmgwkjDjkEUIe2W6t5gh8or6UBbOwBIPFF3dXoN9
5iNojrAla3qfD+By8iny/5W1Tc+99kQhDXGnz+oKE9NnTwUPuBiusr1k8dKqltPj
esKAGC71ZYnY/eSCWCnxIbtUgXntiLcSKs6GVskpiJzzY5G0Jf3qgIWgrJ4eRb3H
LbxEOfaPk6VbtfOh4IiWGweatAUfu10dGyju9Bqjm6M29ooRPtt7wIbYbdgajykb
whvRSDOGPuxO/cPKl0/CW3gkg2Vg16/WozreVqDQv+8KAzvoWcMT+vg5UYjLbUKh
LyqxpHIBIZzAqVteBRVKWLQH4ESHPcpo2tLKjnpHM0u6DDrRJKeY60IutiNw4jCT
bJphE2OATeRtCq5lHm8vJyRU+/rfktsIXIO8s5uOyKvAKkwS3aC7BpxI9Kk9bvj2
LQaqmrj+N9AOThzpUaEb9n7uK23Tf7x8n+LpFNX83693LkA4U7EnWr9g094ZO1Ml
IcUV9AwUmOEEwfhtIGu19S24zHMf2SZ9Mmujgj1pHmp6UJaQ92WhalT+ld/7gOdc
b99BIsveLKHfFGcD2x4Wvra4z4UULkHRJvJ8EeRtJALzvJ1/Qe2yRHpvG+e4GX9F
0FqlFe8R/36pqX2lZdGHRCn4Dv2wZm9N1uv367FVeMYyjADhjb4mp9i8NLCAyK+L
TBWZGZO7ig6LWyLZ/pcklXjJdBYA5GNnlTGOlKuB7OxLPefYeWxs53CCZOiFTlKs
GOimfjV3bvu/OD0McvIyh0OZHmhjwSkKvRazefdxZvFthOECFFYdttt3y2hYu0k/
vsHe5YSpWvE10A+kZnOgxg+QzbxYtzH3FVDdV0HcgOKj+frCNh3VKDLvBdA9yUYy
Xj6YQjfd5Q+zRHy4Agpyyo7sXvmrZfIFUxX/dWdMmgAUpGlMJ/SiFk30tS5BRFXn
4lbBBzvnx0abAqT7gqtWLxQgKLh+FxHBfaoKoRlnn2ZBAARvtRVyWd3GsALc4g9b
tHf+YDWAQn+YWnCjGmSa6wLJEQAphk4CQTc1NYy4SniDzYU4GRRCKOg+U9cjGbUs
u36A/nBhdQ5SmNG9Tn8oK6HU9e7JvxdqlPiIiPVCO8h8Ff9GTQyUg/GcGUZgfwqo
n/d6gBKCSlE8fHwYCrUAsTosSpXv0QiIwUF41EUY9bO54pCebtVLG6AOJOAFLCpy
dmM/5VyuXhHaNFbYHwsWK51BNXe059YEa6F2Yn8w6WbWSoD5NL34yNvzyxNifi5r
OHsAmdkYyMryjVDCJBSeRJVLeJbA2Xz7L6QBPy2c4bkMrOlOjgpmvbWNdsk35j+M
togtPjPeoBsY1pIhRGx/PCEJ0MlEmjv/A7nU+ARR48yyaGKLWZD4OJJry/xfM3+o
eSLBQltnUwaGTcr8np2sEHGYFIHb5nKd+M13q7f6sq0oa4o9nTt4on4i2/CpIeLZ
60mQeKPeJZpdWHKKB+BeDBzIep1w/dmWhGDWKG7PGTNLPkw7XprEbHT1AJZ7KTT3
lyGmccS4Hw5EehDlFH7EKylH7WyzhFrn8iBwnIdwdYaXx+lgLDdIQssrPXcXSdIg
5Z+qdtCjvXahOGdvdzznJj1NsjpyEOI+fNbAc0yDVrLbM/uzWPgLoExqzd4Ofxg7
/bTt4Tcvyt4pym3J2JdimIIKtJZVpIOcIUPUG5M5GiWX5281pl8RoU5TFyXpFMSR
KOHAPUCHVlMpvyjLpvIBetgQboXzOEXGHCN4YZNiN8jsdg07wHWK9MvKFv+kXhk5
21oNbVIagbU3klZHfM4NIz1fzJntpOv/x+cfsxMAV45Rh6QVw8ldpd8VTotybZnn
coG1rQ7UquL5XNAI3mbdWyl5ilPt2cuhUCZvyUL2/+Qc1ALX9+kdOMyUIP0QC3Io
IkL7miTJZJ1evu3xTmxNRk3zIAEX1xYj/fCvqsZxOYJ8JjKUCjDVX32NOmVWrw4K
eZ13hXbZDaGoCt4qwb1hgpT0jN74c+QAEFkQKcdEfsO3kPVjAsDJ/xX4eOGY/Ch3
rtBqdZve9AAZWGaqEOQwatbfo2RT7O79lpePexJQ4ozRRF9SSUHpIJbhyBBSi8Q2
f5ozsBd1dCJE/X2YTAZbH1e7DlzSGZe9E8yPvlzXMF2C7yz2X2irw2jwsFs3sjiG
8371yMb5IIjZjyhNfEz3AdfTxEgXo0JGDuXI9l4napAxjGtY0uBxyRP/GFj+ajsK
boO3Mc1YDPBwsOvPTjOK75yUkaSb3aNgR8EembjwxJXSKuu6HnOTKQy4uTlX4Tqa
eEZ2jvqXIYI3XaE5hfOdrvou6AIC2eFq4746nwA0DNJFtVnO0hzDBLS19eo7XLvA
1lUsVO0ZluQgKOcVS+tekOpHPygdbi9EnQhi+zzJbVa72geQlkMUtV9EEvFrHLB9
SRd5J3C3AqPlNRLxUczKGySJn8HucM/V1ZWVaPgGMwMHNEb4FdPhymJRrZQclwRa
c6MZLmiQfdGZhQaYzHXtbJtEIkL78qlRlijSJ4xE98VSTLiKkMfXEw+lADYRgo2b
yQF5zjC5+N1+tpvDQwl5fm9F8OpHMfaYIDijCqrhvWV2xM5ddxz1o3+EdBQPInw+
tzkiSNYb8kbZBlUrf7ouquQY3xC8Hl+OBwSzLCRDiT3Suv2s59inBDZvkdlFy+TT
4BvXxucwVJLKITwoxR9mJBvwsTlJwFsd/vx3IzlcqcoJOz1s9ZiAgBntNZ3SxULJ
Q2D63LGqAZuiFZ0fdFLzi1MrEL7BT1c7Vi82Svtl1Q7me3/vpjdjvEi9NtMlz440
5E03CVqN4WvmiZTsjQ7MWFP3VzU+JHPWTsS/7BRoD8dbelwIfy/0A28MS1yHVKZ/
3NCu1MjnJdarCX0sTTIjPQARpqFpXEHCmasWaCanp++t7BcRO2isrk3O8TNq3Vok
9DJnOC4re0nfCjAIGAUD035LVqUa7SL/CJ/NUgLk4hDtM96H67+au9tr5dSslxX9
gjKk0iixqSp0E+XKgoZJBqQ3X32QKgrqa8D+OcjQaTDQN0+jhhWw+0lcP30HqH8F
T2izLoq+Vj5s0xoKIO16w+IMxYJ5oxizxpCTYLPkk5/qh2kRvFxjN8ftbFIfm2Qp
9SQLZivBTvI47Z/Qe1vPS1i2+bWhNoiEdnVcmvhyjHYYiWjN8NGA+sRcHpVfcjOG
gRqWAhs84EsvkLq0xes+f5NBFvJaoMKZlm8KHH6ivf7d/5CiGCZQ1yc0AJU7ZyXZ
IwvmYy7icYLqTKozA5M2tH7+PfkBxt9K1bwCVsh7lTlavuJcrpS/VCOJsLur+1m7
b47QYxyzrXR7aDnd2fAUVebmD+KSnoeSiL7+/lRDwvLsO4TpfzXYaXuPXaaRCb/6
9UZDcCLrYI+xGzLiYUksjeEaQ3jrDG4q5qAoEIa9xKVmkvGBseZjCsslOU5jvE0B
bCWUWlAkINHf0t04Y6MTTVcJXNJiTqqZziqM/Wm2qiOExnCCk3ERVGB1a0tSSyGV
Hz8IasK33cI32blLRy4nxutzW/VNkEld+4qo66aqOUAy7tjLlFjk5zGSthQBEXXj
QzFhcjZBzHzMrvxVPGMHrc4+hXDCJIXuEphygMQbQ+6JEjIjZHnhosYIhpaiQKlb
R7rk0nPvzyQ4WKHP8B5h3kI4shR6Uek4ntSHbnQk+77/sQdcmLZhE6FZeG3q0xqR
Koq8NFbDCJ+QzJ3iuab5N+Au95yMrMWoNtWkNtl1aOACaSNALi5WEtcc8/1M8jwx
i4MexCBCxMA8Y43rpefsrYA0WKJYrEAlmMrxDQF5dnDgwhKWJ9LLBTCUboyLUrCR
hTP1fBLy1LJqNM99375sOqfgbdcyHMnm0PiUQg1ncgzIs8d/0l8SDwjPQ+9phKxQ
vvVLPMYW3i2LWBhde+9eKK/eX8B0iQ+Zn/mitnFmyTjDKnaf2O+OyxaX90/D0yhg
GN2MfnsrFJdd8sx4AgWuw1FFTKNi9oyWuqyEHI7gLY+po6unCZXke0EyzZYeOBAB
x8MY4dFV5FvoXQQgt0aK9cW2N0O8jmJ2ejJh4mqL5gDWzMPxc312/LuJ2yHZ6sSW
3CzZPyapMeGnxiLM6tUUTbfWrMF8NdTRB+Aozue2XK+Cz9qscTmb++CZ9czBwtDV
pRNjc+eWiCJ+Homc5UMlZhB3kEjsijix2EbnRk4gp/Pu5EXjrDwF6xk4l7Aals31
2/rILd8csxYW2+GLWfokNN1ssUDzTPiH5q1SJRZWyQEt0kHZEyFjSeyT6KEZ0u1A
x1bsHPj3qqFD9qm4J8k0QI7MISj5rqcy8n6w8TiFOHUsW7T//bwCu34lHJm7WCtn
KYOKGvuI/VLZVxlSGYaYv0V8jfWNslRzOrpyxwimd5NL02BdMt/EBjO2oPFyWrgF
hOb09vpw5J1/lnquSDBFjYbJxT2vxgbOqjQ766B+IiypuwEf8jjlYJJ/t4qlUvio
dc6dOnFyZVKRhRu+FXzX1WqnA1VU9DKUF0ZKnbDtMGj3i8PE2ZGSJdaH6Lzpwpp0
/GVBytgFgpHC5ZyKa5S8ovw303rUOu+eofK+m00DHgGI16DfPqwXELSI7osU5b9Z
r2x+y7Nje8hKetvmlXllECONibqK9B48OG7xZEh6c8MYW5x7/otr7HUPv85ogkEo
eloDhdL46sOoQJqfM8ScxyVKYsEq2PIEpjeFoL6IpyTHu9SXFXVzlIpEtzLLTvh6
35PgBIkU0OZrsIFAMvbAmjtPGct2fgzBPeGEfkF9jKUXTIpSKqifAwRQIKyNIDAN
mlVgNg1tS2/sLq2S7ufzpvg6zZ175MCWY3eJoxroUMgXmcEA6pNlQvBMFnPikg3F
hE2SFZBzrGDMgh2zoJWrXlWucA1/mlE430E0dXZkrDemXQcjcxq3rEC0/6+21yyH
1XaKWrWqOvn0enwRlxeh4whbg04bt64PMA6JH5cLQJMPAQoSAZzIJC+huAt28A6c
uZOcqh0I0A4BMOTNEoi1dKCy/YVvVNPmHOBOlVvdbZrl4KADQ8KyXSZml5NLFc9V
WQbt+qNXVzn7G/KEY/vmvXT7YktzBd4gJZ768/7dq69qDbVw57C2CA7WD7iW6TjU
vUWjeqbJTSXi/6LamnezqRKMbW5/pQ9LZcRsRQYw53eie2HpPAt6eigh5KzKCkFk
/OLI2VP4Lch13CETVTQrts4aEgZqnqm4FFT8LCcE2hUK3YkkwXdd2kiE6Lgq/3/q
jfhlUJO0FBC4/M58XcbHWlHveUt1E+Qp4mToANWntKAajI+O4tFETnqUjEa5UYwv
BUsRM0lzNMZWd8lf9hWQaGEAk2YqYCtggbko2eWr+ZS1H21cYwmFEycLT2wFw5Lh
BdqHdxLXNAQAoJE6LNa/BfZnxPRGqt2GSzpqB/TGP8ARnlFyLJL3DX1qz0uwYEb6
PqZPnrg9BLcUbylXGdJHe5rp8311tKZafGhBCTACkgyOkhe5GQYY/x/QNe35QYUM
ea3IUO++2lbN5P1huMhoKRHszeQ8DJwGMrV6d+NRHXenUZiytWEXPF/xZ7V5KctN
xFc0SYtAo6/jT6sEcrBzz92BuchyspEpOF1nZV8M/LrLF35GovSBE4x42vOm/x+q
eGB/yoCpZlwwRjpE7nOdZwl17sxuO/qAYA60nojJpqDXUY34L+v8YxCORyrU05u5
n2WKfYEH2u0vdNXH9jgAC9NKS1GUOIu0ypYdFkgNDo6n32gedEBkUV95Fgj3LJQx
y3HdASpz+Cc12Sum8U/iy7wQ1tudNqjbjB0uRWui0tvqeOlMTh/KJpMwiKB7z+39
3BL4ZiORPZp8t9EnWeHD3k/W87U2iPeelkDqwgdNDmBHJ2b1jht73qzJHWM0YHdQ
4f7MhKFjN1Uwyjc2s/kLr/oHj2mllRniVgisCE256sitv59IC92QuEqWJovRok5K
JNwbqxEqSr36DI3znV1e0ocYMFzginJlwgVE5Yr8+eYUOKVc/8p0NDbktdNJZUtH
ih/RpJLNWMXAjYwpRYonKyWbscvJ2LgDqqbbkhNva10A70Uc3IEoPHRWQlAevBip
eOMvu9pesq1GutCnTFRtRLgkFfDsRl8/7Bt1+MnM54MZPbwph8KlPpHzats6EOXW
eNSg/rZCvzXV9aWXQXa9podURtqSKvZks05Z8ZY+bxnt5zQM8tE19gOI1Lpk2P7R
GHRadvFojjN7BnJ2i15d6Znk8Djkfw7nQ3SVT2gczSTSV8Ho47Ok2KCMxvDwIA6l
N+O4UeKfA1yvsKYrirgCRffjo+QPNv10uFhcfUH1hAZACuU//fRDHTnOZ3S1z7O5
KVeU4N69fLEj6nnaS/DtznncmF8vv88tjZfD84znFzzbkRD6cibbtIhqUMH7Pfr9
MRT3IlfTQOfmHXGLtkJvHVIRXHmvWcOt+ZWCQVPbnx7Fj9fYnGueVKOpvsgs6wGr
u90teNSlpkYFNNPECOasfJtjbMtPfxt9cr7hl8kfqygbHP3Qtzb6U/OzqsicwK3t
Pty20kf4psnJqc6RJ95hqDeV0PQL5TR4J4/Njvzixh2bXf8mjVmQsw0UmK5pVbep
uZAX+KqX7xCigQKfe9Z9CuCCyHC36ZJJBS80fBz1grZ4RjAYslgjws+tK+glf1xF
i/n2b9/CwXqlsstBfFGoKAD5h8cX8U1kqpxuzie4VPk8I/JxhdGCtfA2DiOfGIpD
zdn6wT2lXxkvUH9vbeQSpnP/ZJclmHHzhdjScDNluFCUW2Sii3Xne1/Wfur8H0Hh
KLyCM+dTEYXCJZ4jhNrv3Dm+fe0RKfkKNU3eHZqBOVkw+sbZXaN4msw3lw1ze4OW
wUEzE2LGYK3Hco8FrBa/qi2Rk8U14SxmD41r1JdG0QQRmPZEJhiD6Xt5MMXwNwmL
C6/r/pFS9dThlKUCQjVerWaARLj8ze1uogo1Wg1dFupW380POafpe9TetGjMFEqE
HHSaJtVz+z7dlSPuSnoPpdaf0TBjz7SdkVfu2hZOD3+U9p+8JJTBZe/lLrm+RwSm
j3GqTUUdDQFl6KY8BizTqQXrE++8eQBTwa6RdCLPc3iX0vldljO1Iw61+dUZSCBH
y+kuPV08bo6c473486mhrvdE2IF5RzF2No8DNxs0Tv0TZvCUB5rLa1p2xuZOtd1V
3bJheAFClR4ogl9tq7IAI4X+DhtQojrHcGb4yi4ZnMkhtAJkynbQf3dIiSbQIgpW
9j4RsdA4S2hmpb9Ki2eRUuA/dFlIemWZpEChVQ+TqLsppbaki7yd+UjV9RHTaclT
CXKWglQKSP+zOXciL+Fc7dYlCucoRJIg3N1Gc4VmIlyfyc4p76Z7n62dccZiUsy8
CLykK7YZLapbXBeLYge95GmkVmfFSPOLAkuiaYlZMhhnhFrpv7Ga32SAMyP5rWx6
RBlzK7iAyC1uSesGVMp4cUlFkKVDzlvRgPSJQVMi6D1rwNVJCgQnrXYpEMpyKKH4
djlK6oIDC5bqqpuc7Ee8nc09sfdwi0aazcI3zMOen4ZlQXedWzrr1YgXAWqkz9H9
REx9TUdWDSk4y2uqzmCoX8Z5Q3L8vRPEzySOdqICAGe3M6alHww48kNN5IwyygS7
rFsY3sDPJe50MYy63ByHhiRbQsdJElCX8CpdPn5USKuUZv83uTj8+kk1Dy7Bbasm
s5lmnVji4m/HjAGfu2H5IZdCxeAn73M7fWoVLQ/CuLqHDkK7w9ExHJiLAQuo2rv9
WaIFdiTbkEhE37VHkVvbCTGNs1sZFw9QHzwUUlxMmAv3DptvtoXoL/0FgKFEN5wz
74K0nzgxdA3waT9kr5c74wZ/GCOALI6lxHHUK139RjHqO8jp4fyZFg0egjzGPhdi
CKVJqCFUZ9PxKRUkGidcziW4LQcHERV7yznc2GUapXv1/hX3W746JbyKpnwspjGj
VYCXiKR7Q/H7mikYoQotj1onP0Jfv3cXMPMoFJXOvDi3YzZUbSZ98F2lUKgi0pQu
yci8t7egdyi8CAM/0Ta3Cqd/RbIL2W1wZEyWqjF5tXYdLD2KHaB2lPPo14vlyrkp
XZW4x59LY6Ndm0Vn30RhEaIobg/AZJnPFtZ0F3mYTxEoXSCCGriggAMSCpxmMb/b
qDx1/wPS98ta+1xC9pP2DjaC/9p/zL8cH2Opiu14HXYMMD39w04mjViYcjjANXPQ
DeDkS3WtUjY5qyA8CM5rsF1vwIBdzVnWEm3rnlCmyGklKkFMqWqTwFQd6YD5VatA
ZC0zv3Umzk9UiLfDhLpkNSH7eDgF7Ca4jPq432hWqoaNSRJbDfTA5R4vc9/osJvI
iGHHmRU2wCPwDm75+Id8FvcxPXM8vp+U7Q+V7waf1LP94TJTIN0Kcez2uZ+uds6n
zpzZinbuzbQCDl2Eh0SIGEgJ9MWPJWJsKUVgqW0UDSoZsDWR8s1FSqUXYjkbl4Y3
rKuWiQ2UfEeDoq3sa8Mo6XBBloQwsxWDT7FqR0JtyJ+UwOSYMSuNOgZoHAa4Ui3v
Fzlt/HaFj53+vNJu0++XRIM59V3SZrQrQIH5Z2sOXE/yQkr3O6uBl+MRFIp/FW5v
rcL+k1Y/QdGeft2BDqn8M/BnOnxEIG4qwhj9Ntjp7Gb6xzQjvIJ80GUqFxr/x6pi
Pe5iDK8I7InBNaRlfr8i/BDYHsQ63PSu/gVBPPY/TvTw4C7zjz6dIOQFh6aGWDth
19nQGWv1Wojp39MuR2GT+sDzNkaDPedQ0yM14N/vEIsv6I3zW0vNaxKbGvg1N8dg
vUpiBP9ssD2ph013f2bbWvpOxxuaGrc7I7r+Tyyc1bssBHtLUSn8d76iM+fv5qe1
o81d9DRbSwElizEnkc+kw96dIxJIJmJCqWf/4LZiBTdPssVbeZDFQL3EtSoAaYjH
rV3OUiv5jcnJ9ppPkljpdItY1lA0IZT1BEwpdHgxkCgQ8kvS5xFLGiEagoYkQT+0
6OubSII1E1WyVueHPmntm+Ihm0jgNo6iC9xnLkppJN9HoriV5wjTkJVV6lMLqEyY
VsJGd70t1D00dac4PlAaz3TyvNLPkCFNKMC3cmrspwnc6ssOSBte/dOAtFevyw3f
uhmRH9qDhbbmtadQki2Q8/tcwRXBnS3HJXE6rEJDAoUvZ3vwnEPkum4sClj8/moL
lNKoHGlpMGiuHXDvg61Z7bPKGKPLScmsFg9NIdSspvE7T+MlYB7wDOUb1aJYH4fd
rlc/6BxtV2DXMi7UWoeyB7vZ0z2c4qRbuNpWAkDP+TSWM4EH7qua9Eazpo1Pepma
Fbk5iySZx2v1Nca+LaQ4BnrvdIPhG21UwsklJUrO3xgJ0gnHadW3OmR5BbZYULtW
5MzZ5krwSt8+D6rv2aJ9e1rfHoWtBYievcGrqR/N7OBiKfXCFYniVa29ITpw6iZv
5ezS/vI+rruwV2dbwSa8DemIkuRZOtbNNWCXfxi1cz8/dHybsWKSjNAocI+l7pJH
NSbafbnlj0fz60QCWCmHkKLC4YeSJS2efAv3kh0QlXJggJV3btJlKNQOdZEXCb2V
GWqim+gfPZSkQL0aI7T/id8epXAltd6g8OJIgsAFEDMRo/QZt2w4sIOSteSximUq
KBVrMFuPnUG2KMeTh3DO9hLSJUGuPiOzDTGsypH0iNQADFvxtPeNRfDXZg+ERVfz
Lcr6ed2gyMsFQ02eNlvGxWWi1SjjmWGF1JK1TqRzI9COpJiLgq1IBPQyjACyrRGF
BH+PNu9XVT4dpg28xDIcEvJEcw3xy4JgAmQCq6cAwli4m36jnSmJRBIDkQhjZxMY
dyzcnJyzG+YFrJcbRm2fJVzU1/uFHOaNUkKY+9GSXsOstCFAfU64RF8yD1xg/vmn
Gftx2Xg7RcZw+G1d/HaoLJi0cWNS6YcKcLYVGxiyEiatVUwHQLTqO4v2lhd4GxTq
sai7DDHE3bICbERCmeKZ/cyQ2mtp8Xe4Wasm1U3lH3y1biK89F9nO5utOjdzEuCY
QnPcpfKk0gLDPFoU25sDEP+hGMSqdBtuOGmhaQCiMyBwKYa5N92cDIAmTIPBsVKa
AQPFW8jkt/2rUpTloSwgN11T3uMv36IOmRg6zhUNQFEg+WhcF55mHj89SW2MzbOJ
c2A7QrPVBDsNe/ZYe64HLL0m5s8BuFV3A6twsIxmE7ZFAmGEqRakzruPUdgtfzQY
pgID3NcGunK0Tm3p5v8jn4G6RoWxdD9H5wLu5rkQuM7Vr6k36sSwrGwl+RMiStfb
+Qx/ivGSVgDiHqcpgmYyFiZD7YqDD8SiI6SkX7D+4JiNojZjZEGvZepv6J/jOOdB
zHXEaKBLiTUPGczjuPOWe2/kojPymAlK5TogbrURCB6n/23WZ8sjFyjSHV8v1p0D
IKyeriENKiD5JgyPWqs2qOcuoKg+4slgqgS53fVdfVkTCcTNPyncL5FhzDIOUhCn
iUmmxji1jDMdUo13wghUbw2VCCnD6o+5h8p+1tIoQAZWalD6NiRd/AZLQUBVhlM1
hhrR9OGecO0fMIlzsHHglPpZ+FzZ2PHxth/Cg0fn9TSBuNGQhFRBxl0D4FyJYqPs
K3AzcTKk/dX+m61tyR7iXztIN3MNQAfIvvC5RJ/kOWKZLQn3V51XyBHH59+aH4iO
nKB7p5l3ER03D+510IQ8Nj8jSNnUR9u3sRPH/+fdcmyJSzCqMtqlhZxXoo/Avbn0
hgej6hF9/0UzVE7x2dEqci/NTxPMZwWqqBPe9bZRJSfDOBhpa7Ipg/9au5xj8ARa
rEw0PtqXopQIfx4s8tlnW5PNebI9vdtfCtLJW/uS/vx+rm535HquzpLGhb6klW8F
zTwK03/pcUksoxM4SqIQu3ogkCRztRCz6GmLLv3+KnrS0NMdfL3zRZ7oXLfVJwFa
X7ftSgseKJemLT/VIk5fJYxNfEQoueTQhhgd8UyV5B0wAAJmAew3Bm+meK8jMLNb
kK3oP+cjh+0oWY3mLz8ZT02qdFSjF3rvzaLWhaqgJfDwxNa93Yx0Ph7jkTedlYA1
/H4DnNnGVE8H/iTjrcENNlqjYVsYDMON1mzc7sknLm0k0pi2FrdZXqPkmFiToPo2
ceKBRzzcQeK6R0uG9nxeDCLA/vQQGDxtxovV/L7xLiHJYEUqcP68tQOeQa99Q+XX
Hoag2mU4jJFW47y0PMt94FK/ZMDnMqClYt36D41D7LG7r83R/bY0obKaieFEUDNT
I+YYAwwgvBvaGl5H3VzmKJ/Z/qPzVVu3rLWL6YBU+SH0wSdDx1io3TaE55wRKvi2
Y+nG3FTZpBsVuoFRh4PldQ6zVb9raMlwNl7I3KQbZOCD1e0Qm57XCeiGDVGb3oPN
3ICFTEev20d/E3qN6TPd/MLzcbjkm8wvVtGIj9LeZU2bx3A9y5K/0bnY1CAdaLje
ZSForkekZi4no33NUP6b2Oehte5LCtRsRiw0WrAzCdbpwPJU9cPKZyezI3SMWgNI
fR6gWgrzr/6v9BUjqmgVPdMuU8XtIt7uzuFnC6ldl4jrzDxnMZ8AgPFLQM1m+axm
oQlUnjSsrr1EZk/2p6ABtdHzY7p9FVRDOsxcahxL+cNTef58iC9slO6lrDnfMhlB
5JryGI5/Xzs5KrxVVCVOA6ZT71O2U0muOwzSKvXddkeaqsvEMqAD6SMkkiSGcxkC
C8NUvRQ6f81oMXkMthIOsSKYGOjz6bJigKSmUrcBRLnBz3UR5n5bgmSmHL+AksU6
w8jpwmihOYwe+Fc+p2GQEhzTfnBogxccoVWGgB3ETDFK0KzTs0F5MkXKcl/pCcUL
sYKZshi726IIbgBvTep5kVKN+x056o+941jFxaeZKZJjGqW48Gy7O28JSr5JOVKR
Z8cBk0z98+jn3mPbvbO3z6U32+ed+E/EW1jMWCdZG/NZNga61l5PMteDJij/3mQu
9mYyiRsmAcC+ENnaUOYpngEqH/v9ii1geuvGDIJCveE+M+2qzMsCmypgY/AmHPub
Y+kT2qGQyBD6DJ7O1HFaVX5VqDZN+xTd80qup4julvXLg23xnphH19ezGhsoOTYb
y9SGvWAEobvDL4rSDN1m/LoOHmGJal9bTb59Du5EsQkwhnpAL+Ii/7Q91j6s1Yq/
51ffPS6INfJdmtZ4Bz8nNd0XfNsSQHHbFYxyKiSSy8dvyRtp7G32OIbSSFE+cI8/
Io+kZW6TkyUaZ7Loyr8ntxsga4Lhnr5rLbiO0c6cvGtQuLa2QFksfNgBakH7zdtU
aVWV4K9GJA5J3pByldH7n2KoY64CEp2beB5byJpMaGpMWEzdcKvGALLh50ksBH1M
Up7h7kbwg+kaFlEiGv9TxjneW3aqK2EukZCGuEaiFJ/f0GboTmLzFM9kfjo3KosQ
IXOcYwJoYmKHRx8KphVeTwz/IfGV4Hp3OJDovvDihiDc85n/W1v7RKbHJuwyTqn1
Gv5jWS7msDZxEHqwH5lmpG2uroc31PYuTKgMCsa7hYRVPNzbpCBA4dtXY7eZ8w31
A6p4KYrU6p3kDk9eoMRNeYI6ythR6oW0Wu82XLpDqvctUbO79wE8jd8+oqfUfKNr
01bwLk1+aE1doenLZc0qOGVFavg4nJgR2CA9s2+emIHOiVO7FS3K883ikW2Ijk6u
7QRc2BDIMNl6dq2J0cfiOtqVYmUjJWEEpLtWeoUlo3lRNseiinbU7AroiXK4e65g
qXVeUptKyPBKB9Gelu4bVpwB3uNlbsISJ+SvSLJBNtmCTnyeVhG3JknPEsgr2Eg3
ditapE43vFoSzf6pAfAjdW4khcjjznc9XoD+NOt6V8itv7mqfNOayl+fMffTXg9X
vSKMsuIw1vC5MBQ7HD5sNXMMWp/FO04/ZdT1BD6ks9Uz5U2+fmi16HvdW/NoIDK5
oPdLAoUAu+ZzNYMPcLOdAPwvsdXFsy0eLcVvUyQne5t/31/w1xElvUD2X4RlAN07
FRlZUmmidH/2QsXszib8rdiNn90isSBLcCmytHkdNlkidEZBWaS0zvunlaMVNe/N
zmSzKTJF5NSgx1HUrQuN5+xYP5982F/w2jiPbsZO3+VMFjdHmwTy2AE2BdJ34ffq
Bkcw0/IXzoleubsD/jOTRKtI3TSyhov0DD3eNm782B3WNEe/sJ+GBZGuy/bWmAM7
ZnCN1t4UPegUTxHoELL914LO1NiNqZttORt4jdrWDWlqkdAtNF4Xpq2OWFAS+L3i
OJUS+7mKHXF7pTSOS8oHCiICOBuaR+eeu5jhdeSFpQOAK563UQzeB3jwmNysbPwV
Y7HobJokIEzsxU7EHjwG2RnV7P/yt4wVM8QwGZm1U85RLAhaBNTKWOpd+qshxjRj
ufXPqJ3oPVTChJdUl3cIBCSdbDsoJW+m/pjuWzTlU85NKpbsf92UnZpT+2MXFvyf
IdI7/Pojzjm7yBbjBpT+mPjCghUt6VdyZ61YaYEDxjYjcxoUTxrTcy428eyO+w4M
hTdSQ3CWohAGt7H/pNgG16QwR3brBu+9APJqdJqJkDX4M9t/s3Uaf9gfEBm8I+Mk
WU1gR7eJFAl3Y523L5bh2qDJymSLikUWRMQHSChANwtOflfjEU/oNyi2WcPARcWc
wsAzae8S7HpQwSRkpjvitX5LiBCeQgVwE63WKhL8dRENi2Z7EWwjyX/dP+nXEkGw
v2tXWFcCdAWsNqaNFCtJGjIm+QQC5T8Uweg4aHatZKzeFftDFZqNrvcX4j6Gq8Ph
wJ7s0i7I26cbBaXWzcFoV+dI7zwehYqgxIHBoMhJdLSmi2zxtiFmNYPw+gj9ZQ90
bC1um4QPKS/fd1vXjl+C9UPIjiWx369pV+JgZAS5LqoMOicnQtGyZjMSyzdYoIaX
lbsdEoYgEGAVE+Vu5Tv8vuuB4SS5wUO0GJzJti5crIIZEovHLichv9j4awdEbrN3
zU4T67CwnkBFon4RJYQcf91DbwZ7KiyyLSAEgGlPagci+OykkilDliFluWcVznFf
AOxX9jx8NTu6GesUy9R9mWtcndLtYgtEQS29Es9sHIVmalYstto3dbsuWAL8dIxX
s0KCzcOGxqwkz6Rdc5BTM3mXDBfSmhHLoY+i+kW2f1zFRJb6MhbzLGRESxVgbRVK
hjei0Uo+x22/WeEZxAfz5mbYxrDxVC8t9wJteqQLklsbv9fzyv01xqoMrj2Z2hHL
C6dXMUhZgBM0dfli1wS2p/GISLHc7Zf6bdo7Mug8W5N8PlnhkpzYGm+x7sj/yasS
YkEBbBlVPvlYm2nlr8mUEqnA1rw5W8ySTAfFwSzy4XtyWwNnsU2uJn7Hsn28Swki
XzsC8Nk6WbqX0jAVLmv99HK7O3pPeZmqJQ2ErCL/99h1MpqnyWmGoRMGSnxiv6O/
mrQ1aCjt5R2YPpoT3eGVSjwYkBSa99qWBY0CQNWOhttUKuzSEAEMs6NLe0djEp/p
Jba4dUSvLMxgmbLj0HepWLm6rdjt+CwM/Xe2CgD5Wk1ZPfzHM+6jOG8Z3TjxCMBY
A44GZdgcI41dKzJjzUNjEEZULE9C6CQIAHM8uzFxccsh/Uq4AmjnmQWQ+7AwApO3
mvZ7gV3eozwr6U6kgKwgHOi6VX6Ah6iCOfdR8xNMjz4zjMTfG6d3QEtJPXZUJHGZ
w21Yb5CFpZwf8Bt1o070gOKMloR9urF+Pi7LkwcAWxIT/lTsqa7pRwSJX9iIGVOE
gJNNRO7yu41y1miPPVsZF4hnD2fzvRwN4phUzHlp2+3M3iL2Tz1WmjXI2157BMMp
+DnaNM2EmKDXQ/5S7TPEkDF50O3hD60x4bi9YliJ9UObCg6JWaj72E+d0byy/xJU
TILgXfr9IEttvcQJg102DZ6HCdPrr46zvW0k6ldjXxcFJcCctjV1V63LpinSYv2B
Q8FRcH8vdMt+iYqJLEigrkBewuTq0ZIVtEo/id9jeeTkR5XBu95G9PjSfMMDNQlT
5Wxb5GJILJtVaXYLHJH1fJdC0d7poUvJS6u3DrVRHlYj6f3euIFvggvYCfigIiDn
cOg9Ac0L+k764gCDYCwXc+tbM6e4PpA2BT3bo8Jgwn3dzsMbjuYviyrgOuIFtFgf
HcAvUfHFtM93jkz+jyCX7rNoPJbUw0AKOMD56q0tSuMR+Z7DnYNbuJ8cQwUFxbXx
T96k5nnkoVUb61h9KN6f+h32ifS7D9fIcqFaiJIeCVSfeYfaAUNalgeMjpxkKy9D
GBuMMURYLA6nUndMNuplUu+ztlh+Ap1QJeExGF5nAfvLbL9bfnSL9DisLzlOdzq3
661zklTAYlTwyhQl0F1vNrI5ocrDemnP5rsV25H76B16gQojyDPHGR7p6idPVyk8
wIs/ttt6uoiZlb/6yz40jLqnAwWmKfe+QhL5kLarIKqCU/5rs6OasNhh8gp4mMz7
Dgr9OjN4p/UmLorIQnMPzoQ8heLMXaGd+GNtgHaFqmFgObEIFab6G3Eyafaobcqx
BpMYr7TI8W3DMnQ5DzZi6nYDwybq0AOrXYIWwt9Rjp7u119+zd4jXr0RRZbDS9OE
w5zoR9npYR6IS64af8Ua1DgY8iya13O3fVbb/eL/FVbkisCQCQ46iMxLO5qojNxN
+N1xPaPd7wQOtXOyKa/1TkazDh6FpqsDoF7PRztB8XnQd9cztxa8t/ujUzGyrOdz
Jquy/7uV8pqw0tFX2ACXACsW6txniX/q3e+ZXqivN7opivjfD0g+0bAa7zfRe0W2
SwsBUjVE+z836tnS+AX3eEhqXWh2C6rh2Mon96YqJwNeyC+MBPSQUkSIypLcUmzw
YBmLb2AurZFY4cFTp/GZ0OGJ4E7oMq8UN5qpsDeo/tfibfLNrk5X5A7nfE5WLSun
MttOpIdNpXx9TpmJmXGCari+Fjx7zHJvxgR0Nj0S6xfsAt00q76f4ceVlfNawl/4
EcWKWMI9dQxS6jM6CK0Tkanz8KUGDk1hJQ0XsEBhmhCa1UtBo0k7YTfWk0+Tx3g3
AkiFmAL5k4tk+1WVEDK7hrbV4KWEi4gVkoFjlq8GjKvDT2nIc7vAlP6dqcpUU3Qf
4ePI1CpYUoPiK8Tgn2ckKoSzcJFHOt/VdJM7FrY84NYztYVpsj26JuBVkFIOcHyS
eZF8ZFVJmVzTR4M1AC1k52CeUuNDYOuSaebfcWw624vwmurLcnp7/R1jbT4y6Jg2
FViotOxJDjnfYE8YdXnUPZrwtAg9zya+6bb+SmJvdcgyRASySzWr4PYMW/WWyk81
h+tZj501TM1s4SjRsnlqkQeDrscNgOFu4nZVuo1M3GRmJMBFLRIo6mYN/8BF00MB
3yDhAV1Fx6jxuDq9WysZB3rPO7gfnACSi8+Px3KMnr83Viq3AOs81rKQRioGfZX4
utaa9IMHYXIrqpuxjgD46OemcYUnSA8p9X38y7mBqhk1uO/bHcGOXgegVkce/9Qm
tSPWzyobXoHs4McdGBfitjAr0Gu7GaH3/uLMK4PA3bR+dA0bex3gXprDW6zMgYKA
kwd8ap4ePQJjkpi5jyJdp29JlAJexOu2/GXh5uJWIgfdz3Si1PRer7YMSjUmiec+
8nkH2kqDBZeS4aWMYJYqVSQMxHW3tOgh5IwIMnzYxZzcWfIXMDhysRLrHkAhsOFO
hVan+l7jRVz/wuAs58tMS+7o/piEXC+ofePIlgp1hlkMCW8/ywJ6Rlx4iXCDKvl1
r8tsBTv17qVfef8bA7BzWCb8s03dpeF6BFHUUeKiyvvgtjagAlLTkvtIKdfGcyo/
D3Fc/UjGspYlkoNhJuEUXlwwPjUSncgEGET0bGAj3jGdRLWhoCXPVnq98wwsAiAg
dMFa/astZHdTdm3TotCvtrlHpa2CWMl+m6LeIreo9gFrD0qgag3Ybcuw9P0ffKib
Sp/dZ/HjZl7tsDp32Ws07dSmh925Cj68HcqMAw6LDAiESELuVufTwyRUW4bPKxSz
rFFEcER+p/PPv7sRx6qOh9pohHnQFz51+CSBtN+x/Sg6QCNqLsPBFiXeAzPX7iPP
e58ZMfsZiJKSZZPY8C67UVmTF0dazk8bGxSAvTBada7iF6spsYYJ9CTQGDGbCm5N
JFzNF3aqAB73SJoOBtimYLKJZsVHa4zvx699dh2T7HalGU3bfuBdSJEbzOEs6e1c
GrSvWFK0pRsoDHxqEknH5o23r9AVyzIeGG8STtW41KyRWV2HnZy2qXWn9eysawUm
+Okp93diIUjuFhiqFL1mHyHn4uMF/UgStbilhl5TAc8RqYStRDkV5p2vKuXrKKnY
hk64yb6jY3fgSH+y/ipQDx9UHYIhDlTYRrKd61DhH6BvRfkUASUN3DMbLlq4Ubd9
/G78R9Yc9br2+mAEzRbMGc0hJ3YsxF92+UcugK3/7zoioQZdkUA5pCgbfdVJrwCs
RmpxcNsDlljFzNjDFo7sEFdNuvL5UszBMewLdZFX0I7tcPCeC1YnK/DRHLKMoRat
p/nqrQewfS4hRgTNiwfH4l1mE0smDeb4FQBrEPqdhMBYI0Q/uQ7wzbjZ8KVVsZn3
kRC7jGLUbCMPnrBWH3nJoC+5fo6DTcj28DA2eBg7i6vG0pshPaboV3Kktwowf0x8
yF0xOz+JUtw7FILw7SW84WaaDQUkFYlKdPyCsYu0kxeyjkFD4JM5/RwVVwVMuGyf
n8HfnpPd6+QIvL04uR35hnsReuH7QakIysa3VV4F1IEGDr3mOorYj2IUJLF7gRtq
bPeu7f3wboXA5pp1Dj0+aIvUjqEG/Kw1MOqqY6EQAF7+xY3neZOIWZHoIPFu/JjH
qWU59xBf+CIaLhJEOKIoIpjhd5+3T9vQg09o+/mrTKaU9boPQ5G2ARnO6j+0GR+J
EEn0wAV5bJ3yboFpfHVE6aa+vF91QjKS7+kVk/iXw51n0wbqYvvHg70lRP6kdsgp
gnhxj5xjTIrLwa3enhHqFuNa0kTO5O9aiofh3fUww2rKfGs3y4QpgH2EaIntEmBd
xevmrLoGif/iiKM1vAVA6Q9H9JfVeEEtIdFKsycwOzsMWyNrmavhLmW/zrdAAqr9
EG7wvN6CoIte8qNfWiCuyJac2To2C3yvE0oAlnNloES85QWbSJyCUl57pe/eAJNJ
nlOvB4ceiFeJlaEVaxCTsSAZVcy8V3xpUsc8HWigHA2NKGuxJjBqoTz30KSmh4Pm
hRPIDlTf6zxS9IvrCvmqWYRAAmgP71xX7W/dE91528RAcWv2MtOOyoWNGKVbetbe
69mASg8NBQWcEzuqp6DwawjC75DW/2h+Vojf8dqfcaJLMoOEQJZCYFXYyUSwYio1
zDAMNsxN+7V62z+agyUisZ6nLwHkfAFkPFmO8+8YYNoaoAtfVihY+EOc/D4DGV/O
HsaJ1afqIawQ09Dzo8FpVT1ycJ+e8EiAIYCt+jw7uAmzfq7AOj2nigwXiU79v8yC
xVL8rlcJoy+NU+JCsqlrhmiZYU7OKvj7bsAJ7azH3iN4bE3haR3QypoWJGSKDGx/
z3b+e7+ZPKN3Ewa41/uo83p0XvzIwwW+JD2HkVFruWWVEBLqj8EL4teu08NDaSYW
6UKbHQZPa6kP3kDApVmlrumM3fxUm4160D3ZGp/dfDreE+/NYK3qb9cROFlUwj20
VJzNKu6MCNXOzNTVlz7CzCI9pQ4s+1HVhSiaQfisetEbILAebtXH2wNC4niVK3Qa
g14uxTJewhtYAjEcc7sRIKVpCkNvA9KQda0vdOsGVg1p9CirS2wDS4MKWUiZrN7j
WLcsNL+PupEYjHe2ONCwTe3oKzmBVQkaWNLZEDll+iOn6AcKnC3PH2zZAuDUVpje
WLjSxO1P3zSq//dqvoZMck0B/klNplNo8Fn/vP9pUq1m5++UK+orIn14ndjW9lHJ
8HDns7bS9GbtBI5wmnLWPNtCLF4L3uzzt/MFZGGWvB9Dk+pgV4P0eWQsbUktZO1M
MN/AB32I5TVrhdhu/JI6lBUc8w474lbu1jdZKoS/q9bVnH+0A2BKJr6KLHzyUUR4
L/alUYhMy5SaZLuIgaD3ELE3L8lqBB621gYAKqdih1/Gf5kTAQjPVI82NbQdWwq3
1ms3DDB5LTunQxI74mK69IIZrOKOog8+ZbnBG17Mg81EntLKo2s20g4JDVxFG5jF
SHdp8ypxNrb3pEDzfCRe7MVfPSxXhZyO2ePQd6GJqRefK5VnsOcccc4TiyRVE4fK
0fRTZRSae9+9J9tBRpNv0AIEslAiP+fO2iIFrtPBAhZV1GgMxC8Ccf9BfCD5p1SU
RHZqggPoOGS3dE2Rsw6Ej8OCiSTx61YEmgz3TolXyfF0jphA0YoFgkIbZBQL9VJ/
EpSVsWTxdVEr18+Q4f5erbKiDjx8T0VaF/ueqrJxUU+v8Jlv7Oo5MptlRvUG4iqy
KgHSvimOrwfdmjDuJWyhpwP1emq37qp/2nwLMBFojLYBY+/TkwWD8alVl9yYj8yP
KxfBDjHdrgsxtDt2cDE1l0QE9Qjn9ZQBZI0Imeo5uE4Xz9fHzf/Xr0Ez236nv6L9
HzIVR1CPPkcvkR1SqzjEzxXvU8dzWga+S7Lc9KhjgWovLmhGS1O9hayOd5CX4csu
DSCE/Y02i0CP+fA5HOCismwmQt2xQ1MaiylJw8lxNVONB2QsjR86xPpeyQcKAzyq
MoNm8xiPzkZKJ+Uzk+4opFJplIvr+wbqtSPxVMyCuMQpoAEcVVzpb+CRw/MnX0lZ
pXfIIXC1iadwjfL3R6LOzovZLcibW1/gVXGe5/GREYW0jPwE+L4GQ4DLT+Ase3rz
ByBQWfdMdPix6EQLpCL1tX/H+Ou8MLVxxcEtz8QDbINOEogrW30SSwQcv0hUzE4V
pF3J6vN/vqZ/zMOIvDrY21C8Wtt7U1B4QQfVXckPuwuexudnEqPlQrXlrc5Y1nXw
5o3sbW+efYvyhkOD670mSM1nSkLXhuprq96lu3Im8QEqhMoBryBZ8vgzc2LYp8Va
vp5Jtv8e229DVVN0SVP12nCqGm7g/L5DD5MjEIdJb3iM/b+r5/Xj083mUGMJ32Fw
LsnTKrMLOlzqJJousb4wi5t0bLrXtKiLWpv6OplEmRLDx8Fr9B3POGrat06FA6m+
oNwGsiDaztM9ZqS/aPVuB1Nwr9S9V1Nv52gKV3zhid6832QMAtiK03gOUIP4oexU
sDQO94X/rzVoFxwWBhAvWx3KdsGihBz/nyrSnR2pl2Cnu4yb0fFHR+w0lixUV155
kjj4pO4Lm2sSpRW5MclYpJYHb4bXP61qjIYfHGkcceG0xC146qxs+DfKVF3faRo1
tHmGsdBSbLwJ6KCvsq3z6tpBJrEkpIgUrt03zSWh5Qjp3NKuuFaqZCKOk4NwFQ/x
7PAD0/OhiHgVpz8xbHGJUtMiyzTB8dwL/kJIcqTQC08VixTL71roOMCI8TDEi0xI
eKN3ahX4bPbNmvJ+hekWTux8oyIA6w9LY/l77uuZA8/pYGbpdS6GGdDnhFPU/VI/
mRQduoIe3ZkDK8lGHjCbas/fV0Z5NKErU/qgrnHF24kylnz6+udDJ6a9JBVhhRKe
y6fP5Wc6kd7wcTHZsl+sDRL3ihlUn7F6kXKq/r1y+gOheMLoJHD/U4sJjtNVvmml
djf1UPtw0J7ZBeqxgDcTCYOCGGMCRZLlIHllGJjajyYHJApqBVmn/6TQECFucXVf
L2IMxfNL78ud6ZHfgn/72p2Y1Dx2XDhiyfjM+r1sZ4npNapC1CqNJ4Xiw41njezF
GA7AoKAaBta60tqQBN2MV+WNfsFe8koIw2rllY/Vu8pcQn8nXzz+ZcLbqLH0HJ74
q1kR/Mv8cz8cKZRe5pyyebCM7/xYbhJ9IVvnd4ccNQBBNQ5fbqiLCa6S3sm2FWPG
Va0C2ci1x7b3BcgHYffy+GqkiTM+j8JhZpjpJXCsrCxbPfk4HhE3crzUr1IAGKob
T00B3A9LedsA8H3ULqn7twHoTwafVagZmkbjoc7lgARbMUv4b8k5t2xgqK6qrc+3
ZvKv4W/TjajK77oG547rHvxZR1XFgn3eDlIi5hR97SdjL+3jab+ZvAtOjYcuDqxq
d3ihQMV79F3/lh1S0LDcxElFjCAqczi5/D/9lpvAb6OXo004jaWeX4uH1UE9t8VG
DeCKSmb89RDhqyEa704gL1mCc7M7TLjFKqc5L1cxRRsI6CXUCrcB7RxxObVKm5ys
g1YB/AWnVU06BQ0/Q2zW1DGF292uhIFmKWkNSW0mU/bdezp85MdIuL7cGrno7qDR
UzBHOsZldrICohZLwg8+DLtI3exgEkeAc9RSaBwCZRFLYHj6C5+cDYE33YljuQaZ
J0au9XopSsjzSXZ6V7zlZjeO6wRMGptBn16GnagEpAOivH3CCHGWO+lVASpAJnjS
43P4elQoDdugLFOSC0AMd/ha3QGOnkQjl8kn8M3A4vkPG0F0sXqPd8M9b7ZW13CI
+6Fov0VVBgRaxq/Ogm6P3T18EPE1/4aipPe8l4ymISYSrjQupHBZxpDK2c4LFp43
IeEBuc1uhpNrqJn54WVzdStsFOWTA2EombXuikVPQZ2QHna+GWtxRxyGtCQcN476
SJ1puPhQr6v4OBhaVQY68gNwVoQ8DbM28+42BhFG5kWgMCJaGB+REpQ+iz/H3pv+
3NKH8mt9OUdHRSdRG6QeN3G0LWaWmkqm3XlRpnkUlFv9qLI1HKOkk7wwd7nZ5X8/
YMnbFhqPSQfHGJ+D3oskaMVXivJzZwaiG6R7VPR0Fq3IzP3HIUpTV0o5s4f13C1m
fdp+1ONbN1b8w65uI3ZjT4yeVSJeEMscVkBoJSBz/OjTg2eRJ6aoqh9UOGVRv1xf
XrnLZnOwQN3C+D2egfg86iIzgtfIneY3p5vnr7ODdYc0rJWMjia4MJsyIoLd3Cuh
kEhJLSKK9Pk4uejvtQ8Nz2osgq/xQQVcMMqdplpsscBNE7fwTX/fzFWkppSMTrCn
4vynveHIpg4MFZLJAQCbST6iVmYEL42wcb1n6qjvz0HSHeTaOiAVYfP9dj42uhL6
xxarXK+ovBqFGdbCErg6U4MTXH29noBCJ/DEa8BO7ZrlvPVT0LNAcbNDIFylnJxe
ePaZ/ItgLDXvVSnBawmLwGWBWJdYjpYAO4zAPYp/EE5RXIfROITIFuYwGbmiakqC
6+SYByCeKAsf6XAiy6rEep5V0QxfHONixywhimK2FDxC/dDLUv2Iqt4yTa5xsUzz
VRfYC/jGJ6MKngVknPytHvSEdiu5SjPz5VxU6HeEyTtwm1w+pJ+7yfQ9YoZQCw02
t0vvzAc/uiRWjQDRFK/3OlPUQivdbx5ncZfQ0wHOiTobeX3o6tT3zTDjfg0rT3SR
1DwCPwDi3AsWkEv809/XJ9xd7FJoYhfKNvORnz7YMg9ZSPnmoLWd3GGjbpPj2/Bs
Vpg4LDYpNAzke4LLlu0XDZMRo8Z/lHdyt7LZe6hQz57joHNvqehgD2FcQ6VxE1Lu
VufGsBP3ZzUO03YgF7f/MsEzogfhH3U0WhgfCxLeDOusO6a4Mukop6TutSrhM3xc
dhDMPBW7qEUtJDcX9DU4XIUwU0MG9cA/DE7kRov9B7/PijSnEcdXl1M2kbq5ioXO
+s/1LuZmmhv+2YP/AMsddmUBYG2tfYB8FEFZZATLTsoNt6vhzZHQVtQZq6snidBq
Wq4on5FV2zmINGycyq+DLTBznLm0uKDvOKSLLgB/4PNQf2rrpGv/uPtyopjJIzHm
wIqXkOjxrHL3fkEGpDgy203Jb8/bu1jBIqP/JgujFjumLmKNB19odoRBBfBfXb8s
ksdQiB4L8/RguI+csvVDTF2uCZ4roUoiuxxfUeIu0OvlChqodooctI2ztuVqR7uU
myPlP0cutMcbDVZDKJeFnjFesTJsWMpD3BKif88wV9Y/CeRk860UO8atKWbS1CEq
Tqq1cEcB53uVmKjZUrj6Qw9Gxcoody2Zp+obKZtj5pNFf5MB1gK/VcdVDuLgmE9B
VhRzuQPrnwDIeaBbztZbDWGIWb/PGrrbiUe9NyXHQS6oYoZXipbsA5G/v4UBo3zy
yy/rJNENzbkdYoH/jnTcZqzMXd/3jtypPLUO0I3tNse0s0x2f7ReyxqXPuUuDztT
LdH1igEXSu2qASJqraHD6VL6QyVyZgCPiHECZSYew5/3wv4sGy8JMVe7CQyJzc0x
jaDJK7cEq74B0hUyXqqO7VVfZGcY/A9sUPUo6gh2w/zNgLJQXZevUCRbfnAEosJ4
eZMww5eCBQPAy7iNCgZcfPRt8PhNHxA9pdw6fUk8jpext1rQZe6avl2pIQorHjhn
qbl8u4sDBIHtuAo0JNPxOtvRuWvgfHBXdmouUMVU0hexil5b6/ppfITy8Ygq+cXr
//gNVwfyCrORNbcwnhWSvH/mLn16NqIOO1ohqNdEEJkwoGhmX9Z5bfGIZKAuYquF
IQ9vVdintIpQGyL73NrGdQyooYtn7rkxQiz747TTpOYtj2L04bbElMyPPt5K5f4X
/dlPNXeU03aw1atCVmu2wMA4viMk221F6e8etCzmOOgfYLFRwhY1mz8/5yTBWVCf
Dbwn0sAtEW+vs8LQcmYLcR76xM2gTzixrZJUsnmrCKiUoTOxD7l/siJm/5qcl/ZK
5fOHYoFB/+MjvkaYU1xnh5JigyB6PTQDbE7NS+q32e9o9sajiziRLX8fYXUP8tN1
sX/0826cns1RgdTPzgLbbCMBf6g+g6nzLD6C8+cLJCIshwtsK3eZ+R7EaaJd7ZWV
jbn9CYiBoCMMAGoECQyWBMauZRtRI4aIqmKnT1WWu8QqR8v2iAxVo/ChWeiOaOms
KGsZnVuTT3jnSTJpKsBRirnBVMni6BBHvrpxcqxZFLPY9u1DKdYUCtm1HuJ6b8KZ
g5nA64YoMJmuWT4s6EI/wakXJoPP11qzXDeVdXapEOTQ/DA5CfQh/H65lhd3sT+g
tcx752TPsgKXtzUPFn49M6+pOSzQ1xcHvUDtmTv4YHmf3ZyHHswJPuGiQpcNs/16
07NZImZ8yfoCrBwaQo7Ad70jwKSJhUdwFocWxlZcPzKebSACDKxOh260fQZxOX8s
jbdkjN+1mZYfuV0s903IsS+gaYJaiiGDfAeLIFNcXrwSxS/XK2lLFkKeixz0tLg4
lQ9x8RQ7hj19xjNauDD3t37cntU0x+qHmTj95HCjy7e92ogAEzLps5KtMV8NHA8v
HmS9B27rVn6jYD8Tt2JeKYCARBhg3++zUwBGgMGr9LW9DM4VErcpPjqDZ24G+5uA
s3IiL4URN0Z7NBQW4mAs7V741svKSU5CEUEmvcnkiBSMc13Do/sH4h5Pe+jkVkIQ
Zah6yn2CDmJoBJP4XYuyCAf4Xtskfrocj4Nn05sDRTNNTwVBJtQ212at8MdqeT58
ZYLrJmWCE6hdQHroNDKsjdNVYvnUghE1gmnp+clyClxS5AlLjeYeJ1UXMjMwFYSH
TCBSp3HeiKhikJSrtKPL/il/yQs25p4RrK5b2WbnyfhqocD8hx8/oqQPBGYvlQqJ
eFYdAdiTzlD4fxtci0E51JrarDA81vUKBHhl6oKC6VYZiT091YhbuYgsiQH3p76a
PbV5bGy40ev05X2p7yisYsjyM0ByPLDIXwCB0YQ4UtmqXN32Owm1L+EvTaTu/YQO
cMAXbVnIME7cNKC82oeyY8Wq9JKRxb6Vk59gW7KMf8zNfpEqIOSRFWvUqEC33DWT
R69SqV18Rzz52gLS4b+dWmFZfOEb00Fk0Efk0NBfvokKmKtUlsk4cRFv3TFcbG2B
Z7yPAV6DNu9qypgMs5KK20yrxnr3Q07eMfdMDhFv467U9q9/0uFWm61WPgRt6WZj
WjWG/9w9I/a9+kWb+zaHO3G+zunj8siP8b0nvpdbqgeTVm48QpxjTMR+I3XyyfMn
zGYuOu/VgD5gWJJDdaBd9sdO9u0XxsF6uvYus3E+oqKcJPvCKhJmtZvZjg+0smUl
6+hds868X9GA7xMF6NGXgCprYAWR/3X92e3u7u8nOtXc+IHI5JizjT/BqnH9dGVE
l4nK189s+tuifhHAhGz1AYkZGyl8/crexCYCEtJmYEB2RRwS9js47pbqOLwyFTsp
Od5Eq28/+7+h2BdkB/yHayCHJaig46em12pDah1m3XRVPs3hoWCWN8bXSQgjJv4Z
kvL/CXl9mUZxKqMs1SQfsNxbvyp4BHGeobsZ5tcJdgF5yyweUmTRQNH9F/NkfyaF
5QSmcuZWDDE2gHeaOWxqj1WS2TM5sX8YYEfCBZHuK7NcFjll16W/YrZSLQkziB4A
neA4AZ+RCzHcmY7VpNwchaAtHBHCvifTbV0YCjmwpL8ynXuXr54X6Bs1wZuSQP6c
T9d9ikj1k4L1vJtnwZKISLNYs1GvwhUQrOSFfUtiQcQfHkfxVEduy97HvwlkvRiD
Yu26W+S/kDS+Ps7Qhd0Io2t33TFwy/5yOoV+LpPVaNuFUDSYa48mX5Y98XqD0I6w
04YEY/rR7/Nhcg4eWD3KkL7HOqeBAYmfqsfc3j4XiJ7vYaOiTc/iInx4y9m+5NqV
+XfkjTFAq2WOigFuLqop330RJGIcl0TnovUngcHBgSewdsOOv3K9kIuKnAg0VM8V
bYgQGuc2oa5XCPAw9MAz1Wzb0JV5HqLtHG7KqXrFUv5B9G9moufg6WZHKDcTZu23
Dp3lMnmoSzwhsItG8jCsIzbxn4boROWF+h4mqbezP45wZMKyn6LjYGlXhVe3C4T1
RWYjOIQ3Mw/MTYvIxO1m5X9Odf/WMHVi/BO13HtJmitjGKQNSP20udFwpqATJOvO
e5uhUOC/tfAiPhebcbomylyoipmbKrOquVLj1cdelibZCWENCDUn6RmYz8y3iSjp
7baw/kGDlGlVYq+3qcMMR0mIB6ZHSBoycExGkesAP+wo12hGYBsWiPynoL2wO0ew
fSrprD4F675hQW5yKNYFq3i8ssRaGL54gTSVw4r0bEj7TW/yXa5lYdqPeDc5YXiH
GwZF/4viLq8dH9g8/SP44swMPYzVd1OavK6YCdkry/tP1WQUAUCdtO9dyGyOHksC
3EG6Xfpezyj/6Y1svls0iV1Uq5DXO6JfVYAXQlXAAdtVtu6ViUhl5n5ew4GlOyiY
k6Di0sDqIZk5fdBGDyLOJTMJAibFcXrb0xlRc5XiMPiJiYwYQmSrMyvqzIRbGRMo
SJT0rhJhJGg64LgstfgqmLqq3dod06eDCfMBeXc1PKWc7FSQmgA/xeRMN60kJBuW
SgOsHMchLZGcjLY0RTORggop0IrPHrh9/3NVb2txg7f6FzIi2ZxICBBy9Tmmgv3O
SajD3/6ypcN/j9BE70Bpj8wuOYTTB0qsLI4jqXA4CBIF+rskDDE5TAQX7jNmBddZ
syczS0rIbB+Pb4+twPc+6yWWnuC9qycn6w40mVW+yOwzQIpblva/oo3DS4t56zhO
w/QiUw2CMerQ77NAS94mMQwQ64FP1hWBudP9mmyJLHFklUwCpWgw9h0dggWOPgOD
sqDxgNeD9zJNuJOF0Dw5yzd413YUUU3mv1wSu/DfmihYtKpienSatTyPXHFItgei
gqplhNh8oJmSyxIl8v8ZF1qXF0ZCtWQJjK947NGE9cF8ctUmQYH07LFiLlPYP394
d4MpZuCqgtbsn4fWjBciYfCYnpzDuU9/AwVRaVwYi045X0+jGcvJnj+pDjkOOB5l
sFrv5AvwjUS1e6lM6oAAZC/3k8EFh6HR5HnwAPgrxYyC+8BzXUyfmZX7z4CdkiWk
lAC61NDsm8PYKz0GpKDOJ453UKyxgJ77kPmXP2m5rcUYu779SaMR9EMJW7QB6LQQ
pcEnilskTFJzbN1eIWW8bHriMovu2B9qjJdu2Hz/pks6PgQ7XrJ/IyYhu33qSplr
/vjMkN17FfylctwtIzasFY/heRQYhP87JkxfVBow/ILG/+KgACcs3WbFi+3naa9I
i2EJimf04bN/vWHX1E/w/bemhsCOVGxL0vgHDdMB50zBgcJJtdwkspmHvCnU1LuP
a1niXQK0cD2XHucHvXwCnQyLwZoWV7uZzdx8I8A5hm5FHxfCp/fAhN0wtCfxSilE
LzEd8CaOYaiDO2KfpoMukQui/3EMtE1vLnhCVlHCtH+QhCmMNKWp7Yamo8Gke31G
ouxyIf124HaUnM8khk8WUnriorzvoR/qepLW6nnb4VVR6DKulYTNJKzdnqTZD2/X
DAN7gRm6OjGjSckUKWQvrjGxyKA0WHUkHAQa5wVtwO6vnpO2o1+xkfiEbhNzfarc
GlEhokaH2ke25m1LtC+GFsfNxtYn3Duo/AWAQlN6Xq5A3b7Vt9duafWbKh1GklQq
yf0e5uYLE/gDKe7yJRfw9jmfiKB9eIBRCwlu8Isw+e20yESCdfQdNDZ9w5v0G6nk
1AmdlbizSVrLY/TTGzr+7/zYLZAosJdJF0m12gxpUlM8hQ6U1aVyYWmoh/lk5nZT
R6H1Kwh8rBf1Pz9xQGkeZa4p7zok5LZXYs3/XtpQpx2JxAQntQOhtcCE1xgNUe2v
ef6tehUabgd4Rol/ZEkvMKconsI4g4L9tUmJ8peBfLK/mvnHBaqQd9jSAl6DCfVd
NQGa85GpVRYvKEjMhgcGRksMVAcXInedctjAzcJRJRKowj8Ged9YfGWpJtehRXEK
5NxQb564ePs9jlUkehBCuQ4NjIuchaJgz8ZJG7Xcq9Qe+g0CEkKC1J8fCVsoR8hY
3XMvNqgIg7TfAHXpq1yVh8WQHiNY5o5WB3xSsr/9bPg1VrBOtY6tQfcClLUq85bq
1gbODpsLDXisgCfjWks79XzC0cOCASxa8ds/BYEgKu2pcbDreBd86lbxl2w8r6iz
s6cCDMw/rn7wSxaHRz5qs04aA7FBdN7QbkIW43yOPo4AMrrEtr88PeowUTpnntC7
l7NPDw/03nwWzhG2hNewGgUWZdetYussiy8xa+bgvn3agyYQzt31QOrqeAvCZLOg
Hn4iDMtiH/usKRdtLSumiPz1V2mnuNfehCpuc4BbaDybdKpIJJhMYI/4KuvfSkUE
HeeJVxJM2fDyGWr65Q5+RkylSsM4vC565+vMZtwBX15t1aWGrjrdj1ow6gG361aU
zhWcK91JTP6NUsksGT8I88bU4pVfwETdDEef7FgRevMHuy5moD0HKJMOku5+SKAR
PInGZHNCMAr2s+oHd2C5ENhyCpMkibGlBG+Bq3PDDBZOFFNGAlcuyMwBc8PxX/Mt
CjfNTuub4Y8Z/FXhCFiGndDHpHERTlmpwMtjzw8eVdTWtlLyomrnMYCyi0/baxnB
yXpMHjNnVifKZCKjbUrsaFUJ4S1lPiXW/I6qbLcloFCKzwU3wkcuAwebUKm3lE6h
Xlgt2o78y20LyhnNz+YM6bPLv9srm1hw8/adwUkLI+X8cxgPfoR1gxptAJ5WwBWW
+3DV65LrCkRRE6aKUNAJhpYlTvJHBB6PXHZVUA+aRXgVNBNbeos/GKCrd5A96FbH
v3oG+lx5aYboNoESB8m7N0p8VUfBK+PZwoNKy1giqw8tHD0KLbCbjbiUo9nr2kwQ
ClXJDRIiIjtcnHR0Rma3WNekv4BMA2/tqvLa0TM0waWb0x0chbUE2UsWFfItPNL5
H02SKtCPmOnFzcryXgHQuw8aA0Ee5K1qOrHple6rPdTTWsRNPP21zbrw5jy9/KE7
VxDr178+8ObQ9Znt3Sr3qdNZuCCTeCDmw37ors5ibCyjxPXctNnUdlJ8EpJRMuZr
HKHhelC0I28UZpn+KlB+K6BS3JFUkKQhezL8YLqdemUkNDH7SxYR9g8h5ILUlDQZ
YTay3jSa6GObjuvxdy3gP46e70fXoGfbiAJ43qfFJ/4MH5Lhwi8hJw9lOHgIQPdE
1kXIT8Js6La6CEXxdVMjt+ChVtL8vlPCOd/PD92zuTkHVs2DsyDHOvakMhTtczkp
kq9lXTPMcFTdeJK0yDWj3W0XjsGKxcmlewkpjXdoTrsKtW8cW7TvNBEtWR1lK5+Y
qwXy+ioUVZ2jpotG73YupXsz8GKUJ7Au5/Nf3j/rzyGtAANkItarKTlnB/xghKo0
spLuSWlvTU+DX0NrFDlL+tPFhnbVk2zDhnWXt5Z1kexhwegqzAMHalqnXnUxn0tJ
rZ+eRK3bf3rVb3D2ZAEesNHCRM8u5iDWwdH3tOFMmEeB7XfvDuuQmMnIl+vSWO8f
T4oNgRTSCvNZVWEIQO05oSTQjlvMbq3sRVrAHWp3Df7fvvvyXnGY1xcoazj0R6zo
KSZmr0ZfNVF+s2FfFYaizN8iS7MitBnaWkcxQfDWLssbPrqYfPHhenYhNHBfJ9et
cKGpqpSeVUoLS0t3Q9OI2sCm1sUWcNVwaN2UH6hlaCMhHb0VDwSLAowzsdk4rX2Z
HoklSue0UC4kwfYyHQ+O+2wRghzO6N4TlliJjJXU5gMN/KfcBHTTTUXTzgVVexJn
b4wHobuwxKmWCVSPz+dpoOkXTBb3XyiG/YdT+qUtn3llZjox0aBR8Ix91w2TbKJJ
m1hlQ3dIkgp4tL9T1lQ2BMu25KidSBz9O18qT3poZXLkTE9aswQHSRCNKhmPG+iL
8xJHzO/ZaOBaM8WQrzmYoeZMASyDSh5LgbPX6MXmeKtsvfQCFKnsU/Q6ST+QsiS5
RGb/SmMgZ/l7GjNds1qyL63sdfsdTwCCHXsIJUaUV4+gghfbOyqArsFOKbCRDHjl
q3Ygas1R/ATOhi7BzAgt4808HhCGRw/1tn/tluu6pjaOYNCwLWMkNVi9VYYG8K8b
0UXbGdCTY6FERiA4DWf3BjfrAxZ5uYJ2WAwWVhZHwang89yxF3CJuRXz4zudof4k
PP+7WCpWFMazloPqofvlgnIir4cmfxn224LB920Wtlo5ovVvM1F91k6qdPHMWHP4
NCX2hPsIbfis6Of+I4J2AnE2e95ztd36AqSw0Hw1sZ5Y4R+Yc91Dm4PuVPdZEmf2
UpOtETJkltXJgChnsk7V8yK9XzUy5VxL7AQMqfoQc4PWeXiEJ37nm98zkK6uaSiK
cEhC5E2VC7NzUVdKs8o0QrWuQCfAUa1ZC3CQ4oW7HMJXjxcwWDnXiWYZUKNonqGz
So7lUpAU5n2E4pSQmVEYxyEVri3+45okD+s2PMyLvtkl6dI6CzEiSETLvh6cJ/Kc
05z2o9HmqELTJo3pxYIxRH7QCxjsBaxjNPo6LJtb8pAzIucuzc2lp5KZGEw9gaV7
gS2GoY7gIz3+t4HlbHB/8vGxtGWiofb6JzoT3sgtkxhCskIF3+9XCUrxD1Yv7L5S
Lu9QakPxqBtxa+QNb5rhgD/ho2a2sdYTQ4t/bkg0KszQa+TMQ3VviGUX7FPBFBX2
anT7ip8pHr1w72DFQpp1QTOjvWLv6+Ih/7jG53Hz127cZeEGhk+oU1ArpHoIpGui
FxpXkJ/ycI1WuCR0bgNvgo//KR7Gfv1X12yJfBYxYW1wXd/UqXBIjXFf3cFu8qyP
s5e1vqnvft+x42SQIHs9PGFH+MntmtqPVFz5mKYlUjAxWZCM/J6/IiomVka3AlBa
LzRWs1HyfZ9fZ8+vjzIXXtQXVZojYjDUghxqIiU5L6kGfvFh+HnOf923xDF5Vino
IGNXtxR0DiLhyxq73vDZVarIL0F3d1nX24f2uy6Qgedv13OUcQWxUDxAaghS53TB
/wz9k0Dm74I6Dc1G5pkk4MMvuD9DCrCB1LM0M6MJlk2YpDfysBUgDJxQlcqcxT94
wHdroGWJVdUixer2udz6aglUs49PkePribX2i5eO96Zv9n3g+k0hqSPFSdYM5jHu
IT6Jsv8s8vxnsdnlo3viuEY2FNnaLf+lKZbJ36/jrdrOhUOiFYW/kR5zs5qUcdbg
vOEIUNXpkzb96Ctwl3UzMm2xCiWW/8YerSLj/Q0dRtpkHe4lK1JButYnd7AmD7QC
zhTRiSlY3WbW+V5OdRZ3hZOJkuL9O7uUvTOVeBqlP+OwDgftDVzk2qHpi5QWZW38
6mfvviwAsdHAHCjZoM6FACajUK+pcXEOzroA0O1bMPlHev4Kh88g7Yu+GUMNzb12
Arh/+6Am3KLih1nbXbHDr6Lm8kkNVn0anoKgO7yLXS/mT4/IH2SaOcGs29z4N/FE
B2xQRciKbHkt7k+cv/uNNQj7Uq3pMm0UPn84J0yoDzQV6rrl4slmMFO56/sndtir
pMYNf0qn+9v4NaiDn8PUW8Fm7jbayv3p1tU3oZQJODjFY6cvW/hQNgvO2zywNDKQ
QYXvCVB8KRXV2+a1qBgLw5aB6epycjgKb4p2FKyMwK+vfoezlwEx60JQiJgPjIb8
EKpXj++P4bn9SCQbvUSy8O/4RMgtnRMS3kfrmFzZhe6gbBADTdNKybCooJz6imEK
zi8LttgmuOJLrfSTXnE/tpiSmWL2h8CDdhq5pt10eGtc73et3eNnvhDYRqLvIku3
yvfilYU6hdLfwz4oxvSzcdxJivSMIA6qRpXfPfedCwevoBLwudgEXPoSzsW35fO7
8U/CSSfEAa9a4xmauRtk/mknl91QdS0T5gfy75mQM44xK16k9hRiqkciLF7JXyTW
gtimjxcAQyJfFEz8/evMuqEU9djb6eLY39gUM2ZjcR0pLasCTgP4vAzhFT8ltscb
9zFQ4TAwKmwmSUwosonIgJVdS9Q5ch1J9XfO1reIwVYlNJ03rQHufirXOTMcJmkV
DNzJDLX03QZpsyEfZ3d+5NFjcaLf/l55Dpiru5+9SY0H90KnUDP2pSbDWyDT9ves
EGohyMzyJ5vNJFWz27igvFDVK3bl7GsqDBoOKcp+tOkAHqj4NUKILui8DEjJbEpO
lNVVESKDEpa6DeKK0ps8hRWptS3Sa95p/l/xgkikwmGxQAwAbTyvBY6JwT7XMrVt
+a6Lc5cUgxnOAma+KteDijG7LpSdFqu+nywCnrYEolMbpf7nRqpQmIHSw2Kh1pwp
U0S5FDKOwmOohEAS8qJutJKDJcyferQBpXhy43WHiw2SKhqRHEtWvoGL9XQnUd5i
odAHlQc6Qd3CLZS5TAw4ROiecNlCAwBgmgfB/w/Iif4fZfiO3H/QCyPxFeGKPxS9
jGgG25gjiA3K9RnbBmYZ++kDgC3eOqwWfOFrdXQHchXcgsLHoFRJb8BkEUItroDA
gwCdYz7rGqYO/7q8L1Eo2HUcJ0BIYEBy5h8YTQ5gHKd/k3R9B9Wuc04ZYqqRNAcH
5Q82n6vf7ZLW2BrXSDXVH9C36G/izcHARvaRczyRUYxJ39VQHt6XuNwmsmKKR5vN
DUPuRC/hH2cjGFq8hYJdYdEtGu9410IDkd9ThaGvPExTr1GQmf+5x7tNtJ4k0rzN
AMvwegCalnMzbRMHUZT7bH0CDIeePj+GSA9i5nJmc7Hi0ambYO6P0Ny1Z89MMHG0
GHAYqfE/q8GtbYdoQoVxlnmybBhbe5QOvoBEyjRnRaLHDpvelWds66Srha1FNCw/
Ve6UgNsjL4zhqrdEqqhUL+rDJMUoAwgpcCbSLOJPG9EwUhS2Wun/NxwQyOxmIyIW
A8FBe5ermREeb6HfUBmGSTR7/q92Xf5+BonljztJOktqtd8EmnyVKnhC/t4Uz2Xg
FcucqfSYtN9IgHW+wC4H32tHzqOHDruADjLAwpke0ybNlWFTMnIl63VEZV8UlP2Q
yHg05bHYsRfWcIDxhdHfRBDf8Mqr0F04kSOtgQoTmvtUg/p2CK8KmCNl9IeNJAar
lSd523CL7bEhqJLQjqCKHxEJkhea6lEJqxHAl1ebm8vMhuXlhR6QVCZC3hDB9NdY
njHp36SGajlCry+ZPhIFI8NPSMqh8SbQBnVAGvt570oHTMcw7pZNlLfHRy1th6J4
/Dlo+EUTzeH/p3fqUEFg7TYfngRl5AjISLzQa9tnSh24rh8ngyKf/1saqmTd7aRg
ZQgVa2+lJDQv8AdZ5+b7d0V4QKPi0ZHE6nvzC7N4Unrfp6eZRfQGl2dodOnuUuf1
PDPxJPpP6V079k89VwBJSBpv4pKfmqWDV8RLBz84XQCkP9Vxatp/JkoJB0p35j2r
fqRDmF2fL1E2vUmghES4KLSYAv2NdQOvxYGcLw8i05Z7JCvx3GhYX/Y+bPA6+4CL
rGBQvjbp9V3v/A3KBScavIzlPzGJGdY49OiDZ7NvEXvlv+6wrgJv/0Tlmx2a08KE
QW/8vh+22B9Sy3oLUqWU2jVkUz0Kft1ZsyLNHQlgNVW+sMQREBl9mHXoK1e+JfNm
vuCVHpOJ9ukK9HhkUKVUNP4vbpPqeiAT9ljsluJW/I/lZTE6VNNbZ21CkuSs8iNC
GfIkuA4Jr9I5ntQShxcXr07HlHctIIwth+M16vUpzfU3VBEzQp3GtImZFmFxRvK3
a47DG8Ejl2gRGM6/cE1MeeAq+Qye6onFo/aeB2psAeSBC3riNephwHsioEyMaTqM
Bx0puUGb6EkvtrklAsZZznjYVTbMbw1+g3SO4CPOuhN+ThJHBOVo2oosAl8D3xzC
fKxyugwszxCZbwbkrPL09HU4asIqCPsaBQobnDq1sVu9gQ+W8IAv3NaJsKxBsWxD
Lrd8DtTIdS0VSSRwrRY7RVlM1+tdxEYRXMREvjTtbOjTaOKApL4tMI4D2BcT65Ou
pxJOExvFBOdQ3c4WsiACCXiHp82GBjH07iLJqp0Tb7YqnrtZQdja76HJv2LSP0yP
EnaOt9qTBK302sg6Nu4LG5QgCBsszWs0THD1piDUH0o1WSPIqx5QUEA19fn/0HbR
9fO6sIeQw0injqvOsEGllY9A8QUvW632+aGDiPhi/BCJieXi0Kc9wsJsTy4S9x5u
+zxp3Ag85HeXG76pND4UJXoq5ej/bkwFZD+rriFtGAboW5I3GnT5QVVuylxFcim/
0Fm9RdJkotFajVagcTio5nyaZX/t8h9G6dZSB/d2dtP84wWumUbxkK0dpCQkepcQ
mzrJFsmMLUROK3NG/KXkWkPGZlA//VQk7B2HlTF9kRwb0e4v4nK9mhU4CFIXwRie
cYPOvEuaVqAGyS3VSApMi+5bOGwXZ36CT1W2yxFSiqj/6Aps1ZmsqmLkJhOjGPfo
Oj5D4oiuf3NMQ8VTslzPe6QbWRDgf46sI/ZrYxdCcjjzkQZY/pD/SVLNu9jT9Cqm
C96jEACtB+RLxi8QNgpy3lGw6yQIQNZTF1EYSkvIjSntIfoqHKHcbamR0sJjgLZZ
RMhfmTleOvuMXMuZs4/Ct/Ai0t4f+RBiymHeB2dv3hbGXkfRuts+jjTYhGnhU0FP
5+Gi9+PYZPkrVY8UYETfbioO8KwjZ0ogX1aFd7DzUdattbIeF7aHChey+eTfUFO/
JmT+T4m4yMDYtUrSV7HpWbCQjDuSWpE7Fmky9NE00bHINAPGdZnOn42S9gkWZznH
6aGDMjQQoEtV9W768Mblw8mu8v8z3i0Bfx9d9fYOF4ScRy2asm3CR53CwiPEjRBM
DQTmzIWVT/FCOUApzSzyzmaaM2fZynRXdVZdUKfIb04cc1FoH2Aaj+mFRQCYp/K8
KsnbIEceE6OM2HSVqd1gF7XBg53nHH32/S3r3vDsuyKloHpMSNcTQSpXaHZ5MA3L
ROo/dOa4x0VeqUcpyZPeo+fY4F+fBnXaPBz8JyDJ4r16ryEzUhXp80pQ23dY1Egv
GHT1DVEMskioIaIamtiTBBuASJBE1nWVi67pZucxaEb5/7/PO9NfslaqqteNDCWK
7GUZ/pNImxLXj92NpSfWWzP1WHCz+ydJnou6utJZ8pLpe93pgT5kTZV/F7IoDDtX
ikTJNLSlRF2LTBBM6O+HEAFUESoOGNjgrQuSuySNFc3cGpT/PBJEKcWJu7bbKpif
5gAhlpEovYxnjzZkYSJy47fjOYxXQBevOYZeV+dPsBXqzhQN9yvA041XUE58d4gO
2J/vHcGeLj4dPnCsgojFf2dOi3oOt6BM6omOuFu4sJYjWZevKPTW3xCge6fLjtmW
CvwMX7E/7u2jY9vJUkRLFAsB3sN7ppZnZ0Xa181bIjJrLIt83DKS5ib683tdWblw
qgXOVdtjq2DVlTGSwsnV3ejf4POB5WWoXeklOC2Wi5SFAQEOi9OwDztLdDssDHTp
eQhs++p1jrQgvux4McwwQU7HkM95E3+micnikXikyDSbAYIIrBuqfTFUDBSJhOB2
Rp2l80cD33bCol00cH5VYv/dhXgKwXounXsb+zZkQ4smTn4Hw124LxPRpC26MGQ7
7l9lmtmJQo+ZfVRNVC26GHuPVrG1yOpFbBHhfJ+djPRyUucvgj8PQMJE89Pyajl+
ZJHXPhzKHbcIR7GsVQWTsz/+D0pA3trlnUcoEEBOTQ4+V6skFQr9QJ+16wSwAPHL
C1szJwnNJp0yck1lgmSkjeiaZkxmPZFSVzhxQkb53FjaXQeFiBXOwccs1cegjJQH
fq6gafSZVjNaidUibkRVjArzRi/ab+5eQZTG9bICVG5OPzHx3K0kXmGsXx910wKP
CmxKkNfXIJck5pEezja3jjpwtozl7nGGboH0vYnCigZb7kakiXMDYAvEGy6ijazv
pkE6nR5j2H7TOjzu8BDK6MVdTeVnGgUcgJEZWfOdbEflUvX/9oxCyDZaukajXGOv
P+x/IAxLPvXZZGY7sUNn7hFr91wsjoQYTzegK8L7JweZIf1bNgG9rlfi4S0WInTl
5MNe8WCG+dzkDGonHrlas0mXufIRklcZkemrAdQc7InJFnt75So8BA1CY9fsoHTe
5FPyD3fgssl04tuxfKQUKaH7lLAPqrjBFHT+zfy2jAsuozqf3AWMarlugogXAUqM
ae9e0jQvj4f39aQ7qT0Ofe7Tbpm+6riAtZ5LljZT7iH+IuaQsXYuUOlwxFmpF/0U
D80Rx6M+E/B4rMJORx/Cq67/o7p8v/0dmNrzB6AEb0tIF8QHYx7DUmLe3tkk5nIO
C4EMwcmOAGk1kGL3BOl67LExKTtmYPPUj/PV5P3NApuwM/wnFwD86Hbq5jN1Ul0C
u1T4sjIyU7H6hAl0DY+5bISPbNRwj+36BwodUTzQSIBHPro9QX2WX/Ltlftchem3
HqXnNFhAWDqQNpBO3qdKhgeVapx5+vmohfV7MWF1aYfLrGhSB+/3HTdNP5AE73wk
rkTs7KHlZ3fDP0SnJofgtMv5bxh5kAIDrp0TyAE0yAO5rM+P5MJijy5C86OJ42pN
i9UqRE47pLANigptuIsgGZa4OSBI7OnAaLJAZZfuwZoNdf0R8d6Dki99iVDaYMRf
KVvWQhPd96X3i6KS4/5MnA2BKjScMTUqKwrnk2ymMMDVrYQcMk4ejq6mQQlMiGzQ
JbJhGSY5y8NVowZ0+HxGtr6rzVPDYFKqPpyfhXkD+VeUkq7xyQCtZFq/qzZ7J9I9
AHmR2+4JCQm6OZrvjzHpUgnkV1fDb/Ol42NOE0BMMdPqJJ5QWoL4hp1U+dkaeYjy
XTPdyQR2MKcixDBdfr6lHtxbgvpQg4GtXKL83EQKh1kWMCogIXzfIUIPKqmmkca2
GT00Xug7vhQrKC4uWDzcDD5V5xmExnZjlFnVRAH2u2j0CTQfWsj+1o9iJPwZNqzN
InN31bhAkGFL8f41vs5kChHEyWK1+l4/aubLtsegXXNK/rXDHB+bO2tWwo6OtiJx
6fGofu8O9PugLqBYySbvDcWnjdC6k/GeoQlCZhH+RW57Ezzah5Zt6j7JUQhOecbO
R9qv1Uw+qPS7YpXPU3TiR3Sx+MuW0LunY4DmfMyg62O+Rey2UR3dam3TE5e3SBwh
oVF8pVL/AYBUx+JwTfRKeZCfWDQ86qORTA6Vm3Ul/SE8cFU5L3NAiY8t1qgLrDN+
BJPvUFgNBIywVavQ4s8OTKxZ+ap7loXy5G6a4NddwLuvRV+sZYojDgUIu8BLYEgV
VH1+Y3zP0kAjaiBDSqlSNo11ajWhsA4rPHYk2qPlydG9kaxkyPlNqcdssBF4JqOt
9uyRs7xWgcdFn2ivxRE4Q9euTi54oMAtoEwroFzuCHby/4KiUsWUMgxqnc9p3usc
CErseth9+S9hrfTlzyd1iy9gHIJvAWtICWibtyx0rYiMZjihPcawCpdwC1SC46g8
yWmh4IMwGX79e2rXlDD6uv1Z1r7tQJT3NZ7sskETH/wKtmYnAzbOsC4inC9XEzBU
hxgUDcWdzwyCVNbArA+yZpCNaf4pbY7+wbyiU1GvFm1aKl0xxCV2qK9rsymhWT3x
6I4VegNfva8ggeEsP/QaA4v2oT18KPUK+IVh8bOVb+/PZv3CnDVfG6JOjcvpPJO/
73/1w2Rpxjs4Mcn2E0Sj2sx4QDEDPpZTNq563vbPrjpixi/O8p10k4mR1eIulImR
Q5W0Tp9AdeBy4+5RI/D5h8kdQzxdq+e7RK/Mm0ZpUX/YPaWy3+ftpnH7VfI96aWP
/JU+AcE+/NkiXTuHBz/MOJ4/m4XyEc0W/Qae4TT29671WYJBVpMo5tdH8RNt/EJ0
g4TO3FdSyA/iyBaRdZ8BUWKIU7Dtz7BN0t2bMBHimtWFfYQhQu0cfs+I6Hebi4wZ
298ZOpQwNBACxAtFvqNpLRyz8Ral8ofs32eLtd6Aqmz1dFfgLSY4QvKXteAzz6CU
27QdX2GD60qQDrVfek9+n02AcpPzkJpP/TmsTG1XFoI88qzcYwC9W2H+0SX9+AD3
tAFuIIBi0htkFyUu6xPysEfFHAOF+bCLME/st3D0+i7o/5MmGEmCPGoUXvldJiwU
twxB7XRMDnrG90qrll3y/WipUVMv+g/rS1D3vpvhOI/61++CXtLaMNVuTdDo/X6C
4NE+u4DJ4zraLcLCessVDhnDLV3xAdwJ5XsRuUd5+dHP7eCSO9mw8oEimFcrzPvV
bYOgL3y+XwhDJ0bVfra4FoE0SuaYMOYgzoTII4DFq2TLQ7JNoUtLlTTaY4UPuK53
njLgnW5yOTW19aZ2JBrxM//ftvrlAVyAy21gdlupmNTOJv5AEaLRic8jPd/h9crB
/P69IFgibvdlzMudNXE3xJSZ5AOVvZdubhoLkamH/0VGh26QBmo85E7fulMmUpTH
RB5SaR6odLxELVeGtqzRFuy8kkEmI0G2PEC/lQJiQ+7J0mTDPyU6LCAmCrz+OFzP
ijjvcsJB6bvPCgH1yN3yJC9fg7kj4YlGUuf7TL+bvUAaa9ItxIU8nrsE4ReJWr9S
CDrcbnXDP1zdS3Ca6hr/L2iqxXkMu0U61W8dZG/fhW56P1xNAWPJY/MwWvnSaJwF
kLEr3p5Mup+54pwdcejHHpBc9C9TQppMNYCXFH0sXMYy3TRoijzEqqOeu/tnk0EY
S6S2X+DiflBRNJc9lFFp3ssPIlb3nmOSpHdPLTMBVFTCJCnH+1Q6a1Dih3kLgge2
qvOtwl4zk8n8ajtIw+Rn36mEHEUCkniM5Fp/amUgrwIwJNXceJ/2PQExRtq+EIie
P/4HwWung9fwLrW2g6CZW9zE65/CsqSuUp9MNavGGWbrEDCgNn+IGNT6TKXElX/m
N53wyLKZ1jO1uHhjStrlWdOWrlTH5V1k+pigjHtjvP6JfnTk3z0UEa8Z32uI+dBX
NB/hAAWcEmXtJiUkqqzjgxK+cdEwpnL6vdggvtaiQHtXhFzfE7Y/fUCHihVi4s+E
uk3wnZH4iI0QxLhmTebVGLVwBzWk3UUYaOVQ0P3PZky6wgPh2xGdaUlASS/j7GeI
3DIKftdCer7TSJ6s4GJDURWVTmNDMu5qmgxelakc1Zj0k2ayrYwGpLoc9g9hTIR8
54E+NpoiPetyxJBA4qJUmr1YP1Ca8zDRgCiwxVTK9sZJp643PF+ORTdrxgQgHzol
dKMKeOAR/BcQr2GmBN9Vso/sa25duPPS8wygjHlsl6zDaYezBeY0nTo965UWWHlC
Kxp0M1Jytcp5zxtFebjW/gIGulx9u7SGK6HUfSiDQL69tdk+C7gSYn67l1kZf76c
1Xb+DgHu//Jo4Kj85BIJRyNA0/sEJLy5IqJxEWStrebH0DKgaIdmaW3b7siQ1WRD
coSzltkL6SqJ5yy9eEOQ2sBq745o+2DBI6lkHwF9+CpNNFkTT1WM4yz2k+u9ZCJq
liZUKa0S0U/Y0zP0VO+JeRk9roJoVHL0Ov1UtcsSB52+CKBX7iUoQUl1Ue7fp03U
KC5/RiM//9gHq9oXWxZqnztighIkHZIgojQOKTHXm55WLVXfEHt8kojMAOJaSOnZ
gUtjQb+FrmAsx3mqThF5j86Nsg2CWHadjNSDSjhQkQxiqXMZmEUJdhxwM/vmJlx2
3m5w18wKCCrDV0LRAKfVrK/sTMWu/gTHHXYuCLkcy7csR6NHsahIwMjoi17wgkNX
IIJ357Fy6LqDrB9LtEK6sBxOCkrzaSkgEbQk4nGcaUdjrME2sM52SCOKVBbLUpf9
FC+rZdjHsYKIvmM1bZw5dmfQNOfAsiF8lBUrb7x30V9X69AYmdoK+hsgJQFdE3q8
mBid6kxi5xBrOjwQmgQw+P0wweXGc7GEGKVk1YKizLadlkGVWOu6DmOENEYTI5he
FTct7u6rvG+pnZrSKlF5m/RhcAk8KbGoRwvxQHU4I6kggIbbIF/rjgAYP74fSZ87
NBboK1SsjGwa1fnYfa3pLAD/JIyW5vZUc7gYFn08KU6ivXQ2SdY0RJIc+1gR+3GU
kvdfJis/D6o3QngFPvIEiWLt4EQuSieKmLDv0s/FrNlICDqarc6LrI8oycYqH7Ph
P6xaEP7xd5RFYGfValuec5vqZgbFh9oBCYxJi3nv8UhPj+6yV6/E/TSuLZWrSP3v
7D5ga99qytFDbxWeSB0WK0dkqFmtHLtAZ6//Qt4E1g8GgTxzY0DV1Iu9XdpjVjMA
pFnvl73Ks8RXINybZPISnLqxRUZdwA9L//su1lv4B9mxfDf9QLlSx2xxP3EzRYNv
U0piZtD0E3O2nT9eDTDAtt/a8Rag9nAz+TAbkF9z3rCWFmGq+IUI5aVhGoclxEaB
u6FTT224jUmLJiLbpgFVcAYZcMjbeHSlnag6m5+6mc8vymAvpZgkpESV/EoYs5w+
BAcm9mAuUrxnXkoP65OLSyuoeRM+AGFxJKGH1JG3odvrvj0kwAlATO5+g/sFaXCW
mmgNTf9EjRQT4qMf+30gKVrM38oz0IpMpC+1EdXQSaG/f7b5EzoG6HtUHdZ2X6Bt
bqhU/mBi0gfKi8uh74wDDN28ezz2HngRLJ1u7vwlQaMPw0bIdE4+NpzjPMfX2E+9
8dNP2SHo667v2f+u+eyfGajeBeDjiS/7pEfUK+EHOaq+pfpogwNOiEfrumhEVfYm
p5CIopF+02lB6IyjICcWvAjh4KS9+KxSkKVrmw2/hbhXlHu4jYROzoB48ypx5M0m
NDCHsbrMbyUz8odiMlaZLtVxlUWBOnzmCtdvJwaE0N7jS3EBiPFby6m2y7EZ+9Rg
PiUYOTkyr9UQORfgROuSvkmiYISu64M4oJJAGjxGyWDIBj1YdarU6uSQxR3rDpSR
MtAWmuibXhLR8tV9lulptBmi2Ba/JdnDAUFqNZG1rnraXrnk5L+mFO7AfAcTajjJ
gFwl0Zq+WGolHBSgljtK3Td2xeqqZgh7N4fgqUkt5hc4BHEeypwWaLefDbarFs2o
O8TFdEjhJVSGWGxB78Wd3WIDgJFDp6WBLVijcdcMcK1LeJo/bDG17C8cyC6cS7/T
6VYAPP84zjyfa97kYQAwgL/vTbRW6rn17D7rK2CpC6X1cCouFSSBck4GwIwpAh9R
eM3t/AG7Kod9mH+L2lUc3X3gfdhp8IouNP/3ZIspRNXBSzUwKrEL1YV5v9Q2mJhg
mDCSw7cqht6epZ5mHdC5+i/6tifi4TlM6aFx0nM1caWj5aiwP7on8JVtE93OHVnu
1ghvBvUgdlwBeDU1jvmz6e+ERLZRoq41VqG1C1gtNvb0bhJetQz/YUCiUXriBECZ
huQNf+5MZ//Fc73fNcJOnPD61a/vqiKhuBSB0XWcKRMgwH89cwW5uDpO+tibFB7b
HVD1hlqaIw2z9kuTWXGQ6QWiwg+ZJ3MFoozyqJm1C9vYFvL8f/x5RlxrksZRThAw
YoCd6wtpqXlJ1sYaYm94rJ4gqzrcUio/ZjKe0jO+dhChhgu98to40MOG6WBrpu6v
xiNRcqq+1T6b8Fr8CH54gvEme7yG7g8yySWk3Cg2yrhnbx0u8QENUjVj/42gKkrA
FKSqpGS2skL/ctHZoIBwZRfNABR+DhACuRA4T3TBsUFAdzoosa6FuaCQtLTAxXTa
K6lADJTn53+o5Iywc7JQowPq4veABNTGlGyCx2W78AM3LHWXvXfhcorxnZPvUVpM
i98jgjKqahaI5kyi8wygFTZHnXKEYV6PxyxG8hgTF0XA9QzQHg6oLuQ9uL3GAWnn
O0HvOLXI/GtWjBJL3WiHvNUIYx/euBIB2w1sy2mTUoj6esdKihVkO2mA/EPsq3P6
JHR/rb2DCI9uYK3IRpFtcRAyW5Z9PUoeyPZVGUQo1b6Xe2SEr8oDZ53qeMkUXsJE
3hOhgAMcJUrq3r0laCbVc4gQhYOwqwHU7fjhrCw4cf70nk+xmhsj5R/woN/JEY1Y
02GJE/FHG1HodDoAcZ8bgQry7VEh/1KwhV60gt1Mp4/jhdicPidAaZZS7k41jK8g
qFyx56vbPbP+LSnbCGH2y8vTy5X2VBb2ydvzgaNhlq66PlmAKclJlg44iPGPgTir
tDfzye41AWseLZAqGcWwoVBF3jz6J/J2DuorHfix45XxbXZLVpWCxjfA7waW7VzM
7eM22kQWKrzZZWCMfZwIxKubroF08/iQY5Tx/ShV/tglQdiELjQd5OPNH7KBosxy
aNrJ5C5TEzXxUyRmkzSrIgUhVnxYxw0tvw4GPIQCCwD8DnZOa3Y/7MZg6bUi099S
RHAs8AmDC4cNfhMxEGHZ1mEM6g+U/nHcjoarIqAO0dGS+/oAsPp83SPhKpZ1onPz
iB85SWN3p465KKCeAalW3JvM2/HhlWpnKGL4ZGnGM//JaXNad54nJFfwnGD2rcvG
nUuxeYzmqPKrIgGymzE5EhZirwKTgSZWSlKLw+eCbrt0YSXlr0bwuDbqXiEcJetH
W0WFaP4754G7TSLJpFDngAow0y07sr2vIjntGCmyDae38WeCvEidWe3xohNhK7Su
6ebanO8VPEz5sJUsMQ0X+1OxdwRsuxz3V0fWqcWFsfMCh0ORM0pUTSSbvePDb7wA
4qPgw2uitSfbi7tTZhp2JH015SiQUiqSQOL9UavKWXYOG8+ZSgDOtuGgyFmPGyS3
LH+CjPEtbPEBy9TWjLWU7qbOPqjdQ8G6G/u9/B+gL2qJzMjiFybTjilODQnoELqj
PZRXq/5ASwAIsHXE70vx4sJU4Amgxysb+YSe1awSYpgx+TOVNF6EZXCHCz/WQQ2z
fmqbtD9CjxeoLORgsSwqWrvnmgGIH3bWxP9JIUMEpJvmCEd4iWHi+hJwKZcJRCVY
qIiXOWQwSVP/yJW5RUZ/1bFAsuq6je8yniF2vWLpmLyxA+/5bTHf6cgx9k383gXW
liVwxHSfS/MBx3g46gdnFLTLhFDJPWlcSOkKiPVO6GWTXs75H+Nw88T477RTQ93k
JCftFj/MhNL7fffWQee1qgETQKd1HnPZVoIvYPjQ0ztOvfwJRhi9ScLstUijrlpn
cvxcCCbaPizuzM6dIov30mMEYbEEtagtR/EKidY51aNC3Z490hY3N831ks7CEKHe
IlPSNpNTIB/pQlyoE8Zv97OoVfpLfGeX500oP8yXK65wRzyKbAQMwEo3C/JaLwaf
j6HyRDiJyFtpfiMCw5Snr5JJ1iEu4EEsKAQamdXhYxeD9Uph6j2Nz+nKG813itxH
NeGmhgsof6oBROvsd7tDXpmjEoEgW/ani5i+KaP7M4sh/YmB/oLLwZvOyPXv+4fD
y3TBjLbVYKA/VZ3rdhNyeL8NUkrkkMl3twQvsK/Z8h7XtQZ/ZgyLzFAp8WmjX4Ob
T/pLjSO6aQCn1V8ZK4xbBRUJHTKquJXJuJm+SOcYHx4MKlY9JKLDWk9Ghtzfxs65
udQOkQBkFQu03Z3zU41rvcqGTgweGQC4cUISyyVoDGdpcaFu03JThta0Jwa1n4MZ
EZQxxr1sPxfD3G1jiB8Dz2FvYuUW8XDxLzy9G+74q9LiJVXFchToL93HdFvaK8RG
2tlPpksftU8J4P2PKwopE0EhxpLGqC7DpIkSZ9IzB1VZoPMbr3cX1PO851y/8yfw
JSO/TsPKMXW6m4GQ+9FdAGsezxNqKcZsxnKwfxLTuXBaiaYvaQFr+zE1EwMP29iR
/zeHjt8R+W8zFozZjTxmy/pmXuJJw9clnKoAkCIUPst8GENa0buLFXXrosJn3kM4
KwjeSB4PiEQJSUCQ8Pk8eHp5GPUKSNjDqrh7QX3RhJgBvaUUHVnqrseg6v7w5kzQ
HBOYzjKH89gyNlPZcYgMjEKIVcmZ0I4eYMHSs4WZoidxUBEzcrorbu12hzkUi2iW
jGNHodcxMxbhcV9ElkN6SXTPJVuhEtowBvfnuqR33KPAtJZSwJH2u6VS7Gl26Eri
e+WZ0AYw1cW/FlGOQUIUrTzLwj2LH8S3fRPme0LC+zyqxrce3OO/IWi+X9unMgxa
fYwpEFwMylvKE5dy2PvlKilRBdHotJsFMpvCGdUobhHl84kN2PfNvNuJDUGb6add
R8RkJncLUefuaH15LAtU01VrGEnmaK3QvB/ZysSn96XDjccgThKVxXLrIeO0GTbz
lRNNriPydNYcHL0CfL4b47Xszp+1phapQ9no9UlCHjtpe+2vV1WT3g4dvln9BL9F
h8nljXisLwv28pcgAuouvxh5/cVKB/1EXGmQcY5+58m7BXfIDZWbdfGIO05/XHm8
2zgao77IniQ9S4lZsOWgPO8bo7r8VFBEc8wgl0Knj735XBmJiGS8MMJKzrD47OZ+
Iq7oVFU/y1VWuz+qD+24rNImTIKBOIdqOWgszWuc4ZRYaVtbmP8WXvVcP2bgi4Tp
Z+4snju6WEbrYgI3yuLBdiDoOciWoHSEZfa3CoT/S0OVK8/nb8nuZCBaGx9MXKlj
Qie6HQhxbkgoto6GwNs2HMqDfI3Tt5GcftfEIify5JI4mZfrB6y1htTBl/SKm6zn
mOxkzxVwJx5YsRYECQH8dyyC3f/pMTPbDj6jvTs/C8x/62zcOkU6SZNS7gAmgt11
R8EqZgbt4vp/vYSH9yEQTOomOTYXDCNaOQAW3BbFNnJIKLKqYqWrcxwGTw28Kwc8
7I5/dp+AHYiMPijMblBuyrGSXQGxHYzvb5OENbLmvo1HzGQGKTTDN45v7Pb+N8fM
5ZyjAf0lbJ5pFdjeQvcpBLgz45GIzFawZ/Xgdfc2iUDhZcX5kVWZeC05CWY+iAlu
i5wQlMJH+rxXzQZ8AJBx5Nde7w+bGb7dv0lRFw2JpD1rooCpPJ7Cs5JeGLRucij3
TUwA5aO/JgaZouyzuqV61mKJfjFH6fZ08YVI0+j0aIUOqM0hqNutkB3kM6HiJ8I8
GN0ZTPVb3a0wX7Z6IMbw51sj8IeV+AGD1WYIMK1JUcFPSjs1lX+zNr4ur2xVgBJi
VtZg017f6C/NsPrWf0tZYGZcVjFJruIl87UECyr71sLyiIds/trTG6xf3YZYwa17
mhxtl61LX/N9XBtN3xBYuWkR0iaIN2hQO8myBSQb5qZiDaqYUQqiGa36XZLQ855T
dVQ2G1xaCLhGwGon9P05YNv9OzscRis2YLOp7Xis+AiPg23/Iuk5+nOgyYll1gk5
W2U1CcksYo1qaWdy1Ct/CkjAKZc6yfH/n6ziPAMSzobArWJS55kZyUjoSspP70OQ
5ZSOffoeuF/7f/mnAaPTfEy/WGgZ697ExepmTYZTaui42waTSekH/sI+4DThdXKi
TnlHizyZXOrc16u7z6byzMsze0z6YU2oviKAOjfHYBp4Sqrr5k/Do/bMJ1IByOh1
4wl1KnSodbkiJPC4FGbaGpEUuUNbG7XypGCkC8GWLSQquO6vRCahDce9nrqivAdM
sDMOzcHInzd+nmhZJmSkCTRhjINjWKCSFrwKdfBD6H1429Y9XyfyDXvIcPXjoo/t
cuTE6QfhdUZK3iq6r/BzkEMI2zAc/2USUMLc/igwRETCbsGbOG410k30RZage3MA
uCOw6WDjJJ2IxEcRVMxuxhFGkKucbuqeycHP7TGgu7f8abvngz1lG4sDcU4G4gQL
7XJX+gIid2eZjhstPhyXCiF3GumGd5xye9G3ET/6Q2LkXqV77NB3NXtpDX9jcGJS
I7VLQEMOeUN5FqXeweuFqs3NnEaDPT7e8SLRNQgFbKY+GFpA1+ByB3taBfGBx5X6
zFXRhwiNQI0rW31DpsMZcoBszk07XMz1kyOgSs2/YGj4J7v1JHXx4uMHHYwZxd/x
SB48LLbsJr2ht8ialhL8Q1Gf/Ee2kjqicrKqPG9Etd/dBEh4X53lEt6zg9BY7Mee
I1YRZ9QOeHUqj1IWiXPUkm9HK5bCbFunkjaUH0yw84OZgsxkEc9vHpEZ1Um+/cEd
cXzAnGgsIihPCVSf7/QusxDcqO9SPKd+Bq/yF3pGJUHd70luOy/yRRl7cicth8qE
xIYAChaXbmklbgubioJTZfY1SbcvbgEdUFu4iHNvqE4ZEWPyqJUKoZdodc9eGY7x
VWY036s637xPsoFeqD1nZBjTbuWbC8v7wuSQgoUEPNZCqyIgDD7x4i1Ev04x33xZ
5fzPq850I6emxBbYwkTFFSj8UXfuUTgerPY7NqLtX8NSAwmOztcVdsTwTfVymVFn
YcsreT6JGj5wM6+9F8YlajHVIwdfkfRDgwZeu0xIXsL1pZr4JRxVGR/vbCuM+RtZ
7UYoudBj8nQ09snVVaX3J5FxVSeMwEkxjc7scf1jfdmxgfYSuIIptk2DeC6Yu5OQ
W80Hf/Z0qgpKT1pJFJXD/K/e23yDCKEV8P/ylURKHqpieXdWsATjERjST+C1RwP2
s/ciM5uxxWBxKWFCSdVlQeK70ITnJrUynM79EaQ0oNFUeEaCaUqVRMChR9ty5Kdd
EDlNjASGEbKcBRyJjabMIXjhvdJTfO1VO2T59jn6YQd2geZ1hMU2vECFtyeKLpF3
u/0k73Ldg3QybS8eiPdmGuvaLY0Q9vFr0HycRezZuDKwLgWW+ZZZGA+IvZBVtF8Y
HpVj1FysAG/Ke4i982ryFE7TnB4CYxfVY9bUKuYS2901cdes0lRl/NBG74mxW2lj
25l4B40R4WwmPlXeCngUBbgK0XnA/pEpgOhGkk9Sqr7vx7AbRmmm4Rjo7scv813Z
FRkbVis+BuEUmDvVg9knq9YVRq4Ydso+R/N29cR/SRXtmPr0Laan4qASrW4wN71R
iWp3EBbaTNtZw60PGyoYqiZKsm03yMVcCVrXAbcFjgLBJH/Nu+9BOgkScPoxenID
m4gPCkDJOAmX5Sya7zpros0GNwMBRLpUdX0sh5zc/EFGq88gaEmvXQopnzLM9Bbm
Gsal2kFJZ/WvqL4hmZw7lEKByKnim1rpNUeme2z42zuaW7dx3FRsd5+ooHAcW6hc
D0kPIzDzWexeUcaKgbzgeEC5oqTGWE5heML9ChVcvnpXKtzkniFdo+wMvloLUtQX
poP0lHuc8UY/WQSN5iwUBBNJ7MzcvPdjIu7sLT5koQYNohgf/kPH1WIl5ABKFl2l
1h+XJ5KCFcnzh6P1sJSK7M0NixD4UfoYM74Idob0bKoCuqEehT6yC0MxXcUsoP4U
Zg8FhMu4ZJccOuI5s7URsXGcvZkE9LBvSm/h6QCaIVD4B7MWyfeSI+8U6oNSv+uV
V87le+ote+JyllPpoCgrVm/XCbiC4Hh+AfqHs477e3d9p4GltMTQbiF/uc9SVl4+
K7oxxLUTW4+29UASapAB0NikV9Ja29RYwfLPKnxuJH/3/rfU2CRhE6sZU/+pPVGU
V+/qP9E97wx9UZT1XzNt8f6medrPPayng6xXmz+6gEMcoV0gWStQglDCj4+7TpcQ
b8NSExYYX+Ou71GNgFi7vxRrSD4Ljj2EE9eMoiAG47BPZaGkdEt7oIaqGqSEskgg
LG4bNxCfJooo4nGCusNIqXZ4P1QedjXHchYQG5MedunUh6BXZyYlxVzozqY46GuA
vFwriv0kao8SOaFomwQEzYpajn0Tu5o5Ghzl6sr81zVjS7za9dhgWiusFYk4rFxC
Jha3QRXk9JnpBhjEL0mmFijIyxSmBk2M5G36PDiMReMbqEdnJBzXuNTAjVTJtOtK
q/c8/Hf0n0V6JtHlEYfVkcqapQut88dBiW1wv+FGdhJqJUlTo5c8c0RaD50zuPpY
vVHdkcT0jLRe4vNcOibks1UaBNgM9QyGuDb3kg1ndLUqBytG1CSvOubj2Z8WfeWh
241OU/Ei/LsrrkwFVziKVTjmpjb8iP3D4n74r6WOLDi5auwEej1v9e+YrCEutUvN
Hod13fXbsDww67tGQk8c47ySgilkHZcw6v3dG8bBLbW9AIeM997o4YytiHcBVSvD
g0SZxDqJk/+twJhLMJMHQ8wkXRpD9trJ3ASRUnVpsRmLrFeYMAFn1lBoTpaOl8nh
CzA8vldkcaA+kN1vYQDbu3M+CxSQhpQnFkO0zAyBxabcJnO0IpC5gAenN3XU4xJJ
Uca+b3Nk1q6FuzjcjrzL3w7FObaDXCVAprervO+K7dRduhHF3sPh31L8r3kVFgnj
HgnHodaq4cC+WOn4fVkZuEkExilC4yiWO3anNNgWLsNEMY+3yq4APy8QV9W+oWZg
B27ZXBsAxiUYk3QzZIwIe4Sbc8ZvtNBQ0NKaK+bNJTHg0n7uXm/+wOkncvFMjE2i
gWr5edCFRpSOCX8V1FLu/41TCMfq3FANbK66TvjTDxs60vvMpnmRg5aQKgCZmbEM
ESqwIQsXL24chshDgNfCt3Zd/J2UJFRX9uo1ropKzpCKRV6vJFhf6DUUwMQ7rZZG
Ri1VvIoTyZkuseM+JjgripfwMAe2T40XihvFeUhhZ70UHPXWSzR1wdGkn2LE4k5a
zyt9gwJYmzkVYNtITmc4fT/v4rRQnUT8n/tiukVXEsdo+B0HeT0CIjQ9GN8C4Fa8
FU+HwiawvQHCuFuq99MsrE+43GZOYFSRUcpcCBaz+qAfTpxITUuIUVvnNOlVDVop
Sj+/s/RzEEBybY5yukrkaU5YjI5ZdIji2zA08sCgcvDww4gpgNO+G4zzQqe0Gh/U
RdmZVuufHk50Z4w29OHfl2Zb7ulfdP192WTOui1/uNfyUWTddiTPprWT2AKi7f6/
xNhgc2sd32h/rajCTNwbicV+nfmrVQCZgAni/dJ0LYMpnP/7nChwoyWiuPuLOn/h
7hP1rCjTtqQuiF6ohaZvGBHb8YosnyMnNv8eXk5Rpb39V8Ndxrm4Ec0cL1Rd3tqW
tePpCfXdUIHaFJNhPtg7ImfmdDtfVJnCA2K8vinF4uJGBb22Q/5YzzD1R8TLXjTv
KsR2DTfIFsJ1EWjF+DiuNFVPa+jKaXsyjMZdLcf72LIxxWfueyb7rfFERYROj4q/
iRtaze1jpGSIA7x6GttTHeDBiuH0tyinQZZyaNj+wknHZNFSpDhE0cwz8OezegRJ
svh8M2q+sttqkz9uQus++Z/wKT7rsCBy25QBkCY2MjSbifYD/pq5BqIJgeUp+N9J
wkRYGYk8YBwqLS9MN70uFn+FoNTUPk10eSo0Yjqxs4SfUuv0RVoVzGFAO8Lc0gIU
8MhfxXi7rcfp/thvbHKEIHjegV+Ezip4ixlEzG9MWphm1TfNyYfumqrxc1Ki9TdJ
qWU4x5cC1MrrLzjZq7S7FGBAhRCLoVryScvsSuBCC17YwXE8EYC3m8AhFh+cr5w3
E9T4lfFzBtuX7ks8Ifo6xN8g9d/3TtMCHL0pjpxhSKedj2NAIGPDWeQfFrx0Tt+i
U/OZqcj3oFd4I5HxYCspjgCVGAZ7LZ5qzrPYebE4cDv23shVyj8/tgjcBLGUfIGR
nal7psLm5CJtOEPLno4q3Abo8Wbwlb4Z9X0qBvJ8rxyvLSL0G2ql1MTFjgL3POmg
lwKWH6RmC6inVUWSAFp8KtETfJ5br5JbUDha22HBuT9UX1dXThFmObEGMiBbg+/8
upgA3BJe4l1C7truymhcE2BQ8M/CZA2JPoM98pi675Ce8xn0hz5bWlP413zfP9H3
M10DUKqkALKTsuww5wKzI2G9tIMlC1IOp5x8tYt2pZg5GnqEbL8WZ6sXlLkPFP2V
AwMeGZB+VKGPKn22jg15xDQmLjpccmRQ4v5Hoby99vXSx5ElabrkR3oJf/gAiXHD
L/FfxobY3cwcV/3EL3yxR/Zc9oFVn7pjrzubBa/p2zfNKX2XbCIHaKmdBeZ5PKWt
KyirKJM2aSB9jzsZTD5r/s1m9LgwO7yNT1OlrjrnH7VsdqJyCAMUWMlloqn+4/Hq
fteM+gUHwZLWSmousTQg2NswO7lwzhKZigFvuP3uW1U7UhfhUPU6LyG2PQSDg7eX
SLGUX3vBo3yz+p/rz5g5ruHrK9CRfjLQBTtC6Y4JQoaXy10ofuJYRE2+QWq0xe/p
KpLQoyIeHfL88CCrrOMUSQr7xVAC8LrHnsd62/CQgT5r3VUevo3pUhFGuph3C826
oYU8x98VVIbG2Hyfb5Vy69Wqf2rq3r8FYkvmKjurWa2nhRoWxcjW5S62rwTGEdGl
IX4ytvEpMaJLSDLR+eU4kbvI2Z61o0e1z+G601NBJmgCBFxJdVGVkrBQORvLalWm
4QkW4+HLOx3XQ4YTxVpPVjg5j53G+9KMXQZD6/m5nxKB4Fw/4Q5KUvfQF3xetJvb
mG844nGizTvqEJ2A6H2b5Hybn8EA1KLPk9LzylF37y5oWI/bD3zqSg1+yRjWC4mX
hCmkHclVimJm0T8NzcbQma2Msqk+JVQV4KHe4Uy5+Iy+2UcyiWdZYQvHgYOZVb4L
8WFrApSUiXJAOTEmMbRb+EfNRwCL9Gh5LjK9udEILIFHdByVmntgbzxd/TCEX4fL
3kHkcKPjBtyIqSenbQzk9T+G8I0Ear+vvKIPlflH7Uv7EY6OPysQ2i2STCV2KR5W
pkSwsXwSaIxWyZ/isgQ1Qb4YgmQy+KjQp/VpXOM/UBerEVgKi6ZdXSKZU+Bq/I/K
ctj5P/OMiNGGtzb9OQaqPeGsVRJLWKBBM7/IL+gkNuVx/90QWSkNpXzjiOL9AFqu
viYLlvQBeSN9y0pRti438dN4KLleQY3DxzkUyDLwVJLHJrreJ+Er4Zsl3tZ0mRWY
cbvkuikrPERkExz0kPczovcBb00vt6TlzsLJhjCGCdPxlKMzImCntb9OP26+G7/p
9DUAe/GQYLtbegGhYh2p0/PQ0GcwtCLRkpBzweKh5Pqi6qKa2N9ad8mXmIxQs1AD
vovbtKioQDHn7LjmnY5Wok/zz720Ui0dcnPENr08oGXt/CkLYyXs8rPYHkm+KGiT
i6tUaOKpTqvkmdyVFeh5T++0IxM28fHUWUOQigRxXxiFOAGfxRHFcbnoZ1s2p4Gw
KE/Pyn/2WGgzg45YIDsRMe455Fp67tj3MfKsqPmcdoOHW3nxRq/mloNHnUOl/X6o
7Gwurl8fJYUkwfzS9FftC+QssLndWG1hvm8S23tBRn47nN2C6fm9FRULll1vV5pS
j3jSH8s7mK8PzL3jYF420wHPo2nlrS1MpcQtfA3JuekiZh1fxahateIBDxRig/Mw
F3rKAr4rv3DBnTWjTnpgyeI9F8DorgnVZUOnN8/ZiIOpDdpTLt5dGfMltaypclwS
+av/0m09K9gGp3UGUaaLEVycroXNetiwnUeO3t+KY7/XIxty9LWUpqJ3XF6qdwdm
i1nIKv6wOo1uBDh3clmCV0ZQGv68V+nS+U4TixecNZYtXhmKJeBMlfozglHcFOfJ
eCmZTkPs0+RB+vlAqYTJaSbiHPEz7kFNaEfAF6kfmgjFGHQoYlhtDvN5o/3AhiAY
LO+UnZPvUnrg1RTdghfPHhbCA7zEY/+bx1VRPJ4gc3rIIyccqlL/3WT2WmP7xoJT
JryUN6vBf0BeDpb3rOH0i5CEPxMNlcE2s574JzADbEXfPUjewZmPJ+2gLQDPdg7I
pRsUaeGSFbfEtwFywAEvI5S2yKG6cfdyTe1opkoxWJWhKOUmC+ZqIfFcDcEZmvt/
MZQgEbaztRlIWoSnKGrV3J4zwSmiHV8akVAR027oIeFYekpWMJG+JQ65qdrAMb0X
DY2ji5M9KQHzb9jttoVLFbrXHpL7PBCRXNEaw80avv/BxVuHsBqkR2zFsS46K1W+
72Ckv5CIdVHSx+71cJFUJMsuZLQUc5kW4QguHNxRDeuj0Rrl+uxz8gXb3IWjuTwe
fBu6+XuHPhA/hCB4BeLDYGasgff+vUwKaObTnpPc6ywkru+979J4zuUBZKc+KuLG
Kdc0zp/4xA9GcOrj75QygE40uilbSal8vdi9pOzQ2W1F64bmmWLpkzvWXlGItW4M
08W4mmbTdHdsYXTQr/srd04cVoKCM5sljBjNmAyuXPa9RjNtAs0XHuP9reMJRz19
QDL/BlQbauwsh9IPIrc5qWf2CY63mCvEmPW7uYWROvo4XmAl/SPuWyuqs7bfHs2/
2K5LnqLH2GOtUrbCdkDOcy7bjRz8Y+7KQq5UeHLS0hoPTnVx5XseDsDJqjW2g4ZL
Zw00XzlUkrYOWgu+H+Bqs+11TlsMSegBsL6RpRkPWNDOSk2HSiGB6zEXiB/CUHl+
S6WBMY1k8Vp1J0CV3orVk152eGVJWujEV4I6oyECXPxqfmCLGTrewlRDu4egqthV
6nEW2m/J2+3aaO2JLhEmcY8DYLxFkLuIHeOglZm+6UeYDKW5oNZYU9Cz4fApf6Du
7rMq6Zmz/g3l5vYKcPEoA9PjXf7HEVIuv7KM8j4UV0bgAYUK5hyS6kvKtV+qjlgA
ssMHCE9JCc1mrVVKgGNNc1Lg4xo9Oo7XsohX8L9A11hh5LfpcgETkOo7fdtz0OCS
YqPzvEtTN3NF6oQ2EGY83syWhRdqEv2QJMHNnZ7axZdFMYtrB4jhU7pTO27m11fu
QMEeuiBci/3No8MzCprKDIhQYQobgz+yjZJP/UYJcvuzj6l1RZVO0Rw/TRm19/5O
0KsZPwhke2QDY4G2/5q67kkAQsGofEWepl0rBxkV9uCkXniCSJ20Uk/50JK7rm8r
pbG64CCsV+jiN3wLeXwnxI1vj/mwhXVFWAgP0j8DvgH/tV7isZvWeFbSz2bdvors
TevCHD/o7kH9sN9GRvDng/icYi5CNZkgJaP89cOsvg7jlIe5P3VYMPIGUdSvyv0J
gjSXEzG2BiJ0BPXaXCsCFRn6UAIxqLpvpklzLlJmMuEl5C0+U7cYTFLGv8mZ5ltt
eS3D2fkX1DS79pej3V5FUMLFdujnx9Igq/eeLRYN8dvP/kDDVR7b1TFnfEcZVxVf
Q86I9qu9p9OoSsHXKdIXY9D1QfL3a7znq81aHO0Nt8prqOL1wolOxMQR9GBRWRDq
2O9SCkwHcR02J2UHqaOI/6Yw0zqEEDx9sigjfwFm6G1MYKaMMc8no1Ija8vD7tXF
uq9NfSk4YbKPFTsg1s1aBEkgXRY655ryensV4x7aiI66Ij000NQD/bX3ev+1PIKY
OsxWl7W3pDYwU5zT/6MKT1roTYLQdQ5yRIxjJZBrU5WxsIYpoEX06KPL5tO+sdjt
7Nf3mLuHdINpFRSBo+hWGg056B53dQheK7RW1AN7d/xHiD+33JTRenvCKtDpiChV
0QD4q8tOdp6xN66NmYPQ//pknPunKa9pJSevUouFixZe2l5Ui/lsxP+pKGjvqdAa
QONdCV5KeQsUzT6ihUVmQUDmFovRWeFokQ0dDAonAnZHeCOcqLSxri0jOPABbltZ
xsYV6s45zsNpOoo3XsSIYAg1cDB4g42FQlwJQ+TowuTF7l3NzD2TdjCqJL1pZ8Ct
GxJtIdQHEyUglb7foNRa5n0S+g//Ag+4eBu4v5wojLUY7P2Y1z0IMXXeH2mEUlb1
TeOpm5tSnU3EUvRiMS7KEdL5+IXhmGm+AB1DEFyoCQF5CDOQUgzyvxTFNVHW52K0
SdIzRtLiZZRyk2NRcmm5sw3b6nS26RJeUQsWtlUEUttjmtOO9WPsmLZMcm5bQwfh
AJVGP25v+WE0mImxkrn+ZDNSUA7A1lKSaFmptEhGIXpXWWaPiWRhIKaKyXK9/9JA
NBuyHPwALMOtiZqawNm+Rrib7CFYd617yalNWd2PQoB49dRWajVvp65AawyN1sje
SiC2XIARd7KzT3Eslwa6J0cBAf5stFcFVBhha6gZutHaK111VPhP9kI0n9yZpC8p
3QA7SGJ5zvntghHRn4mmtDNh3keiFc5eRodrZasJmtR9VsgOl1vIZ70fW2uXBm7V
gleYVFxTHQyCdYOzP1pDGOjwf0XhzpVQPibLyNt/yRa1NgdZ3GRAJZmvSscVyq7F
HkmFRszXEW9wR2rC7ZFkS0ZPBO/c5krqqRzQ1gBvcbLV62SwSG9MFExMHM4aAikL
G5AR0BLItNzJDIMYxnzCiJdxEFooH8N6EY+8lBoJSit1TZ0qqCB9FVwaDZ1Xh9em
8fWTO2Wuzc4g26GV1LPk0ritlxCz0tpR4TvRjpMxR1k7SAaH9VCYg5QRuCz44kJ/
9/koIjLmIlpOrlTCxBFvoFudjRehOPgM4gga2Y5GSZuYC4hfO06CEoIt9xgrGwid
mpL5o6HqDvYe4SRtgdyrrG/YBQulLyrxy/BxoKPjRYikTwwCuYJqXcUjAJTANljr
7smCpUdffyCZFcp33U5rO1vFRp45/9xO4BbeFpYaUFTxi8j3jMmMkB8DSWrPrxIJ
woD9DVCwL07BWo8fo10H2Efdo3Ve6szHYw86/P3h3BQAS3BWAmGZcaFdiDqyj8K7
JRenk4NFr+l1Cno1qMCFCPECSMy7a4qEtRhbMCwkDxmVD+BnGqZEz5zRdX5vzUSh
b9swG9J24nOK1ruLLHKCdw0/zDdmvPam93gVh7rXzby5265OKHw9dxi/cjqs63eg
PDPThlc1Dsd9CqNlLUc2/VtJazL5wO6T9bLfIWrGOTVUNAFol7tKW12Lmh/vPdGb
ha9aSh59Do22NKvDpbaUiPdxbRl8fFGGkXLcfXXmRhPspH0z37xvU2h+3A9FhV7f
u6odAGn3gXAw/KHNPLTvLOLmRDILpmjCG12tpncv9D5ZJsku6u7qjryQzYyfGYX4
7+JZRVy5PxuRYnokq5KBTz62xN7fgNqxDkhU3Iz1VLTvSakD+so7wa1Nf6EhG/TW
68NeMcV29nZrto22KKUBtBifIGpUSGym9xcy+7LD5WOYdomSXtQSf4jHnWbdMrOf
jd23CqERTB61voFQ8J8HGv1DhLGr9RlGP4TdylSwgTjcaJWPpcmsRxtGoZ+WrNR4
MFDF6TY/BZppm9c0qCjvFp4vFE188J5LKmf79tyTemODCwgkakb6x6CEo38e16hU
EJVz9Dth4D4WbVRzqa+mrBxNmPw3dPRP23nWgpWm5oJH58HDFm7s2h6jIDnfxyL+
P9Dh+DEIRIWWzucps0SgZfKP/ZQLvpCBSdHc98X9z3L9T8sDzwch49CS4tg1GpBW
3RDJs5KibB62tOC3H7OHE4Kb+6kKNPWpr2tflH1A0/nWFrilWrlhGyy19cpYoXhF
ymWEugx+6BM/DXiwDlMr58iL3de9rCr4JO0s4cGlNdnmtTHSZMPE3dVW87lz3A9e
fwwNhZLEZrk88OEoEwmaZbPAUQF9Aov75/PzMCKtjy7HaTwhPwbVmnrY7A7guRDU
we7CRWbmIj08y75hLO4pvPtCPBfzow2Tq1MRb82xJy13FMaah4eemjMPagGetnVF
qh+SHtSb6NquQ0BZxLONcdKpqIEatGDDLeKY2Y38u4QetZGoEhpQEI/fjpfitzO9
DC1x/WuucQpc8Va4omBTAS7PJDkYiZuSblsbFLd9O9yQAer4ooK2T4cMRnrtWcxL
AkP0CBWmj4dTA7vkOE+DUxZrBPBJtjMgD1KR3vfXBDphGStUHexDDOLsnbDqQ30Q
wsIJPJLh+xjnJmzbCGl9BJSZLSUz3M3kOTJzNyuxBG8wCGwEp4z8E9pMRtd1depJ
8+wOvwM4dgU23E4Fk6533rV1Na2nsTrAZqZjxsmvjbINfqCrFLqPlGWwsB/ws1uC
GpS8V+mVMIS1PDyEk9TuSIUi2wQaXd/mYLZp3G536r+t7fWMUf1SZ6X/7VO2xW36
chtlpI8WCLBcB/48LIGLqGIv3DAQkcKl5Y0cKzsqbEV41zNQEWyjctPpplPf+l1v
cPv/BGnZGaV5eeBTBXr70KGanSUxIzFQRwG6JspKlq0X8w2NwkTq4wmdH+0sTjVc
IbdRnBjavGhJ7YCwn+YYsfM140jfRXqkJrs/DghDl1dulp21Uo0K5UTiXTsmmPFQ
pQTD6mu67M/g7KHkN/GDvR72nTcheEu24X3TUJZTHtY/gGHUrn3sCl2lejxhZNUE
HvGcRMLaUUc4kO9OpK++j3+QVsnxjoPAp5aAaEFqmvI/lTL2tns0S2p0XN50xPdo
tuiLaktpAtVMZ4V76SBVHrSVjArfJClihhQV2VpyHB7lk9VGZ8LoTgGmUzymcYEu
4/TEoIGHDoW/SrYTYPMsZX2aObY9sz2WieRFwbvGPZyCDFBYX5oPG8GnAJq+y9f2
rSNJ160KtS68Pz9ODGA99eLxiJJa6p//qWLfvwFGoEByX4arP2IBwhnHAApj3HiG
DwfuWm5EwGCnmTy7lTF6uZcY+rL8EgP19DE3G7QdFQVY/tmd350qH9zVM8kjgI5h
1jSdKimKXPB3q039mh4fMrWr5Mw9w5vEp9mA18FXDwYdz5kTtHYYkkay/Qz6gBOy
l/jOF5UGuJNvPKe67ckJTVHEn0kKOOI7L94a2yyBSsclzRTmgONee2L97ixgmDQF
eKYoW7N8LGQHNQUghh6ZhIlh1mfvU2yhACM0eo4M0kCMUb6Y46AL0reyL580sC6l
6DMrEBQJexhtNfaZ1SW7YE6vZXpxQd6beftkuUcOEcJY9I5Ki4AWN84ryK7WkW8n
ZqH7nJf4LJNN7E1s0+zlYLtLoWSroesO6K/pSwFpvVlmLTJ6elf55+/TAtz3kiwm
JhANVkmA60VaSChOs9qIVr2S/DdB8tdLZmw5XsWl3B0jRpHURrv9tg5/dD/s0RTS
t0wgaJQvXiF4nzxl/OcMAEC4c9q/TdbDwYhRTvLJTpAH4hja3Z7jJqn9WaoptP/g
buY6J3ZlKMs5YJs1gRWIB+YM+bMPY8kG65qG8aZvxxtpmmx0A1ZlAKizRRy632WP
+Q5rmfBYf1L2HiwHiZRDhi5wWrYQ9XP0xAL8P119Oiq2ehD3xsfnX0SvbqLmZ7fI
P6y2yEbUXhTaGcvrP6kuj12OOQFe/ATD2SOawnTbPY5Txbwp9fOkMOg4Ud3H9O+M
AelyMkByaR40/Vq10gqyRPp3NHBH17QIgjNFPcKJ6345OyaQUZqpQ2FNs2sXFn22
yAppEOHZCW3Ls7t3tt8I4zTB6luTGFIuxjXnacU1UfUW+inGZ+Z/dwVkGAdgMxZc
vZQk0zUfyUKf8FEcpd/C0CEVNrLB+jzbZFuJ9xuFyk6lkx1wD0Ai8DEg0Xo2iiU8
31BHQPluK9xBgRPdyY8KqjSR8YsQZbvL5xBu4p7K9HhguKG2iod+to43TDf+BR4b
wJcw1JHn19GZmlmxVHF8Q0qFQ+PP6qOA58Ota+BWKoma6AV3aMafATcWGVEDBfIT
QH+dTuer302JcIFP5VyAszxZ7vm+cCmq7vXSjRhXeXvq9EiavSAZC52ciIux0M1v
sCAx3KBkKY3ITpQXn00+aHjRPwGyneOi7yq2lqqnWDuF3ghlEFY1GC5lMCLXb50g
kI9Yj2vHkd/uv2mgg8PDME1XkTLppSJH0iVevEOBdEecFbcS13MQm4SQWJtCs5DG
sdJ1cXu1OqvcZu9iajZWiA8P3j3UpLK5wenvYCZ0g2p4wrZYM1MVlzom7NEJ4Ogy
4yp4ZyXU/pzgmADfgj0CuxY4AxhJUi2n1wGm3ZbqN+TNk0rQwN3XvX4+hMjEShTD
AZBBDQto2ZeqNR21grXSROqDbh/MGLWTpX7AHoKXzT8p9u9UB5YBJgsbzT3QpS3I
PH87wRXmDPK7RY115lRiqvh2RgH3Ef9rJaq6qShw0PXiMxcvkcxpG5ml4g1uOTpJ
kE+wHEHg94Z1D5kg6ZmMVTCzsebnMymXlX2dVJbVtLLSX9t7Z5UCrIwHeQf4Gcjf
BQ9i63OWvTcLJ+goou7QN4l5TSNpWTYXjY5GBEVciDMWXkPGvIBGwSQso6aoeYcs
RSEHmg8tlYLLHtk3QRghXQzp+BWHluCp0pRk6iR5TCWQM4fT+b91z/pJ1YC9P4ui
FBx/CSasr4XvUZrEW4wZTys8/NDR2mvXgP/2ytdVRq0Ud4XvdkKt4V2xZsK+Fzu/
Kx9ebgaSiW2CmwXFgZhbf8Zso66rfwl/OB395q+7G5P11CQRN+uxNbqKmec6MLa4
CZ3FrmBzLcWKgLXVoRTiWWaA8rCyuFMCJZHAQo2Wa6nj4CwxDudPH4ygtxckmRM8
r0ztvdejkeFgf/5xlgBBp70K2wOcV6Owac6NKNj7RMGZpXrgRM2bJsmlRyy1JTdh
dg++enrI6N2oDx6T238mONs5I4ief2UYGgM2OKSuBamvQ5R/sonC1Cy5oG3zA0L+
aAVN5fn6y2BbhBSdHhxE1RfGeiEFoPG8zEcH0cDWiFyXKB98Ely2a0rg6oJKdQMg
PjvAcAdVT7VMVk9DA24OoP8JCnLSdJ2fc+eqvyAiR4fU6s29+m4Lt8I6BsZse6Jr
ZtMbQTH5TPEeBzd7K1XlvyhjGYz+7xq8p4oUIxp7R37YQlVumpGmbnXi8Y8+roQK
Lrl6WaNsCqJUiPifeEmQ4OIa9Aq6/SkwrJIeSIglDHcO8A5s+4qBCMaVcvc1wwL3
4nFTjV6onHi/RNpxeA3hVs0OsmE/n3lJn/UzuWBEMVofy1RMHfMry0ctbqp+W7e8
lAZ3IXtiamIu5BU58UQOAeq+lyq5xr+hYg3dASFIEU4OIo+LRxjxqQoL0hw2bfoG
UIrcl1ECv7qbGYbudshSs0ga4Tg5dWsxry44qvwhaCFSOKdsmJAVgdWklczdvgZ/
bQwu97RXdrAnByL2sixUC7TpbVD1vTUd8l6SxbuYekoFmK5FvanyOo2P25S2e2WS
J+RQLl7rtyHGp4EsMSZxsqPi+S+MprI3yyfrWMqdptG13B+HCleMm4gyaoEX5bWM
tS+gYkRoBTZC3s0aAUOV7rhYFlA8sZoFE91VPI3XCZn4jcc5YyoCS2a/72QI4Vju
qvvKY2J0ShWNsYvQ+83nbFWup4MVFiA5Y9RrBtCQ/XHRXqySP3wT0qwl21VMIbuI
Hn64aECEQta9GXtB0xagJxQ+WKSR05KJ6eKO4clfbgIp9JMjE25ZQsIrJOSXPzVx
UNtGONsiJNmh7H+oqGZt5MonH2DcHJjtm34F7gi8UugBsj3bvU+5RWSQnTVCDGOP
0B4PV6vX0MmyWt6M24CCtSli8F1p/oUHwBmROXkvOnPqQ89BZTjY2cxLGRbtpBkg
MxI4C02ZxJRmpwuho2vGaTtD/ICuYy8DhHyL4JzmVpQU8zG8p6llfL5vGn2+8Uft
jdB/x0zjVVMDASBfpshpqedpcDurnrGUWHnoBRjhBLSqc0ricjtHA+AVEwGoQWFQ
xGzQADn4s/jZ8tbeGyNaGkG3cXyqVJsPRkI0AgQT6GMT8se8MUzjpSa0j6HTTppj
E25vaPyu5ZPrvDM08mV70h1ry7/03omRNOkMa1eC/18IIlMw3x5v8NVIQ71WjKlk
taxYt3DC8nwLSarytMxnUEEV9QoVfddrFNLupBkUu/MpctN/PqarrTTEbkrO8m0G
9WVIxXKKFerZb9gQvg7jz0J7leb8ojSVnGBaezWzn6OcUu60rga7syDcm75jib2w
ACFafCOmQ9bmUKWs5m5dKSMnefLZwOv0l4FJjOXmx3HL2hXFpWI34+xIV+VJe0Re
VOahSPYHp7+1dHoksEQxZlnVZ/c99FhnK1X1ZrislS36ojBrgVxbRWWaeNLjZJNq
85B9HZcVLB9I/0cv7DNNNGKhBzaF6wf8eayVB2eIwP9lgAhJgZ+dSAH6qKo9+rsW
WCJRSELrlJNbc+EYwACLik8qX1+kVB1vvD6H3AOwfz8lLpZpxWEST8gy0HEwO+C2
H+YqJ+Rkr6pmJWZQEcbGaIgGUq3dtVsDdczWMuwzh5ieo3PWqCXiu5WIc8xQ4yAn
oghTnfm4xiGAoynRA/UFgGoF7bYn3FQgqp0PyuUr2leD5pv53+P2NLPOWiFPny4G
E9bo0kwTXHZPsARoYc2C0sA/XJU/DZLmQojg47Oo9kCb5GbKH7ibz8BgyQAenoZz
lTgH8F/YRiPJ4FLjw8shfN4O1KNGCriTNmJzE9hCuqVtH5e8f/wDqhcMh4wwOfCY
XJsXOYc6hxmmXMKNx2Ue8LUjLhBROV+QvsGLw0vpbaMoG5JNZiuuS/IYQVic/NTv
0a16uIzSoogcgKOo28m9XqH7gdX0YLmdTMlN4wRrj17tuwVYEWyL/QtQX3vG6iLX
r3spwYP3+W1JbYl34SzptVP6S1ivaQ9xAnBkvPezG9ykgXS7JlT2DlqmYDjp47iy
Ch59jDNJRp2HdYb21F+Kj8JiZ2NHtBHvrRvypO5uV3or8iAQqK9OS0DlpwwhM810
UnHrWBJZqT+yd/1eosJBSO5yguuRoW6OHoq5wE+kCYi8o1js9PUTXwaEj2blLB7r
244OQ9Q52iYR6WHa3EzJvfqIl2ScndAsZZqlgeUJbUvEsHuc72m4IXpLhJfKjVs/
O/HgoBRqkS9O1kMR45Kn6v3JJEv65GGZyoe4Fb0/UGGfyDJd0NjDZfWEIB+FK2yK
5fDWv69ro0/Fj+T/7QF3OOcwRi5qJZ05uJN8megZTaod2TW5J8AjVPztm4gphaMF
UWFU0xMtIDj/mt57SvjeSZOrVdd6aQh3SCLIHNEv2DVlakH7p5TKajpcKSYiSBqa
+IirFfw2RVwhKJRpmVwf549nRDxa1vITwEhItPac2E46eE+P/8Rsqda8lnPXPg9z
NVQ+bD6GybHki2r0dVpQv7ShHCY/iGD2Itec/0Rt7y3yYEZ5NR1i4L67TNlAnw/4
MqLtspfL0Lr0trkG6PXMjt6Pn2QZipwqfiz22q8a5EynlWiM3/T2yO+Daa344Q29
VVCz66tmLUlzCiU99Y/YmPw0DxsMwd+s0ikT6itSKNSqEiCHC6B3/bEsm6j1gNm4
R6UGK3szAeUrc/pNLgHmFVNI2BNcJQF9Zk2DfdxPd/EJ/+nP6RA0sLFg7wBcNh7+
++e8QksbCK7QlRH+PjsMywtsg0PFWQaC3nT92PHwcULJKGMUu4ew2kqB7EWOYIuS
R7k7UxjG1uHw4h269LN+pEwYCbxKWeUmscKGkqGvVsrokGAnNUio6sKgZmQCgHOu
PxUBd8dMdJD72HtZ6WeQ/cGnCaYs3qYxW3OfoY1Ct/6Ei3bM5B1zCHVO8Xem8zjq
SZ8M81uEC0n/Lo65LfEjHjdx5PTR6TZxdPjL0yGRUjrWgLA/T83gWdH/g/09IC96
ymCfRcYTP1bA3eQDnus1evwoBFxuuuXRekmmvSQ0At2+7FbAl/mYCZdzfsqu/La1
AMBPn61Ap4ZsO4qKUBbY6aF6SLXY+zGDVOptis/3guy/surx2la/c4oKLfku/bUI
mBo3sFy5a/AL779lXeEKBSY56qyFo7fscdA0WIW6PMoiBy5NMtoU38mJvMsLdASy
u4aBDniRMSWgL49+km4DMHpXf04nt23mL21D1XF0IPbDm+YFyugYGg8SwoiOKvZi
9WQDF16PlNNrvIycun54g7Dj9s3aMe57GYkwdu7mQAtwrCrNx31aQpKfIN5P8G43
+73r4TKJDEJSOmJyNfu+3SUmXjsYlZKpnvdKqm9RWYYic82G/dkzfDHUOMIKOBDz
qKJzCnVlGSVOMp5dguuj8j5P8HWh72OjvcJdagGEmP+CUma3MB4GEA/SCRVgp4Jl
5ZLj1HY4K9ibUhG6jgHAKczot95StRwbLVUHyc3aLeBhlXq87D5N0LiO910dkwbs
sTy9vzGLXqKo94oShLdmKhY5wg1TdVhXsHPnhPRXjlMFo6a6i/5YevWV0J8kxOWL
+U5iOXqacg6TyNVdtIvtYkx5fY3YOYnVBuMe+zn9lZbxxzVh/9xD3doa3+Pv6+no
0u7YX6QlEaLFDAcTzbrdhT9R71Kco3DmLOt46kq2GURvCr11yHp4Im3TvBQwEQ0d
iv8tvu0MFpiLC58OOVYo7tkaJCF653T/mN45bVv9PcRqke7/jsxrdeihdAOjR/yZ
S039kOUfBV78V2yX9fR5XJWbfjrbvMYmXkFkCukjZGyOXTEPL0Toqyo05JVxvxws
H5mjqRy09FUTeQgWvTQQLgNRK6UruWuIcb6wOvZ6PmWHCAX308qXJx9c9HVJlBqC
IyPs5savms/rQVDDPpLpce1r7ba/WtfPt2aku7l4/BNUeVaqQZK1JJjNaLsdqKPL
RxLiMG4UArpwzsQ9N17Az758xIXB6C2SR8w+ILbkMyAlzjaCWMNRFaghYhNesk0c
oIE/L7lUrATdkHzkerMartsD/MiWRoTzS54ubEuy4NsjSAK7i05pcdfyha3djTZX
86pqE5LW+XObGGd3oYHU0Sj6Pf5plwj/UA54JJL4p5s4BCbk1neYBHNXR+5iPGvM
f/9vNNmTSSbH2GzOwAgfGcqlC0gnmz7EoJfWGGlFW1r3D1fv7bAvsWXKGopqe6zZ
KfEuGwA0QV3x6F/CrRe7x+gi89+UhnPqcvryKD0KLODbEbv5fhpwevGlO5QqopcI
N9tK3Tkc2W4cq/tzrN8P8yPNW4bGOFuqRFDLVVYHNPxWYZlTfXSjK9ADdStRDSC3
ZEX+63FvXbkvjWfgLSgJ8Q7+WOwRI8q1wzr2dP1NDDuc1BQh9jWFj4fUB7OETDjt
YghSu0qmGqDg+5XvvW2nCSSNz7sjhsvRjSkFF3v+SeKqEk3yK9E+bgchloUsoJCh
rSlw5Y3mMwmy7YeB8KLviTqYlg25w8WuuFSBNZjWU2na/waVMPq6j9Mn9Vmrxqci
GycVLggMdGtjiQbisSSi5CQuI+BzvAmllLC/rvT/ONEgownfLqZIruhDstz7BpdM
qtGh/nKKUGQOOt17nfSQl0ZgxxN9lC7e8o+5SEHjZf/0yuS1TAcGEhpt63E2fjW1
F5YUieXKtGbgNp6oN0H73dty2Eu30eIVuD2nyot2OLTxZdd48dwvwVcnwiIpqjHM
JiV2ZCEVD22OFO9L6BfLYZNaxxULFq1k6mHflMxdDW+JyiXTCBNbz9ri5+Ly6QVg
dZmgUYguSyqUIiexqT4TlsagovaIjUjTIrjtzRQrx+ztqDDSlfpaSPaEy7aptUPx
ohAqL1RG4m8Xa5kG5G/59AViUV7BZ9ZXzvra00qKg6BKnZi2POIIKvS6LygfsOqy
wGij2IhZHT4QSR6uRRQvJVYfeeqYkm3Ic0dmGL7+hzwzhO4aWPSHLxjKVF8E5Ib0
O2WCJ+0CBd7r7yDzm+BVQd5cdX7DLkR6sInb4ZOmt+CFY/xG5eNz48FqWIX3n3pZ
ZmNU5n72LRAXXBk5mcgHujH0b5j/um3ngNltQH7BSApWUNwgUi3/ETZHwdE5clnD
uDKtHBIZt1ydgzHB9rucaa9JFYyqnuEow3RWDnr9UdwLWqpYJlWIma8KVXnH+eQP
LeAQKQ7ysDE73urgshBguKkaaic2WHYmmoOuJpn/tOrQQpjPu7gUgEYuMMTFtbTo
kWs8EohWSx0iphCyHErV/+K0ES2MPrCwsl5V2h7KQS2OMtm2FpnTryVGLqoAB3uy
p5nQyCAaoOWD2plderI+wwEtwZG4BV3yDt9MpjtUsYCD5ZCrH9b16bN6aF+7XJLW
++k0l0STyiuGxxu4YSzdsUukDyU7R8UMqZstx1MgQnu43wkUkMRUjFnSN8GQauG2
Hx5B8EXmUlTFu00D6K+bLtmtTBZ7tSa12wlpYTFK3znEdfQfwmkFW9pFeb10A8dU
nIKnF320aqKoN0xut5VTe6pu6uKknGi33epHvS46J/0R/GZGxhb+RfviLNGvndyq
Gxgx7fsiVojxpgWlIipcYlS8a6J9vMS+EU56A2+iSam3Z7G0ST8d21Imqmk4PfKg
GtBQdj/8Cspep9KwXdmAmT2CFcN7dBxq5WqM0xDdVkjEYMTz4ARSTCwnjuLcy08g
dMjbwGKohU3qv2fuSu9OMe0oGz8lRceILqMM1qzx5dBmk8FiAoAeQbMWwJIOX/XG
78WBKSZU6AZKakJPRfqLJzWbc/kHDtTZLmjJa/k4wmgBw6Zr+gvdFWPDe4bIYCZh
uluY1SXl4d5VCMxtQxOWHNkueXQB5SuVXIh8If1ZaOaHB1vEvUibfuzm0Sd+yJ7j
70rASGMYXVgwQRG+rpCEHcrAaVhxEDHiQFRQAYBu414cmd1hlXyze860Qal8mg3F
MujhnjsYvN+a024AG7wFvsyO5qtc7Xx93iOYNUvB/f8owXE+i4axZMUDAdHAoZeD
0kNVeXu2yJVpAuqqibcee42e5VDChbJoQ1IK7xHN9JMZ3LCap12308lMvoBzmNdP
sT3lcc8vOtIxdwzSlh40wbzLgoPVdujQi0p0UH6wqe6ldThvtB4dhBfmgFIxB0YL
zSwPsmiDhbG7oqE/jaKLY2R+Ibke2TeQhPsAgP23uQHlu8+NLQ83nmWt/OY+a5bb
EftmdOjMRcOrTRVU5pqZnHnC4qGss2COTVwwSkQrYoGhAQbTOdXRsSCAmDyYW5fh
mIrQOaC1iQY7z1ZlCbBLKKGtZ2ZB1LDk9UGFYGppRldKrksge/vJI02Nv6PFJAgw
3kDYx10hGd3Sx5aGMM0L7yYZvTDxRvDAWgBygITK6JPXP9CS0lOcVPjdovhgPYhW
4nIpOCX3zhogWaK72cn7tPih7yp6+uLrFuDxCfrvKKyZJJfQ8u1gUBLf1IXciZPk
dWAmXdHpXhusGLnRV6dtnzOt51OpVQPmYeBvmvtnoE3EfH0ByBiIS7TPBsruLN7P
QDEvPyWJ1BTYIvKAH1EqD6yl8qph0vuJqtkj9ijoK3ZGX6MvDkRzPWhWxdtEkCQf
ujoi+MXyslBlAt8sg7sQuUAQClDyhAyk13Ju7D+JYlQHO0UFn5X48WzlrqqEGXuM
3s/iKPIdsCjbuE5pKV+Dg1RfO3jL15UlCl0pdHH8XWEFHy9Sp5uaypz7zbDp6jS6
r1/McQFJys3YH1mc3c0gTtV263FzBr6xUvxkk/NH6gTYNTYfvCGZl2mfvGSWxwpC
+RYvbxICTYmpGTz9YUvj61V3lcEfodMrHOv+sbbxEAnozgX09oGqrU6LLHKQ8ZE/
kfhZ2JnBHrCTOFRo5fiNDHmMNYyJkLTMFbRrc2W4LPtRoC8jxUvIGJCgQl4X2nQ+
GdCTvJInWHX80EpJgVEPXqzkoYVC4Zbz2pWlQNxpC+0I7m/s8dVgJujYXRLkWNLl
ZDiohqmPPjEqfzaY8WRYDV5v0l6bWu0TBDHo6OUqDTL8bSRKrSK+VhDeOWcwvREx
wYgQyDEb7LwTRTbvfKm8mb+VvnJlvAtdRSDVwqsErFYqB55YcA6aMf+zd4XOmT8q
Iqp+JCBW0+HYUAcIuBuqvYbN4G1lmXFUoKIU5HwLqdkxmMbaSsrSLpzbk9pzpI65
ygmajn5y8CdTsUVoCK6VGqDKUr9raoi7lxZHFpfKkFeRwkAEIA9rhmvvI2IuHAIU
cFXTNhcurK02R6s+4g3OKK3iy5iaevG2RsVyojms5fVwSo1DxfiTWGDO8M4QZNa1
Z2xnTX2Gduphzx54CPMJx/AgzkO2VdALpJwPYHbbcxjkW3UYlMC+CVk2jFYlNgAa
mSj7Fs5B8yBZykZINd9HBJ2z/eS70C5p9XZDvpG/whlH6eAlAZkDzQhRl3ijRgvQ
GH3R3Wc59R7hmUUibB9dU6oLlgTbnRlz3qS1A9xZhhlIUAHeevdfXCLKmk9wBG7J
a9EeKvM856BxETg+zve0SHXMFfZoxT6eeYm3UV//HQIK68hoGGrW33YUo1uwAOMs
csFVTTW1OTXp8wdprOszuHYMr3EOgkgIkxdhdhX0jEqupV+hz7R6PVW1e+3u1jBX
f3H7Xi6VXk4eUNtazI1CSff1sy4e5uvPLa/gfkkmEx0b+ukAzyHMuBr7zTGGAt8X
Ial7c2XiIbOyZoKamlE+YiWNViUW8kEL/o9MHgJtdGd39ArxTpR54LwJkuHILN7J
d8QuhSR2pPxOmIEBQgclE8/E9uSp52tv9QleAviLYXJpJbpsMkUopOCmc1sCs7wU
LkOp21nkhIqLtjssnnwVXM33+m5R2BB/L0ZelFBIeZX+MrxNUqmpfxZEjCZf34/j
NThMCZMTaQmkoPblbX3Ufu5LDOXWBQ6swADicTcXG1GV5TzGhYset5NubSYSwXdx
aOc3Zf6i7hmRXmrR33ZGEYQ6Y8MZUnIiwvv0nFYnXCLM+/WRj1s0dmCEo/YAlmke
1tdY8Qs3JaHcL2ZxFL9HUq78kbivrbAxnX0U23QV/KFtRryoonmmIlTR/LWsvazt
s5M6fL35LGL+gAuCf+Iw0jC0NdUn9ULBL0nXD2Y0HwaouUKmUolNaIKleUigVm8U
YbEa1x+5Lw7bU+AtzzI/9cEzTloJv/x04BXIumZXuY81JcGD3ZCNM0hdTBJHr/HH
cnCI5qinSxNbyop8f6+uJkD78UzmHTyTSQoH8lfYSW5ahtQT8fBC7A51iTgwUhXa
eOvuXICNQ0QDC+Du35bS9bRcirc70uHbbJT4oDdZgDPSVCYS3jO/3suhjf6xgZtX
vg0oWVyd/QDJ0By9tJUFandOeUwg2bJ8RA3WFedPfL6tr/WMz0fgfzu75Y2OXgws
mWjL+fk+s21UrXpmZiYSGmr+ijsm+LThZr+LJDGTXW6ue4VvIDmXBAHsEAkwZ4Uv
Dtohe5Z2+LvkzyitoQVPmfVZa511cvWv4YjyMrWtj8/Q3p44qW0bSRCoh3R860DD
pvoPoP9c8bAcTb1yznhKAMPYnz5ejOqI2fsySSS2qI22bWaR0at6kAQLakd44ekm
pMHi0GDMOyPHhvL3A0KdDQ0j3lxYTBoKVlh4EqQdQ081ltSaXd/61lu6w6eG7shA
NGmcoiRmvR62DhU6sUFCDugXQTUmmsidohn0kdW7ouhn5gORheRjjPpEvWQI0k+O
HDAAt6HjTA6Coh2TYZnwSWVuv6smtqtPG4OdZMcVa4vhZ1+sPwykMJ5oOLcEJWrN
WWFkP9yNeV6UJmaDKRKLsRw8lZcKJbVKl5WY4vr8Dhub+E2rCykEDXOii1oPqq3R
nX6H0CeCIQVjXaQdG4fCpRA3JYzs2KaRXZFhsRJPrAIcNQz9DGoDI0TSP1v1h1OF
mJf9wW02WnGmp0XkdcWcNwjQbw7Aw342xc84ZD+dRpsCdT0cEzoFPkHbJdPUX4QL
zHGzLpAokMwRCG7EWB8VkqDrH/+jsibYPCpknAECMHnPPe3rvFxzSn/SJWOaow5M
DPVYj99myr+mg2TnuqsIVe6yEr0tWYopGXBtii6Aa4B1h6z3FaRrT1pa83bEtp42
7qCP7E4eD/IwLwBZdGNBC2/ZxFdgvVhQBJTtif78yBIrgA3Ma0UxVskzkt1cz3OF
MFsb0Ez52A8uNPWYvJwPZ3cD+YSk7P7f6gZtkuMzKRlP78hb9l/f61Lvy6ZwlkB6
nvV1bXQAlgYAwbjeW58WH2EJdmwXoNAVaG0YcazOsYq98hTaw5tiNWCwWPvhxNmk
LiuGnEvhaKNMQmxFgK8P51WTu8U5DQYzC1sFVHO6p4QOjyN5rssbyk3R0QEazvoe
bjLM+1kULq+ucj2m5X+Im3YxQ13W9crLMEqW38coP0Y8rIcioOKISzGuuhRA8qCm
aCreU+w8k6OlYdJPfKdmaYVejH5gWxGs/bII0St5J5gc2KQPptX0jJwpEjdDiJZj
w6SPZGF2bUCI1UqPTZWmh16lic9qE9PHiwIvLO+TtBjALlcXCCR9yWELB75Ly10s
vxq434JeAj5N8B9Ug2V3VD+CxpGVNJ1T7AdPoqZ0Mz8QnEOEwx9xTLHmAmwlr6eq
70CnzOdBRjlTKPOBbbWnfJo+Mnus9lVa73n/+ZIjWD1UIP5cmOPG5so5/3jH+IPI
ojXRaNzfNo8APibjHsfJ9rwSwrbCy8E931bCPtjrjCrgdbF+v1uyb3FpcUMmsiNa
7w/qo5MoI2c946AdCkL5IGRMKmIaKCfP7S6f6ByXHukvKDuNYTgQPjlQIv6IY4Z1
16kFKHeQtSUwg09LKWmi5OrUGUdNj7Gj/nFJrE/qba2H72/34lVN8C8+gw0xzeYe
9dy/uqGdqn5ORNhQ2U2E6aINqPAkR8ytOJGSHV7xYjo2Km3ogCN6PUaEKcFoD+Ga
kmZP15MGWMBUZkPkJ5tYsYwvOALZrEXOEE55I5jRg2Zc2a5k/FNH2vfR1OIpBFnU
zUUaTUwWbK+ohR24jUcIIZR5QoGCbWfIGAOkFtp2nb4H1lctsRzez0DOtEni3AJi
4KPkeEpUPdAr6OlJJgyoilXPRr+2xd3uuZscfXLPxXbK/OGqy/9Zr2oGLyyL58B2
efoiGXtyfXF7GCTd3LpFmYpzm1W6f7Tf/yxgtE2571NBYPE2kgrYKHq8i/3+XpRU
qyp6/566ze1DW+fov4cy3eLBilfG7H1z8VgYVd4ve+FO8XgOQYe1JCZsGaNB3prB
n7+W0lKAP6gvhmUYxF4EVZoUhx3oqCrKFqv0DnE7yUbdlHbJoUcQsjBYWfOEvvRX
JUaVNgelO9x9gv3eROMS4ECUTAqZ/Izunx12glOLKGpYtdzMiwPFMDu7xCqyGIHF
rXP5w0TAFjyb1L1GkbnyGKZLiAzzUSCJtnuEpbMxfGG4r6DK0zSE+dp4Ioo27SjP
2w/IOGJ/ICCH569Fvw6/+Oqjoj16G4IS0IpRXd+kkpT8OaHx3QX5fYdkQfBl3+jD
LyRihW8bU/RcBPs6vO9xBZzC4yxCRzzzo7SZ0Bxux7tk//6prAF+ez8B2YVSeSQ4
NXlzzL/AC1TWmzHf31Af31xUW4U36rbtP+g4gt6KdpvrkL8ZAlt8OaTmRvehnihU
uyDQZVq4T92FcE2zWnovKuxIr6mK25aRpB3v9Alw3O009Qke0WhPcnZuajhMQVhy
dCAwbev4Nn7g9CDagZ0c9VxSRwxrkqVAnVu2Mo641MunH0hmDD6n96qvSTzR0uy8
bWQeciJV4oEG6GirFiXsrfuF53e+UOb2KwmyKcuOhu5bL5qAnUeMjkvQj0KuHuEG
YZwq0xZGptEsTJxNUu2C7xf5mGxM5bIQWaqDHToA+DjahtioqDQJAhv2PwY6yNpk
8OjnxYKKaEvz2FD1Lz9ZmUiH1vZ50Miv+ElaUULznharLUsSK3QI+QfPcQ8ly1Ud
3onRiSWhfMK6qHLXAPJUgX4kidxiubcMAaTjIN89Mx0q17+Q3r+aqbPoqjh17w6h
BgBNSf6aohmy58j87yFTCRusAdUaNGMOxmLkxKRIwqVvSHfxN9KhfbpuHuXKmk0t
E5l/2gpUVbn4xJ5BX6d/mKQRjyVc6Lv5K6qvl4hUv4U1OMoxSdkBiEgRdaKC+vAA
QNrv6fKjpFBf6XEjxMTET6kOXiV/sibiv9csV4Ik7bAWXPIO2E6PlwU75R+l9gpC
oXK0Qv81IiPLExea564JVgvjJYXGYvkzlBBtBejIlQ3C9PZ17fFCyYhprQ8qT7Hs
epjuEisZOvIs5EhQvtbOkCpzv+OBmGm1g185/nGPIohGzheUjm10VHvObkzHyhI2
GFQaimgltmhVbQlbpDtqpzWI9j9Gjp6JCaBKwI72VvW5P46q2iTpvKPRjoZP65i5
ueF7xmRtPQIgUke4Cqp5X6P2fDtXOU7RfNobO2ql80ELEffPEKgauyWypDhtbfMr
MsRR3RQh9yPwLFqlxRaPo9+IIcQur4c3rnBoSDGEp69sM4WcCbiDQe98x7uv6S2Y
Z/Yp5GkueuGAKgWaiXpNKOcg6tpPi8TL7XAOgQShz59BXC7bL3O3MD6/NwhmKFSt
D2plyXYRlRFR4uG/OYvpaw4Eoy0CD1idLlafG3TcG9f7jGkxX3iat19EBRmyqV0p
otQrllHqhjik7K8fFweXJvci6Qy/S1dp3/3Bgxney52xt7u7GSwgnBrib0OzDATK
ZJi8uqB88CdwGwkr3vbUKD24AkjHeFfMFPaEWRr9N8OyNavN0NLeqhvqbQspwiq1
2QkC7qOAontSN5wbxQKWsgIVV9XjuAubBOuVDjegpT3ajun1eoKTM23O5CC2yNyR
uf6vQj73Ywp+pBzaYEqyj8M6r7TkY5dKR+YCQuvlqbtzhIQHH1R12kbqn93PlA0s
rZYI/279veYeMZ9115VQ/tVemz/cWK7Pn5VZnaT+0hkNBor0EOK/A8hXAO7h5iJy
9sckscDBflHzkE70TJG5ktpzc0bYI4gK/Q/cKqyGecTxF8Z73o9a/113mA1xbXwk
kzm6iWqoaVaf78sdIY5MS9O+cxTE/3jSZrrwa6waWNX0J8ahto6AB/2kKckXYAk/
QfgPzZbta3YaUoFhIUdQTeWwnspvdc4UHrdKVozUsWWbeDOPL/IpUnnANVcvwhRt
WY6VKu2FhQ6Bv4vuY2XrZyLfAAsFpMamj6//Dq7gcd8N7KC0bESF8vIiJ9MBzt/1
cM6yNxnX1mHdzjywi7C/7eGNtS6MdjMJF2WTS5M/XlvL1RUoe/vjlgnknzAS1VZ8
1UyW97Q4VdgypGlfJRJK+tugXQv2api7f1ORzSDlUvwe84qRfD3J3p7gq2bl5UTv
Gmg01sH+JHwm98q/uLN06xXS450PICy7xxBBcPfVIosjepqnIFWugtVvuYhQneXS
Xo+i2KFxf3a/NX26gNS7sau2AQoDYJF8z0nuEdI7mfC+4NWTd5GVvtQXwecyGVuz
8WLRJwagPv1WJA584icsU9VIk2tY+t86n0mz68TMA5ecaWQ3S5RSz79G7crVYB40
Q2uEQL11/2Gge2bRCUNaiQgg/YelfW1ePRWl+dWyvbQXsASVPjO6m+4bgc61pD53
KXNolH/841JTqxSYrLJ1Z3Wguw/Q01ewLOlx+qVAoFaOz/N25ivY1L3EFTk2pyej
I4qoRVX26mN/v08AKlfPVHoEWIsU/NU0xhNq9VihzyPYLEf4c9cbCE2YABrK5YwT
w5vF5uaz9gvmaIWjcw6hHAJFlMbXrivTDa5wqGyGbIzQJnJ0PRRVp2zKHxWtkUOZ
myP5eYtU3bQqHZvSfb9dc2lpji0yOtwEqVXReXgJ+1LDNVaLUD59YwlMQw02p/bC
I4MnkIcsRBPCzFeQjSsxL+gsoFJcpXfKVj9aTONnaLC1VeyLSEVYU1Dma930b2FU
droOMgeTlfeYlr3F9F1yHUC4ITgnDksF0xHQa0lEsUrj9P5DEA5bBCf8SlmYHOvl
PpJN5+ub5UljQ5ge8EyBRmdq3yW1cptQLT/zN5+HUe6+jCVMowpIhhJz3Rpt7hdp
l5YsVRl6fuI8TMnhTmnc7pMLm+lUCGf6BnFj1DMeivf0jrrNT7YUAOVBtnvsD49g
Nyq5rQKdAsxTpAQ0XrMyMCksTsRnHSZh4OznvMzjWSWLDaGXMPmRcnUrlbndDAKW
Qg7GEEizSrHIGZrxCbOb/GDPKO2/GdFIHos89yDlU6UHPO6c+fv7OI0IlaAG+v6q
snNt580JjrFbocaUjQ8UArjOkXXe0I5PAoUIWzqjQfBt52MdQT05tH4R0G9lm5eL
6UZVfqRnXwPvWXZhZh7rDuR92vIH42MdpPMuh3WqpqpU3YOj89AKuQa0pXMbm6Jy
91pHNn4FXBWo40bI0/67lPO93acWB6U9jkidCt+IFgvai7tCMdcByZjSjbdw8xK4
HkBkL2zj6eYE/u844cpAhsj4x96Guvhy3RNkebPKng87AEbq2EtnLkaE1jaWNIko
1SZIMAUseNtXCZMdePJqIsYW00Xt5lSEUTmPRrKbyB/+R817wTOHVLxSd/YsGVW2
s5J5FB0jOmvoybXJdUsI9nMCNaB48/BZJhXrOHeJKks8FWonLdWBVaQS1GLslui4
qvgT4lKjUKHwn/nJnRiiLxJqLPjmVyDh2uQxv+rYz9AoRmzgDOxOEI0kAQVCl8F+
Oj2eucPaPMdziPsgujx1z1jApsY4v+1390WaZj3woRe539EzLA6MaLnjXaraXkB7
cDxGHd0mHNj5XrUsESwfG4M8rZ3OzN98Nwekc79qoAH5QUUMzcq06D2Fv/0vzQgR
pcsZBVo9K2EStzy9bEQewtahzT8cfoqKtnKrxKwLKz+fwA9/lJFZEzqoG7H+BEuz
UGRWbnl43Jb9oXISKr00a1Ct3NpxqCwZssDnqUZgwjVwAgzkUNHOt9zTFyaGo88P
TJynB0IjlNdlSFp0eitCxGddVookoDxR3V0COYnJ1H6UamWDZtIne3t9cFaYIKte
jPQWnOb/Pyz6o2qVZIh1BQHDiEDbVa7BQWKhZX9WzH8+qGRxRk08uTz6hZe61A+l
dkGR3pLVvnuBQnp9JKw1NwAVbogOSaOomctyD2W+DNqEGWdW1+7eA4OM9qN7COal
nHQMqEAe0XxWJqF98c39uqvhz+LMbm8nYd2n+1u2cULBeDyjSBFVNif5YvacG3T2
XS+RJjTNZ4PLnp/PoDn+tvkjJBlKjmzZgxYdGcNYK52vmiRnvT8CaybKu8UuInAf
2Xe5WN8O05yuc71XkuT8jhD6lPihBnq909+STghi4scyTNryNV0afl6+CM7jR1KQ
48UhzxeUFpSYkGaM5AVmz6rd3AAJ42ACftCConkn5Fve0ZklD2hLwgFkKgKNXzLg
NUouwtD7SgEji81tV4oldZnFVtHXrCI2K9C3BJhETiYHOrnNsbgPN5AxoaDCONrD
9DJYN7T0QjDrCPDSI58zMNEWVt06/RU+MOrBD2zs1yYrQ4TlYsWUdNayaqWvck0e
sXzASA03muWwG9f9C17boR1bKHaLSbWbnpz/kMcmDolb5sgEBwvAjPNT3g/bMUiS
4ETj2uBs/DTxU6i3OISMGVi+IuxAvvTn4f8xBYiQnqibySF6jkGtVnIgXdOYNb66
63vjg22yoU9UH8Y8yiEZkF07VuemKhCg1IKcYv71hFZkiGMXm4tBo9O6/G5EzWqd
Sf2GEV7NZd27s2roS3l2oP97CnV2wZFrDmSSfTo7o5hoRslvWcdrUqtIt99WZ3PA
b93stqKRXXQVy9+BTgQ/JK/5nJM2dcBwaDkyDTFpNbHb7co/vHj2RcT9/1wFYklL
+PUVQeFYSwkuz16HY0zYh3CWyGuFkxrwL4Y6xwDiDu59Mf8AsVfJzq3R6JsL3QvP
yKxPc2f9virEB/PqrTkorSHXc0wfl+AQMj9Man8iXnN3Xr+XouKPC3H0N1xwfzCj
akTpk7PLj3/CKdayaiFy2XOi6ZfXlTyvMfAAH8ERIziyPyHUOfl0ddp1L+IUTnrv
Y3FC0TSqXBPQq7HCV1/0tWEDCPtv1ooff+yxV7bPF4/9lh45XEi06tqxD5GGSnRA
euJYUJvlgRmwdYu7bNTt8aJ2l0eLdplWMOS7RaywPcj1fPonKcpCIii5wTvEv76Q
olgX4oi6Wb6UUMLNNnd0M34w0+GfRDGBHLBmn+Yf0l6DcjcMpQgHH05OEKYCy61Z
hg8FaRVBSidORQhowhVZMLk3zfZiBCNS2uG+navS83X293dKMqIpOuIl8qJqnioX
qXFm4Xv38/8JCdGwdpqq6BmnTvt21h1BB45fFbIp1Fbo/IuDuwRjv2Zw76MiVtiz
UAFRcwvlbwBljaq0C8ZoqWQndYmdJZY21MghWBmAWxUzWL6icZmZP/nQlwy/bT9E
qwVcY/sPxJzBMP1A+IRy2nm3QILjeZO4HXRuCAhXx6zjwUwJ8VOZ1cNBetusKcO2
6M40Uwh108a/G1iKlgnZ35Ijnev6XxrSU8lVo4ZDvWtCBIgLGapB32fmz9K5+k6k
WhQAXBlks9DQlHDInWbAJ67DtprgmlQ0sLyM8At0tf0r25kUZmDnBQFAU8dZuOh0
USygOFVFzC1dCuHJC+Tm65t2IpoA1gRA4GQAYVtQYuQec8PnrlcqQAUQej0TBgh9
o2c7G2lBSUcEj3tSDavt82fGTh69zxzyJnfPIcd4Ymh8XHN49/aNSOF637ycOWtx
ktT1Tm1iAVk133M2dbi6+Fv3E2SBYIWObKBlI2Me5gR8/LF64j+r3GGBM16fHTjH
qXhWg4MxPe0kXjP+CztniB0zwpL7KKZxKaMpYLr/CxWqQOvcXYBMG4U3DlzK1BDr
P2C3WVPTKWCn74ZMheo8pQh+m/nnh1DvN2s2AbLj4SfOuggG0CIwETCUIvuXAowR
ENK0CQ+oKQr3Q4i09L3Banynhk4DmropL3mojlpWgp7oxRH1m8S7+8USEI0a3BXM
yHAJ5tRwAAXJGNQwtbLLOZSeEHILfehHcIFdGQduFyrcQGUpYuHOGQH7XYI64gfP
GdRuBqfkLevzRFcvDFQvVJwTsVIvFn/rb36hM/22LyNXCMu859L4G9X23oOT2SdI
H9ksF9aKoGni+i9JBtHo+44/VwYMUN2uAEFbydcJY4XFfdci7m8NntL8G9pJjUId
JsrUPyTzgAXnH15aGK0XpzVX5+zKKKtuZ2XNaISGbqeSkhpveaHSTBBApAfgQdcO
i8mwsWYsH5mQqRhxLesWwxCD1x8RHaGTz0Uf95muA0Qe8dqxZn6/30bsVc0vM1Jz
VLk4wUu2QOr7Pto1lfukiLvhdXtNWT71/3ciWfN7ys0chvdar83ifI0omh09+Cx6
rXrfndM2tPwkVeJJRDTV90Su63ClXatRUW4ATy0EAq5RBYqLDjfX1eEomqE+174s
zr3VKYGNLjZMHx4XuhQWpgTCrQpoHHz/rE6d8aUUFRC99p3Vm5xeOa71L2fv+Brm
dj9V7pv+k/0eyLogrtO+XaBRBBxPiFA3lm0LbJAcmRrpO8qnbXkSeBoOiYXI+cad
5x0zKfQx1oE4cbUoskd8JF6BvgL9j8E4J4ALJMgYr64gphsDXyb5vB4ImJI2+TYb
Yb8f8NjzHsfKSD8zBCW534fqTYTxtBzLHDGXxNM1rwSSUhmei08DBXjIJv1ptyOa
v4WXjdQ8M4GrD3k8mJ+BwHOflXr30N516OeGt6P7lvATCC4ChjddTn2KEXpJdILf
SDB8IqdLeQln/uDRORIRWzDqjbaTKy9H4KqIGZSmGVMVJMDUjYO2y/qv6HAT8K1P
wZphAShx3OOQVV9+gpHBz6eLxr5v7rrIa164nM9T91rFyu8HfGHJHRctwMBPu3PG
LJy7D/Bsucopfa3nV/Qac4DqhqTdq+Ab/janecf//kr5JNMUszPdRcTrtsLa+AQF
9xw6pGRQvXX+Ig10oHVuCIyAdh74PxpJCe1+2cUcH3n1hpOJROnm9rUFVDFlC5QH
lsbhczzrQINP8OoZVhjOvE2cVwxnjqpJqF4vcjzK1UggZ1zlouBff7aHeib0sTsj
Ty/p61uREQ1f/2HbeSdn+G856DfdbVr+sGc+LcXLYqT0xdAracVJOYcHvBi2ZgQp
9cHW7y0lsOvA8KW9XWkjZxnqTFD+aZMzJGkxKj2e4rTI3bOnCnmiiz4pP+so2bDV
c8uU25jQGoWvn5wNBfisCUx2P7Yn8FD6I7xblBUdspySVgKiNKiPly2yOmlU958g
HdSUgy6I4Mdk4gI8b5twJFiLNQxxb1nRdoUENK0vST9WNJj8OsgpbvxmPqhLQK5Q
aBunurxmLbP4puxMHTJ2RexeF+UPNYTvw1dSeN0Lz75WDhrvddwP4yvyENUQPd/q
AeCpUdmYOS/Hzm9pUjIGE6g0xJushpuXpckcAof7W+xusW1EIJtvAU/JDemjzgdn
9RaY+TQa/vNKAmFRP0BhnX2tVfqd8GzGGqNw8lnQhBZHhcXrpKBI/mTuTcuGR6qM
9ydduILz9JYaOjPjx8VddZw2JpkXrXszIhCVoEuPMNb6QrT3ZI1+t/GnR3q5o99c
ZShsrtWrBGYFIYkHUMoKNbvMQzxqgjD/0HI/nvUH4HWJr//4oRy7TfqKtHkSZjjU
fTTZqyjK1buqtJ8eNACthMFcCX3dTsbZAgBS5hRgmFzgvfhS6v2p6vg2j+mqzNd2
ilkK42mlLeYpTbAbJl3V0s+xn49IzhLjj9og5p2pUkuW1wV/XU4c+DykXC/85IJQ
Fyu/Cxd+/96ixMDfvKK+ZeWErd2Udhtqg1tvuggXU+2sCD1NOui3wjmlog8IxZu6
KuR3OGAAVhlhRjWCTimLphf5vFZ+4biwp7AtG4ofFFYFxdn2Bfmz0vFFIQS8p4hu
a2rWYABC+8OsLN+YiBDSlRq/ije1EnKCTmLSVLfUZ29Yke3xdW3Krs6priAQc/UO
L0VZ/ws8UJbuloEuxu5B4pM/8DYeNIm2Dd7HnG0WYjncJLvPjo9KqipQOD1SLiM+
/jjtBp2uJ4t+CEHuga5fiLnxZBtDro5+6sgW79ioSEimEHgIgmi1umTr1CE9jTen
Dyf13/4KLRPN7rZ38wnEHsOboRiZWrXkBuWaVYp0v30wMrK+qWYB8FzTiKAu/KZ7
m3lX0qSQzHTXM/w460RxWD1mC4czF4VbhBeENwBhKSkvoQx3Vtd3S68zTBLRQ/nw
9V1Lwyph+gABIJvFs+hr8j6g7de2bikeE0Sv4LJBl1JKtWzUWgx1oJFSP9j+xW4j
eyMkkp/DQhy2m3DFoupmzUXG1mJne4DqCNFkAhfBqHYDFh8qVN2RTbo+vBuEpR7V
3+c2FuZ5vvTzyGwEWf1gOOtK6zVn0n9tRiLreBKsyFxMOf4kAkxDTWK2/09VhFjD
BLC1k8jCd9mhcyfatgr9CKXk/RECsueoc2dytZYM4UEh24IcUHyJADdB0fgOSjqA
n4uD6Lx5Nd0GIkZkRRQzGYutlwwu3G848giGy6RcMGiLuNlBWPPWGDo2Z3t8E10U
Mn0YgF9mq8HDj7Pn95ZrcNQOnufyzif41zD7VTW/p6BI6k/YkJh0RCrDQru3S9mE
HQOdaEHnuL7/vBJtp0vSOguwFPGjF+Uv9OMoHOdTTbC8coqBte+E2bH5unEwaVLl
j5gE/AjPyrdQC8qtJE4iUjbG4vh+hXPV3WogXbIb4vxVcRfofn7rYyI7mVcLEome
qDRQzIE0Z5hI1+nqPmZzjjCLMzrdR8hUpIXWjeR71hqcHKHHbZrMgMzY210Q2lgP
q/NAi8F4/NWQ8ASdgSdkvkQDrGVlAJHXZ+tSEKJG6bfFoxqCoZGCfQrxbd5EYW2O
DsxwqWccRq4D3ILFrcorxPGGZ1mIDPMZnHP5S95mBFiTKtBE1b3LXhARybXr/8/R
3q6LT/0+OXXPUKkuqW6BVQaGkGpElKkVR9Wb7HpQNF0sxxoY2vRlIdX0iNtBzASc
B0IOcAcwBbHVEAAtGmBV14KQ6VDQoBsD6h3mwzmgzqO0sJc7fHmK3i2piLRAyw4V
bc3AMDX58mCAIiC6bFJnrKBn+9dpoH6kPFguwpmYXdkhokcpEiJQpBFdwxTR/OTS
7KiLXQGvgv0UporAaHRMsH7oT9E/IQ1/KeQexBmUAVXi/raSSH9xkkGYZYeR09eF
AKLT930XRas9MwKgX6KS+ohjZkHxCeGrx3Lk6kZxYDbavVqKRaWdibKJ6C7ildo3
aktZf8x5nbAObpAPD430uqoj6wlKlBP69adCJQRWc0aEELR9KoJXwihSrn0uAvDS
PoZ4YNEKGuJs+sayQjO3PFVe+5VdnYBGcPm466VSo1Vhl1dwav4aSmoA5oJycd+1
qpKb3QmuAHNZ9ZMCyAUm9bfiOCxwtCd35CVzpG0Tb2j4OZONEiH+spT597qeZx0c
j3O6u8wQzFWSWU/7AafijErDECQLwYYI4gesbbC0eUXCNFD4NHilQo2fblZA9sl9
ka+EciY9xGOofpAKVkndQssJgsvPYKTFZ3S+COMcEPA0oeDq3MPWDjYVz5G3IhQt
IgwQrL1lzjxcqD8LZb/5TOdITtzkoSHHNFjr56okjdyEgd6vXjUb2E8oiEA6DcIk
w8wrJYNHoiv6sdzkO5Bd8QIn7syxHP+qhi99PWlF+GN4jJJiXPUy3CVuYwnmbk7k
H5SzW/FO3zyIo25A5wM3CO9nswYLT+2MxlUdhd3/bSFh9SQGuDFF+BdAVwI5J4/b
ZX84QaQg6luOqm8fjrFEU792PS7tUwit94RGJP9kO/p5ci4YGPVokzfJlb9dXHcb
TmD1P0wl8RCg1567Z7pFQ40LbeJ7jfP8edBGUQXhvl9zchHNOmjEmCrwtoQed8Zk
DX2qmLzar1+jz9i5NjCy5lY0Ur0/5mE/fq+ZnHDSDpj1jJsSwIj6d6pBIn2Y0xs7
w6XyDn++cz+HRoAX74qc3YGo6bDg8iSjPZyvNDkP/IhBrzFsrev9fKuUNeh0zIQQ
PP3GG84ZLMDqS2YuAlBbr0Yis0F/lNGoEEDr3IKRnmCKSja+fz+8O+qg5Opvz13B
cHJQqYlqeN1T61St5TzjbY1JPv1Ebi9VBuUo5NwAWGnnbEkTkscybHGsaiZp8/1h
mc7ON3XNNg/dWgcig0UPiq7nyJV/HovCP5FPwJwCd0D7rQtYLbw0oRzgxepbSu4G
tKuYWJKKtXhtMUKBYfmx+3h8yWVoWJ2eNxaJaWUwOPwaJPJ/iHbCledj7SzqtUeE
jkTBBuSjqmUQY+fxI9eyufHQSLw/6d6Meg5gdplXS74HHX0YspScMKMDyHZPI7/p
sUaNYjw0yimH0+8Js+0/ZUHcFTIIb/4tUMyq4HKQrV+b5G5B1n+MPIh8iTd7JRKo
38hqIgnpCk3eu52p7JQPWxFZk4rEowqeAdINETjWK4aZXA9Upu8G9BJC/eSa5/H3
VvT8QaeT1YWhmZh6zXQN1+3Qa7cyeOkZjWvqdIS3zdHrOk66te/IS5oOVMiNU1oW
zmQQlg/5NoX0/IfOzQjuonheAZgH0cQO/Ou1SeaWcbZp/KRe8fYzb5ru2S8nXwim
8E+7Hotw4yOJinQRziTgj4ro3KSrUcLTDCBzanKJBQc6sjq7Ql0461Ybr4C3PIuN
wlDjDg2U85DmD6IBMX2DOHVGZ2ndl9R96xCZj0jgr0H5IwExF9CwZG3K94rS4yk6
51QJfTYDQJU1BtnZ6/FKD65GB09eNegQShWzhXdRM9yUxEpFbD74WfENuWEFoGRA
KT+toGryih4BN4ttTwHZUcQNx4GGAfV0H9WhNNPBUcvlbLAmC2E/rSjF3E63itkO
a3r1hxRtzZIMGZsrEnZcCg7nZYU9JqMjoA1ogth9WK/FAxYVwlwo+UD/D5jjvVmv
Pcgto4OtyZHMtWKcuy2meapI1ny7YZT0xAEawf00ETKY9MOVsCmMK7DRVZU+hpJZ
JZB/DiIvW9LJTJamPrZFQ63lU9nHWG5fSa2aDwhC6myu5AIiB+dlHwjGPpFf2RDI
BYUYm6jyawunJqKKP8rVRm7aJp8NhrZEAy4KF9CocS2JzJZv5DikdN0wIwSECX7V
bOuBqDCNBUo7KJYa98L4vEwvNkVV/L2/soACCm6/yNRYIMy3IIQIUY4TrfmdHmKH
iUtI7XKHSyHX2s1j+9A+a0SIzbad8g9LOsPzio0tXIu6DmdD1+E4rfv2wckkHHKY
/6FaZXi4mWTX8v17iIfcEhNCf9OGvnfZbHU3SzTw8kJYXw3kclSCdozBwQ/j3bGP
3hu+UiiwT4R4iKH/UH3kC1YRSDXt5baZ+visep7CT2vRTUFHwtb/vrN7UJmevuCy
GSAbyQjFK5R16yGWxbC5V9lmllNd04uHOPQE+uWjEfnru6U57no/xskv5f8ToTqb
YApn0rodCFudMbOSXaNzYMg9B7Om83exm1yfttrhMqP8V4rxYMiJ2GVOw6Wmj8H7
tYdFUt0/ph0TDn+Ciz7rWSdRLdMPg2089C9++Sm++B5DNf6Dyzta8gnHw2HvquLS
CkMRmVpIkXsrrfnlIK5ob3cy+H/9k214HyVXSllyRZaz21nhMyFHjbPh7wgNfqZ5
SJa6S/zOzjct37PgNm/W8JpLqYXKkmpC/MswradHMsMqAWcrVLRNXoI+ia0YwhaX
sYkjq0n3vBwkzOdTW57sS/UK5jxExhosXZvowxn1MwbBxHqK6YiwZ9iYiXZKbdRO
NvX1r8Vrya9dzGdoAGqYh6dWVeCsUDnaGj/cCtH8Qs8x87xGb6cPXgHn9kwKQLMp
8hpU8/2WxNyzMGdIes9jb0Ab+i1uRMWqEVtmqBKz7VW1mf99gd2Fxts/C69Rl7Un
9NVh5R4iTvsF6jMfIShJ4ffNeuk7EPsqiFIX+VrfvQsXJZmxuA2LjINzoDbE3bkh
O87/0EUCXXqMXaPm+3WeHNpa/daEhqIggoF72hSfaLOKy2a2N8HI2eeplLR5pjm5
xFnjJ4PIDRme8gbw9JmtB12AizqlQGlkrnfwdm8Nhr0ThKt+VxSDSFpmy0U93TT8
SLPbSqS4znBlXge6kWY5JAARJL9DA+WssVlGN7AekziMNKU6lo5dSr9Texqm+uxC
TFtCt3lUJLaJ2c4oj9Yw+l3az0pVBCeFAvBx9D1PlOEFXu+yfOL2A5B4qZbziiPX
Kab6KK+X/FmSmOfOsLPeMkj2bPZ88GjgkhPmCDaQTjBg/rsHmeYvzCDwRrRcCOQ5
xC/VNMRcLcmvLfIK2L9s1QB/LUPjrYFPpHdJwGwCz70itmzN48x2kt6060mqQYGa
RY18lpZk2HK/MWGaD/AgsPn+mDHqzQl0iond3OY7reUL+YxaKRvAGZ/0Dv85meeP
kr6crhBCWyFsdRtWQJ2x+f0AOzsjg5NW4HAIaavClBxm7Q12Q5MHnzrQglW1p+Cx
chzz83qVdi6gFYaV2yibjuBIeF+Rdb9e2OEO1vYgn8+krPJrWKAOhZIcFzx/CB+b
dwbOlwjzHCmHRbiUk/5Y5L5YfIWNcscoTAleljJeSJ8TydDk+G8lmswX57FX0+3r
vYlVoftIxVVaDVgV0ySb5DQFfR7s7UQKJ7Ec8yK3R2d4Djni0IWOkjkeuyRDGfJN
lZScmM2AVjmK7XcAxJwf3Rt+S8hd9EcCcVhsZpmhKjTSKJuk4Cu52StCWWhEM7U4
geBJ0JUJs/h6j6db+oCGDPM0jsR4shY4R8ECxZYncduWbulF66poOUdxOLjWcUAE
kLZ+FHkMmNgkbeujoHMtaaEy5slIstaB4ycQokD6EYM2RXFoGxcHXgWQb16yqM71
3A1Rih87Rp9kdWl9BfxW8J6VrVfC5DwkR9WOthfjMJAezKvgsq5GSNHQqgtJt2l4
EL57R4e2GpmEHSyTwMwy05hY74byptsAQqndkdIsn8wGvAHXwcIDDrwMjoZY1K98
5HXbrD0oucTvCZKl0n4td62Jj2wOwsWib6NK8RoRMCHM4z1e6w0MTQwkqrEewLBg
PkO4KEnOHcJIYQHf/AtcRP0tTWJ4+iXXfT8meNDqLon6oubeu3UiNBOw6iTABUNj
uvbZq527aTVpDN9NaC58HvoovqJG9DaX2FSsXvNAmo9luGUFgXiGWb3k91ZPO+XW
1lcZIRmGwM0DoMRlbrWv4mlu1jcnSuurt3GL2xXbEAmSyJmlwzBYM6+SQ8ZleuuX
Iw7SATBtmuOWWXoVtrYeTfY4oQ658ZKSIvCWpNdJch5xTwXooX5rumQzmXDYM87s
cG+GSfXmXiWhpal3tZSYvdtYeBWyZGKqrYlvrl2A6JYW/P61PPrKpA3fsE+mgRbO
XtoRTNh9Ye2ebcwn3EiD1pviPHCy+IwV/ADMB1+FIhJSYaqHtUuBMkozFvfszuLe
8D1J0GKmywrnbsmCse2Pe7Tx6vhl2hnyfyuRUn7RdnvX1mln5uB6gJuB+uPApyi8
yhGcjH5M0MjuxInbvwXO3a2xhulnNazIy/w6zcnwYeXt+Z4KJP9FO+feZAySYlzB
em1KV/u6XyIzcsZon3lctCYO5nWLnW+dhsgcIwW8fDo4xLZW6whRzWp5V51XTimj
kqYHlxiGD7WLuTER0Y6POEpzho19Qz5xsqmjKoGIB7wRnSNqxfXDrleSVq0wfRE0
ZI1EJNr4JEbMNfv6JJVm3GGWWkOcJYauEJLrNEYSDpfDaFkTnWVwBFjJve2sSgrG
8017tMXz8l65+Bs6F8JlXdK20d2PqW+uKnLCnJi1sZZ27W1RZimyOZVioadGOkzM
dTeHXOBdHYrmdfGDBRhi9PZhmGmyJ+f30RLPizvVTNRxy+FPDL0V8Pk8Wsu7G/pl
77f7TbXQVJ1rGw3oIzUC0UXK5nkJvlV0s9RBbJLM8bMrQfZ2u8rd5yvh4++tWTtq
G6o+K3xhtZ0ZuvIje0Z85POzYHdkwLbt2zTZqUqMa2fY9CCgCOFPOHKcSFqJZ4EO
WPr5it6zKAKouTMt5Ay1oTiH12ehlgSeAKQbMXR0MrU/lyQrOIky5oAzjFVhXlmX
EqYWMi0KvFupN22v2KIjhIlp3AO2V9eRimCb4QL3o9syJri9GH+fuc4JMAjVSnSg
aJPMxEm1TxBQ8MWSF4+PzDglzENkc50KUH2Ck8pGNKo+3j8+OTOesghEjTr2lVUj
ChtmC8OvGvANd5HSDJdaxgxM5Te5Ido0j6Htqz90OPj14FfpYUdgY2LhukVlL3FU
2uNT1I613ey8fkTdawckQ6KS6YIA8W40XOgSTZXkxGNXvA5M0cjlQ9ax7gJJdGrA
7gE9kf7vqmajq6iYVsQoSXyoqRPkUaeHBtPXo882ZxBulmyRl01LyhGiQnsVikkT
q/lGWq+VgX8hq5ZueiOk5fRA0s7+/oPgJNyVO2n6+aSZtMz3/yt5B2cJiSErUrkh
C0mRneX8cqBFbXapdKp/axY1Fkld2zYR8oOF/MKPHGGIpXazYTZ4iOXK4AiYXRnJ
eV97jM+m1DhE/U9xp1hSgpKzbF5s7OnhVuyIDFEF9tcnqmNA0JY3iOHPwG3wWnh0
923W7CTFulvFcZ2m+VQqwwXMmtHqN3qi2IxyBtugdXBumnMBYJTJHZK0ZKyPZMk+
vdIQiNKZW4Qdd/nfW8Edo7tMfO7qA+ZdNifJNZyh5S81LruSzzF2ps8RSGgnu30N
1WEnbDe/Yqu1PMCH8BkuqMlSKnwgSZCGhDqeKUGvdQ3M7CjY0yOFLW6p//+WRWTX
14djYCqAg12EHQ4F77VWsEJ9E4qdfS1LRC+rB6aRcIlQT3kt+nsfXMmQQGLiHTrJ
GptEsSYFqalU/YRNd1CuV+yBMQdhDUGig7hhu8ZdTVNUIZmM83LLWD0OKtSrw2Vm
Fumz7SLNJPLj5B8IJ4oqqPqjXjcXj7oS/RCywhDuqtJVAYVy6zTN1M04mQ5HELbu
CpnuM/lUhf9BOsBXDtEmmKtpgZILwO+mQ8U9Ktf+j+lOG6i3msy1rwYGWe1DseAu
jPiF1j8dR+WK4MWG854V4B8LEn+qx/NCKNsK+SokRl8Kg0fHddlE89qDPymJ4u/I
mzmtliNupFSZ1GUq7qE5V2EZ1dHfam5ke7F/g9O6eeTx0IrLio0RlYiXHWh6D+kj
AoanwfQuexBzrWIMelOCTusHsAGEoaiUTMcI3Cx+fjuNApK7Wzl92KztZpEhbM3H
e14AVpIS/CKrCe77lmM37TkYtdd4Q+WIld57dp9UGMjnQFGnkEK1X5Chl/s25gMB
TbN0qAIlPlT3k/soou6IUwkUWjASm160FgMh5J1E6cgGVsG23Utcz9KTbyrjqWUB
q9+73Dll5tW82gsPNP/BpQcunWjqR9aLmgL0aqvPKSVL1jjv2x7q5JEVBRbiCSAC
wY4ttMSk3wyc6JIWvJGE4BfUikwo1ejQOqhxOVabNR+uSxmTWjW32Cobhrw8BrpY
md4qTH2tuej9QN1ksXE6IvUADdJdU8fK3I7EvlmSQhfJsOUzh4rY/+ZCcv7dhfEV
3Fb6+5QnDK+2NL+M1+8pF6a4wdRdskIpEbhol0yu+MdDnGiOLSns7bamOYccCtVN
9T5S/r8FujtqTfdGmoj0xkNaSgdNMddnPZMozoaH/o+Ww+jUcMILpjTHgJZd6Pk/
P4Mhq2tGTxO+lI5mr375Py0xikwRPeUqzW+hmcNelBmtKyz0ESb8S5pHe4VZu1RR
7uefdnlivmKVNMiSckRjYYAgs6s4AQdAuV1cnLGUcpjqXbAJW0V9w4hTpaS4QGAk
Cj9MTTug/OS+v4pcUXJ6cWo6BnE9vsyAG56Ddtfw5xfXrzBXdwApx/T1D+GI0hH1
8bnhx94lcFrc77gTGv4L64CLs29V1zj7InUTaEO5vNewNg7izvZQQD2gBp/Lr6Ha
QyT428KIgWCgnaVI9ZYriPjsEq/3lrZYn+QqzQg0t7K6FkFDf0rlgc2oxua3QdQI
cehGab0hzKiaw/99r/Wk+FtXT8IWJknWhlyMW7yVxUT33cKtnC7D5CvsOI680HBY
HhXMV9oxKC/EFgWfiTQfT+7hPRiRFtTHafxG1HVm1cL2RDS54l8CiIOMEbR5qlyZ
k9EXfz1UA1ha9mG4hSLA/ZBmtQ8CDMbTBi84UvO17FHKslgRAtzufbQlcNwlhTmg
Ahga31LQpbEGvoy3skkN+Pe5YlX0WuDTT8N+ZTR6B7/0Dz8MvDf2ijJpzJCfTEcr
w4HJGpKA/+B7ywly0VY510IrrcTMqPElQjPg1tYNsijSCJrx2gU6o0HlD96QKH9f
muBO4a5pXkHpeBBKTxX+9XwJybA2ipaLF20I4TKGkf5vAWAUEn0tyalEJ5B+x4sh
jKD9vivPgR4LgHyRGnMhaxGcTXJAJj9xqo4d+TBZs9DuVJtjQqw0mXWlmSRdKfrG
LmPrcr70ZekOABxRwd8KrnigU2t9SJWDTpjVoZHbjFn9LwF0fiQ4/Hfs6Fy3ZeX2
WDNsCkFPkyRKt04QRgmDt5SiAJu23g9/Kq35S9Nqw1+VILYdAj112DMgdVBJZWrX
Zqe12T6FPMGgEOPRQfrrO7l41P2DW7IdCKP5zp9sgfV4+Xir9gMN+Z4LCld0dwTA
XMoh6bwqXaMQewiNZsp1s786lbBYd+p6P5keExG9m9Tjnm1eXG713NWJLEBCxbW7
GiUyWfTKB5bG4HiMkwlkG44JOQzhojbz+Ovx/YhoLFN1YlQO8DlKDq9yawFS+DfU
Vz8leQBPztIXB0LZERuUAWakMr9ulnYu444DsnXha+Fflt/s9X7UiOWJauQ4oIhq
DWBVbS1eyitiDUI36ljWgsh0c7vov5zakSjotdTdwkYb4WETVp9FhqHZq+4ZuF1M
f3kR4dfZqEKbJpT+KQ5HVm7HshFIfRENqzGu54jkVeYcTLIVyey8wwG8UY05ipd4
h3Gjm1YN/HYDjJhCy6xHTnYac4/G6BEsFrv21/oROqIG8cqVOA9dZZsSnvN2NBwv
TIOuevO/z1YyCp/odLXn21mnwCUUvagWW7rMiuuPf7hjoVRwL0IjSMA3MvRfcs4g
Y+8acJs4mXdwTDcz4MgEfldHUnifs0/jlYp99Ghzf3HfjypDRXqwzSZ/4uuVhR/I
YFHJJRfMr+ewd1qM/mqEPudXKjGOhsdijUvN+rtcppisqb5NDBwpllwu4+7g6tJW
1TY6Gvb1aBz+MbsVOxmtUGYLPE+BYByj+p/5QgKaCnstBJdHf2cqKqIB6TUuL89M
cBNfniqsZUOAfOIu/9vTzY54lrLBQbYdh6gtjp4m2wO9Otp0RNgvsygF+VmJoX+s
GINK7HZk/7p2Dj2jqffp2n3D/cANN62DyUMDV7thNIJONNb2Z+MJC+hoj7RgOihp
29fQePt0h09eLQFjioAPeVt9fMIaVMES5o8x2vaaHVLi7uxPt+cdVzA1rbV4urph
NGkBHbTuucRTX2zvuOQRG6SeCUTvnfxAQZbsM1bJ2ePtT/KGQ6nTiTqk2WCc1W8E
YHTmKUYEvGT5hDQK2RUfnhdnxn1YzWvDM7vZ56a3DXvS73RpRy5jJimd8b03NyD8
wGg3COEvcdVDz7piD+yhiQRB8trlx8F42VuxrQkYdNa7GVVTn9sbWy/nZGNnFbx/
R3EYseWJtSOyGSkLz5LTyRZU+B3OnazNqrIZvUfPwRU1gvQyO+8PUrYWYMGe3UJj
w+Zi2uk5f0ZzsozmrbAtD+tT4dBSDUtTlCW6aNDZC/ZVhtEEOLvXAZ54I+PumXU4
bLvG8LAiFxY9bgAmFZAyR43Y36Yq4C1rawcRZyMbLPZfYtH2PPhjhvSSCHA0vlm8
OXsNGtMDJdHUHObL24R+zvh9qHq98TK33A8uRhrCeQsLkCteEZ4yayNlcbtXKbU/
aMHhJvp/xjXIL/MphvoBvR/pAfew9IGxFCd4oy1x/UmEnMFNYlr+9DwkChx6lpeT
avG3AX76/SlEEEtfBSz23t9wNQRJYSA5qwHPU3MpPUbt0xmkV99vIMktLNYSMP+G
EtMqWDES14Mzllf1aMXKQ8LZv0cVX0CuNSMG1fpC16hVs4zCso81g2U7dzzJtXXe
qqBZma2kLahh/4oIxIXxvRat7ZzbM/6DqIt0XMa+nZdMxb1v60unLZr3pHiP/wlB
KYS5TAsLP/igGIjQZf7qunczEPvQXpLl8cHzkHG1obrhDGzSiSThwDPBULOG129G
6v3mvk0FfXOSnbQsNlHhwQp9DWgEqkf6uWnmJ1v+vOoJhSbT7FCqQc+6KU26Hcop
YtZ7ABAhj30MZr7lI/ClRr5X7NxA1Fo92MmDNYd74kv6mMTbawYEw4sv77jOXkfU
NbC8AJnirCmts+qpX9gGb/pbYw1liaEDaIU52iTM1xla9OfUw7riQqHGs2Gr3146
zYGCHQxDAJwOvRMcm6QumXzGyPBCpZvaWeXGm0VSp/ONjAttaGvoopGptnTAG0+5
9z7RgbVWEenqDs1TggYDu1boz7L/R449hxGGitV/yFSzWI2Bu78JfJRFv6oWjDtB
mXJWW7i+7MVWL/CwkS+rog2veFbpMEo0Z62Fy78uD3yXlk+x2ZmU7Ui1NcFT+bNS
jqk4e67Hmm1l/nBc92/ovDgWKmkHOhZfrTlNGc1fTK/EyDFwaz1hZiVpQDGAj38m
utocQqzsjsxX9NJiawSOxBGYgmwG1DcGVjQqFaIivwlBGU434dcg5LMx5oKiY4KC
kuEIDn0UJ5BNt11N5kRRzhdK/8D9HU4czLA+rqwo5yg9aH14JF4STQ3K6cUxUrpj
1rT7oM40HL3kXaswg/O6VRfi3lQ+j8dZnr+pfOLKUQpMUZh0Jj44kBVKiVArGR2c
5kFtZy3OJDBcsEg0rEGlZNyiANr2fqr/4Ai4Z4bpHIl79KLRm4YhQDc8n1fh2VTE
KOXtaEFGol6aeyMyh9cljOTMZlShJtQDSKNKJN0hFau2RWQML6/cA1LbkLMHPqKK
TUFZAldYgmPxaU0L5RmMsJghE5ohm5RTODW6ojO05hbrmeP5RP0IZIw+6TlSmrVI
sGDWPOnMlk9bfJLtVVs/kF3hycsfkgnwZJL+QyiDPv0CpBjvEQYCwEhvIPFy4TdK
GPcD436a80jVal7jN/KTI8WXGj/8w7bAEKS4WMItDz9bl5S+7L2ycv5BkTWg2bDi
50AjELvSaBqjeUZ2MXbZ1V/FFZ4t0H0XtbI6NsaFZuGqlILCM1d+hV10bafuLQAy
hAzl0amh1QmmrasYfOxBNhp7cLvg5d/soOhuI84saAbjNE4LDWtcwbCx3CSO1OPO
Was2i3HR/kr/cLnMqsB7OKZOG5Yc0bHdWAxM5vkef0bEwyIBEFQNoqgWgxRSJbGU
NoZWLru3kqttSTRRu8vedTt79LVevajtmsbOTYA86CndU9qvpZ/xKKh6H+up9oAd
5+mnWKJddJGh+Ekgc6gyBSy0jLb2k1On606OP7LP1NajIkm4+jTtMqzEUSVM5GyI
v6ENijgZ+PirH4AgkCAQoNMCUGERdoXv1Sop0PQNfUNrWkLu0xInRpjj4AYjfWQ9
ocAgboCsW5vyelLQP21HRSEnrRjiW0lqZ1awW/ZgQe+XhBe9j4HqAEM09nFYWKJT
CPIolWOHxkHJQ6Ba3HqPRK7ViYhfBizrXLCGF5ldmIjvvbqLoTsZ2MyRzdOyEP24
X3pE+VIvZ3chImFPP56sLpXjABdNZ+oX4oIgzXcfi0LOPsyG0ssaguSDEs9AitpN
WYYgDydtgezc7lS8upP6lfqM1Y6lg01lCjKdg0u/lVCO4KFDDrII6g7znibaoyTY
rGbv7eZRtgKpJJ6qqSP3eWJBzSCeAnmxKoqcC7EtYYT5VTfQfR27JMoH98vXt7cA
jqWMkeULAqgEBqUPBSEse3b3/yeD6BVGcssKgvr4ZyfC9V5WvOcU9ShgOjlIEmbk
onHqy62IidW0uKrmWCsLN//j7P+fKbDDhEvdYhriW2ZB7kUw6SFo1J+XPRq0CvcX
SSjm49UNfrsv4DbQCdeqkjfcY6ZHpPpfUWYiMRUfY4N6GO8nPvelEzTThVO9Sasj
xEBvRDMC1Lfo3JuoEql8Mw+anWOxYH782urIOF1kEX8vYVLKR8e10lkRP9xa0mUl
AnFM4Rhfw0HHPOcscAoFSpDHv0ZFEMuRGnuFIRPJL0UAHe8AVSAyS2t8tIB/hKtp
yfuZbZsKFk1xWfIgd9P049jd5hvYllIdxOogJautwtz65LobO0k2HuWZjtW9KTLf
syljo1fE75+4eSyrhQKByQhVaw/HXBjn9VYmrkynHyAqFpLO6bXk7Dhor+4q8NFU
JtNdUsXcO6kGSEBRZYo0hXlTsr6uUDcHkT+8099UmC6Jo7mi3OCDPqwna5H7JKm/
3yQngmKMsNYuav3TPNvzx4kmr08FvpWgwkq+bw5Wr2aYsOArVEw+SpnyU6ZEeH/n
2d8L8cOSEoiNK+ppIIFaCCsyE/nkLLTt3AzZYEzLVOzC1tDZNetyusiGlkyZQKYD
xnfL+pI6noBuubyURdxv8Mnv/m6RREK3LuZkvt76VC4s0uq6E5DTF3PhBOhboMwH
zssx1DqxlfsHjMIsCsUxcsv0JrOcnJFhBNTt1CFC6dPfRAg49YebO/FA0RLQ8IcU
PC0The77PCLU6qXN/fuVuihl7GR4GD4/IMSwvveSipeVQv9mb5BOTcsXRlXoRHVG
O/Ml+S2RcPI4MJnbCOtmcmSN3XmKST5+A7Po5dw2sV8qSd1Edwiz927yPq7r53cX
zJFRXY1M9DCfg2VFz2cPjha1j4CotBmn766D0gM41RlIijPoT8yYxQZkSypkctvI
KU/YcMf8Ikoe0WjIXevyZeH/F0whIYgEB/CaAF14Hg6BRqIVG8vuYNI12nNyX+US
BvlVjN/CKXrhmsoJF5KvpJ+tvFc6rRRzT41FIDF6tUDxc/nkU8T20TvxW+syu5vt
Vc9/PsWv1b3kpcasYqHKsnnssCfbHMe7uqWYU9EOcNrwQPU+6RCKNXNrYQTVwc4X
v/2rsJsrTKsCwA5JOK4eZmktgDaOxBYz83c28Cefcqb5yDs301QjtErYol8oShN2
kqutwvx8y0mmP5qBV1cl9fyE32jcdDw1JdKRlaR+nlUD9vzzIRsxsC5T1Z5sgLCp
0VGFXTKFnRHkhKAMWm8ZvkL5sEBxletjTxJLLUbvPv1t1TNWUrC6PqU+Wnlmz4+0
pVO70DhvH7ZWAPIECOEiZ5aS0buVITwffaopkk9hcBWzfozHT8yyqde9a3xUHdZz
fjUi7bO0rJlpRB7HqkRHu66JYUWJR+9k4MMQEWLaS3kSkIBb9oSB+RlX+66jRKY6
+gpHalIWEeb9KvhxXDvCTRJU3jQgnzs04m9t6ZVW911TyaCNu1oqUZYdo+aDiZnP
XvgzhQSXpZKW1BwEq+p5AkkdYnEShpA/37Q3UyCrcLkig7ZKz7q1DZzQyuYHUZMl
uMkZVv9cuNKFPo4w00fxkYjLsupPD04h0mUtc7kiYvVadBZj/nb3iip7aIdw//2C
DEi9F52AMbyaaDXMyCAG6JWAWZzKc8D/0aOj0N8XZFCGJsAfRmgmZvbXT6sj5fLI
+Ry1I21XFC5z5b9Kagv3zDZbRID1gi3fUWofUMiEDBt9Fmw5AhdjC3VVWbYDk6wB
0Tkos5xruCIW4+qgkBX08oGC2kzhE5ZaUgQ9jlNiSYLlcWooBLsYcbHVW7zTo9Pk
z7kFa9r2ZuJ/468Vn148lcdMIeUIeBSFlAmbuaymELU3sxMuYwGetJS2uTyPnWld
xF13xUaLZP7BKyYB5WWXVFazBtDwrusYv8G8PAcTSE6mrOsQjm7acY51/Edzw+Z2
JW+3CHicGJW7zFMSAaaehe2WUv0TJl/QzFW3BvifXvIGiKRYI1SpUnjIOC4CgBlu
vVME0Upo093WRxamZqhoeCCPJ2zn2HVKYLPcRwrZeKUrOJY581JSDdpaiNpHAGiN
G1jp/BjjLb1f19YmHd293txGgX76Qe54rzgP25fwy6DtiybZdZiQTtXA8Li3jfpv
772EFn01a6tvRhhNSQDL0eDm5ATt8IB+y/oSjB6+aQGK4CMJAhCzS2pxaCnoDRVG
KuqF+tTHJPQvdk/l0qlVnzReb34c462Voo9RyIzWBJrBAx8skFS7NoDjDdHYWTMc
PBpLHir/YdebD0CPnP4iBRi30NkON8T5V/RRSgLKWmyOR2c/eDPpYNn1BfV8i6Uc
r0rTYcLTl8iBAlirl5Vt/V1JnNUcYe2BQYF2bJ5TBoSxRa2SoGqvK2gPtNM3LJne
kKlNd3n/OjtU9bqeuqEgGgj9s1Sa+c42IULjQ//fkLrksKj39zkykrP7FXNCNVEc
sosEkjXhfyhAaF0rgS8KlHzABf6jeNqi6o8+HHJStjC0k3VJZd/zMhKwuxj7iv1t
TKaxpyCDxRpAFeH9At1ZGTnUiahxwUQX7Q8ImdK221qZdB6ZyaZs1BMf4jIf+gZg
a0z6Nh4A7nLHZ/MbdJQSUa9pHZ7QV9fB6UuuhxxSMVzkj0wzN+5YlvfMyx4ZOvRj
D/IWLZjRMrrFi/kw1nI4+xwUHQaQcbbyX30MqwfhhUft4+4FDsLF7yN1QcThu4wu
pGw7oCWG2WQBM6XCXBeq0DlLdS1w3DsjeuxH2ZLju1zITYIHB/84LhgztXSu6p35
7sdwGp6H7EWfb1If5LwrTgx2C3mvJ4j1HeEHPK+mGl1LLea9V1Q4W/P+Tvbacfss
Vn72lPB4vGhdkCMJLag2SHPYhbGpoQ70u1zlYICjRIvWeCxI15Rp5OdIeXMWEnUn
K2y9LhvKk63TwgGRgFPNBXsnQlyKdm8ENBQcOHl4F7g/gI7Cv8AmnPk2Pzi5t527
hNY9bcinyVkJDinOIihX/Ar9skJ3tJciDrysdZG03krOLL48sfjQzMA+MCaF6e2d
9Xbdu0+iUSt9KoG9juZznT3tbMx5gbkrTP4pA03JxQBJX+nNTRMVl9TQ/ALpxcGy
GTy19FW/i4aHg3lynfZx4mkrSXbwYFFX8GEjSis+CLxfBKptv8NsgTkC7ddlTxix
L1M3h0TGVUAJZcqt0fqCJN2pjP2tP3QVgleaQyhSNcx7r558N/HArJVViy3fXtF1
qeRPM0i7qNSC6Xz57Bbhi7WdOUHkAQ3cuixK/MGOVATAKvaJ47OLXX99q/LBfQ0j
ECPdweu0cS7Zmkzk/zPVjX7XG0XpDiL0dYyqpuT/+lH3m+fOALT2j4U2WY0ZLTro
l/H9CZm1sLqKfp0s3VCWLYISjcC6B3q03e7jo36Ldiqs0uSfGeeuQvMUFu/0HB0x
Wl8hfbjL6MsH0TvAS1pJcDBKabFuAVnT34up6AUXxtXUigMOC5rYUCLtr49q+Ju3
RO7O3/DEff6D6vCRGNJx7WSklSo82RUyrdeUHzuM98fNDdQxb1OhraxmkIIpx1OT
UQuHlaRDVQb7rIVYGBWWelYx3NVoE11RB/p6z/MGV1PbaBphUpHa7tFBgU9Ao+b0
cna62a6yQDVAJEkyJpNjYhgGxvjP7Bx9cUlZeQcEMWM8l0YDrh5hDxihF86Jo/j3
JZ48S5xIlvuIBdGrLJD+c2gM6R1namI1Yq7ef/bVXQtC3J81vWwE2h8OCjsWQA/G
YZt7626VJC7BOqLEnreNSpuRQYXN4nJ7Nf4F9VNT3iEvgptSUyYBHt0lj2D7hhuK
nksKW37x6tcbctH99dcSbmxjRAZs8yRwnp0Cmq9zUbV/QPAYiasgx8teXPmJghBU
yITck+ASLJxdCfqMI9R46ScT0iGYkwqZoQUWHcKUAmOCTHWyQnX2Xl1X+MFI4221
Zqmq5yglzFi4irBK5SE+3B/NJUPEP4mp5UqCFE9fMP4zFn18nntLE7W+eUTXku5N
Uxvq2rgdFEjHrN1NaA79NfOHMqWawzZnj5UUx8ijPTsoO56/NealOqMgQKXECkdD
l264WRfF8/RmuTlINyV2W3GFOeYTJF1auWso8Qb/gUmiJFiQswv3vNytXQTnCYyY
Y2at4NmFO1jLxldIO6U7kEY5Av2qQlm4Z4SJe+4Vlh+uy70BTvZhNs6WpAevOoKp
XiZPqLlDRYszY0kaCP3PveIdDN+0/IGsuUopNaKxPSeZzSxqq9adm51Eow/muGwh
cSgtBpeU81OkzlKyiSjIkscUgQEgKBWYLv5nZ6LpOb9b9Lhhhs3VVuwJg7afVM+h
X5B9LFZzabuBgzyUd0kscqgBb23OvqOdpbW7ucC/CWS4MpMKOIKWrPUrgSd0fbfm
EEAiZ8HbOzcrDoONZxybJfWW2P2h8NaengRw8v3JuNd8Tv06yctCmLOF2WqiXDuj
YBMqywS85JnqNgrKfH8WqV/1TOKhLQ9Mzpeuinx6TS3LXoC0Drep+vYE7VWdHkS0
jIFq4GY8wCGf48bW/ewM8LRECEgK/JFii3TqnULu8SPiUT0qkzsSUAnslnVNp3nZ
94lzPjE0bnDW+5gKKMvctHAhtfNEcGHwtPR3CAj5J2YOticgHhvhmBYj8KNjUNEr
Ge9BbwHfZTonr3Ia5Lac20ymnPtvClyclxrW4Cwrl8os1UD1BETukxhK2+aDdKnr
MOi1Igvg+ZOQ4aAZPIZDiDxKqHuSrZ/yANTniOkmFZPpGQ58kG+zbjFMJrrCoFFO
AEX56a3m0JJ2aMBTGhCOzKIs6+toRSP/kq8K5LApV9yJmgSh+S2Wt9JoyypFxNRf
0Emc4MsflDw9uUgFX9chC2fccSVZfcJGLv3INxyE0RlrzXpVujqtzZMLMo3/4md3
JgdwENNeXTXrmYod9q4k0grbN+G/XrThBXZJj43AxRyzeGiZzQRoYwXpsKVNvHUp
jJWwLZax5WFmNuGe4eq9rlOLcgVLRC7WmztpFcClvDJfM5UAYG18CY6nnsAzBubN
W85LTrAT6Fkt+F3IAgM3IT8dIfg0D37vRPMjPS1jNQ2pl4ZMmMWZ2GaoQ8sSVuBl
AdERfufQaZnF7pHLv0KNJj4ROiB/d5/hdLln4vlnYHnPH94vXJEKGrYzAStDunr5
ocG3COrxv8FsyqwZu2dGWDrLOg3lTUWeCq+BQQ+wkuknq+ysIYS0wF2t0a0egANh
dSlHp88olW/mgRURuYKT3VTCI85SJ04XdoClFfUbEd+219dne+8zQ5IaK0J+TTPw
LsJxDBf/xLx5d8MOxoupSxNjgOu+aowCSdhS1onuQdoxqnQt2FjKoyXBsAFk/6Wk
t7G3jNcMrlzuB6x47Cks1ZbxqKE25ss44vCFZzt4vl98N2g4GzgdDzRrfsfehG9S
t+k02HQeTh+3dDUTvuIE1A8ybiS7HEiu+/ktJG8FE+6XnwyeEYuBJX/rPxr5pOtp
h9Nduyy5JtO6ecV2uySIvs1UhhysLyCLe1YyTDe68YajKonIknYtaZJi/aBAKT8j
kjP5T0NEHv2s2zxvaQ4zJr2lvhU+b4P6OmnvxKtx14q2cnBtuIpxHi1NPsq+VSh0
ID6Es4JIBJC5LYNwHChhOAbpVJhGHsnhpJKQh/5f2M0FjzTO8sc2lD3wZg3qOmuY
Fvn2dNIsLvaxIQ5tm7ZgwYe2Z7OqDdDFZ/B5F8yIlAwGlnA7YrH1JU5FCq0wr46U
+iAS8fFhGHrwKOYrrkJLKktLCAf+d7qhJ6mHHg5VuchWJfQyZodqCsvfP1kCeYvm
ed88H7xGTSgb5t2/Qj1a67/dVDmzn98dj5uyMDozEVuGPU8UAk/Ledo+2FPtQ2p3
iRA3kSXcrInPwG1fXyqKmP2ikL/tRytegjcIGEHTOz/BoFGV4ONTDWYs0waLLBRQ
dL23t8JzVneCBiTMCdgPE54HL2LnosSz8gCc/iNNVBDFAh5VKDxFrdjTmbrwEa5T
eECxm15miutiuaT6w4QJx0K8dv/EgC3sH3DSZSe1msqtT9GVOBiRarVJ0PP2WZJw
HXkhAfcsAoYr9rjc2gFXkn74C0kWCZZXW5Le+pN7lnfECEPoR5A6eKVJ48rSCiuA
0Gn6GPPldyqOu8GLWQY5koocnDl43Sqif8tFizBHt5Kq9rx3yHo4em8RITLpM1gJ
2zN8HnE9guwl4okE82/rZGpbEmWml07xNekr51+sd3Jxrz6bCkpEr7eZsFH+2hBm
42Ki6GBYUHYao6ucR2QSRtu95jsyA8yyEoeRQj/GhD+K3A5ZZSr7VjsPESC/c5Gl
/WmqzwvbC0JIIqSsZF4JLQ6hF50pUTuoeSKVtUPMJE+17Yy0qpoCMzQQ3X0AnM88
CKDtDI+7pqQIU9U0E/25edYTPvj5YWASL4cnvavJfXOEtcDxpjsS+dlSoaY+xiKS
ylGEOvIB5Z+IPNS/nrRWeOY0uAWmZ0idnReWrpc5hc48wRJQ/7a2apsW7p2e3Jtl
KjxFxxa6IdwvTPQDc6zjVGqR6ZF5p2JdV1zrPgCMp0adaewdhXnE9w3UsYLq7YQx
MCDEjmiyBaDV9/K8yxzfE22ZVfD6aMr8Igfd0KNqVN8/Z1bCVORwPCjqCUt0/kIu
vk0qOhj0bRtsfy+eP5ZD4+9tHs7IDVIBfz/oc9Vx9JWwdhgLRA3FPR1t+hfJKvM8
fLAq7dFFes+07Cokw0zaZgBaiWUbQwaNCkHPh4d50GfPbKju0wtZl1ZA4o+hXxsb
+4CK26Ca8R/laOXV67LQqrnmnZho9eXU19J+M8O7nkSGgJekwBXi5Sr6eCkuRtLk
kA7ZGc4EeB42yYwSm64uPeulK8t5XbeslCQL3nZsW2MI1k+OF7Z1jV7JMJBO20Hp
nh5R3jqA0qVmvt6wXJpCYgdtYdu5xYZUO9p5riPqCjXtyI586qnxmd+MG7djtbyU
3qtZTiEB4NLMqEkdCXYsH1tSlhXIs/mJGmPYJNESVncrO1qR9k3J0r7iBFKv1gcQ
hCLZF43NyQ3wCSVfTvEZ9jTF3NIZybssybVMR8+6dHGnPxSXsIa7O4L05yYPDFUI
540b2RqRlR/4QkB5SEzDe9wJYWO6zYfsqpgtBhGaDHMymK3D98LnFc2jj9ZUhp3P
urru1UsnJPCE2RWNUbMwtrXtwRxGgYuJerRZ2L1CCUE7jKM/tW0i056ZXblrBKKg
WqL1h/8xQ5l21PaNawiFeWVxm+hIXLACxDs9/y5F8pPb3huu605BL+/IK8UJsALK
RxKjCaI3kkITpZUsMrjhqfWxkTEmB/INwyE59IXvkiafhoRgjFQ4C1dt4Kq0Wp35
XJ0NS/HlRHXSPPdKzqHbL/ErHZdm/N2e3hnI52GzwM5BIaeD86GVj0avOfksj2G2
2Gmon3E2YIKbV+ZBD9GFpjdwmArLecnpetyMM5GfSkoD8Nq48c/lYGyAOmJPw2Lo
0ZevZfAuwYFM2ADyce969uCDA8uQgaLogwukkdwqJvyMqSZhxMH3moY/Ct7SH7Eo
qnE7E5fsFp7ypezoTXOBz9et5O3yERFMrGlWzVPuknQ/A+/iHibu2aZCxhmgzt2e
7HgMU+U0rN/NR+MBBigm9IVBbJrapsVM8vvfjKon/1bQR4SQc4Y8ii0ARggAs5gu
7YAWFB/Sc10NvvnBABd0r9B0Q1sanx5GqZIAZVWMZZwuuOUHYwuJMTO1gedRQabh
PVWc1T1omsK12aZR2xmxDXniPF4hvnUwhKAXRhxm4PTJFZdvXng3U7wXg1O8qWpX
zBbm4hgU5Fu3PiYO6gUj3Hy9WoE/a355Au6z0J0WyB3J/oLxfoLKi2Q9Dyc7snCZ
knuYIvhrrl/FU/5Wu+nER4h7Ea9QzWgX7m7sJTsDbXilZsqBS188+dppETh42/xF
3gj5uxFpRcrPcgfUVLzOImmZ1pWdRhOqDzYd/6qzGkiAc2ns3c1KeYw7FkDg1Eby
V+YrQDxqGgq2Xe2oQLevhtcOg+QxFKXMwu4J60tSZkbZ1TYJXRg2bXzdMuPK9WIG
zit9zTfiK8nJGoNd1sucBWw2SxQ8WFEnIQsgAlJMn/Vkohnzd+mBA3wYy//Bpihz
J9oqZMv5khXqX0t9fCg0O4B+j32vMMaW0yHjaIK6/UTPNnkdnIf7fvtsXUAyneT0
fX12B3N2ea83qZiHkyomS7nMRLDSmjTvLwmHahIxmLKd6qA96BfSKFObaw2p4n3t
XZHTa3nDa39/SPtHdP5lpzM6o1QoD6JWMI1r0b/90N1yC85IC0L6SuS/cZx3uH2C
OR8DRqvAv4o/doP59I62lR4Zd9OlRKDwUYpHAqti9ohF+KZ/h0XLdu8KI4DR5Eog
cJ9KqGQSwAGLI1UYvENGzFuI7o97c/WDsotp5ZHv/n/HwO5gvEb0IgEZTBXKptfC
H+SaLzBqVJdXk0ZJQY5Wj+LszI1aTwbhQzBdFLKegD8VRjoUYPZ/KHCHXBlkGJbv
NxaswjsEtDccGJBj5xlPqSunedKGh3/MZeleGYtydNz1vzqLQStLS/rLM8Pc4R9m
bloGyFPCizUZyg8bvsfQHTiI7RNk3VHF8Niy6STfaNKhjS+XTOe7K0a378jXJS/A
SXa7eCDsfp4gzDotmyyDg+mfkXaWdZjRkZToB5u3RpPBMRnl044q5aHnfydh3e7Z
PvrcXsPMrCHFJ2nq4eGB2GA3yKVE7MYlDePfmYKpuMsLSX1C1vg5dS0JUTTE4AsY
9K9DMFqnrenegnmjnG0cQ5s9avog10k4XbGHMnB/qnwAXURlhwCBhHR4/5o9eUkO
URQJNWG8cuTjl9VBGQNadK2VZStLAwcJByBudvMn3TiUNBekNTFuDNpqf0rdYou4
f8s/MQTR8v7Deh9HbyJXgcsXv1aTjRd1aAjCDU80yPNxwHKsJbZFJlbkUwCuE5ic
kMCVrv8f9WIWDRJiMqckYLOgf2tgE7Yy5XIHOkN+hLqoVbZV2taAUoDyP61avr1l
BgKPVqCUQXqho6fUqYEB6go65wLR4tXPZv6GAKVY8fdy4cOxoOiUxPyyN/RPEOnS
oNvdZE0kCAnJdAsveHtuxMM/AbrtEYu4ku2J/7HtZ8aEFFZoghGYeIs+Ufp0ETPZ
aQ6SK2roJLZP3F59P1k1r4nQ0nCmmBGEameZ46pOOULa0fjqIOXfmvIdbhxuv67l
EUMjTDzpxtDDg3MOxfbVxepDGd8eSf8isisJAApzJbtnUZBtTLNYCDlKp6lLBJs/
LOh2rh19kJsxSEuEiVlxxdBX8OFZbRFHjdADwleKqTKo0plmvg0NeP/S0p5H7NA3
0ykZ+IFfnJTsJwkle6v80v7jdazIOUNtLtwnA+wBTw3tt1JE+y9tGLGiRzVBacok
FVzCLtt8qEEpPQT7tqw5fb8v/peM0e/l8PJertw8A1Kc11ha+aXJJYqY0ssW3YFA
vKWaqZTM7D6foKRBq4i3slXGBtVqEkRVI8NZvk0g/7rYuPREx6frOFWpk58YLyzZ
kjQfD1dKldTi4Wb6o6nBtWicg1niFp2tU8JGxSvuC2wEntKv32QRf0uxjhNMf079
UEKKp00RWOFFLt7YZcUmfRAwutdW7WeSv6toVhT7Wc+Blh6enbQIsDvJcqgVhxss
s8/YZbyYQJUnoNwC0YrkM6lRFEeGi/QcdY363h3kordHPcTc7rAomSpvbtNzXurs
aTJMfzZf6masKd9tKociyPgMwk7tf4l0BUxtCs/gXzTzkEuItrIHpDZ89uKThOED
3dZb1/ZZPZst7881Y+5wYVKB6zCfE+GSgPFucRGgmGdVvNrR6pYxsTj2IPiu/wl2
wE1ERGmYrZ8yVo71eov/SHFgvR2ENCLYHh8caqoDdhImJB4rCGkh+ANHGr1YsD01
lzRL4Pm91SRzpstC0KqgDI5j21O1pwvMEs9mr6vSwPLBWtwFL/YjpVE+towzspVJ
mH/VAWtHm1DGi8BAwyaJMhclAzTNfJbZbnOrJpMrZkaxpG8ttSdGFhvLdP2Kvr78
+JiQLZwEn9V7213ZtZgSUfcf3pp7em35IkEATmdXCO29hkUeqjM9JIrZuaEUn7XQ
koIEnsToAxVxTXf2tK4b2qXc3usaDJ3wABfogEcKB/1nn7mWGuh1hEmDEsx2Lqiq
neVwuhXTC1ccBUdMbDHxZkD7OzZummWuSf6bgMh2WjahM1O9qdwJWQsF7aIKul1n
F5ySpCP6IqiWAEh0FhcztYjKWfhOQpWpGHZDeMvKRF1kBNZjOw9Zskk/05tFtQB3
uUmsTTaMcuQommfuU+sP+cL21lKnpNcOkRQ0fQR4CcVfPVJBpeH2PE1qQuztPTue
WLrXFPVHqmFhJPLz71KSH9HiVJQmjCsSDkLDNEUfgmbdncpH/DM33WbPJwn0ksFq
lHMKuu9Sf9yv8SkqMngi2Cb+mxYPETrqg/DcF8zCqir1wIBkUlmq1wQDMZ6BK+9y
T7sgQyDz4/Ii9IulDDvruFlml0TWZIo+k83/C78n3eQxNur8j1DilpLDfrZ7OJYl
PeeGr1A27E1Q8znRCZHufV1vV2yjHWygAw78Nilt3sPgBlR5c7qw/BrWKXDRjlcd
bdvF6ZRanyZoGnDUyzgv2Au2Ngm4XkzPVsjAbrkWuS4qRY1X76j8vbRn/bx7TnaX
mjOZKf6/+gD+J2c5inzpytsNZvf5YVs7niwp3S0i+WKyOPWj+29PR/quKQCKlisw
iSrknw99PkIL8l0+YOq1A+Y4m868bAUHNeFll0bx0bX7nEc4jRYd1Xyn38OXC3tb
hhSDOSJXut63gSSPE6pFAco/bH0N3FXBM+Th17CZb8dCLqFdMXr9FLnF7624sBze
YCk7woMitpoEmOSWkWvBESs3WQa8ghZl286MSR4bl744Andv22Zorc7hhk3L/Fb2
cbR2XfAJwTtyrZD4x7XsHIbq2XLJFjdzdD/dPffMJonn+t0acNERkX0LWtUm2m3z
U74eJE/HZLYh15Wb7G5gxPwCmv2YXcsQ1QNE30QWkvrdb01nCpbutJg7vZqKI4qe
huKGU3gKURtGaoALbAgGx5SdBsG7IFqC2DiSB17BMSVB4wVJ+ZK5sFMA44J5Mgia
t/8SiCqn3Sv9uEVJAwQp0CYeM9OEDjo3cAv4xZeJgRZvncuVjwWmJtJlAVt3SROF
EfqsK0p1uWMq/9F1JruMMnv3SBhBvzDSo2iClNY9Qc9KR2t1ScKUPoNOtwaL4WBZ
m4YV4I2yQIGygsx2vj7xNTkdT6kNEVQ38YNw21c7Ij797TymydbhLnDrGg5Ko7g2
P6JhUTpxhU2lj5WoQE43Egy6CqOhSQpJcjEwiJ4HQTQlr1c3xOfn7aPDb3lO5CRp
GwV22O8/1plHIjEIMO22jqrS625+9x6bIyS7CO/XyNh5/9fZE5gtUE3IpDFSaV1a
K7KAr4yirj7p7IBz5seK4XsrsKSt+rz7+Ml6s/OFN0CG/zdAxNpYbNYJ//WEfTFY
nUvVchptB1chvjqq731DX765TNQzI65xFIRrGaTD3wiYnOfgFRJJ/NXfnRYxnbKe
+YexI8YuCtZb+bq05FFimHZHyvRS/26DYRwAXg3/nomLUvuqHddZdpSHMkgruf0b
bqC0uf4sv9UxIOelf9nLWLm3fXuhCEiu0Jnsjon1Zd6riVPkgJMQf46uWQ3PFKgJ
LslS/1KEbxXpkKnEuijfPMiX4sNZxbz70Y0cpDFrTvWoSihUgblb8DaXIlljd242
lQsQ9XUOKFNAjMfyd8mxRng0S/Wg+6mJw6APiaS18LY2bkuEOM7BMfd8d20c1tKv
BQXX7S/0uIWOA6J9FiWDjvqLg0ZdRjC8Enh4DlNo6ZTSughmUzMO6DgaU5t0tO94
7WkZMLMVzrTRe0RIZ+koxnaLO+We4u4H1b76vnhkL2pE0KSsfEpfDBF58IATuFVK
EitXnf+sSEnD9weV1XXJXOKSMOq/Gh8D9bSOicIyxXsU4SjJ4OVksbFs4FSyI9Uh
5I0PMX5E05dicYVYsHb89L/kaG8/uu786gkeEK+8VmjYUfOeqTjWzhEg7UITKH7/
Bic1e6tFCsBuX8mv4GpgcYtnvIElXB3nW6N2Au37gyzncokAwYuWXKX9K3eLV8GZ
De4GrIqEObQx8T7Jy7XZf0tQWh80UZGi9RN6nji3vPv2hiaptrx3PsKv2S4KfaoF
hLobNe0LaNhr79Q+Xm9tlEm5jGG0OUYhgCTw+sm+CPrwrMh+V7QVVetCkPPzwv1t
Cm+WkJ7V58Cn4bb7MOTY9EVBlk20pdcpUzaqmhlNFLwnd6OTyu4m3eFwzWEb8cdn
weYzzudcnvZEbbMLQgZHoqjGxSdjdTy6qgT3L2xwegQhlfpmraWrHox5dm3U0Qdb
vzMDQoPQBp0Jp+dy9kqoX0Ehlm816R/sq81QuGTgPuJWHi6MSKe5X89YMdCW6J8N
iemsTee70zDNM/34OBoXVnf+y7pyKK4//e1X/77yvZoPwu5cRWl5NbAvuxwRnhtk
zJgHCEDDWP9P89uFMNz8BdykmR13uAAvSp03MS4qnhFQkIQi+qLA5yAr0Zko9LjJ
gqzdgYr0CnXEaMdYXNP1WXpgWqamLs+Wxm7eWzL4a7JQ3zNRr2tHyuKWYItyV7a3
0PssKlGVaoH4dNjF7mZVBQwcx+khyFid7+n327gCD65Y72O1s9FIgXbhpsrJjq2f
Zb89sSQwnl+QNHT3lTZ/ST1ahqFn/hDnS6CH7GFb1eJKd4cW1raokLopwWHGh5Oy
3U/WLUUPoUQWqkXCpZhKTPDzkbsulhHDuVCebNSOPASOujzEy1SgDLUqfPGC79zz
+w2sOB9y8t0CasGPKBxy4xzk9ZzWm/DQ9F5ZwWlsQP2AelFLxPTn7AIXWpZ4rzBL
Z3pLE4KXC8wWh+tXB4ozuzzWningXDBKx41kH1eLhz5QOAH969yMnvHq8cUng9hj
3oF7iVv0oI598mJYp/xl8V7Nk8bQyG6TAJ8k29PijJ7SbtnpGE0IZxCVDz7nxI64
CH00B4iwfyziWYnVa5roj3+Bp7oD0HWznvJf23xmj7TeIRobz8Bsrx3UR7a/yvM/
gtLs4dyeZCHwefMzESgXT/VbB47QWo4j2SMyRdghp5AQPAFtDSP+0hf0BxT7R1hV
Hwi+lWM/IV13qpJ+Ph+lyajeeFzeAXwD6y1rtiukgEDpD2VRi9J+dahMbpsFtKFw
dpd1AKkBqtb5gHQPfZ7hBYhP46zsE0bdsYANC2Peq764WF6O5l8vhuQa6vdiZCy2
RO17xG/OWIGQNr9Bb4kU+Oc258xUMJpTy9k0Sx//51D0K+hmhL8shN4NpAMhJNuM
xhMivusIL9edUDDwSKp7oINXc++mzpV+PGYVtgz4C2BQxraXH4j40yGllX5b0Y7Z
Jhx/jXNPkTzhqIJjqGpruKnJQZJ6kuoTb6oohlPvpzkM5Z1mz1/pDKj3y2x5J/JE
Pl/spuBkJsytoX4WzmvMGTpwS8BFMM+bCY2w5vljygvBL7tfa6hGETBQUyK5PhXq
1Qs0d5mN1lTJpDzF7/Sv3c3rp/rHiUqWQ//mpNMqMn/N6HSKmUo2JcJVE7Q2vlDk
9boct7DvLBoWww9bipCw2iV5SR7Tot4Ai8M3SjvMjxNjHpN9+ZFIcD/LIuDfxTf+
Adlz+gbNycD9JGhxUKxGHjynNNfGO32/m/HOVD6VfqVdojj5Xhl79vqHSOr1OSow
naVQoxFOqvBqzXh7oYCkB/MtJnoxLhH7F0IuxEowzxYG8Km9DyTI9bC87jOBIyoF
+ZPGXGQlFW2hwpjk9wHTJ65bUPd0m0zzrBukN9zSYhxNhE/1SqVeOCapRMl+v4Up
4GH+9qxZQ2Mm7lbf2sY3obqWzHpInCb6ZMKr+QldrlXflCZfeXy+vnIID7d0WFPK
VtdFcn228LJoFKGV9HJOnOMFC7DooknfJQem19wcF7sVyFgEPl2HJtTAklI4zNjF
BUZ+1AGK74kvBZH4UveEpYYV9wE87lqLZ2GPARwKBfANl71NbV1gbaKE0pWrj2AV
WazJK71yC9IgbcA48d63kXD8uyAltLrpaKEzNuPqcrrH4/QaC+34f7M+ceHxDEWP
gMI1doXqw/KQ7LisxnIBRUV6ia8+9RFyD1+9o7c0shrvpFVUdrOLT2H2jUfOUzhN
ca0ZnBtS5FwHkHS7IoOLHiGf3V/UmJbO/QTwp04pk5h4ZP2ejwudYSDeh/bbN5yJ
vDMoOzbr1N9aoHgtHG39RN3vUZOsXVw64SSoEKoNvKGxXeXqUBVIHX+2JuxzYPbj
TY8qJY3krNMxwcOYyRJdVYHXfqoGs1Vgkgkgk1syDEww3BSPUyehMb7Sl0XG+yz7
N0fVPsCGCuO9yERJRs+nOxYCmi8Tv9/DIEBH6lRj73BsoN4rYTAAmpPfGFsFAIY6
E521bV0Cj/fHoYaYCjVH2A6qfUqrIpgphxiDa0VWWvPRbZLcc485wPtKXWQVaRXt
slweTNmySKcp3H7TGNc/wKZBdEsG+BE7AzxNtKR9BYInGXnqEVHpxp/AMpF5+cjg
z3MHQZPOJuveqeV5WSgvmV2UGKmEYZi+UBEk+eEkPdDs04qfz9CSouGjD1JVXbgm
83uo5ZO5CXBbG50ZSgUB9vQ8v3mPVCx7+w1pRLXFpkliddSmHfRXepWcSDKjg4au
+xsKnBNN08Dc7Juve3dfHsS5kvKkYxtSAI/r4uk0UHASm95ftVRfOPUeJ8R470rv
o6uhIxJLpJBK93PaSMXqifXnOKCLwTKGqZ2iK404WDsuByxKE/KEWBZY5wnM//OJ
fjA0soQb71aL1XNRbqw7phqIzbRL1YLUHMIlC92QT8MqMw1TaO1PRz6zLNwiPOCr
4fu20+uUjPEDfLBdqdzZftNmtCjh5PTaUUu8l5O5xf2+QlpYzDfmvk1FbacwFArj
qGtbozn9oHJcF6O0aV8MrVWI5wm0ttfJKJYLIyExt6evHH1tFdhdk+3WX22v8Fxe
B/AAtjF7ikMFIEZ1p1C396rD26zPyGf61RtaoAMAiI6xMHCkMZcnlzgScR2BBrt9
kqY203b+PJsKHmitH3fJazS84RLDtefgbkvKJFF3WFRZT/dlN9XGGuuzXBEE5WBA
a9iAqaYBt5igHBNOwMPMmGEXV6WgCBU66lJ/ncsf5DFj6P02BjCr3YkXGLvig/62
vFEKLtPT67SVndN1CrOgIvaRFOmc8pKZfsMixeW8fc/VRKgsC7B7DLHx3WvkyXJl
ZMSq42L8bzZs8BR/ZUprrMa2LvDABY9HrxY8Gug4z4FDdH2kMkJxxHRHTsINPF4A
0zl8LIUOwWGof0LAiVMgQUbmMJ3SmFo4F7B6Sq6FI73F3Nf79zHO/XBgfqavj1/d
oEAQ94IEcSbuGqOctbGdaORmDvPVO+zrtbtwXXh2Rc4k14mzSKaF2cAx+/+ZAdYR
GlKbiPH4JL2NVYn/3nTrolo3s6gYBT8doxibUCaKBSFk/IsufvXkYlsHf/sWBXcC
IsOHbGJuaGRnfekUuBvp/Cz7pnPuB8EbvCwAMecRzqMw1PHl86zQ4uLTmCNb79wW
EUWnHbg5BYW9yNQ/qpzl60R1asgaph+vFHpQM+jMCHzZlyBkhCZnHkOBqZK3K1zH
9m7Q/C/GRmE7evEq/t9RF9aB6kXBxmlJOktue9uRYChBHzWG5Xy6rjXWeJc2w+VG
F45dMJNVN9rBS3YBnG6oTSeXoDCxK3h9tj02eocWPt+HIYsnqs6hHZbT2cXHQTJq
y9/S9FHhJ+hUWydCTjAI0jkgB25b7wdh024t/KUUR8lbxxy2DYZLbVrqq8fyW+GC
Na7+Ck7H1w5LkPs7SAnaRdcXnXhxwEpy7FYGViLUV9bBI9yoOvLun7mfHzZ8/3p7
acTc+kSKq9uydjpo6n1eslpC5GKR/4/ll03rIlBv8JErcmxpMwCGvUna9+5PlzBG
JfpBe81zNeWBlZ3VA28RPk4NrmugwzNAO6AIGR/T+T4Xd0lYvwMaArRVD8YPGBaM
GlVLlyxyrZcesDYnHXQunf/cUoLD2U8QnOD8KdZTttjrPCeKD3EKDBH+/oUG4F7r
FY8Z+Ev0MiNGs2iHh2dNqBBzdv2fiJE+OfPjgaCr0PWu8nxI5tr0Ve19L5DM1JjW
dKtZl0Rb/Qp8qcA4gjGiprdsB2mMm0C0FQs7v682Hfp3AUeCrkCLf907y9ForO7V
ZE3DSM5AMIfkXJK7FXnbiR25p76BMwneeBSwYthOGQHUWfBJnux9oaSWuDW/hzwZ
Y3KaKcnZjCalR/c9tbKHtG9G6kpaX5HW52b19buqWx/nXp2bJFwKX2/Qs9Rhe2SB
ZFEXiTCNQLkUZhW9E+FNfZcMGaHI+EBpiEkqHFqVHP5x/q9yvTJ/WrNC6hNVyVOf
0GgOhbseqSRja03LR37GCz/P9jTcMZWuyAVc1RSKAagLv23Eul0WYJRmNqT3v7fL
UJplg25j0uRqVK2j1VK6XEQ3ObKDpvUY9nEprHr0VMOO8jU7ZxS5vmwe419rA479
lbi+WAzLkKbFX+/Sl8ITrnLHgLIcIPfUmig5FyVHfgwnIfIn+8onB7mrQ4zPlEMI
Ij23l8LJjlge6gq5TSQ5Jr2dTVz5cjjin5ETDzUl8xQYsEayMHwp0GAH00WNRj7Z
IxaCvF17IX+g/WfcHZbnw41053UYaLaKP9caw6jI3diafLjBQh5PHUoOFp/cH2tA
pk2TWXrsStalzgehVY+9IcAzLx8ylsk74o4IuuKo8eyUQaAhps3f/WrPubfNWt0z
XyUxFHiHAXl3knhMhiJSjoxyUBaSRzQUCR9Cnj90Nc1gHSbhYU5TByX78+1ZegwH
bM/D1Qvpw6T6tkC0BmiMn45jUCpJ+ze+3eeGP6rsHdRFb4iY+E7l8dM4s3Wt1bfY
DrqauPdLVUg5afZZLFijlWrvig5Z/PtKIMdLOLgQTRgpc1CLRdKLzIOFzBXRh7Sg
HlqvNCzJyGRWtgp0f4KVvGfGpFCE5Us2zVuIy+k5v8WwZ3qHniY1YVYz9zFsKvhq
hItkA1CgBmrf4TCke0S20u3+tpPuCDoKmKmuJ1GynxXg1UWgJTf3kgTXmSkkh/hR
/682ioKa/nUaT7pJrmqA/4+jySGC2vumLm5tDZsMspj4co3t4M/wYfvhOyb3qSaP
iYiOKsHQdWFmZNB+D02QZNxKTjyF/V9l2hwqX3bIJvS05etLdb+VaFKYFaIkErcN
sLezjMgZT77moRwf5Q3L13cUzrEIdBhzcnlPPMCoRUc0mVsmSH7XHvlJLC0odbWg
Sf+dmYMj+OtBMcbwwCnvp21h5qPYylZLI9EmHtw6LnBL/qmWVW5ElBP5uy3OupLK
sxPK1taxHAZZkkEm5TVxV1HATRxRJP4AT/ERpLv9taOxCSUDoCDlx8x6dvne59E6
SGXeFwGXK4osj4FCjhNnhMro+hHsP3n2APuhz9FswaZMGT9cQNkNBL7iUUp69SCz
p4KO2aAN6C8B1IUduwvKL3BZL6hNsu/9oQ4no6BY9kchRkxh+Wkk1Ej+xo/6IL2b
nU8/k7GCen0+1Ms6hGINBZuIwhOD/IAvfDXIWIAbzFbAtD81qEqyi+XHZcLX4DuB
S6Wb/AdQdmsIfNdxg+kEWXyq0wJxyYP6ajzvCiqB1C1PL5ql5DI9nuJtustiIBzZ
4j4JW2VG7yvTKMsC/yeYLFMZBTgEFul9oPSDlojQt0XeKW5kqaJzcQCeOXgzStXM
pMyGswi+GSfHYermIDCiUtBZ0WbtsyjVxSrWvFTljxoWdOetM+cAmb9UVlzCTZSw
6bMSPXyaM5vlylYFljWeW9RAWeOWWUJD9tSmX1AFLYo8o61HBIWRH3kWNcXZr8ax
0GAMfmD6DLAme54ako0xzIPYj0jPg4m+ZPOhPji2a7abr9iIPNNFR84MRsQIUImo
hVLa7HZMCr+41eyTm6LVFneTyCCENrpSDONBl4BrkQp/L6QTQvdF324zM5c0I/HG
LwQsv1rfVk9WqcVYt3mebb7GAqCdqvFkCzM83kjwa36A5QG30GPpdJOZKeGzMs2Q
yl6z4YY43akgIFL9uHMFv9mq9R6xd/v8ZPWPVladLMgo0oyvQNc8IynOxzSqpxCV
L3lfy665Rx/2qfhY6JV6ESVCtPFCJtGdEhJhRSf4F3Knb1bsU9YsdEtMLt8yx1Xf
S1AfaWxvPm3vZT0gVd8MvvYXMUlI4x3bWUoOf40VvWnOwet0XezBrzTz/xGPtnpa
U+Fu3sIUSfBxL46CkbegUXLAdXvpOKfwnW1IablyXeJEXJA+xwmVu0nFSFjEiP5N
LcvIiPYDFySjtw3I84CEsVne5lKy5WedXv/XaPUBAzeZPI7SfvMoMJejxBGLh7UG
IDDx7tFQEw4xanXEckyZvIcUyjNlDYUeyV8plHB2X7/phEFMIGVY5iLZsvRH+Al7
Paik1d7JZ4Ti2r4YT5MaPIBmvg7zmPJMcti5IIrW6ftd3ZBFgyXac9TdzT3D4izm
+EUkT2GXpIhOI1yCRpOhY4lfMQ1Xku1fs2Ojc7m/6PK/2JyJAsmXVrlAzYdl7JTZ
Q0ZlkLmtP/EGoqUhG/ZbSF6SNsLiU7K3TTSjUoJ9DrLxYW5nRI6zWrlbDlA6G3+G
Ow5JP6Kf47KSsoSlPiK6N8gy7U1ZGo+QjzPMM6rbFEVds94TMhCx1Jc0CZtUC4q+
X8Sy5z4c0hvGY5wN02W0D9chB1WcQotDaBFUM1yEuwXaq7stNZECN+a9gTbiAMMK
MbAy1TKauA7OodaJJQw6VZQt0Bdc377fd/iKJg2a0yNeLgF6DqvPh7brBXisOJib
5AEmsqRpXNvYvO8XzA/8z74pPeeXhFTKuHAKCvW8vBCLCsdzehiRe+22TDyuEd5k
gIEoCeGVYSg4Jb4SwY1PSmqgTdX/5jollL+q92m8cUvth0W5/vg+eaZyQGL9PXx6
lDeJCjGr9SYe4Ih3U2DZv1+sNY3rSlNVO37IhY0q4WhJfb9M/hNZ8AgRc2487xDn
iAtGeHMdJ0+qVYJ6PqIu0lnpcPRkfMmloj0CSsm4e9kTx0yeUxSwbd/RGDY2oh5h
vHCXay7VkU3zKZGf1WV9HNNFtL8/EM2GTLr80zAYHNO3rU90O+hbvSdqnpwPut56
3O8fKg8hMcjOriFuhAlFII1XYsLeVvOLSDdfec45BPCXzAWFq6EPxb81kG6G7Fme
oEcor91hTD2533OOyr2cguGt0S6O90xd6mH3ffif/KsPZvqNhqEz9oRtVHP+K0H5
HYIq6XiOH4coE23Mm8LdQf0xDeMoqWUaJQjp7DtIo+hX3Sj2BGy3gY/6hueCOcLp
ulsOOAfxiFzWw1dVG0SU6g+DREJNwlSWkkGa60A/3XCYIe1f4R6WeqgzWOuzhzGy
VONhiLR3PAWL8u2sD3NOUbx4Zik4TZPLUE1EYVE3Ucxe04m2YpbcD34J2eJOWFSV
jeBOFvQTihaO412IvYEI8G2nSHgHMU7I2vAbc7xOeGdoIOz0pEnFcv1RxzrOe4+9
NsoeW8OUciZBfKK2TWGg6HrNRf6rKRIoL6BqRBtS/yQrhHYNIZXoUDqciEihcQeR
rcYH2K+UoCwUGoEHzcFJmUlLw6P4ttutcA6HkBYn0Na2kucNKjRe+J4j4YZSqrmQ
VnULgjj3JCpv3EJQsJhDqWYAMNMbQohhWTqbUTIyZvMuhndbfP6AF5nOvfnKs3I5
PTaKkv7hyY/4BHjlD2N6TODsQKfqatxBD61qv7+85SZUvlPXsLC8aFIngsWyKqps
DopC5tDOMgAH1LmoKqh+T1OwEAjMiUzWtmnlbtnUXxvIS+37FoML/eiX+0aTdLeR
nx4gGyeeFT7zWu7JpL7UogdvuhGJrfr7yLltXek1lxvK5SfSYgyesuHQYlH5HhUX
9vGJDQQkBye3KtSQcM4/m5syBE9vxGX5ZXkDvIF48w4fcT4q81mJ3gYGLCL7jIo7
YoAilxPxTgMoxfbnEvs+NOHNFw267L2iozmJCLMKwNQ51rKnPKrIou/H2dqPUt/z
/oRHEN8A5MwIHXhIZdvp6zqvpjQLEcKeK2gXKtVpaC2ub0BFHA5HaQxj4WJ6rYmv
r1vV8C7UCwh45CaQHpadKZ3Fu08CYUjSKHWmvfK2pXxZ0O2w1MUMVuGqLzwDAfWf
7YLfqAtOSk2+8jH4Brx0VLZ48fchsYCJox2Eh2empHgIhBzoqdGzyuNVfoM63TLQ
qyQmLZJKcSfwhES4pa21lV5w59s5uJ9igf/YU5d/MZJ4usbE/6sv+TH6d1jqo0jq
uHm31cNdcc26LbXzgHDDbol2x2ZetXtVCz+6Gdp6hbifEmxRCXFOEm1a39GH7yB+
wOZNSW6RsKpeDrw/nyIAknwnb8YgFmDwpPBaHZeD7mWXbAUERShjmmd6fOOCEWZH
YiZV0Zt4YM2rdlZTdIDzy8CUtuFtFDTkPhqfyBrSh395MmzzNqCVrD/uO3MlA4II
M83IK3vjWNe5zGZR7CC2y7C8N/XWG3WdTo93L8pbjrrp8lEPReTv8OIIttl+GXRK
cAwJbNByMc44TieDFqTNPIBs9TIxCZqOhGdKcm6trKaXDuoFqRUbtNtW5hSQrUVa
5d3HEyxf8iXvGjGwwCEkfjmMbx6uEMVYGum0sP6m3bLJ7G1MB7xV6ZwV7QhQzedq
QC762VMbKzyBKDw/XHUOwSvZ4mdAVZfYlUFMI1SDhnPdYFP8Ievky2kbNcFccuHx
FylKv0UsCgo9fMOcWRV0Cl8UMTrp5h/P8myq6dapk8YoQdoHDSkQfM/eXoF3CjR0
Yc20bP+5ntpnezZT9GPzmex47KXW/xlbtys6r2vFGiGklPuZj66iIVtkLgVjfHLR
jwl0zj2o53C1Sw6E3hvgMt37Mnhg+O+11lF6uY5SXpMgrh3XKnGM1rbITmy2TUyq
k4paD3EpC4I6tN6k6v8lwWlCMmPffm44bA9fq4CoucukUx5zSMjoOUDISMVhtOZa
2l7D8ppVlflqwL1d+NhYEb6YvZObHfXjqvvDV1kLrzeW3OOMk026OFacvdekr3LA
fqdqIrw53Zeq42fIuemoS4j0fdOQxqP4NPgBRY6Dsl4RjVlY+/TZS+REyEMekohS
x6kuN7k1kwEyLJWooe2YxUbPji9evEhC/oYzeTvlWj+nC5Pp3i52p/Nof/dvhIaZ
XX2tRVXWixG32h5tgB1+2j0suMsWSEFRnc66aLys+yNblltWF3AXCMy5w0WzeY3W
8MZxMGcvmPAb77P6T1tJK8JQXzV/X8kgSSNGZfX9IGO4BwkFPjL/pGmaRn3eE7Jn
iQ16eFxQ84xWvNHZRDZHhL1Uyl41/L0JBJnGcqMasZgvf3vcLc+RUi+HO+Roxx98
y35nRD60XrVbSDA//CfeTLeUhLFfRfykdaPYLMxE1aHVnyHjGbqzoJ1YYvyC6eag
1ZC9sHKW5DDUcj4cfhuM1B8Pwy0Ieb0HRhS2gPmB/h38NxTCQANVtKjWjYgxhVMz
onjM+SGgkiGdpjSohK9sKuz6VrF8v+dCavTkIPq+W0LdqKYHvCtL8QxEPOIoqkb1
z4TWgpSwWzkIvA8RzDfhlJytpsF2KT496bhf0mANOKTh3JewVZf0nKlVZDFLBL+X
76smyxeDZ7Th5xu+a8aIR120ReCHUwWSfURiyQbBCplNxIPriaUNOkhtfo36wJwf
Z5tB9etQmlffGtfc2mSd3XZpieP8ZKxpUiPFGpcvzXgVOYKSjYwOyxgci2PJekQc
SFCYbtNYo/PQlgoLV6f4kPaExn6zWjTD/+1DPC6/mhsABt1QNM/hrcOd2OivKW7U
mN1aIoepXL1hdIrR/9nCdU4JnVm5vgYHw1G5d+6t6z57YReSuDpNxSooQD66Q7Mf
j4rEeigcSVwJVVidLtKIxzdTm2FQ4P1PeyFQgI/Q3xreqtidoZ4VWIa9Nev8nBt6
J32tfFSV8/enO3IJjgmy9IJVGFEf/lbrZc5mx4dmZodKhrw8ywAGF0kVEI79sW+a
thAXL2SmZHf5JO78N3/MRFkvA+TLa1gDXvsTZGGfCghBiDhdnkKtNWCB04Y3VUe/
hj4kevMqG+Ru5NSmQWKmB32KGp1NBmfB7IAlPKNZaYRR3NPOuYr43vhW9bddVyE3
Q+4enf9GvgJrpORMEvtiLh+PeiudETHl1lkPLbtrZpmlAbG0sTzqKA2fvw3AyBe7
2qGlssH4oALraJiJ9VLtIcalcz450pmjYNE+QgOwlqtMv47ZCeW55VDVwaaqUKyw
ehjcRhz7fMu6c6Lc6xnSBZ0umvUT5tz1H0RZ/rW9hKhe8o5Ji65R+CvuMCpjn0Hu
XffbyBeglugJAflGU09xWKJDq9rgLje9d1fZjZ8ILLQdHH7IxkigEGRMSDwofWXD
l5Zyc27deh0NwUilisujZk//LmQUmi+KeiWwp5MZGJ7pKfrENEshpO5fG+/DFNBX
nkZV44VCNIDulHKZj1sn5qLiUTDrIx1xmi+z00neSis8UktqnA72/xWtdUAoypNK
dQUX4QJf94SrOVAR/oBmE0URAc80hJT2JeI1zMR2WHpZikUV5FBIvuEj1l7JjNR4
+bWxzAHRhkKfhEtdS8ZA4ZEX6OCLds625DYs6GHRVRKs5gpf7YQLJspTWgL9IDQh
4ETRlTMbSlRQIHuoa7k8oULIo//kBOM9YvrmgSsUX5OjL5LQFGSIafLczTO6QIIf
MNC7LcNSY9RvvYkeN86deTsgmpck/WDJc/DfhkfoZNwd+GfXRR83Uf5Y8lvKPdHt
Q7DpaAFOB0EEAl7v5JmYPl6o9Y727pftgT/dzijUNQL1PHhrCZn72guhTZfMu9k2
n/Eci4xkfY2UTh2eSd/4TAziPrdb4l07TwgA7jAY1n1TLzMzjYVkIy7urWWL42wo
hS9Ovq8QxbIahE9p3TqXhZ42pm7KTi5243lambZiysAQtXmEo2+bu6HUkTqFNBK8
1ib5sY4GLM0DVUBr5iONm2qJZ/Z0F+R6V6HjwrxQ8h9LzWsXDFc9B5eVua0hkmvN
R720N75ArP9XuT1xvIahAZ3g1h4hvvugjI3I8enCJDi4/iNmzStBMG+GseN4YPch
sRmwOiZ7AfupNHepDsz+307qCOoztmSZsroHwYjoT81vcL+s5DCNyMpf0zumouig
GWgDH8SrM+JR/jIrcA1rcH8Z3i0VUvJ5kKzSp3x6sWcSq652LR6+rPsVzC5ZTNN1
5eQvGG9eZ9Yd2EHwQ/7UuXJ2G5SAW0bnI29fOe68skIYFCg1aWClJw5HXfpRWi8T
53bzF8iWN9FAO15DWq/rg0VSyPNjQxwmJ11z17HhT8fr2R6oDujmZ8nMP6AwC8/r
qrtG3yJerMUar/suT+afXJcwyJgnqY+5G7xWzfdgxUO9RaUytkeWZN33WHgDBPm9
zeQDPzPBKhOVzJ4GI7s/iii8sSz4nr/6JYv7i3mRYs0cVQYzAX5j6Kzb/G8Nwsf7
3bhLdWm2hE4eI7atWYBChAkCjDwnAoqEQTUSrqKxhXWoBJ8orP/Oi0HzmZE3f+1v
xXvLdcv/s/FGdNVmzIHCJaCLk9c+UUezokZhvJZFJolePNGzalfx960AH3mu7tH6
wvsVSm0bJi59seOOXRzRa6VA2RrukgL8C73g6B4qWNIh9k8cbxxdCs8C/zVTOhuQ
tI3mn7daSLwE26Cc/qNnhJgNnTq/ZQIYVA0wZvt/9zOh/ema81dZhbYM0E8V39g0
Tqe1RmMXe770/4f3jI12ZMBp3lcHKcoFbo4l11NCE/ZFjIcys0VkGQ5vQvIRSYqK
gX8bc5U62RcjiJUaq2ganl95pxDkDcE7kWsRtqGpXEOy6Db+Ph4LfRxX892rvA/t
HJpei1hhXC7paYiDlJ+U2szfbAVboXirzvJOVQl7CHN0RwWUPn1dNbVnXAUBqAle
21UOy8T6jwb/AgWqNlk6Ymfe6Rl5wkpD1M2pTDo0peBPC3vbwDrG/JVjpmTmP3zG
spALvLd9VVfnnvpdnQSpg1A9oZsmfkycjMWIK5fuD1FBGyIrVFJ5AgnTP6vzYDJr
gPB55h9RPkf7bmABhu7dnYQEBkTDH308uVO1xEnNygqt4RzZFnyjgZlUQ8/WIMDW
d1QIE/3g4BqASZIZIgVQ8f3uLw5HtN4hFkeBQiMLN6GVS4CZioqA9UXZOMDj0ErO
OWjkgS+NWOXHqwB1B0Vsa/f60FJleECmwDcG9VKumFVANJvQ38GAqF83SFC08wCI
yGuBgdlGpCsoGAhqZgVIMd3hAVZxcJVt+0ZgqNmg4u1T/BqVXDp1c1+UCOK7BTpp
4VexYUj6bhZsse/lzOenD58I2RtyT/ephVt4Qtv6Z41Fz+2cdjnw+BgeOfd7slaE
N5KS1657pQP6u5E81lBl9OGLe77NR0woYvlhcJAzk8mAvQzLqd5hTmXHBE6NMG57
vcqFR1B6nlyZBCKnViqu0VYNvAIWl5VCCH/i2J3yk4HHB9i+COwi/EF0iv7+apAt
XrKhFWN/2uzg6zQpEsxedE3BwqSUAgk60hSJDGfNjofUKDYrIk9JqmLHZyz8Mj9S
8QrBAVfFpFDNrmXWBIFQcU4WhBdgf7Sf8yVz+zlarxxDflrCPjn54YiOi1QQoPyX
YIGKl8mt4Z7IFaVlNewBVN8UgCzYCBf7HrDlIWTPyx3UN58FDP3s6+csGODExAAm
TPsPwlKgh+aKDFd20oOD8/3Vb24P6bD5ZKTV5GveU8jIuVXT+bqdmDLb0xuq2JBq
8ri23goyiSxd7VhVwXVq8WNVW7o5Z+djMlgw/HujdSxwh5Vbdb9jGDjXjAgheI01
ADsLmHnwHDzt3d8YR/R8kwm+BgdcSyJOaSv3/L4B9iOR8YqFxtZ3674veG6gr92k
Bu8yOyGjlwWcYx4qY43f2HAX0IUFz2PkjXPVVTYhj3j0rNqOWxvjiCuad0+hxWEF
t774VGqXLDFUxoMDQCWo9baxbeNro0klvoaYKgpQiDMoZ2l2i64Zz1ve0yt/cRkw
Wa1+Ao/e4I8NMfOaOVU/7zv2W9USmelR1GAzEcOaXMekceiVGag3lhFJ023Qb7PX
SXEebSfdpzc1/OCm+xUs5LCCdzOBTp37xM5NlmFpzjGHDvQiA9yCVgLm2Tn2Pff2
joCl1gCbMS0cDXvbUL6jm76GURB8UsHifeHH46LskDPq6CXXdHAxKjuvSAj51ZsA
z/NvRe4XDZTdjWQD+pPojJLQz0qKvrS4FnGSKIZlKFOQo3VTUBLj9xxxH6XKOBTp
PcnRQxGohoUynnXxQZXwixQHe0iy5rsfNhodKr+97VqnV5UabBpaPu+ymfHW1qns
0gtxVvXFTpFrOE6MsDJUQA3nt1ghg6RChEePmzLZxu8854QrI4fCz0W25k2WWjX6
N3+Mzh+9dVD74TNAJ2sFgrJVXO1gNiQfIuTrZXafohcHkm4+k9i/ZN4OrN03/Xbz
gO/8RIXGh5UU0SlOtvHkibk+N/sa6j3ez2hDGCnpaTLixVS6yLyhUXjfQURzKSIX
OWdgsL8lVME4q+lrKkR5xKA0yh2GcU5rXVT4Twh0wf2gx0q7r/J8Rz/kCOzjDsmY
+vhyGkLmnqW3ivCohBVkcJdGPuZPP+XUtFYppJAkOlpEdu65egcYeGFjbxXXtoVL
x5gaGXubvtXlcaQI5IJOVzMn19Jd3E4e5mu4/v35h0h8pdIOcpieCRQg1TmvTSFr
8dDSvWs6AJy6IbWiCxSSLpi2V14j7TrOaFY6jOlg+khGpHhcfOIOsXkjKlWPZCdi
aX0BRWuACjVUiWzXhT3/MFQqbzXykcUMnjyUhy9LZgPZ+YyqZAFvViOIji1CYBiL
eiI1xwc50dUMH5qpAzQDbHSTc8GqAv9Ib/HkjzN77T8TK8clqNsAoSuyK70ZXrjV
34g7ccGQB8ESfAD5a8d6s4G0jbSFq7QUfz2X/ig5693rtYgPjtblDg+AjEy+Vpsd
ao6zxAKpyU45OZQXaSV+t/oubncJgytVRKtAtvcEElmPQ2nGZ7fngSsCl0NLaytB
nmjG4LZTgCnWqZexQE4lDDSMrBGnLJnt02apbAcjomcXiZQi+nY0izXgNte5dh97
t5sPbU32HNOVD2uZxda9NrBLHxhzAjdTzkQ63nKTPuqX93d/97ILu7PXcuKCItqy
SAm4An1TKD90/OhMwkWzMtJbOZY+oZZSEEppfOw/QNl9cnCvOzcagM8BVzciJi25
Ti9VhQLovTgfjRSltekmLQlSrmkFx+EbxvEVOIju3B6PuSpboEg/5CsUp4lw5iEQ
6TAJAnEkhdnYl4qUREyF6KFhpWhmQtgfE8+BAC7wx+AG7LrCAiSfL1oDNup7c2dr
83YHS+tokg5agebpo4q7GEW5bRvi/zb/iuxcOTwr9kf3xEUrk0RAmHy4OCGrnfKU
c97lHrwFo0LthdCAJ2xy1T9Lz+ONayiUFCQiPnRIEREAYc8RV7chwo+Zf89vSPk4
C5KNpuovEuK+JkmuJOWgDuG7CWNWQYErAbX4LMljYPxVYY03vxZE64rSnSXnughc
hxVu2SQ6Rq5vKtybl7v0xypN6pWZX7RJcpdgou7kagkMTKTU7KigGJeI+PHockGM
LqBJBpgRwP1E9M/XEEd7ERF++SVcMpZF1h+h+auEOEDqYKu87shW/rAEaguePQaU
Ej21BcMS64nKsItAhndn7cfq1qgQcbfb4a95GrPFGPco4AkzbOqsL1GoJuxYE3Th
/xhfLxLdMGCiVZObcxDAPl8GjY/67rd1fC4NLDUUM0OTdMZCJZ9sbNsjLz8KNzpg
G59zRvVzDXcz8rlFpbVEQscLrwRGPxr1U8F8+m8lOuD1eiyE72g4kYIqdanGYY5z
VUNtr4gOdEsA/JsWQZoZj8mfLqeG/9B1G8d5vHMwucg/ys+zxTyLO2fSnakz2FPH
s9rHL/DKy22nI5nmQWbCmVZo06dVPN4bJFyYbVpzoXpHpk1eWhNCIK22KaIk3BwR
DqbkR961ZE9pOiS2ToLHexjfafN04JsJ7RwAJw3d/0INV17NemfL0H92b4o50UfM
jKuVzcgGrOTgmj138e5MPTzrFSJaXjqgu8Q2oozpZcTGg45z7JJH9N60URcnwOl/
gxey1lUuALMEv7Uhcb9X/SPtdWdBG4iuQ70rvlLZW2Nryth9OmwnwaswCWA6t6wa
ylhPYFnt8CC9cOb6u3PiqepYyTW8HXlEUGIV9QKzblosReTW022u6z5mlYHdRkGU
XDcOzyu5mx1vrd0rGwoyuuaikT8dZE01ES2GdfIuXwtrBzT2jXIkVq+JpXa+upyk
5rHO50i7mW2M/ToxIJR9d0czu8vSb8CcoJnR/FzfmwVRWQzFrgYPTPmTDUKlcvwr
zq5M+RUvZFqWYyfFRVY6s8/x8ykO9jdAiJJhkkcpBwzv0B8X7WRQXK7YRg/Ts8aM
BBQgMbbOZtfmtxoEMst3TS7nb/4YiiDRkgMRRQELIoeujQbXQ12UoXOoRGp0UInu
epbK4iTZ5PHbYM0WZ4A/WTYqv1qOsn8OxcDNAmQGKE6zq3KcbUJc88JC19bMHJCb
emrdIUumOunP1UoMi+PRUxwpB0HHKmHq4aAyee5s2KYbw6r8SiHB45xxtLpWuJzm
AcSffB+O7zqT/AjZ4YXnpBZMXFQe42epWzduyW6L5wuBTxaCoc26EhJhVoIyApRu
r1rbNur/c+5evEFP+jsmIZE419SFJ39jOab7VUO/mRe6RZLXoFycomh3muU78L1u
SMIKZ0Tr/QQqLiZ6OLjbH2s69CqEchFkx3gdyS0FQzBAdcMrxOmBPZSo/i/mzL7c
2+UR2oPUzAEq/9AUCmY0aWdCIuAVpw58nIFjDDzC1jxdlxiDs+kubu/gtYSHPOvH
qGcIPHsgwo7HCv779c3VKZOafUqjf4V1VjmR/0bWIAn5STeotRlayW8sB0aJWVX5
CIp6bTMGA+gukRaiFx+7+4K9SpH4Ab5lEbHnMzRTotxlfsQWLNvDeVu/XdBrfpzJ
jgtW1icTMmbJ2a89ebTUbBtlD3+yUJNOr7L89gGSJHBrj8yFS7pZbUlgTjiPOWMU
0Vk2RQny3BZjc/PofVJxGvEiPDgZdT2wlI2F6e3/k8QtTzeKsvfmzKruczovm17S
wc5p0X43+DiGCL2tvP0Xg5rwxQNRlz8lSg9lJ2ZE4A8Kj3NE8swV6q/vfOChz87c
GVTzOIDr+qUj0CVyiuPLpjpu0N/sA8H2E80A3o/O6LsuTfRtVjuNBN+RpSKvXvUU
fVAElLzKmMbR12RehQroD0B6wt3BbH+CIJVLK6IaW7IKSFe2xhayIE35vi72vJem
o1m9k2iwbi4JboWIVodZoV8nq88vH7wFRljW/QKTnQXBmTpSjVD0BpQ7OthvCdyE
RiFpcfALPXhYV34kHSmRvkvjPJtM8lfDNx8aScF+dLeZ3ZGGjTQ2rvpWLe3bEdm8
09oMonlKRo68kvAeEt80o2AiAqfKr7v2z2RRBcFK6vCGacmmOBDwaMNhLmmU9K7W
NZBkT+uKg5sVmYYSG7n8bH8o99ezfKbVKoZKhSdQMS/TXfd/TILkRSALywREiS7S
ohpU3sOICsVZs9/Yd2xxjFKsRdc4k8BDgtNHLqQLe/ldTjONPInwS1GALSTed6cf
xLY8s5njUhjCPt/TCtnFRtUmNQDp7JMBUX9QJ16sLYCS7cosgebSQBTKEjhBQzn/
FltlWsyGUN1y41x67VLseJjQYGXdhdZdc6emE7g5ybi5qs+Lc0PgVbO8NBqaaLMW
vAUt58HXHHF2RucUweb9r79pflaGAGqMiB+owYIJHDrjILUPXEXVLZf6gGsTJWS+
u82FcRovgxhIk1VRMSRT9u5aXCtqF1aT8qslh2rNSi1lfdcNMMS/oCuUcmy9CuND
zCSS+ARlfmp0rKyiBg3udaCTyCDYyhH+GyYwcvrjMJ2Km82oE79a6ksgEk6kqd1p
8uJWYjufVqRUqEoVKGTf2QG59zb0WHjLDVterU2HqlhBMkRWV+246rroSDPjeyri
U3oCbgGoLCYOYK0ztUwo137BhOYA0FRf8Bj6Iu3kIG53onQ06LoIjcVAgZZe6ZEd
2Q8dqae1RA44bw9Xe5ZP9s3pBBpU0FHK3mabw4mqIzdetDark+Xlg2Cb9GSEWbip
cg7ujb3YE3gQ9IkPxGDF50lN4Da7U0T4Ji0GZmqPsDKQF2yWnafC1FT4wtIu4D9b
XA7p9NKsFX9V5jpmdLxHk2xeEHQovxI8gKv3ealXYmZsK0PgA7MFjfjvvWWgnEuZ
qUsARIs8pUUq0/xAsL5vUi0zSnJvYY+7gmy6byVHIxU0t0Y8BYzxhHxXXQ3/OQsz
8z0FuW6cN6rKh8lVcEgLQHlmmSvz/YpKFYrUj3jXZ3VtAJpI/JUopqJ+gkFa7wgU
F2iAlxBElZXYjZQFzG6r4vIySUa4LsEfqDKHzhh0VVdAHS4CeEvyAk42yaBY9kh3
/Kk0385LmOnRA64g19Z7z0Twj9E5gS4dSX86WELoeiN2ZBrptpuv3SIGy7enOg8q
zgZji6b5wCitwtnYExh8gOZOjOqqPe7YCZ8h2pyejtsMfAd5fTPyZHxpTguRJOxS
H1tqHtiO5a9UxgtspV1WK2qUB/P/Q+IkvIz/rMZigvY+eDtvgK6r3rvrRkJ3e5SZ
c70ZoCLtLmRrnWriTYxDAStIYFpDQsCHkx0bl4dEK67euseHc4sHv3Bpo99rdOc8
Qn8pt+gwmScSop/QUhlBBfzXUsO8fwCkapURuJwEhuRYrEmI4eac9Ta0Qqe0GhWx
AxVFhMiJa+a4dFSo/U/M0vUmEUyW3WWSSYbPWuRyTcf2uCcsmfocQiof+sjBfcSh
JWftsV7rCmIsUMWaWecIMatEeCIsw2a7c2DbeCD9gkiDHg5SNwei7cM9LL6s81CV
39qorzUOaI2KHi41ypN28kYkkUqctNW30+u9oVHA5KkguS/i9LdeCZw44vYjdq36
XoARy+wJpV+fXnshnRhcXiQYxmymk+3HMfSTRr2LFxCgA/UCfLzmrKohufBw8Lua
sFNEuu1Ll4U61feqjFwaNUPHI1JntCGYFQ7t6/sh0ZN3UWEvqcxUIOPmQ1vYrBzh
HfWMBCdNyt/D+U9Jizqx9ex9HAoHqz59SpGkARwHVh8nXIqx3q3MUYoPjVQ6HIsL
uk5ljk+EBswLJR5PkTwf+5/DlLdUHrU/dutQ6GWJNcEPd77lizYliv3R2RCZzp7H
/DqbZNx5GhsU+kxRooV9dScYFd1DixrF4573xCYgoa/VKSTp6P/MsqhYE97TZdtn
cA9/ir1PM4xoy1CTY4A0L/MR1gr2s67P2TJ44C/AW0IW8htGBikQsnnhwIGPt+sS
oZD9YuIXseuOl22nhaZJDuXiTU4J1IO+MFR4lWkrNepjYzSL9y8J9CpWHluawvCS
SdPOm6OOCTn3zFwmx6Nv6rSj6XZiQvL2nAiV7l0aV1zY+acVIO2JFjJLXQn/x/tx
5W1TrJdksRnNDdMY68XM2sa7JnHeSKJyXlnyt4g1lJb9CGyrLXMxY66jTM3R2ZL2
lBQS+EZzljACNLcBFM7tIEK4JwiVElRuSY825EW/gwb/xJRd9BaZ4EfkFGoQP4Zz
2OYXfBWcwilneTLUyiIy+SANIsiQMS8eMB6MJi330wTbS0QVLLQ6zguf5VyugTNS
ggJvVU1wxg9zx0EUQyiDlL1Xx3fpR3Ti/D7zjVH5F3zY3fBzJZUIr0Xvg8RqJ+pz
7VISU9qGQLKwEk4eV3sOz4phuThMD2oiGqYCDpp5QcgKVYW3ngozpqP5xSmlnBXV
SuGoyMoi4XkwHwSgy2e5uIcaSnBZCigPX9zevN8lP17/68nrv1JKsHY68o8cO8m6
beFKnIJfWEElS56IB8BupQ1wnC1y63Q2Ulxx5BnKhyDumInzKpsllTsmI2NxpMrx
Su05P9HYYLq9gO95qFg9j20JJtvA/0BBdYYWfPrP1FdWMAWUF8IYmC3skgNgVM00
L+u+mf9ru6Msv+H9H3j//zVOI97Yf/bOOsmUQWELDMlsQ5iHq/5k2xuBWSx9r9L6
6TGq3PSj/JLzVxRgR5D/7Obz9Hb8J5k95gkBDIq/aWe9p2iezG2y8F6rSG4t2WvU
zNuJl8zCfqIDuZjclPQ9T0pRNFS/jzzj2ieB+LaWS82kxsBiWAXkIvk8/ZQYdaiy
LHGpVloQ0oRe+yr0ANihEHw8nCzuUThNWWVZdTrCcaS4B78biZS3hd0v9uuHDEO0
/GYUt9UYgdFQz9I3zuJGIWFOaKdwzCWkJKaN9a2qJhVNevQ4VNcDtm7epOyGQDGi
LsukgUmy/S+YDu80tcx6oZ3zfacYW7RDlXA2QWm0uW+XxEUYvVa/1l8ouzOtjOCr
KlTYJR6PnmcFUKks2KX0sQsAgtu1PmKGklO0q/KoQDkKoL9rXCX565lO+FyTnLDQ
qmLGx91gBz95/PtaG9VaRyQBKpZNGxRFAyX088SMpYbsbFSYxHHZD/gtoV/yuOcP
vqducQZj8PBaNxeDfuCHkPSnMBjG3w6TKq0pFjTGZx1mOBVLWUkiVcTLQDTy+h04
RPB4thu9CWzSRnTkF8YKbWR1/SO8qem9u9p04tgSLnZchXYizjfyM1ibGEEO99XU
LDUIGAVQUXroibpVp6OnqJm0YSaC8E7AAkLdpTOx8cjgwgYlDlMuyb/Jv5UZXksP
rNT/dL6qt8iwOJleJqdoMZxz20NYXMPisJDY5ThiY0Xm7N5vkisKksYyI43loBtG
9HxQ3kan2QzhFk7D6vHYPrxPhCx5Bl8Vl2SPF2rGdfuzPCAO4K7jGKXVDGTMq6HR
sO1nHGwKAtQImeUnhZe5k70m/+gAb3oTtBfPSKlN/xRKdvLjiflVo4aU0vIKf5Jf
kFolvQIfsh4q9iI7LQc2D6NWaSnoypVrRhXqG64SQvYMPF3/7NNskrDpiGTVuTQ/
QLI4PQvUDvweJhFyikV0MHrj0k4tXuU/I00H8YxG4WwibYUOEZl7KJ8c7kYw+w1M
fwcY7Q4KOMvt9IvNxvKTDBth9ExeMNqWpgbs9LRVhKJ8jablIQ+Nq0Li++8M/vM0
0PcS2bUu3FDqDUJsOZYFyBU1OWICTJDo8jB7hqETRTUcOmDi+AQzztWt523Mj4O5
/yMkWd44gz3By3NotNhznnyZbrUINLk5sxjCNv5nw3UZDm9QVNoDtD/IhaIFAdPM
Lc+NlfPjXy+2ZDrErPhxbulPdtDHuF/aMce9GNoW+oF/6ttNjd62N0ZESbn0EinI
lpXfvgfcrZNUzUDmA2MjWRBWrtt+lngfKLlrztLn1WYMYJ8wR7lS6tpH2ad0bB2A
LVdmFkH9m1C/P/V3/GUMIsLhk9kk56KsIr8/PEkagim0y7VEkimeoYm/h9z1FP8p
ONBXdl4C+2ibr1Hq8AaLBcLmtQEF5uKkd4ip6sFfVovVeoXWpLWOdbU6Xg/Gl6Xf
FLn1emVSYSU3UpiAMm3Hgeu0INpLTZuQV6YrmosypzKm5Ny06Vcthjja5KSNw11u
WbxU1W0AppthgTGzxaywJ2YI/hn09h5u5sG6d2mwkpGNUHbyRXF/gFC0auyVAs68
AAGccKUOwoHDqlIzlWaXkSYmDl/Ky5NJ7FPRi4S7hg9fzig1n5whXqI3JCZ6aiai
VQVbwYJiUwhp4JGS1UOUlnterv8Pn2/JnCk3e9MsCuoqhGCe7UlYxxvTjzJWh0pK
ziohZuhRvXXSxruigtBYkT3QboSgAZM0crjNtZpuaaqzI90CIgunsf78LAhUqz3p
BJi6D69omppMJjpG+FcGsXGcbeav2c9k33WhT2OEOOoUWc01czAC5KQkyauKd6RP
17KcuOy/33AF3HfZxZsMFaYvjByYiix7m7OMHhYu9OLwCRG2MMCJ5yL8jMKomb2O
n94g3Iw9qTsdEvioxp6wrXIi9jJxfV2mrYNDd6dJ1fnmbboCMYbw6BXFdMxtNJCC
PZhEgjHhOogipRa9e6WWLG2b8r/zk7rtKZM+QHCqvCBDTlfprhMQ/EEBUQjUUpdJ
0AglbJ1IF5OzNEIz60Pbfmo2EoWmR2oiGEwClBTRCdstMwpYFMghxS58pDtZVm7C
Iitm2PAFOnqVW0coHB/t09foXRUbB6p1f2z5a9GJ+QR1ACENg/oHdJHMKC5scK8O
1MP1AK8NGXnIcTkRhRywMczr7Bt8JlJN9TuUbfHfdG+QeRXR+66o8pBRjCatesvM
QGGFqVJIQE5d/5skynC5lNuJOqkYvpYm9dSJeHMFK0a126Qrnc5do8yqyGjsr0z0
nlnTyEDWad/s9SH2g3J9m2IBFtMfwd+OHS7wymvnnbkwroEO9Pp4T6BZ1dvgP92R
KOYr+RTpMK6vocPm815hU2EqpIOnruzBIzCzqoufUiTCdGbDOuH6z8L019Az3gEY
hfti9lwS7Vm4HB4l62+dcRKhiAmbOHxUXkFZPqsR75WgsjHYLOUipw9Rjj9A6Qd5
T3qyYLHk/lxxYC18I9DnKFuAmRcy7dLCk8Ecbs/AnHZGrdiILIIs4+N0RmusN9Kv
JwDKhc0slcH/1gUz1JV2RGEj3xaYKv5rwIdEIFBmJaamQ3MyDDKvrP4eUzD9fbp4
q7I5NU0RAs6gSQ4M8WVwqElxSGUsNEneVYCrHRutuCVYjzZdjQ+7XczGPSl/9SaZ
7/P+d/e17iQMSnynqJAiuQU1njPnuPm3SvFMaQDevJVVvZfdk+uaqECzzTfmgSaw
N+bn/416OB3k+2o3vxORkhk9MYDBzjGsUc3Xo5slchzc/F+WFUaHnLPCfvx9JcFh
wVpD4XD3QI9HAq0v4Ne6JYYE4o915D3szSTqmRsEn96g/mKLhW1nSlmCWAwJScns
+sQCFdaJ4zP8UtlsVF/dKNvl+yCKU4uB1UltY7TFJrQGHJGury7u7FQNX7LMrvOO
wozuMZn1KZNaum1T1B5Gq3JQmKiccglgaRWv5KQwaaz55s+qiMXs37MM6T8TRRft
1n6r7E/Uc2PS4lBSIwnkscdklWXOXtImwwyHSEq9MnkHhkDKY3rThRIIMRm0nGZ8
g85Pt/i3raSmRXhJgxG2PnC+I65474YO2HWKzTZ196snSA2Kvtm2LyoLSUV8n6Ro
l3hPx4qjGA29sZiZeGa0TPHuhZUkNd/B9FmyhRQHtMUSVeSY8lStH4uKWR4ANVSe
SNEYAuH6PfgVCbQxv0FxP5jac9dIKxXBLeLC5NGu+KgBQDsnlI2fViJqnUNgNBbo
uvyBVZk7xINH9uWtFy93kInCtlOJ8mHVyay23ut5j+rybSKMgvHJyyA2dk4+pmGx
ZmsNKGfQaYqlMcxj/8tcG9F3wqA81TvZGaiOxuFbKlnIJTBI4ccqArJnNI6HMcak
kaytDfi09vFPjeYy+icVagiqrwnynUAmf2QqqNj1WPXrZ69dwc9Q3oPZqiQb0qfS
BBuMHfnL03E1An2U9FkvtrePn703NItyM25Sh0UG+1ytUNPAhDxYl518Qv31oEp3
ZKypzVQG/tlA4AXaPm0dQqPf8oNMp9HIMLtbKgh5GWHerK8+St1bycH1Nz+17AIK
lnyWjm3Y3hoW0GCvgR8mG757Rmrapjoyj1ryjVmWZnmI8QH3K20M/HXs/GDMArBy
/Pq+Pelt2uwVlxjoRp+n9btjNa0slKqrynRA9Gb1PVTD5eDEBglVOMsfXUA3T++2
OHoO0wiaOoj5tTa/VQQPV4FE7J4MgHoMaib5CRRAdJayvPy7s9Ni78DbAtf99ppW
zyOLJQFwNOB24QlAZVf1aCkkt+ygurdMjUTeIb/ISVZQLUI6HmCxG4mm6Y/J2qMY
jPADjE4xleNsYk00If/u8AbpcOLrmRDmwdaTvSc7bVxLxHMK11cJ2A7nW7m5niIX
l4+DCaIeHSRcMBN/e/wEtyyvZ4MHiSr9LBprm9Osi77GsiGmnvJ7MIo3eD3oidhw
IC/pATZPyJ/DyerZCagu62Rtw05iJakhtyrIyLUa0zcGo+Jy3deC5yQj4vhaHdE3
u0hwFouiD/UsQAMwZJBk3cmm4Woc0NOBjigeqoJOXui0uu/GuLxMcObtQbUYt/br
Cgg1Cr1uQFTCb+Vtn1i5oaT1WG1thZ1cluhqUKRad4KkJl3eVI+DxqtPF1SotP7V
/6sAFTvA+nMRTfggbQuJmag7/qSvzys+4gNcGnu6OyYbbausbOFwSEzir9obu9F5
wEx/8Mip635VgMIor6097VwV4rzXMTon53AOZjsNoJgWyB1ZbvNHxcoFcz2mdO30
VOBglxWV755xFyCWkeNivGgJAHLdOCIvNEhovQpXEHQP35I12MkF2mm2QOPxeB/Z
oN3SXFnoK0jIEeBbJOd/IVfM7l2d13oTO+xJ800+5m9ONW/H7AosjvW1WVV5X+Eu
rmlm08ieoBH6floDXzUJPXQ3ZyK9f9wc963VI/BHrl/R/6b2VLhCeV5oKdZZzoIA
CS6WEAKDKtZ3ztPBLWFs1imcEoFknVed6qLm76xh/zFyOEG7D7g5ElTGfIO2OZEN
Mtwg8mCwPGmpn6+ZUUWVaj06xh4doqN14PqqZ1yRer0fUVYaA6r4Z1Ob1NyAwm14
J3viBrPev1sXopdjrWp5uUYPsIyJKIgIOdI7FK0NwVAs3QoaGfvM86eD2dZKsLG3
Zs0ys/vpXWPV2HI+WIWbeiPKoKSWKsgYIlLrEoXn96bmR/KrktHADEq7iLuZXDcp
mSz1sxap1Nvl43i8WGj8Qb8Wc58fTsbS+eIZzvWlZgz/6PZ9BPUJjwXKNd0tPVG3
rbuLA2h+DwiYGF1s472+B+auLFqjOtWpulldjDfpCGI+CD1wRXodCTBDNyR4MqOO
xXTZcMULMm4pMj3eSOBbck0e7CRQOopfCeSEOE+mBd/wuKvsiYV7lMMYM3NRJjXX
M3EW8vr5BziTU1U4JXq3qOfsKONDZc+L/tgSWhgzPUL4pRzdcoZSMKPVtZZxOpf/
2E8ybKMrlQE5x6mfZdJ+bpxmV+/jFSrCe/Hjhyadk7fv6fqcmaMkv/1Yfv79zRj+
jJ3rFrFTCptsOFlUJwde5gEyEp5Ap2Q2jIkyKdESoWB2V2CoxPXVOZ8GSZHJer5r
dbl6QJR5ix7KX+1vFxycdI4igskHo/mQuORcyYL6svdL5wXW2grMEFry+ECTBcKP
3lYqkD/CvIigeYpyptv7gec4Yiyb3JsfvSvd95BlHSxla2I/RJ1gO3PyrmeaN6KN
7kCSuoXjKiQmYg08jGdGpw9bQhXG8XXXA1uI0ZqzBdqe4bIn1dntl1goc9hUTaa6
nmAdLrM+bHdP2/tboBziDvCTcphxc57E7YFmY0rcYxbFY6CFPfyobgofaTkuzClK
gQ83SAZOJS8SqPwBkJobVXAfJlF+jnF8jZIFZ94AqlMIO/8VtMrqdxeVa6winwFD
Uutfz/m0DEVHILjTKpizF6Xt+AsVEBNuAEH9u4kZNXlhITQB800jSEhWROIwHa+C
2X0o9qpkH92Kb/rk5GKi1T/G+s8xdSNzl61v3L4bo+BhZWTMsHDQ3S/cHOrVVrMq
0RAfFoeIudadyiwi+3KHwOY6T0N5UWg0DJu4KEFAGONW0yg2AU6ROsxCBVIlmgPV
uEBGTqXruVZJcEnLvc/zf1ChpgQi37TezcG4/h9IyMQdckY446sVMc7KySKglUWn
2GK3gzNSSDlqz39yort1hYyJCITgDAzgc3MduAeEUBRZmsIigkgEQVjGXjteAA7r
TFXzlMpkJN8soDAFMMczGDv/4ueYhsuO3HlKhVeglezAxsV5E663b+7IkOusT6R6
7FBmTXeBG38v065sX4bqLRcotign26WHrK9w4G7oGnliE482pqKyqgeFRsQ1WcFf
3mczJAJu2nZe2mCMGQcWwJfX2AKVxfSu+zkqUbxeS8jlvcvsmvtLp2B+4b1fQalo
snXbdF2cnVdSaQHy2XfFkI364dtgzL1LpHws2v9AZokTomeTHhfygnIoGVW8jRub
9Eu0ruMgaEi5+s9lXhourVaJmIE0vijdL4/CCv2ssAPNjxZUY0JPuDGUy7AJVnFT
BRiOc0Zjjq67p6lX649faVmbCQhsK55EHPOlh278POKstG1oNTGrGNAWgnCUr4Zm
Rb0lRy98hckPe+V/qbXS/0OoFWdY+DmcJMSqxEl1/bZiZ3PyK0/e8sAXbfHQshH8
RXP1CKGfyBeJ5J/5QmbpqGXXmyFe+eAAdv7g3DPyqGw0QJQu2Bd8DNIietrYGV4t
4Fd/eHJhvn4uH1CBlbQzaa1YJ41nrhRlwVmCa4kqBuiLCfy2wMLaVr4+Yewohj/D
2HMjMDDU6ldv/rdVP52utZXZ8FHGUFlcGPG4XSnLzS9ZK4puaq0NbPpRDAUUha/+
VmYJkruakQvGH9rLCiU5zGLcmd6vOb67vbLea9qa5g7tHX1XlTDeZUYCBQNNeOtZ
pc10ZqHvY3uHFfBMeIxbUxjmVWQnvex8eqnNRwDq6EKZH8ux2lddKFCHTeTn4hNw
AwJ0hZtgrzGej8K6RS98s50nuortyk4lkinbgWrWeOZ5ZBHX5doOr24gheJ+Ty7b
/kFpSA3FGMKJzbZBBjVcwCtq2ai7IkAVeQdY+h2yWcMJeXE4RaGzlbGFklS3/a+Z
BFFld3sLvabk09PqAsRf+QwSkbXb7k2cudLQvSNC1WMT6Oa5Cazfwo1C7L0amyIc
ZLRUQnkAJ5MsUO+AJWwa6e9pQm4DgTmIiLCygpbVx4tvUQhDLOwsriosF4QAe4UV
Kh4lbt+Uuhls2BsU81wOS39qKSAa5mUaSH0kveeiB8ej59BQfNJrAxQ7NSSCxkTp
eoGen9tXonZOgOFs9TgoEQooHS6b//EjgBUu8jc5Q7DDloBnPErxbbGAhP8L8GSg
DLBZNvclAEzoEzloCDTyARskar/6sgBCZqfETJ3F0oWwGuCU3pCkN48I2eW7Xr4g
NNpGe8yqU1jC3LV/wkG59xxwBtUvfkX+PUqo4DBOOhbrDQY31DR9tYGfmXoFnzES
dGYG3FT0n4H0kX2Sk3vHMLg3eh0qcPyvbk9OMmoI4pSH0RTyIxrXbCqVIB5X7B9g
HLjwsDUuDjOj0EP1NmdGLpCy/gjsHEWN/pKiGiUrOuLddx870xrjt5f4ix568kpv
Hv16YMfBJgbiteMLSUG0vaOgBSwzqLBbs1EVTSQtsdXi66VyzcwABB4sXDFHqaL9
9jvNsC6x44YW8W4+kfwrgbPv/Hzn9quzBbdbfIgd2V7btotvryIzvdBfuVjMSHy4
z15I9WbBkPNklGiZDCz8+QTS1WgHsVBSgofO2U0Ng4ImLZPOCdCmjkulCTc4NDph
k6NiZUKMjyM24essCBLFq4F70FHzt8+bj0ZP4lOX6nQtf7oN1hjIyxtN3OZGylcT
/hAE2SEgIOcymyBxSePyZDtPKWTefaIKQF6Gk07Elc3rL03V2aOewSahb6gJCcXU
9Ba3w9vsZf46KmcVBXVjeCGh8T6ZL2XPlAouaBEThrYKZQDfj30eWD5ljZD/hMTl
NpQvJqIHmj1GpLAyHWqGIIIryGLatATlXNJfkoDiEr3D9dq7Tf8K3PSy7VI0e7jP
EocQYkZEcQJkFkXPXFZTXNSBXW5k7xr4YBbVOxTcnsdMdtDgnV6vwnKq1XK4gnJF
94j21xjiWovnL8qqu8/OTW/7dGFogK8hH6C7vq3vb36ZuQKXTXVMJL+EpARUHPe6
F1oYUSAPBS1R4ZD6o3epzHskZgsLxmKPlFEihmoQluhDkoNc8umMPlc+oL3JIliZ
nhe1U/54I4LBIQZYZ/IPPkeIlUuq8Kd5F/J2qlmbkazTQcAyBPnBH5SG3EoMrBG5
xHR+nhNU7Pt6kEB51HFkMf4zuWn9vDBzY3v+icM097VD/bqTnZAoMRAu359NeRvH
uJndNJHXVHktKG5igNn9y9dMBR08tgfaKNxNzHFIFzbkadvECHuulC5p2qhoLl4i
++oDGtws9gZbEcRpbLPwHgmyPjEgJLj5FlXCMshWhE6sw9nOnJwsahMeUgfkaOih
VTZJLXQZgUAilav7im+kSAFdWNf3hSV67SP/diW/iBzbr5EM2iShcWZSm4kSealY
sbw0jVcjMzgo5fwnR1Rs88AJg5QjrQFWSHWC/ESLzl6CNLzqklju+pepWp9hW+fT
vWM4LNZn/7zfmRf1UwjWWEH1sE7hJRbA/mNkEKouj9JXrn24iE57QYgdnUc3lpGe
0j6YiDYlYKfWikrzDfJ/hx1+nmjnF8dScc82cr2O9auqZYSzkrH83M6earhS13zF
W3Sc+G1Yotzi9nsp/W7BubIYdId+roAQF/FOWbnlWIBYfzlhzVVSh7JNUMEFg3Q3
1Ct4fnJ7baptN/ZRBK7uKU6KVLwOcZU/Dku3+ip+HjTYwQtE11RspjH1N5fwxZ1s
3p5pXr8bsxcHRt8172qaoNRkcpcoUkNUttDuuKKldPZhzFsOJ9r+wqQX/AzJ+Rqj
1OWIR89ZcyFIQOsXsWfMiNeRyYoVuPENjuJGMSXX6cZzWsQTeZV3/RhWaX9D9+Vj
AGsgxOAW5VZkwScpcZ6XpoHOM0gBQ8tmPTMQnmZq7QJ5Bc7wtjFSe4Ipx9WNwITl
eomQyjNIgfBGD8Tmq5nuXOnHGoabkcBytr9S5kbU+dt5X75CFiF2IGNYEDTUrHpA
a0X7Szvz3yxoPTjdFUU80ULI5cxJ8FXcNzEcVnkpxf+xbFvH9GzvC6pkxbfX+4xn
b2NBvIxU0APgRC//ykmDcwlAlsQyp9stUCFx/Us1CgfTMdC/LeLwzO/nOm5inU7v
vjXXADDC6nkGNk2QJl1ZbA8/GS1bou4WlsOz3MSWxpqFfMGvl0I2jZmC3PpBw3vs
gUqkkDniaNvdKuKUKL8tW8CbZeCyNqEWb3kgCg9oDEhm7mG61Un1748Nq+2IRI14
B0lnR26Psc4lMKB81krDk8hLSOQzf7gJikxeuUIbB09lNFKJgS11u/CnC/hgytcs
iVE5ZOO8suZN1yS0hFg6SOwhZBc8rd71T92Y+OheCjQFVoNyWj3/ArT0EYLLPqja
Ogqp1Uq1c/y3IRiJe3pdilqVGZvQsvVfcffgpx++nEaXdhtwZBZo8q/fGKHZra72
UUggp/Smy7t2r2lGTWZiHSoawuGpINjiNMzy+U0e2pc8QpWssNUXp29EVssyH6hu
D3mOl8c3eAyZlpLDQGu4ZwBrgG1fACeh15/f1Uf9q0WYlCbW2sMnwKfqJmd6BGxk
irkCD3j4gFLAEdJn2y9I+kOz3ZB+eIJlsViL4Tutl15PFbZ1c9jjwfzhp2N7LTwQ
9HJgpHiNCPmQenagzz1VcOj2YPTZykjnUtTNwlJiZwuKCit4f5x+95rgxsaeNPQv
+4xs0kkOteU9dwDxpu3Zp6jLf75uE3+EPBzK9PAK/L4slOMGS457tn5pZ3fU5emb
WGw2hKG9E80RFQVGvRrgwIi4nnhUiBA9xdEB65w5xJ8xRQ1lF1zVZgC0sl4UEJuQ
2awXoO55n//NuleGrpWGVot1X7ZIs8f0/0F7lCx4JDCOxWKBkitV8H6y/yaF4lLY
RkI+V0B+4laLY/weQgffHwVmIOgX5XMV+DP02sCslaTkE4ADYioVXijdXxtfdK2B
blALsibhEcSgq1BOZjydACvG9dz3YzKiVo+stColji4a2kYn5eHFgsWrGjzlfanX
LEXpYKt4ZiLPVe8Z7SFHGGS2MUaQXa6bLGEhUFeU9n742SFUQXsha2tRaP15B4hD
JktpIu9FUdfcxVu/CarT2SDfVIIMEq5LdvCMvNwJQrEp6rfKM9j+WeK2VoB0j82U
6l0UFHAi2SO+GWNXLELp8dzl8vdpbnPDvlkfIHlWf6Irk7/RX3XPgNZ79ObKACS/
9NuMkJ/3AoFD7o96vOEFEPIBSSO/Yx4JTjhcFJsC5ABEykJTKA/8enkzmeqhXX9e
B8vBfhgZksUUcr/YHKu35WKWE2ns6GV5SI+EhNgJliUOiGfOApxLiXRSr5q6403j
NEFsJDZCeB7E7ruCVP5AkRCvu/Y2/70sIUa/9zkO8Dg+cjgSw70CvF+VYoaHedSV
Ti84n5u6pEQtp3IMiJNSK8gYURRHMAfoJh/IJ6Q4MbfhmUfAIdqYtsJQul43lVMC
FyV4PCUxEVC4EVYBtqLni4FAJJIzhC1LEfk5ukVa6G0cg3hvFSbuuZTurUe3QZ+7
9e7lFyZ8SPzX5OtpePzS3RXyQcyvoqqxhlmBIQNY1H5Yt1H8O3UbLuSDvG1qdJRJ
1JKry4k1Qh87LfBKByWq3QkEWL8CM/sHZKKk7jytaF3/l+bQ8nudc5z82dELiKCy
XHWgI1nWmYUWGiSk5+x8EoEcizX+Z/8DmO7nDvN3h62v04C/w8xJLywq3Sthwsud
Rhfdy1TCALiveehdMdS1h58JRCKJXkgtjxa6J4XPIRXHA1DWvDCmZ//Ad4d33+Hh
WcbPMEm3qjxDd9njK0rwLkYOSy9EQWaKDoxnQ2u0f6PsQ+a9JG6nx40ZjCNY75vr
Ook3LAni5NJhpRkZ5Us/EerIi+nTdyuKXYwyMoYV7dflU1aXKiMuUq4ZjimJdUKM
/Aa9cg4zgVU9gUT+VJ/F5rXRqLBbU0SYBDGqENVeo6UWEFt7/ShlLGFolQgvNG8Z
jnkAu2RjrSBvpxo0j29Bl+n0OAXQXMOxhI2KDWpUGneODTc3uUfoTqklWeANoT5L
BAo7TDJAiDOIBfjsU8UquELdcHGJjEc3b12MfksfrzSWZioJsTP0JXGt3HOHKPx5
6vkuPNxBrfjJbsiHYMpALdYcMjwftshzW0+DXIckHHxZOnYKxALhEreMZdFlRUhu
WDJ2ijm0L9fj1r2AZHvtPSjC47f9l1QfDmzzSvkCprBIOqg/4RgBgn0LEZBuaK7G
MYZ+Gq+9TXW8wEEiqtmEoceckBMFbT7NxxEWFFrdk53UtrIw/an2+ta3ElTaG7VZ
UordurPQOxVQfHT1RCoVnFn2v0+8YxfNSYnfIVr8bsqxmG+8ycx0EQBU3Jzw++Fy
21Wbd4DmfeClgbhqLHL4Xf1O0ijso847wgoiDtD/yXHon3xRu+wEVcjpXnD6wjno
ktyR5qBowLT8OkQQWpmepfWuuLbb3FItCySFE7t2gkzVKo3vX63nGacsSKVHzNY0
zYWqzHjpL/Alc/1sRD4VqVs7N+2fwchbJgcw8L0n/T2x7hbjKA1mvF59Us0/7cHr
PWjwtMk2h6pEtzKkVM73VnmmcpAyay30M1JbdoXigmHFSAGYB0aLsR8s7MoWOZUf
LlHPqFzlM5TjSG6mATDTrydeEfDPJTIrVPk3AxAow0aGJNAl0tPPI1ma9zt0+L9i
gKReAV06YApicJXc+7PLlcPqXu6jHqF8uVNFkaL1tTE8R8krReO9sexlYONZhSp8
zA0eF9krGcZlp9MfTm2PzY0CHcsKzFL7Rt/ow2FjvB9h+T6oARQbQG+jZAQc/0OI
LEt9JAEYDoYu7ajxiUukUU9arMn2DYufI2JPoMroJ8vOu5Kxgx6xLIk2M6kISyNZ
R+QKYbSdkn7tA4By1uZenjVc/yO4ssxABLYrX5dfRE67FP48dYV2zOjhmt/gtClY
U0kAnlJ+1qTBaZJlo3oOtoFM09nV5j4DtydK+qOeHbiOdV07OdlVFIQXiEsR3wTu
GGn/zrqGffSbd97fjGK/+bs8Dv/m8UTu/rdrdbiXwIxvq4lnMJ3rxPT/G0pf9yeV
qu8rI4xCToangN32fBYh1Z2hmHwtK1GzSVJOB41tlUD1hnpUQWjcUKjCABS6qrRy
qOSdoX1XJcqj5XiEY4kL21JjnaQgqLTOb1znlDGbvm/LD99s22nY6CkYmvwGG08n
sGgILQThqvNjUT69u/N+dFGT7RzUZQmGCB/f9X0pnkplLrufLPaFBW9FNS4zhQne
j5X4Dopl4PiCZfu13+mIvB2dfKq1kvFGHeqNXTMTZAZ8ZILNaprCov14lLbuN+YJ
mmlMKmg6CkdwvGjAKPF+B9GcocI5XnJ9YSbmZ60/taKgT2V9bUwUKbLniTDLI36N
2+cFpO3ngjru4s9WFDTo3lp8Y2Vozo5A2k7ziukMcwYeiPP5XcCgO8F1B23xQNXa
AIe/rnxPEkCKA5nYhEjC3D5IT91sPQMa2jiuvUMf6LSa6g3KjLAEqnwjLVR1+ohr
yAtejmHHzMfFCNT9NTHpP80JYHj+gxZwBAlcQb3CcXnr8H1SSvmlqZaNX9yY/Dav
+edDg3MnLh7x6cqthYcXdININd202hFRyfSsXkZVFAGhYEKao/S+GtqGUnW36VXh
806OL73o70JQWOdemd9ZNgNF9QFivedmr3UKN4nSHXSPRQ1hz4wnRduLYqKtQgmH
DN5W/ry9uOfsX02gZADKkAn8UoQKlKVUJYmDJYY4z0+G8Flasi5sGgJHT1oxP8PX
g26B99LbIVfsckGBkrHl+hlzcKA239V+4W44dDDDV94weYqusePh3CfX8EAcTnXK
CGhGoLDFRsxuR7929aCAzuzsNmdFDGL0NRuO9Ubei9g9RsKORcxol1Wom0O72NLg
c0rs6wR2GrhX1QE0pwPmo60f7Is2IC2THCwhTUipPER59jP8nkg4GU9E1wSDVChC
ZjDDE7Ba3+P/US7/D4sa+Nevyg3i5bqyGXEiQ3lvvka5oYbSNAtpno4H2odFfXEj
eCWDzksHW8Hfw33h3Tq34rbDjXHybP5D6dyL2i1WZx7lUSjyfPv1lCYxFXoClmrZ
oKVdQGr1umG5jOAEMX1wDSDZ0mIMUFGbnvPrAP+D+UqoVzkfbME1A+4YEGqDviJb
WdJnyM1TCxzfGJCOjfOPbXwiWzMidEn1hXYhTXxlSfCmJtXLq2yzskkGVibdaSEJ
lYWNF21gynOxluuecl17gPsYzufSp92bdSgtUCg5iX8VK/R5SHwxdaYclEdh90AQ
DfBoevwMV1diNWCslQX74YB91Qo6XRJa71mW/rzjN4UrJFfYdV+8GlEwZyFwSc9J
S3690YhET+q5zn1AN+/fvzVymGj8TCRUJd0CJxn0OBdHGYC9q2v38cyNOs2rwSTv
WC16EAYcd2WReh7tAQ2Gs4zv2LvQsadBMkq0027HrPbrEodGEY2UwAEqk8XIIEZ6
t43og3UIN8P3rnoEkMBHlYJwe0PSwYDxcXpI+GeuP6P6xjWG7PVf1yK5ZM37QP1z
IUgV90oAssy99iPfTBk6hicuo7mnH749fekBgvEUPeHueBleQxqsGR+fVhI2ruaA
zNJjM/c7t7PwQC3k4pZcLItp4FmLAmNGKLz3pwcaLaHOhz0PZ16wckMxhoNYCWly
Pau/dH/S0tJKnfqdcJCacB6jmc46c2i/qHzWo1WIBgTKuGVZed6bTNrnfQHYzwYz
52P18vMhn0aOhwXWcKkitDRtK1im7277w4MC0YXP5LHJrrukAfZPEFm+6DkPu+7j
v/pbKuwDAQVUte8I6QAWL3qU0ggUunSX0femPjL3iTmrfQp1nWS7ljz4Z5N0tbyS
nBwtrsjm3JUk9FZMG0n534uKGmy3Y7KkDXSLXCmpLdpnq+6Vg67ng2XcAaVCLn14
08BgL/rE9wscsXj9+5iy1OjFPgwWX63Czs8OLJKbtY+4rZ5xX3U79YKD8xdvPwxw
2Ui7ERN7+LQLFLVzyzYzGEfcWq4rJBfyKSMbpdlk327ftjtKiqgPCRU3aTrxT45g
nhGFu7bMV1raJDHqYYQ/bvFirzsYMjuARIEDcJwfmSYm3IMVtSwo4ySkRn7s2tui
xN/91oCW8MulkXTlCwZMKfz17hntLbsgTh5kZ8oYhwjxlg1SAjCn1u0eeGfXnPSK
Rzhcr+jNCXlEMU0W/wG0YatWcFa+2TZkt75mCDhCyPCupeyTHe80Q8nj0cBEanm6
kr09a+obgIJGEX8JEXVK3ukVgZ0QwPBtw/u3em0JH2GyFQF5Xg3idsYOvgcIZcZD
91pCp8EUp70cRbvvjrvfT2+jOj8hBSliR6jR5Hh7INEtJPUxK/8d7NZ0YbAcxPsR
OkAoTFed8KoCee1w9lgIzkZFT8qUnY7h624tvUjVuCaCdZQG0ji/lwQExKa/giTK
oo3Nx0deLYXugiZvDOedF0xe5OLw3SEeCa51DV132mfWpNg7u11jZvQShSaU24zv
+q6eJlXIj9hw4deYNZ7xRHoXuvh9mEQvu7iLittJkVoSygenTlbVVzWiX0t4+tm5
wdPKQREyeWMbKgMVNmw63YEwCm2uXbCzpsrLxCgNZuMZrfWrD5eOnmJDHhKeAhne
PyheYYk4ug3mVyB6SrTJk4zu+TTtpO9FKx3F1x+UsmMFcDFaCbpzg1u5AjlBSWS/
2+1ecMXx/er0teWmbRpZN2iAowMKNKd4tT331xdgXI13V59as0aWJw1EoF/A/fuC
4X1yp4gJpEB6k3/ypwkG/xBz1EBo0cfOYU/73wITETXpAZR3+UgzcgDXUPUKquJE
NiGNu4ZrChSA0VYTaK7Ig/SIjcfWudYyqG73v9i0KGHHhO6SERv6r4BPoWa72zJx
Q6fPBhvLRS5kdcU/wVZwF2gEYBc80HgLKLuup5lbYUsWfDWe7VT7ZUtevn8wttVo
TZMHnjWogpwxFXp+rzOwU5LJN6VnqKkhxBuJoVYkbbila4l1oKT8ia+JVdfvsxZ4
Z5ZQyHhgCimbbPMSpuLgzRblIncvThVI7iRJssHDLuJoeg8zMhAetY661M0Xujl8
wbx9oexWtL7HrgFgg8BD4nxlPy4dtkCEfQSWNsHjRgfoh46z1tUs+TMTEjeUo6Ut
gtfYKip8u+xDvrwjZR97rwK7v+PAMZ6y6DjIXrcD8vbGCrJcXdoPNcspX1X854xG
uKPQvP5YIai9mgSwpJsomYoH1UyzWU85sZeWBLxFdw/AHF48Iw2ehVzoh17/Cq1p
vNH1wHKrgZozZSImUzBZqArLiutnrXkB/8gD6IkS+a4kx6kWwD/1TtQUYSYPKT6c
UD9DNwNJ+l639U62N33NYjx6eidasD+GQy7fM899a6cg/ZZv/kFgChupscP9TXyt
suJdM1J6h2JT+Ajc69bgbpIKyRFA1r9dyt3Chsoaj+BcTWn0Q4s1kG/fHFeH6yVa
hdNW7ht9xoAKiZEyW+lvRRFIZ6SeF+EvVMFzrGLec3wOIAIbKk53c/AphHQiiE/5
v7uqcm33D+NtAmO4MusjbgKOa82nmCQlqlvzivmTVwIUC1wQpu9I55nk/Ll7K4BP
/rGJ+vRdJ2ic6FN/U9U91VcpVEb9c/WEtLoQuKZWkmQMhBjlTnjfCQFGoyg/qHDc
eZZwmgs4c2P+v70UwrEPe0LKr5bgpQIiuVVNGJmKajAiiPXzUSsol3u/vuZa9EYp
9RqxJvDYJ/5cmbvD5i9qqA6RLfahW9SxlB/z7FyP3CaojS0Zky4/WZOMW6fiUdqV
BT4rxU9c1KJDiq/i68oGelI0mzFiZZFn7jvyLCYU9R2ghaRLu2B5uCHnHTk11yk0
sYArjj8cHlfzs7rzYVjmcJOUfVhPdwqyGOldIxRPOB9hh4LLbdmAW34+1cv4RWpn
cezVuH8iutng1EmWi0InfUHDXbhnp6QWxuU9Tbl3riWf64/+coV6HR8hwfoS+AY9
FGj7dIJ28DTIfZ2nUtB15Jn8dAOWZn3UlX2tUVZ1habvte34yijlmFWEgq4ayZXV
y4n8Gnp4uvNyWM+yNqsA4h5iuXeRho1VCtoZjVAWUgvP4Y+yMJ1OaGkSZBOwqI4e
akBvuS73tIQBUX/BqUvf4TnoavAJAFVtrUvV8rcfaCf6/kwjr0eJG/TBVUrd/G0x
30KBcCx1RTBziT0/rwqUlMGMDIp+y+IdxgdVwhWlCVk8Mt5xtmV3Sme0KKhx0kJ/
AlDMZFCb0C3uxb1sk0sh7WlnA0TZePhn4EhHRW6jvfWx87q80T79rtVGOvQOH4mj
94RkB/g3iwBBanDekiM2+8c6MpxLpubHG4Y1pKMkg1MH6BXXtSa/zyODLP/e7D+B
uD7qIAmaNreLp3exZIpj0ldgr1EaewfT8sgUynHSNMt0OUNZbR0Q3FUUMjBc0XjD
NpibfdM9uOAk1TprgkFJAB3f7Ob2rr+ij/3oIyAZBF38SIBHdGbZz/llP0R4i95S
dFrXFW055hpIbAOJ6ZDDWjlMTfR9ViwtCUjD5KojukQp+EGW/n0cNx3rnW2T0dBD
s8VRLpF08z1VbYAvufZUyBnnDFdczKdhe+JsltxPPQiK7dcCZFZGzN9A81j3Jwxy
OVhAvBtuew3BNul04eFV8QfoVUUphJk1iC3qpd9OuoaA1+6ndj5fh83ATbqAWPAW
FbQI0k/Z3yVvXGSn2JiYM+eEMeKH01o6YMIucKAXLvc4pN+/MWO+hHuVS7oa5+ek
NufxfJcoqcTLii4HKQs210O+o4jND+61+4RvGgfMgTcj+LPUoDtK5EQUxp1pWEkS
u3rJ5i/Y0kwBC64BdGp05Gb3fC9MhlFDY40uCjYJft8Zf7HwE8E/OI61OhWqbeM0
DHF6MS06TPRxaft5ZDYml4CSfgkvHAU4MOP1L9o+u8wgzrA+b4uazmUqAJKxGG7p
QQndgWV26+hP1fTS2+Fdh0/d+7dsAFXkno9TiXptaSxYQzkfXfdTOtz5H0zIED3c
oBiA3sgETRorgnNIH97KresOZapWGwqcHSEqiUluNXhcUUvlMquSFVAbp9yo74Cw
plhxIXpvATuOtFUuryefKUlKG8ppcSgcjKlLjQetMshuu90iObt20Eo0t71T8Ozi
OOGNzgKCRirdvGAgBraMOZ0hlXJ+VVCKyTO2IdgVOK3sWOHwS+1XHIbUQ6rZ7hSB
pMJKXTJKGp3aAwadR7knFJ5ADv2D2UZaF2Uj0YEgSKNCJAzV8AIR7W0fAFs1UBpO
KIU1oviJLiVWRf14IicKHQfbU9rC/2C/5op5zn6xz0aQQnNsCvhgWZxZkxzwnV7h
swKJaiVNVjDISdwD/x9tiIMCEXKRIlugftziT23Z7LKxvCqyisoXFjVo0wQN7YYi
mcSjPexEV3atTelOADdCIqJC/PR4qeB37LnwS/4FiF4Ao38fRpXcCpb0Fl0wjRmj
wcJfBqGYuSwb4B8SIsUKDuUR0orTpbLUpLqQTsWBZ5nplIktunWmKqfER7dftp0k
9Lduck0qozVIbgpCQOg4rsIrjAG9zPHgAVB0klBidRNmBFj7/PeAiOpkDVFuzRY8
jNfw4g8uaS4/quHVfacyclcMD4F/vRCG6kK8AS/Fl8eFW/sSHDmZi4swTuGyr5/b
wKqE606cJA6Gyh+Lcn4BffN1rWwSu7iSwM95dByglSZgFwTmzv4TlN+ZjTJ7ieMY
gIq+NJBoZDSdFTMn1De5JJ925HW57xH3DZy5LXi+/htF1fxMKyL/RqiwuPQD85WO
tsH6HFNZrM9ThYFl35llgtpzLMJxnQ6Pr9kHevl2uarnutMzIKA0lc7YzcpXogFC
Lqwp8siyzMlqIcsVSzCtJMqWmCgsCZYD6FF0goUXh38h1vB5gkBknzC5jgwTjz5h
1Tj8klJqOMhqPKSe6wjmLqU2trccrIv7oUEfo7wat+BtnbKI/+SXqz6X71B3Rkvs
P1HdqEB4XGpLgy1/dNDVg0VVOXjcybUduP0iLREbq1wsKCJYDZSkI4+Zn/E9llJC
3GeYBvJ8/B/ciSvfLa94phE1pgd86McEgoC9pKw2aPXE9Mn3Sa/gsOsNBCThdVlN
bys7Eun/EFHqbeFAbVjmR1Z0w3Ar1NZT2EU8SC5pKc1NQFoRPoe8N1I42OZosh3/
+rq35WmfjIFkeCeTJnwZUZ/glsJPdZ/hF2XSGNpWCaire0+ozppRXbaqwZ0TiYSc
BbCnplfw6nx/n8ytUrhF32PL3povl3n4WtXi+F9MTsZ64FSDghbENvxm1AdW/pom
yNLjccJPvsoOdavqMS1WYfP5M95H/L6bhyNkh2wmL/w0P1jwxvtfnrcX/8JQCo+t
/wcTYMsukYAh2jg5fnA9wEfBKoiF2N7KytvujH8ZnBnLmbI0FobDb74RUGa1MNmA
zRERzt8d4fVhsQf8BOv41LbsXYQHIzgRuApLYMqx/jlP55R9f3rvYu5dpBFbpZ8b
3NWkXecKlx+iIkr2oCxwpqaekTjDMymnKa4VukynKies8wCC+sTkBjmqycQuX+it
vqb4+niYhfF30T1ra15o4RLnlOAPIOO1FTjO7ILBnxgEz6/6AK0h9OW+ybExIP2g
r9l4c61oOHYD0FtJy1aoB+yI0HrxW0bPjupH1HFogUXbE4LQCvYGdco/g37CHPBv
hlCM4ehnapLJvzEO7ardRMGAkJAw/1MRMPBbg7xW2HmCWeYw0XuH9AZ+EsQWty17
83XNB9XKL2BdV6ljqAMX8pUR5isXLjjZ30WQYHH6TZt4SW0iVtC5xc2GwCX+e0vV
hhwG76KUjTkSbjMWMnnKNjCa0fMdkDph8L9YhqHvzV+TCXCWS3zkNkErB9tlzP4L
GyVOV2tpVG3DxXLpFrfNGMJWnf0QZzd97StqRvHr2Vo7nmpyBWMj1CQTea7S9nX8
RyoM/hAWy8l4FmUSePl7Le/fQ2pxyOkpT8uc0OgFuznlPISTAHpXTVzZO+hn38a2
asVW87NIlxiepk1SNZja1g7ZUsXg6JjmZ127jV+iPwf7kKX7OAaWPRldwy4gvPz5
yWX27CAVkSt8GyYHEQmmYEjqtO5imT/avfcomoIUpRmOjkK4YAWYOL8pBr2ui0mR
Mw2AECIWLjzw6ZZ29GC25mra6n+gIivzYZ30UxShFOHXzefI2Qs3EYTrEQmUcw0a
WECGh7kaiF+dMbrjAbe0AE1KZxY1bthPYyLC/GMg0aG0E8IJ6WlDxYcbS+0c8Pqs
XksPY0HwofRTqzWfrO4N7Ys68+SQxSCvFjusgvvNbTf0bd3y95LRRaeH7mpaMXbf
igmxPXnCwgmK2u3V6zLClpJGiz8pb61OVv7mEiBgXmS8Wq6wUF2c9Sj9fIe8qfx2
iy7CFkIn4wiPuFicylHEBwGIeOStNLW8Tr+pcwBl4D7aXv264ItykGjGGq9lig39
sWEv7ZKpoLujiU7reRaTKn1ZlVEAXhfMy11bohlGim+kPpsjnSod4mdufK4Zxn0U
yHUv5yscYYHp6wK3Wyu+I5pEbkqn17P20rj/0Th7Oq4YLV/yvhL1ffAdWaWgZExD
+40xp6FvS0DdnEMme+oxNJycSR3WpA4wmMc+i5ITjwQHzUK0xgFyzAg7ZS4k1LVh
NMFzZSzEzKbOqX8lUx03is713TLcNPKMRh+snp2aBHtidmGgv3t2L/TQj16xVw1+
PsQtT5AFVpq0ld0sTnyPN4cjvNFTfsz5hlTHhOXAVnI6R0TYXXLNWhrT1WxglRFu
D9BxDpRrfQBbZbJiIcj7gTKBqIkVPyzlVbGOb0U2JrgDYeWbymhkNH4hM174ydpq
HZc4JH7oSFJcBHUIlIad/jj6qr+l4KHbujPlJgYwM7QempdFgCIXTnu5ELsmD+Xo
xo2c8OwFe3h6r2YShB4SyB1a/oE/8TjMo9gDmnIij/zOGfEpzQd3W3qKQb8pPcuZ
YlMkshpI58NeE9/1/YiJWG8mFSu8IeJrWfKf47JzhDYWYCz/hUKyFQU8Lz8kdiJJ
lNUKFDD7n86EjKAX/s++IiMGgsACw95rXpzbn3vaeVpY/UkyTcy8eneYVZWBaS1c
8oJLoLGxmU6oEENA2qFsD0M+ZblJfuFntkxVeunE20YizAeJaE+kUUaw7eFvn8a3
Esl8sJdr+TUQpJFIcsJcQXpzWxz4KfWptRt/lsWarTlVMPdkEkb9jvwhpreFF2lN
AimOBddgFSNFIynUZnthKArD3tBTz6DIwY8UKMYV24S9zWHkDTXtFhtNfzt94i1J
wZGu3gylJ327SFzesl/AYr7q3aACfwh8X59G0olryV4NI0261z2bHh3yJx/h/Maa
WGRBL+Q7TzaAqB6TW6CD3tm1+wOt/YcFra8U2VGJZrJH4qnJctr3VryWoZgiuxGa
BwUx6RHIxjLdvtLJTll8NuDte9GypFxM2AOraslDylzdaVknCFX8fYsnTk0+AlJU
72kpaO+6sNLkCh01d3Ze8CdUknQQxZ1hIViG6ne5mwEELiG781NshlWK8LAOZVAx
xrFYwoIaCVfOJDIAIOJ/9YBISPZ/JuLKESRfXJ0MKZFSUflGGcIngGUFQTM8anX+
pMLTDsaqkK0yTP39uon+OC4JmR8VBU83NdaF7CaXmBT/yDxuqRxXhC27rsxALlXl
/PVLQQOvErl2ta3t9flmWl4Y5m8hxI8r+oXHH8sd1k6Dw+qu0GyZ39VlEjgodbga
oS+EIPWQnGnWX0KCj3uWRryxl1ACG6vlmswlHcfrKjrqEskXwx6lXjxuqVke5J49
ihmDDjrx1V3+jMxyYiqbnHFzp6ymX8d3pzCGxXC/c92rQwfbvoEGFKJWLiwGzrUJ
Pn2wrJ5UM+mHPm5Rhtx215ZPXXkHsr8VrpCVzo7U6PZUKcCPRPsMGN1AnozFqK9w
TIm/Z9OB3zQ9SzpO9ChB/Rm4cHuzyNuq3f+uod47hD0AEguLx4m2iOOj8hmz0ueJ
NV/+1wHk99ugVqbdgyo1+ZVeYxy5cCDSWR+vNaiC5BDofREj6gwp8Vqb9g08kl1J
LaPkI4QpX45dMu7IsttoPP9FgUvVhHfM+kgc5Grc41cyYxc3qIfUjvJBPEF+CFH3
B4ZptCtDJOusQVYP12BVoOlFVrY6cpIb0Cw3vLlxOiMXoj6UDNa0c1xiHj0M/vIv
SVBASlWUH1vQ9WbFJmNyd+lMT5KrIpHqibZ6JM/77eP6C6DOvE11QeObwCwyCZyN
EctQ3CYKfvwo7wEYDKsGGahX2gqTK4sXR7Trxez4P7JaRqNBhXVvJfd6k21uYyM4
7LwZCgkpHMhaSMt57fbHLQ/uqKQuwijGOd2mKzxTJD5DL2xkUWkv0ybMX9Dr/6FO
VL+ImiwszfLpFJai3Fd4Wq+yW/uVeY+Yp840XSiuUaAeP4uOIGnqt3H1MDo9AG2w
EHbUrV8yMMtRFXQUkvQ6RlbYhipRSzu5HFxg9kKpXXZXDFPorAOmL56PSEtIKS7b
qU+zON1uXVfqIOMim9w2nIRZLcKuz3W+lMia86l9tMNSJp0KsmU6Dv2ZLl7pAeZC
OzBZmhEbIbVaZ3SrQapR9yHvCU/lkzpyOKBqlUyCV4MOuXm7Jz/Uq3mJbN+shBoB
ZqiJr/ASRspBWCBRdEuFm3JZmlxLFDqdvUn/oUOVZqUS1r5KqYmJNuvkMFju9Hc2
TlsMqWZPFrZaL1uOO9ixSkCBPsqrF2VuDQjDeiGkhK5DyVWhgtR364JDEqIaekb/
DmSORUJpMs+qT9tQtdkRbECijTk9KIbg3BgikSJjgP/5xahEF/h1ESIMnLAZEu5T
ImSJX/DzbcgWO/mbH8Mu3YxBR63jdJ8B/2dvh3xy85++d/1OXOGB4P5zjjGA+41D
DlC97wFEpxtz+3Yd72BsmvVDfQeEiqY+bi/MOrZjQK0ZlHIOzvyuWRmwh4lF2vDc
yvY+38FKzOxbtMoqjWx1KRsyMAfwXG+MTnqylaPvewDTCqTVBOkmjvPadXzoYKNO
AJTYoSLveSbRI2zOfDucJ5Mey0wAeEDbeQz2GOZk1FwRLPpMzt8XNewUecalR4jk
Yb0pGplozOS3z/egonzwSnRJndtrxDA6oFkDoOlcHosMoRbEpV02Aa0dXOwuBqXk
KGwT+VqX2HQS13lV0xntlHsfBJiJu9iywyyydCHATEspk2D1oG+TdsrQBLZwvZ3M
XyksSOAgv6yMZb5QlsOwpJjoxyPKY3mCiqg30aeA7bF0ISdwLjw5g1L2aZ7+u1ai
hSw9bsHYzJPXcshYw1nbpLBftwD7VEfvoyg/aCOzw4HJsKskU+rE7odacx5/UDA5
IZJ89B0MND7fRFlh7ygaJYEnUnJbGVF/gRiqH8dhQtf+DhGpy/NcJXtDnj60jS7Q
EYivHAKxKIdmoiEpOajUnfMzYxJieraOIoi4E4a0UyamPZkgkUigIrF7tVjTW8zS
mEmKnSEPws1T7RnKhror53jUvvP9s8m7icB8Y8e+QVQskJgWgseMI8KFN0CjpQyg
jM5EiJB8r64Oo6sssk+MwPgm516y4EldJjq3qpRdr9wSrsJg8iK2+z3FiOY+xSqd
Lnd20fS+AjLgJIJOmHGdN7hstqYfJsrUR/DcJ8y7LmxEpaHdk6i+1+PfpKmEFSs3
cWLDdO2afS6jW7WTy4ClxmqrCQeaI6LDD9B0ZyJg6gYFdGFaK70y0QF/+L3xyAhQ
R3YVxTldKPM2EUNTqRzY9Vg9EzGPNw2FKfcKzpC3E1ndA1Ub+YKQ+EL3gVQL6UBd
nzLHc1W+P6JnV7PehKOg/9waCwQfwIOTUnqqHxT//jtBOzRyGc/PPFasiDaH3Npe
Oii0voYQU4xvKVC3pXEl7h6tzchakGULWVfTsMxVMEDQpGgnAP3BnyJVXSrsP59Q
tBCXfMz/AUfUNdGrY/hxxEp2IftA/dMflpYZ8c0NA3P8QsF6v5FUMpRMAfZTggzx
q3LTsDkdnd8Vc0asQmRFt5+WSgVrRcXdkzZ+NpbOtD7+LBy/haRvI0VBuMCOUb5+
wgBQlMl5Rii7SuVlLRzp/ZDdqEYdnqMFrC4iHxhDLCrgHgoMk/bsdZJ9CCScwDfY
2/n2V73eVIAM5BFVavcbUcx7Jih6zH5KT8QeBY2QOw+9wBjl8J0DxaxIrUdFPo+T
jH6keU3cUSNtrY1U7mSj3QS3MQI/xreNcpG/D/Ktniz2/Shjg+cCjSxHJjVpeRFY
2yNPC+VTumif8KAdKzqkyNiZjrEFO3439eqcq+7eA03kw5+g+TJ/ryzphAn46DJZ
PatXytZwpSSE0Re1vmlRHyvghOss+q9u1tWNgS66CVfAzJzZfqx7DipwpPDpYFHw
lvytOSxO5/6MZZ7LAZ8zSN2YJO+IwteGVQgTY328xbgmxHirjQxJcuB6/tCUY9AK
Q9Qhw/e+9Wwk9B7tPwpueQlFlON710MtcBx3Xn2eM6Ft45b4XrQzfL7y3D7icSg+
iLF+DK9ZnBbJwXzO63klbY2U6nhl9hKYB00fuYZGUQwY/f9ybSoKggcHDwfzAYCS
syaX8EgufqxAqiWqTT74RQSbQkUIrahWCc0YfV8PZ4YyBqADIE+cM/5DwMH/gqJL
4I3G9L32+0K0ErKJ9lf5bPfnRJNymMW3SfsuzXjMcM5SC7lZpfcf+9dcf89ySvxa
Up01o1xpeUNd/ZGrRAiCfy7jz5C6z4AgTSY67PtCWPUHjJxsGxhpHNEefcH5gu7E
XpTYuZkp9RbXVvm08nnUG/Hu5oPMsxjLFOcq6hvkwuDl1BE6oUqVEzZmyouNlYfQ
nobCopMtKgUVJKhYU8CZc2iMzTsQFuH/Kc46O7kCevU1Kb9uqRwwLXel3sjevx4Z
K/tKIjmmzuuSBZRQ+A5TeVj8Yj4xq66kdzbfOqujtMXTGzxG1A0mb91/WoqBWjcl
xg5koltVEbfn8lGRd3YC3K79aqc6x1aFm5ZXjq+SFHpzqGpImcRC06g0zZ2q9Qnf
P2Ml3NF67yUNwimgLEjdDsEO+syaaRqI4LbPQ/eo4PQLqskzVhq6uyH9Heo063/E
L33zGVP3i7X45QHaYznQ1/Pd8vO6YRd/b4l0Uuwb9E389ESvgCY9Mr+N2ZkGykih
pQ8OTe0pFwDn06uqLK4RYfWDiNRQfGD9LtNJTsQbGc4u9Tog6BJ7nXi6lBIu1+pN
ON71fYWuGaKAOKBIAJrjDpI0VMMsaJuIdRMChHiC0QvLK9DlGUCVMBztHwb8y/Y1
LsoO+f6dxx5L/Iaskmut2gmBDn/b9ORPZp/RE0z7UD3XEQhv2Jw7ImeMTBfvVcfx
lhgoYBEt5B7RiexxNIBUh+XEguc0xroCMjZlbNUdfxK42O79Gx+rGcScgyE4Bz/P
F4xE65xJSe/IFYWfD7rUTBHcqc3vFN8PWG2UdltrKs3PnCjy8A7VStII3tWn/e5k
4J/D7ZMtDJPESVsQULquSGguTbMkbHYkluedkdwpZcbmDbi/cHPTEPzfz0ec1ulX
Qqv65E7ozgaObFRW5JF3j81JNjJrzmk9t1/BDIsshDkCJSqC5SLN0lxsbAjla4M9
+oJxwuR1i/L/r1+LvC+PkP3NMcP+KOeC/HpmJwV1XxC/Kn/ghACCrYvSXZQI62kj
g+TQfxWmIVC33ifFevhtfs/eYtFngtU7q4pBlmfnhk1DJPMruzK9njoFf3fGhM0l
Zg7E3oczSxJxyVn7DBU29Tkl37vy2rrCq/kZRrQHB3+rhAr8N/E3Ku0bze1I0fgA
KGLnczdLVH9X8YxTvZoY8rUhwdHUG9MWnZY2moTSzrj1G71KvI1T0aKhlrDuMCv0
g4ecdCuPA4u8zOTJKrnbBUltD3VG5zXp/Q2C4mSMov2DUtKa90GieW6CvG+C2E7I
fXTEalz031NH2de7BAeEApNmglIZqP3JPdccUOqDOrfOyoOBebn4GDhpIrIbdiyx
ZCnLJ+Y59cIKuhhIqJBuFOxfG7pUy0mYS9TeHxD4o/2h7PhgqOsWo6B8/zrKHoWS
tUcuyf/cjXKbYeqTuchxv9sGLBJc7WM1PW8MFaDOpIpVBC11RLkOkpRm9Yx4Pgl7
QO/KktlWEqzGmQD92q5FQtEGmH74e0BDdjRMnIqBfpsrFeJ0DXpzctyufbrYnIRu
aNt1nt28hipIc0ybiba8sERBSL5HckxwTMGZJPPFPgpJmvTjTeoJ9DyrvxVcA6RJ
+wZpCNvmtzrYPYsRjIULqNgqPQ9DC6Pnf5xnopk2IVlfk0d3WyKjOlUNx1DZ3CPA
LLbTeAc4N4rMBy0fDCtGS2wfqYknK8ejveO5b9Z1aNNFrQC+/xul9/E+poj9Shny
HNfwzCZUs1qu8ZAwAv3dSolB4GRNn9l+Qwfvjq3XCTb4dIEQRAvcGxYCH8kkpQFk
CUuc0rXx7fYmpBdzZmxtuscRvli10uKRnStm+9mgdP9uwdwodt2/TXaSxlKLRuF0
UQrGJa50SYN6kHPb9I4Xmect/NHlOgx2DlIHXQIdXv50+4L2gNpq/F2k35Kw5HB2
Vzl2BtqR5+dULQvTVPvyv7WngJMmxgbvNhovR6NH2dAGwKM73hiP3t7dLtAH5csx
JzOHW1OngmD2ShcSgJFZBFjv36TIxKbH6+T1xDkxiS9lkCT71kh9kYMjNiZmi9qd
B1ykprWtwaR4hg/Mzt7HdJ44WIRJMfCJbJ8LsYCY79WSWLu85ojhVSnD7T7fj0l5
RodxO0YEMbEKzAaHKQH/YZFuUOnZ+Yr8iC7EGfoixqojrIc3rdSE7VfyxUQWkmOb
DoJSm63KbHZ9Jgwphlu1K3NN5+iYJJmalwfElPAeEUp8OL/LjxYNKDbWfUG79Z4Z
1EDmghXgI0+2FUHOMpLfK2BM9o87hTjiWRsxjbrs/JNSuSkhWain4neiF4lgThWL
SyKTd3P/mvCbyRAlL3uDjGmPaVNANa62sGIc5mmEIyVMjIlmyASGI8MKiQraIB6k
Fgk3KUSwMJOofkgtJsjKlIMgpbR/yMrjY7NTAp0bAbIJZPO8YhRkP7TjTabMC8AT
/5ESmW3k8r0+qJsW4NbBR1Foe9xWvv7gsxSAuaIWTVVjcH67BvfqKUJH15jJjIXX
F8puaNCzfqZwsasbAPVd/B3Q5M68Yyuw2ZXXzm+LgEgZa6CmeHiGxVV+pkIXJHRO
NmZgIYy5CgjROMp8JECfvGj0V270g6ARF7vZmIslZC+D+tyEKlmZw4i1+ZYO1f/j
voTcsfD/kyzxrSV/bK4/eKVwdOaUXuFw6ekcj+9kHf2XTHarQ2TBX25VHKnDfXt0
jttVM1OojmnriXkO/ZJ6MoRLTqciTSlDnZX0YXVVr6qkWbBO5AsYVNbZj54AxvXX
ZIZ2W1039XyThjMEmJBne7Kq4CiGpgpk2P+MQsOuOnQjKSw6nnDimjWtld1yCRdo
nsgzySSi51KjrXnPo53mH1hBPm5NblAsMZz88VRTblhF9t5tk8dD91LY5+VIxwCV
N+lnmUcpEhKi6hEhJBhNyL4QbRJYxaflhX3Eln+Ks1FtSfPz208xfJBE6xbi859s
LoCD67284ulo/PT/IsGrqwvYGJyFNOhXQRv35jD5KP1P/mFh6LDicWIZSeM7Bs87
AO7LQpwx5X62s8UawjR7ZEmyihchZMPaOyGKVHWXrku4Ju5gA6SWJkOBzNGN9W0q
y86HM5zKvj8Oxe5WSeIpvqURzpVeo3BPBnTdAecm5UkSlAaOHw+JfZFcz4AqlEPy
RkkubqK4UdcAuU1O4J0JIYe/7dpynO5qoxctpDxDi0nn9wEMaOwfopSgAP1F+50v
GZiPBkOykqXEAnhOpQoeb/Hzp8GAWIIgimDTtXqhfFQMoCHqZgkpxYosAOrWIYgC
MwCAesFAkmpm7Y90XznrQQVGNWb3xat7TitWxY9D4pkiryR74C1lw8KqJE9x955E
jVlK1zFYyEZkImNi8gMyS9YL8PbLBQa627zpr+Ky6cDkfCSEViKEYHt7j9ABEWaz
qCSuKBoUxUe9pV4aGYfIRhYnrMxCvvaw7XVuZpRFDU6DQjqS0+lfEmIZLtvbT56n
wIGQsaaWv7dTcaCYlb90o5JJLq61oR6ZVwadS0u0XXiRluWs0ETCECrLGv8BUdwh
5m1LUFAphe4WEjr1JA7MJc3DNX+sZj6JhxhKel4LiokDRFaW3E7anFwYFH0lc73s
a04kv786DwZmCIs0Tr7axaf3F2guQWIWSJt2aYEPyv2OU6f2y7NAhla9K82xisTk
4B+mbnAsOGR6320L3T4mSw5xZj8P6aHVII3a1St1ZM9Cz+WqJZ0HstTtRQ9281Tt
r9LIzUdumhmszagORu6ZNkoKKL+zXNmCHgXzOwzdELFd8UzarH38VVTnQwC8UADd
mOUXsB1Ixs61kQvDtaXKTruCCl4XiuGPw5OnUVcLSiznsG3D26WMJhUJHS0tZFVy
xOn9hlMk8wAmSBDd2dDzDiMEXHU7K1o52X0W3KmVLWdsqKWQ2ZV/LdNs4cwo9oVa
tWKvOowV3PGaCsxd35lTnDCq8x4MmpUW1iRxMVH5k9Di9qJoLxI/2wZSaHzvy28Q
NCYhDWwegzWBUCRnb4RRKQ68NgUlRPbhtiLXMdtx/TYQq9CbHV/KQpZtoxj6QomQ
Z2nUViX9w59U2qyvbbz7ThV0KkdepWbWN9sQEterm37xRwgIIG5J4jW7bjDFhWcl
KEGyxjMCT6138m4Mgj/xnbn9aNOdXU97sJec5hnROrIscQZeFS2xFOsb4NLxqolK
9VITOa8eBYOPxCWm5/UzjcAgS2FdlXyyOM3ywEaXE2LKlLbTZCtH6PHtbjEpmerY
ydN72ab2X1JcmmF+2wIdJyXYucPPfjTmn7FtHFMnjqGrlhLTZSCpHMlG3v12Hgyt
22PeNkejw26geCdXG92gCXcVctTSIH5GYDM6IRzB+cIcrYYG9bclSuJHXSaaxr5I
PJSX3aznLI1G/9rahM6y8Vh/sT70OH6iqiBO08TIaJL+L8ojb9a3PUtA4w5bv5X5
XCVDDKoPp9RUP0YwkCaOEtBY4SwyPb0VePrY0QQJgYNWbsXnb6PvHieImRNIXy6f
uCtBB8hFiVapgqX/gjpR+AkRqUOb9HagOfuRuUVYK9oIfKs6aQipKEq/tSKiVfA3
nZm+rq/gNV8EsjqhksG7gG3st5Xyqzycr9mGefiLcv7HCszM1rJCgzREhyMGPJgj
5QdrLw0siupYeZMLIeb70DbAWWWwwRGpWeGpzp4MSu7XVjtlERSHdrmNcIGb1Qge
NShSeYcRCOMvDKMajB7Acefg1W9S040WPsSkR4fO4DKTMAxg0DJ3dYvrbkRIEOHY
4eUM/5tQFCYaChXpaIWdcu1R3ZGZxOqIkouGwqUh9u6zw41Uo827RdWYQXNLzSfN
g3vmdBRQIAEkT13m4E1IRwpj7A6iiVJ3Qit1UV7Cw3lQn4ITr5XMfQN7zQEc1ini
M22+FNA5/nr7LLZtU+fleazY14Zx2b2mGBpzLdUoNG+9eyOaNRUnDXBxbO/rqENW
Z90yzdEQRyHVEGHiEd55lUq0CS1tR/TM6GighcnaLAp5nvTs0F9McZq/VqxUI7uU
LM/erCAetomDVBueG9xvHYLc1au0BPTrfRyc9+0WF8E5ayKTt5FNyv+lEnhXgXFH
RX/+y8N7K9nKO9kWuKdVBs+WqYVH3yj9qAx/twBfXvgyOGn6IoQMa4eCpRJFSP1b
bzvk07p0SQCrvfuEt5KwXiAOuC+aSByRQ0lv5mStCFqVXmdmQ1VSBvUaipdJWiYu
jRrxYzUxADbv72/TxWX3RywUzkiUkxE5r4wC5ShJuw1WJJmbuKWH70ccnLBBb5R1
DtK+ZEhKwiSApFH/Bmo156VeW6dRnGSU4ya+VVQxzAFpZVXF+Zajhpmq3/UBMynW
ztKyoObkiHPvL4Xr0t4Eze+2R0yf6lDnrPFGwP4QPrM2QeJMVzQI7C5qx/Aw+rSf
s7jLYjE5Eo+g5N8IKZXQNi3l3cHMdkJH3UZyjkLnTQmU4DPLszsQGHHXX/LnYliu
cHX9ysahJzctPVDDslm6Mq1dPyhUtCnimQ7378dghZ2r3llhAKAqEgZvrehK3M2e
Ns4RPk7hdWmS+dEapXj/MnAxPIftJA7L0CqDm1+VDbCVffy3fK1OOmEJPwBQqHG4
sHs9Zvr5B/QLh+YpgD9lKGC7xaU4kISYCY+YCe+x4L8R1P5spP8gyxl5mmOaQ4/9
Ee3wl6o/hxVrnASNzu/mTuT2PsBbzBxV0BuQ1Mz39SpeF4HQpHhCxhyfbWjOvUD1
q9JtPNmqTxo4+y+Y01xzS2+fNRZ4Z1m4SyXkcGsrqO1JwHQkHV1hCYuUleoZtmbX
odgA47p6eqRahcffJn73K37aFOx/YmE3Zlrn17QQzrvEY5PgN0uC/+zACHvSNQHO
OXdsug+kIReTF3sUvkAYam/7rf0YXwj43JELChMWDhLFcEs9FESjDxeXBNPutBpV
1HGmxDa18UtWbgO2PORpBkVWqzS+lafyxNtkP98zkSJSbxFwZFz4XpNHfyI5MPPl
G6kxzj2DYf2UkIUcYWii/EgZbrA2OhzGfi4ADlMyEA2pueNqeZt1ESLtV15JYuyD
nplLx7RrY1bFGK8UKEAMb4YXPmwrZpGRxc/TNTwuGVL9HqXEmeyCwddn6RWhsflB
46frFtVe/LfQ7k79jIwxxxbh3rdCS6eXiqI4hL5xvF4cpepVkqtgKqxDArp84tpg
Udq+2Fv8UYSYsX1hrt96Bb4xSKQrCgDGTP2w6yS2k5Iuxl50i+Wz3vEDF8sPIt3V
AldFclmNShx7CFfPSa4jk0veNKafVYq8eBg4jjzbN/rijuO+GBEJ/1JYmtio6Emp
9qgl+3b1nWvQVOmmLy8cotSV1jKweyE06kH3ZMLQCvJWdltvVYDwYvzfvDMl0Fo8
n6aXVJt+4kz2n2w6t26k9aTkX0TZ5v/DdEzXRWvOyoG3a++4ywXSj1q2tbC6bkss
EfxmZzBddTGbabqoACQNSrdBNfmad4VoS/QgVUFz4rU9ZvJg+WTQyBs7huY4CZeH
xDam/pQ6b4ziL88mFx6R42iDibtpXUoaz/pbuWOdy4I25TBvjsnv/CiGJ/rKJf3B
gw2hohwQ3ugKWu9nPyXTDgLs+HDpuUzBZs79eogWXGFHQdipiE72RrKezrYsw9QV
D57EdmcFMeFpsawA+QUT5sKvn4deHkx35WRUMghoxZovPSCODNhyhcb79UqxR9OB
CrH4g9EsiXzcgjhZgxYxJ3oyeA2Lko5RlhslgILJnyOctG4Km20IsqlYqB0muRMi
SgM7MsQMWpjHrRsi7Ej9zgDPCTyyTkvAKXZ6IeoAMd3rsfDLCf/Fc0iOXeRQrnYH
pbjhyPu/7nj8aVZKfp+og09JJmrI/RAfPArME+4uXk5taL5qXl39t1tL2X4gaFQ6
qx7VthzhhVcBAxCWWYJCVPE2JzF80pG/31XCzDbF4atci9ejDk1Pu2be8MTshHpa
tNX/JDyOUY1CvLKubQX3kB1zII/9zcOqH3hXlFRa0JQ6ZW63CAy8UqarzwAqvpak
+dZH1NWbBfNAz5MpB6QWTenI5qpXuvnHMH3v5e9SUt9qbZqN9xS8+agYS6ud/72d
rXrKNq+D5+wUiRp9W0ns5ejxl3Vj2MGcG7Pl1s5OZ2sfd5vQCjCmnsTpWkTXaI93
lcziMDFyVYZ+/SQaYcreEPyXbIeY88bTlcMS+Fmahm4chhqrBrDLS808Gf2zRsvI
55cJLGbp5Y0BDPcSPauBCVJJ6pvh4OH90HjiFh1E07a/JayrnNHW2QdJFcsSVluQ
iKZyitMy2Ah4Dw5YXQZwoy+ap2vKi7fvntpSD768ihbIYi+5u/B61eALJC2P1FUq
koXnPpzjmBu2UnTcujpRtCfBwfZMOY63uf1gkAcbxVu2iWoEYxR/NP+LR7fk9LTv
gk5xWMA3GjnL4NbpTUlklEkQs485394tQP6TSjVnGaoG0SxNF9f6Z7DkTmOYXmw9
ygOr5vkT8wGeRWRC+lMOfnKlam3TbBCEIfwTc+l7MHiFXCRaEqLN1voXzTEHAbqk
FTQ7ukARfV9BuMugVnw1iwS0cVOvuOsUCyiavBs3dxoG5WeA6/5V/w8BNl1Cri6x
/KlznZo2r/pgRm+1ugisygSutDaOpHsfv9T2kwwuzlQop1RzNzEPytJLQXF+eprs
ciUnPkpcP7jZo+PRmSBz8FdfkhiT5kFE1G3Rzq7wwOguHYEcOtRM2nsDFklVooiH
JWbcPMvNm1bLcMCwhdhdUV8iMEzuZaRLoU9XAbcbqg3YF4MsfoOVuTQhiKHVvxeZ
TAJbmL35IVmEuaBVT3nhrk3Ly43d7KUiPvmJh79QfmOPT8lku9qUIvOebjeWrgvs
fNFqP4L7xwCeHgfMUKUQN08y71ww51qYutgweUgeQbrezp5WfLggTwsiAWNuY0lJ
eWe8Kuc1kwMobmd+h283HKNKJvnLknpg70WW4JENBUT+iie4jUmRm3Brt5FhNkr6
EFsf4Tb8wlS8bLCsOlMFe6AKCrtjj3a6EB3wUZs6gSa8zsQ7/c7PjsSMDcESGm72
StevstwuQe0WziZZM3XfplmDgs3AvsbSLYytnCmwQGD+tfPQUXmTCxJqD3dqLoUF
cUyrNxDg5avu/VBqbBcLOhqBUK35OLEB1PvgOwkMVx4Rnd2gCb9lTecPWEYB40Co
DxHsfnoAxyqPX4lA6Hwpgnqo4l4m9FC8OixjLl9oBAIkdCm+THiOkk2N7hssfeZj
WUfY+CQ9JiVS1GPInlHBqI3pgZSZGGhY9VO4AGS4X84d+y+viBq9LIdH4pN0PyH+
NBgzICAiIrh262SPYdypA8va4Tn7leL5iIlYbZLlTVAkqXSo2lfe8pSgdAhccvTQ
+uswW2hYoD9XpWsCOqe6c74IGsdaymoSbVu93Git5TMygjl0eT+/9WcJxApTf7LQ
MwFOIl5kNuw7tjPAHcsEcsPW8Q9egJDgdfvFJ2Gxo3liZwr5UEru3JcBHlf6cbL6
RZAhTDxxMIYkQI23ZZma13HGlQZ/2oyO+GjZ+xmw01mmCPnkqy/tLxA89W1QluiX
+OFpJEQp1ugoiDyYm99s/mqe+2sAkFrlvaN4cz90OwzrQ4HfBGyQyTcA0vItRy6o
px4J6mGtegAorLABJe/HoDC6WbhW7xd6iv4w1a8Jya/3HnVPOeCf4BXnFSbfXA1x
g9HVCuKMkFxVM4red3dOuvuwdCHtikmQqPNyd6vi50Lb4yPdH2wvXvb5DoaAeERB
jnY6FG/8UO5InCNy2IfvyJoORA01QzhSA6IfHGvRClfYFqibvRk0/U5QyoIfikbE
k1YYbZHi94qmppxe2kjUl3+JU+nbMnuKe565W1WX0q9LNIOWW9nDxoWuFvZUH7Jw
8PJ17s40/6myBRDhqf/0EAJSuFBPkmfilEX26j2zwrL5z9XmpQQIBW3fW8I9/qJd
SS07wLTmPulBm9YAOsyD4Lk1ccQwejj+IbsPkW2x/kNVIf8tCE5O5XBlWVbC+gsZ
g4Ea6bWVBDuiu3j7WMlkTI4WWfA4rswtBTY2VXxUzBpUBh7zUytRtS57w8mQcy5f
la3H8cIygB+eT0eiBe+tK2oBFqedMUhbhvNrbU81D6AmdMc1FzEmKI+Deq2wLj3S
FAnkvrpG62/bg/2rCbzkLI5j+Uj+8qoVrQ40ZT1nbmoggIfg1drye50HZyNfoyvH
wp9pPD5O9BP1AvZ8C6Zhzgy4gjUdICwDso/tQMeq2VYtjGmuLmjer+A4iSZ1BZ2+
HBL5fzyK1nlxkCynn/zFYXWujp8/pDNNm8s05vWve6gtWnGyqd0dEUc845MmJ/6V
QdMFDbEGd+E2kpyOYOCgTnM1zJ6K8JbgBC+Ty/IguVm4FMneomI/ySsAEU6s2OK2
PG8V/5ha9QF0mJqnwvsnVBVJwsB4hhWHipAuR8h0Qfh620E/PGtyQs2iF/JcDTck
zgbd5MFcuBbeP51wqW3xJggbuzOkt1WWOzTxQl+5e8W3ghehkuu6WbU6xqMiY8sx
7BmCyiWWQ0MtSJSg3vAUgiD/AWaS2q/3TLE1sn5MRDfL/Y32RyrGUOznobd1T3/e
UqW/dm9vBNbCr7PmQYtdKL7iCTLEhmEMLrzctQ8ifMPpf+T5iRtMZ7pcfgbj+YQt
3wpii8FRBLTN3zu2bfb/4vcDamE/bDyvl+YiL+EzxZjQZgu7dnyt9pgvejYDUbeS
ksFo4cO+ZNLFhrVPIXMNsuvGlvPu2jxYz5q2mrZlzUwDWRIm/5GUdrJB8b6SSs5F
LDIkaBANKiwxMdkR+f59mso2cN1/tcl6YOsNXUOkzZHs1EEjDbHrIXw0k6hp58cU
yQKwnGaJwFCAL4RpZ6f+wt6BdN1mFvg/Wtx0IsMXJhzH+ZL+7j2Rd4pESXVEB9Kn
Qre2NcHZZ1hoSBfT3xZmlqBcrpuGpykD1bvE+N1UFKk4qdinp2YX7xJdAnm5bJat
AEe80A4U79HFfqQi8ghhVWPKywjxOifYRMTjv30ko8OsR75DWfcfc5ONxK3ZQNI8
o9jHti0mTbeWuzKGBKzcihMlO1E8M+6e9ccoq6pZuaTBLXwim8wv3e3yYAJGEBeV
hBLazFoSR91fTKj1UaKKrtRQm7betMuwe7VfQyI7WDQVoGmPYDbMjz7H/vylBzL6
AfcWZe5/luyUKc9QIuSHT/ZUr5XMca/fE0eGiYvVqUGBKWaNACSkgRYZ9vVI/JpA
VVyEf/+B7vWsMLzUpPxTSe9bJ9itEGd+u5nAPKdpeqZVAqiT08T8RXharRGScDgP
X4igpqD49wLeO0nUImQ8BC8A1pE2n7+GnCsZSNO/y0+5/T182l3MwFwxOJPB5Qti
pnHN/KdfjhJ8PzkQdl/5XQteBwtUfFACLQtLdqWfnNfOoqltY8t3I8ZYW0DrMUAG
ZUdEbRczgmC0ZifXdPZcg6Qd7XhmYngsRXxCkg5HxahX3Cq6bLXYqoBswrun9i3J
1yl8UdRZPSDpkJy+sNLvpOZkxXUxO+Pd8vBRxasSH+ceFKkK1ytL79Uz0+O5oqvv
eCabesMr6CDyhfgZvk1dKi+RFPD7xlrVyNwhivYTLzuTuaXJ+v4027+LRJ7m3CHf
mbhAStZKdFEqurZltpHjfgOUO/T6bA4Ogf3kfG4biCEao17C3GSqu34m6+zO0i9I
W4W8om+2U09ZF9XXFcjzJJFr3xIpDHBHMfO4daOITjc0zRKm/fEbQdKi1NPaIn4P
mfbdVYVBn5M1NbrOhzKwpDuEa/W68PQXaf/IoAJ6Bsd2yGYqCKh8912eOdWkLEtV
PsbYO4rXB4WfHGmXoha7NAsWYIq1177XI/Dgzb/J3qx08mYLseFmRHELh4zNgj7H
sa6Es6ks3hbYmoyonGnLytx55l4krequZf8a08P+szhW5yUGSXGhVgP41twzC1Pe
9q984gLOVb6hVcoAr/ClXxC5G6GOk590SiljF+HFuObSFasnh4x0elqXgI/D6NNq
n+BYPL6blddiZ7wogv0RgiArwT1zZVtKqo7HcV8lQ61X4ezTCw7cVIURcT9xsXds
GjvfQx46bNrdYzV13/gaC6mp00C4ldCLIGg8cwKSj55vQMR6W/1iHFI1KcCaj7gY
nNkn5H/PrDZvnjOVKeh6QT+eTg3z583EsmP0PmP8Ajz3QiYNKMq542dsmlWSTKcW
z0/iZFUWcG1/RN7gwAiw7xbpG5nL3mdBny0T72+hjBn8LH+OOMYhkFM3TiS3590f
4czOW/u+x1soRxCFtxgUziMpPK9eKv62kM1XT4iKuPKHjb+uIeXdmyq9vGAvIkyL
D/zYFh50BK/C/1+I9vNN4coWG69JAkCkM4gQ5a8n9W3shN/028h2SVo8467rrzMs
SAoPOo7JHDLbUdp2KDjJYgVTuFD/IH2BMNSz5LI1n/r8nSveHqGHREfhHgEURWwV
veGmeF6VtAR9eaoXv/2U2L4WMDzLdzLqWym0P0LGCi4Lha8HZs9dLwrAXgfNV+DG
YxNuqjlrCQLGxNor1tqMdVDQTSXAe+pDBu3VXgKetJvHUgi5xXs5UN5kcsiLEeIn
nRBJGI94WkKGJr81LD10UOoiLQHDPIqmyjueGHdIPgvH2hUDpITZ7M5VQxSZTXo2
O/Tc5qh/6roFhsQkdyNaPqsdLtT6ABv+mgZp8Tvct9BNh5dsW+RspZOKB038JFBq
H+7C1dH6EvTYyhLx1NspxYQJNFU1xZXyq1nUXobMQqfy4hZOEzT7vz+nyhlYSPZE
mt5pnV0sm7uryCip2ogDROROHOkbLy9qh0NY8FKZH5I1SV6UM2hbsG+4yiBLPw70
12cQ+e1QzVZLyvBH6LU4dDmgHwAPbEsKlNNHVuD6xffLM/orKIKQoBCW6Wi0lLlj
jLcCr2KauHVhSGoexr9P6sHNDGQP+2koru+x3oTM7hCo1nYe+ltkKR6bHZNy3Uv5
vhV8rFhiLiqUZrXFV2HwnMm7cZaqoCUkr/wA7Zi/tGxV48dCG/FeD2G1I7wOV0J2
52d8TWhZe+ul+Vtfk3XSF/b5Ccssei8TzaNa+D+k7I9WwNxhlVmIeaw1WtciUmFF
axfpbI69v9rXEgPQ8YOSoKXo0/gImRluXxQegcmN+inGZqZpeyYWZqYtCggjcWyI
enj7ABNivvQ/ToSSOlXlMYu40qj4qMEhzv0IG8MMbGjpIQub0hs0h99Ghq1EGsFR
9uBOr6fXLoOALQGx7MJufNjowd5zbpYS1TOAD1nPE/SJHC8b5fJuH+hv1TPLL0Ui
/dX0eUF/ALVvuBUVCIuRc7+bKzQwjPq26G041hnhlgDKi5HW/Fbv4S/z6Kidwj8l
pvj436Dvkmr3ZP8IyM4rgxqMZE9bqyZMbWJskzaE4LoDUgQTR7+9K3lfDZroTrZ4
wtRv4aidZcPFuZjO3ZeExwWwoBNvT6hQArqJVr196Q84814EM2BcEW8elrsyJMoT
5hp5bj/mf0lxqnDeBYH0dtrjBoBqnsRR6Wf2jdTO768328lIVEKTRbd+zx6YBi+l
1+Mj/GdZPh+7Ik3InqNoyOnnKkwiRlV+agEmYoVjWnhECASu7HXgw7fhfVJqAhe1
baOhZDsm3K+47CE+B3VKXNmn6HZXUguDze/gIsU5H+Cx4T9/Dtsw+1v55Dihjedi
aP7H9boDTOSbu999ioeTB9ciLgo13cctbhxYGN7QFysu//ZeHEmGfjb0NcLXMF6Z
qt+qFvTX/vnre1RMn54+11lxIiVxJmbLx2zfOyckDvqUhhJLM6y8PSVWGWhD+u8D
VANT2KdQg6p1n9Y0smiNzPzWk6Bx22IPSToboVsE/GbA1B6ZYIz51ctS9UJy/2TA
3wcGZf+2xvR8GafX9FfqyXxa0mFsymizKdfAs9GE9JqIkOpUb+3XvDhhk/uNwWgd
v3ZbvJ9+PHOlDPUnVaWp81J37VjqPj7Gtm5Emj4p/HESW8aNdzaXfjLc6FNlMKGI
vOfPSilUMfejF5QMhnqYG/irtjJSJ69XE879CiYuOh5Gy1sbcrIjeS25UNwudIOI
k49pF5MclV/jvLFHTMDA6RKW45IjeGGAnFQgvZ0KS3fakMGZaYJSpmeAC0wV0Bku
rkZGl8ypB3PxcV0RgF7XPvY6Wj1/ey9QlmwEYeiesAf4Y6cxtR+82nonSqePJadi
3nHDlmw+ieKhq4iyV3rP4kBkxrdqIThRNWm8BXlk3PQxVkfnbe+6/Ovn5PLRXwiA
3Xm+XCYDtKwpvvFNSY+KfrW/8wOLpC8uQBe/P/LXUOpE2iBl7tfOk8L88acxp09w
CHz7Bv+btD/ALUYruvrjtDmyUcxjafF9udUaw0FZw5XOmxpG/PeZEu43TH8mOH4s
IW+S/Ti2LqbahOD7M12xEUxxEsKXZSuAqHorDTB6YdkKExPG9u7qDPG5UsFqU4tb
s7gWfzkZCvZGoB93ESmXa2+pFh1dCGOxeknPDB2Hus4AvaR/VZa5G/zT7U4GxXA+
g4EdxM7xPXrzR+DZHWXCaYLuuuNYp+N0z3JQQXfszgZwl87Tfjv/C76++jP0Cb/1
gPVo793tmlFwog2yt6jwLj/BoU/XaoFcBKziSZq1sb0d4PMvCoCOYodvyQSXdBma
C1Ha6O7Uvc50il95voEKUHuYBf1e0Q5x6X5jfyq8Cz05Uv74weBYyOKANRClbO2C
3kDaMubCdjNerTLghAEHjjq7VQqGejJru8uqkq9RtQQNTtfVUNHVuxZ+CT/i+SCy
XfTYRTQedn9b7uxyCfVS4/CeAWL+gBcLuscwOHi5M7FnYwGr34sHg+rHVvwyBg/3
1U5AIapuphT9NAfpo6PIHabgBj3FUIEaJYqrjXn9W3Sc3136ciVag6/26Q+FkG5A
zRJqFdgbY09zY7DBLBrwJDHVc2M7ATxukBhMwNB/lp6MjxH9cOF5fJZYjX1pTubC
V1ne1eRH5X8vj7bVFMQplYxA9uBIe7KuCLsbAxkZPtcM8NgvVGptYxGiXv2AIPWD
wl3F5RGmu8ywkUp5jFL9aHq/HFd7dHBSNYuci45K92cBC9iKeRXWlDGiGyhzNOYa
d71TBRoiCbAfUW1jsv0gXechQCYToytpRDPSSIshUJ6Vh7bUdCdNQMIM4NzQ7gKj
Rtw/S66ORs9w6o5zEVp2ZZmscZA6IHAgtWALrV/16Pe/TZtbAa61zeybYjvsUi7R
Pel7fNGaeqPX8c9hu1mQHeUEQPcj2MQfjKMPYFJ25r4GzsJYB6yeEeNTgoYBwyfU
PO8q66LdL+HuFJ0Brgu5W+K73yuCoSplV621HofI42bTgnVnNAYRB9eZWI2KhUPl
G8ogG3DdSUDl5JIrPsypiqeWyNsJlUUc5ITmjxJLhDd2FNKyMFTbG5i9vVK4mZRq
wn5cMeffZa8YxwBTM/ZkxZhvuC3wCrwsvubl5LoCxDCXxYTyymRCzi3e39gS3koz
YejGguV17zA1265QALafMTg1ZbK0okV4PCFzX8h+de4VVZA5tn4ok4DgnNpGpw36
eHaQ/R15G/fX4Xu6+nNy9GtGf6zW2xtv9jh2ewYlY4DTc6estoX4zDPlRYWUAlH+
/Zyyfw+1RZ6nxpUQ+pyxZY3jWJ23W+v2C9QVKJTS8BJI1QaXfOz4RdEDpqSe+7eg
0GMp54eapC1DreFGTKf3MtKgYexUN74znUzZFmOMvJ6OaEV34en1F8V6mZK5P8pd
BK/UBdNI+sis5AC2GN+XzVN3yAPRkNw2V2kOuw64KcA7YfNrfuUYGTt8KA6iVKPW
R/qJX0IWnfTQ/dBEQdqXivVQcom/PZnVNOKWq4l62r1alMQ3yMX0lXeFfCbogwoq
vJDxufHJFi7+mPyb2V0/oEIAcsboQPK4QjJbSSIC1t7ZxwYMC/No+lDS7IpyeFsP
fvToHF791molHpLlX6CL/VJw8sPPCLxbdYfS6CculHrWGhJ/6WTuSfo/KrRcIw+X
fFVbNBby8jOFoXX4h5fYYi0ckUV0Hr6cq/sW745gqDUDc4rjCaDwuDgsnpsg9Ucg
NZAQapsGAgHO2Q1FnfxNaH2QHrPLQs9CAyvXzddUIf3NUGRdRiQa375ZRgMMLFRN
rwLPLC+i/YWYFExuEq7gwEYyA9qf0BCVFWzOwGWVY4TxwSRWYbXpmgu+DNHNloYd
cZfAthynJF6OAv1e/Y0eIwp1VLyXaY/YYvFUjwN7595ZmULExi6NFeh8aGW98AnE
5JBNYNQt507cHlutpQRXjq/WrbOx216glfUYZXhbyxDiICeWW0WYo0jilS7EQbJf
jqZSBC5j90QbOErXuumuem0NXfvJKwnLfqmM3w3XuE5b/ucscaTa3bEGlgD1gZ77
Lsgrvimedi7XFLUuPf2hm6z4Kw4pJO9xL4D3vODkwUCpihsjTrCtnm7sc76prU9E
i9MNHlbs/93/y47jek40o9ThrOPgMGzbSAP9xg1i088mR5/Le1emrcdc0FvWCSww
TIjXDbsiiaF0/eSSEmlomphVG3eTxxLde3HVe8kEpfiCEEFJELsne2u7ZrbXs/6U
7kLyK+cof7Vsy3crMreMuCyjlun7jSyqX/1oiScYgiT0u4zkIz+6G23YrPRrvQMl
2/1seybYZQbDwVAt+lWuc0ivfYr30ijk0pb62GTd5cp1EDofeNIAdRJkNw11u6uv
bFtCijN45Wwg1yIGcY83G/33UiAiOm9Zbxw4YGr5/HH/TGUkDPMnfTt93FeNPgLy
j4Gk5sIyaUlwj2vpINQC6vIguyaTucSumibENCNFYmAr3y+em9Ar7ynmTX8GDk/w
3bChiu3oVygM0EN7PqfWK+gY+szewb6grY0W63fjs/NUojd8C4zg3oWYLl1455Tf
fuTv19oFkiILkraklqwAOeJU3wi2txiVSRRDv4KAk3gRVuftxQK410BL2cuZ+Lij
TMS4icd597jVuT54b+U9p52YSrdzs5LqSiy/t7QN8neT/fJfXC1yjqjO1F8MT8z0
qSULcL1os2IBd7zxSTBcSh1ougzwP2K7cEoC6eXL9maaLdfosQ/XaiUv/TFzurHI
g59V227q9ICD9VEcNoK6KivAF+T3epNzXsVeJIcbxUwrSMRoaudXDPqvuG7XPBYt
gEynstGaSMVR/eixTzh1G7C5j6it1gHpuZ0ppF1/KzowRGoRpZGX6yzWqA7c3JBJ
goV4Hwe1LmPE5k0X8VUxT5uLVr/e12Qmh5Ofqh9UbWr+0pkVOul85BRDBO434D/E
1JeRoapjlVWy/ts2V9eNYcIPGQQjph96ggWake/m+kAROaJYgemytxvPJvXA2QqA
MrXTPYTOAu4tfNKPD/likQ76xspsr+GzXzNLA/1J8+wbjeVABto1sU9t11nBMjb5
d05YfZwg4kB3ZZmw1OPaxOHZU1VLJCh6E6M7IquHe7kZAc76Enf32MBlE/O1DpUe
1xq9yGzbIDCep5RVv9pfSai8ySemgrb8TBT7bW0Hv1Wde7sItMaukmpy6bCAoVNZ
0+XYjbGSr+BnWp0/fUDqn+NkzF0A8uHaIHSaAjtTj9S0pQsraVGKt11rX0hH+3cl
w1KKr0JALPOb6gNEqicthvqzFqTfCYSnq09Ac1wYF0enQakhVWbmLnmFCedcADyT
bnyCipj5XXoy6t6Yt+MzNoM3YN6IeY1wvGKIL9qUmOfC2CrBV7imqGj8cIa797RF
BBqqRTJpSOfe38U1A/xSNnPAvhiCURbUZo3tma9HyeLKvRo7TBKGYy4E0eaHGil8
LkfDEPsVU9MsCT0eee/frUbeEL/XNzZir3w3LtS0Dfnx1nqyxSB/T/3va3Oi43i4
T6FRMwAZV41lQuRJlo3uQmaAK7k6kwsXXspWc0wcea4LY7Wa0GDnJW3E2vR37j7R
F991MTBqF6chacFVWFifFtcvhBUDI2b4419wFGPQhQlUMdbe7sEhhfU6dleE/SGz
nKjO9M7ws7nv4NN3BzFE9c+NVoblx0iNTCmvEtArtQgm4DdTbOx8+SyOtmIAIU2u
UP+JliYlMDkITmMpt9migI7sg/ZKAIPa59FBS+LuMI9e1ieFN5zrIW5YoaS0FyCD
igXGlf9RoGoM9tqFaLT5EvnFhdr/yYtOg6I18jqP0xxlN7TWuz72YFgk3TuhXaOR
YrRnVDZe1YCmg7EoLC+2rfRZEehxijEe62h5ks+kD4RgkogmNpW7DaVurKrsVANu
rQSKgrCLoqW7ufT7SxF8aJOgWLytOfTaAx1GJynV3COvbekZ8DDwE4ANymYS1tB3
vKKeOWaDv/av0n31YzqZJ9NYepIkYhzv9z295zRSZLYusfDAL2fQ8MutBPPl+lcn
Bgm7fFd2dKYhsy3Oaz6+XHhOVvO81bf+CygKNK9/DLYEFZI28Ta+WNr3XUNfWuJr
zFHy6PA+/wN3Yxv8ZOYCg09ZOxb0cY7B/Mkzp1fCu7CGxdf7ZMncFoPNfvL/iLM3
JUA6+scaY1hm5k26FjcfA+Zq3pcHFA3U5VO/92pQx/H/V7pq9U92i67mXMIO31+n
uK9I5lU7gsEYKsJ7pFxcGudveQtFznIfDsggS/K7kJnn4UeY3TOpNZp5ZiTBOaRs
rGGyFrRqTawcdLicfU/IkjI2Ws3KSrrLZfbss4168LvR0p3r9nWNN4vs776rfRY9
DreqZDgzYPawuf3C7fzrPRSO9KiRHIuElkpGepg80mifvsV1Uq9RJM33ypmqJ//m
ncxxwI8pdd3cQ9vYZApue0aULfZLRBWkEaqNlZpz9n+6bHz7Vc7qiDVBd8xatPQq
8foBWJn0rigdzbo1teE1QUds+UTdHhr1ON20nQ0OuHF4lqJUuaChmVkBB9ux7bRh
lXZOH1uMUXOqGJptcjdXcpbJzZUBre1IfpjZvaXNEANQ0lvmw46Sf8NWjs3Mjo2f
20RoN/p11V05Pz1oSPpcbdX4u9jYE9B2x0oegRHBmq2rwVtCrFgbC1s3/MF/qeeu
t/aLKCBr/sn4MtAknbDRh7NBAaViAtQZNLYS5fos8+pWotZXt5hiFglJH/vCKbhc
09SEH+gqQbDUDEXoRvxGQENXEl9yDGE8iU9F/o1GqBaQBj0nppqab3W7XKQeOjOl
QZ0fYwERl5faMwCwW22WqmNk5QktXhklZwPSMkjlAWS1KT6Vm1jvkdSFQZcnJ5PB
3NVm4+P/tFX/NK/z7NoqFn+DD2OIGSYCOcp9ID5/lY+pKxNnNEGf/+4cju8Px5we
kr+R/6OK0ZGOHR3rhuv2r5ppVLg2BFrfm038699g2UqNMDoPMae6thXIEUmx2PEK
m+q37uHluOYCFx7cveIP0kkszUmmMDUMAmcWQd2VJtmzzU4ciIZHt7Lj366h4bou
zDgRjpBLWa5IafQE8XFF+YeXFwFQ9PJo1gIAIvwH9lwFpPHR6P9lzfXILW9XIyyo
P6Z//xJmKQ04GTswq5IjMTuqW5kdtYquSXidsDKtSSc8We+fM7rHmrPcYaZj+7ce
9snMp7tcDqRgc9ofFRCbLlG3JA9JBbXVI97TMNaXY3oMtmINIbz3LfL/D+5+pJVq
AapasgkM8BrWe5FCOdGZ5nztv6mqwBgTgPG21WxeQDLj/OSQg0fcpfm89FeoC/hZ
aLBDA8i50GH2E/qg6zo6MIxPJMojSRk1wngUlfTWDaBQrPSyjMovgp2d5YipRMyQ
goYinorWTfqdNW/3Ox0oHVa7eujC8UQfRzwG5lFEw5TE5YhAUyUx8KvYzQbu5MaQ
MVY6klYuQTfo4AfIWiiNiMx6rE1PPHYuJFIm03Ud6AwOKPLRSpc5f+Lo3Fa5HsOh
BnnenvFisGaCpcmvftaWr/jhEZLSGd3beBKwYx+NEGHy3rzkVh3RNjADlku8UDIk
8bpWC+Xy3W8tyaEiMApDzT1A/TGK4sFx9Cgc3MsYIpWRYSDKmDEw/wXQoT8OKRnF
YAq5RQvtaxu24iN1SnVF8bmd3aIIfEgrpKmdTho6uD7KXyDa/10wJDk6AtJ4ktet
CE0VVhdNPbYRmx73loKh20xSBB8guOl2PnOjX7qZg/HTAaZakgGgAM3YYhVWPt9P
sUB8kfK1qEHnWekzGRbM1Gx73+H+g54VyE5D8I5NcLjB8HbSljQF/i1NRoj+4p96
GR+fCbNW+FmBSZF0ouZcauVY7Ecb0i4Lfm1qPu+btjRdZ54DgltPRQ9GxRpC8JyW
gpHuLtpK+Rz0NU9U8YjLS9DFprcp3rpmGfTVp8HLcU4BArxCQx7CEvIdwT5Ua8Ds
qfVLsCg1vwCLbAiC3I3fUPTP4ZbuAXJBUI4f8hZcYnk7MA6endPZQhzf4f/SiN1m
1ovCUZofKRrAeejGi+kGA+Co07mrfmJQu0dBtYbvPdxSOsWTRlgDIpOLn+qJtO6f
8ZURVpMkXNLTip1LX3uYOjUj/c580ZFEp4xDmra7MrYYI3EsjDaJNWcOYN5t/lmj
7qik33xTv16CKyWhGzJUsXaOONr2JtfJ9xbQ822q9eKD2U27b/6VBZySlDFjAas9
lS1d1ThBvtbbKNJWOv5Oet4z1HTuzSVSgTe4BJ+4av4nn+GgmqKJBx84wTbaOuM0
ymfoLf4lbJhY7fthx9EwMQ8m5zOXWZKndLLc8ybfWXE3LfVYAcr6tFzJ4P+8G7lZ
rOsZYMPOUpzjtG7ZSUMEbRZg3spzGTPfPH3hbiVZk8eOggwGctgBAPCf4u/3sRru
iteNdhwkoCS6CaGhEKi+jenAM5n2mv62QJEkIw16EOOPAeIGahWls5o5lTDvE2Xq
MZTZKPchBgkkzHkPp3bjYMr3A4qAC9Nfc990PJhKV1SpCqimJQvOtxsB3IS6x1Kh
QBniNxPSBqALKhr2hBhWiXxQGkhlHlFHd8DxA0kq4UTS7xuPW0Tqkdrv9/fJRepU
ohRWGx6Fe+5ASg7a7AhKViJvgbc/JbtYpYyrlDx1tJF+jmjFKhCaGl3E66265iWh
PndEwPaFcrt2tixUzFCgfY8N8r+iY1Luv1GnlQgRtPviPtcAZBfDMCu5GB7yd1Oo
PuTzY+66oBndssnOtJMKHYnZQHhWhNq0KhwqR5fOqp63vkAxVCapD4FsY7vA7qdP
vUlVxgTaP+eOLqgdsNh8hc737euLvmdaZsZQqLEUCHeCxM/uBjTPaSDHYsM3pYVG
E065VHbaKpQ+d1XAUaU8uCEAacZ+bflNgAo58Ztgbj51HS+YX3to11SsQZOj1IrE
cWRA05ZHhpFJvoSgmt4NuLvQot4wAtf/J5mqa5JLXv/YRHN4U4gcOjNtLPkfL3tW
r8rtAC9KJgIjYMilyMP3grOMXA7NkbtB0QUidCGmyhi2LFsp2jX8tZBNTb560WIp
gV9yuKXqIJhJm5iA9eoh0Vfg0np3z2zWvxacSmvhBOmCLIYCbmWrwRAVQLzzOGBh
J/VsTeAkr1ceGPAiXieyM/Q1qidcHekAwXfFQ6jWwgdjXNCGUxIWsSnJ8tiYds5z
BkpLPYQDKDTyveMds+kD84LUuawl3CRF53KZMLiI8eZQ1zaGlZu42w8YpKSyOlnQ
gX9MoxCdPNLXObZMdTq+0JZCj8KChabYsyP1frvDoIL2SRUHKN/k3zwOutUqb9/P
WT/Hos8fnsxJH4qGf9GsioeSm47OgN0avYDhN+nEhnzRL2RAQp93MLlAuT5n1wJC
SXjiYDejnfNeKqXCDyivyj3H37mUyxYLJ8tXGW9QUUDdrLpLVyO8xkW8SnhySRDP
T47DrBptK8jKarJ9jt4jqWB6q5pjMh5YMjNjcLPaO4W63gLgR4Y1F5p+Whzk9trI
XuYlskEyC14Z2DPjNOPQzm1++mJ5uMIMcJ2KdFfedxA2RbUleOFKOyOEsNBGpJi0
h+RsvNmOkDgQrnBNNUaSvh/2Uj9YmrLM6RdSg2+2hH97h6zIb+LzLipCrSo5R1Ll
wJzh2OKMMRlWwngN5c5fmHWRX32s33qor+BZ+RSiq+9zb2VzVWlXXbmzd5BSHhPs
Ecmhm4mVZP+tBUrpRQfyVku2TwAY90S72FMs4yfKIza+2JoubPbPIZwsU/p9YEuw
bq4ntRWNehRJVsfW82SS+JoOkVUmsA52YCgeitcxEwc5ilBtFv0DURIE3W/vVJkq
EYsGLGJRNBQC9hszllkTLAmtRJJhQQlwqmEdvPACz7dPAkresk/kaUCdsWahr7MJ
6cez+6x/TYfbTkK5AqEw80qxuOlgTIiWsAJwITe1Yf4CfrlOtpSWkCNOHfDDJaxY
XNNaPywVY6bRheZXnS4iRSLiI7DzX+uUDdRNp4W4aSIQ8IN4dJJj0VjPFQMBa2AO
HHHbXT6VjBJaFSiEzVn3LYC5fYQYioV7MRQzPJrV1UhCV4Zq4h7Ta6r16FrsEhx7
3qvesFXDT4nufxN4vuE3E2rh9SzGanGhcmuUKQYVTNnrYpSNJbotCE0cffCrAmmW
RMk9JZSSOMM74aUqZbLPZ4yx0LWwJox4VqFFQyh+leozldf16AOu9clmJCHa7uSW
bwKqLzaA80jk1CekaFY0OLZAH4wm6kFlKXB8lR9sp9RqTZhw2NXtgtlZUNIpF3l4
XKHkxRedJc96OCJoCNCwVdmMMJJICvTCjluHoGDqgqJh7JHRL5ZCNAtGOv4sYHLf
qSwTOTus9tWr40f8xiX98xjsOdxfyHSemcBLBuo9ayUuupqE395OiKeL4KPTh9Bc
1FRzqP59hiNBFBmVKICa6mzYCNaJpMHAvT9xpBjtfUm9u+Hv22WmUD+CWlbx82l8
ZoeJmJkhAnQLcp59wrWJt3sZEBY1/iR5/8aqQ/4b5/8s6FQ3yM3AjcP83VHIaglF
LeT4UwjTWgr2/nAA0rCLTQ8IE/X2atgB7BVvoA0sb9YQoW61aab39m6+Eqa+SVBQ
pBP/RFFnmdagi9IatAwrp0wbeYWPTexODdr6mpYq8kC1m/T6sMjfL6aDTvOJta/X
cG+0D1BEyQVdjfyVhFoS9IJoIc7DhMvTMLjVPCLXAJuqJis0p8rCTcVIb1pBwjRN
T37PDJ8CcIOGafMnmPCwnb5XENDry4WeLYtHrzHzbRgEUiZvv0ANE/nYPkheDSxH
ZETzPb0QJm8GrKgp16xbatbaQi7P3W9eqyRe1oBPsbZAzhMcdjpjpSGgpQpvMoDv
sNt4jHpMIuteiOr1EJXPgmY0LdrPKm7nk997TUHfrmzB3qlzV9hfqnIRFnb7odpn
/ONpUPNGLqRIVMAbfEYr/n4nstnw8cXKXvmk5whXiAbumc4gAiVL4IdLJuIZTNxc
qAKh0qBmmkE0nRL2aaRF9sqqqeZSg5d7cSlMMfiEjPpnqYyfcK/tWECYA1ylGjac
liP/rtIs/3r3BDwkiwNcA05avpftDQuadD2JBi7guQliatXPF8Jov3KWZleMXoAU
iXxO7k1JlBHlKvewfmeUvE2G+e9gSdaqrczIBiblDTCLQFzEDJWgaS7cvdLS7yzQ
kSuWBjFd7rZOY+8R8f3ZO2mtixCuCtNErKUNpTQ5mYo69Cyh2mibKkuyX/FmRdIU
ZDCWe2ndm3O96VqaUrvzT87WmM9Wk9q5QT8nHgtqzxDDXRGhVLqKRSuaUvW/vb1m
hrvf9pv/k1PNsZGQC3TWHEMeFe9F6gMWqO0u1fEVEscFZLANa6FmqpB3xHIr7qZk
RzdC2x/JgKrZOzHCYddU6QNuGY1Sg4SJcFJJDol+kC9okAF3IDdjBzM0IPg/dUgk
0XpBSEfvYsbHkTRsuMIrrUxVXHWwADfUDxUifVOXRD9w4TUe8lNPTER1aOzRmY6h
WYpVZQfnU0N6O3kr3GkfA7W7dP3rsHg3WbqDkKpucFi69TFA68pqKhV+E6m47zs7
iPIbmwU7yffXr3nWHEVyyvajCFJux7bAnI1DmbYt2ZigvcohH2RUY3KacLOIkR3O
XQ5to3wcAQEqfjDs2gZsXpEfxzJmaI1Y8nWdp+PUx9TuY2f7b4r6kRz1gOwALhKL
hol9UloPVxmnEZO7l9Nzpn0BdsjXoCNUouj1JjGu9OrBipI6WveHB7NPIw3FIrff
PyVlE/vdomy8r7ZHPspCAwUwXapOqgB8+iofDbnVuvquaKpVRxfPtaQD7ZQZb0hi
CIa0Q1lu+GCJZXTlkWj5tUK8kWRuT2mJt73qeUjuEEt9G9wX6ecXb40dt8Nhb9r5
/omvpQtmi+4xwgu4nuug+MNZwLYY/Ml/OeUWD6N0IhWxsmPih7j5s/AkTUcQfMYV
Qkd1kVcyAMuldEkr5Anc/5kX0dPXUR6LIKv2FsTj7Et+S9AFq0pyTSs10UrOcDLM
at/NwqCd5qL6XvDKTWYLbEW/k9xdGn7veM/8pt1YrpgT5AzsS5KPbCSTGp0SZcpk
pepezNn3A1DzBCJcMociF5AtOUhy/01XAvdC/zic5s4CuIZxZkC3DUIkP0hccjwX
Bnhb4Vp40uqqCjwxkp0TPstz/ZOjAJWJ6IrX6hvpN+2H0o1aU9aXpmBwT70NzcI7
s4MWEYHhOIPBi6Ve5tDvd0SgPzQ8VivcF7vBdbS8dmffRzrCWK2o8boLQbgP2+Uo
VBSQQHMl+s+9vHF6/8p+EryF5YeIvR0XytX1ORZg7O3gSOVnAT/4ppr7OKVmvRlW
N5xY+EpWGi9KSs1tlTsXsk4UuIZB5FrTNbuiC/8q6IuVGSZO+NFKozWGMQJ3h9AF
IPWSohx9nwziTu2ZamFZljKqkgSMC/wnORVYVUolqv5Xgy47Th3d7LqGNQmr/iK0
q0NL62w7cT/B/GRYqqkCPrO14RqTSw36SCOvdCnwnbES24HxpYJ9cTq2dq84Mw9b
zgcK7O73nOw87NeYyt3CbxB2048vesok8Mf1t99Zi601BARPqEBKaS+tQVDLiAXN
EvSKnC7pi6AuTGhT1jsdphMOkU2PctgI1Mn+D5sJ7P3Ec0FHKQdQO91UH9pf070D
sJSBP0wOO4dnMFIgWNaxJMJcE+v1ySB1EyAPnOPwShiRQOkF+rbVyKY3x2eZh28c
hrYIM/Twc5hCN+tdRfzBc9OQx2LzF6BLgTT5D9okeLRpJbgoZPUTpu7893F1pWSM
BAtQs1ZpJDGQfCCzub7CSsx2F+huSEXTwDFdM8RKbp90Y3atgoNWDtuJ5d1cWxsH
LmIWb4/tsCY5acIQtS8sPVA5yCFLjUBTkYxzM9a1z8BWLxnHMF0MRhUbrPIrZ8L1
1//npsh/RGt1rr/YNkzF7Wxb44xANz7j3EQ4hi37Tg6s5dV7+Jonxtkw59jxuTeT
oeCMt/GjkOdIGIOpmpleGspAFn83KhPIZyyBj6Y32JyxJtA7W31645y/XZp1uX3K
76ioB1wmn5JaDNbXlcCa8FuSXbQVNrZQDcgbCRNxMEXbbevIkd+1KG6cFscACC2W
lga/RDijWVwBWbMJUzdZ4ew0H4Je2PVgrVdUZyZ+cYVeAemsNdDhHtlMRjHhPJrH
6BTcY9+LMYwvc9gkJFikgoUvfC1IQg+CTCM0JvN+BY53TA4uSyWR1gu9s+PQYJvt
kLyeVF0/90TeaIZipjyz/z0FL+PNosA73wDS0aTiwjTr+iPlClLPtLVTsx+iu/no
WA70EHhqiSnwIIsI8dFg32A96pp+umj+O/nBouqCDtiBpeF5xRZhMwafBMiFFg/Q
qRn4fiYmQYBpvxlpSXJZbT/zaaHpPUyVTQ2XUtOUWmXjRMhI/q3OLDUzUieM9Avc
eSMvhgQxoHxn4tJRcsedyUyGMRtgGMvACWDJL3DuAJzY+eWnghkeK6r5Jq9odfUy
RZnhi2CSoMFKuelms028btvq2UZWQMGaASKMs/9coaEATO0+Z5WkSdANr5h35wim
4sUJTCQGG6T89DQ+vlRD/ZrK74eSqzxcNdJfdqpwMEhvUIhF/3qZCl9DEosl+99s
hyM9y5ZCkagFxOtH8L0Ojovg80B3ShPeSjPmrvLaS39Z9olmU/xgotj2ynLAKjCU
cEGaVO1QKiA1KFZGJBskNpR+4M7Ztj1GejUiu6S7Y++kafEZyjFJEy00f1440WLS
NWMzhpW+xUXnkfl8zI6Jxjh+VmPBDjLPqq7wKaucaV7yxrmFLEikET0/DipYWdZI
KYdo+tKGlV1UJpYa55JkLgbCf9Tv63K4d2RKwsilAS9/pxajuGrVOq2/RL2+Ka5a
desC5aa8JbB49fU9Qz1ydz0hI1eQcGcGg5K4UF/89sDgUcW1ZjOux6wnVoi5BUtg
BMBo7Q4aWCTRgBbJpxwssQIu6QaSgCwzJkGfZKjNRK8czi/d2rodUBmVO2AjkfuH
RVN4ztaxHiWJ340LT31hT/yicGezFCfDfnG0dmCMhC85UOcyhqdkQIHlJ0acgRHn
2R4YvhNEUj4W5kwVEDJArhCy4LNYHUmLIhVuaUM4x4TMv3a7ybee/ojnUx5Grm2U
KW1pFpTGI1T9JGQQu6c17CfG/lGHGtIF1dEdWLGd3LAUW/8bJORAe/J3VtNmy144
XcpvZ0032KbIDhFhWWPpyb4c/YP/cohgY40AAm4GwZuFsc2RUw2UMlWBq9UkAdlG
hmzFTr20HArVuQo4f3i+gGU9Kd3sC/INaMvGlr5mvqJl4lZR1EwX6/8IOk48lGck
ag0ZSEpGqMUx6sYA9MnWvb48sQ2X1trAxYpPBTkOXufmNF/BHEbSzXn0374EzPwL
s9L8B0yREvn/XbQTZIZRA0iIf2PggCawRJKcmMsaQ7i4UD8TzF3iBkxjlVIc3jrg
xruqpXjsr509lMTPDeAtZxlr7PClEesrj90pa1JelOY8WIgLj8twqOpjpfUQMwNv
1n/95eZPADcAMBUtYTGfeXP3dPHpajyLmIXNdNjHEQaMJUZXFvor9l6/05PqNRr9
k9FHrDMbMFaJOvKkZqSRoVIyhMgiehFgHSoQFNIxm4RqNBaIVUvy4rWlkz1B/dLp
vOeaMh5lUylZHaKCJZlY+wfsYAchG/53Aqn8MrwzDh2LKhuHGrZs3Ux3t52qhDgG
afH5OdHCjD84Ic31kmQeNxPcQf2141zKmFIL/SOxyc5qkl20E7bWP0Nd4tmkVLSs
uy0iaMFH+UiaGC5I8nWGsa7JvtW1MCMpFiP1WldvjZ9TBzJoiwR4lUMGlkkPpXXU
fH22rqzol/wS4OMfnlYAEp42EmeLJIvGELgkACBIPCzPTGj0ZTIZUZqgNd1X6j1R
q2TB+5UMQ7xRj8konep4JiVIPZpdhesl2lzSD0UbWGFcC9x5BLwsrLjR1kWB5fby
Q7PK3caPCTH3Grv5KiFkoMyFe6uxiHoU6TN4edOUg12K/36nwri3QodZTTIuta43
Nl9bwMqKlcUvyZqgcqUl6/LgXzTUi6seOdWXCei0JHNHMTdCwUS5Bv33kCidHq74
8fxDF84+Jah5137VZ4THdglhslZV4TbUGg6uVX5aYa2Y4Bm5XrJwrqtMqyqv+qWU
Dhmelfl7k/9ev7CmWnXck16Q98WlPCIu7TOWW+SPd28pIPnC5iJRQEepJNXN7Hqv
vpImg+LBeE8ASC5FwbHIp47lUhqBGecqmREyqSK74Dmbn9u66AopCOoeiuZBKoGM
hfxyXYxUaxk41uzXa5Y0mhGbpB8vuk5ico1o5wgpR31cyJ1lAYVkiM+W2cWIOMwY
RDAXQQQRT3nGVHLlwIn2hEBBRMQAaCOgYnkIQk44k4c1Jo8VnyAkwdY8OzuGQfHq
JXX0T49RyNw/vIUSnjclyWa1X+4rkpNEnlBPFSdJyhsJN533CC6zRDoIodtP6cSN
FBXhSrmvVJwnW2kM+tMcpWnIxtxtw/GS+zvN3Awxy2JoznFAdLkuq8uF5l1ogKk5
KUDgPBI3ihU70eidGq1fj5lLdpLv9yg2YykpKV4cToGNwyrdDnPkShc6QFBiwge9
LKDFjBCQixl+HWZrMu2QyC44XBFtpeIGestOGILxPjnUyRTd0VBc1m2swrBjWvBQ
+Zt+LyjrmAWnybTD0YA8MI2WCbk6/JOfN8g0CX4MGogMnrXHqvWadz/2MCUV5M3b
jYfLF3AGwu8SlLEN9jdFEJMim0P/BpkhyRp6tAuwxnQtsnQQ+KX8SPY5ZiY6lI8i
IYjQcQyMTY7kSQReFurZ30YpGVGpMpW1OnUlYoBuglVAhluUjTdSmrKWWMAiT0/O
kNBs5cznU5dbkO3xLGef0a24d+dGy+Yw2R9K5aMrdiTxFLMUyftM89n1OFspgN/U
KcQsWsJAYx3KQPpPERuZiukbckKPs6YNOCuHMezRx0RcTS7XhzKudle5NHts8gU7
YQT/QQqT7BtuKaeWSZM+JGm5YckQHVZFRDpuWErwdVPY2CCCQgXfcsKR7MChAm83
wAuRORqesFplP9Px8YF0php8VsPztGyIngVtD/FCagtHr7t245fWVfQV1ybrQ0Y7
nEr1k/Ku3stLUcUAPf9eEoCl06IbgBEsOWbhfVaYYACJgcG46sNjv3zfODemp+pU
c3Ukrsy872BCzV/54n6BAmGYYxYB10bNqnZQP1tWyeo9CQ2UBhwEzL+jgNf2LzEH
I2GDXD5U1Q/YPwT/raglpp7GY2SnNJ6qnFwMtw4SZjS8VyztCcE8czWaoAezqegu
ZErDdC8vHhyqOW9IDegCpLNLzWT4tarpFRou/sl/v8hf9yQ7ZrswzdV+6D2fTMWv
aM7IGdGAFBqLC4Os+fWDl89Rvv2PobgdVKxnaI8AB88xu4cZxAKSrpZKcZnltS6Q
wFTbJ/uVpLczC96k2osDYLPLXBgek4zF4O4YKOmnYXoDizU5M6el5Cg2OeFW2Rwb
/WpSJy9+cnA1fwGpcWYTC6K9+5GBAMbWjEb+Qg6C3b1ucW5TR3ZsrYxAveh+6TLT
LToxy5CtCfVRrV8OEAuunSHIl+ioZhLfJXzZZO0eKiqaKl3eFLFZZ5lWkmmsYkpe
PpW4J78yTYjczNpBHHHgjhzzosj8DIagT/ciuHa8IwAqpYOK5l/MuB8Uto3zgPSX
11N+fRwAIecu0wrSOzOqScQV7Ywg8P9f5y6J0p2tnSllSoZEb51g/+1rRREKQ+Im
iGGaRswOECdvT1YAwti9UQgPBuVkJ1Ie2iB1i/eXaAPwPu8y4aOm0UQDYt/EDS9C
PYHhrk3E1yvuELMPeOP4NUgbm9eiyV7Ir5eYyg6n2GyKV3Jq1TUgvYwqiX5+MccS
2IbsiRLw47Rpjz/uDRv1ls8u4uvSTRqw1RTDk691zm3QXkL1TE3SxAAmKbyqMQto
wqAcCqXJDOzLBhzCf6Db++fwXDKMS2fTDPLz+JI5PfIko3Fb690jTKoGXnDuvrmy
Ziv72mNLfJBzUULaTNZ3gE74+upvAe7ovo+prsCJIoBGgg0xWq7vakf9bm72BBho
RFwXusR58n9b0u8y8rZRQrGhXKnan7zZQ5m4n3A5vrZLFI8QTYi8iaFYP2HV9ozz
/vYp8alOoTQIf8F2DYWkpwg79IiCd4JXWIBqyKqs/T8R868n2IYPMtjaEA6LJ6Mx
tYs01auNGTdGyggQsXSYILuskSxDVkYLmz9yOZ64bdV066sVb/LM1lFdC95axVP5
6znF7csTyYNQ/p4Ek7+M7863PbR1htpDmZlXQIHXhM0WzP2eL8freRaJwHJPqwaf
kwDghAzJP5D75XsLjtrCJSwi7NriDvGlRFlgFD5N3vYyHt2VSbd0gi5ZtmDjANFw
6HKgXS/i65Pu+XsDtCUt6fyt4VLkM9KBdR1QN18AnDrGbg7zXSaX4xs1Bh9nQpCw
f8Xc+aQvvp6wa+ZQ++UT8YBRCYwHgYP5BYiZJN0pVjGIsilRIFRmfqL7KDYrLBd0
hBooQmmTj03X2N6CYP0w3QE+/yICfAXAt411P7fjyTfmu/6iCoG8GNxPyUUt8vGd
8hPkVkDa3vlPs9QCp8akTWz3XKLuDtTaJxJ1Fn/H6hHAcTsRRlYKpSi/oQCxjiyw
8QqftKG2nLdo9AeoxdYaEBGCev+mQ0qbusvWbrRCDG0Q5olWnny98+JSTt8Zumuk
g6LsVLmiRRc5u+uNcqxBg8vLwV3kdvo69NxjVDxBzsItfF89hE2o95MkFsa5zTpt
4xWnSQxBhVlTQS1kGf+ysZuKmYURTyhPbGT8Uf8mD5FJ0w3kL3qtx6qAzJZnupUk
JMrSVI9OP8FnOTEjkGfNzmZhBNUfFo8sEd9R6VQfsYd/5MQhcV+uGMYQUecaOQhf
ml2djOClHZvkT3ndG3poYMviMWcqrHNjuh9rioSYtydvZWm5d+4g5WQvJf9jf8K0
Pc4BgXNNP0y5N/0js0SFosJvIaPPZNZszelQ69q1guIG6qKT0mzIwWYY4k0eNdxu
0o6q1CDqWY7BBsVH27Ak/I/81PArj29lChaXucM6PR9dMCjIh+E0ShhM7JWLakuV
GF2lFGLF7An6LaHOqlu9QZd7Wtu0jgjjRYqzOsolzb9wvC1MpYk+kpJhkc9NHO49
073JDWMhLQydK4fp3gflbl4cveJ6cJvIenjamo7U3FAflCshno0x6KvD2xaeZi91
WUhB1VJKcdFKaPy+03PI1+jZ/cgJILxsE350QmqAkQ929z4CqpHGQE3Fy9b+Wwbk
JFPbCo5xAalut2JLnmamJpJiBD+LuJwo0BTa7EqN3StEUKzvoHAcluHiphuGHDRr
7wkX+aUXjy05sUvP//K9fXdObNMM9iNnVoXmxPlX5KuW+YfCUE+6h9RHR6/qseIR
nT8FQhCYOoKVzg98TlJM9BERZXBeE3rrX/UhipXxsGFRuMdb+RZMlTtMob4BMQnY
YmeT7C079Geg0Celv6bO+X887z94Z1P/0biOVYteiY6pcj7ciF0vr2BYIVO6Wr4T
NgK4R+xi1f2/GPKVpuwwgW6mj3dxm91SgBSRZxpeg8z8Znl5/0kGXX3PH0FhydFH
c4Vwv7svUOfHBmCSa11SKE/7SUg3wIgInY1WMQbl0PjFaltd33w9d7zxcBhmZuH4
+g6jKKuGeQrcY2lXnl5iPT63g2FqNj4mZ5c0zFwGxgB247uqP21MmFeOymUiQWtQ
9kI4aRQzgMIIXLN54JQoW36opSjftmQi+cqKQc9ZR8+8xqR3MUWcrlpFElEtaIdA
5H036NX+ZGWqUbCAoXuEGs9XQgGYGdDwM1nxc+wzBLXkkC3usxpnILiJ40moirN3
wGCegJV+DC/bimdMrObHbPZC+hYjk9qppbyLBXUi/3VtpQU2BywysG4IUollQXGo
9CUAynFHRQkWlhGKX//Pi5Vlz/gWHf0IG4gtiaaP/VlEVvHZhFCDmen3nfFO8AIx
YCE0bad8RZgj7RXUZaTiU/mpirG0xzCUrTNEiVr+mVj0URenpo67xmJIHhLHDGPj
X5jSOh4JOu/b6D2S9AH5OCOfrAoiyn9aTc/ELov0vWGdYcwpK297eqOyk/eQq8vR
v09w7ZvhYwjArT7j/SARbd9qISmfGchSewyVViovoEndgSa6o0cpjEh+XgysGzl6
XBQ6O7zMR35o9v5p96O+kvhPWsIokKqpVg/s1bn5KvazU3YBI8x1gOCIskOkJdZK
UoDCl8uO5qWzjJMUArXm5QT5qrMOZ109HjmG/zLDsZ0agIDDOJI8g5f9nohDaLEr
6GvWJ9ZLwdnabcCjwPQAbshgVidOXzV9diV4U7gqPrMOJQFoZPyte7nX3hqZhSsh
Ww/gNq/viZOBuCDGYE09rhRTy26dPOPZtAl755qfQbG3/GRNbE0HEl9GqFuPZM0b
XNGjCQ+oYi6c4A5XD/hQcH4gW8CoSKT64UnMa8gOwg05n+aHxPiLy4UcmK02yLLz
7Ulfw+PoKY7ZJ+MXC65TNMvbAHcUPW09Zje6DoOwl89dldCTodGK7N24F67Abm+f
OjkjZUn5o+JkuTfwko8dMwCBTwc8XviTx8PLn0R4de1rti0RgcHPblSnVzFGBGLu
LK4OdgRrJp9S3JpoBoChRgw5FhW/5CkWZj5nNiz8qG/bCVYGLpDpVKxSpKMf2Wwd
/9B4KCV+e330m55XL0X4gd9w0MSKDybYu/sd89PxgSDt3b17m9ngv3TFxurLnA3+
473OkaKN2jmI+Yc7hVs0JFzeH4PJe7vULaTMNGSC9l5QYQG8MvRiVUvvbdDFvDp9
ikoKnvo+3OY6Sh8Nw2wo00T76ZqUZMaYKofA6KJ7BMjgnSpNeyJq0U3PQFWZ1/Da
mwg0SrCxHTS5emVJTfjgsOC2XIVHaVQ8Q7Kzk3l90AvuhpJYZVvEoqUAH1xg9gWb
TRetkhqc13oM2fAOL2UIVMhfkMsWelqv6bYGRcuwFW1DPeyatynmrxMfco6S6bU2
SFL9MPwiLnwT0fu3DOI5Wr+PoB2ofvhyzHKYZr6+8VXuDQ8QRtsgj+Yvj3Ua5VEq
ubfUVULm83/1p/bBREr6Rzbn/fBkc9F8SMHq6PdGQxAWeJhYY0XeeRqCv61FtVZX
HewVKfQYLE1bHNjcTe0S8Ba5ZaQ7NcE0uzPJg42NGGlN8AwOx7+BrwEPFDm8dMeY
HsKa6bKBziShVRLwa4F+uj9kqDk/s+xtnL+HJmmFi64gEbTCKTHRoJxzzBzEpQpx
cM2szOwhOLwll1lcjBBjcakv6uQFHqBKyVdVZ8/xTOT4E3Wy96jLnqX4VMk0vHHF
GzsG9IrohnQSbkRST9YsLEFLcolDLgavNrV1qIKGARcWnEQWcFgyLjQz4UXunQPE
0sBMn1pIMSygoBPof3H2NVv+mbR/r5HmyWjWwWDjlaa44kX8tpOV1m2F1zmUFAhK
6QuknMCVsVN5HD9CLm6epY8zIiGep8vQgDbvCo7ZYxmQRGltun9bNTlDGG3MUafi
5cOAfZ7ahpDcidDTKPtBd/4v4ynsnQsAVBMMkqek1R4HvWnYS9i3aUJm0gW18rpl
D0OjPjgluavIsaHUYkvEDOOSwNCnrTk6M4ku9lOmdZ7Ir6a003hiMDroTahcBQlf
1gy5d7WpArrJ48ME0BCTCrtfU6u7cSlc+atcG6IB6/fyS59kYzbNjvZOUdJgHjC/
Pl3CoKsWJFp0Rmw+oMtRM0dBuW+UIiEjBs7RJ2FPAZGgnYLAxi7e6IRfuCTt0Msk
mB9DUlwPaZhBCsr0gSpDG/dUFoPSycv29sWMna/rsZYsnUWC5kMGdI4Ww/YCkVep
JzN0y+C7UmXBs9ijiq4j+tuqOoyzanoOOEVTGhmK7du7a+MSK5MM3PNME55/qBJg
sty538UGDz9gasKssqLPq0sVZtHXgZNSIMrYpZGovdvZWALq2chGzY+HJmAzlZID
8IfxtuLiieE6VwzgckL2Rou/3XWJrEsJD67Z68mtwlZTZFo6KV4dZKwqEcY+TzaL
++U/fUgFDVngBrXnJb4ojZvpHYn1KTdMNbK9xFTMFOvcD5ccEGFTxUUWFUJia0b3
jS4nIr+kZmCj57bqDnzoRBaKQzN0Q8sU6lCrr3A0dCi0jnFNEIUSdFB4ZTtnvV+G
nWjc9AHbXM1xO/bJRu1Eq5FNjglSdCJZM/ITrFWlHMX2WE/NVXZYv8X1LhP/1Ij8
ZnZQxOSquny3gTQwmuaYhCaR8yDnRq3M9tCTA9zU8Bsp6K6kDDits29+/87gr6XA
FxAylmy4PEW+OAkhu840YLuxg0ux086zM5EuCkibK7r0AuYzRoglkyjl1Fp1QKm0
hHY6ZuJ9vBeYZvlknkJCCB0onsvTNf2qZEIn+973pMlX/UNqty28hBoXae6REHey
3sa+oY5Csscj7SepGlM8A3oMeLVRSGnVHgZQOVzOKY3dELelqZwQCflQEC6nx2UJ
LskPOVOEFfpxHzU9n56mW/FDcEF2ZcZ/z1cgHjXp1icOnSRosxH1GMFDFFwD0mOB
aYyMoP5S6bGOseAvSwJ7ZslVtmsgpuFC6AKWZrxFMyeKeEOpY1VyinaBl9bcGr3l
+xSucruM8u0wQjSB5ne3pvj0IwoYbMvr34CunANVyE87WPulutyVk83ab/16MX4S
lxVVClbeyM4+az2Y3xE1eCLUbcELBu+mu5M2jH+PKANjR10RnaJAjpIoiTz/Yn7Y
2dTVRBgnypOTtkcZj2wV0GE01ZE0YuJlBo4s4wNd499oZPUdPwWhyme04TR83ZD0
XMkD2n7Sb4dEQHOkfB89Urg6s5c6HunCKbUcEChaW1sUMAprXPvW6p1E/iVNTLn2
bcSlYKBuUdH6x4BeBOah0STgNTtx1opWxz28/o6xnDyflhOXIpxS4xGU2xBEo+Ye
9Tw/My6M3fuGoQ/Acnjnk0jnebh6XN58K94F/ITYX028usek1oUWlyzI7SvFT4sc
Orx11VxoqkslEona05J6JB5HAN7HpDhUqXgqLfusOmTYPYxJRLqaaV4qppDht4FN
SgXJi8qzTE9hTQbgi2i9CF4HwGL8NH7HUExUIq4fnAOccwu7tNRkLHDNXfaaxb+J
0qRm/A0U8HtN3V6w1VYOixwS1VHZnt0I9FCXb9S/XsHbjrflTPH9NLLLyLnwuH/N
Rf81SQieYHQ0je/fip5fjYaR0Wj1khhLqXPOFEoHzo2R4SUffkJ8Hn2zG5OpHh8I
TsMYq3aQFdQjhwpE+hqEalSrgQZ/Nro6o6e3jkn9LgTAJOGCpLpwlQBVKbHEU9QF
CiKLok5can9HeR0HN0Jgi9N5w7oFkxTAUeSxdm6DtChTu9R+I+JB8wu+0lr3jpRj
8Okox2ombErThW7tmnp0Iw9n/1m5scWOmZ7FnExGXDEBPKChvriTZcv7v5bSmkb5
eN9kmAtq0a3TMG180c9/4Hv0bo0qZTDDudjE0hO+pBjPHFrgKdzk/DvV6B2HeNnQ
HlVkKNY+cumPJhzKpyaka4N0gb2d8K4+8SZfzqYzOfvj2lYGHpIsQLXv6kL63JYn
nKFW5sk07cpXI9yGNGJ4zT7xFic58pyetXP3GMe/BsgDtpnyS/yUJhLLQl+10n4W
NesbmSI16/w+fekhp1aG+czG2gaJnaP7+H32Arr98usyVq5qfIDo1ooo4YEVNoSM
Gj+GKlkSLtyd4aC38pQ+pTEVpx3qYKPVUJEar9wrc54lQxMNYmhys/Em9Nj/FD90
0waxMqdF1QSoF8tStCjveVHSXdMKT9ndWsouLrz6yjC+z7WnIOX+e9GyzhNd2BIq
sSjZ+kT5uxUSfg0Y2AGCkTr6uykBGyt8eIU/qFgnHP2lkKrU3ZF6KkoifHIlUAXu
PsLQgCeaxMauxOpGn1HffCdLSM/fSglvHX0Uy1yo4EK/AZFmzxITP33Q+mdddt/o
ziegLQXbHT77Z9fEa/Q10P94HRrzZDjH5t+O/nuS8+ZS37wAFJ7TJKDhGabVlHMe
SBazNiLZ/Z+EDlpgZ7ydFPTR6AmEDT0Zz5Vi0HWydr9NXwi2WWL6rfqhuWXNvinc
F00i7dJqrqnTGdisI7nkllb50ftS7zVKKpH6qaYWwIAP64hE2aRWntTRuxdt0Dn5
bi8HdJciHcJMCFI/NspExw41VLe/G5PdeH39hEx8PkV3U/zXyQfAv8oG56Z767/m
oUqjCSjuLsgsPwaghK4EjObRgqxaYX7GrfWnmQISQhdYTibRL5IUR+728UFVLSpy
VgJJDkyUDKcv11fQrDJcK/SutWfJSqL2xotML7rcGVfLS2vbktOwlmBxMccw4DFg
Jg/kHbsed8skK451KBgUdoHhOCu0XlSHOZKRyBhftgrkrS0VA6Dck9wOgZtDuMXO
ti9jCEic9q5NswvNedxlg0Vn/FkdKT16T1fom1d/gzSgz/O7eBfLgBrQ2UU5JTUd
pF7trscSk+3CGuBtKh67VEsc9CWQJ04FC51nCW2sTuZtmnJAhq3sJ+WmmrkH1nQM
+7Om1LMAXAcq2R1gmOrPpPbghfonPB1C8GZm8cTiIeeiKdJX1nDjMC2vqH9clAPa
lGIg5kElHufGKxPmtlp8uZdaWAv+ptTuMVsdiyLC7xnvSSMb7TwiSKRV3SJjEpsr
yPGaNToMWCUOXqCE3O8i4LtkYJaguBmHCdAatDY4fw89RjBRuGWDNGcsT//GVjt9
EWPcu3spz59c93DPnHt+rMtBAOf9kmLLC59hPDAB8TOhr91/00sV/6E8JAgUgOz7
hyhBWirL+xCSt7QcYwhW8UxgVNscIPSgnFb1rqAu+JawhDMQZFJ1HdbD/8aqIDsB
z08ZVdNTp+87nmE7X7pRLqgJauoC3v5sBcMwvMeTHfUWIM5yBwbtNTsvERk2tzBp
MEIMIbnbstiWA3I7K0kFVA70etKW56ZavwX6kjlSG7y277XffgDrYMUBUSmjB7ZN
5pN747Ooo4DUZsKVvCAbHKiX9PxQuwNqxux9ZXMh6GRGLf7zTbsx81KclmQG68rg
2Ayj/SezRm+o0oLKPhRSl256SuG8NxUDk38xG1tViwuX6Z+N86ayyg0sjXvsfEEd
xxzTjdrEs9s2MXCm4vh8TUpssLFxgWG3Rsnnp4jO44lMurMdy1fjzm5n1hBKrYEl
A2LzAUihit/QTLRFa/8e+HQOwzvH40DFMRHRZOHqE73/Ft1G9OdvFU56Il9Sh94A
PBK7wEe9skdWe32sIIt7Oq/n+fkjCFIgTr8jNHwrh12LtxOUtCsPBRXSNsx7fgU7
1PqeS8cH64ZUUG6+vkjU8A5HBBLVUE1/LjEhv0UftQ8h0QkVt+zSTycUm5I7jvf0
Lz5CCqDVW2HKaVXeiyFEjl3lJgsqyowFrgHRA/vfIdEphAjuUqsHISi82fCBI2gk
gfhvreETkzd89ZAFZT38hwPrJzZzKo1Q19TWRYne43Qhakw0U/b87Hf9WbMnZnOb
/33XFwVj92wS3IF9iOHuQQiT4ZKzU0Ke6NKkjAXE5TNfXkVXbA82NFiQJPAHp4LT
1ZnSn8HSn85p67OGYe63Yg5i/Kj6dB31Q7x6uRAd9w3WTr0bGdInT5GAttlOqxUj
RJsdET26LR1hQWCb6rwDCvZe4HrX18TTCDmUQR59RY2pzLK2i05Op1NB1phENnn/
Vg+WLiI47/GSY2EN7QfeQWxFc2DSeZ8rnnDuwxfVkSferTvYVGnVcPHfX5TH3gwi
MatP0r6GKB1Cwg+OZg1FPrUYXLkD4PUt3QUUNTyOXDPgmez3ZeL1z4Ry5p7ATUtD
nUSWXr7DKzogbc5fAI7QZGIiERcs7Jb7wucQ4E0I/XKapQKfdY8Flo2GtZDi+PVa
CwAwd8fDT09e0xZMTYabHoaZaxYWmxBUZCpARl7zmI5e2fG0a4gGXmH9UpFXYtEd
4s7Gr1pnQ39O0+k4+rXdPj6s9YFmSikIlq0pRVebGEj1wFMDCSzOkeQSaVDCI8UC
U7PHrAsFLPW93PoEvxeg+QWhRaEAUqPWUkhYBGA6SJE/t0Ng/JNMO90CXGeMUtXw
hrvlagdy0PPBC+9vnGQGqziP9USUMgLu+wXK6vyfdVeenNCQF7/mS8Z9hu3gQbY0
BVG0o9d4QvpIco9vqzGH4Ju3t8F1Xpb5YT4wivKz4G4xboT5p0XfX1dzRVFnsFBn
R2z611FWz/cpHpXNXPk7A9+bLwYBhZ7fRTu97k/E22AkhKOVkuTS1tH2icB8dGBY
Qpe21YBwq4jRTtHjj/mYIiwPG4LqRdfOwUC7YE3rfxb4KFhX9TcuX/54y9WL0dM5
A4bzOR7WeZi9hnL/zg3jIRvi8684dNFqfdk/yzQ0WyavO0/I7epleD+Uul5Jx7BA
2IaSCr0Pim5sbnC+t2isQ4BVJLJgE5aKtZpCrgUxpaTnK5qYv4zZTaio906Hoeaz
Z95yiRbIY6m8bj/WWWGjx6PYc0hahXTRdhcVs1iFslJHovpF0eev3HOTuhe42EgP
ihwwO/5EtlIiB/5oQYpbrBkGugfwzWHxcOLl82NDCuVUx22e9OS8cnXM+LLjK9xK
OWwcxqUD8oO7MDd3hUwM79xz1/vZ2OJUdFwI7qeNwmo1qQFpiyf70M6IOW4dTSkZ
kk+1e8SGa8W6Ek05tjK+qIHiK14NNZ/4sebgS7W2APxmVBPLAqI42HXq89OXrxU/
/WSMCvvqrBWXU4MRBhqRNE3vFPXNXn7j3WhDgxVuOWSeY30F5cspEECopvvQCul1
wqiBjdD2qmH7NYLC7SxTio0Y2xOdzWWAO0+afEdlPm+m72PkGp9Wt9FZJ4RPiG0d
s6gcVN5WldYTFAOnrDtk9nbYqMYqNFLVQztfJ60la6sVf16g8+OYzkZRu0siSKpo
h1vUsvuQOHgay8RRjywqDWK5jHXKKhlyhw3kOUN8VPNi2IYeuFn2UzTw+1KrpOxF
M9dNEDwNZuap13kcPXMex8E32zcFs8HpJgULyhdEthzeP9jXrEYjIi06h8aRG5M6
KIIfxGMJlg6CCSIRyQnPmhaRlnMC805HBS3jZJZEXy7YOH+vwtkpE9J9nH2MmRBM
cQKX7DKpzIEs8ThZ7LAId8/G9uEjR6+P/xhsKlKFUYIhKGG7TH1ykT65nn0zTuoJ
fG89etdtK0q0oye2kdddwhvl01ETfmuZ+trY3hRfgkENwCCm8Trv3TvcDAuJFwRY
CkdVRfwejZkf848GzX8yNGkHhRGUNTM17xW6NyKjajcowSy8vEblM9iCg1FFTocB
96/Hsmdhy6i5PqpFpqv9XCY5Km4xKgThnTkPqJGi+qEbsTWUnT8kJzH8+G61K9XV
Jgwitgwib0z3bRZAU8ogvvwPZIZViDQOoozb1sDVAlNxpHu2uPQw2u3MD9WvX4ot
8hZMRO4EE8VYe2+qS3tSwgyS47IWCbdNGHU/Z8cuM3VRLrqLeU20qsC87COLVLws
KXoOUSaug0pMfj4BGWE/YCoRryZsMcSsyGhs7Rl2LKJXOblxxcGJPDLoSK8tkHmW
77j/vMNZ+V2MQbifmO0YacMbFIooUDS2uk0y37D/3sIaTNboOR6ZBtibkFIUEjg2
wC0O7xTVTkjKTap5mgZjGqTITu0b+cODBZkDcPSNszfoEGq7yoTlvz/uq4yOJGug
vm68CIymUHvn7vI0U5Qf7Xg71TSNtTOU8BjURzL7gGedcCOWBJpXn3Wq7OWN+K/i
TT/CQgVOA4gbj9HH/VxlgggnKk56EbuxvwR+dW2bzAUg2SvjH+wfDyYy4Ddvh41Q
PjzEJBHH1YciiwsCXCchH78xhAF6St+QFkDd2hSvLWi/xdwd5Gfspg8hd2EtrG6q
ZK9u0dV1Lk2LrYJI3QaCNsH/cmLuoowVi5U1s/mp6744YdTn7piZ/z1Ue6C7yQNP
uWVIz6BB96MZ4rU87eZ3dlGfrhT1skiWJ5hsjZT393caWlDtx4Xj1qmiybiH5O2o
GhN9zgM/lBKlpA1BMPsKXL1guc5mpWyQCA+soGFDDDaLSCvvYvlYU/Dvuy5lgN8s
AvfyPUKWB/bHOEka6qe1D5hX4LU1M3uIHrqlSotYqNiCmmj1/KktczD/YWnm3xxt
FG7vz2vcYp4C6aLegaQCpi/LsQhN6wznVsgLLib8ZusKfU/wA1+Fvt7JcYdxuqSf
MMN9nLmARSv7F8TWfThOq6Rql6uxhq8A6E69DxBj+KKSLTFM8xk+JwMDHZmSCfyc
jJ9MmKI4Io++INqwISSOpdzDDEfQwDCtimU7drRgqN6g5nTHRENYEzl5kjsHRFSe
67CTKGA3NCQorwjbJq7ZqELawsM4WQXq+JgwNuekz4jiNTc9WodbILKwAeOGR6yn
9a8jlbUKYLJBfpFDIkSl9uj6Zp1hzDWyDRjE0vI+bvok8VeQaWa+cJgeBcANXM8r
zGAmNmxwbp0eL23PhN8peRvgkbTWIUz2RymwMzoph5rtKns0zp+dUWw70NFesTUj
vi2WeqX0PEjdHgl06aR3ezL8cJK1CWMjLj4Rdo8AdsHCYchIAYZrCgvsFJ6moW/A
/MQhTcJCWBmjhQzpHsl7MBy4rNgtidhAsTFmEWLkp4WA8z8WSldi6e+/JFW8B/80
UxSGSPdMFryneWSYwUIhSbU7XyUKIyFWY7OmlLIEXY4NPrlq3V1oxEDm/K/gBD/v
k3PV7cqa+Bpi1w+x8ytBbZrX1xMdeE1d1XgVRQgVed5e/Y8Ed0T4UAhADoAJp2fe
ZkD+Jc/IuD6UZ7z7KPqYCnb1+Ihtu/dfOFEfWK0yGASKEN7XoM19edmkxZaZO0kt
blHLna4qAq3GYfW623Vd+t+vBqHd+nUhsorlcGUiPVy4CO4Z8Y4sIH2IdsEUfx3U
eONkARrPNn2Q6vDk6pTC0elLLTP2FyNxJiqD+DnWhH/TQyW5TZp+sORjrPQ0NaQz
Lv/6Y5zP3T3qSphafPRTqjudM9/+7XcvGv+vWHmBoaLDwfWKkxq5AbjIuuAQnDWs
EoXJgU/zQ5en/MIVyS2bUEPERLbN2O8UN/WcmhpPtbI5FBRl6AYqr1PVjOXgySAS
/ssEralnCao8zIBiVQftjpD98yytvsH3B5/e0ijg+7Hlb0Klfuh1GjdgrIX7Y76G
kDzSKsHa7McdqHd6S45XwH3PPDepft8e9U/uIFALGE7g59fEwmqyP4pYyOrL87UG
uFBfH1gXNd9qKp7fbbDkJAdQMOn6mzUFPQHpPc02XNhVQO6Ix7ow6XXX1zlVnvL1
/hYLbZeKANvlW6Ry6VGZ8D7N6Xe73+keE6bCiyEXRRrahnM1wMs+GJBczAsaxyBx
la+zNE63wuGYdlXuZnlGMFVbVnuOkaNJXE325auzXbyPD+nSyLhl8Si/bbhRylo/
75Hgp6TtAoN69b+foq9ZuaRjC3ikRDJHAxuqHmPyHijjPkBi1e1ct4FL8ru+LN4B
Jh2SkElYBSZYiNPRu+nxk+Ht6+5LQ33Es+b99kyg8RXZBVGC2ApxfYxkYSUuQrGO
3yR0rIlmnFLtOmmgFGYzARyT6MlUqWToZQxDCy8nNoea4jDRjr4yCZ+0GyF9E08n
ai9WRTFxfLNVKAJB0mPwLwM5UyUhU5d+N2KlzuAr0MVTrQ1twChkhzbQTSY2vmsj
/b5BH6FUWX/3ipHh/P5ZG4Ry0PY2EA7gKB0WHIapLHRplArUy/7OQHsBPVo4Rsf/
R75zeS1HoKuffBYpbjj5mJFOg6p3v+fj6Lm6tLweRh8/7pp/CxbujjCP8ukeyWox
k9Bw+jGXq8w0gyvDb+ee8QjYDKXKwz+J4WCbvhRH2W9oJySmfysAcqvt9tL95txh
spEbjv0jZEDvZIEPXd0VozjHetsCs3flfM8nGjaEeVH9iErqz4BrjTpna6+RSSjx
IuWIGTSI4iHCDFMojybFxWOkCPyPCXA8MQQQZmL+wV1WsVV/Vj6mCRATFFoacdHA
Vb8t0VzGjCCsihTjwweaxvM5f61C9dRfIwL1LyrpfF6YTuDuATAu04gRZZT9qHY+
qeeEYKdlFP2jN6OtSdGDmSUMyzMCexeHOyW6bRATH/pLXct2ZVbKur0NcGe5pIkb
vAcIjbSTGjR9n7Ki6ql4EE4O/D6iG4+RvUkCTBZDD8JLBxfM9oohjgMT2ZP1tuuF
6rLxTL/qRfOirRCxYIM28QeAPdnCDDz+UR9N86PyJb8nuFiIL0y97TQl2fN73zhr
T/PmWGoMX2Bpaugl6AHADdqG672uYJBw2jKqRuCWeiyhOMSSEF+/rl2fYPKv/lqi
oIzl15hELevt5NkdRbUPDPv8DVp1SCwn57c+GUmP0jLIM6rdFQZ3G2EjtjIz1myI
BtJySHLojoroRPv2UamW4RCeqqOue4wNPpGmT4QfMR6vvOgZJgHUUtnSi5EuHXHx
vvwWxbi0IUcT9aBpZiIf72+180z/KAfOg7B67bHSDKIDKg7Tl90CHIEsfYcmL0lr
HVbP/9YCygfUEiuiFx4h1DzJYanPtejnPxcKygzdn3uBZVWJa52rSnUzXp5I6CEn
H1UD9EFtsdl4AF14u8AgxxrQWgLHYQlUn52qyh9Ql5AZx8MgPkMEeNLQQ5RUWXV/
f3z1cDcFFQbVplYmtu5xL9oTzJtSCdoe8SsCsevx28iTd9pcn0mYuxKiC8Fcf3l/
D8t1hAQYVxGhit89glLxf6Ia2GyVy3Oq6ozV16SV7ofmvjjWquvvqpjUkKcuFFe2
1vkAul3BexgK8UgULhm1yqBZLzD/htCwu/od8mn7tQzCXbf/wSj/byORrIWZ3wjs
gYzcw8EXdojlpDQv2GnBQPLEuR/04bgrdswl8j3tJP6trB/LtxvV+vBIEw5wqi9p
1DnN9XizrbRDSQe2VTfoKzd0Va+vBW3tVBc/ia4aK8GZK8VSQuJOaIyiuM+wemR3
xBWmNu51TmzFQ9HwZkzF5fj/IT0laDstzbsfAf5dVIxCdOvQv1KtZ1zESv6/y1S/
K8faCS2Slo3ibuZ9ZXMcEajYKQ15ppHlPSlKwFhSNVf8iqhnC+Vvx89Zkt4xSnGc
q+KtUB+eKeUwV2yoMAtFNJK1wX18e7ffIZ3ydhr2sqU+cNHtl9Ro4ieFC38iEU/D
2VHIkOIKWTPpkdjkFNOeN6iMd7SIhnqzfxMN5dt/ldYSGh09tod2AcDwWRl82JmH
Dr5IzYVLi6uGEXuEV5r46+SsLdd7CqoBaXPu28KNe1iJl2Ywfohb11DVj5aN2nff
Hh19DOs18sih74KxTWRvDesNAjVi5ZBXiqDx4TZaA8GcQvlIhHau9MufOCERoDkU
WTVRzA1YFO+JwSwjUXuG1orBSXdiCeG56E3rtF0pwverRtsXCBQeWVolsa6gkPAj
vsRxbauWZO20/ivkAaihpDh7AGAzTOJ3hmM82Vfo1hiNSw3Lc8XPx6kht1j0FvPV
k4b3udK63d+TkYunkk92u0RraDbwt3S5RhmFcczc5dM6ConXfqRZIlES/zH5byfd
BqGhvEhzgPo4Sn7bgQIPQDsXfY7F3VzcuOazsOoGjyP+o8ntot6FXZoMgl8q1sMK
0ycah2A2xxHKLO0BLosE6MQjCh95P+UOjvSxpE6MwjmdNXti369HkNXcFeuCa07t
EUoHOz10GBC6GDMrjTkqYiwzXVO0jqHJk0tktKDjdyVb7QUlsExxVVlFj51Xlluu
wOBZa4dFhqhQQDbPQfqQxPDe7S849/EOgojeIMZzzqXX6Nc8cGHpoYTh+i3xsoQg
eW4WN77TLxSF46iLCINsNlWqywIuIsIkJyVRcpwFKVqWjUUUCQzHNKnX5nyNScWj
C/3niTfozEFhoKdtwJMT/thUxGH1aiIBV3jzR3zs9uAybw+QpANjte69QaSZSS+8
+fHrlCoMkn4pOgndiSHD67dmLUlOcC7/3gUnYFKwvennih8r/A8oZXz2XA6v9Loi
dRXp1mBs14azssS7JBrSCugfHJfYYbkI5Q2S9asTiaAuElZ0gv0isumLjNilUblz
CBS7ueVXgTyOwZOj8uQAXF4XmbS0bWRQdlkdMTbVRtKGJA+sQWSKj4HEV35Yorzk
/UCHfbdYfoi5MsWNtLRXoer9E3TLy6ViVRvBOzm4C1BiScy/BzoEWzkxLZe9KzhC
hTKZgaVhTrqQ5ZnZUU8V0m5liOjWXODLSaGk4gnSiXqyepa6G3vFa1QCo5vixduM
162DPgVbLpGApTZ7FJeQv1bvp97kcHBQTffDshbvtnZYnAq7e82nvX9wRjjNDZP/
WQn7seW71m5pUzg4kBsokZN5mrPgivhLs+mn1i3NDE3L1GXSOLxxWlq5ss3wTJBp
sECZaiuc0FA+5nRvu6ejdNFeyDFMj3DpmYR3ilM4EyCzmZWyzz4N2nJkC5Jbh09q
9DM3HEN4L6CrFq5fqnb1Um7nB0B3AXKxl2JnKNO6NnjA5S8LxgHM/53sZ+ASoPxA
pA3gltfMPWU2ReLVUS2t5qYz15EgQlfgcCYns91zcAvflBnSt1wq/rD2q7IiS0Xo
ZTxlACBWvGPi5DZWh05sXzEnyaJiTOzIb+4twkQ3HwqS/0U4UI4IdE7P8CE8u91i
tkm0o0kJvhlJ4kk/gqI3mgAPziR5534DxODYO201zXQfrpVHR+ezxUdlkN38C260
XOmSs/9VUrGXX9NALSH//KpP6TAEMrRQfKzfHPoC2kSaBXkzA5QCHJs+Ck6vJaU7
Xf03k8hJTTkkY7eAH6cHHPqezIJfKzHmMGsXKH86OmUM/DqPt5g+B5jgHJUU2RBV
cISazBPrn19epEJGOY6DmE5wqeJZPOKMzfc/TgpRv9RznDaXahjXnYpad6zYj3KQ
MrA91J2UXmdBku6nPJWpU2u5p9sUSzJv/+g3QuAqbQOyYH8opeTzrDD1lfZfTXHm
JD0qbkBeR6aDvooqcCzopusrQFVvzHc0+QPIop4vxpsw3wHQbCWI9XMaiTtNvZJl
YwS3itrvrSiePt67RjJ8TB7e6z4ONtAJYU5sftpYBDWq1/8HIe5urpLyhZ6Jgoa9
6lVtWCJyzGiu9BSdZmvzmJcisynCfkC1/xePbPHJzUUtg6Pki3MSJTMeipe3eh4n
8w3TIfVnJlOWBEi70POLUk1uTvBvIOHeq8vLKNVOaNnl4TaGxFXQXlfsdvzJBIOF
PAZYutexG6EAg0kCg6PP/zlPEGFTn54w4TGFmm1D/lfZmsJLvICDhsCkHTOcoFLl
QUyWJ0FQlfAcgI4pPnyWjV34W8meezUe8Xvp0pbq6Ex5qELVaYmy8Nssx8l//9v1
6uGJHkMPPHFXyVZfPlXH3QNtFhn4xcWGj//0IrZro/o71zWuajhsZoKAqBxfEInP
KM616uoq7PRMy8ffl1Wkflv3EijaRrnRbCNoV//eMfqbBGK6wIQj8paa5N/2Mvhf
TQeVrXvY6orgdlDWfHEDjVUEZHGlTuwy7JhPLo7VVcxGHNHQfr39m39HN+1Dcb1p
0WboBQoNyeKjvyAkaEfJlWpHpIzBlzWUxGcjcVBZlxbmAu0xP4P6/KXgzsSkCCuc
Z9DXRDK5MXBIEBU1DvItIlVtZXH/z+d1Z22sqKBsNp1KCCy4AgJTDwJ8vuVC+xUg
FHKlW7SbMBXIEuRTKq+RNHloFUNDGUZeD5mnXHVKHA8V2qX8MVLcVPxVD8Gqgm04
ZfRK/eCxxWeTCCgFpLXLTvS0mzeUw5LFQONup0x3YkbXwhZx02xjaFL4wGQX3kRR
2g0aRUjdVBmoJFXwexqQxonNKmqQKstk6Uykp63D34eOIbbIhz4vNocQoUgB0qC4
XopYRo6YXaEdOC8NcgzD1XQ/mkoqUdQCjjUhxWXX8CiAMzfBB8nw9jnijW3debga
OcKxrR0SBg0CYWNTpipUP5NQl+ufKd43ViDGMsaAAymRHkB/AM/BPrJZMXIB1Iwp
5n5pZAIftGFjxbCxEQGc6CxLN0usS2SfJC7+gMWsYiMO+mEx6BNPm+Ea1hvONUJD
ABaWE03g9Sh+46QwOynsm2K3YXEs1qmjKpxNjASNQUxW3jO7EF2IAKunjjVb0kW/
jM88dN+PZa2WHbXLS8Ya32WYM1H6Oy9R500HTj2oOaMsWDHDQ2obkOqpE4wxKfvX
/r4XkixvuninLXuVQpkEs8gqOxCLi4tNto0S++dBn+i21gT1vFf5wvdgPBw8bfin
Jg5RX1/SGLKM7VYqe+aJJwMHBMVx71W3LF0y1FF7TlP4YHcLysmRNIJ9cWy0vpCj
uifR8eKe1Gu6lYdsytmyqRpVX0Jv4jug1Qk5jN4YEuJtImFssNMydfascoLkR5+Q
Uzo5PShzByYalGdzM3chzLLwiFNvifY7YBumpAoDUUubIWkvGw11eEUjkEsAvjX+
TiTeVQo9+RyOWSA49uXeQkr7gwIzzitirkZ7otBw8wqGsVxC/9wiY8sBQyMRyVPt
DDyXevEDtoCFndaMqiN/+U7h5DdO4arzYnnpBlPMBubznM8RAiDmHcEtm/GtnC3L
23Y3SRprPVushUxUvVOX1ODOFck15joIWIFRW+jhU7bZp6gi0EE89+VsuXOcdK0c
I1I6DU+mBVl/DLoHzhhcThLfjHnNI9rtqnk4DTnZZg5Uk+L6gTWX6c406sD24oH0
5NfKdD3palX2ImoSDSdWg/9xAwE+SiYs7Qo0onwUtV3Z7w6FDzXMHE39+nXOwBBx
QNvPL+egRn6FhFb/kPAl9rpDsm4FDMJ0rCNng5tvP4IQHOVrYnOTguxRlJkAmUNx
YZcTnIn0MeqzAb6NxT2aFKQ2V93ehrAf1iy9OAvTWDWJBXpenOJwGKB6jfkMc1zf
I5hSWak7S3jDB63c9s8UX8rzEDEPWjQslvotqGEfla1k8kh9xpAVTsdSdeT889mI
MaAUwQ+kdOya/IAM23GA4PpC9Ui0c54bV0eEfq85ik2HiyDJRsORWlCmqcgFv8p+
YaTYzcIRDCHJXulf4XfS9556iHLtp1AitqLXaUKnK40bAqh6S7RMl9WgP8KbWyOs
3SpShxy8jqjVYv9lJPRFyvIXKTzpl3bi2fMjdItes/O39oPjW8LoIni+2+LYYp7r
EqDpe1bBzyJ+0BnXhgmJgI7Uy/pFaWNDAgmR+li6c+6bSEqbZFXJuFwJYWrunrKw
XBe3GYdJO/vYMQbAQhcfdzYzaC+zL4MsLtxDjKFhUBZn5E7PdS4V5QFY8eU7eMAT
aVuCkIgJAUjbm94hVEP3uBrgQPlJP+ZlAwjgCc+zzY53esmyr4l1KEDOkaSTJom4
MIXESg3agexRSsfYudpIZThwbGTHjv8C7fh/VzocZFGfb0BX9bKhJq19PRV4F1nC
G05XvM+DWpeL/qPwsjosQoCA28pdKGOD6s2SffWSq97gSqRBHnAaQXSiW1SCNr/F
eTIfur8lYNy+AdpwbiRZD//IGgSCKEI8KtD5IGDTU/JVJFCQXjUHjDy4zf4BlPSU
E3S/HzGgOrJKGiK8J6YUK80/2rZV1pRIvC7G3LD3UyYmVM1cAAvlNnU2ilJLoxbL
IPyYM4P89p2BVV6gjD9P7TEp5t5QUIr6Zm8TPYikP0AooKV0DcnkSr+QKe/mzpmG
YJl6VRww8pv2Yt1jbKr1R7QcPqD2V5O6T3ptm2MAP3VdoGJXD8xuQ2ejJqxJUluH
UkNfepi+CdDgPFQaPiJ2oHgt60RZ8lFFYuRcbJP+SBGxWvmxHTQ79jPByaJ0JNJi
yCsvDjpxkwT9semfKFKCTHUrkKm7TlBWQyTt3QDUDtPbPl3sv+5isCVeQk53VwWC
NSntir1qT6gH5/aBxvEq+rEMJCQSUW0Fb8/g/UaRHOMQbaGvScmIm0Gd9dBtPvLo
ec1PYc7a5Rg8HG+FOwnC1/tMfDbQ2j5vu4OMzDz7bhOoJ4Y7zDVTh2a/O0eCHCdi
hmeAHrbzj8poNQb4ZlSb2bYjrQb/8L0WC/07KeCPDJjruApcfODtTDpbpvtjtOri
HO+mX3MhDEOOIcjglomgN1UCH77islnFD840Gg0YZISrwitkE0YIIH+az4D4lESe
uFUkqMl0XxMIXGnAWBWug7eptFpZOgDak2MXi8QqL6It3f9kO9BW3Un3jljfuPuT
6AGUg4HTJeHoc7CBpGTKllC8jc7QlEK6TRkohtJMwvfKqQDnVFzWJJkyOSLyDREO
aDEwz/UtSVE+Drsv69QBWA//aOr4BbjzRQd88tHYKaFUb54tty3/tQis+4vygSWg
EQ+T5pymfOyw9H9UB3RAT5rjzNybAOr/irLIBskTN80mAIKEgQToEEUuAig62djX
+/eYrAvhc/QfQWsZU2OKJFPi0nmpyFeinT71JLpX/qZ7ftQ/2WTkGDqq33Z5ZoVL
boYGH4ErGX1gnP4oguOsW/tA+e06v+s3UqtDyR4aSse8FaGBdKriYwbWxKcTKo//
YQAhoKiSq5Vu+kRNyC9gsQGUmSeEluEKbrW4sjsjLFimrLFNbMWDLtedGM8ijcbX
K3ckCucK3eyFOcbhdNTF8RELHZqLDQryWPM0aOWVe3oKx8MK/+n8kRpSVofCXZzr
HWKHLS2fdQAsOTyq3KiVcpc0D7K75QVOVioJQWFtrt8oM3FziOYHsGSk/6bqI5MG
Vhw12gHMn9j8a5+gIdueND5TqEflLpFE3bX7ASlWnXVSZqr8/0dobfwqsrY0qV6n
k1Ox5Nap1kq/qzA7IuyvwyScfFWO6YArgIrMasEJuhA+6Dc5GMSSaa9KURN6N85H
8Kl6/emN4d4YqQ2yMKUvIH6xpcjiQdF5wkQlq59cCPWnPwC08cpj6+H/h9ldLfBT
/ExZgySOLPUnClHpISFfNg/q7DBJx8jWdv7+kSb5h+DJw6/paCRH7wFZAg8tXCei
cT09RXZkr1JwT/XhbBlJ/6BfAycCCD/p7iFHVnhmOHXReEk0kkJn+tNCEyFXzd76
1ifcDqKsTtwMpKGKjrWoIulzVb2HRD2qiXhKsMXTNB6twYfl/JmnooRS7DXW9OPt
EpuTtMr07xDeFAhSbCmIXIxdmR8Bgdgb51pGBXoGN50Vi/604OP5YkFZt4Yhtrs+
7OAJ0VYIroy1notVylrecuoCa5yOKeVoGj7IqxEPU0leyYe5erPbAcJYS5SmDU0i
juyQH69A9XuB6MfzkAarilBT67ytOrIB4Qv+zYt3cXDTHZHRo2pQyjF2KT2m5/Gr
uNfMsvWcz+33N3YOde60FAqWdhHyB8EH0PRaj3XH+Lv6lgJUvTvn6NBbEUwjFn0m
DyHIqC15pelx6DkcAImlga1dDlQqPKBVpKMJa5PR+QSlSa2guqTCRkzfXxhT8/Tj
Q4CIloIvtjqpbJvkRTUzGNLsCcyBuAt62XJ8PG1ZDn1GXg1T2+YZC1D2QY/zxGOb
NnlzegTbWDdRbZuM023+EMiafpmHPfm3j1++VGF/tGMMg0bspwP8Pck+8gG8/sEY
lA+76tlYwV1LKz9wm+WtlvXgR8CJchvkIf4Tcxz/C8q7gWhOhATOeuUExqtd0/9p
tTukPoMST9JqyvpegmkRPjnaHNUnQMZ69S/VzLBByfOT393XS1l7rZJl+OfmcJCj
8O3KbAo3ZwdLycm/Ct2IxVql3dHDIHeKzmkB7GIiCYmKjfVvApdk3XBKsAEGLcJL
cPvwnI9Qhj9WuQOeD5KIUn4nO/Ao3eFUDgf1S+IFJHeoPRRbz1g/peFZcL531yqx
q6xp8O/KLHg7M/U4S6ITVEN6mgMLQ2E5X4T2LavlFZ9P3ZiTq2d2X0kamPdCH29L
Kcr9x7ytaF31wPNXlP24uOtEKqP4rptRWdB8saUxeTYzDmPJE+cdYi2AJtMgqXW3
v9MthkyX/8j4AJukMShuphWpDEksVZrtUFSzPmbkRjojVKtRFP2vGGUFctluZGxx
ndbFF6Ee+qxzTTUuDMvYFi5Q6zNVCFQT+rdIEAuMGFIWU955cjMATdwDIxcEF+UI
D8X1GAluPe8TBEDzR0y2QpeOx0j3LSoQtPfva+NdI8RgF865W0Rj0FAeeCFyHSNI
t1y3LX5+5e7E0obkDu5AvCyYAjAcCJjubNjRdrGYtApLEc65XKnzOG89VRVImW0W
Q5+Wrm2hv7Idh01EnDAlfIJipBboVJH2nG2TfsScCAWltWbTiKatjquaNk7KE5ME
xDXi+YdpiRvG9LU5Ji1MadxhIN7bell5YXZ9FCCZqsSRULtysEXr7SK/BsNZ9hUE
EfYHrsNXzHcnDTRvTsu9HHlRNHqCu/X0kLxV7ym+jqjr1qmwRSsNBsmF5/BzUyTS
fwg2kZuDmSL2L2yJaLJTuWuzDHFjMjnfGbQfUMn5h72Shk2KtUMvtTniSM9YlooI
UtTSuTO1FttDXiUslI2CJiM4HCHV5Q7Hc7UtoD2AgwzZEnp+Cr+o3sx/ZevPrDxr
zstzPIS5pY9UjrmftjWit1t0wEAIi3jB+qRQu63Zik90gPn9A6mXZAbWe0Y9gCuQ
kWQ/d3dbNM4NFb9vVrUxVEbHOaidTsNZctqA8SehRetRYk8vWgDzrouBw/4ylPtp
3sMfES6ErR2z03k6U8y9GZiVYC9OI3wZXLj+5j6fxQ2FLhntFuzywBX7JnKdRdg7
XSVPDNDaRWaXc3pyoCgCYPxHKR6bSV0fcoIszYDhofQGU/elkSUFwFq5KI+sbcx4
9oOS8J3PjKAogGBW5EVy7OwigFZwxk3p3uZJD7su7cDI+6iuth1oKFGuP7quA/IO
U21vJRuPFSU+B7sWnjSJQIKHChxoVIXskAhsiF/0LJYQbJOgFVoX8J61UwnoOGDy
S+rPnfWHZhGt0JSJ5ODJZ0no67xdzddibdUO2DHeCUq/T6iLZWyiCIwPtZn5KJj3
IjHaexF3pDuVHaPwBWW+pO2nPc3aJ6EPxl7aAppa1Lej7PQBHevtDnWVO9VnUUvY
IlEtKlnmrsmSj7qJWD7JSm8+6cv+xtrANJzOrrxzRK3ejMf0XBygzETl4hEBmXzO
9TpNOFgZFJKoQl+2yvR1Jdvr4daUuCA1HXkM+9/TjrpUR8899ZBXS73C6L+38/ev
g3FQDwQQGMf4kyw0aCu7nyHdrY0jhhtxVELfsOx9mmKoaXSDv1Weck3yyABkuOrN
k3q7wpVKviUJhSrLU//3BZWpI8mwy0GAwA5gHsIoVltPtZg+uZxmaT1Z/cATi9JF
iHpV4Pi8ZMhp/E4pHj9doIbgzcpGMyDzk+2kbg84Ijpg+CHkIUNIiohyJ4nYpAKs
x+nb1kv6hdMcSWlPM8YpQZs0qVAlpfWRA692BkZ48FwZTJQG9ZJwb+XprLoG64o+
CXn/xPGctE5/CuiortWU7Ixd5yfPeALbfvhFVOtnL8+oKclwUUA/zYPrgCDomKkP
SIwsdhuhBUDccUtcEgfzLh0DVJEhwlXwuUyWv9DpiLo8FDrBYNueRDEMcJw1XMm8
3IEuqYoZpG3i9xt1AMVYQFmfzYPtaaZ1a1Q6gWDcJUvzs30HNWpLiKoiMSDQ5g67
IteOgzCiUTzwKtwz69+7IjlovMHheOjLvWv/yxwpQuAJ+U/NcInzA8hamB1VHls8
gr1glQwVhfjBzMXUOfmr727PJgRG/d+7fXLSjo1SpZkok87M8RSI8ajHElzxbFlC
pXuJypi/bIxMDJ6bzeh7tQnnyFvZTaSIvRdenYUiomIj1dXQPrAscDHUAvQGrwFt
/ymCWUcLjhGkmwvoE9+uKNvVUOQiwnl52X8n14Ilo/UOsb1NFxur0LNF+emmtcWk
XgZkCfLOZ0lclkiOHj5bVt91Y/4nl1OcoaAe392ZNEXXzbtKyekgY4ecn9Fj/ynj
82tFWUQCHJ5NPXOuDE6bgFGZZ64MmB9xxWhlsXrxzyUxWacWQvfXFLP8a9L6JtEw
4XiCBGJS5zQj6y0pyJapk5tDEDswSBOBRAiuk2AsjdnDb2j4PoVxfupJK63EVIOl
jsyuwCwfYtdFmNkqm3Mz1HSNkb9MKt5apfnaLDWtq5s1r17ZBfOfCapAiE/3m5Mi
lgXwEY2IgJJyhQYcNuH8fBVDYT6UZ1xqI9G9JD2XljeotoPYnaD8PFfzr6nkRGO9
vULP23zD03brFTXfxPlPoeqNghT7yhSjVTAf++I3b8VLpNLIPxDp0Qycfw2jT0vi
t42RG7BmGgxi8cz4gvshNvXbhmVqBZnRGUFUZS+qznKk6Rjv8sd16y1PcMTPnJ2F
NJ8D/g057CF1npJmYX6c2RGVO/AIloQlXLK7SpcXsFpbZBByNAXuzjr0uKCaZvfY
iSSteBh2YcZnljMqKDhyf06Kt3Ps+6mXqkbbMOmCt8OZXNss4IVv7xohwcKDfM/K
AjVBxoUFpD+gufz8J1mo//GDnuNFhbBelKOM+o5L5so4ZlJsCFlNj66Wix1iPMwA
shVX88MgW0Mk9yeTz+InDA8GT28GXh1FtjJcHMsJxdAkfe37gTvYRdpSQf4cG8U2
6XWurFPdl8G5VnZaQy0i/6XtdmmYsLgWh7JlceCdQJTCVq1K/aidKBLqWFK/8rLP
RdaRFBtoersCaXSQr3yuXvSpgsy2T02Zdj7ttYHjMV8LwoDDJA54gbiePL+fsPmK
OLlDswqRQNqh34x54+WfNQRFCe7NLLQZg+TKElTPIbaHUaGt6v25jQbGqMIFTxEc
zcwAadTxio/3c2hXpV8Div8NpWXDpy9L1ZI/pqM/vRIxCzcGJV4ON1yAgSlDWYTe
OCrVCTK3q5GxkjasQsxUZ0G6ucxg4wF2B8csUWr9JdyGGBIQeANtKXsevXVZ6yvQ
AEOFwHgXAmYZtrBqaAW3IXOkboZUblgLiVa/Dsfv+ujsjF9C4im/tkD543b5Bu5v
KnR19dBk1Q0BQroMLrRgdLAuWKBeYlSq58CgZk+k2thPoz3z0YjL7omwqLwL9pCd
Ksjd47eCV+XWsuk036kGI2hZhKpFEbe9wjPwUqAexc4IIDenGU6f4unFUz0Ewu/g
/s/D3+lIR69FIwWhhcqOm+jMOuRLbl//W2uTRO4NSPzhZKIvsi/LphkuDCE3vGzQ
7OeH3QEvqmtl9YVExdt+7fWMnmivcdUyKqHSsKDduWws7HQo7kzb6Y3TphA3uFFN
pSaE0l6lQ7+hDNhF/i4wGduyATNBi3UZU+I9gqJDgB8rPIUKCXexqHl1jE1sDjBh
AEhDQ4sPk5t43MUj03bx+UKqKzGLtuHPaugLHwWeh/htdtmmuxsWji8gQqHKSPKn
Ob+F+SbVgsDJk8Ex9I5FpkqRgtg3vgSBzW+R7JdzASdaLKaZLMvWEZVlznwm9Pi2
VobmCq9PxPFIkdlGjJRWYt+Qq0FPJWRzcj6E6c+BlgeCTiPMjEsjL44NubFKarW+
2tN6s5lhquzsu0Hs+ffKCWdjoGp5+LMXkQfVvAoI4Hdn70I4NpBMLYVArznqAir0
v5aZoWoMJO4b0Ajk+qWwnlfqIYByS/2PrLoECD4kaKnCJC/jEbxvx0pS/dWXKPFI
G/pAYeSfQ6vNmS+iHRgJxcQfzanomZWmWIQqg2Y2iiLbByQ7cNcYW1MD3Cek9OIS
npqfgFkXtF+ZhjR631pqIVrosb9uxeVxHq726P0BJ6W+SEjGdju4dGmd2kZMyy1j
fbsVKoJdy13J0lVzmB4YQYjv7bvski2oC2t7uE6kJfIZF9N3g1rks4LPrwFgxbrb
Yg4c9FpfF+PRTIXMc8Q9BYfaifTdC7GOOM1ceQGngMadc6txafSidIzGEBua3VrH
Q5KmycOIltgxmeyJhDtckKE4X8KRhOVb74xQf7VtSP4uRIHRHsIyCyN+VLzdfwgU
ShfvVSaLF2B6f5Q1D7+hAM8DMCHpLq5v3cPBW4jLqAaZxYHefDae0/juLKFcYd9I
XM4BLl2ylQtPHsUD5yb8B1MfvBwn5xcicOBCIVCm0aSCdBei60Tt7P0Q0+Pl5XpQ
0S+AknI4l+0P9Ns05Bh8TQkb2/mJsdf7TxdwUBqCHtwUjC459cUcbfqD8MjIuCTL
/9bCIv1Hl3/PnRtVOvksBiyXrK/wg7LHpRHW8b/xY5GFpUtPXo0mfrTJqMwv9TSV
rhR0V/9ewn6OdEDPQSBTgWZLVtNJkow/wncY5JcKMlH7L8V2YR4hGVbZT65cIpUF
b63a2n3nQC6uLJQ5CQAG8uoqW5Vrp+fMwhdpBabIEqpbVS5PWLwN1jEkPzrUCWhS
ZlsQsjdpflJ2RQOWMp2XW5hylUhdk0UE+Hx/gWdlmvb3xSJNTR2PekIUqoA9SjM6
5DhfESvuaTg0GYE/UC2WfbCfzPUxYjbyi1W+2RZEdzS8NY1pIXfDcDloUdW/QBTU
M2R831ZqWxXaZhtXSCsv3PLHN4nxbHvfzNCJfQpFPl0/ilBm2FBse5ee2Qp0fHkA
7VBQAInOvBqzD/2mapxIlwB+GluxEg7vbzASvM+7lQQcgEW1OQHqwj+JUi3voxuW
hPul8KuL1IHYyVxyxUlO7RTOV3JjO882Q3pgiQK3tC6mYy7iTu7EOVkAHiRKIelf
CtsycKbYaKLl0an+YmNutZh51yBat/ZS4VgZHmFavLUTPjC4sDbw0obgFyN3ehEo
cEKtN1C+at9mkCzeQJWw7h2W2K/0puNPA8fCeJ4SgMge2zqDeaUPcjLa+Hp2jayD
Gm7FQJAK7hsk1S5fl/4VbNgMYnZDYtVJRVQ9xwL2ImZuaJWaaGh5EvCxYDnhHbT7
/5yzRA/y/eeLmBN84WEPJnSEWYkHHaGbwPkqI577lyIj7Ve6Qr2FKrvAUAogXapv
3uwcdbfG85fkvT1JqMf3rxD4hb4ZGqvTUxOX10HpkqxZejSNR3SWaq/FSzsYGxYA
sNd9s2YsPfTI8WVGXG8jK7WRR918mS+rQ4rzpE5+4ZkG+HwLUkPPMwaWZKT6+Wbn
p7OD1uvFbHYLt4wrLCbVbjbmc3gtYxV5NRU11gI/P199QQD2mPIJ4Q6/tGGwaiUs
A79ALU8KIsFAYwQlcJbPV+5J9kQx74A7deZh0e4B03Wy3QZIfiJCftJTbKzSDRbt
lutQ+AygwUQh3wzSrpO5h8pyd4ai9gA8aDjsfz0a+d6NY9JP6qJQeZyD+E64ZuMl
Sjh3lHPUPEQvP2ifmhq0LNSQRG3kDIAxxHAk/1t/tDePH6Gvog3byeTbV73PkUMu
F4Meg9GmxopIcrITw4RjVlFkUqkGUPV5dQWWnLLRkee6XBC5vvTnrnoZg26UzZZ/
zwoQjj17VjzaHTcoohUSkIamEXYiRQf5j06ZAF8kfAi0CSqWs8qoim15M7WbfTXw
CRYak3BlwzZn2SUXNc7fSaA3M+PrB1fnTT7jq2SH1OYQLo11pWQeLJYIDlWz+reP
wdCy6tYtK4wVZxxGAuvacolOCOLdOqqMyImY0+jQfpY8Jcdd/OTQ9aOlAYboR/90
ukUBD2+gLrXrRHqDivFkbUWeSD/hHOCi8ntsqZFK7wdEWaYG/OpA2Jhttlv0CvMA
wGsxhL0nPRGRfLhiY/ReMFAmjBE11hjuginmiIwmcFwszmLiWQHvsjUSvSvVsm7f
aNJu0GidnIHWUdrGlawrvRH22EbwPJn3QAERGaySVC4H8smcj9eQP6kGMD6e3vue
zNXKUi9AEaVf3px047s3f8BGe68cmZu7+/Uiiv7poFS1nBCtzJb4BZLUMP2Ad23w
2w3OZMvMuamD1lmcHFgTRbRULtGTWzr1PYgLT4Ey6+Q/t5EJz8G11/2I8LL3wNiF
6t+e/cvIpAUaV0k5lFP0ZSMffc5epzWnh5x3Kn67Txmeb6LgtaR1LTInq79AfRRx
C/y3ZyoQHxtxaLXvx0iuhKSTSeTxFIo5oo/j8YW21oMuytQwDoyH1Pa1Y9aVsG+t
NtcoC387MW8jCNOH1kr+XneCM4wMe7c7EZz8vUJbnSRu5zTtx+sWNB9vLLVwAGfQ
Zh1ozsMWP3FZIUbaT66dAfFPDqFnwjfSDPnAr+4ikUtGRlk72dRckPqeW7A8w3fb
MLRcQseB4A64VABOODUPp4hDkDRdrbgTwLJAs/U1ySb+9NVfy0Fd8IwtSqj2rkgQ
yayVwU6kg0LjpVc1OaDJ3vj8FAAyR2WK8p+AzEvCP5OoKWcIsbme0SozsFsLfHlw
lJT+7OIDPrKkr4t/RTnFuDPwWDR4cFA5McDu2c0BtoG3YVYr/YinFT7xIyXC4cbn
44nas9smhnVvOh4cmAmRldSwshScRwL9wjXgnqdiGaQCTFVq/8PprOEaOHazAumv
N4rAIoPa2GdB9EtZkHIPlXq2IfFR3kzBJW6+eVL6p2SOIwnsZmygMyXjR7oweaDI
eq6Wb3i3hkIYtkl0Bjmt2oxmNdg6XyLrh9DdmtuRz/ZrWzZqi7ZXUnvS/C4apd4g
wNvqGoBB6B82ooxQ/K0eUzarN6QKdp02araPIGfHedUqfqYCaFV44JOZO6ENqERY
O4+Tf5pV1KEl5cq4VFFjDXnwALSPs+OEYoKgbG5mx1i5kNvsYKW+JsY5j9gFdDMW
fUZaYpxBa0Eb3JvLJdhV0ToDh4HYuGc7jOcN6RBmt+nWaejNtGHZnBHFquWqKrM7
VCziSt4Tcsn+2UNlpqhjQOKEc05olMKZsZ40QokSOfw/yP+njZU3AtXb9ar+D8Bl
ZydPDmJ8ze9cV8OCyaIGzenTX0YkJBB9a/JcXfP66QzzFxRV4t0v7LG4o+Ad5OrX
y3u435ol/nCRtoX+rkkpfVJDnPu3CzCwlUHvrlhkoFy7uhKBC9yNeFmT8ha9z+8p
SoxqAwUUPjFOaGVxZz+dq5mL4YTYFXV/cRgBG4/fv+6E5MwjXLGujdpZsyKH5eRZ
xZtYWlmJtDURiZ7axTr++mxaceeM5VD6e7OEDu4jtDSphUHA4QtE3vZOm9n0HNlY
UC7+7NmvTL/MWTTy4g711NI6/c41CwrqSVwfLLKTdokNe3mxt6iOmPSWAc64Ek9n
1T4sz/Y0wC7C1fyy4towZLAwFoIFEa5XCyIjzK3DBpm0dqXJ0p4NQWCpqb3lTixf
bpMZBjysumdVZ0D3Mr81Jql66ctA/GbXLAekY1RhLCdi7Doojy4h2Qbk+yOsHFmY
SOfovuTw1o/G14gTVLQu8nxBOo0AhStATpCwd5K9c3W9ndJ9u38bs2g3ZTkQakBP
mkQjL7ZWWb3e31INi6tV1i6CTO57mFZtdyCsuOfe1ZeVsNUgviPHOwb3gMfsuaYQ
ZCW6ga1FJEa/imsvAKEqamY/qeTV3cGuOuVNe8qhkeojb4+SN7s+ffeX+szEUh9z
f9peZZu3QHfj7Px6WX4PkRgbXznSz4zAHUqVMB3CkKW93fx0ceE6T2gwSOQmX+r2
/I28qsQmWa37UJlBY+mjwzR9DLl1X47KN1RTl40X41TMrk4KWGhUnFsRySm7RErN
t1dGA20/5Gp16TCYIkVgIgKdbCsChOnWhaZTJRvsiajGS9gKSXSt530ERHl8JkLq
QVeu/79vMq2asglxaUfjrtRj08efvjmzfAc71nDtBTBxVCs59zCQV6GYKyuZDB3u
3LgSFhnvrir6KPIz+K3kWwNKq2PgWPeBYBz+0R0B/6y1nnujMTMQoFaqYMr84g6A
cAYief8W5Pm+B7PyDJK1mtgP12bS2bj4wVx6GizZY6gcKN3anztKLxstDxrWtJla
SgwGUwYXzmfEQxVbLpOaAK6VOzY+BGp1D3Obq4S7y/NUUH0dX91L8NUGC86iWcal
4MPSmQAFKGOLLZO8pZYmuPWg1DH4n9GZiq3C3CHjIKJmHMLQUnudonNxzOTPgEnF
/B+sOtQvM2FRpfKqI8PdOPCztHBlnwsm8JmiGazZ3GW3P1jfybJQVnt7AskzBOV5
CmspPrgCFoDrykbxWDH4tB3F1jncCQzoYtsXQm8v0VO6Ziflqk/dnjz+51UWdW2o
bqU4Wc1sQlNsHQokjX97KEcH7IvifQnCK0zfeQvkkgyYH55NNw/RiE0UhG3nBzdw
a+jYAzMXX9HdxyJUOR3eZRPXYsVY7GkMQvsQ8sSmGgK3tfVd058QD0648V58uzBP
RPOADnuPDJJwMwj9HDEEARUFYiJbzOZtRvAYxyPlcbS8V+rzuyI+Jf58ZC7RhD8h
P6QRTJLjN6hrsmVVI8H3ClM1mTTtRP8p86gZ4BQWZDRN6N7JgO6Kc1mbJtDHnzRZ
M/Wz1wCGIERbIVMfsuyNB8kdnbPNmDgGSlKNBY3t1y9DpRKLZgZ/J3d/DaPlkF+e
uMd73C+wkG3K9fLcaAUdMEynVC4XW8xwkJxUor4d1MKDCg+27GoJ7MnVKbK16knj
1rfVQJ7xru1uoqyDuEnPM6feN/6eNz5JYkwDXCGxSI+SiFc+1abc6+F22tC6ZU9h
WV8ZAcAfAt1f3ngYMoBb89L8HTjqN3kO1eBTXjjDhxF5d+o3EdoSlcH/desezDMP
xySL3ezLU8gv9G+bGi7fm0cvAz59CPCmIAtvzJxp1/XRr41MUTErxcG3Yh1fpJXc
2uu768fgdCE3X6lZJydc0JoRKufNpvPy/tUMbceepA4l0laC73ZR5i8iKcHOk1BW
0auEoG4FWC8ioUQsSEUsmqPNhyxXb82vQzB2CdFnJoIARhR+cKIyiqI7kfgKY+zG
tAERqv34lM/eFxWC2Y/w0jMUERvzROv6DE0quBBDAPeQEVnfscr3xhZcoe5f1s8j
N+dA8UGig7tReXkC2p6Wgfa+biWmP06JK32VUu8N7wHTh2Zqb3qmUdIjdUeMBd4j
Nxs3+raOhxhUFqagL+m3K/2dd5QqQ7IeDKycn9QsBRjMwGWsSMLIyPNaBbs61Hhe
BhUe5zwGmn+GYBIWEQD55ZG403ezm/oUm57C1H2kmscjuQHXoxZlsK+sUNthYRTu
hqQi1Vih4KSPwVlZFeYrYGkaC6Z6SBswWQS6U+95x/JMExEEJtp5zc8l3P6/2wUZ
dvAqGWR/SGDK1evvYnkWj5Sl0NhCFCM9+wf5U9u8pZLwWcmLUITJQCfgBuzFVuTz
fr2wnOdUbVsXUgl3qW4eBskSs7Bt5h7l7s8DFP+Ztm+g88dZQ6CN/SMIoEBrEnl/
iW1rIddzQnTTLvIOOBOaj6DBWWK8FcNGgAXEL3lot75x7ljOYAbN5myURPESzQ4P
jaGf5OUGdAkv4aTiTTMGXz9S2w4vCnjERlHruuTW1/GR9o3V+/hGb8y4mQickIy1
FMx/SVGBKCMXxF1w/EIc92L5HAQjIBuw3Iq2smBhxrF8z+5KDeB/+HOjiJjpT8lp
hQfH2R7B6nGeaxgz24CCl6R8FUrSfEYGpyUG7NrL6E/pLaSphqyijL+8WM8iTHic
GLN3b3lMM92kDc8WazYmxJm/zSa7uzhh5fod/hDaKyw8HjyfD2y8v5etGPU3AeRI
BvXnVU/jJxF6qyc/L/OcXTVa4UQXnoB7AgUuCvqebVToyNXpVijq9EK4s8sjm5/q
nGicXoprpJmSyJCehzeUgQpqqztmSdFRSSemO4bIGOfp5L0eS22Zw69rFe/Ztbje
WbGiocg6eP8Zofutmh7gxJqLBqS1XI63oY7Mn/w9cpu1RIWG9EycuqoMYJUQx+hJ
G1m7kvQ8h5hqdsOxuyLjkO3fKMt34raxjt3b1ni/kewrTpK+fyLYHr6xLUlnJ3vW
Lnwe0XmOESdyw+ilDL0SJ6CQQhCQQRqtEAkIlu/f0I11/MqF/ufwRU7isKyCCYhC
4XGSyfplNneGj7PQTrDGF7kejHlUcv0U+RBF0za97mzilu9U9crz03mAHUzghTgI
1JArtWtx3pTwBSyzaelmqpQJRAteBkrsnpruhtyEslxAjq4DQ7lgG6Z96P+Ud5Dy
FDwcug939osF0w4AwNW9uM7o3lF3xQq+dqpjMOBReLbgVlH6FRrkMpYBJlegrTUR
wx4AF4MSlGTbZH2UVGp+kWvhZXR+izJWUQMFnyEC2t5NRD85tis+ABxwjWJzfhRu
xK0o/s8t6aEz7ypxIFv/q4gb0kvZ59HRLlpVWjCXOOYQo6miA/GE/hPOvjhdK22L
xANH3XlH+0MZg4m7edspgF/EBBYEUWH4OFHMdSzK36vVxXfbK/nM9CAD814rLupt
NA98Q6W1RcAaYJ79tNNqY634ie/dGeHJtG/QWDIzGJw2VRzfWRFbsJboBWb3c6vr
l/1qexc6rrfAQbmnlJcTC1ILJ1VzgfbFXBbdP8aF1kyeMTs/XRg8WFkkYoHe/dIP
C3OC5tvPZGOYViuF5Xu9EjCFo7aKINLs1YuKfa7UN50w2KXxq5KXA8auBocVJblT
OggSF0V1344EEJYOgOFNxmzxN6c+BwJOIwD7/D8iLTxM94fcbIsZTogonEYT1D6T
A9W45Uf+jJUf1waw6NIrqbOXKMoyXNozzIXNdrFcQ1Uevm8uqSf1JgJNftEz+LuZ
Av07AR+a44UQukwNcAtO7ayv0i6TyDiM7iHrVQg/8eqhxbm9N7S//qgGfBCtsJc3
jNvoMJD9R73X1d0SUMP0X8NmtoR48xU1fToH1ohndFhiBhmFDsc0v3Pi/r4cFmtj
4UX7XSHWeaP1FLEBOVtTArF+piY7em7NxuVs/FU+Mdb2Py1a4pGGMwaHarthmlAT
r4CV/HL+4K89ZMAVuBGQq4pdGSzGTolnNzPbzrbQQ5WpIjwmGT1SJkQs0JgoCNKz
vvQ3dgFI/ifSEaTyNyBnu5S22ZLjD2DHdjzjWQj+L5zsYGDi9XE44umNRdpufV3k
X/+qtIPWZLukyEVPloTZxhiHpko4ACXgZlbxl3ZTF9WdiQLfs3xzgnOutOQhzwfJ
0dQH2vBK++dZ0WUEgye+hmK+u8NT+pHoYTmPtlRn7gRpESPqhpdtnoIc036+f7bg
mnUfilM1KF4Z/ds83hoA5wFd6CoiZsMlVd9cwGqHUre67qxDrIJL+I14yThMnQdk
+WlQ2VWY4udiOH5F9mZIXhi2b5+npGkGIXQaXTaVrVuhprJYa4LUf3UFiKc2usC2
R9871950ZTJp5z9Q0J4XJoN4pZz/QzmGewmbF68PgRxOf+V8eygImIXqjhMw0bTd
s+7hGPjfs4BMRAg5ZZGx5jtamzjbtPPscno8Aucs2jc/rdK7PAY2JFHTmVI1Fojd
lpHbdSPHsqO6HyPJzGRYGHaVe8m5CFsyTFpMeUwaHxWcJuxjGn8fJp2Ja7cBNdRV
llMtlRSTEuRXusUe8RE7PbQIt7y1AROOGByKmNlpp0Yd+ux0Y4zjWJ+C35NyBAuj
afRow6CsKnzqk9z3CmFub4AySwjQeWyZr0vwQM6KRQGbOzGAHJ8+3aSKqz1VjH8R
9YHy27mrTwXu/8WRja2DAABvsiyvprEbkeVYXipmeG8VSaO9HfH7eeOmVvVGda5O
DseUxBq4giLDbYGRXUdccX+Y+jhHy+3ytSAi29pVU5ZmVI5kbOZu9ieqrxSegCSB
EANu9QPajjQPOF33/kwwkCosQIZtUgU8c9Sccf7FmC4Wd/2182D8b3TVjuyTeI2R
arWM4y/cbBsKvdnyw/lGakwZ2VtWRvEo5Z34zUX83ZZnmYGYzXGNV+Oq3Dm2Cpbs
mr/TsCnQNE45uTTCO/78BlAf8NMiRM33BRAHVLlR/vUpYh1+y5bgsQri7nSG3TtI
7u/sS7WsK0AfdZAKgW2Lh4x66Zuc7/WNWhXYi1N5oVqsBnIE6sfXAw1qNUhcer6S
Jpmq1LHK/pHjZ4y2jRtaOAnoq4K0H5KJLaFCGQdNpzDK1NTQL7QSI1NtvlRlDmpR
Uia7A8mhpy/itKtowh/9yWBZLYpfDzmUqw6ojlcHux4ta/cZjMPE/rZAWAneYXFZ
I/9tVkI4SJwr0RSutJpAAHwtPTSoWDCq9XcEONFUnKeAyGkl5AJr27UqlitjaKUR
W/3v3rhEQXZ2x/7N2/o3/sjHV86WuIT+hYtY9WUjnUZ3Y9U94kIU0e7tqcNSi+At
hU7YIRTcXgRuFLaNGubu8dluH0+dNkM5RKrdy4GWHvFtoFA33yrZ7Gtic9b+kZ9e
TPEkKTZj1gnU5Jn+SaMShXVBB5dk4msuUPtNmIfyQV6/jRChaDEuT7EvAoKmXtEA
fDb/HxR8OmTuiiyiNl7TA/PQzU2iOhunaRIzKdu0oLebqRpJIu3LA9FIzhRex3a+
C+EgaOO6HVHD3ja9n7LqRj18GKN5N5lD05sEgaS9Eb99dW1L9GdOcxMQ4zOARw58
UFjd5IP270da7F3zkDGhsX+Nga2P78HwoELLdgNmcI+Xv64Z/chw20ncW1BXFemo
hWjDSj5g5IUSn7RbpVUYy2z4WWZhOEThR6M0dPGeKO+LoB49CtTmc6G5XgGXZlWC
5+yENmCjiPOIfyfoZiAzFpfsEXp0Ukpp45682PdsZ0DG55u8LikAqG+9IfagRckJ
VflA8jHmrCC2ybLOuU3Dt7Z2ybVR5mwo6bHXfbFKU1AtvkFakHCx7D5BBOoffdX1
bb0MTHrWgHClBygQG1jzV/aEm9eZCPKAH8Lm2wbZ63DvAdtHm9tYMvKEgyqG8dlM
Aq+940VnfpehZtrSKu25+V4Zq5efAjoak7LM1CbgRjRtmv7Uv2bvvTmqtvx6rn3o
A4ZlnxtWmKgdk849fq8gpDV9OY0dp+Pr8hIajfTnH+HR+P+r6l8W0BXUh+pvkFjo
aMgt+QkTsLvJeaggZ3ZqysSIZZUtd+ZPA2I1a6uCTeaqIC2DXGIAzv3GdZ0miCPp
McjvCWg1LosPd2SuQvNN+IU/s/5JHGHs/fS4ztD5gaIv0K5alU9ZxKPT1BbTwv9O
nsOdN9ZiAhu2ZVV8wYN62XcT57gyFelMIwz38cLETmz2O+bSmg2A1ZDn3C2SkIY1
LoaFMAxEqc45S8bUbM5jQGCNSd67DRiBeK4eGP7wUod/sN22lRse1U5tJ2mAnDHi
3zjrdOqoOlUnCDLIdGCHrW5LUszWV8ryYhtxaCaWCU/rXnnrPpF0uq6Q+f7eDTw8
AajjWxpternoj7WrSTkxOcx6PNLbl4eijo2hKKwRLHrAvKG865EjzKWMEa6eO8uO
9hW7t3of539kkkuNIQeSJf7rKMRUAWMO0OoWHPFeOfBMRo2/uoTzQayiPFOC9xIP
yXRQfWkyhX2tz/uQovguev5N6EEapgn+AReB5a4dD8pEEiGkNDNMC2cfgdfkl96/
/SHGMTF8MkJ96c5BKOFdnBiQ3QVEgOI/qCISqJ6tKr5d8B1peVQmY0uWO1X4XenD
oLcqYP2xiWYu7/qRiV9yEn/p8PhAobWiYksg+lJxGIAxw+pldk/G/lRsFNIQqoRD
Rxg0m+yiEjkbNlGvMVW1LFYuTN2VN+L+D2GobllxS0oCAZgROFBbzTC52VCrRt0x
iXrtnLYbA28C6Jt1hf7nZE90oRvjTv+443VLMj7MmV/3f0m1R8obmywSk8Xz94hy
vKpjEWsVvDKi42t8eeAtCPMaeVn282rVLaBrzYmcsyDC1J737TeuNSPqAg2w8LVU
Oo77fUuB0e9Pu1nJe5xpPKE9Xdt+gnfAslONu3J4CmXtv0q294Jb9ioxaf89J9Cn
yX1VrGmXnl26xdFqYNwDoR1mAlYbnHfRwwcBvs7JENyjoeGL7X8svSPEdVwjy/iF
ZfpwdrNcWd9fEaQKTkg7VhrmdWt32YHRnHyL46SGi/quC9vaByZogYPI+B2lrLvs
W9UIYG3mpDd0a/017mMAo/gx85tDref2Pp3gECIa7usJQ2k4V/AGjHSf0tZ9Fsrz
520xJSnldAbKbGc/moipveRpLwhcqjCxWf+aR7Y2nyWgVtdcu3vBZtFZo1sVfcI6
v7ss+xX5Y3jC2DysyDL4raI2eE6gVbrxqBoxQtK2MY7ECaiwuAXxV35ze5J4N8tb
3bp4tmMKwsgEUw3kz6NU5/F8k1/e7/Serc/EpVuMSmaRf8SEAQIQ7tY4xLzq62K9
0Now6AWJXiar0dlNPLuaEh1heAh+B48vG245thuUTWz5uLBfd+CAkLGT+BceuDZz
48LOsDiBjw8Vv3AnaH+iAZ9l0LjkFaxRzauvHT8XkwqnhgVQKG96FXOIquHgV4xR
AHwQMSicUyCJ2WY2XTiws0O/cqF/GiolahlGgjFmuaHPxCQJtb0ca3V/z1K5IBMB
X+mwAj6VoSpnhvkHmK/BmzUE4h3VRh3SjK03e2V68OtkkCln5MR1VrC/NNcDcLp2
/0rtAY26zoFqJ/3rDqmqyChqxqQ3F4FJ0drKjB98JbQD7bdlUJZU55bj1qcrDLLs
hQ8fzpFvEHFF3PyBK92wmYJGiIwi8Ik81HxA2CwdOkWPolsjhJmcyVY8rUOW5OZF
U4vRp4kaTCUSbX/EQr64IBf0KQwuSju/oYWvz6fiYczPqHt+h2/i0MKFEXWYOcTm
/HuSKgSXBPQ0o0ixaCRpQj8mk9luO5Wu2YmrUoy2T+HrZq5zSELALO8nKm15XCfR
AAvOBXep5O3FVjGlTDDFk/I9PW8+SH2Jp5h9MyRypQLWHN3NPZLnboSg7BZ5wwte
4/aC4fNcQjwBQRm0CP+LCTImezf3Hb+UTL8ByRw7cjT4jNg59u0gRqkA+4Pin2Ik
VivBjQpayaCo/csjCDdORD6jQRQ5FbR/QSQl4r91OoZ4KTWOLDUrZV1A3msIWUQZ
7ixsC0ZJogvTJgasrzOXts4OvIVfHCVj9bzRQMzheTLXLpkC8vDLp6eAu1Orxnhn
ZqlDW8pC25kUaORQ+IxqP5DmQGsTauxDPkzmpuSFrCxSMdHC4E+fUoKHCqQQdJSx
CefLshhfGYxbV72/TFtzG+hZr6uAxJ8SJMDMNyvmB9OQrYSUOaVbAxU+zSzvApty
7YqTSk971cLpQ8c4Dc+ZMLpELbX2M53st7hvOeBsco8YbIj5QT4FvoadpAe5KLzd
f+nGbrqWLLkTt96lWGDTUDwolDCFystP6UHEPikkwM8q1DxsMDftkK8QiBagXNNN
BQH/89zU9OGP4rL9alwwh5dNzgPmvp4AksdRt69IOE0jAfZcFJb7F23K4NH3SzNP
L97xx4PRr1Jfi+mMYBOY1w88asD+XlXf5OXQjdYwxXSWGUrI/kgPWUXpfAbk8VS/
ehYvzg/K+cmBCCH/W3G4JN+sCqSxgHPoqmZEv+sQsz0ZMUGfae9AKJFrlaLKyhsI
xMVe5MHhUZAVWL6vBfufOzcCpbjxHaViF2SEFx6IpYYghnLsQDpSp0ZtQD8J/ck9
NM3NVq4uHTbe/D1BG9I7/EfGQ71w7pjac3l1aa72KWA1dzAFQbp0c/szOcklkgoi
8CaseQgXg+H6xeHUW4LdjSG7PqOcIiUziHV/aE1v/9D8eTorbCEaGLQbp8QR2k/A
5XXGM8xc3/tjIbPYzpdj4hPBDcEXFjyv7U+jLnOlVD+Wv/pK9MI9o3VLreVbm0bj
4UK1f3IM+8mh5JTd26T4Wkh8+RdCw22kYNiJemrIsuyHHfTaEDL5iTFr2cpJp9kK
NNrp5B6DGsqs75NkaE3HoCZPvSlnTsOCVE8EGPyNVFkrlYwtmi/r1sptH7D8eMh2
U84kF0X11uwheghvDDjTGpt3PQ0Ro9lRf1CFxzbvkpMjvHJJbC79QKLNjEcOJCFs
DOZ8QKLHWT0zIU8nGsWtWqHkR7des8Wm4GGuGFJzbD1aoX0zmL4B4r0U/oOpwKFJ
dpfyyw+TSLYPFNMr3H4cMre3e33yB5/FnFukuFx4LoqmkQhRYtNlQ3DY+KoQlC8q
X/asVE/Rbh5S8UyQAETQ2MoqXAN2EOGK7MRP+1VGL1jwvmDd27sOpIxqckcyMWE9
ZmQHl78D1gsKENUHu1plzl1MLILM+QKL65pudUms2gFKJMzeUINXgOc++c0v8GXU
7d3NnMHVNWs6ogNhKxO7CF0I2Hz/wLetdrZx+LFsDf20QIA5xGmiOScX3gZOAJJX
FH5ahROjx5zo36UCiDh7hFxmYp7F69udTL0sQcSU/mVZ606hUOTTt5vGucU84sEv
SPgAJlmABVVcC/BDLH3QvNpzlfkCCuUS5qlIV1Skbvrh9GY2vlorTKtYhfeFzMNQ
SZAJfg/+i34S9T55w4prpn+6L0wJ5rtsN0jQnhSemXg18x3osdIiBxnH7eAAWUrg
oC+N6ajIgYBF6H7/jdYVm8c73gLkCArI+lthUI4ErSAr8oeY041lx4nadNQ97lRq
nC/O0r6J3FyOcn/8i0CHagDzk0vppC1BeGlQcv+egV0lJ4Iw8cCSIrZIL7evFSPV
btPCE4aI90nB1ZkPiIF5ImwgPk/SUSjbzU9TPy8HJ4Pb2WIJrY7f//ZlB6xUnulF
g4svMhTOMIb49jW9B/GTnqTs6k+UBUvBvhUXml6YXM5CRbQlRg/FlBFGrkPUqpK8
TlhoX54dBTfUSonlNM/uTHyYgUPd8kerWvxrUhmB2SJs3DbsMKHezipjYxjyGY2a
CS1IJtskzxUTkWcsvZz3iosfD/U4gT4LEukWlHMHYcBvBRLVudHquZppeiMty+cA
etZR3DoQuR+Gr8xLJtLGAK/hcOaTsxzSh+5yBrzkYTc0URdaJqomCyOKK9vyiLk9
reNrw2NO22O3nE68fHfULg5m1EsogDZsQSXuo0R4pJk0qSBPs3mj86F5Z6NJxVvu
/k1/mig6+nX5UGuZzV5sktDkRXpwaK1MSVXrl3tCUVloZFXbSoF6QQsnptaAnm+r
f8IXi/0ctottvKloYjTi3hLoHYnNvrJlcbWOnQGXmZzBA3DJX+xWaU+VxYFdHu3l
VVeohOKk5cqfPWa5rnKiPG6qQZU56BDIovJLlBLSD2lw/r6Zd7Ub+ZYYK+f28f2/
FgSY0TVQDXV+r+OQ/4WMvQIRtMgGGTPRhbOkTCg1uoxme57xUCJlcefJ1KXzOUAx
tIuE80yYfnAE5qekV6uhsCKWsc2JHxz9GZeh0iEj8KjN0r+2kvhKiii7x2tzG9DQ
iTwtfsYqo8gul9e4PnnUnzpZvXH1z/F6Ee1cq4EOB+MlrC96r3Czli/uCZJmo1pG
7CM4JOPZmmj0c/7tBBugL4rK3y73wGu9An7js4I1d/+8g+LmOASDU6lnN5T6OV6G
Ru/zqCxcY78tjCoQpQBXOnTdoiGiIB/+mDlkCEk71C7V6HTxJHdtORIq42fuqE8J
zpvsIHfzJr+YQPKTyUo/4IFWSVKlxXAGcmRa29BJgXTs1NfW5CYadi92PN4bpSDT
L/XuqAXK7g05hc3imLd8KA2Z9xqRvmayUSNZxyfMXYXAEwhhTZILBxq2BRaszaDN
3+QdwGicxaiZa5T5h2WefAYSXHWsiENOjjWcUBLFyIzTVU/p43TFujjJZLwfI0AA
q6FHwZeDcYSfI/0Ktrf7rngeLk7rndW671QsiNFOYd0icyKnrrA30IJ5e/aa9FsD
wfaRrnnOQYiTPUuSpZjOq8qo5BOtoQr6rl0Chx/gik2TmM5+69pviBZ5AewybUxJ
cSsYV6a9V4PWDQ4pr1b2Kg8t+Nz6bPYEK4kon/gRXAOdbQ8zzTPJHCsYvUGe3vXQ
/n7r63pRtNLm9+FFm1bL2/5/76KqA+qdR8CAsfQaSZQmEPaShDdgOwHkuxhywc2A
csSqVjtQZz3AdW04VlSmLb+yFP3z3/hsuikLq5kF3OaqYwbJeoFOv1KVbX3bjPP4
mwofdL/Dx7zKm69YqnexYOXbcsYEIUdFRTRZrIVUSuxPmvO8TFOYiZjhE8xu/J2L
kzxMRYAT/jg6r/uSrn0YvcQ3gVI9V9B2avsurea+e0jWoqqe1fbOer0XavS6u9U0
oI60/eGRNRE0jYOfqGZfC8JAgzJOT4zox/Fh51IVUE7e89vLOVROpzcm1G9fQ58O
dZJH7S29qQPVOI0IqLv1eOJhH+8Ac86dl26XySQhoJM8R3OBd968+s/RhZeBFma8
3NdwSbUqMXV697GnPiXYjZWBoL8d0EdBn+D+W1PpdUC2VD/xh2KJp3N5MPasjFLg
/uvOKWAD6Pj/kEZTZd9j+WAhgXHpAjbTbCDD7wGyE1DfZ/jWn7DAPrKCHuCghqkp
38Kc/cZ938QeNoB0brif9ecql6w3uK/Wy4bBFi8IuH1Fm03c2w7tyu7IXsWBFV91
cIFhmZRMdoxEhNurfdfKCawFGm883PUR5zbXwso//8v6CLRsZzq/80dH+aNBEuZF
CCKWJSawuUEkh5+300X3MwicFLhMBpE+VJeVtoXPqLEAQqnBP529fWFynWvF8xf6
ryLUMYzjJXnJRc50HDLe9sBVUHONGDuXJ9cJ2UCYlsRLVQUnGP2nv+XujOkzTaJu
2fwF+0js1zoamDyHyibhD1yTBRgB3LLaTb8Kbvxj9iUcAp9SFEIOvkFK2btbu/Mg
xNvZRewEGsF33F/Jbfztxx/KSrsNWwiGmQqfpJqGnJGP1hbXiFe/cRh5q80I4j90
xWbqnnpHJd2cLeUM/XTuwkQvBr2WSqnCBxUtTzeQZOscvPQfRV6Bd60oJaqyK/mf
AQ59eF1CB9VKw+N56ZoKfl9yiTysEmrCJkcr/qnRJY5XFAvr4u4IGpvjFx+XImBp
J7gyYNVJUytQ6/WlqJFbrBn5ejUtbk0jZRsFFmfffnj7YXbThqVI8hsS3oi5gHQc
KVi/W6r4IiUJ0my29RJpY3iWoFcVlKq80n+WEYP/lQTQ3T4gcXvA/9apPoJM6cZq
fgUvDnvtw80M2eSWh2EqzlNFO71y9m1LSzENg5j/3gN0WKJfotiUioV2Ctqc5Ocb
0Q10y0Vngo0WakZIy58i/hle8WkBzgWeSBc2Ijzl0LXpZewB55Mcj70wXhnapVVw
1fCp++9pn7ID/rc0b5wHiFiAL4grNzrjKp707sqAkPnpGYFcXjzBCIsObS4ofajZ
NJA9SmRKGukwfkZ+XTIe4p4Rfv7PSCAacmHmyQSemxn0Kg+2oNnkGnQ+pNffNwsz
RCPhrQJRBt6Mta7HAhPZOsBx3xH3GC6rR8ZX9sUpjmD1Azwt5eARA6ngpoD1HIvZ
ywRY/7nmKw80imC9mnCIjMVsBCTVr6/Lu8BG63oJM1cTz9jNhvRYHDF89NwFH7XP
iX7BUZIxfsYjtP5Okq1Seq261HaqLlPn7W2TZjNiZQoxAIKCsKUaMOoScwf47zV1
o3Md28DOEjQC/yCsTrj6x976I14pO5ropdtJZ+9aVgHZW4c9T14ARMuekfbQ8i/I
B3uV8esHSdelZtB4jxUGmWSyx19Jz9ZF+dBOGwMs+Fk90/U8vuS5x1WCMCHGoywd
3CFuS+OGZcwCrojMYFvbBrBDGvZVuU6nC7/B1RdYDMNgfOWQzFtGt+wwP6oSC7oK
rQLibsIvqWl+j7hYRXvuUQAqptshIdZYIso1gjEwDRZ4f6rKkas7WZR3sDAKkpL1
/uKiBpgNZXn3F9B4vBkAuWskhyeMfSxqWHRsVpTBsnsoJycRG4DOvTG11ow2TLiE
E4TjlIBpte133R184XC4AlvoYaQ3iEFfuUz7YeWB5xUTPlzRRZdzD9tfXsPRHASw
ZA0hYSJ4t0QoKsv4Z0Hcpa3nqJ6ArQhHze330XXrRmUIP6vcAMUY2fb27Qmo48mz
cemvGfFYUDswMysWht+SP+/eseoSPFEyZwOG+ZpQpOwKLDnbfIMBL/r5gK9FAOhS
N8gZU/2URdQh7/plp4YWJgtsSF9Hjv1Q78p56OLolQuTk0RQ7ggZcCv2PlbojpAj
EG+vsH9vQ9wQloD/ZobaCrdQcjdTFeVtfHzF9vPuGcc4Q09qBjDMWYBk4QGQrSpZ
jJb4z9b96M4w8IyPOtweokICSsbeMXqC+YKybrk6SE4PUpX+oMlbDXn1eQFHZsAd
nPa//Z6uVUNORP3GCKcM2s6sdJUMlpWpixCHLiFcZD4ayN+lDbvMzvqQBOMb0+hD
8s1wOEakdjPYeZV/hGYgDVBFGZQ4ztUAUlLYiQhAQtYVFkef6omsW1IaWiz++6Pd
Zl0UUehAiPN9bYd6q+uIG1QEhxYtFvMtziaKUuBYkkew6O7lUcxIrYEiDQWrMwxI
K+sjCssOqdObsxuYmESIWtQDQ3hnaLOAyloo8oYfE/Ko3WNpkz5/l8NtJr1ndnhl
CIKTG1cm+QfJpzSEaj1ossKeAHHYmtpAoNO9rV6sDP8eUQS8SciwWhc6kRLDjsyE
wUFfvC9aMnf4n5YUxi08RCnpbvgj/jpVJVKkbtBiyYOox8ll3suu9/9KGx6UnJke
x41dNW/L4nvZFvxkJ4K6LPtGdXbCFB8Q65WMBMxBdC67jkf7ouD0bc95gRCSA7DS
BMInXoI1nI9M/Mvgoj5gNPsdCu7S7sGlgQpQBlDF+lvan3rRdUT9kUEL8Bo5pccD
o0THOLtKPHiGJgeb84kMVMmsQUjTJ0Qs7pZhSRyvdfiQevb68T5AYLA+f4Qa0Bix
SB/m92EyvgOuzx8VbccUchpbmjQUmXWQOAae/+lMxOgk9B6KCtcfo5y7KxjOjul1
qyFkzs1QWw48U/nfDpg+Iu+x8NunYOq+IjEWo96A55M7SQie54ComBeRFi9AdHwP
8fwP+EkQ9Ir8YDBTCMx/Fi/1zIiMx97IA5aEGAdj6sGYC2VbOEeVxwOwL7doRMUM
Xp00p81xR7RktAE128kGcM0zmE6LrgkNzu/3Xvi+Sr9LBUquNeUh5Dro1Bml8SoP
p0GOfk0uAA8H17shv0T5bmfMESvtiwVBowZPXFTW08mXhI9pQzR936wRrhWF18dq
A/Fk8DBWH9YJLEtxW0Xzht/63cteNcTD2yZzvWB12qHbq1+2mFp3eqnLP4tL49T0
/Oc7kgZgUa6Q4rmw0QIu8DgtL65JXy6+p8tv6s75cuBQR39QIrvNFl5FixJ9W+94
8B2oEsghqR30rRazDdQ1JillpO+UCGJNOBt+w9lFo8LEHSHU8O7n5BpdvbdBigeH
RPpB/0yWqozTkIK2BglZOfMnCsR2DXXiQ89bmE2n9i7MsHOmc1zgl60awypjmqS/
gJw4Ky6EY3NjgSOWwgEofpAqlEV4NUFHt07cyWHmEMHduTKhg096mSOYC9O1yPed
8/Ab0p9PpZbewJM2jRBJTv/WD2MYEcBICS+g8oPGpdl4MctCVk2Ssl/IUJffWr+2
vFRaUFClddN5043m8Ot7gmYmTul3t6XdyXXdfL75u4rJXF/gJZIT03xnRJmvwqo5
GVa0qcWP1ES3cjCgtwdQK/EXyYHoLmeajCR1Jom7EzFEt40g71KvH6U9L5oIx5QC
5X61zvLyaKtoOoFej8MSp/N6tOF7dfe5kHWnPikpwQ8+RnGZrdpy0mdka5ngadGX
0Vty+T1P9a7p+SgdSMFKtU1yI9Z5R4BCTxwZNgg30R77HY5lZLahYf2UchnoUq2K
NpQkVdvg7sbnR+RiPnjk/3n50B24VHb0E2gYlckV3s9cTb/uztIYnkMDEKr1znH2
ahmRFmFrPyhMlC7K9+X5ahih2i0pxbHOz3lPtwC3wfeKxwL4zBqO1n8wv5bxraro
ZMd3LM5TUfSTZd0svYQhS6saF4pDzk2cgoj3L+fLh2llOX5sClBxZtNuD5a/Sji1
JkTPfQAr81tbxo5ZKdlRLiR8JPQc+pfFe3sblUcOlKo5cxytWoXCZhUQ4QJ6ywPv
1fJX3zX3wubgI9oFwAIvxXFr5gJkuIgMFrkpIHd32nAOFSb0dLUN/Ok5OaBVrKF1
XZmTkMKWz5H1bVr23psgH/+USaLu5wfHEC817EGEl1yquEIE7FJGQbq6TERUZTmt
jDd2dBDjougLk7IbWCs6Ekvgl4J6FpXHFnhi1mtF9dmISrvMGIgN5IbkR4tDfWsY
nDYx54Ro6NTYS4QkYD7ecGFpJYvk8YTFHTIbhyAhQESO08EmXhBxUUjAS590gLFq
EcCmHMQZR1A3L/haMmb85Nc+Ql7qkowXKeGRUfaf8KwFqpAXt+gsp5rpjiLZ/dD5
GPb0qAXaRsN/Cf/neZt888rIPLvceA7orNPcWM7B+y8VHuUR+O/ZcAVrXUcMU8Uw
ltRHgKAIs8uNCUm6g9NiNAgSI0X6aTILAJ5X4tbK1rvPGwdWLGKZD3aP6BwkOYMF
vLYF8nCEl2UWgqKyEIZCdTYWcsIDfvQLTGSDJ+CIZRtLmNWLzCTlZLkMO0saUSV8
UQBM14jsvCFibk+LiiqCi36QpIIr7YGzT0XCjqpphJgVVa/z47UEIODziow7RKLA
x1Evon/X9UtYd0PjIqDgMhCwbg4q6jNfCqGNt4waDcHOdwyLJHqxI+d8DLf/IOyM
bB/xqyyPKF19noviI0dBA13dvNy8Gdpdr+G9gvZmxoKZ95AbFZFAFILwfTx+uhnh
Xl/EBcIPH0imGhP4E2OwSLc5/DLtIvFXhGGK2zVKKlMmP6ujBDjgUxrHMxE2/tPw
iGLMAarGaRi9lksPZ3tCGvHXFJRoo6NY4cnf3038GFw1NjpbpYL3Ee9GrHbeM8ra
VH+h4YaU+8cYkw09PHglDuGVpXgI5ALn3eDbEkWGknCNkgi/r0DxKFzoeun4S21r
M6EPZ+thGKZr0n0S6RawT9kJ4BQiG+ZBD2Zs+iQVxhlsuBg1sfJLuFDH7OzYO+pc
kF8GImOkefBDsKRmnZUqnyo48DVZLgZHPN3POO+4VVxvzS5+CH+Y7tsmjlk0OtWD
FykiQR+zWQ3pdRbZk11f9S/s6ZV9OsGedpilxRBOsPaQ03K4B28yS4sz+K3TvnyF
Oq+6YdwbSxCdTOxjLtLeQh+bjdiU4MYZGNfkD/psJNw83a9f+I3X3Ze/NxKgV1rT
4SwGrq+I3bBYIhwqz5Mr0JWS0U0/BGZ/Z9toVH+qxr349ptM/VQqwAZ+5jwl45kV
y5Yt2S9EfQ6mp9s/QwuW2mYnMeibrSPWb3OiVKrM2/WGKpckhfaJ4mcHN8Giye4C
KtmLWFEEYalljMcKVuE5Dz9UEaQDi5MffE8icng7+b5INaIyaUzkcOPuRzY8p2cg
0hhJSRi+AsPQ2bPm9ZZfwIZyngsrjAZnVMkT97fCxNeFA2xHu0aHqdX7+j25RVkc
3Pvdw3EkC0UNZL9LC08Z8WcT10M2XcTCqPOwMmnLlF2PYRQcTOVWhZNHDUQq0bNU
DL25bwt02bPLuWQ8sOCnFUAEHnm57X3lwdJrxETplboOf5HcxTrDk+NIL88zVKbu
fOgi9SUOzEsYr8tgaMJKxZBxFLsiWQ5sGFdUWyq449vTgeswJuuUXHVNh+FltOxX
/1K//Mvh1jMGTDCLazCg/00Dzt2WCMCBEgxt/Z+fMgc0l8OSIiH67DqN3wA6ge/j
DeGYHt6aLRfQz64HllFGb6gxhjprtPYUDrjNTcWcEP2hL/YfWjn4kWilIOxJG6eD
lwvIClclUjd5YqP6fmXFanVKI5nXuOpCoZvnRBxYHSqMoP6t+hyVdNUVKwSjhG9j
XFHb+QNNAX9+wfyQD4oXSt8IQTYphnhFRrW4IHeRsuUt5jSBz1GiNrMidyop6wok
blUtKDwSlP+aJsmvBQajoBvqQmlIY0fKDMvArhNDqQJ2TvHDuxfxygUWQyVB5Tje
YF1ZpD8o7r4K3OVadZVjvWu9fSy0wmFm1X+QVo7AlPimgSP7hf+biaBjQYmWBsFw
zeh/a7/vUxW/vRnLwRmONjr6zC9tHU0mPzyVSIzdYiONoomM7m7bpqQ6kOKUKjOS
WaBRHWCRcGyW3dqLtqGWaw+vXl3kFv64A3ba6uYZCq2k5iiwmCcNarI+G2HqyTqJ
XbODfjZg9vJguL0KK7H/nqS1fnJ0/xopxAKl6EkYrp1UNI7iwm4jCPLXrHSmfnsJ
CylHCi5vvqIxCKedGf1GIf6mTRiyUSeAAkJf7J5SJ3G2VMsnTJaVO+OZtScu+q+n
QFbkKD4eD/AbWSRLZA4Ent+TOrQqleRsJMnmz816cQJsdyX85W0AMCUXvkejh43y
My+9rFhgfw/cF3Yw8FMmoUTjOiGiFEmpqW9EqCa5c1p4ZZHtal5KAFgHgPNzT9jZ
b6lCyzCGqO32La9yEUYAYCt4jev/bFf6ewfgaQuaLDcHws7m8+9xDH+QMMCVuVi8
mBFg5pLXGRXhsAoaKZRO2EL2KA33McmS9HuVWYnyJhSyAXoVmM3JdOM3HuRCYByL
Fz0jA/BLwSy4GOdxEBhP0I3ZJszkjmxfjZgRqFohyfqy2UvoUqXczrnFwBl27vVj
o55pW3sCbhGj4OmzImhrXKexz5hmNZmq1ToHN8sBgAdIxYggf82iwxyl/mnfa7Cb
+1f+AIauR9gs+fg4/mEBFmPLX2Tj4AysUxA7MaDTWT25aDibdOhDsuaJWfTcuKFh
01ldxF6T69gBKW10pSMOGyOyMKJvbDinMyuGp43Ob7Ivuu7nJUllcbCZpJ2E7l8T
JLKmgpdjSfgFEUVJjdoptMOeV6mYzH7CietJCJjAkoPfIKMgQIUOHSxtG4yn7Om9
2E+hvhO5C6Y5hdg2FoND+ZOi20+7muIgSqlSZu8uAEowIkMWFPez3nJT/r7xK54G
RTFWo1pzT672D7J4BS1V+GgXKG7m5AcSP+xL2lsuVyndOv49oeOZcdyGgDqIUxVH
Z4Le7NI0oR5+eJKll8Ak2lCw1gcl+o8PNeYx28fNxeQdFMacbp2bpXYyorVX2Iuy
9VIaplwlcfAKFELqocSlVOTY34aG7ozIoOmXVTSjTG4Jy9yiiF9dWTOm8GSu6w6h
Cay3LsvDk//SZlUlNgcsShCGVAKfU9lWtLsfqNifB94+ytoo7vfaKPHmjbqsBB38
Ewkfa1QMwNWfsMdyA3AOZbqs2OCrj9+TUcLX8g9L4+lbOsEkKb4j26h0QO04ZZEp
oJV/V+LxjqK+QfsabxAB25wlAdwTmdaazjMCIpVtnOPwDRpQWlLuE2PNshvL5Ak4
MJ6J/9w+ljZ/Or1ApcxAUFpZ/bcQ7XSqU6AfXDjhzPYhqRSx/aW/6AgMwyEe0pKS
sveihFKErKCAq0KN+4oV+Un6VHoOjs4C2rarybMWe4iPFgv7HGPZGPI1tasv8mXE
4syRlyzlF+t3rG4uM2zkOYZO4fy/TXheixHklX5QhBTer5aR/lY83ZSxlFzya/nu
QJ7hquzY8STmnti2BwmPON63hxGS4hMoYJdr1XWn5oDKG2IGNLjb4yiyERO/SYeh
7tvvdMT6Ov4TiN1tGOqBJ6A2vBIuL75jfU/6aUAEggwKVAERqH7GMM2/r6qh+1RL
G6ljIF2vvg/gxV3uKUDOI2JT7rAGpbZpLMDS3xiaXzrh5QjOdhf9osqJJRF+fdo6
1hZpX8Y3RW5ZOb5OGg9w1cYo+ZnLOMXlGTob6jO1gI0tsreGE7JxqlBPxMPpZdUR
96sGxwIov51foevHue4rBg+3o2058huu6QVojrDV3rIJV3MPJUSM4J8rzsf/4kz5
pFiVQ7jtBir/hbvgkhNLvRRHh+72FHl5qi3h4wbbtn4o6e4gVkC57uC4hHwGGbLu
FTlSRGwWQEtuWf8tuy/xB5vMzAYNrLV+xlt1xckfT2Ap7BzCMzaES16zGVuY/qlh
0WsFEe0ixxziGDOFkLOhtC/XglAnkxFbxwwZhX9f3Vlj5sDcp0vo4x7VmAHOUfpV
xBRgg5KDmWe44ZzdXjLCGsPnTcl6agcvB4EEiQ9Y9KHDiJOoqUqUWBNVexsjNa2c
g/uTL9DmmVlHz44pvrZOsPe7d9nolbdCbGJsaGR/nQDybdbIJD75gI63pX7PmWg+
FVRsGmiKw0+5+BD+l7N9owsuJsKnQEXprhleqCFuwHdTD4OKfTcLRps0F4Ap6K+8
6DQzeP17ODLKh/Yr17Xz84Q60pukIG1uKnYQk6aWyuDYMnV/SVGRV0vKH7CMqXsi
sGKSowrNiUei8x7kzX2YQfzSVa0OSh07pqDameBqkeYWDDsvdVk26P+ttySVcqSp
cLOOyWy+A+HNXrFt3AWxRQSxDbCamWwslEqr7QX0rxPfJENiltLY3hLof1s6djjG
OigmVxyRzg7ppnkfnb8Np+KU/5oiSzim2gIwMfRmAIgmCXzUXItfdrKEV4QoAbOE
iqNVyGkyEWiOZfDykTb93z4vuv2i34wF89RCRZfLTqJtYms21jZJsPWFl28yeGOW
DqNWMU0qhou+hY1F1DpzVCxXjPKuTbXXjPMwbpk4z78bYbBYJwUBoZjkFDkxUtsv
8zWpfrtwpCzaJAOPoPnXOh9STh5i+2wwVF+kdpBde7ci0VDxLPxeDGfEeXi8WdtJ
Fgeh9cFfrnHocW4O4NakFowO3eltuf2r2vC2/RD7ZRww+EmyQoJk+V+z8TPHCbks
7S4q+bR5fpmYt2H6/Nm2tqjdiIBqSzQ6PuGRNVkEIrteJthjzzPlINc+4pFMnLE4
7Mr3ke40IsVriglJkpg0X7Ae2fxwA0QDTsNv5T8/+JgC+rn+A44SGhq6oq3xGdxo
eyLfVGLa35G1gjDct/JimliiANG7EcT3RwZpcjPEfqbw3uE/LGI6e7hKC2nkNWPu
beRRNHy260Mt7Zn+S6eNa7dLiTYjbnvAMdBiJtXdPGnwzA8tk7bwuvnpTu/vK7j8
MtcAtM2keSVirBg7DDE6PKuBa0iiK/qzXZKIo0Nrm4OR+2Vrn16UigHDBni2NqlS
Fd0+va7cEbeoT6myEHTUkrLY3FUMnn35+GhQ55JCEERJ3YVkwfG1bZHfauJYkNzw
9X3/j2wZIVxeb+qSiYI7R2gOVKQbgNbSQonWTmVpSFhsb++/XsjbDc90gsrcPEOR
Qy2pprsOJzPIIQJ0Q8aP1kdt/Dg6dE9Ojddcy99oOJGf5X1QGcfrpy2cRLzNQJkL
P9iUDCfJ80bTCz9fe7XYuFFQ833Fo5P7XCHQPnB8uVKe6DNNZSx4BzyjKX/d998M
KqoXLd6FArOAxH0c36GcOh8hIs9L4PIZjhLCo0dOtmmwKYFiViKLq1+zsrHEWVDD
b0QrF8fonbhkxssKXX5/tmtvG1S8Tgy/WIxqmBrV9s/xTRIQiBScse9XPnD3aMuz
HmIbpug+7TTusbS3vJFi34DN4g78by2R/1X46yde1shbOKteRlqKlP4gqNB0MsBQ
w0crJgsO+W6s/yXoOOW+xqhPuvnt3UF3nBPr5gyZmPNaPsZjAQmL5dmSHDJOuRg/
AGFEkVoq0AgYtEwIG2CbKZ0u7kqnWWCHk/l9viBSBaEJJ8iNc3lK+gOTZj6rjvgd
NWSyo61ZNXoLgC+Db9eS2rXD7vu9+3hybx9vPyOUZ1MgobWDx7UgB+Rs/pw55Na7
Kmnigqda9ezmMOgAV+zW1Rjoaz6+LgXlOYKs8WsnR0fadAB+gEsPWdil4ppF9ytj
RFWKIEy42EV3oyZ1y/D35qYB/Ko8Xy/BW9gY+dEkZwW3yntcY5nOIdEz8c15TPFW
EQDsDhJnCEjVd+0tLOZxeRlKNzcpc7NxgXHASfKUj0OItDj7i04s+lwM1emuX92Q
yKFpmjbq/VUr6KRwrQi2laENbrc9vIyUp3nW3KnfC5a09DtDW1L77L56I82Ayps4
s+WVjeMXyQlvhAfpSV1lMyg3FkI/hsfYeVMJFUKCFaaUYO2EJ3OVwtY1UCpW2njT
xGmfWycMqXMDsSu8RC343mIxcUukNg8pSQKvtLlmt6uM95OrWyoskFncbnxrsv1L
9/47w8iv+8BTl/iTjp8J56NppydHZpKxods5JYsROhB0b7JQTES+HteALo7Mzws8
HXC14x4QtCFbLjmq1BZv2S2txhCvYaEVRKwaY0RRxHLtrZlgR46ppIG94jogda2x
ituCZWjPfQbpKLxBA/5d1U534B6W4Du+YrNPgNg1nV8VDyILtRinEQraa6t+rktW
nxi1xa7nmpQDIbNh1kvSEgDQaapqQUheX9fkM5byHESpr8Am++f4+m1IqwJRyNlu
VVYeIqOOAqac94lmidvOKSGSAO/H12nzDGjvUyJEj+j2plChbXV8vw2e6rSyEAFW
hRhcMMO/lxll9513mPZZAwX2RKfPLkn/U1w9Z8GWgRPKqufc3zLf5Y4RLRBrYr06
Jq704qVQMiR+Ztkxzwtpo5YzdoarjFKInBqKNoR115A87bHh41BRZDKmzsI+wv+m
IFzp9TofiNbVrOiheArLpuc6xjzukOx7TUr5L+nxJZKk4R8BuCA5dN4fzkMghiA4
yyHxydbykpSO2Nl4nGPwTG/VQzavX5PUMkPDdIwmIS77JzG/PAdnXuj9LKzFFrwG
PKNXZ/tg0eT0NEnAHvVWRMvgqfA9vjPjmej/6bK6J5EfMqDdzpJ2ALeHFq5k6U8n
Wn9i1hSrNF+0XJExGioLnMDu+bRk87TPDTQ+F5dBj+YlcLNWgbdqcCpLkgMpogIn
eL/R8HthgoMG2LNcMDyCRi5ctJ7qSod/w1AzNqgmJi1DQYMnMHueFnfFWFtdntLF
Nbvzo4SqaP/czat+6doUsI96Yniw+gWJLqRIYFKku5DxeRPU1CoSAqsUadk64Du4
WpKC64c5V+sCdMn90SnHRRYicvoXg7nZumtZmMmFx0fyYTkUuIgOM69Y2ZL/3gJY
0iTOKEWK6QyzrqzB7/m0v68ntorQbEa7xTweEGJSj0+jgEkqLV/jqLwOaYptaoPa
ilNY7WjB9g5Cwg4zx9YnlwG+Mny1dzsCkV7JbDFUgfbLqz6UWmOCJP/mC0J7XVrH
aZMuyfH5Bn3HJ9Oaavq9tlkchiO6URB7gBoTncYr+PERAb6O2ihHXf3dvjO8UF8u
UPAbyJLpAEhtQVr5CQBa8vwnO9O55wM73zS9/KYmw72o32k7cnFe67FmcYDzQX4N
w8KwMDSPTb409Mv+XNRJQHz4fjkPa0fLkI+1GnVYKM69W4zoDwNSb7Hg7KzKROZd
MnbGLf875Ya0MBDZ+Bz8ArO/WR7TLeQuDDAw7p6itaixXxxwoAeszYthzKbi7jha
Ak81oc7Eo+eOAqCvUpDRIc95skFzzHbNZ1KtT6c19aLTqt2FApddSkRhMLGTAPj1
60jeWm0StGuggqSf0TlT/DCEv7qpdQGqMhgov92Oll0rwOmUcaoO3jRLpyRDOqmm
WhUyrXP73mXD7EfKsEuYTgENiAwFQvnSzYdS9ivkOuE6FAqCgr87H+C1MCb9uXEf
j5zXzGDrYQAQKVdGztg5qpiueT+Tj4J4eI5TgPHYyLwWNIqbcZKhP5zL+7+dWuc+
JU1GeRAQdazjR4IdGTHBP0THYgY+Yf7Ooame+iPsCz2lifsJFL3GkoNsTQ9ZInGl
C/cjQohJ3S743kWJWHgwfBP96wCZkgnbSgun6Xt+eVESNzIcu6+zZDiLnZNGF7sK
apymjiQMa7IzB6e2zad9aE5W4qC5X82yVQSLiT15Ll778TyGGMs5wwF6FAmXZffs
9ubvkqxt05mpMZZj1aHpwWsMY0rfOFakRY806sOixWXM67e+er0x03zhGBu6NNmU
uuMWLsMpanncyX0KhlYUCIR10kEQSnmxs/ROuwsq/wbJcdNyDbK8bBpDgIdCz/uN
dSUgyow7n9EBNuGdL/Zlxdv/JZR3vRYkD1FE4GYpSs+emAYvJJe0QE9RtRiXsDrz
DgyfoneYozDuFTADfbCjFZ+v+HgOr/eH4AWBNU0wNE52wFpR9jFoKG7cIjKn9rjq
35Z3Im5CdIQwXzj6A2uCexBbuQcj2lkU5vLARvtm9gtmimCxjNg1WEiYATi0YHNO
LgkbFvNH4z9nWWoXoUHqqvsJ+GRinwbY+8FsgOTFc9IKVTyXUJVEA5EHX/lSQnhe
H0Toc/AH3U90bOxn9o3uefES0Pzs0G7oQF8+FAdCR34gnvjtpAdpoi5YCfnHDp7h
6UvaWzoUa6gK38RWs0Dzpcmn5379bdOD7yf+pUpLUcBqKNXDDGyYPn7tG7giG+OE
92zReYcDC+VTbFPPwyt/fJ34xZCb2DWMyVJoMxdC5bxikB/CTozOv+RAaLmwUTOi
+MAoU2TtAm7fVe0rnTAcukoA1E4Fj10BczS4dzGe2ZjPBJsbIR3VuTYz+IoJdsDB
c4/6xJvNQ/zOapx39e3v/4h9b9ZUic9fjoXTrlfIFKBKKrlcfkqFulXy30CeuTAo
d4RoTT74MdxuKefXxulB/G1I3v3KvQXnstAQAcIadw9+W8JT4LUvNQ6ObnXDtmWR
wEF4fSgpn/0ws+TGQUdHAU3YONDzeY1SfdQ/x+7r/Dxp4i8NAK30oTC+XwHUTY03
IwgkHu+xwpJVP537FrWW6+nKVRUYkuGUloTzB0zx9IKVLQxLcLa+6Bqew+jsaCDb
TvR3P9qy+/VvB7tujQ2YNnSAIkqDEuC0ckdy/B79jz39Chr8vAzd071WBo1EDBO1
asfZOddbQtKoji66aqNmi0i9v+5pjNouoYdp+RDK3tsHV2DasmanjmY+2GRjsNs1
bbpMYW9DycqqUbRu4iIS5LPL0mNUgIyG+7o1ZCgnlYtM379VoeivfBkPpXTKQP7N
XxsN0NT80KKrJwW+LZK2McOzIQG3wwGDmtXbUpLQIb0u7O6TNJXQydilbv/sv5h1
iWkXlGT820kn09CwU/RJKIa2grB8ZFvZlgzFMCD1vb9pl9/r25yvWuxpPiqS4TvJ
zFMTfWVQYnRsH+3fVkUFackst+GugIECwWti6id4IGkSp2yjOP/PIR1tZB+838iR
AUrz2qS1JYtBuTfnECD4gi8rHjZ41miuzZiTr6BYLuPrLczMEdkMaEaRKDqmMz56
CLtfwnMGlmQIAuwDwgPdIz2ctB6yQXjAFCmpDs4c3vkB9IOwRIKwNTQ7PzbOEbz+
e9MIhHRrvsG02H6DF4I9LiX4/zGyOFIh+V6AsYn5n2LdqMn1P6JhFldQtVhxKqdY
v4fNNh17ynmGe38Qz7OPGt9vLjMDUYmPbcVj0FPsE6pzWLcIbW5m8iiZ9ouv4K6E
zf7WzmIwfE+iFYSAgEPCrRvxADRAnVVi+vEC0gMDfyIGcrXomOm2aAe4DzVgGfBx
qay2lmynWEXkHqSgi5/H8xBXo73hSj6M1dX5cibVmWA3ZqQlwWED/iZUrjIQoQbP
d55JYpwrqEl18E0b0rfCp79cO1luk4CcjcoKHIiBMNtsN1p6T2eIkq0/LE1OJDR+
V6/7BfM62moKPLNuQOG/pEOKlQX+x+FTqXqomo4ir4sCTpDkklmd55vU4M9I3AxC
yAbX2Kc2xn2ibVZYn1UvjL4/yP9z23hiMzaNx0MpiqV8d/NyeSK5/n1CEVr8/6GD
AoanIDII8eF0oJVo19FNOsSP/ajDdJwE6qyVcUBDqD/OjRNpAMoxSCGli1DtZCnY
3rIjNZOlpuw/wHZRUT90+rNbyx1X/L5EjFBje0bNrUU+JMZpWbJNr0VVKQg4cfk7
tR2YoIvh0gRYbgPX3IGHBuI4cV7F89pqxT+HSaqcavMBOazFRI7HXcorqH0zkgJi
SIcYmwbIphCZaO48mTpxZWiBjUOyxQWZ6AmfJIORj9RrjdpX1YY1qAZQu1mlUbyO
fGGl/KjdrN6O5826N4zbcNax9vZWJqwM7keNuIJruCs4zSjB7O7ixc+cMNLCxjwt
YzQBL5NvyQOVhxC4LTBzO863+Ud/kiQTTVW1te4Paww7NayqTu2VYcL9hKm3dz4E
VVGrcZhhB64vDNO3Iwq65pYUN1ptwk3P8RP3fCE0xMB0jlyHK24ocndLWnEc45z4
znLtECmSGt2YSPdDQ/HM8BdUaIB1l2NvkNhwCsdscyYv6jcZ0hvfIeleimzJeGt4
15AGxEjY6W7h8LCu7gLPIrhr3iD9LHqrLOD5Mpgk8ZLmAJPxGT+Q/h1hhB7Ibalm
ox7LYWHUXzZNVXg+XFYP9LChf9ouIJ/rYUX2NtahzAhNZVs+7kk099RrN5Aki1Yx
frYAxorkmpTHv8WGPkifrWlN9DN+C3wZLZUjvl0xNLyzX411HT7JRyN0ik4Qp/Hy
0jqCa44O7HHAjag4bJGefvjFOjdjfamaDxJ2mor5iGniCGoW02eT56WiS3E3Y1OD
+o23a/XBbFfLf/AavftQxZuIC3iGP6TpHMlrgfSNfosr2Ukr+BiO2JF2eoR6N/30
auI5IMnGvw1od2ILzL6kmNQXHF7yvrzQ2u4K8zjZSvmBT2khNSLrJ3c6b16+a/Fj
8QlZEpFwMGL3n6UfgQUwn3f8SsTjJ0rJX3HEdbEyNCx5pva+xRD14i0mJdDTUZVw
rGuQ4JjrnI1bp9e9sDL3NFDwaqOFMMlgik5/ohbkJzirhw0mzeprDh1/BmRQ5PkV
e3j0sOfQw5+wOQYWC/CT+ALFiXxDSpv5cYaSLOZoq6T3DnMQxhsle0NfDoQdDyEn
K7LZVN/r7qLrbR/TgqdWY4T5BA8/Enuo4CYrCCyfpXPrxHfQpFX3KNbbOC0ZB7kO
o97l64XZ8xd0U3wrwbE6a8ohKmjUYJTLyMaUmPbXOuLdRl3q3uHog+TUivtRUh9R
YOp/cO2StipGvaDDvzkI/rxN7rz2nprjVcdL57h7lYPbx07ZVEisp7R1C2DAG4Q+
purNHZQRrVxqSbUrB/LO2OcH3EKQNhAd3lZ581j/gSkiuVVG1yHQdryl4qm75eCO
eIuS3sXnnarzS+A68Kh2d/ot+FmUl97T73miEnnQPq3q2ilKjH2+2ChebVYK9Clt
/MqQjw7wnIGxaGZVAwM72ef4wax+XXOsfF8LwdKCYGvI95wqZJKATG/Cg4yLsYgf
w26QPby46EI9yA2YeCLQLQqWQeSEy7IzSuL9mNquel0Ln+T/R8RfRBPw4/S7H6qj
sYJ+2ciE3r5eSHcvfRiDS8kZHIG34rLTRHbBCwxND63HeJsa1BVaVyVDzg31x/iW
OeSCXMhUNnU1RoGXRMGGx5Xje0iYzhJcenrJZhZUeI75FwNm1rzDeBCya26cC8uA
kJcz7NX1qJTwSTkwdOsH+FidKQqJWxmJOXMmD2zq0mvQ462uUtG9+YGTk5HBGQoE
peEEs+mQtQUHgn7g0DovhEQa5gx422vK9KyoB1eTuqoSXdSczsPmvzNQGSFdYsWK
pt1Lq4Xsl4LGr2QudGtWrVx+Px3EMZWnG/Ig8CmtzZFeeFcEKnpl9/4wCac+BmBA
SXvA6Kb5PQ19EBIgVLaYmMMBp7C+w36tS/5A+dqNUrzvPoU3ph+wiQrPRV30OuK5
LMqLes1k1BJJHrd4hAOuaTZXUovyVy5RIhbFbUOlTrrQSIhvSw4MRfxCy+5BNs3s
qsQTLlUaZUU6x7VUUWt9r9SkQF+bAIFQc4/4c4H96FMZ6E1v9E4jWA1e8f6gg7J7
Y9hLcUC9auMOOp6csoPM+ffTDVqRBDLHBFm30EuR43AxWcigazKTOjM3mTaOWmfl
Oi7UyQlhq3aDacErRctLYx/FK0StAIkt6G6JESlSTiJeAg3HNaPxnUcEOaTM0eV1
gybqq4myLEE2NLIYhYM/5lhISQNnXRw2hCiCx52YbH6byKYMKFj8mQMzdsJyNqcF
YiK554PDfudMiDmXEH0eJRqeRbblMmRPBX9zTbgHEvVbzs46gnTWQuTidNJfc3Z0
0mi/W/T7PhUDlIAyUfA1WLoFTzdmU44K4zm63mXU0/rtvS3ZscQNilxuJ7IsdzUK
Aw4lEpzoyZlYvdHeIhjOigFPv1gDFnHbx1jHHtgazbjsSkI+SkaQF0LaHuO2sTCc
ckHgZrNRKt8p8moGAnmlHNj7GsmWJNSPCsVH1VJkLypiCxHigGKmsEREfKnxoJbN
kxLuMdn/6K0AaWWHV/1rJNSmDFJSJn55S41vuFdR03znb3TBHastiGLGSLBhOJo+
BxnGvqr46y3iFgdggWBXL0EOYq3R1w2MEuqIHCtVqd8k+kgLybfMe4sX2PgHpzXk
6q5o3aTMm7KMF9qUrrJyDcm5dK+RQrILikaD0Sp909cppA7Q25iX8caBSytuzb4v
mHK0bPCJq47egchxSV+C2QtbKEF8HzZTKz1nuJyeUT3boJ6IIA2yDmgstmafylxl
P5EMUq7Ntq+7xnTI1wbvgHhnJzNMaj/IhyxJCCIRi3GGGCcagUWphKWEPaGTZYss
VIHSesTWEmSQbRJf2wzfei3kJjoBY+jH7Mm34NC+C9aQtdx+cKK+ErmC0OUstdB2
4FcCafWzvq0CVDpyAj8A0xkf+KsGdXSK7eeEeJedvm88oqkQ/4PUrENfmIFvSDIb
ssN1DTw7/8YxgIE5YpUXypCIQH3y57OoEdJbZXpe8gymHwiQ9ah8O2UX2Ad1hf7S
bHrZsWSjTxHfnyF55bmdOuLG0mbkL8jSqYmbBwHoypAXDsQbQC2zNy8QX6+rXQs0
BWbrMYk35vLiEFgW5EtwTQJ1YySeqIc2ev9K81im46mG6JyyCn3xEySe9RZbHDHt
ibmBpr8tcQEYbfCxDym8fRwAYvbrXZBLYBt7TXvp+PI3m44tD6/sJRMquFBOci+t
36X92D6B2uSscA70vZnbfkFoUByt0xRuAFKDF73mpHVXvcwBLoFEYsRB8h5GGlqV
Zz4tf8sqnsL3mWL40OFC3bdfrS8vrWx3B1zI7wh4qP7JkWdBV/by17lgTyjuL6LM
r6paTttIvgsO5vFtHvKi82nJThq3VPp3DfZlMkQdVSN7XB1asgN3e2xsKSdLM+E1
IwFUblg0axizgySybG+IqKWNGUxvlOYSwTNVqGS+URtXUXeUIAb3EOvOwokJjD5i
glHeRgsbqmuhrsmiuyNcJH52Off8OwH3CeeVxmpwUeAb+4M6G6E0h0R/Fc9R+WYv
DAEZjb2K27dORrGfuuDj6lP7lkhBUd9KXSsx+avEze4u04Q9UJ/fQgwt+xrm2rQ5
GK7ix404A+ujaPLoEG3Az1jfPfpb+Vr9JYugHXazAmJwphkfy07vdHPEs5+uO3cN
sT1zLCEQFl0r2mQol1I+Ar+ntr4+10ctUtRy7BrKXFB6JqZVWSWxh5RvmcRXPuQ+
8Rlsp35TgFe5iYPYbZdolszcmr9QKIrtfCqLa1muiBn24ViK1qtEtfpjz26bkjWf
WQF4nq6mjFRC+SXGx4/2z19iWOfQVh0DkUUqfKx29KSgvberLbEggoCcvGjK0Yub
nRXKOqPCz9DhjlSXh/MZj90836zbLBTk+zi7pIZ5UFLL04qjiySFCovHob4WyB8/
LSSJT2eyhEOJgyg2pQ8xSDd3x1VYtQGQ1BKNokrsmHc9BQJfQZNjysBa/H3Ww89h
3uL3zU9cCeUYhML9xRVtPP6gHbuFUGOKFJqm2MHyw2KsdPbPsvH/XI/U+7bxrj2E
V7K7jL8wWbiPYqXrt84Dm4JBul8UD6dfyfexi8OuvjJq7fO17ORowq9Rezwn856E
BlMUqMcwm5YrP7eI/qT+8Z8ePbBwZyh9bnGhBZEntPx/+TpJPITesIKYPjuZ0M0B
tIyhowE7SKEcl3QZvH7DW5YyznI6lOnvhdr+tQIonrtqNGv21nkVjk5ViTm3y/i6
+fn4P8bbZ0N/DT3PL8DTtCadp+aS/pyRxtz6j2uYPcTZganHaQEHnfpeBd+EutdR
+qQzzjOSkzaAwH/iJiMEmbTKSBYzE57vPHeRiiQTFwzGZAn20qQSgIL7a5aWb86p
9ggsxf+zyULHN32xG3IIv4tpwFNTNQDFvc/CKNuo+vxEDxpzOgf6rKA5sxDSP3yL
1oz6LbHqoUWPcTFkkjibzmA9YORoWFcPlyxhZdrQvNu4qqeIB0VV9wJhj2lVhMNS
BbZYFk6WPT+4pu6bukwAsHjEaVihYMKHD0UZ9/KTPrNazl06H2vWJo+QVNa/njM4
wY5nzgCvJeMu3HaZelbtuBNUNmGYuzH48B4DC3kLoFNe0G1Wdj1Q7gCbRZsA896Q
jBRqpnuKW/2MZhWBR2fPAw0zd426KHlBL+uspZ8KGoALFDMX4sqb2v9KFyhJDzGh
ldgTDxaYa4lp/w91RhBe8TolMDk3/ukN/M1GreDyCkYB6Q0/iMrgEVmWnmrBQwjU
E16b5tysefrzDAcEPUFhh18GUp6484D2rAuMdUWTUqckf6xatZXzd/xbpDamIiKC
JU+5Lgy2qFH8Kb+ex/2BTOGBUw1c5BkCERJtYvQ7a8CP0R7OWaIgg+y1QUla9dFi
pRITDDWGwnFMx3k87FVoha3IQt6eR80rFvnI0KH/D7f7A6JArqxCQYu39xBWtpca
+bsJtnel7QrhmqTRfJjJlQSOLehtIYDWv3C6FPwUH+rqWV2uF0JdfJ9BGrV8Jccs
D9uZAY5sO3DDa8XnxBSk2a7y2XGQst5LXUPAce71hjcDk3Y9GzpQVjmNH2cF3O30
IEcKGtSx08skYFWcEyHXDkneav+QqusOzhJSyGf6B9vyzV9qfYvWdWJ7eY/EHxe5
Nh8Zm/eujlIe3FAAaJSSOmA79arofOF2O7RQhALYWuG2WKwLrrIVICy5mUsed4jd
IMF01n3IL5nGWICrTUXZ4WqFsfVfrCTtqD0+RfV2V2ToogYYudydwMOFiWjhAZ2U
uaI42znNgi0YUJwsXZ1WmGxFpEB4Zbv+Y+uxkH1E+7ibutQ5UehlLraJaTqVYwuJ
nRQKd1toPcEcfye9jhUowsrCsD881WD7IWbvy7lNk8nDRHxb8mMIariULGReJmBN
Sq45FP1yuJrVelIG9YT4NUODLOoPLRcZspAm17dYm4Sg/kyIdh6NAv3tYmHlJd2Y
KVU1rUl2Bn+qpElpaRVVAl+zx+4DHG9GzkOZvXtpRPLOqQk52RFV8U6q+kUOuYOo
F+CnIRmlL4b49llbm3ehWwq2yQ+9pHoda0N2DPriJYUVhcXkC0m8hU1ne5XHBJWZ
2AGnEUysmVNvYx3CJLsDcYM5MuZtLogEUR7o4iBaCrRhkoAchC706EM7h+Ycj83f
aYHyOOW70dvbG/dx3h6YcEnQZUW76cQlpbEyfe7gJ+AjoHHBLL2FIevtpjEiIttr
IzABnzOGKqgEQ3EesU5hhIBQaD0/ILqy2SeDjrEI353n4hlyTMlrorYWXMoL3tj9
7gjfrz6EEo31SpJvolQ6JGmFIBKy6oIsGQPUuZyrecl8k8NPR5jfTk0radsN/5VN
mbKQ5xNSVTUrQLbv7OVoC1u7ALEn17F+PbWjLqe5WulQy3om3pVk61YUTC1dHgOf
wJWJ1FXOovqwbj9qidMj0439QhSKYrcdPv7tSnzupBry6+kqUqwkek7sdRjM0yN6
NnC9mNpEtl0W2b1JHfbiK/KIXfc6B4VEXDnmjwaUsTXSfNxK/IZG3CwXzLMIikWo
OOSyb7Tb/Ixx/AF1kxTqvmuEdr7y1qqse+zKVviyENEYByN5W5f5tED7LvPqE9xm
2hZWvTYRIRKkKynefJtOxWMdnIidjs7u4vpkcZqOHvdrc36H8FsHXk4m6+8ouRve
p58ZlURS+Pk6QfaLtgO3ukodLTSnHx3brgxkJo2KScnTZsMhTICUzJmkJaAVCRj9
iDzwt+sAx0WqpOuP/iFH5om2L2pb7usZExNtErrwE4YJ2WDszZRRuPaUFbEjb3H0
jcWqr2PjrGPQYLN7vekD3QKewkxIbLYFfqZd2itg7Yj3uDkLzkdkv5yc7lPOBbq+
3x20BAFN7TD29qmEgtBr9RXUI+m0uktEp4zptmTQxZFJOpcicWqDtSjbxQaxirgP
ddtanwQ0qJ1eOxDWJSFAP4pEyoPNayWhIOPig0PLKz57ilYfr+WNqICSkxk+7bFJ
rXeyPoKABZlo7nasswTVK1o8cuxizltbQ/7pOP6dpNFqV1O9TUhQzSKo1v+TaT8t
0+fL/Ze3S5Y9+nRLoVPSl662g8Es7FPyysSeyiyjk5wrw656qm3GYgsZUJAz+OeA
9/aNgfOoNZDUwg5kwZjTO0EP+Dv6P5sR3DnRKy7Bav/FOB9ii7aOWWLMIW+flLeB
RyiosXB4SQ86V0XwAEpNht27RH0e/60g/ZBboe8wGr9WxQ1irFUbmO1etR4GmuX+
WZy8WX6aUW6NIzMdqd5XLVXNCkIV0XxJzQavQubQ5S7aXJ5/c/6kRzY9+wAj+6Zq
6pv5w0B1mYXIBmZ+KuVWO9iv2hfy1ZXWl4lRPA8pql/HNm2oF9PjYvpmXO8x+UNL
qUOpah6sgpsry3YfaeCGm+JZp/hbrvPA2DHGZTb2RLCsvesudG144HNIICmeQjW7
vBhz/N83Hg6FTZcK6M9FYt/IoSCEqL3XoAjUd/IiVkpoYsbu9b/5bdSv15R3BxDA
M6bNFzkI5mb+7uWkjWtcHahE/n1Kc0F/t4BJV/qwvNGnjBFR+8ecCSHOKBb7yTHC
Ecvn15cJoUEQ5fFcmc9DY6vJi074kzd2IG7QjVhk8cPzT0x21O9VxqlXYlP/8Jiv
r/VKIR7TasrLx9kXeOcxLPckaIU80Zrvc8hlhZRQvjG1PZ78N01d7eQJ3CGSzcGt
kyB7EWMcuZDq8ILJIrYmKfPO4tHEAryFFavuexu8b4vnG/nSqNHMXLrY/0dKC+nH
LmzKQi3hW2Ezjh8A9W0MKxhNfnV4529n9G+xPICOlBWcSoWRA9ilsqMC1I3PgX/n
hB/Ca8Xi6fBn+3pFz4EI0Ngp1guggKEMgzzXIsmJXd0kpcpbYnhICqA5e5DhUccJ
tKGRERb33ttYwLZHSYSoCyTeVO4o0D2+4+1OrKtddfy7S+XMayVdFybEmSjMCkMZ
dahyDAQiLANveLeXkPbDL5DziPiIzDJdRDSTszWBymVXFjsEVJ9bh7YMhW+OcPB7
yxgmbHik/hXymKCqbfFtCqLVL7jpOcfcqdM/ng5F3man9QgXJsKLfjbYjig9SgTx
H2X3OTM3dV/AXtOzVR5zE2rqGNCdHuUUaCq10EFsQWy0UZDX8JlXPQM7LoZr7/88
J2rNONuvQLA+n9a1GwHYO1g4R3y72vrbbC0DWVSSyM1mCeew9czhkfM+ZzFcwV2s
991QSIgAEhCyTIFpluyH/qvB/DHKQ3gTCRh00bVKrAWEDRuxPspy8SeiO6GQZ3Sa
PzB8qUIMF00blQsuJDZ5jTxAm44rU8X+aIgyK4ykeOPnJvmkENAI+wUhM99NgxZW
wi3TTvMzEv6pvOytuYs45IjdUvH4GsQGwlQU1OFrRPjC2KpX26MQjl623FkZ2qNk
blV62/hMdiNGUz4ag577l56kWrTb5UroPAyrM6nq4PjcVBR5pCTHwmOhtHMQ3gan
+1HHF/4HD45vAO1UztugGFbPvRogXYwJhNjoFgzbiUrEZcUmf8BITPd5LDSEFLaT
rXyKfLsRAL0R296lEvhl6bhxratBAVbrNQPDSbblMHSlQEZIQqNDiKfP4InoKkTv
L87mNaFH9BtCWJcdKch3twM39cGC/LLQZ9xHZ3pt6ANQmI5gtb2Le3zj43p+VXWA
N8UccYWxndrGzCHYCLvqkitJaWAg+LgNrkGCeYUqKyQ5QYZImwIRjUBSBccgvGKU
bY65ZOXuKLOGoYFZ0vl8RpBPmoAfW5K4rzxutQCEwn13fY431dP96aSZy1/vSxxq
vILE7hpuzd3HW7RCcReE/e+3qRl50xP6gBpGUk8Ncom6ESiX5d0uTthZ5sZTygWR
R20vyRJoCs5eOJszG1GxKzJ50IdwLmwb4/oOiBWE/XtTZfcEIekGEJ8ZEB4BDFQV
f1kIPPpo1+NfZywaMjdcNCX1JFfHmCyU/2je72OPi/89TubUwSZBR8QmLPiUa/NC
P4vjeO0Y3Nr3A3nyu5C19M1BYIKWyjHfngg9R+ObwoRRD26tl08T3CWzOqYZU4Km
j0yE/IMOG6oodVFYNa9Ojbrhcj0NChjHLEsWJo5DAYRSGMOMkzfsp4Gn6dDILsGL
TYrRWxLaoOTNsSwVMobcvqEgwjxs52ShKTqJtuZW35+QXWn3LxiSFVBAGubfqJGL
7JFx3CXex0MMpUycTkGl3l6z5F57EGFNkMXJkzBKo2DMgSvvIJVXQw/bMVMY6Hnt
KrXlTBPW+gKSc6qRukMWsbfsr8GW99AHnXYWv3rMp2Yr0Bhp+Vl46FQl018kVYfV
bcYcm2YC6kZFza86f/CZoS35vlLGZ2MxMFKp68i4yhEMx6NDPs9LYTaq/Ouy351E
92b7v6liLIST5Bi0Awk5x/xQV2hx62sF/mYsdWpAVGQ/8ncZsdRGh0XAlHQzNkF8
oVrjWaDAwbkNf/eXFmdCHbU/yYTWr9gz59va0GdUbieGXMtfKX7YQsYzIVKdMQbG
/h25U422Ld+4GwFF82r0+Y7ipI8FaiF2NawNsIdUWF2sZkEOIkaeQo8Swp77OcpZ
S5DW6Xf1hKKvqOmpvv5xfKLiSCDvFPt+8KYduQwZ2EEnO4qAykHjgWqfOzR2MxZo
tGp7nAn5tBfFbIyNhNyAQ9rvZzjOah38qx7GyirWSbTV/Sq0nhJmXqA5YWNd6gnF
mzygKrAQPqxiCtT3FaWBGQiRVTKC8rnOiMerZ/UU3vRtOrLXFxL/tNJ7f4IKA32f
tVjZ9c6tX8pQrthM3ypt+oLoBnyMoirDmrWtmvqZEHK9V2NeANrOWfO2OWZkrfjM
VSLfTulOF9C+qIb5dPRrfyKle5lILZYcUN0bKDNaKVjaM5qlLkZO5lWQaosEqvnK
+N4y7QiouV8qU8JA1wLYb9n7lezTQW10SKvJ2lcmQ5yNbTgOCTmLHdlGVCVBPAxe
5ASvOuZ6btIFszBPLqA2+Oq4eFHqI2ucdvKuStJx4C1uolNnl8YQgk2yyMFdFMxp
S0yp9p5yPLlq2QhlQ0A6aQCLV551YkOobxMR/FeDRqgnbMzklTUFeEM2x1wI+ZIy
LmSTXSpgwWVhCqbeQ2a9HYACX7Ol3d1XhxuH8FtTm7l0tmyZDsdDMm9BuDcHCs6P
562YqCRFRzFvM7oz5mgMVM6ssBduSUthOlOATu7dWmVajGT8lmOsN9dTmtM8Jj5d
gV1XRB1M06gJD8P51Z0WZ2n2mnUxduHa4kDmsJOdHg/dc+sfefeyftDvWcfZF7Tc
dE/W3KiuulEG3S07jk+U5N7X3wZTTSC0ZFOmhs67WXcpEoVm6WW41gKR5kiMJFcX
6uPWiE/q9TJyFFVoYJSdWCNBF/ynvWwPR2cgHakGfDgLIYEqQ/XbSKKzHR/e6JMn
NRsX9+Mxc3gcd6IzHjccrkk1Cl+ovNSNiAe3cdP2c1Mec1ehNhKpTEnTgkfgv8Nf
Xa7RPNA6jF7Bact3kO2w2G3LFaUBgPZQvh057q8dEdtcpSGgJmTauEn0uBvny0Yi
AEMcJLJqIAnoCk82nEd6aR+WAWxcY851nYiVvcw0eQdg8JECA3teMgXnosYLBQnp
urS0IoYhuz+MftFBSlbdfW4fI7NVJEdinr2pBZDnTTYe1X+yUYYAhGyNfqRB4cgW
vT0ge8YTRYla0bMU4dyvfS+WNIAiYLMB1yMCIB4zXlXKiB1yBefw000ZRn6qvlwj
n+SagduE4g034HVxsYliWcmXeUX+5ic4asu8MG4Fr2uoNb4eyB74G26ZhFY0sNFN
ZqWuelgfDo0OUeUxB0HioKLo0StDe8YaSiySOhb85N3b7WP39zPz4BXNQnUeBoiq
aNSLJphOaVVviVFYWg9ZYwJOYAgDxh1fQh469TQwdMkrEAA3WS+WXg00R8VmBtEr
jVXauT+d4ywjv/SV34oua3cowY1vgFlnzFnAAhdFeIQN/R3P3FX4dX6oIrsTflru
XQ9sDMC8MDIQxbCGYc3kOpIHR5fmM5H6JEmCCynmGl9adQUENTNptEfgzbm8MrV6
8lpuXtZuhDGHkeqbsGBTY8F/4GBbUFdXN0ATA4hlKBbanI4OPw6vVqheb0mWyNDp
8pI7mWXl/Sl0GS1IRYEbimsLsPbOUXB/7OvROX6WHjBMEb1WvNrt66N1VKS4Qhfw
6BdXWPosHXH6iDNfkJSMbT4H44SUU38rAQcK1YzhfmjFj7VnqySSlfE8+J+dEbyb
CtDkxXX55r7nffjb+5y5rryZuIVTdIYzcngp3C2mZfASCIF03jp3n8S0GIc2zPRg
/+N3eUP1M/BYkxBsT0i6DBgDa2S7mGkwqIz8btIceZHntXCSe7qXoS7oJlo+utdH
bNbOQfVmcdKbPzAe7asHkPNQn50nX5bhgC2MeQbZ/kvohDj/0RLyGh2YTAJaOh92
lsO9F6cCsdJFkpxbvyJRjpeqyxtb0TlaRJ+4UAHVN6zawSGYmhmUNld5pge8owY3
s15qy2xBIEQViXn/vjJAddjrnlMHog+oRoeg9/TL6T8ubmdxBkR8dGYgPgHfUqXa
JhloDKIz3BCX7Y7an8JEYN9CN+EJ3XTleIrKSxDOS9GpKEF5RTgnXaM6YSSTJnFb
axgOmcF8aANqoDdHvgVa5CmQLFz4vVLPjxPGbHVS7aiKmxAh2Wm1MPscFQRH0pxx
rtwGjDui4Lmcz1UGOKS+egF+uf30ZvjxZvz3Mf7CMUDsgEVzRWPqis/f6gFDhrQr
KYU7l74bXr05odsqzyKxmB7R6fD7QhAMCV/XHvnIJD7UJnWd976nDqxE4Oh24LR7
UUfEcWIIUNZwUEQO5U3jQHYachPcnVuZw/lwxf+A0GYcqNjvAdxHfC47d8vYuqEV
4hfOS5PXbiYtREDDGzU6ty+7Q9mvA5q0pGxpB7uHiDQu0SKmOVqf6ye3GirdRyp0
6ktO4Un2tvj2/5YjbJSLZqwU46Zpkqp2YHsZV7EuqplTMXwEQXhNB3Md/KxI+Cu+
TCZw0ZvUnY0jrBewzcpQT6UMsu8pLFBstriRMqLlbhL2zW0n6hAIiB/bInyKLvdE
A0HqQRKtrccSYmAn+1zSTfy3xxtwxLFxTMhmHgo2of5pwWcZ58apIVKRCXDWkqtc
jKIF9MMOZ8GaAf8EeeoL/335z3kL2CXT1cp0JUHDDcJxxaQYBVlWMN9090K6yrSY
A+38XEdvfrq8Q5ai75qKW1E2hfirIr5kFM7HyYiFj2TC7RFjgHPPvBwby+IUglZa
Cx+tq2Md/w6Vx2p8xir3EQd+VOlCKfYY7QUQUKNI7DH3YpDu4KQRC73dI/meK2CO
cXyT5wwGZeT//koSdwdaeWk6RT9kUTWsaf84W/rsg5t+GfyOzYgvWF3LkzVT8DWS
yLc/gK2SHoJB37kQHEiMuU7qVpsH2mjGqGaOkw6arwNCVkvLHOEuuTvNzenjqPXx
SxT1cR/jrYOKGT6QF0H3DMVLYj2m3mauH+Z0XuQ8EGrEkdjWkfK3Yg3izC95dpaD
uETDoPedGmw47RUCgDEP6M/e59dM2Qw85HR1wo2cU2kLPqAuxuh7WgXr7lx/Q50R
g5LN6FTEK/sX6gg+PiUYtoiDUQkE/r/saPeZ+lXNXAA7Gz+HOd3LuvZqJ18qOwr8
gvvJ72ySrdYTmNCrCTN6iOvVOWUKbzUcd5X+6aohLrhXxu5Q3Gf1Cey/+3RYDzaK
+qrcqw55hun4eZw39yZSxTmQ9suFKWXIuZ+125jVKkCbcoEF32kbAU+NqSE9wJiH
77QOvjgChltKQTS4jNKBEFx2lNGMxBssiL+cXkxAyAwbDkQohhi+ZAB3AH27ilUN
MToXmhf9Uss7oXqYrdwcU3nPyATCtYEA8OUQScla9AwYW326bfjn3FVAWmG/+Wmo
KeteTcSPaJSnf7aIoNbmlquBTdkvnLiQitueay7zyAbOpyUyqOJ3Umq/etzVtXfr
FNtkJaxnHPYsWid7RJQyRPmpgh9vecdnGtPO6fi+cBneHakr0t8trZStDyj2NL9T
be+xJO/unP3F01EUr97uMuLddeu3icaS7pVUXtDAmf6Iepp62kWan0+ExrSXtLaa
eEPz8qKywJiw2M6yNwM2KKUDv20D93NAMBYtg2uqoJ9mS+bQZ9LBo7ZDciBNqlSq
Q2RNwxVkgWwJCB1uEL8h4TlHxvrgr8VNwkGsPyHYf+I5VjxRTJmeEpScZasZ3Ho1
9v+0/U+V6vFWR1w7JrloSyOlCZc2vtoBRUdvflMc2TXzbdrZ9Nbr8+AMgou6w3Sm
lZWUvbao4DcCxExrS+zq7Y0yosisDnt5DLvHOFK+Ois4nG0k1H5e0iqrDfeQD5EN
87fRMLg5iF7q2QLghaiVOXCw/ItbSSJvAkPGAjigieI7dOAaRVnuVze0ZVYFMTXy
zwNoUuBnO6L93SnVooDswURmd2KHChvLgbVKNYgyTfjCAhLkATQG9wNxW9k7ky/P
jEB8E4X/RGxFwEdYKULrUMgNn1NjNwSSny5Vcc6NQHnhngn8iSnzHxxJz2nWKXAV
E5XowGuew+4G6SMRLss7M3o7B7L/EJysE+vArNwITNJfS7DH946QybZR84er/fc6
3yXzGtJOwNBtzS2J6E1kDPtPM85iIPgp6bzxMyjlwbpiAGaA9BBZAwZP0kCXpZa6
2QRnlnQAgb6BY3qKzbNQ43Ww3opmp5CEmjsiWVxKZTWJ8vfIChlhmT0UzSfeB0jK
SZHvc+gYdN4QWqz4mMZKUb2lo+tBC9NJwgZdtKELiSNiqrXOcCOenuIWLVr1esdF
6m3866fwKmC7OdHy8BzkPhGFDvR8jJsxZrVo80wod1Bq9raUttq2nW3sVHX+LUkY
DI47aUOMoHnG0Jv9WoOXiIQlWYDTSA2Mt6+LMjfL4aiWjez4vnGpFcw+9O8lKMYg
Ri1QoeL6hm/jkY7mj+eHoQN9TgAfaS5cWuVBuUqxmkD2dBBv+XIfxopgRSgsAS7n
flucxDSsHCYN071VhUT6jmEHrXj/Y7FvSE6VUjH6StOYWta6ynxVqZDtu/O0xCvN
Qb1ooLQGTptKziTmthioafLAy8PGkq2w0DE7WIQHrjfPdeWMqmGF8vOppfZv6/3i
oceEiK49hVC9OL03oUaLzu/xwrLXFKHw7/KT3mFiqS23ttk6wf3jYabZ1GUGU8kH
u9QgR4orcgff1XFvmbNpX2/usq7nEE4WmBX1FAgzcReFeJcKfCX5BromYFhuIg0y
zEEVW/Pdc/tMGLPTuYFuni6Cv0GPo8Scsg/vFlDm2Qp5pFl/DFOfrHFleg4AL5Kr
QtpTam1SGB7WmxfY8f+UZPQa3cGjfaxlqv0jFrpBBPflVQ8pKBD52JiEgMwvld/5
qLz8B4cwsP23pMb6h/Wx/xgjHGNBJm1r2pSm1ffGhpCf+7PppKxKl9IS9xr1K2sN
MexB8pQjhauK3A2XzvBiP7gRjwUHIz4YL5jwxWL/W6M4PzqHS5u4bMT/2b9CKzrH
ApUXHOl9dE+yyplGYZdlpyxi5zk85cz0p+B0++UTY+pvbshhoYTzoDAVGnuiMlqO
dsqDxn2soUmdYo3krmp+Z77HaLn88pbQOBkJ34OpcPVebSqb/uLX6APLI0pLZFpv
4d/mgS7+u3HhCotQUc4jj7BEEuH5Nnd+NQisZ/1vya3QaZg35ddMs3558QIglrSd
+dv4P86SPkeU7oH9DMsMpaXY6MBEcI/rtJYPw1g2D8zP26aRgYH+w5cN7F/v9+PF
ahCPOduFRRLWxvzV+L30eS9XAYYgVHSHdFgSxdPLtTQfgrz8oQl8N+Fjx5RcrVwL
KFx8m6nrGX0Jzn4TkhwcLzu+rgRuO8hEbj2xI6VzoAVCHJI4k4IRLjrgRHi82PCL
7XWvmJFwcSVgk9ruD2Offf3w+qxkcFrN2G5qAang4gdPQuDEVPvvsPghyjwd9hbb
SuNUa2d0lBt0rltsMOUqsU+lVPE4bmDRqmzobTWuWM/kMAD2XlTnj/xvnLdd1ZP7
KtMzQ7dzmqaGotIF0umyOBUmkQwt4sQrNaa/YkAar//CmJoLDb+FFnbnzS0TmfNZ
HXUN1l17jRvzCOArJjX40sJdmbNW0q8VvImG3xD3y7iYXCDXrc1pCyBafAnmiOSj
3v0JaGJDN0Fp92hVnW/Y+GOPOCQYpjmd1ttSsgJlROrDAtVL2mLD/07SyqDC0iWS
BYu/C042FFnjKkE5Umbx8q4rSYg8kUfGQ+/eXTc5j0UyWheQFX1iR/gJT6SDDvYA
+BVRi+uFgg2Lsg+rxXPyWo6VY4j7tz6FvFOppDKc7RIComiO1FDO46SA7CTQ9OlN
2t7gmRBdzHWwmioWifdgYNfkMnkPUxSCO6480/NFa3PX8CtL+XYTCNr1hl2rTVX6
VNisq2Mr60pwhy+me3Nqql6iv/RSZbLZoCtN1M0gnMxzEmjDA5FXQGtbcHAC+rL1
njO8hKgPaAIZ1++jjgGK+BNvIjgAZhDx+sGtMmoTbrObTbS+ICgwJhdFArEsIWtI
CjM3l6vSocVgFlSshfo+QP38Qp9NyosPUfV2Ywihk/8eic9tr3GWqfk63aEiDE1f
FaPq17i4RnJuow2ql0nIXh5K06MM3TEt19Mjcfq88zlZdwtjkZ5olNBYTxHaQCT3
rM/A0uVIxLv3Ul9qs0S6s2n2qYLuxyT5n4ZoGp+hs2c7SU7g0hMKxRctLsqRPVyH
nPnJg3bsCkPrQ6+eLtFPiVYn0kPKfvLwsyY6klVYAdmgi2nHD9vME5JZJoXv7pJM
9Zp6qbPmkarYVmcJO6EQx73F0bje0ljnMupVawYIbI7uCuk3RLuhGj03ZEoRro23
T8sR3MGDFWGMfoYqRNvbUcyiix8VFQPysYm79WzMiymXRyxfGTXXXaCF8xYBvHfe
OEq90qHzKelI6yXiEhozWq21YxUz77d5rx5smg04+BgfDR0LyLCD9l0scM9GQ6Pd
jy2fJlIjxr4kTm0lcFaAFU/tUgd8ygm7cXHzIBka0Y/R1BxNAiokOLoQHj4zVSM6
skRrYxBJfLHIhJPWY0lEqmA7hJlEyJilD2xWGq8xzJc94+sq6SoYya8Z8HjAnurM
4oLeGscwUHg62meoy4avDoQFUAL7JQ0mjFYhc0C8FEpx2dredhWfnzKTgJx/INiH
B5xKLbKAcFgGqf7QYERZZeeYw8HJPWXeIKZ8u7iBQD2CPsaOUVrrZDVoq8SyRsmL
IlfYoZr2XS0us3Uwr9aJuvynetjggqYwwNMj2Ciya+C2i4vTundma0MAr9LA/UyG
i/HwTbxqis9pUyXhlbVPpJ2iXo95JNy9YoLVogKjYb0z7RzeRGayZGMsgcUaiBsA
sDtKd9qzL+cuByv5hxTZMnJMVR+MkUSadMC09u6Bn4idw31QFXVW9bH/vdIDou0r
YiGCqDf3yJJtDmi+Ifo9SgRgInPRJysWhd75wqQor8pLA6HwPUbv8uy8lvbM9haz
/+HnrWzwfOL9BtVp6picAkN0yIYWEwhgJqbIfE37hKJLY4o3qcKcRStpEFs1wlq2
hIUoXMQSlM46+rxjLHc2e4eBqneMW2BNwcF1RykHJJM8sjsZKJV/vw0f/0hb61G7
mDQYA1sj31pOdcH5HTCDn0wS7MyXSh4ehwvL2Wm0TYAAsJ5AmRrXFA+QXiL/nUwL
QwVDXdSFKQ8xyHCV7srMJyzep8caAeGEK77b5mo3Vl9vy8OSoRUmeOtok43utqw3
Jw2PjRXmo838oXysPF6fWkxfeKpzIhe8ps/ZrmGEHQGGVGy8qPavHL6rjyOj6gJI
ivUdgd8tietzyE6GuVWtV+JYxUB6bOlP18UYiL+5MZiYmNHfbfj6NcLbxZnnwBib
eK2938hbz83owS5M7z/CVyytUana3m28kvdLMsLavh9Zh17sh6VYlS3CQA6dvHsk
CHnWg6eOKReA1SNOzICZsIU4LnTdGoT4a9RHLcPZozUOczbrGCppK900KFXByl7W
Bg4qiaZ9OJqlyo9jGysrsmk442EMLVqaNm3Et6/1WTBTB+abf2qUBtD0U7JmCuQw
pIoZsMG085iz5obiuGWtEzb5REeCzIt1IuBVDCC6VOURfgvhWSzbKXQGfQveNGJ+
T93ICFrNqQfve6LvZ9eMLJu5QRCW73AFcvKSpEv4DWbWIKIA6vr96vwq7aWG+DKd
PEmA77LQ6vh4uCgvNbbi0LTwFawvLkl8VZjgmdh5CYINVYkiFDXPy+Vp6hlm93pt
7T5DXJKeH81R1DDN/fHS0GysyB4fsZtajy2hfyqyYClUVOYwDwFIRGoKSwzApec1
2T93noaOACukXNmZ+3DNxd5lYACerGqaAAtVlApp4jT6KwOYFT0vHx5pcXO6dD07
zGJiL3Gs8kyEuu8zD8c15blBjGkT4y1of4+8bednNBUHtlwfDP5qZSI+fOKZut4P
o0ss225PNKs8FWNkaqc2Iw06LCSoG3S5bvV1bPMQ2mPbBV/X9g9iyND8uPG3VNv4
oJyuVd+Ln4fO9SG7IA0IB27bGxD+A1YPxc9v/fUO/r3rn+kOotbQ60LGUWlQM4Eq
OyrRwlc65D+pIqLBabroUiV2UwvlTGcm8D8xLYa6zqyzrQCmORVn6nNBdPt+L+AS
NsEH0Agbl3uPO/Exy9Mx61aRmGEG5jxDEsyLwmVL944DqhwtOzI39ilVDONu120V
zrfbIMZ/B8BIqLDgjVRsXX9GtY6WWE9VWPc8u03yGIJFznUSKwnsL5OoUWuc91+Z
/j3weTzoYgO0snbaZXq3v4A8skkQnLOW+Cviz5YMX5F2rP6p3SRAKsEmfCuIzhAe
/7/w/H4Fy9YQdEYt0ahODLvHZBEOkLoi47KQ2Mp5/fv9y/MPAymKVVXRNsCrPI1k
e1rFhfEn5+QUvDO0WSNXIS3UBw+LhIQRgtnJmsihrZUruG1q/JAPeqbcZILpgRvY
/PxDoaXeW5BP35dc6FTSmT8PifkzN2ph2FttOwx9uVv7qpaKwgiCseAxNMZ9r6DF
xbCTE0EUFzw2veb9hGj1TQcmUdx16FR3qXqYmYwCbhk8TYgAfy/R0zIgUzpw0KDG
CqYGX849EClLpSvS674wgpyk+m8pLL3I+Iyy3wtDDdstkHFyIMF+C6g7n5JCKhuD
A26Td3DbxJd88lQXpApn7VLm2ymI5mF/V7Wko//emUcgLoSSNHZbJMgXsm/cEcBV
0Dt3t3/xCgNeWNVmrJ2fw9mv+RHMBHT3Io8egHrkDyDwLDhXSJ6MVseJPBhFVnI5
/9vVfhysgs4giVhm7EE6hAA0f4BGbDf29dkz5d739CudJpr1tbYS6R/aBlO9mahL
f5EFV0aAUlJ/a4v0O9SBclrFUg3MFHM3m7hsvGCycGR6DSXe4Dc3o+9iGFcMVNt2
a/7NG65guXQGiExKRIlTBSizYbnD6DL+QmJZjZ63f7toceSYS5SUSnoZmyyjOYAm
eRMLRViq+oGbIE3Sfkk7+52ce18tKe6o/Ssbx90PjSBfbBKDoNQK4Ql//G+7MP0v
nmMDU9k8gounZSX3+5SWsPB6T8zrt8pHmFydJK0noNGYi/FWRuoiFceAfE5Pk0mI
lDmkNY4WsfrQVqM4Hngy4kzr43JYF/HL1n/NUqu1VUwIIjdS416/hoKB63eMoFZO
fNrTFIFnS7JNlngwu0/BJefwul/7LVE+hycbg2ksibJaTxBFHS2QP61mqWo2jSen
Kux3mD+DiLAy2vpgWZkJ2E1cI6NS2g+970OmPo2OEoz5Fj7DN6p4W3jWC/24czJJ
RolPmxCrboYujmoBExL6rnL4X7zqQO/XGa40WEMVgkIuZRmtcqnGovoY4gsvvEXm
8vgyZbzl3AHOJN053PhwU8rEnAkBvdmecm32zb1q1oPUlDBidmx7E59hDmY4kzYD
qYTWRk5OnHjZHbBrvldtXcEwc5UpFejdYQ6Zu7gnuY9F6TnatpL8UerDN5TElO5T
kezWTHP41jhqVMkO7KgmNkyE4u0iWfHzH46TloENVmlogGIlZAyGJNjMIjAs20D7
PqoSHYn5FGOhetyDXGrHU4Xku6X6EECfe7a4VeGm7VD8I0uStDAKryd2PN3Dw/Ly
uHwzOxh7CWIqdDQlF9yWYmirZ5mQI8NCHD/0hh+f+E3GiGEUl8/3uK7dkcfkc60u
jie+cOXVGidZDrt9uWEfwTU/SQJXkUPOnTFBK/t2LrUq9IibRj0B0QSpyCvd4pne
AG0XgFDtWrYKbgHmMafh0D7Wk0HOFgGZyESVDohdHpR/vO5Ay3nmDcvp1c5z29kW
pgOYUTRDP2GlddZHo20t12TR4EeswxS6XPcCRLO0ICeeyF8pf3oszUbA0B38G71O
lgnNOExVNc4DFIPqLBBq6hi9fo2eNA/S4ETheW1mYyNupuNhXso98+lZzQ6CfBmV
i1Nm6KxMhV4dR8lzjLulNGrSnd4c7kGEfOrCNayQcsiyRsU8hUdb0XfGiFA71xhN
iRNsuPY/VxjI1dRNQtS27DJAg5ecjLxzmyzMYzRRcOGOG+16U06mv2vfGYqJoSvJ
SM3bJOJiY0ZxHcGi0BkU/36APXpXP21ylyw/y9nz3MeFacfxEH4R/BO0lK3O8uzw
8NGY8Z/DZWEoeRbEhZDrU6HU/EJ0vGH+rneD0KiNM6ESoj3/6K1g5vCQdMSavC3a
HL8yosHhO8TKB3mUkgmNfde+EJhWC2fCjz1N+r8OiGEfjcpiKx1Ebg81k9emiEDA
qx5+V7cqa8xTgNenrNuIAqOP1yNlUkqGFgwnLDuHiLzhdhjktyx5G+R1pGnnUKQM
ofQ6YItCMxa8dCFD20BUfaDAq0DEkdWzntIYOmvJ8eO0ySgt4gZEDKh59a8Pa4Cd
wryXvWRuA9YhMKx3UidO6v8ehqp25DniWrBWpiuD/449B90Z7ER+1ykQWKNLx9qX
yqYH807MrF9n7Vd4Ois4BTpQJ30zvxVk+xTzYPqlgpS1KD19rtbvPNfOuc7Lykdd
k+uEZpbhuYEiLmCwWj2T0cqdoZyma9MaHNDD30CHtAm848gjTe1Ov+N/2psFtL43
kLHDdQGm6Gz2vL68h+40VI1cbN5zg5tG350wEdfkRk8NhMRJFYvnM9nHMU+VvQYh
+l+A1wjrFoMq/u17k60ANiquYpZ3wGW0xkaUgiV1odXUXG+mpdexvtHTEW7CHB1F
33KUU3mnYKk4Slm8FjPB0NyRMQOMm7v8KQyfeehy9+c+RSld0D7b09n+0ai+nlZc
Dm8ne1FWElE2W2exsQVM8sTc3y+vuoMF5EZuixM5KfaOtCt11q0JqU/TMLsqaEpo
4DhVxcWIjKXjOSI4CKyPF7Sb/45CrZ9d2XxyJasldlrimGXVYgRo1nwKHFr/ifLH
irkElWcOvF3VyXvFNZ8/lhm8qBMajyzrpvR/lKimN9UGJpNxE9OPqt1XyqUOfOZs
9WNAKzyjnGiGuCT2w13Je91WO3RAE0OKoHI81Ka0l4q8cLzuXG36QaZ0CapnB+u0
e/Ze4XiHdJlR5ukBR1u+yojGMEIk18yY8XrYetIqyxrX+QCQFZmJghclwNaCSFG1
uOUXQ68XDrdt3S9fOHED+xOKP4qr/FlgzMXKpTfOTFCDe7Ml8U0Qn7aL0XKWo+Cz
jFopFE4Rvu7fWx582p/sQGYqTUFEHd0+CLPp/Bqoiv3hb92ctKXrQ003hBVYwxZk
5OcKe3WdjyNd0cIkTPkKXxExUevQ4pwrFDdHKH//FHy7VKMzXo+DoQHjvXGFxAsd
/n9Mmm3G6QSiBFwfKaHAZ7gF9gjt+FPVqnwnpl795eFdv37jn1j371xDYKxvR75x
HsOKWnpzckEmwfuIg9wxPjPcWWmpBteAdXEhe2Dxuobg1iBXldgOQTFnJNn9QtMW
DWreVkdPjGyf42S0gAsnnLvj2BK6L3OMDBGOogV39pzJFAMTrFUjvvHJjL7soIHM
vh7M8xn8UFhusYisMGumz3qBCuhETYPBY3pO477vk3mfSlA8zrbu4cQHIDbwiA9B
3gFlmvQYYE8oVNIC5Qq5X7jGr/O2FdPvu36hdu4Qo+AtGkQjMDOjhQMuLYlJd+4u
1ysZ3tpi08k5vXdR+ioEhuJBx3G/yd+Dq5m4nAHN6UA4fGuaaC+oxGpE/rOTZPYD
LR1RerM6iqOZwXwl9ij49iwoDOFvvDuAQFzvK3/2FzdW6mebSNf9nQP2LU4mHBnC
eHpZ3yUuh1rdj3E1DnVAw63Lpi6Ls64LeZj5yBmZKjLIQdbz4lVEIUjeCClkw4K2
dkMOV0xM9+43myZiAj5iUUwU42z6ihcfJGXO9PoNjl/gh7uWvPwl6hJKZ9vEdaX+
P5Q4a728thW79SAfpo63hXK3ELe9KwYeZyyj7ihj/DCEAN/dmAyn5NbQTQxFmnnB
V49xfQ0RnOXhK6WplWA1FF2+jnn5j92f4i89Q6kSiUQfi6AKAxtrLo1aw3G8AYzi
iKcboSg5PDQuXvMFT4r4FIF7PPlVuEQCnq9JyP8JVYBkaVAeEjZUl7Z+I7q8dLtT
UMvBDsxucWaj/xUI+Je+aueu/zJIBbyZ2H3lf6mys+UdW+S3NHv9W38Zz2q1UNym
G0kYmkJMqvIHrGh3airEI7tKcH/tnf1IxQMc4WU/a2I38xwyw4GXTRIhglPGEXt5
fVr6/zkWFOgNe40ROgST7CEeqr/QqGGJc7gTSDS8SAmpuOC2ja8mqSooJbp19ZG2
J8yAbtrehjMkKLCQtqSoXZElIxs3TAJddNwihR6W7Da5JSt1V5ClRUfXq9njX7WX
/il8ceUiRxP+OnfjO/kxEKmi+EJLfwMxBI36QsPyNv8TVsBHjBT63bGXa65jy4G7
I9cVKtPLVM/Thyh2qhU9boNfGuAqCrJQIKt2IdNRW/gwk2xmEe94AUG7nxTJXHhG
oq8ScUc20BdOPSmh8ONaeuehHo7yPDaNqxDvLMoevfflOj4S1o0owW0Z8XwgFI6K
8P/WaWkNoupXPgZ9s9zQTUwd5glk6YqDfrH4ReAZJ+TNAJ1WT0/O6FAHJ+9Aq2Uw
4MJe3UfvrVejSqYl8mESajXmCqnD25oguV8pWzV1McMogdf7sUufD0bnXk3uEdp6
NO0nQYYemVkPdinWP9tLJXMahd8hDgDNwTTZWEm7+isCGxGobD6UsKT0bWnovsGW
jOczMTXvej81aFUzlJG0QX1xuZSuhTgrbyR3Df0XTjMgnvfXUae/mwYdJAtXhFJ8
cBKsq/uB3BSlZnaYzJegSFhj91xyA9Cpi6GKybyEKW7yIRj3n9270TEVcmc6/e+Q
gt110af4uwohncCLj+7v3/chCuwgs+QxFx4yznFzhOCf25GSiYZyse+LHbxO4FtF
qq3ffecX6yFR4ZOJsOFs3yApvW/EOahuK5Vj4lZ+MwmjKXRyJzxSFP8SAj6c/5E+
ylWg/t9WsTXgoj+3kTYbDFqen2gk6UQwJjel/FXewHzDaqtI6M8hR/BlWMI0nD8x
9cf5tpnbQ1pzJPPDwzumdmdPpB8DiGUQ+sWyn+NIWNQn2MwzPzVczKr/wL0TeSru
o0KJA5EGT8SNhMu0S7wxGW6ngkMaxMR4IqsHZGAM1I/WoyMknXrFmdlObJ10v6KI
OOKL67MwdWPyHWO0p/3DX9XTUHas9mog4hASQkqqXbAmDK9tGTraz3NBR497N4W2
SJ/ccENk1zBdAvV7fkafDTUca9wUliTmvwR41OvOlDjkOUPjDkPOMJsjpO5+lW6o
jxrAG8+V7qpsn7tZK1CO6kPR6zpg0RquTXePF7V0xrdcWxra7IjNsAORUn+nhbl+
06/VqGWoUAJgRBVicml1rh/GKpWc/EdUFwhjzNiEU89fHUFp0eKkfVSZ33wFKIgu
+E0UBSxJJbpaUBSITY6zg39vODh4NG39jqAWozZhe5CCmE6Kwbp3E/8nS+t6OCFL
+NLE7HU76p/GU0HFf5TbfX4e1SHgWK45QeYYBY75aCUZIi+tQmpNf6ykwfMlQuG9
i11pCh9De+11GiSfWiRoNPYsl96hTeXQbkyphiaNmliIVIwZuFfCdS0cburBnmem
gK8hPF1QUiK5zojkgQBKgUcn/AP1NJIowHgyke3rkzS+ZcIAfhpG+zc7MVwB9aOq
cUHVEpkQ8G4eIeenh9ypRokxv1bMmEBq1x/d2e8UjyDYNpPYF2Ud7PROjzY1DXxd
EtTMQu1fWU1uSZWkCxFJjtjDKjxG+1KxQG7uTqS+sD5Gse+0D5Sn+RnnsgajPck2
wOnP0779BWddoJGGiRcF7b/++yf/mQwqXxyt8bR1zjdFgm6rPc640GTphFfC37J3
oVTg3FeZjpFzAPHwOa3E6HclViZAH0IxSWHG7r4BN3c2OSAprX/XXiYeyjntwqpY
AxCzXm/k8rgSPfeByanH/qoGdDEP+Sv318OuhHDUPN1ErNYpFsNkSoQBo/2GoDbF
2l+GjSxn9xfdtkR/5JxTeoAuWdS4tTyEMqZnp95OZr8C2rvII+XMKhKBb30GdKjn
ZvWjI6v4diAzROOXqV/zSKRnQdoI4ieU4ad6W6doDJCCPJAOdjvhDffeV5sJ4ZtO
J1ge7oVOo+IGGDf0fiUpkXBhCojJQbFdwgwsqorTI9mhT7U012Q6rZGgZBo3zhDX
AkgYTvDrZMlS/GXuVGydPfwo4F5sTXzlU+9rrtDl3p/IIRX+R5oJTS51xkBG0IpI
nLjUB/e1gPQoOLdNmJhZZ4MPnbdPiZI4PDYtUgCbwnvyM0NPRM/EdGZDrvnCrEV6
IhGYlY5AmFDVSUi/mElCoN4Dw6Eqz8M9cRn6eSx2CYyWCRfjMnfkQ06At3rJiDzb
b+vOlg84hDQQrXlQkVKiLxYTq0JB+9iPbDh2p661SBz1MYrWse8ZQm3HtvGR0dQa
UFP7cAQBRhxhZKayun6/GbmdRJxFHUwl20NxlDyUeQkHdLu2/wI2p3D9oS5A1X0X
dvvSxu4Lrk9XxOXlghqJhg7itt7WATc1Rg74EP5HAYYW+tgrdKgah0vEaSQ/ePpa
QxpHr7vnePOP8RqfVI9O0ayQ0Nz7KcfQNtooCiUmZ72TCiomS0Kcyni+H7g60LMT
PNL9So1IlubrtTluoVgUgmxlD14aEVEvzhYoD3AW6rwPz4DcRtdXEnzJn1TaXNtT
hzGNXXPX8yrF2xhbzwNljw0tT6YD4EDCyubKYPu+GfqHl8RMI9d1QjY14EkqUK0A
Jx/mWaUGiV0gfUp4JBAoGLEoVFwmJEE5pCeUEavok70OnMXlcQkSAySlBSqP3nuJ
ckMDwyaIwH2Etz3GJr4+0tjozOv+2JYOs14KEvrbviyW9K5uPevkvhHLyIFiP8rs
6doBYSyqSdibMFphBfT2a51xhYdAKt//MXliixwWFjbX6GaBpba1MKZuTa9geUF3
yR0F1z344U7xBWnPqVx5r+XcO/zF3ojIihpr98h9u8WT2X1YPF9JZjJu8asPeY/o
XQXzoOcTQiLLlO6qBOAQ4DNClasXXOBgIgGHx+fzf1tF+7PMkA3mKk02BIN8U5D6
E0cvIDThsAAsKue1HUhkXDXIOBfmZ0JkZMroYByYFKGzGdCJ6bvUOVOXAuRcuB/K
GKT5mcRPs1NsSonA+QGyFhjp+oXxnn6HYOZkueIR1RY0H9j2mTXCMNZdWtcOnX4e
IB5OckbtnTuRL1Xyx1fZuG2GEPSLajb6vaXgiw0sWfgIvz1+n9ZE+8ZxnmHW/DDh
vjChPN/W5r6HIOj7yWMA7kDbQffffA4dtL+ZD8f1JluChFWSmnsR9qQedoWd7n0s
Wxfr7yMg31v3XQbTRBKV/OojHydsvfS3uSz2g+Gy92Yc7J8k75HpjETILBwiod9z
xAPh5/hCO4A7iEoGScEwByNsXpd+2C9J60lh7/tSj5lv8K5ctMvn+eEWxn4c1Yzn
etGdeOeaYP2lzA4x3+rOghe3CPo0ftcdN3lHukqrj9jhkzZ76MXy4tJNlbWLqSrh
TIovfL92mUNsdXBPqNChCoBs0zDV8cNHvRRAcvbsV0gB1Orzp7sipa3BiOLPFBDY
DHW4DhbAhrPiZ4agB7wcdl6bDz+Vfqi09qfPkxlRaH3ugMeWGjwxg9TqEY0t/NZJ
gEC1tYBurDmF/kB+Nzv3Tzl9QTtHWVI5F8DST7EXRnqRYojDFOnzyU/o+3kVrHts
IJD3+muFDm958OSTVWcz5/hspB45FnzfhWt5e7QejZGku52rYMvEbM977y7ZP3S6
eACP2lSt0vDY3Z3mYF7ag8Rt2IPHSwv5X2JHy82IWurI1VjErFMRH8zf05QaprVD
sEpVUt39yaWIHqA/cB7uiTjKvZi34pqQoJHCJAceRqOg0ijL/WZRCkXqbXX+gHsL
+ZHVmWqjZlFNSZVjirFsbcOFosjHhMowlK4hvu/Ye8iVEIT2lrLGtTjiLMj4V9Q9
I6uICO9uWDpODBi748zoHTEVGblGjriaMKGZlL+6ZCfuus8krgxoboh1sUHRTKMT
imYRgogGUMwTtwXeCzI88+gYYwJxeCZyp0CnC6eCH8EzIHv0uA66sDG61LmRvyMC
NjdxOE1e1jDDtE1ymN5/kCNlO/feIQALMZVO1zvDU4bpi3ruyHqnCRChiI/Hdd+m
wr2LNulWuFEBwx/7S7nI/ajVzKMRvpzuIjRCOhx0z71sgmQ2GTYnIgmcuWmiZ+e9
ovtm/R+qD+XCXfF4eTkTXxyVgcWu7Y86wz0ws4WcuitSLdWgmL0j2FP9EnfA8D+l
TSsucsoYOF3GuibkAXp7Aapsp6LyB/8K9a3xgrsKA0WRDJ0NmY+u9m+8O/SK3qjE
i2JsTZZmcfDQaEXr0b1ks1WHlDC8XF5buLo2X2gDdTeP4A52IU9K1e13YDIpicWv
FdOGXuUmET/p4MPff/dpLTXnKHOXZZul/j99a/EtLFjfSAZxdcJQWq/rn2DmVdBT
s5lZytg/GOZRrQcrYkFKaBCC1N6vE+LhYclHAM/0vFQjK2gbdn7IpL/RQImI4QKm
aWf0hIRW6AdBghZFz22ttIJPbPU/xNCamYB78h9hAc8+/lgi7dxCOfIlxBXad2Gx
rXRwqMzaRIIvgwjT4hRTwnoUfOywHe+ndFcnreNdrNmOyOfAHcllHzsvMMSA32nb
MUJxZiYbYA43f2Og/9nN0sOhrAYUhYyO7hxiwBRidtRpJbhATdIAKNzl4gfHhJev
IjJ2e/LiUMjWNgRk6p1Aw/v5Nx7ZlYzP4YGkwu19G6uXSWlTuSJhvDc/Yjn8GBfP
DXQv+L9NHvfNKfdLpMdp3vi+l0YWwy/+bt1ztwnsCktr1K2SMo+WboWxvsMk2UNR
uODqoF8abbX7IDQbbOM4wP0fdcXNZDQvAbyJ/P5klceHoNnCRqqSKRfsPyrZt/EH
/3m9ajkIZiv5/apkDTTwsVHP/2Eq5XuS2NZtuV8zLUNDJwc/jhVxP3HeCs05QEex
dKfiv6ASNNCcIg+VaH/z6rnzWTEqIThqgj7ODukvbEbkHIW5Tpcvsf3Hwt1B+O1w
+00y1Nvb2Fwy3bxPQe5q/RKhUFBYD6rEcpFNp9hGMylmDEqWQ9jwwEogVHEFIEUP
MRt5Hhvr/pkJ6XRNdxp3iZSTqw9N8RzSgUGZb8Cl7XsYnK3wQ1JhQ12k4vs3rnXZ
2oDYgFAXdfY0+TSyfq5L4yL6zkt2BtcaOSt4/Jr7bczeZr5zglVEbODYuBe6x5Kd
aUB/CiT5WY5cZIX3HdikBGYNrR7VPWyy0OSxlk8GheOOYt6m0DgQ8UNLNwQqMypx
Y0hqq5z4PP3lp4M5f2z1an6ZdS0vxHig8mRWsLKfd48VczUdcW8hAHliqOuqPU6/
cT3k4U0Sj0rktR5U0km+EaOJunEjRlDXHxsSsJBIdGSY95L22nv6BNXptQhbWdq0
HqK4lNAUoD6qn5YXHmeK3zcM4qf+CwFJXBv0qG/RSZTsBhcHrt9bZdiiovm7st+5
n+QBfbIJo45IID7CVQV86Z5j7HIZreG/HuIwX04Cwoz4k5TzIB0aTnXe/dkR/8ud
DHYbn6McJsM6SNDqETpK/jCXif9bysGjN9PsB0y0zPRocZco7lFDvgozqYWuyF63
733D+zkPyO94i0QvcmZRIoM4SZWYWYfRpbehIv5SlHCmJ0BFPNz9hnrcRbmV9Y2s
XWbS7j0S2dKPG+gdIYOYMdoWtQTmjUpq/3nDgIDBQWAzgC8qyXz/MEC8r9lWRD8B
Kw/BD54VVQxjPoeiKn0mGfbdpDd+4EVhOym9+XNOTLFGlmz5V0hkVCg+t+LXKVfm
AR7f1wyfnnfvum8ma4nqQM8AkU4FADw8XBRX8RSGiexq21yQlhZ+IEgCdJCzoXyY
Pol5JK66wfQhEgwRuOGYG4Mt1+B092jNrJRG68FhBR49OsVk4PdoGetRDqwUrWiS
+oes13whELla+nTZFjwISZt9HXpWARn3OVOPZBRjuW8YbsEKFm2OCizcRLc6KFt8
2wYJXeJfn1iJKjm1so89ludSZOISELIogV6Vj313x84XEZ016dAFyWnH7NYgeBvu
Jn0Yy44duRdEUoacgdo6JlPFkU7h6ALQcaaalbTVy/kVQ5cxBtrzwjcB9EIT7ZHs
5n5xDZafbrs7V9zTZVdRPAU8CfihW1K49lzcXZdVgh9RkkfU7dh9XTFFeZBVunPf
+1ZjgZNi0zdf6yyalLqlXv7NGDOEtJsE1IZ6zejBFbfPufOWCQY/G/QGTusjmkiD
VHCgVR2X0QvJXYYxd3+sucdFE7x+Gx7a7QsYJTMsMtY1QCLYPX/Z7Z2SUEWQUeyk
ifOf59wM8UqTxR1yzwqkgHWcv7GkypZP2DwkZkHDRkp+NgMqi98eduhRJKZadcX6
RGS9W2nA+POwC+FxMK6Fjno7wEvkTob6VVAm5YEeFQbVzAtsSyfNwfiGzIFKxwI6
+unmzJo8trxJTgTz70udV0AsiwxU1aMSE4pJ3YcG2nkUE+bLiWcAwrLXBipz9jf0
4KGHOaILIAmOUP+A7RMycvdLXOqwySuyo1ld4hisqkRs4uNKSfTC9Fz5rhL3G5Fd
/lD2hLoCithgxgi01qlQmyCnEMF03BFfdxbNFhbqO5BunrixuN+vDCdCcsodTT4T
oBR4Emo7FtJbccpj8XOuGeD6nu1VAbSV8/52sjF+LV2eAJMXV3KT4aRRGMybKIpz
6uBE8MpQET3/uwTtadFlmULTpdooBzhJI/WdemuI+aRIq/NvXhbrw4S1JhKlKTyd
wg7/NhklvQVCBd6PpC6KdlCjDUFWXzG5bDEgXDabw8eO319RlLSHvbti2b/hA47W
XU9B6a82Wuyh1I9s+o9wrGnGJRvl90j5Y4cMBgScaJU0XzU8cnEH5dmrExx4c2eb
mejPxMVRX8BfVNCaKeAQkfr7c5N8ehez+MG4vOvoZmpvRTLRfvjsvoZipCdxdSg5
YwWHMZ2LBTr52KjDSH6lFRnr8uDfn/6995TNRNv9SvLpV+x2NumSnDL1KsxHndJK
1+4b06p6wtzXFvUG48NPpuzuRWuUNgDcb5W4YAI4p9m3IasZxSOuF/UfFVR/yVhV
qIqJ7zcVDGFeficJ6uewlR1w2wtjmovu2Rll3T3/lm34fhvt5arHu2mYgtJuEV5+
sWZazRvoaLVkHtUndYzV60S+uSj07B9RXTS2KZ56y4waEebxDQhoox4NrGYpIs52
+tBMiSn9fpS1yK+pVO+r1UCteoogpaRdhmfIyDTFns3vz97z6qE/notvxc95vErC
cUFEdVBC9IjSh3hNjn5YFidilN/j7RcaU85MBeeG9itrIXfWq6ZY8QPhiL1iHCMW
iM6wClYQrt908+dxTPir1I6sxgZXC0q6cjtdSyNZF5SVskI274XuwK5+WrrVifCo
xLgUf13h6BgpnWmE4wfp+T1PYz8unmciIASyb1Z6IeJCOMM8G3qNgd/vAXeNqDbn
It01QziC/AYq3c1jsM9eOyl8KJnRy6LLVRVUE5LgIL49h+HEznVf1B6KTQlQ5W9x
MuWunzn+Uk3f5fjtZjgtKoGLK1iJgQXT9PJdYS5ALXMRuMZtWEBPr2k6cpynKTrG
HvSNp1JITYRZ4sZXOMf9p/0CO29zaY7HvNR+FAxIOME9gZibsiKgmj5eSqXxPzGc
2UO4sgebqGP9AjXI1tpV6x04CPrGqOphvGENx6u5jfdY4z/j/ea+ow3TiWjPzNH7
YmEI8MubWAh2sGb5lfBfzy8e6k+x7l4VxSAAgbnmTQy9Qe8dKsFQlxrxUvNZx/fd
k1zO8+nLTdmSjs71xwH2iqW2DO4dQtgrIDWYnz9qyt6A9qDZXeB2qCxfY0b+jFrY
96SftWHMR81ouJmOKTyjbak5Qx+NaxuMZh8lIa6Mt5dyz8lq81g2EEyjhkLS7F66
5H/vvVFSZcP0RmzDwlSRPcjIeYFMgG8rQqHYK+ao33mKiZNWxZbJcLX64k5e1CQt
epgDXMeC3rQ/EHSu/CilZtHOPFTeqnMEejTAPB30P9Hva6EU5dSl7G10iwGk660x
LodbGJnPuBr/ih3O87PAbd8mgfvOeV1a4weFTTtZ5bLKgResdhs6nhDTZcpIHR22
7S8VCiZMp5cZTbvzXREoOaEnfCyE7Ao0Yn99BVJXs8nXhHqUR3FfIpKRwecm/6sW
AWmIZatH3yrQNtrbdT/oXlp6xxUnBViATWhi3XnOydOhAW2uvL+S5//OwQMz78O/
MzdrBkQvamymve2S0AXfDLwXQ4TpHlX3bjweKCbEBE0KZpMXHMM4g8fjpreww3LA
FfpQcJVffNUPW3j3F0owVnzXEAGZQrLXYDacGj40ye6XIxDjvyiFibd68uzdc/xY
VTB+49HAshqBOkRMadGB4uB/bZkDczAlYDZ8O/X53xL85RQR9rOBNm1IWnSjJv8c
lfw7czcOXpy0kRPurhsnEWPjvX2BpyUkIL9tXhEdh8oF/ZveQZbUr7R6/y6jtxy7
gveVf+7GPNHYRQuwG45SchifqLWyJNi1HQwORiSye3SJZ8EKN5TlvjQUh632GlZK
b4fKvW+Wo76Vhd9tMsME/2DkuX85f/xhuDckJVQGuLNo1AXCOTrL8plkTOL/b3rJ
RU5v+1PVKztlPbPz5IQP7MfprnCulXpFDcCfatmf+gaKUXcLjBK6o4lmD5W8Yy+j
ERJehAdOV7MlTFEkiusOwNO8/VnNVXh+oBZ4LuDw8s+IzGMIppGWK8AGSbyHSj/w
IkZs66lgA+Wdt1olHk7CtSFJOgZFm/6QilLXvaosnUJayQEz8YRJafNuyzSEgBOA
RHfOMcDcWAnq128Ici/X5fY2Trep4QfBLsE+1NGmtoqVYGvKkvktHWwefq4qfbSZ
ij2+x7t3CiNCfhTNv2NFEFMXxOQD/3O0camvAsQxhaGz2utER0UOORkvD8NXDmkD
fCeJn1WlLCwJkuJYw6WQoHIRZ2jsLH+yrZ8gYdfx8U/G5u+W7KKgaxoLxhnp4Is3
XTdQlbGROo4uafhuaIScrzn6yQ+qgaNjLAZ9Mb24TLUWsNpS5ivn7+UZdWpharwg
djHuHqkAIU+BUcA/Y6PFw0us4u7Ffq3WhooR3biCsUQ7eQW10PmLFSbeVgbcRlUP
pMj895nyUkb35CD3CfeXh97SRjUA2D8yGh9Lt8WdgKIdyRMoeRaSVXMxvJuJI4KR
Ri2Xx06G5RYlKbeha62NYeZWjQKA9fnuE653E4m/vnzwiXgxgiLb09cT2JzxTG5t
DHTg51l11Rm/kOgMuXS1G1koMFw7hOjf4CUPLig9TDPeaqJVMny8PNODmYJe91gr
unt33uxp9J1pUUw8MczjGfz+Qf5TjciTej376nIqXmEdEHzUcMCXH78W50gm9DB6
qdF/5sCkFEHsZqi0vFy7Ohef+CRqXPyZnA15TACJtCVJwGTDTDxxkXbeigO9Ci8R
3KCAm7I7m/uTM7JHFl+Hnh7fNRcRGFUUkN6OsBpuN16aHZ2A0jzfMK678BjXxg7M
z1Y4Nt+WrlpgdmlT21pI7GS0Y7W4gQAIKcDXLXoIkvGfroD4go7gkZNvoT2oAKAE
+fus1a0mlmIjIv0EcAkKcnoJGz9+C3mp1+3QfcYM5Vyqb+rE/8g4Smx8G8TprOlA
eZ+WGTGt9Q6p8Am/2WfpyXv61oUGkcz9xSACLk6UByGU6l4pmiHfueMrX/hCcje0
tTIWvn6Yw/fpXCYsNwoJr3XDgoJ43avP9zrnyZp5MY7vJw2nZfmzAZXNYG5ynLJx
2jwH6segjRrp+lVAZFtGf337bK3DZC4TLRlWTm26unxr3QBSuiF3/Qzz9QPuPk0t
HPocNataVaI8yLe9RspTPB5SMcBsvShyWN9JlFpDQgLpsrw7xlqExSv185rURf53
Wee4TbUqIp/+TCC0hSDMV2IYf0vpsZfgab0Fp/MkpBv9mVIPc6DznJaf6B7ENTPm
Hdy829Z6i25Y3+7SDjljk1PEFPleSteLKhTKIPYyDQhCULPF9nZpgXfJo+JPvGsg
0XX4kY9+h0vyMUoL3DbU8rvbn/M2J2NT+I0Ns6Zu6ipJgYlbaiIJ9LxBDdgHXsv9
CxtNXCKW9KxcCJ0pInLQ8vHLDmVFMM/ZiBQBsW6L07QUhIpk1GtqsViAzom6Yf9T
KIDGCWsTb5yt9rQer937l4dOSPnaOi0+/2ny6kMVnr7TcaZfoDotz1zAVfDyR0gA
QqCWohCvVghhUn1p2JOIQwWDgg5M0fKD31grLq/VG2AH72wFXtQGIFN6uM1Z1mHn
3ZiEaast41pNIUNWZ00y778M7Rzvr1zDUR4W0SBPDTOKwdr09J/8oCejR0ypzSdI
ukONYG5cDIfy6yM2zPhjE6FZpl4Ik8WU2HViPPyVcCvPdi5/Hv/e577Dg/5gopUm
sLG5KXAMtYJ9z6tO9j939e0XSEf1ghOoha9BuYTHuG2EKO2VW0nyvAb7D7fh1EIV
j9u4nb1/BpvUvgvMHZ4Xsw+mGStdvBciOmUl73w5NdNE6owRMYezadyTRAn9ipDi
2VyUadQlYu12VyXvz30Xh/HSLV2g40Q0fFpnN7C6vYlqFcKqHeg8l+KOtNWtEdGt
KSgglJuEFOaqX7xKdt083GgvFdEk3bz25u8ynUnNfIbhFnK6Yzk6GYhYHvYdZfuB
IJIf2qlquZ6V+0o+YLY+73nhk9ZCSa353SmvR/Gn8geKX7OchYwk4HLhNXSFzWpf
DI7dCj63xlJ0Zun4rRnjHJQCzladPkDg3A/xY/AYJkcvuHFwUBg4pSaYLMzl2WyT
ilCv2Yo9LroAKH7hxe/u56m2LAC+/Y+7ttfzcdvr6IU/IJM5kAu1RLCr2V17qmjJ
2RAVNIpel3qghVM36tSGyA6n0Ks1yRshtzw4flFvlpyUdaxDogHmmWdsOcYPsSEd
Vo4DJrrv05711dokjM2GVGjPh75ApdCtmuMUoMcBqoFqjxz1OeJhpfd6FJWe+UhW
eYB2nH/1ferwKi8QpZuCYvS9jmez7ScGLYXDr28Xi0aDEWA7qz9bSN5GyTjswamf
zug6pNd12cdndwuoFH6IuIEBG9KsYyeRgwRPGlsRmLj8ooZ8C4nz37W2pXMY6jq1
5eVia7qhAzCUH8SJapGVk+hydXjMdrSOQ9R4QdX8e2/3GbfhAxparOMSjsAURfCl
IJYDPS7e6CZTsV8Mb6VEpCGqK/byXWOQ9ugBaGYWLUtSeNfHORSHM2JUb19636GJ
L8YscvOnIEANeZp5M9y8B6vST68kez5flCn+DJGs1n+1AxJQjhU4DkqL756P/o9R
TQjbjVIRPk4rfS/2s/E0zT6tflXLthm3y3ez5m+mcVPwLlR7XLR7L4h/dvs40Dcq
3fyA5MEq23jynT+e+765UC8a6/bjHZSfbJfRjOpQM3VXPtQR+URnlHokQPR9XQya
DObDBV88EdyZP2J+2c4Ws1T1APAEEbufa+niV8BiqFYRwYVzawbiOHvS4jGahO+9
AeT/7f/XtsjU6JcrjSwd0bCTUI2tieZe2LNIEQCBLwU/rilV+GZ1dIZJEqqSsIIC
GMTL8nYpV+M2Iv2TYMSBYRY9jgzDXL1Jak4MNaHzhcU8nle1gKIi5+Zh8vm+Xuam
81Qi8eJt7GfUI5tB2Xtoo4waLJO4FPoFoY1zz5CHh4yNmohVlcXgxIvOlXrOSe2Y
Me5mKfgP1K6kLk41DVI/WoDSgqAHqkOLyZd7jg3Wf9dGQ+6eKTWVxSqcdeXGit9h
hypuef5dXIJ4cQpMB+7hlrWsN9CY9ixqnTytPjh2OC9r4oYl0yQoQivbViAOLb40
i0W763tjf/iNI94eX7S09odSjqY0pEKzlfuc5i2/ryM4wkcbEwY7ZQH7UpocG9DJ
9mvaaG8axFzaBZVNOqq6zd0sWP8ivQ/lwJ3gH++oArM9swP/R/lUcSxaEXW+rGR3
JvA1c033BgNAvphVy249QCPqd1qPSYTmPWmXSlzTYns5WReth8/ZaXagF7h8EvPL
IOke+EIO9uavdrn279hqgZIR2LGk3H3LVnpG/CBJNSd2UnwCUapKTkDfUT3oOlJ2
SOGFFVYym+SY+bYayV/RkcUDndzaUL+hN8SyJWfGfQk0gYLit9/NhHhmHswsE0DY
SODpTSgkfnVw1ob9lmwRBor5lalVDZ5Tm/3DpFKod3ypwxr6wikx2JKcICB8ZcgV
SOJ9wxbr/BPqRsgu8Wr02D1D9YWMOxnAP6nbMA8yBn0gjkZpsn3GnDFj0yS+BcEN
cOg4I1eAj6d5WRKWLUB8An5wv/8X0Pz76mZm60wicCCzG3M4zqXCV/kWJXla8En2
vyQMB6LCrybq9QyVGvu4YkE+1cmDTiKTSiSJ+Ge/dpxoJ50nGpOJQHIfJUu2u6tf
UMpDbDnMWTJ+SUbHD+lnTB7ssgZU6Cpp8Yd904U21X3rFCS6Wv5NFUw5/cAJh8LV
ByHCqdn4MlFy8firwcx68EiaaWw9VJJioArfVlZUtuALYJpb+KSFakk4NYhA3xAe
gZMb5SjO5dxry8G3nWJHu8Q2aVi94Ml9c+1NfkgbmPQCuBsgj8kgmzvDFr1OnFLL
oEbsl/HR4uP46S6bCtO03LutmeXu/kgX9upCX8ZSoMCcuMMj5WmtgerXmdRWw3M+
F9DXBTbNcROIejLTiYvon1Z4/7ij5gSoAku58rkYym7oFhv8d2/9zicsXPMtD1gp
BuYkihH6qHqvxzGOCqN5FIsXVqI+U+I+bZaBYpABvvDYFeYlUKPU86/3KGD9PwK8
RvBki/P2T9e++SyZrGr5ACP/Csj5aWYe6gwkaCcrpxxIq8sczNMs/yuIm+yagxNG
qWNmuc9v3d/VQ7USZVrR0vZ+Knqw0wOXs9AC7VTpfn8t4nKxU6R1FP5qNR5CPiGa
0LA+vq/pymw6XJgBPK5eXhOgpKdz/26JN0dzHPH6Ok1Bx95NaOaa42Wisf5TP+z/
X9xlYqH1QXK6V47cz4rqHukncijt/ad+pl5qkZGc/knLFgB0hx0x87BRB55RZig9
I3kxrnihXJEq61A00bvgu9iHIjo9kKijqb5bD1hx0mfspIBLb3j35YePd6O2AE2l
/+lLUwnhgGovyfJPSQH0v44Ati4G2RhoMYzhaaPss8yzwCR6tLdSV+hcdigLwI6I
2V1WiOHmBy5NK08OMYjGsdDyLF6qWcko0VSuqTiOU/xIR7x0ND1rnDZlEfeMaWIZ
lIyy/rp3FP989e7oRySrBfpZLnm8NtBiecBYfAn3VDgJeD/e0V/rcB69M7qKr3BT
be8X7I9UYL9Aok+UA0RVljj1q+PYXsVgdXtkl5y3Hs3WoW1uZjoD6hE7CRkjouGi
/fdh0HCZj7FtHhov4wd1b6lEeLEq0LxZNns31V8H29ghSr71p7J8qQJzC6gcfDko
HjKlJSuW5ILvqcj1kGc1M2ft6zpkW2rdgwCCv8xHb9i6iO3z13jWLQiDId6bpH0O
W3eRvd2gzAWLDLMuevDF5GhHjucW1jV+OmHs7SbmIr1roATGL3SE2uhfFrrRaqk8
z1GFbb2fgGnBoC+xrO+drwtmHKscCp7mNr6Z9dguQK3Tvm9fCdmXONZ0CO1rsZu4
KwJAqZZet5SNyzZ01JC/zqPK7XvHa/SCm+hBMmSajTPHE/Hz1ftIZtkxPLZQ9Ba/
3HZKV9FNMThzwJMfAjAMIYkVMG/7Uj63MIY339KEdJSznpkXwBoUlr0R4q0Vxx9N
mKEMLRRBLBrrbIaQqtaJbWx2DENTOuJoCgy0MlZtfMQKGscQq9Tl570rENJkGSPr
F4jAbvONJlNJEix7Y/9euQb1HfJrnPLrS+OLLUAxk/1ZEyJp/Ag18w7bwWYD4KDt
YYEFNPFPYZCg1hxNUkehgCGNXGRltP5UcofEpW30sNKgch0oPNpftdCmW73OcJ/C
YPrlDwkiH4kVkJy3PsNwjx8P06r2g2I4IZdOEvuHELkcn19vQn40O9keMWqr36il
Mays4oYmRBXKj4LVG7+EsNuhzzx48j/ERvZndbnAq/zFLZYL8hkd4b7Fz1qC5Mri
OavEZkMBZEzzzy9iPeC9K0fZeTHEWWSWvpNag1RuXpMrmZqWpDy90axJOlRtTLPk
1r6uuA4h5MxYHJjrjPptyq3JsVpYebanGTnPsJtb17nM3Uq7MjG91QUhza5Ij9W/
jZpBP3KeKzEM9JJ6Z7R5gbhf5EGZwP+XNOV5u6oF6b5D8OnpepZd2+5P1kuzJwLS
gTWZ+uHInd6twHIGBxxPOtRKt/DlVYc84PNtBMC2/iAbvsZRkpQmTzA6aQRAnowm
qyipn4qDY1+0eGwmC4M/9CmIDFEr5Y689jpa/76JUMiZX2GA+RbyruWMMgPkT45t
It4o9J1byJhMgdrIP/WQq3ADj02CR3W5W5loHD/rNQM+V2ynLkpGZF6yzI2IDBmG
hhT1lPHSfML0RWThJN0gPlCvclbWwcdnTjBa7WNCgkGC8fgZsDa60X7IhBGPkvaC
mrl2MRNXUZ9JMyCMsWAkaMphjKps2Bk55/fn4TEeKZvOKuhYh7HxJbRTC/y9ijQj
iT/G2OpaKmMuSgsNZEolSA8+vTG3T9kSqTNqeTSE0W10IFi3mdpRdpMNinJA+NKn
f+v8KILw0+21hO238sD3muml6w+hWWdz6FHsbZoHhM2Gr0NuKJ9ZcEwSSjJhh0Qp
DA6YT4/5F/JedurJlxRa7NBvQElGoQ2FT768aohX5sI3sbrfhUR4vTqwl5kukquf
enHyai4vQ8Nhsz8iC1Yv5lYv0cxoHOe+DEEaZQrxg4HvzcsbBqst896/asdmiHRm
Hx/ZWjkUcWx9bqNaQT9fuKgRfzzLHdb1JA0HM9GhRr3UBEuJCYoa35v5OVoSnUfA
OaXaF//Qd9N1Vn8nElgeDcbs/IZJlLmyCjSPDNJnaDqy0iqKBdJogLDSamqPbDxm
un0z71U3weeBb2G5QBiHN/i7TLYs2m0dsEzC98z0wsxG2GuAeCEP7svnjVVWvz6O
t6mQpqZq5kXpufpZMhOCUcELxLp6xjhUTG1rC2C2cseCqR9xCOOmxhvfk1+q1OQP
Xp2jG+mrA1a7ohZC8Gn34wyHE8S8dhOZdhQuoMq4nH507zN7ZUS8xhPfQENfAEVD
jJ42egBwbAr+9+rvh3UlnCr4R+/Xr3faTe56JlSP8TgPIU+Wdaw0fLFmEhwJBKLm
R3D/VrZ24PEfteIZn0xO3M/jutWEvRZCUrFY5ZW72v0V7UTEnLdpoJuStVc7bqvF
4NO9v45KS0SQvZOfPw9/3Ux/ANE/X/o77q6MPFsfyd8RIVWfwmf945zmSZ+WZe4q
5SyYEsYpFz4Vxz09AK7Ft0O5JS33WYeiiKeC7jUqlryD4BFl5GZa7QlHfDQc0iEk
j5Wgco9qWQYsn/EIWdlJGlMsAtBguQQxMp878jLBhF7iFDm9/8aekAbqYP9dNvBq
ZfgZ/1VWvTd+7SzG7Z1f9hQXzMpf/t71sU7L+zQ3CEE+e4m5BQHYNAKh74JdhVh9
jh2wdHkHnGrbKRcI5K8hqUm+8IbbyFX9ceUPrRx3gIKiFlTdJHAbhRONLF9y6+KE
gk4od6QQ6oV/DuB4tdtKH8jtbaL7R3kJYCu9RV16GF7DrdI3GWX0xHFjRBUQXnaA
BYgtfRn4ckCUUMp4EnIwndj5ke+jjwyH1pja0i5c4UkS8EaK70aEPotOt1KKWNzP
F+maYuxiEn/sZweaU0xUYT5vhVKDqCDI4RKyAh0kSnoEmpiHds/+45zcyja8oWfm
I5jobrJMfdAoYC9IK+SjLR9UYOFXzm0azmCgw4Fpwi1hUkvU2aogpBs35QRzADMc
+XEqRrAlzgmcbK6kQwNGAFXq0lL/4C29i9VlG+Hd0dcH2+AONLAsCxLytr9wKKjj
EVfKtkzqPHe+3sy1/rIdKBhu9YZhHMw8eOV8sHy26+F2SrMZ4wqGPuHBVQCs8NnU
+sBiZCsLUoA+o6o7vhn0HxkTZD9D53z1AmYWw3z2c1ih2+ZfylEyzxuDigRq+5Cs
zEfRyGZkN/sF+Yuxp0bYStqo6MNiI2r9Zayqu2+unClVdg08x2veQPnootUyAKnU
T29vjCnj2qnWqgujiKgGNdx48dwZr3K+eDZ3oahEO2x/Dqe+r2cPEt5UiN9UrQzl
vIvIsHLDLswtuJffCO/GL0BOW4XXbrL47hwBroI8lE+6xdF4me4a2XDUF41va9ce
hObrqD8D4iZrM9HUbuM4dEVz+pAALC6yFpxf6J130iOBx0pQbGfkqdFMqeMDyZB+
QkcmeYrl8CwgyDQnnRk8Exft1y6ia8D/CIi0uDajxfxxScb+PsNw/qgLQyuEnLj+
Nog8ByjB0jWTS7st6DlcFbqEJ00zanK0BMThsaG+H4qT4+iC7qnI/g3SGCT44a5K
gYT0P5GNxEHZxQZ7WOlFKNk8muNSwvXidxfxak1i8L9bAb8r+8FmXVZGKS9rkHBz
8x+vcbrss+WmsodX2biDTJ6oEqiEfNmwOTut8KsJecEn+pEOnbPTswLFDJBMrVJu
fp7Xi2yX9e3KpJn9503BFKGV6xSYR8VhnyKbZ/DATJzZiwoMP0/ymBha8haR6HA3
leXEbVaV7eGBPFu7VEhKi6nbvNie5a53jqebqMeZcHYZLjDNHTv2ggJrQgJCFAF2
NfGoozoLjPtdZjRqEuZl5JLBfjanfFjTLiKiE1T4me9TaRBnXg5tfAi7K6C+Olx5
BupyO/CRttflGHeSmo/HOIlnckf0Fv1q63WpzNI3QfMWX4lNd+YiFfDzZsZIgx/1
AuasAhbQdxH/fuUmQHZib+4TeydB6/o6Z2GOr2rrqIbbF0hOkP+uLmvQeSwJzG8z
4VeOVreaHu9GuJHysiYRbk68iqaaBVdzEb03YuMQ0FsYFsMRZ1oQTNtuP9CUa/50
zt/9VoaIVUWoqQk1toPpe5Fx1J61EpwdAiuXHdPoNoazc289dz+ejnk3wNM+UWKT
vihQjwelGCB35D8iu0G1XMQed8jKO2bZi2k1QpHWuk4lcuc9dJypTqmhFkeCSYMV
S7UgKugdPQDbhZNA8ufsLAVI8CP3aRaN+cx7gK0EJz18QSrQoWMDweKY6QRHdSbO
yOuEnEAwMyEoCSAkkISh6xEiMgeZG9+wNJywyRwLoSdr9/ZK9vwHttx9HSkU9EZN
rYL7OLNmLAcLBKNFlzftr86Ak1oWBzKSLg0LjsssSWUocUVbA/f63msSpEBGJJnf
Xc//HALmkn5FPZc79xr9huCGq8oh6J8z7QSSgeg4pqq3VtH1efq3Y1EHR9rElqTn
P87mdqFCfLdFEQwIeKJH729FjyXhTAHXWmEgr/BBc/ZYxnkgpOIC9RFYqLA8G2Ld
9u7ry1puKxA5sWUMZT5qNNyyX7h2BDfiBT2GDiyAJyCODkKmVRkyijmR/iT0AeyX
1t+q3cleKAEONIk+9ikm+3NuRb6l5dL6U6Q3Paaoc7XPCBsyC01fP6KCX3vQaW+5
dLqUK5YOEPMLeHrof+MNM9mfLy2TXuNCnvd2em86ShzgOl4ugp+WoJ7CjssBSCfZ
r0S61RDrtCvMaQRME9cN67iTAyLLIWtsBYUkLRsV9gkjALqTxrrKIXC5Qih9vYMQ
tACtNjuRy2mizLUVqkSw97uo8dLwbsJQqIhUqwAHT82g5PsL5DLbKbM3QCs0jU0v
SB+FZ2yOfLJ0VBGrrNjwyxlrxkt7vuuPVJfQSxq4ExWWpVDuzwIK5R9pDBP1wn3j
FWcJE3LNgcrDOWB6OCbcFAxiVJkPWR57FSU2uJVq2sSROxwnL3BdHk744dMlnaAu
ODHYY/Yqy2y92PqXCSv5WoipnnWJUxi9Z7kJgBbZ/T42jFr+swX4sIwy3VOH6H7R
1sSVqt0no4Zz9sN+E9AVNEY0OvrdPvLZkhvByHBQy8u5H78EkvXHb/wEFVLhLq97
c3BT8yhfRKV1g8mZSrcoXBSk1JSH2Zr49SVJ6yoghg7SCQL0rLGM5EJmDEkbI70w
vTaxFGWCR/kk2oMoH6zctqbmCZG8RROqA+3/yGUHKSolIvuOf6G26Fxp0S5RvMCY
lRCHJrReAXJgFW51qa8eFuEs30hWPPqmnamM2loVASGNLhIg/H7nWgf2P2NAMnww
KS665ZavmHOBv84+QFFPYWL/J2zs7vRHMw/TE4aXBkDGJnU9lmhcco+XaZyK+HYA
LZ54Y/7TCclgcm9TvGAPZsIk8JKrHm9pwgzvZQzvsa55gAzpsAwGaieyhQENUiNw
jGgWtuMDNHO1HWqNOKbQpyrzpx9fzaiFyMtRSK2dzD51ARM/zi9YtcGUeNIzeVNM
PaXUA2kBktM+HnAodCq/Kj+8rbkw0niEo/+cayHQNYfuD8GSwqVK8Osl+eQwEthS
qJeWj41v7C/ubrsGQdAj1XmZ2oJHq4wYVJ6dYy4P7R1fp9n6AitLkOEHj7Gec6wm
1pTTpBgG1ViW2azJfnRe9vn15HQnCR/dk/gSsm62SFjebTyy7WqumGgcX0M/mWmh
Jvw5hj1ZMt4Nyb3s+xmj9RGIpXUu7U24HfTQrRbM1jsn1dNH/4duACTODQIk/fOJ
espSM2aF/GLgBEj4ljwjbcTQPajRG6pgltFnyNmwGEzuIMpue/HhHCCUUVBuxNVq
5gMLlbe2AwtWL1QhFo++jFGgFJXHfFRe0txkZfjmOpxKxSM/YGwt0DoBzAWdMpss
YIFlLieZvR53RjYB6kw8KDPNBL+ncDseXqNGaq8uK7o4Jm+Mj6pIqew02efvaNBZ
uuOlgsYZu6fzFpeoopl5sxopLUmh0HtECly2uKCseWrW9B/ILyRQifQyYTgAID8t
XT7TqBy+ereZG3W8UEzMABjwtmVAHgBWDvJTtQJwa0ovqagnlsPZerHFUXTwtmDQ
k6h7KQzo87X5eNEgk29YYDqymqjY7Hob4dkDFuuz4qdL+6lrexQiYec8nU7ey7l8
rbR7bby8lNBq93n2sfeD4iXSTeR2lPTLfTEuFVeM8IVf/SKCRkr0K81IhgjM+yNf
pmqNP3X9lBkifn1xHubRw0GZXjdW9IcQJbAg5yR2jF24Q9rustlkiRy3GEVq+m7P
1XBCpyDcMoEvIsQxQ5qCE5+Y/lsczMwf98evjFYRke+jKWtkeYeSzNsectdNbsJU
6X5YhqJA1r3/BVsmuwqRfe5RJCdTSA5EHrTC+AqCs/lg2kmkjkzkXTmyg3E7Sy1H
I7Aw3w/nLJICnTo400W/yylgtzQ/y0XeqebTbyLqCSrtqSj1DzzZcVdD7Z83crH2
gdhOD9Dp1ISgFLXH4azLCn5h9CZU9mad4Hop6Tigtw/PRyDZOSttCrNCDyd4+nMI
ZaVAaeFeDLiNLNO+BaUZAWQsh081vxtOb9i7R9AR05alfNewuF56kVA4dulR53Ab
kNG1exhMs5BfxXv4/mMvZOh24IFreo2bEbpPlZNPqFImpnbc6HUKTpNrGuh2isBg
H2kWcuwDngKD6IAqcAZqJ91MzcdF+/vmH934PX73WoQzopVFeUj8CRJPleEoL/Vc
h8szFtgpzp0Z0ohEW/ObKbE16TP6TUYRhxrwf57gCmdNO/mcQChUbebbkSp6CRSt
94jSHVVf6OIugrDmrE9bHiUgFPknVbS+F7nM+GoesNluQhXCrpHE9HN6kXnnaTR8
KWh9kRZXaq/kHOjIHr4CqqxtjH2vpbRYy0KgCArznkxzUnnGgagdSNHFBpAZl1Pe
WQNE0ri5vTDQBTk5CqXLDzh6z3rHSLWbywcqi3SOYyIlslaqih52W1CJPrFqm78E
MxJEkyogNOK2Qd1V9N6qSvrFhC19ft741qO39KAX40NS0MGTPItByUnvJwbT1yHs
qyvLJ1oM6Ltl/oCoJEh0vLh78XEJl/GUDXAsx4LcHIeU5+PZEq/La3HHaQxjb7J8
gH7JXClCOw9u9C71V44vZ+Uu/G+QB/xJ1kO3oKzt4b9ae2Xf/ARSgzfF+1/vqiHu
dR/zcU69Ahyk65Jft2nhQqg02n29XpJ7f/XBBo32XK49NjFL4vt6unqZN5GtM3yZ
nRUpwXAX4Nww9wr4kmzSArPgN+bWUBRtNFcQSH3N6oh8ji/H8icujE2edcVePbof
+r+TAe/diPITYC7nn/YoRQbO0gfZ6d3fYYZPE/BYwRZ6pq33aJOnbd8dyJqGPRyB
AK4byJW03AAghC4vc/2lvXZvB1ID2b7nFcOLjRNTmDzB0Vh6hoiOHMqqKNHCb5Qk
NWoSIsfQiDqmoe/qg3AYZNSFJtpMEwCAM5E9zwnfliJm6pS3FKqXdBELozHdU31o
+B+aLsZ4hErrKh2TQZj+o3A0q30MpNLziiotptwOep9A4rNShOF+ZqMPa7YOPZKN
Qif0KmeyTFyijDv7ASq1SeSLv4l4QljwozCfS0343gDypAM/VBohvpGDP5ACVsEZ
HattMlXzcQPvFJYUh1bS5+WZ4V+B3Tiqv0XDhel8YCkcbLlx4G27Eb3MqCfQtTS2
0qHMq1hfiGT5mYNeoxp0wngfpU/So0+ocJALAwpNm/NTb1s5gCfw13orzPIUK7Qn
Lz1W000oigqeUb9/vFWZyZM2UFrsQIifnR9y+WeEpI+yeOo4CsMEM36nC5qU2E8x
YmQDriaqfLOai5IEclthu5f1ZJQdugJd9TtIOZJK6r5bUKods5Q+Ne2zV1OVhZU1
/vltGkHalQ4VKzlZpB0R4ebdennuHkw/mlyE6e416kRhtGqLqKMjXYXCL0/He+BI
OYGi2HdvRSN1HbPcVKI1XHx+F2CP0/2D5BKURuIUeZHkrwS1+4Cx+kitLmKa3rfI
3+u/323WphWut93704SP3AoR5PBibJF6DThQ9m7yPwBzZASu+0HLr5phmTBL1qNs
Q172ESMU5wSwyuLQt1FKqLiBzyYzv8f8M1BCYS3jtDWkZLgDQw0JnAJGcfjwK+C8
vEWypQXS6nAqFHEVEhGl5VlqBBg3msRXp5wdyTYrXIZoHmLCqlG7YIDgscxU5lJd
V8HdDeJtwGc2AiRlBpKZ25fg+wwY5akXRnz0hKzcCLECdYihZaMBy+Q8dftOU9Oc
nO3D/dk4Iwe37YIYPVtOEv3b25ZpEx9oeR8BRuNmkEru0jvtV75t/tMRYIAkhevQ
WrZ8YcE0spHyjOU7/zAVapYWj6HjpVZ5vbg7DsJB3cuCQRswenjR2DpFExJCXEa8
sO61kUivCFR8TUms1alY92c21SIhDg9yq0APKPZhlTFEmaVRALFvQc/fCJ1LPm15
rWbjUwCBaa3n9QQhujMXTvieFLa+7j8vY8DWa5ro7OFzjtWW/OqbjEs1Oo6ntFri
KQYKAyy6XuuU7ubT0bXs/2L9ZMaOwgp22mRanoDeXlJgw5Xk0fuoFEbHrADL4SRl
coO/QhUkXC65+Ao/919Hv8dseEEulHcn80C7i1U2dIz/soP0EZGar9dzoyfgIOOq
tUrt5vqg3+fKOAQ/hCYuYWeDpArmXaBd8hqAeJ38RlsHVKzcpuETCAptbkvu+6e7
pCth7FglJTWmC8N2EyMzz+MgqGZOZpUyph5051aJ+A20Y854UBIfnmlo5vXZmHqm
H+oqqq4u14pbd1IBAzDnHktyNEYSDyp7mM5/BScoTRqOai5zelbqGH/n3493m7yh
uC9tB7beRgHFWAgBqPHO0YJSSbXiLlD8/Ik+OvuVOhZnlzyY65+hmgUkk4AFEhYg
rvsAry+QB1Z/Ku+2B6MUjsHaRmoxWNogDhmGG9jdzc/GAb9TFefympbxYJxtNTcK
6RIBEL31tEFIQ2EJqoVmtc4crJegKGJwC8tjlth93iyTSk7OgcgbYYIjXDixKy4c
aJYGAaKtefBZt3OeTa3hrWnHprQtULBRbmcxMEo7WO/amMSnFIhhK61WOHjUhLFQ
zNRFKtUfy/l4YauSF7LXDGnMCgfs8qKc127eXutIGovNAiEkmLBrtIunhBlOTvkI
HYb1dmdmCMCutOBjqDOkzOd5PImil1xUvxK0x9kThQomNEn8130TFpN+Schf9QVF
/4WJcpTaQX2y0ymXREI5RmD+GFcgJt1SYZDuYSvW3xP2OX5BABIg4IWA+HzG+rsQ
Vj29ZGZnwx280R+TCy11zYv4NTJx35gi6CulkvFU1OWRkyUG5RNDQKkMZVycTwB2
Qgar4qdELYWbEHzjFVWhgJ7UdPIWIHC/ic9OlIiRYcasp+eEkW48JKIoGQtJCFgk
CQzd5EOFNl/2AsriPYZj0VwQruuAqtb2/4wGSbkVl+5rDr2AxRhouicK7w4kmQdl
Fs38LWz1+vgI7FeX8hTSpi0GAB2GtVZs8hgL6RqwCQorcl9qAwzerNjcuqMoYXS8
qQBgdmm8NvvEcvN1dJZ0zqRabBEEcQ1wyxqAJBzAfKlA1D1FS3F3PaE7kDNOUnoN
+0mg7PmumKaoDNXtjuuMMuB6hvaX2/bhiV5ZuRNcjjiJj8yFc7JLBrcwDdH2+xwz
aLxSci3LPCsitrgkF6VR3L3gJCziFb1bAJnuvmcIY3cGrMnELB8bpyRKsUnWqPuk
KXW38hc/EEVOLJ2k/+OV3Kt8qR7T9LUMHuNhcTH/G9H6EEHm1aFza2vk/0c+WPdl
XLbzS5GqzaQFVfeR+aStHW4Obr2l6lNsERMPycl1L9brKEjkbH+bWBFpQK3TATu2
Pj+ubF06B5/O2W+7jvTOzChkC6oViLewuhHUrS4fpfRwLoOod/RJh/TpnEXHpNOG
zld1x8RFs1DXzxRLt7x8PLM15qTBR1sTidKjTj+L6HL2BjeOQyKoKq1FZrCWrnVB
fHchMYOpUXc9cQADnWAMDzHAsCF56Ev+9EMOU6lBw0PSMJJ+Wp2i/1dY1X35ptLH
2L7gUU6U5isgXohbkQ9++itP1cb8aZy/hs/yPhUBQqaAz6mE85icE8X/T8SvZHC5
FMy7Wn9yYyGb+2D1ZT1lNMctcaKNCFbUOsRGbwwf/4sIjPAVcquXSEo7uwExVfJz
WpYAQFkeTCx3yKjb8D8ciQqE3ydYCm2fm5t/JL/56wI4sCHwjYVhE7zmLTObUxKx
ixGeHEPHLrkP2jRaj2xPsk7LYnCC+fucq9gUff04581VTJk+UvDhAjgaJgZaGs93
HLPr/TPdI9LJbMCwTONy4Bh3UjPH2aqR57nv7Q1Icyhl/ZeRPO4Pz6EQZk1IClNc
CQmweHyx3U/E89smeWLfZZkR6oD97gFQI+0EnybhImOL5h6AHK6Xl09OQR7Cu1k+
klhzgkc5TIXzReIiuPBzpT/q0vl/T1zUMP5kniHhl6EY6MLjkGwtHXmh2Ijdvqmi
m707KjYTlbApc6QksUGWJwGWF0tyaGoZrgS3R1VsXVRZSNY4YBiKBjL3vM0KpNjO
INF0WJlluwB29YXtb062EYd7Jt/FmeUBKESOCTk2CJpVI+0kEY6HSFfLIlq/zpGD
pp1KSgRdsry5inxWu6xK3HfAq336cX7dCger3mkN2Dha01//qtxh0NaROgfCDb6O
eJfBk4t0eUKIjnTB9z7NNd+UjNkq/owsqe5EeI7KttKiBzRBjzpsYdzg/UR17bgX
xYDZp4ph4C13740hsTn8CTIZkYDptwPjTkdDBMAV9giLUstIcpHrFh7LtgyGT+c6
5IwIOh2tXdQJi2WVqiWsit3Q9qdgL6e6SB15RBATGkBQgy45GVST8x8tZA//fWOQ
Pu5lS1uAIFhRtqtT85VYmEJI8YamugT1B0lT5I1xQoAIG2V4Yws2rfXvIcwxpcLx
1c0n65f4gQFDjiwUfLVPpMZ8NI6xtMYB64NB/ZhBUye5vg7FTbZ7lpKSgdwzmCKX
iuIJUSIELZJrM7iUs1gIV2RcoHO/QweU1RIrb2IpeLy38lfswWeCVr6Jp0VYOq8I
0PuouK2f2jaOfJfcu36n1agIyGdrP/cdXywW4LvJM09Z0nhj24Fd86xOq6D0XGX6
bFeWkmp2MSx/l4rvS+TuOf7F0lqPRSWjgPkRyqAPdh7L3kdphHNNz9YCYLQxweQD
ALaWvKGWost4GQ4trAO0jHkA057//atPL1IRpXAVWLA/DDKlCYF3urdaw+vLRJx/
ypK9+8SpjE3NRp41b6Gi8NjJxDf0W1f8khH/MVok0fxVdkrFY/0JiSCavdNmKmdF
G1Cspfl1fw/hD2OQBFBK7rcPkuDnUmOSfTUcnoYCT53wU/JeNNVCrOTBxtOKIQ97
gSRI1D0hH7yfNPYpUYPbfHzZDMTXmq3sLtbRpdGCZmXtLs2RUdd1gXxdFqO4HkVW
USeG0/7Q7g8iP9/9B447c1zeJC/OaGrOXnocpiT7g5AGPnZ4QEDgFojwxcEM/8+Z
yOS0Kj2UmH6l2lK9kQibgPJoCAYpqtGqrgRTfmDHnS+HibmXG2MDABpuV3z7Mjv/
N2W7rFOAtGP61hDKoan0it8C68FzrG5PHJ4RXmscy4uNnZ1t93S74+UsBvAiQYjh
sym2nUZZPg0yorkKJ46jSFdvwrsNFrHBBYJZLxLHH6tcWnq6zTF+Gcg6L6MtGnqB
uT4h0biZMwz6cg7/ZYb17LwU48g5/eoPh6B208YrzbugaNJ670i5wtz8aRUAEaWP
nmqu2F93whl1NFxbi3E5VWaVySifXnUdtiRpOlTPxCtoCv9LLwmLZ/VNsOtKRe2d
uKzg5KVZGYksPiyCnU7uFermRXX7UHkuNmn6MPLlU8X3f+b8Njme5Md0vka8IG/y
EVCE6683pRRYFTTFsP5eEOsvWmpolQX4TtYog5lCENQeX2nrj8EA3zrl87Pqu2Uk
RVX11DmG7zopbW2GPZ8bDdLyGvpWrsqBEv11YAyyEMSGHCHZ88zAWRxAD3IxMrlJ
e2k7yNcJuybES3CjB7QTRi7VUp8bq/Er+9R5NFepbqaeQP44ZOHp4/LuPfLuODhz
HWp/1+0OvL1IZ8Nf1VTIK0RKJsawj4T61bEzZqCHksb6XFsBkwi/Mm1ZB1T0dAh4
NHs+rm5tikEwyCrpJfEhjEkA1gqaVPPdhuN+D16JIc6G26oLJLbg1kqbDvcv2qhH
YE2Wv6Iy0hgkQ+ouy6OHuEQ/SutyEo+l9vco5xeryhRDNaJ1gJPsBeTE6PCEkce4
3G4bOS58BVIY2+vJeiYyh95vXmMzZGzQNIP9U0WeetzKuVQ2xajXj9pWtvOmTQ8r
G/UC+58CQzM11on+nhogdQ2ixmvTu1nXmzwb9XgZCYzleydSgM3JX+ECauY9LILj
GGGzu4pxT/7TvhLH333UVQ40GmwIn2AXJxqPjecjwifPrMrD4BWALEQdE/ldjwwP
dX6nSkGiIshtUjfJRG9oStCUBRVO6eQHxiggTO4N9fdaw97Puq4L/oJI7p1JyM0E
h6wnWNnuipXvcmrHA0Ich1XpjuOS7rC7IzgPuT7TqzUAh3SjkC3nsYwkAx7nVqgs
EW5VJxltQU3SyJiERAwcAF3dARQfsQr1aNQvykmGvvcRK55Gd37OJUcz8tVl5o9E
V/t6rg7/wZHbQWEJ7ql6R2KSaB/WKs0wHaf9NQszG2NGFn4a1GbOrJu/xzs6t3ei
irWF/9CdIDbRPouBAsye92DCyCwuDHBpKcqTdaRoU9aOaLSY8xoO8Ou+XxzLSOiE
scN7z5yWiahXnmL4O9sBBrQCOpxEfYImVGWtEXK9vYEoJGbLVXqHC7orGL2Xb/2Q
pkRdaakFqowzZrpCj+jdjnAov9/8+DMOO5MJXwDlrha5XsWO0iqEtsUOywB9G3+H
DbZM4702LZp0Lt+XoGquNKt38S+n3wsllr00h5irss0+EBiOR7R6Dq+8UdmpTkqD
IiV/WjmRUYIcA8w0NirK+leFSWtrjtOzy0F52qqeHy1X8VIrkgy048JfzgwRJcJP
EFfpS+l0IKyHGs9B0+FotndpdFF0IloBGn85hitp6Azf2OoqQvftTUxzeUh1ZHI2
92FelAtQxBgBHdYsq1SfR7xM4vAkLQbteKzsqE5+AUMNZ0o2quy0lu8ogHvkUfYz
o4LA/pQbrOgSH3NfYYA3J04YGEGJL0op9/7bg+JOX25xtJK974xpcJo2k0vr2CS/
azzGmI2r6yV1KjFcEA9TAnJjnZ0w+XzwvPfsOrI03gXX76LLRnO16Q4BiXPIvKPA
TOWRI17Er/f32xSQGF11uZDl8L8jxTtgT+32gpIWbfm4UKDDudhnvxnsAdr1oNEt
sLV+fdK0D3dUjdKBBT48KBjwFuGffWDZw6CaRKsHcvp+XdzpJKhRKZD6URuHneUx
WSncCuSYM937XmawIGS3MVDcFSo9Lw6Hq8n27rBSb1DyvtPo27ut2YMvN5c/Er+N
j99oc2Qihk9GRxbnDzfwuXcFW3fWIOyzwij1mVK8kCjZKroMjPgKDOhYxpytKV4J
RyPF2rpi1t2jQ4kyURqvPv/GtblYrX9vPRPqwvlsUvp7gFSzcgFbp4OTOLzdvylB
GOgLdhQlmlbKdSyVvWGZxHmkVgdBVz/fCaXf7kmU7dpDxknssV4dIXNqf3qmoyPh
hizOTQ6mUwdqSm0jtcVXzzgxzcH3ok2dFTt75F/gNPU6aeYtIgjroBK1jRpk6uPC
wmRDNbi2u42L0NxVeNp+vT2AAEcYdnIB4LbJMtxKPMnUsZF3F3vf2cOWRN3h7e/Q
iN6qOEA5F6UYxUFWIgOWzyHKi945ddvOPj4ZLopQ+xPplpR88LURLDi3b80UGxRU
b9R1cnFFkvZLvC3RIc37tIofXw029vc37ES4IeWHnM++wD/AIfCIZqF0nY0RO0L2
G6ajPuJ1OkqP3BlFaxX2jDwpGe7RcuDK/qmrlNzBY0MJXVYvDAtXDiKzgzD00UxM
y5pnObtbayqjoeoy45SmFuD3IleAWiI1XncPutDeGP8iLNNaLnF3pqxk11jneQvP
6wdeS+eyxwdDVDKQ7DQxOhbUZ/jHgMY3j/QBCBbxa/bM1z935AwhxKjs9aKVb27S
POjcskrrU+ia6HdkEsZ0AMldOJAJtOjoMQhvbgxPr6zgpuialPA/KcZmUKIaIlRK
wM5V3D73L+6iBbTOII19OBtQluao5jSdHnvvlRoc8Tc9OX/+ZgZ+kC50eBU9bcnN
rfdr7mV7JiUKrzIgpi/au/WVk9Hs//CieqGVRox7EeUpj40vMckRrQ7cHiP4Xb1L
dSobpPQwgD8VYTsfYfu4izcIgZgdHbSx1z+U/KMkbLKaeBeUvIIfCvCukIYKLrvk
qZDY3ekRWZl/rW94fGp6StaUHmCy+aI2muRCiMMCtvUWX1J4d9jHqy1/oq6ms69y
U81cXBQp9iy5viWPBGkHLuiWDhiPxGX4wZdx/ViDDEch/7dxx1rRtOuP9rAXPicm
c2CrkCt0ASTrjkI9lQF2ecde2pFDdat8DrPE2Zw/ItTvpjUz9rbARxxY9WV3gXg+
Y+yQ0RkAR19yQh2mFtEO3SPY5wP/pfzDiVBmTbPT9YKAXzXh6D4I3W9E5845+fID
vLd2//3JAUOIRmn+Pw+ckhIA7zb72WdEtJVIGXJ6kD+jSJhZsJEcE5nnOArtXbHf
28qozinD5D2inITNL3ciwv7rhX3vYyGJzJyJzIlZWR96npNvhQcHojQu6yHCxqAj
Xq5APx0hCjfrntJJp1dzv0We9cRno4I5vURkrmsQNF7f0i9n55LJWBTkRe30gCQS
QWIAsPSPKs7+kRgcZc/cSaa7+43LPk8hQ3QwbKHNFXKWl2HuwtlTb7xbJr22ylCB
ZV26u199h2R/e7o3POAfU/J5jY2e+/+e0us4eZ/F7vL7wxfaiLqipKbpm+D1PuaW
t73N1nle2ota0cmjtw1r4PuHnReeo9sPNHP9SrA3qvmxPHtavEo2tCzUrCCiyJlJ
oQ1evSw2sBXG0/x/L3WOwFHNHeRXcHP5F9PLgGX1byGH01wcQJ3J509XreDLvixn
8Jux4iw15i2mGeJc72bw/raSUaqllMO/gpVTjWnv+uZ11U20ixSNPX3FghKa65h1
pV/3DotePyEZgKwso4a+63sM0OAvcyPlyk2Cymj4ijVxFltqPIvDy8p1+EK681Cv
89ItBb/54g1fdO6N9Nebu57HkK9tw180RbOSr46xK/2Xw9H/rwnVKCYnx7Kdtc6A
JNaqvz8vI2OfEcP5scxytH6GVlo6W4psv233UBDjJkytHlSMrL2RX01wVC9Qiv2j
HkR0Vt0ogDHI5qKkKG5DqoyIWtXmQG7dkGLC7lfEASUnt0o397p65UXbwClS+wjc
HgayPEY99KOnL/+lT+YQKlRiTUZ75eRd88mnQyesKla8V2MAK6mDgws2oZpiL5P9
A3217uSzaPGx8a2FBRgHDzXcMdH7LmOS1p9YtNkECGyQXVt5j421Pkwkvj/Nm6R5
hdcxrevxtD9562/JipfoeBdelrYDt7K8nEmobp3yhuutM86z7/doXLpznOXY7BTQ
GlA3q4Iz32H5LY/chsurMVyeVii61Lavcbs1cNkNLHPmsQ4ggbFuGa7dGpWekl6y
N2yIjN4kvb0SaFA5h/Uh+aBU8YrDi2tAJNfHPdW8YYLfsqobyTA/JGejpK3fcnIX
JCIu4L4M1CiEhkVnOvzfrdtHfuIZMw4RnA/kXzE50ZEieasUFB4FaTc9fI4DPgsF
KN7rRMYQg7Q3eO2Ab2dhT/XN1rpfLW3kIP+eWp9ti578JlRh4xXtp65B1tbdy3Nh
S3g6k1HHvAQBRy8/xyTJqZp+J+C2q1PsHXrnNox6yV1Z6kgslwddL/JqrfBwYyMc
QtE8LwGf3gJdFIg9R3uTNSa7mtdnJmn//ZXgEsTcqmA8AfcP45UPt/RIHSuBh5/F
1PTGotUCEtUjnaqi8dExMfBuVZFNeks+O8jPuWJOJD9Nk8s5vF4vnQO9ogr2ufgL
1GkpBoKM9ueSFJ5scZPJzwXSNF9YBQ/RmA0DVo2YfrlMF1N9m7Y4vIIIo7xDQ1yw
/b/OFC/LnySIBYZ+/+9VCg76JSA+je6REHsJVTVS/pXOT7EhXCGouRq7GJSt5FRe
xUo3TqeGspZmw1E446jL7YbIxmkVxkDZyGzqdpdba3yGXCKHE7l3NWOyWxh9+U1M
uV8Q3+DtJpysz3L7MjmCTjnZrERsDmJjfEYVhEL/H1y5rmF1l3q9/x5uhwRzIic5
eZ3C7rOrlbrIAo8nCAwOryPWLedkRcjygsdCmrG+AShgwOvco6ZF9XzrwopcB6ls
nhfRjx2qjkEzw9RVdbnl9TmhBOXQzd/uNzoj2yFxDlyEBMFcX5uJYPthwdt7X0uO
9sjnvYPY7vdFi+LhoIWwqY3lZiWjpG+93J9ueXMkuyrGKW+PzlrvBX4i27qoO0jA
ODWgi4KDj7G4hw8fIUMltEUTjXBiflNUnM6Y2V5vgCUMh5vGrRzSuvyLQFO8PGVt
19rNBN1Yqal+xT1hfq7tWvYWUhs2P5SklNL67XGTaRdKHWUvMKp8AZogjIMT+Mma
rjmoRSjvRr8Rcv+6QPCs3SFZOk5uS7ruKIC+iWNWLkYTiG+gnxc0mduxD+NUbovi
a+uozbhGCp2IazlQEomYwxkm/l8JS8gHeofSKFm4dlNcMR4v4REn93qdWZSKYkPR
z9IekXSgX7Aerx4O5MTxILYK8BAELao7I7FG56IinUzbagxYbuBxj16HX+6OtLvB
38I9iypYdJ9l0l+CTWR3FIAAwB47AwWbIGrvgx14KGPaZqSPnh+X4A3y6QyV/I5V
SF5efj0ptHN16TF58vg8d86QKabunyyKCo+j13IapeOyuff1WM97KL92AYdweg44
6tsq+oSILXeOwQec9SUt8N6ktH8ZFykusIxh+DJg+t6rTG6SEqszM0Wq8T/HkRS6
U6ll8vf2ZoS08PcJN3F0kI8o6tacWkiNEHZ1viw1SqOE2iKDRWRDf+exXD1zeTSY
hghjHrAjFFIK8dsroceVPPJr5aAbPdG6l67ffFlTzbxn4DNKT3EKd0PUuLDJ59FX
B7mdhV6AP0Uj3HtiI7qTI7vyHCjyRjcZxYuvpXpnNf1Yg62XQZjI82KmhYNr3msZ
U0sF0x315gubDMpO6KyXaD/CC+2Q9jHxfEiGgC4ueSeU437qakE5+YlK9AE7tjtx
n1FUFtzKLNRTp/qXAeJBAo/A24YcBn2GY1jOb/vVwSeWHcg/+DVHpSuaN0XXE9yJ
FDJydrHsRz2mCPf+pOPpsbTyzz1Xwgydab+gcGVeMGojEspUWDKODh08JdnNKxix
ouhAsk13bnbOqfr2mwzCnmFAIOl5wplr3MKWTHSkiGZIHwsoFMhbdqvtwHCKoWcz
k6ZEEgkZhCPTk/VeigxixeHKoIgQRnJwW3hMiXQXFqZuLozdBbV46E/9PX1CRlhQ
sKYTQJBd60+8tJ9VbddUZp8mmr/8bOVrEMNTxosRhVQEb7VazwGakQeYv9Rqu8DQ
Yk04DIWgJjxN9HgbEflhO6dLYa1J/6otzaAAwO3qKMZeHjvnne9povrF+zrjvouK
MgWnNeomhmkC4RMtWvF3gfDa5CoCdkJLiU7EE3EKAFHXSonA0UahqVref57u1N7o
rONWAImkvb7tMvEbuG4ngLNZRJsObXhu5DPQ16386zUkwjjWrC63k7rnP/UL7frq
XxVPBs8hvgLcSF+gSd/LrMuYCTEmxAy9MCZwCuOsdgftm8jO+07PJa6jf52li+X7
z9+85+A/usdTVROXMUqYnrecI4tE/7eRoKLN+gmAijF8U/sJCfJTxeJXnOUTQJoM
Zgq1w86SzKHTPavhm1NlXyRONOzzjjtvHOB8sPV81vTWYvKIIsPEN5r48HEJZ1el
7IstmAgZCxzuenVmP+qLPUE8igQWTKNKINdmMWphe1ZGzkYc5AhPg+tRtWw7kP+3
mfObNLqZWANMAUrxefH1e1PdMcBFYchdBCivKFSjNIYvYioSUh4XE7jGFbtYz05M
LmUYVqAXn+dRZjY/LmkfCWuTvDKderzH/9P9yFTt4VodRdvt3D4TCddlOsHw3KjV
gyAZAkThgsb2N1VKsiLp9WIGz+4tHoRNt7n92kN/3l9Tc6G0Try3PCq9Qd33Wc/e
NnfsDFdKmnb3ACwfK69c7Y4hkD9l2+pDcYBAfxVMkukUE+od6cJSFPPcQWD4HOX3
SHOi9qRsjFWD7s+dNXegonqEfaljZwDNQ3bnY6rdj356epr1Bg6icMlXO5ZPhn/R
SPcebpPxiDPs02FaLMoNjiiFSajs+U4xWaW3aC/Y5dENAuVvAnN+591z3sFXcGww
WbXD3bQSa9Lp4HSz/J56gTCFGydxM3EwPU8Oo1XRFlXn4cSPSiBrjRsjb/FfX2Xj
SkAzxPWGTOG3OZCSFn94Ag5uK1jq7+xo8x58BlgZ02hPdgOOxgsBVUMnjSsXEpe2
B9SJ8xqg7aZFLhIllvaH9ayitzEjLcdt+qRfUZiifS4an1yEdAkUDmBX5kHRISma
ix7pA0NniDA/MBGTqD3t7lAD/HVZLd6o3PYHGNt2EwvHJsPH60jxzYuiBD5m/eKE
Bh79xpmi3gCTaObs5U3dXdYQib70dQsVTriKAQ/svogtTjgLhiJIltNQq+1zCf8x
UlsCxVDINET0bUxhuI3skCVCFnB+hVYsGQWPRwTXDsnUvRCv73mRe6Tv8fC1FZQM
bp48NsctZ5aNATJWLmAzs6ED1NPsfX8mVcHlkevJWmsEX/eTdcegRUVyd8RYWOd0
vJAd6+/2arvD0lLiR47sTpg6xOhIBdcomvLsBABk6kkN0tbjzT0arIcnWg69ysav
88lqzlzAjA5fMIHgz9Ui5oAijhCwWiFiUF0Uo6up5Bxleo7zAi6XBv3YYLv65mQk
VNEzCEWjRbJR3ObJ/AY/K0J3ehMOzIllKQGbDet17Z97xxPBSi8c+M2KSJ3qPjUk
EMy/gE5IQcAoRn6Q+ntJ5GkmXdJo4A4kNCrEKo5YwCGm4iTaIRyZGNtxBYKwHW9N
BsjZRMXMJ2+qIhkeUQ5g3p1vWFyguHqMF7226q0E7vSKhxEMF9+7hdM2UFgIZjdH
+kTSi4TlBVXtIS1t/Q/tQ/kt4wPyKh5fEPwa7H99jN90Pwvx7sDivsoIDXaMV18w
08W4JZA1TAe5SCREVDqwzDgkfUX3Z1Cf5id0IBfLycMHFhKUWS+08GQ1eX/QABz8
bUk/Hfnq7CVhmW7ruY84FpqapnR+32wSmt1V2cPxL9vxKO0hLajm+tzJWWWOzF3l
CHYM3IpIgfhYI2IkaNUISzkcaG1IMi9EknJ0XvauyIUGlxoEPLYkp+gr/CaVMVYS
IuIBL0LCxUzqrw+0yPJG3YjK8BaZk0DLQMeWJIfYx4dJLXTvS6tAkM3xWR7lzUIQ
L9VKpafiXMSwUTbqzfQDEaEbvnLa+8GD2Mm1SPZRFhJhyi3pLrDHXYqILh1/qydM
9D7IlVSkZWdViOHy4gvzaUYjSQ9sspPgDu7Rga2oIGXJGOwJ5Oo4TLnvAhTrUcrP
rIjF42Qz0YEetdEFvFNQSUH9CdYfw5kaqzmqryA95ZKiaIhq/sxFFx8t1yv3QF+7
RBkFUtKSc4qMirjpx5uWyLUCfLkk4nMy3Ho/UD0HVwdfGstpphR7NZGg5NyZqx+A
oBPX0RSaBPtLBkoAXe4/T93nplkYYdelnejKMjP8dOr9V4PqtLCb3weFSCPR3u6H
n+58+BLdVqnn0aDqmGp6cZsUGjEi6W+naQ09AMvTUK2y8OfPZuQx1/RlKMA+GosC
/vHTovTFygfLpVxoJv5oP8P5x6hLvMsQpYSJ7fSgTQTnrTHRjSGx9paDVX0dXl+Y
UcQNlWKgERZDkoeWblFasEFjVBl2lsTwkr6pXpanAnAk9L+OZLOYUa8TYXVtlFm3
gswnOAkHKeCjDYuKnfNTfoCj67o4NhbhPvDtR2zXzSS7pbruEq+esYd9zrS/UBT7
QFbIavc6eC27umb0uA9+WS6ejGIAf0hKT1/BPB0RLGhndyCvfBedKzydX8DCLSDO
CLlfBrbGaD7kndQqfjzeKzHosUUuPxI41ty2JUaD3dCNG8QFIqKjUM/okjVktV2d
sg9zCloaYinU1jKrQnb8F2DjkhIVi4fANIWmk3znSHBYS65N8+AzFFgev9q5RA4j
pK+efDbCz7/PyC0/5HsBtGzmarftqcdmZ+br0mu2XbDQBT8q+RcYJiN2kevDME2u
i0wXQ+Pf3a+y62lnIDSOzsG6+whvuDWP78msGrMxsdNRjy4RcS9sD4DMqpnV5tog
PZYlBOo5ruR0PZEzyAc9vuXsfEN0XBUVX+8wObEfC7gJ7qwENFmOnJqTGhBu5ujW
fuIyyBE7D6L0RQSpyKe8vqQf4r/tGgCOSTW9I16eBPB8zPFFugaVZmlC918eNqK6
Rjf7P3BwuDwvUuGnM3yJ3yjLHYlcESQdxoH4H6+b+oyRZ3hK1fWpVnWfYkHhWl+U
773Z/rzxczHTahhZ4b9eLEAsJtirYnT22QO3a6pE3icsfF0LUOEztO9BsmjS6uA/
AV94WiF68r/1K/F/iBg4uQkZjMSQG5REk9lxiVqLLjHt1zXRcGQN3bWYYWU8l9Yp
b0MvpQzaIp40vfcJBEOq4dGZdfzwNChe5scXDNcdL1bSvi75YQ8gQLRzfhhwn/cM
tYkFLq+cFwZSCglroYcqkQIjGOrEvh284gxUAfZZeWX7JjZKBVCzk3TieL5geIRm
4Mhcth9l5QGZr/EFxx782XzSZFDBip+acxc4GMBzXM3td6e3gUI/1lRsXTW18BPe
K+UNhAuu10ZLP6blAN7rhrq6amgKYZjE0wmjWQcdGvUy99SJ1Ogsu6abflLLgG0m
KozxgmE4neoeW9mDtWkfbjSuY0AEr7g5K3ibHcUxIrWlYLQ7HdsuM5DJHIRawvdu
UpDI//umAb3AgGWziKRggm23SBDA58ryZ+w6RwRTc51db7mJpP6pF224AcTEw4xB
snvPsyusdQ4FkFlaXfoItkXz3qXoqynQGEBlsSFvYwI1PDocZ30kI2HyH7J+HYW1
yK4+eDkQk/zvKyhI+8ac++ufUJo3StRU4q/9Nn5DdwFnbITXbECuozRhu2NM4vFR
itryqFmXNzB1fg4EY248xyv0uM2oOm04u2I/kcXasQZg9zG9iLAjn6/4JAVnD+Hi
/z40FC1WZoHJvwxKGPVLH9dtu8aBD7SfFbmIot94F6yRM4BWUxCZPSWexyQRPRUh
YxRNlT+//oo8QdEPzJFz5vRyZJZWUgmGHzw9X7BbaczKNYHl4R8hSnflt/l2PFKP
z7JenDv0SsiaW1O2Qj4oktb76Wpv3hkHbOA3d75iPzFy9wS5REaHVQXYXdyZNAtZ
136+2f6+327fzhjG00cjVYL9nWRy8CXIuKPMSQ1UKwB3SS/uXnQqyOwDa4ziDBp4
Kp/t56mAMplewYnZOkdvORdWQB12e/I5mecPMluol4HXpnxY+THeI6HsJXgdGf3J
9XFc/ncWqk5wSrzR3/xXHpmHtpWnzkbvY5xR2rfKs5NqFxDA/FTvqmikdqI09lc6
kUu9SOty3HrOHmHrnSJ+kO1EX7n07EY7PdwAhdH3J29bb1V2xJKJNGm642/xLn0e
adds1bdFTnM8sGBVvqe6WpxGoXLslNQ/xdtkOEktSRWthVpYZNRKOQz9JkFnfSBd
/tiV6imt4f4JHGAPPaJf/vhqkgnS2QTAzxm9yXPWQzEiz8+xDZx8rpIoE5oKZoSN
taLXmSRXgkwsw0BTu7MsIie90IRZVINbC9uMaQDk+o8zAY5ElUc4mx7IOVX4qcKN
uIHXmZLxpFQie16TJcth9ZtAj94V6ghVwHvSLz8ZL3IW8IkPM+yl9YZ3nTi/4SUU
3zOYyrtijy85qYaxg2yYPCyy4/gaZS7/56/lAeWWqfZQfANU8fpnvx8LVkobHbDW
qbnaw+OWAurkyR6awdMc3+qvf6nSBFb0fI7/ooYIAxBfSmg8IxXEA7LfERMfW0UT
ddIAnpQuLTxuN4w1sVSQslSp/NBlPOMNphfEmaqYe5pdSS5hTRpGQdOHcCNZg2f7
FS6ZkMUZUYC4xrHW3w+aotu2qaTqIs1jGy9gsoeYXLtpwKPijRvaTC41p+YRM1Bg
v4/EAXURiNoMV3KGlgKn1zPeIOSBZpeYKG+jXBDld+gG+TcByS11sZ7VO0y0mHQq
XMunam47XrT+I/wpDVWnmCHe7DjXhBY4F5piGRDhfHssFzvL/PtqHjwQ5FEkhYMr
nNwWS5oCNze9IxeJaRGf01OmF64M4XDnnZTtM54WUMYUo80zOdNvSYxCIvYhegoz
2Jh5mVXkLYqLhDWrS1cV/tpevPlK336xujM1cxzwJRxEPlV7yU56OAalwCsn7it1
NALLGRzUBYcPMKsQ5nB4JBmCdAEz/0T7i5oHULKweJPG7Ao3FqkkPJCDc/FQp/Cy
R33EMSvpI9VaLk8SC0BFRQejFYTw3y5EcC546yoGHDZsMZet0GUqO4QHUNWXzs2s
k7PPY2GUfdCbROo8Se2hgZN6igmqp2JN/oCjUeesE3DpcUQpoaZL2QWX1jxXookR
8d5EHiVs78Rh5XCkzsrmL2ndqfYtd05R4Na4cWS3WehK6qZ6wXK33QcFyskS5ohH
uJIu3vVlkFU7AwQmHqq6sDmIG+/8NT3bxQGQs/UpIRNSV6KaaALc6eDe3ujstqql
h49aAmDSJ1M/z5yUau9BdSnnIDDsVXArc0UiOM2h4jDAACLuezdL9Ew5PScqai3N
knRVHbEN4DGO53uxRjXuCjie4ilaq7NUvG2/Pe9L3vBTcSGfX+Ti6G2GTEgzBmO+
7DegLFTanaUkjBD2PoJIvvLjViGgLqO0qiB/uHLnQtTrIU2xrNMgfU6KCyu3nCOZ
ia5fUHOVZJ9nZgyh1RgHRPCieha19ZDvv0nrPFFThzqeypgsx+DUiTI3pWddFJty
Lb4CyLV67D/dm2DIziJjBrrTqCI7I98UNfE4F9iZvjYS6aDBLCBBF7IJT4K03RSn
h3WY7d/rH6wYJpNwR5ftbCyVKSgmUVnNcppa45SVaXGixYVbu1Q1IamSnWpIviUg
sRoGs48/ei6o7OIhS930Yn+8bkm3eK30d/9sQS8MS28UEoSSehY6wbD73rzKMwbX
8+mZ8lUJHNqVS53r5meCyvCDKNh6wHl+VvLFLO1R2cUDLNXoBUD/+9sNZwD/Iloh
1nhR69VsQd+wWe++ymfoNeBPf0aCvGuHIegE+xNb3yJ5bj8XrmiqcFIw921LnG0E
u8hlHX57UvXPX39Sa8O1CFk65XqnTVcWwATMvHTkr1S0hTBMP5V5e4u8owaW2LkW
54JEVmL8v3GlN+M3nwjO3l/91Fb3dLTJ3GoEOQWQ/+UxQXqZdSnrkNz+P88NygsH
rX3ayeFQFooARbmPyyPgS99YDl0YCZAzGYKd3o+BY8Tk4DNtXIRRxGLbqEPsnD9M
4CF04/OTF7KV1ZADb/9iz/ZUjJuwJUs3RpIvAd4R2mttevFStbsIaKUgU3HlGbEP
YA+/vmQcqOlkWvGeGaqQ1XZ01fnT40ZnkwCTWexpSeY3ESi6ECl7WhXmk/t2t+vn
9EFDpbq0dKCBcX4mZlSEYVLCuBGkNvM0qTZRtkhaFa5UB8VCSj3q4X27m70xiY4Y
UI/E0wkQAsAGUV64s3LfP2J54biV0LzlKI1DiwUpDUiZsZeC5PLCqknM5Fc8fDj9
px6UrnEoWmq9h3XD3NejeUP/Uzj119kpAiQblKas4bG0Hm/kGZsCYosCi2AGDfqH
I2KmIkzKxElEKg84mWOBBicjUA/78ymXEybf4l7WLkB0awbsSlQS5LZu/utu0gPm
tCLweLOuSY1p/1K9r9O/N4WWbQ5td0442cGem/wBx7SX5vazXK8llaioUdB0c84f
hHKTixPA05JONbjLbcVpb/Eeiqr5mbgW2bljvXRaTT3oDWDwo1/gVXhf5vyvk2H5
nLTxbwvq2M9DT6tE68nD3Mc7ngmTAFKgFdOk4gXRyAuvEw7CJMdmhA3mnE4XvS5Q
NnXLqxBXiR7lhUuNQyi/1eBmf2NHTnCW2CB8HSMzvq2mHLZFIQDfn8P3pSDpca9/
cFXaOhU8Rz3iIRpRDxhXdgBp3P7SLgk8mUnWfLqQyEe6KbvS69+P+9TfzNswoNkT
dwuHT3NeXoA80NjAAmeUexUV484Rg7SNdafpT5NDIoRkO/sXYFdmanreoCbROo6X
35Onav/0+jfNlnN8oy7wcssNIkKL/1RtRjuiKLz6isL1sdt5F4pFTAQT6Ko7I2kD
2THD7erQIGlY2UD3egSOQcs7KQhEKmDcJFOE4rnLjFZ9AZdmIUnuPrWqnUYW7ZN3
DRR3M2czKfJ8nSd1nH5DAa/l5Yh2yd5+YjA1P1gYwU/lCPtrCBxaiwj4tPXSMqM9
uodtnF+Cxv/Zp3y8rgPvDYwt591UfhvXEJu8ap3xG7imK223xa1SPQrtkuuW8y+N
47o5arG7b8Sg//u27TYgX576sMs57K9dDdafbYG+eQsfNB+LEi8Yfx10Qnby5sjU
szD/WZKmQ6KyifaPuo57RiNwbDMI+kBooz3UPMN3sNCBdH789V83df0nTGM224Yn
TRkW5+7Pxb3BrueIo5rFqqPPayorvBaPGtR8Zt+iVcMFr08vNaixX+IGOJxDHe/a
Gwns8aU3My1VpDpKyWiLWRZlsTzFO/ovC6nqpHTy4+xxP5jwiYigB6Zo2RLNcNwi
pF8tIBUNiqhFL6kUS3+xfSTiz6YooWxghTfU91E+6dePPgH2oEGcaI2U+806M9Vx
NYySfg5SJ8k2cbJwvFU4fjY1FiFRl45xN4B8LaRcKaG8qrGvH6Rgk5WJLU/GpYV2
mTtFmZi5rgkxhj3t/pUwE/9OWQjuJYb8jHsZrIZlxi2YywxRo5Qb2B8ChmnZ38Pg
fRQRtPa11DUSzPLgpmTWhGY3pDvPQ4PxcWYGcXYKPBjC+Z0ohIcJAp3XSiIoChWa
d6q5zIbVcnuidSBGaRdpzWFqhla8F0G+qW+D/gl2GV5eTJtSIY0H5v5wFTa0wbLJ
HFTpZT+IAXZdyXyWa+qh/l8zqkuanrDkwUAQolistCElSYUVxdpBd5bl7LNHtigi
IZPWcg2SqLiLMJSU92ono2K1gWXm0obFOWmOziqPvBoJURiA3coK7HCPoyBXlvzU
s192n/xb71Mxy4mIYaFnecQESkoLqL1PgXLXv+AJz/vVMTJZZA5EEkb/s08tE9xW
hOjbVD+W3/QPuh+wVsT47iZNfNIq5KxKF35hL+ori+gTS6hqs0fY4TtO2cLsjpYc
1OUTSAKab6iflBezD3CWWWw3M2Z8UeybHh57nFVlZI2U+vxx2iP6upLG6/rF4R5f
6R/U9frptn5/2Gz/7VnV5sgxbcBRO6lMUSA7IX959jrAiNpX+vEsnkpJ1j0vIxTp
fJYMshZ6pQSaFBU6jEOUVSULJkJIKYCk7jn8oaobkI5Y3k7Zs3lqGgzCcBU1U8iH
l8iszVkr1HntDOG4PA3cPI6+oMtlkboLPq7qn5sVfgdmnFSP4dnIy4h/FMSXgdAU
eGd09wDs3N0FCBSIakfYLs8i7xLXUOrimwZpwDw8qm+RwUwo/652H005hrEzI4wP
hDKTJQp3dHJxeyFuhbMshQ5kLgNayiFO++h/Crz/9AzlciZNVeZtKnStv6zG8lTl
OOsYViMhpSrqX1tz77n3nw8ifY8dXe5Y+RXxb9wFqqrCG9gFUXHT1P+OOFnM3LWp
w6GHjOu+TBZOn7NVQw5IqcFFOefUFRfuA+K+egPteXDFbVaipTYHLWq3HtkRJ98B
ZnrU3RFsvfwbAfKk6sxnPFXwh11IzCAy1b6jbVetjWPP7vktZTX5+bT6taN8045H
rHUQu+RYNzSKaliY3eqZuF91wPHa8ntLGf7rhpk69BWyCVwnDThg1+sdhRtXCTu5
DEItCOs/YTcJrHhU4GZK5SsxzHV+m0IIvzGf44QVL/RnwO3pZaVHPgP17ldpEzVS
K2GWpjHJlfadpeTlu6/7sAPl9Lieu5w4jBdSSdNhDX3ubRl8LR4SNQz7KzIx8dZS
wNAnYvJDRBcYb5jqQ/iqLRXd3zLjow6fP+iGzOjZUWP+ZbgyqBk+lIvXT8UHuZgN
DrDxLvIrkm/7loYhC77/HKTudu0bDzmPJSbHo3+9gUi43MRS1NV2zw6c3y2eDXl0
06rg+M4u8dl1gOfcSzaOLEXtyC3OuBTi6wlBFSLtLUmCxvuQ3ssYOggjc8ILnXLo
uZd7h+Lrztc6IwttOFuXgphc+tcR9m06/kZzEIKdtsaNQt2CD2ISJwBE1Olrqgp1
n/VXGXiALFuhFdkZl0WAv6ipe2OyZCCITkai1bq5X11nMNMT0zmygLmG3PjYefsx
I9cBWdlrgpo8+4No43OuRXlSAu6A+Xi8Dy8tcxYNDTgLNrqua01+fZSbNOk9mhcl
YThhzI+4zsweY0+zKVIBN7YvKuTwx68zJjYu6VrM/9WTgActhnF3Q0DAck2vyAaN
TF6K2hrfRrUTbtf8TVTXthFiiOt7wlrM1bFDs+rrU6b7/TK7cxVEuTdIHnrL1rXV
jEnnR1o5FuhTIraDnVFBW5bGsI+fdz9YhWtTdf66mWXS02hJXvKI+HOLB/sgjwr+
zzrL3qAb/kBFYbQO9iZlGBLHSwaJ/T5Nk34LKh43W2hRoIU0aEiZIh/7sS6JgDtZ
nU7Wtnwq+O2/tI+GO5JOuvXNSHFd4S6I5MBJMLI6jQ3UidyO84U7FSlOtOiagfNP
xAVvNtMKotAnx67NgQ0qq3/uFq0XJVHaCFoxqMuIMY3pomiarMBABU27QLwXZkIS
cU51xRAY1AlF9Cs3KVB87LPWSut3wLm+RKlfRN1ZWl9Mc87O2j1lT8fV15NWrq8d
Hi09HfBAVCVv4XJ2KrgELOnQMBtYTJza9l5CSoLwipea23gKEhF2mKihXxxO0fUa
ChT0ezzfNd0C1VE8Sc0/UgEhe9L4OU3acrjUXjpLOzb6i07GPkYxpl0pgVQ94Yea
vUcQoWoC8y8MoWBTgmfBNtAhsaTuUhaJG8lIkEc3HHv4XRWDYFFiTHehcdisKqd1
7cnfH6NQTZB7xMl87uTBbbW5CfTUJh5wXa/PHrkoUwOTNyCR91J9tDLGvGueIioz
9ZguuWcsK8rdNUXgXF5al8Ak6Xmcqa6lUIiKM7dWfkNQBPn0JHPVrAPGueZlKGKp
0Hd5CuB83ZiAVtLtl1DIrDouplTZ/DFMey1EBCVXilRkfa/XQzbNR+r2+Ono8xrC
pEG/i40WTpPY9Rb4ar9YeTERhu1GOIaqsjSouCQWiV7SfE8F3vOcxxy6Z3sTb4Vf
fd//968sOHQVWIxhd1CtnTzR0sm5RlXr5Xq+LH0H83JjEQaANvmGnTu2g1F29XdU
btnWzZ+rhnpAEYThAz1DxvKXHV0Fbupv03j/KPLjHZMV3G6ADl/tcvGDYtrB0s4N
bLFhuR1k6gpBlkeS2sACE6stn7ZAGfQ+WoDg8eSdrgCO8FJLBeLcl4PgBGWbzXsZ
P5moWXmktE32Xax5YaqQNJHlxtEQbJxtYo/W8rNdN8fFO0SUy6LF6esCdELKmr8P
MNlo44wngRJHwfzODJT9syvrI4p24yGkBK/7hqxU7UqL5JYK7EM+r18srrwmBb9j
M8zdB6od3zlkmLlyB/WtN2L0/5P0O1eVefHo6MriLdAi5/pmiDuWTvdQns7qDKB5
iMwwQKLSGTsSi8hCOTlTo+MxVXMwwcY80W7449SRqlXQbg/4CUmcvn/b7qNckMa3
WnxwbehICA63/VwNfDkrmizHGs+yKNqAD4zC25PrS+TBo+nnH0ynq0SZ6ox2lFTD
kp9OdDh/MotvVG70cPEIRwjPlFHN3GKKBpu4KfoN1X1OSIoxcwFRVcA3ulOXFSfD
GmFXob8WnQtxoR2YQsalarl3yPFYSPVe3CnxZqXyF104QDbQsU0Xn5eOwAxTzuqi
rQ4VNc6PWojDxpGfS2Ch+5fC+M99WuwnPZGMwsaSv3ll2ilHKPZHk9WYCNg8NDq9
XJMkjSlidmdc7TMoeD/ba/xwW893Bm/Fotyjjyytk677ikSiHc2l6RoSalXb2MiU
vkvlsq2KVU1AGxkjXPfVJQPxOtmoTfpManQmQ6mEL1Ici4pQ9dep8vcyx9vPgc+i
RilhoL5xJ1A8sfGgWp0y7L7YmzXYZNuY3SKybQfby2PQWLgWBrzoQne5ZkxJpB/g
GStYaeM9au0qoGxrDtWLzsC9WtzO+7DIOe6VGwZonymYInBXNWPpfTXC9GfsZW1f
4ZE9NesImHGN4ifbVEKy0A9rewW1Wbio4x+MQP1EWvxc4qC4+JIP3d+jpQxukuru
PcaCfHGeTwFd2DUz3Cd1ZkOQ9DLXafI7LfNLbWKaqGbD1NZmm7e1cTtZM9nM3B1M
w4ols8J4bQr/Kjc3CtGQY/l4+twgH6ebJuNIMezuC44kM/7CU+IQigWFvGkB1ldX
50guF8rVO8iDv9JQZKgjHTWdkMi18qyfRFa21RHGuiVmSpRzStWv5IV+Dtl3t/JW
WdVK1v7RRfClWRvaM4tVdXCGS2ClF+1kgzc91974lVreAmxak0DAqu3ygaRxGol3
x/RrDfGPdcFeHJTtY9bXxYU1AkEfmXZ+2+CEES/6kEzQAlab3aZDyxY8Lo+3FLQU
6n8wq63NLeCDOcoulqPYr0bm9tgElMBSFfm7dNnRUB2bd0ylIvmjAauOiStXbxc0
dA/SC8CWMbndA/AymgDCm6+ciFdAh0s94Jhx0s3GVFauTdnGtsd7BQuQIp2RYU8r
NoEuhEsaXy4jtB1sEaZ6EOpNhjcpWo6CIlA4U8D1CDf9V71RT3GQkjT/sSS5gvwz
+lqobp+9emlao6iDdBoV0d6AB1iHKZ0i3NzH5MC4NDlI/W3zc/HboUj12zTfWmW5
7Qsc6q1DvK6nHwCp3I6tT9oFIi9+xrlPOB8PS3wdTdnFec1qhOPJec25jjxAxnnL
S63gvLw+zoaRFh0v9oGwqV6wrjYR+9BEOtWuAxoXLirPfNFPPRQT1w9yF8Mk5En/
0cwr4JPSg3zQu4Gqt0c8h4/veLsJa36R4SSpRWmZEo/Mi/R/WkTS+nXskqbjSioG
KrOUMMwxwhDqa+OB68R1a3Uli1/PNtcv7URFiAU25IVLmjStzLEI/P7KZlG92n1V
/sLXhAzE3PqhxLe6IYzu+kFNgSShKyUN5B5gP2Yl5NZK7kWRyJm612XQA9iJhk0z
eIbE5CgGhW8iN2UDkIscl04znMH2fpvhpKm8uhwbLPyWDWsIaPl6XPnhtZn6PN7h
Uq729+buE3Hfne/rNby8U2r298uRXvXE1iq6WB3q6cM2A5678ZZJHRsKlQB0WbaZ
hxbcrbBiHWIbRRwfeSqwoeFEJvrhSFarDzthcYiMdoefJvxOG9xhanyYwVpZcXsV
j824s6gw2j7Zh39iaOeLiQyoPuUtTusahCDCMvJmXKibQoWQh38nwlJbXx8m40EH
6tqnmjjwjcraiNYvy4c4ALqUW6cSOUk1N19Wbin/+scVxXHrtgbooSIqoRUTQb1t
U+22HzNYQPybnntRu/L6+2+MxoPyo4iUYHQUMXVFBN18RFuvTeRbeTLBsbj1zzq3
Cbuh2D5ZQbyE2ox4e3h1FYxyn8kthkfN7fafq/c3sq0MZGljEIVDJtBMiziaWf3u
LypT3WIPdkz0Ah/QifmwwEjzpTRgpXkdeNkNJRYe81EZHJdEVty8uAqZx4qRNx93
XIWm3jjbTGWPbV8685Ezc74rx39YY2P0B3/xClHTQ2OOi6L2JMZs06aAyHbKH3jq
59SJeiaaCXW1BTHoPyeEv4Qb8Cg4P2l31Ko1mE0yFlHlN6Xny80qfr4faewME4vE
yp6AZTDfF1539mshlfiY99iHWrUHtnzGzLgPEUhaio5OKrPgKRviW4yWpb42q9Q1
8rjoF1tjH6tHyL69alC4HVc6uB2hvsTwUNYxvAbqx9E/JY3OgqWGMzANuSsJiQlc
Vbt3U4m+ix/z/bPPtdksgkE9PNmrsgJaH4bFusZWy0DYF3+tWWEWgNkaKUaZR9sG
puwm6CRrO6OzAwtpzYnQI2qI2OKgY+nD8rmJ+suLYeLoMtgR89vFzzCs9jGAXmF/
h6DDO30k4O2pcu8DKJlJOkHfwPTi1KNwzWJwczbl8R7kJmSObcBjI0oM0HmgMeme
/HLK+9IVedFd/eVZs9Ck0MrV5L2ISYlRfTbK5YEbNE7IBc8gNuSkCgB8+pgZVJiT
YmfiCM4slPkbCQyzQCKWfkv9PdKkYAUSkntSkE2my7CeqfPqfqVASg8yeLKInjoo
7yi7VNxdafezcWFx4NvJLQZGjmz2j0rGTFTgn+THIth6L++XhrOV6Amo24Uicuh0
FmrbCGl9VejZkKhhx0uMvcTj1ijk3UDh3h/ixeuuB03gvZktFywv4EY/HfKvMafk
rF7uX6w6wUzHXC3LbJjceYKCfDt2UTNaosrKahbl1o2uOI0eLM5mGE+aFz/3Ril4
iPz3B4A6xb2xufNk0ml8Y6yuLuwi5IijI8wCRT7Mf/ifhPhIIE3+FgrgDXSF8prg
YWf81obZI7g3q93oODs+sT9w4qQ/Jdqm18c2bzLgJk1Vrei0BV/9YmB+SdbAG8nJ
h3CA6suGbXXLwlVD/IGFV1rOflAR1Qtq9bWTNn86bEKR7MTWBBEzsaI2v9LThE2P
3QcL3vqa5+qGGhYHsQqfebhoiQcBZbhLDWJcfVriQ5GwFaLbKdZv8R+/VG9MR0E+
JBOtP1XZpTRep82h/RNiD4EW3p9VA9Q2X2qI1KNJk0Phya2ZTXKoc2OjTGyxftsV
FKmqMhx2/CGTW7GYmlnCKmfy5pTfVL6R0ZkCF7k5HmMkhZ8t3RVME8TGirfmsSER
6ZEdypVg1d2DYfywpoFWkz+weFugTCSfzmPJsWAf+KmkMEiQ+Mc1YhEYMFd6bXgA
/3pmv2FfCm5+Yx0LQJG3MAaFF2AjmLX1+CP+zTy+i17S/II+1CvAtfYuufzHCXgm
oi6u0SARlGFACiJJx7j5cvL3rqSnYyUUbtkbWQxvHPQxcZAsn1eocOmEtP7hp1D2
q0VLzjyog3fgv4vx56PrTOZVzw4FP8o2hTLi8tkAoqeKmJMU5kIpF3tgaY//E8qO
zJY4Y31NOGG/16HJa24XDHZ3nQKo8/CdIxYGUbSj3HLBR4ZGpNIbwZ+Wx9YoD22l
WFs7SlyJ0EIkeCKIvV28fS51aD5jJQov8blV5pyD/04q88YngCa5Q6pNokX8+ifu
kkN86cJGXJWYLNTaYYQN0v179Cc9izJIAP+b1ym7Vf14L3mNNY0gwmX82eEEgs57
vC8QUME4OCt69RowNozshY/JwEWeo25hoQNYcvJ4yFf+iS/2pe4iiP+F1iAnVYSU
/99I9RDzap55T4q/ZWMGdRwuyUC5xpSom3a+3Gy8/1qFPGwxg19WtaRmxsH2i/Cb
moYOdr+hTGcKn2ZSNCDzblDmw/+iUMhhmzdPHbWiVD1k3GzKNJw/r3aj6b/Itptb
Yw9+/flBZLX3StuJHptEkA5y1uKQQ7X6ZlIQ2LBBo0THZbJZFrcn0VdKLy46h9mA
N3YWawRK99P7Xovlhupl+OtjRCoPSY9ok/B445PAZ7kxjYwBdOPasoekseJM70B/
zlqQI639Ps9FCwO94R5dlRa+w59aNsqU9l64hdajddY3RQlo8bayfwuOLcyBuTUk
PfdRYf+rNnXv5Wacl1YDw1bny/3qOTh6vEFaQjB1X8mynFXUtGGIlTebKZ37yi5d
9dcJ9sfO8+6L9/rKiFqjSvWKI6rSRO5O0RYaYPie1i9J/KrjVjpR+oG/V0Vofi8P
St+yIN1lDIYJFImR8JpWzzBO0OHqbpKPeu5/Frc/ijZlMAVSGzApGgBGCR5CAwkG
spmrfFC2fDGlf4u7f050B0rLd765sDTVf/9r/kj08oXjTQklJcE8crdwP/Vp3bNj
9RxLx3rwTGDKIYe5lw6p13oJTikGMFfhSvJh0u8gPLjXbcHkfk2hTxo88xJNqxQC
fIs2xH3k71nDqxK942HqK1BxVSt2LxWtUDbLBYjGi7UtQEv3hqAyZ6sxW+9NE/3G
lpt6hVb1A6Mr8wAGIt3hX3TVyH+mKF7HvqHB15hbrRMjiPAyTgY1LXniq982iQ/u
VjFyKMuHk/YZ6Dh4pVkGiTHmJousZUFqRgu3OwgeCkAGb0+anRkJkxrSELaatdB2
5RhBLe8/SBG8dBjkCc+zwf4vCA+M/W592fFX7woh6m+5p3jKAvYyI2Svrp0yaCYZ
Y/WNKzgdDyHCsuy4zIxXMjPnkv4ZSPr4H9o85ClIKITzzyF9fkLaHt0daLnNIcVn
cVc+a8d/UA6XxBLO+m7OMqUE+tuA64xl4Wcl6zPaYcrrIdksOoJ4+w27qECO2ktb
OnPkHW5UdZAWQ+D6ue2Rr8bQCjRE4pVurV6vF4BqZJIbQOufb8F/zvAs8pUmhdEr
27ZQ8+fKnVHG3xwql7331EvkM1wnIw/nmIGnBUym3HCJDWQtQ38n5bBQYaguAnO3
nUt/zwmHxAtNC1y0EnTbaEYpCt0q7eUmJE0BpIiuGoUqbpyNJ1IJEMIG5yw+C+ip
Us1k+3xOUk4G6sG3fWLeQO7H5vC/fMxVySGtXQ+lO4EDf5dpHHDfbKaUaa4oYaN/
awNczMgqShbAv98g2DNWF+YlI8nswbYGxYyRaqfO5wkwAh33dmItMp1CtOZF+G3u
QQ0rjUygBvHI7iD83tDt0BKNMtY/DF2D23NV6lV65ZCMPMU3dciZbPxDnlo2kFNB
x0UxhzU4QGnPpzUoVQ2khodEMc0xUxzsFlpuiV7jWhz9Z8A2o9MaVpsy5qcb+qRb
jKUhGzh/hVa5C+uq3jbrJv7pIddwQk3Iy0fzJ4UQe/9p5kWaSkq/oYu+GhiRKhVY
9XTmqwHsoMqrviRS7OclIAKNJsPLndvu+T94Qjshs7ggiHZjiNfeIj1j5T8wt+EH
1MOOxbwJ+Bu/6BUsyrd7WChGizvBICLc6GjpJeYZddOFODRz7RoQOHhJz89RmBWU
DTKklH3Dq5JyZ7IVK5oHmoIFecx9MiF8v2Lan6EHcYWEefL68EocogkAK9gyTNqO
o922IUB2ZNvWm0r72Nvx8UbFs+55Miw/glnP0RY0sYyfocHmoRb6SppG1gxvmsIt
M1LX3+33SCMAtjqPGptaDwFYSrI7b38499TFFBnyJLQduANTsICi6GduuAf3Q+n/
aUIIQMFK7YzVxCVQbi9x+5D/Q5haqGe7WyT3x/DgTnBwhxe7rlB3EwiY1njw7EA3
L2UxgmdwWVGBaGT7aTmt94rINN2AtnfkyHm5zDaOuyAxLQqdkVGVLy6DQZNH/4ie
JXwhIF1+ht/gdacQSJJhUTZywNocgWQBDoS1rQAZgmJswVzVEUlMeCbYQo/0OtOT
aDFVlMjMuVymcCTFyyFUF6txYOEgO7rf/hV4mmIoFl7CnyQlq8w+bTCTqgT3MWli
9LoT9P6vBC6/aMZ2/RRJHSsTg+EaHv5MAcZIHh1Ig4pS428gcc1LkVK41FmUyfPz
qnml9F43amierl+VtYrJUfezL58cbWIqLMIoxAUkvZ5+3nXBXK/2XnQYbNkm3igY
tu7fdq+zLGaPri6dJEFYkeogXE9Qi5jdWOLixY9WwQ/27b1OO+ybi9o63XfCyRan
t2w2bbMzmr2klstXHUSGgtaFd3oURwaTR9gLCJ1DSHckgSreT9ox3t5w4mulPBv6
dhDyPvZOkFB+/olCrQC+Do1iSBwMski0ddRJJrkyuiDYzz4Eo1PqdUUeg3ZjozEN
NL8nyufj67E6d2nn+IJv50WJy/R7eFZ9bpYiKhWZsDgOWj+bHBtI4bZBnaLHq0Am
AVYMAUJAw2nml5DEpGlRbShnkbPzOyYxsXeUyhL8v/ywTfRfoF/tsbpcfcqpgdTb
sXEdIFdSXNY3iFQ3fzCxN9fdjksYL/y/V7ieiuJ7ANyZZhNezPfAh/MZrR23QUr9
sUmQMzm+r8uMDFVyXPYpRnTp1U5VXm6730NiPJQ/pe7BfUPNeUpOhMdA8CWvgYfZ
BoOmMX5ZkdxKxAuWCPXtsUMrJ2Vm39ax2iCDHZYxAV//wrBeVj1dcqTtjX+MhLoL
y81okNMyvx18PYBy63sW7IvNaq3yhqFYkterkPobrdX7YoyzZgJ7hB5igkSQe4GA
xxkBNkydp+yXZhEeYNIS/fCWkJyxUQWa+9KOnKUjf6cNpfMnggqW5UNH+CC7Q0s3
LxwZG05rFrmYqnXJ6Dnk+tLvGXfFICh7fcuSVHraYxoGuigZB98GqFk74ru0L8yx
XnOMrd9aHgGpDNA9l+GuFgpGXm7it9KnGxJS+24lVx+AUh68tej16ELz1/Vavt0W
naMuel6fzMf8mOf87JFn1fmrAIw9QraeBsUGBrUI9ijEj0tl08rp68OqhZ8TgyET
gFDERWYKQ/ZnhhsBObpcddIQ+pu50+UmFGO8PKbSmTPunb6BOmuPYCS4LNiw1x5A
LBTYNUEjEs8YNKHW9XGoruT+9XEgI1dP1/pXOFoNlDFBKsOFlNioRg6Be6CxBjgO
LyY1gq8bpDmKUgQyHaBBcPJqtA10bfxkera7EFNjj0ldS9Nx3K98kaJcZYBtmEJm
UXJz/tHD7Jz7lesZ/Lzqvgrs2tB6PiLQLP/M9NGUP8ZcqBiGcdFB3QctiaQhk/8l
NXp5hKMxZYrblYg6IiNCvMKByDbjzEFv/40xocC0E62GqyxqjxQy9WWDthiItIgE
0ZFiuJPfBA2ItfqQ+5RPgUeAxaEfex4H4shju/Guqs0ctFozRp2g8EryWjrcJuLN
i8CY2bn2Qpd6rPWrnCoE1MHBdZzIiSlANjuNfdTQLqGT/ju6vBRs6eXrdAlcq0fi
P0T1AHSvidrXn7LIqf1apfCbplBg6vVLC+ojplLaNIjVsVYSXVksw7UgGN5Neze0
N/rFXIhDWTOyPXnJ4oVlOP7ZDP6ngNramvd9dhD+mIScbEhvtQ+lpSYCGck2W6wF
MatqcJcNoGc3ebioZ/rKbBFHFT7Su30UAWzyhzqrymhUmGfsFX1QefywEb11uAZ9
av+GoJ9pyMFEc0F69a3cLiPFjLkkdTwEtlffudL/dWelGxp771Pl6VqzUTi7XgJl
bxrVD1+KUPS5gb++uilT1T4QJ02CgpfMnGfhj7idwA0qcAHJUxLg5GFgPH0KKSnE
UOFHiT1dDB06eZ05Gek/8gkZgRfUOQlfHWic+3BrkaICvWtzwClQk//HnAQrpRu4
cnGq8CWMMcRgViJmywQE9OIUoqN2NF8JcsFPd3VL7FqTxOL0mQnBse96NQ6WaUN4
VfGFjO+4oaK+FMu2YWfsaCyNywixh6wY1CIP/dWeBzNFGp70OVrWo1UjoPyl/+V1
DRxkJ6BcDPwwLvio1WUO2g/sTQ1jfdi3xAVs3Q4TrHWp5kYVlnTQbbFErfglxbiz
HsCTpVq/V+x7iwbxCHs9D3lN1v2OZubq+yIudApaMeZVBdZgT4PlW9OKPftR4+nG
VL30IrHYz5PeaQBIYmm00W/iQdE059oLQxx7YYPnqQUIg8dWj5ECYj9LGLyjxA66
PmEh5i0lcAk/qsW1wErw1jasq3tLLF98RsSs8hHYN8RM11khwmjGQAg9A+RpdMFx
LZ4dJrfFUASam/czcsbN5VWUke08WqI1fWsL8oDMkvTdGaIBJvB0lK9Q1jbmksuC
wUkr+QYTX9popwWGnOtQVgLLgWHJrVFVKBDiEuviK+zr4+D2ryPvsJIvbrU6g9mO
t+xWjbzhYkPQZ0W6ILArdNQsUOhibUgroz+q28d8MnfNB17EvGo89h+FZSOpQ+50
F9SzgNQyGYbzuRAIsGnWYih+stVSox34lMhIARcYIQXN8eJEnxPAzJ96j5ZhXnir
eERB9j1LkrdvJyJ7hThEEm6YnmExkJVu7lUSM44YG2SWDPUP8RZ+0dAZkoUcT6F2
2HcWSCki5ybVZFPgd9yUo57usTLaxBnfDdV8+zfV9d3eEm2/4ymErXyEMZkNTouZ
FegZS/zDuXtj27BYOvsAu9maBU3No300fh8k3n1pIr15o79rQSIrK9gaJ3BA7r4Z
H3/8oQPoPUj6iZPIcLUJplN/LG8oqE0oBvhVfn9FhJ71ya6tDuQmwkRi3Q1gt01a
/JpNysIhctxHhS15tGF5wQgGsUtM/bewQ67HcZzADqXvGkk4ks3g1t8AGx6Ven+x
SMD0GCJKeDfdOvM9IZIe6arbY4g+Xfh+QLv+m6IqL9JAzUalmT2/WX8hbgcLD+Kt
lFN2CZ1OegCKpAurLFV3sC3EfpLm+6iUMeeO07ms3oqX0Fu9ns3AnwwdORW5NFlu
wxdjK2pHPtCho1MduFnhcVV7EPm9sG2ej/Gu40W2KwpWhcefvomSPDFWUO4uCyAd
3r+wJfXgOMIkgikb/YVXviPk4jOrYU2PCCBy/kz7suok7snyOW6P5FQkKspnr2Oa
X5od/sYrgCV6ei8k2ouNuR+fSfl8YhFlHNDag6PPzVwksUdBTwBR9gvBoGc+0HfG
UJPjm25fgbpD97FMfjjD5JQOlby1uNt5ewhsORUfA5Uzwjy5QVCo8uuiCLiJMEAx
jQTf0ioSaQjGPSf3Y885oLduU3lz0PK6PYoSerCP0DHO675zu/2F0CPlyKqx/Tiy
YZK5/vBixY+6CvTk1jwRu9NBjK0KlayKGTCX5RWDX/zFJbYUCzm63qI6qK742D71
N+GKEBf0NPLEZvNBPBpE4Nfhywr2J/XUyEybi20ECOexeSJELImGkUKytrhkrNgc
xxk5mGiC6SCO00hsdT5gcK0rac3DiWZTRKPYh0y8iju83P2e0TRsefYmch/LebP6
u0Os8m5Se9f7Ez7nhlulXDRaXW01D4+BJkcLm/WkiEbxxKYcd4C/z0PxGhltFPjE
gWiDO2oapo1z7UAtl9+jgHmejc5VEfopsDEcRehfWpkqFdHQuT80xFZDA1Vd35Ig
RB7t07Gi0mtVAgj/5cPQkLqKT6hRd8+hdGSImv5d2hJKtqOr4XWE7MRml9eEBiuc
gfNbsRHDPyL9iwOqVH6WmR1HYMR2gbJtBATlv7eTjoNF4nl9Lh55Av/DV4sStf6G
tj676Q1XUdVJ8npZFjfCl9kPur8iA2Y2j3qGOzuLsTxp7Pgdt4fKSVQL5oBy2KG7
HlINtvV0leY1OToHzkm4/0fDaf2hX/mYKqPSScVDAh5Fdc/nijCYMkFOKku7t3z5
RRAwGRhFClmwHD4cW+UVfMaUP+m1yBkFpwm2lRpVJ4gnviV6tFU5pIsLN6DetW8T
fu/p1WSNWaH6/J+MikSEY/di+NbvcqAb/dN5IhqAm03ANngG2WmrIY1y+ERH4+nQ
T7BOOBoAgSIgxK2seEyy8Zl9rGdd6ppou0VLuxe1TEoekaqWJGNiA2pIpG+mJejL
nDZcjd/966SE6/4wldGVhqVf787qBgH+7ga8jH4SkrdpEyWiTOWTRZL1j9g1RdAR
ESybECZy9ioz/s6Ry5E6cMpnSphORB6J1ETgq7xY5RJ5H/+uTs0qTMqarZWWYGjj
anO3z+qS1ljjZKnRZ0T5sZJWziStxVVhi6v6JAmr5uPmKv1x55EpAo0Q5/BHgldv
BINBVFEPr4GwtwiitXFdry00BD41+URR6tOCHVLwpj2vN87lxWEHisBSDKeR+Uqw
CJw3prET73zXBrQJ/mWXWQFxlSEPbOfDXz5fPqRBh5EqPt4ojngSEWCfRpC5SjrJ
MU22Log+IIBQ2Q4fLtTZfmRBK55HcL7uCzV61POuIEkjrNFwTBnaQHXrLqW1w0mz
DYrWlq26CHuWwwOmi5l8hKQqKod2rpu6i7aKeSVg5c9FGRzHx9Coa+lpGeJKJsFt
RdKMv4WFy/Z0nVRH6Xd1G4dK384lFm/WojOP6kNYJR4QGZJVksbcFNF29zPklmVI
NEl0j45DDgmzbgMA/gDBl+JPJ1tNQBjkj/XcAk2g0nQii2Q89lPuEf6Ctv0kAd8u
37hCDY6lHWYcnc0UDyLaYu51eBgxMd6nePv9mI+GzLelZLoZOhwQy8U1BoWZ5ALh
F3NCWqeYVzDlTW7QdZmVR5wyoGoKrL455SYm7AFYegBFGKWHdrC7ADSi51xM01B+
DSwW1R/iA5EEl3LXgKoEIBKBzGKXTJ4akAWtji4fvd5pbZdUng9AM6Amc9EwpHBN
XinMgPDxyDJEQSOCknHuUb4ri/d9tFHkjnKcGmzyyQhECnrtQvJDop4BcOJhEPTy
66XRxhKnCYh5ZXmVqfjd7D0pAjL91AvAhoaSwmApE35fOHB8CMemi2AxqzcbM4+5
XczF/1K52nP3P8eIl8lFWR65GBCOEKw8SSHJmuL19KLjKZ4g7XRZKig0RQc/30YQ
Q7NRJCaNSeh0RB5p5SAqDDbg5Ggx674kfK5yQWFllDxnmTLRh89kZOa9ChgccLZI
FXm0I8atIL1LFujz8+z5vcxz9g7rDfhEaWlPUmB4/mjoPDfi6MGO7wikEbbGT1s0
qd+nIT8mDF1LuUWCWydpxrX2u5a4JYV9wkprQ1MJPmUbZTqbZG+4rrzjwBkt5jhM
Tt2PUuRGU3GVXAv0/W0yo2wre+I4nKxP36Qg/awiyqDmBoS3nu1vtUNtAe9TEDXw
vaTDUHXMLw2ho5w4dddJj2Tlx1ug5p/gbpxOBQ2qzKhW21JNP1AkiYGZv02w84MQ
FAa+sQ0KfT/wHs/ubcu12IPzNg5v9xQnfjIYvxkE8dylkuCrl00lqUf1i3PyQPq3
stTS3RC6Ecx1yk2Erv6U0nRdRV/Q45ra9Y4l+xS7Zo2GRviIHxXJDjqttLKmaBx5
jn+3pc7t2sN4SbzNPOJNCN7Hxq895J4By8J63+WRW8SI7InH8IxZL2+LiefuFFfR
SjJlG+xef/6fDOjI7fpu/glIas3fb8TWu9sG0YImmh9YKCj4aaEJFbOTqNIX44gQ
ZBAUnCR0/5F8CSp6s8xbfgFXOtRMhLghYCmV7PzTOBCwomMVMm7B+pBPeK66IcQu
WfR9aL0HvXDJbxylt19nz+pE7UNn42fHM4laWe4Z9YaiPV3VwsL0PwHCXUOrd2My
+Qv4G9kH2yUzbDEW6aoCTpH5z7xHz4rV0HVUBQONRL/w5gidygKWEvUmcpaGPobk
rOX4tYP/Nyweb2grxN696V72O5RK/n/S4mTrauZZVdxch6sZCoF6XDFeoDI/ioG3
pLH89QRta1WFXYHlLpdB5zmKcXMcxAVFSmMGfRwkNY4JXs+6u/tf+8fMkEfenXnU
CH4OmWvoo5iu5Sg66l3sXC1mYcDzComcqOThcNRzn47Ds7Pz9UJyp2HkdrnOhVDd
OzONeS3VVCGPpBGQVi0Pq3ZnOd+iz5tJ5Hlr3TBs+5QWNf/tWMNgKjQ+wdiZEg75
6JdeVqyNEP3hsS65fBn0DxwjN1yG3O7L1H6rb1IxRjhL8lLG5i0dLwFKg0iR7S/j
G9Oyx361REzeWVK8EvjhBBsNhWWxzvDPAyzDsh5O4pJ+R0FoyeK/Cr9mrowWQ4ad
vD2hQpNRcImwLbDbYzlE6EomLkUF0bLuZoa9zBHV1V+9iUrzvcffNBYPVP3ER/uv
UZQ4mTKcYG/Yi9btLMz+W2PgWNh/KAGcgxBq1/rtF4Rzw3iBlU3Hx5ByOX7f6DME
T8SumlkNnmIu1TTi2ct6lwn46fRvHOhKBygA6sgZvBXrQ4b0pb84M7hZm7IBSyf0
7t1Vp39Yor/PBfIsshC8HY7yCfNFi8ZuCK69n4RmexQV7A1dfMlYt/2hk2zG80az
Dxz6wZuwgO9wVwsWFUG+16VFElHJ8iU8sQLRjeL/2CQqNUdbCwhm7l9erYUDyrRw
UQe8Mnm5CLDipD8m2UvN3Xz2FPrz8YwB7BvQpYxXgW8HlS5gBwDd60O8zY64lPat
7gUFX+pa50CFQ/MZauZICzlmkB+oqL1IfyITEXFZiFgZZPzKF8i1BFF0NO8Pr+0t
Jd0Zlfy4uAyr5DIaMlHf2osPQFQKIg3XhXUA3NA4dDv0/DV4LInK4x1S6YO70g96
oLqsMYaFI8W2rtU4BClErKdpthq3EoJUl+78Ec5/Sco3CSoACDiqyUxWpfWe54qb
bsJ/S1yhKJj6vPsnODcGaRKI3qJPB4njjsvRy+QZ/k2lLYRa3qWR1URCVxOq95+6
AHKVL/RN28/S5+ShBQgFBztaWZgFqA0oeklZH6d2/MoD5f3Hgo6zK/VWK4xIQv7Z
1k1/mXh81bT+wyzdPRu9UqyGOlwPx84rQMX7OSEA2ITEV6u7SntmZZe3K2QcO3cd
K/DBwzRnqXWA7RyHpnb03gjZUvPB92y86qrB+pbaHakZl7/V3JLikp6H5edz8RN4
QOA+ArmTK3M+OzL8pGOdYgaPNsqRPC6gssqeewf9i3kdQ6KXS0J7CXwJLcqolGId
jl0iFqw+xKyfcUs+KgZkeL/BryEXZMtS8hE/AFZ88GWKNYPlUQZVIMMs/1JzBCyF
sQGpI8Dto8dqKVkof+udWcoIeOQquJnjPAmlfEXksRuG7WC52qAbw4C8k5cVwCdF
1n5ruOMuVHgwp+gv/NeoQAbR+bN9++8U+KunBhOi9xaIQRLWbgpVRQhkAHwxjiNJ
ITziZychcfG1UEn96QrnXd/9Z44+UmAI7jkejWIBMIrVR/9evY1A9rPMScpBU4J3
Tfbhm1+Gc/Chrfk3YIph1YLem3x/Ki0hqd/ZVemC7WUONtL9/GEunQIpHQZRvOyj
DIkmJLegtoOiaaLFchV95g1LF9B5zq3zulXH0n97wbE/C+qdkyhzjIUrk4L8LUUu
WrEWrFwGSdDJg2OmlQfJtUZ43/39XqEydKlMifIbTrNZWn/HOZsdpRtmAQ8+Cbye
HvWPhqTBNei+GlALC0SXoApAg6HRMIq+T346e2393BZepo4MMN9tC0PftN4zts6v
8x7z5beImOiyP7+FDQ6nMwIDUonKJC36OyBpho+MfBycPBzON/SNAfCox+H4fZZf
0yZmMpUDE5LNqb12H+HQpHKS5fYbGRGyRkTpdn0H0e7Hcj+phz1EK5eVVwCC5lMA
Aj87IMDJdDbMoqK4cNSensRmwYYr+LIs1kL/5yJ3qsXR5OL+rAFEAeasHbgngxer
JmaiaB0agbTvaV/NwNX+iK+oCkFkBpCTQ4PS5gb3DDg5iheiot6vT3Y5TgwTkYS3
liGdemHhPbmBFjxjapJtvgbtmVjASNgwjcJ/cFoA1zOkA4f7JMJWbLegmTm7c0yc
Qn6AkVkRvYiyeQuCYq4PaKEx+oWmsEUkZ2yfq3shVCjj9zVv8VFLA607o0CH960Z
givgNiAi8M+WfhPVrHTvlKGuWEjgVDkrNx3VS64kaMgwqSJcRVsFdbUrnSmbNDZf
fzxtNe/etf0EyAZ8eoKbINjhvdVdpTIwQKGsbUEXb0YJK1kV2tE8wAkfOZx0lgaO
rklPsvHRg2SLUDewP3X9IWXZ16X590t0k0K/FgWBOX0llul3UbmvPDCdUFoGXosQ
fFcfTpLYz1BZjU72pZwDoCfux+9hc509MpEBH1zAP7Ak9U2WXRUroyyLW7FYl8bI
fgK/mM2G9JwW620j3XYOUxD+0CnSaDfyXH3wdOy2mixVVSXPTCLycnQdINBXkU7a
rEP8wp9NCdiLZicYVNY35P07HoxNedVwXoaKS23PSSRJojVq2o6Vp8A2JNxqbCMS
/aBLLz8rngWDLnBtvU8nQF6AwU5iaJSV7gXuQM0Bf3rjV62iQ23q6450Yragnd8G
bLdXNOEnu6Ca1rTIufq19UTF09f31/Bgv9yIObJnxkzJfatr98qQ8x3It0O5CN0w
vpVK2lr16j/Lo+FRs5jF3S1xY1xIwQyPaVS4trRfxbskXIW4t3/fGKI/Y7Rh0BaD
t5EPNygQM0YphIKqeJxofOJaqkU1AgBNJ0D1HlUuZgueXLsGhwTiRgQxh/68hwDO
mF2NkvNi7AsiM6XrvKlJ9+tmJYKw4+J2x/zNL1XhFlu4VvKuj7OjAj30b8+F+b5z
rb8F8RoM5WVcklyKaQkM52yrsMQQLa+LJr9qubIX+pni1bJU0vqKfxROps9XqXgP
01m/bOmmvMrJkm9zh2TidopJ4he+14FjjHtwY9WpTCVXHzc6SLFNNVwBm+PqXLz6
BW1Fu8ZD1AdqMPyCHPzBI23Y50sMuSrWFkAmSdFgkYpVpNYhxIsmyODajkvMpAw4
h+02AmD+0hZcoRsDqmk/cG1iol4+Sc84PZnTDyMU9p86+CEM7rwrsW53sTXjq8KY
ybrjEcjss+WC3wnPhiLo08hBYPNVIgG975q187pL+xwCx7F+wBAecY/8rh3tt1GX
idVNq+2yhebBA0vsO/w1XjpnLQUi7dRKtzf1IJj5eBXfHh6tJMCEwQyGfmZ/cSer
yWgFD8LSqo+okMxLE1vTgVH9umXvB8NxFhfTfMUMVfzVcRd5pwgKDg0Jr6IJOXEd
q+zV3u/lUzMhQUvK8ArWhqN5NY9/rpZf7p53b/HK7sHZwbPO+3+HqqZV4dvDjtVP
9HeTX3549B7ThNBRj1oWVaiwWbxEY5vPTIRa8BPAllp0iYRWqvRiSDKkFUo3hCwq
Q1rEcVACeGJFEwYEpAh8MPUrRaGiGZejAeZ9ylABrxepfQY9LBJ9EpyYRUjRGL81
q2hxwZyEjgbGVdLTbizFWaY5/Wpz4Xgv5i8Kcpnbe/oc2xSNF/YKc+aclk2J3mGg
3PX1nOw/M+gtDS8V5Q2MkuZ1IAAMVSTaVpFazLR7qExILlQdYwgMvaEUN17o/5xR
UWnePLLyFzSaCxxsqPLLI2Df/MWEM2KOTJXT6ZmcAXRcv4qGSak4MxuDtXsqlAHB
xKilduiG0QgJv7HuM3ijD81+SlLjb0ZjMId2UlVe82N6Z7AydpNm+Pbsi+pDkpmY
rX/hMhlf8WHYdJDFDXx/qLakL+ugTgcgvCqjTDVXN5/PctVeicS7mYX+WVBRjN7m
14+7JuEWeoJ6ho1vY/quh+lnC4BcHQ1TH2ZG+vj8KC6HEINsqcixgplRtyHwY4zn
kWj9hPot6W35LXEpnUCETR9/wr6Sjkfy8E356VXi2wL7tu0nBga9/3sVxaA8INhP
i1ORGafTrToNzE/gqdCEbUF4sQsfuXcoLyasfhclC6Yq5WWRDX7ohDb9wGzMt+Gu
JyQUH7RhWnKFP/3jRAY8Opc9x1vq5yK91/EjmOjHR7EeUvyKe/nQFV/e1D42HdhI
daSkuRq9pdZmfyEgYxEMh/tHBeR9+XJ02l8sGpZjO2A/u07N/GMJQ+Up3YYWSVV2
FAniFp9XqJLLsXtsn7fAsfmeYFDKciad7xw1CiTVylJRfmMlcWan6zLEB0WBrDnB
ogVMheIIC5oTd7RXYLfh1AwIhIMK96jqlM127IXG322pIaVjfvXAnzOSriLL0IOO
KH/xf2Qk6QlGMITV9N5nLiug2u457iAW5gPkrBVfN0KmClprvKk3VnFTAqaxNmwi
WTmx0nH2YXgN7xEBPawp0f/dKEbS9UWoW+cpbnmJ4ojYcR7nMMBag8I+Qg98EJbF
YlsN8s8RkmcInTp/1BvnbdgYPZLl9poIyqvQqoUO4HjQ0pHgSYnIJAQvVZVAT8qM
J9btrSdpv5SSV4Nr4SBpx3nDMvOPwEn9VHRaCgyH5IXvf21TL7TQ08R8HuEFBNPh
UkjdT/V6LYAtdDmNqQVW11v0fDJ8cZZL+YL2u0igoY3fh+EZF25H94XJ1SJ1rM17
6f2yNNIlp25prE0tzqxh6KMiOhWDMikM0ByE2Fj/98PSOEWvaus2fciLRk9k0QjP
a3YjUQKOuXMB3z+hJqcUC58fSdNc/VYKroVHt2Vvh1rBkD7EQRptrn1GG3nJv1Os
euf7Tpy0QSTqvVmtcS5HZjgEXKFIOFzSxPiXXuDV12G1j6LyTdJFDs2zg0XfGytJ
FJwxmkZd2NFtpVGFfdmKVfD8B0+oBmHpZQrbA7Zbil85htlShmzAfO6mJWgME6Iv
Se78xsTH3Da4kFrHt6cLX7LL93LxbJidCmKK5iTB5s9jOiNw2fUS3ACnszGmExqJ
p1RibYqLeuaoWiDnL8HEiNkFB8u+KdMC2zUq+KckD9e40Tiw4EF/8lLdpwaj0dhg
GZ1TZPWIOyHPQJF0LLPMo9v9vjN+0i0tgWtmN8Eq/zTNMd64ZjBQgj54OJubDkTO
hC5/5IGYircHyDD/QoGJqP+mKUbfysbP8mhzOucz44Ym7dC1DlQQEX/J8ikHV7/n
5nWuXgChq82AsqYpwNSOFky4eM5ddJvWlzACaZPQIz5fYGp79VRJF++pWufWZMHB
+z9uX4sebDlWBZ++YkW5J5QpkzWw/XhlDdBjb4r+5CPeo3rgCLF4n18+DoSea0EI
eUh4biAiL4ZzVtX0Hvzqt7rJhvw8OLpCiN0LsK7t9d7ZTMipRjGGClctS2G7FSJ5
hMHpJK66M01HYqSE6uoJQ+naOiGgpbgFIggNZE5awDHUTEI3nmkGYdkh8LzSLbPm
+H5DFd90+GkTl0wOUYkYj+oTT6nIKabfSLRrL5NBs4vFdSb4aG1VlkZ21aVfb9QV
YXzlsmpjhk2H99BoK4YmDDiGRND/ibSq19D4G1WyCubOPVOblyipkSL6XmfKpcuc
0CshqKjF4UgqvlhxsXCQE7Y/OCQpBEdRJrRI1XHfIkXDeaDpY/bb0C62rLewEP7h
RSBneUV6Mp31nkcr9H0yN/6bs/+Icys9oqLPsSYmv2X2W/AXnqueHz/YFhGGH2QD
qleglGeok0Ndo+d4dnf1ikNRMZsszUyS3wh6bjX2nJqw5Q5z86/K1yxNOp4vVYYE
qE5zOcyBZ1utf6fgkFRwdW5be8uN1e6fXJK9H5Qbx5sTp0BjpQ74lwlW8hAY3scG
a3p/u1MZX3CMDxn4gA78r46hiuY8yMZyldjVChXKWvQDSG2hNSg+KXQoAfLXI4fM
K9ZnLQf1lWfYRNjsvbM8LXRa2Bm8QDrRpdwgVowhMdhzq54ClngBH0ZIoiLIOGsc
m8bii2e8aTUQfVkBmn7B0M4JnxeBEc0AxORrx6up9HcVBA7OSKsaCgd/N2Fv1os9
/pm790RPBRzA0ARNePrfZEnh2IM87A1wNpUgGcAN6txeK9ylQjj4W6TfcY9RsIg2
IWaiNjH9O5Ug7NCRQTv0y2YApVh3jTzz9oCMgvR4yy4iv00DN6fuJ5uj4QJUvd70
a7/ZTLqI3uivuN6L0JqExlKQAliDdmB+yoDPscpm/IFXqGh7k6ih+Ix33neVUUVx
v6jqDVPIDe/+Rhol7Vlb/4ERmmwKOfZ0UDlXkRxJOFctC9VvjPvhsL2XMJEfKL9S
RAtLY9MPYBQmRlefbJ9hYdgs1cRU++HKQUuSB0jLIjhGfUQh3dYW/vF3rAmb9N/C
jV6B4ldNjtdbMXEzUzLZfwrS8nZ5n4j8odVWrcDaQVKkE8UJ+P1zYFSvrH0lWy4H
wGviB85CmlmkW5bgJA8fjfmwHA9wimF5dTdwL3VLp4RE9mvurpjsZYZ+xvuPTOML
31XDAN3VnyXUpEvk2FUtQK+Gn2AY7BsVQPixH2FXEErhGXDG/qUYUunRjXe0EOqa
4LiUNPa6cBmCc2FhtP/dXWOYWRVmTjENfpJyymkLBaycP69DLE+xr2hdcR5bL1xe
N2b+Kk/rIrbc+YJqJuCQIfYzjONov1CXnQj0L1h987tX/WWy4X+W6JvQctmzb5wR
zQFCZp8muxHxE2DeNzjJtaome8PWSAk4cE5PFXZXYUyXejLOCaKY6lup5uWqU7bE
CAFVSJd1nk/TgEnUkkRTz+gbjTrplRSJkxLWWywdI0uP3VjOGLUg5gsYZYIDeAdw
R4v3z8KWOxDG3DfNv+sN4K8/36grgYC8MTRIfCB3KS0tB21p+CORZzFdfjp/f8s+
9+mGoluB38JLGBPoLoU7vx5KKhjUm+TBkbH/3wzaDDkZ8C6n0hJdqAuR/Hlj7Nij
auDkr6e1/CFOdzkWkob9BeEN0VI5+TVjZDJY7iG6XU17ohmyFCnPz41TTSjN7Anw
DsgiwUH81+NJd4brKddJYUG/rgeaEjrl5tZdBm7Bn157eWHPfeN2oWVa/WZ9IUVj
30IzsfdW/AVqw+dijweECGZ4wwy159F/QYXSIuz+egvNxxBg3jMdT8OoLge8anb0
vsDFanSYeRkBKY6s9ZM5fRWreX7+qgZMlhmHdkizxH/VCEvN5mE6cVvnpZ77TSDd
p0HjAXtQDExDkhA8MUi32C8xMutBShDHEr/TrHl/w+ms0mpgKyBaJgmHlYY+1Nx7
TownY71UYs6rA48aiZo6bMie4i4DWb1xe7uwhczGovWnLhqkvEFbGXaC6KtOWPqa
T6nxk/bKN0jwDuFHhAXbwdL/kCnKmn2yW2pImhvaXArfSeGLCyA19+TfzSuaGZuD
50x7s43jykQcVFi6LeCyzTu1s64lMpLqeR0HnTvjPASFIQrLpBXf7MGnkSObmZF3
m81FhwfIVoV1s8V71Xzi9V7JA3H7Dk9TaPIkru+7CuZpYHDn6o6h2vrImqEWQITW
z8gjr/1U1ejLicTgLUkszYSIbJ7gUvdMPJArxE/2cCCUvv06l6RIrXpyoiofICy6
YM/nI+34u46/jxzKIp3+5CQyB2/NAOAYRrGxBti+drNyvLrD3YI+ph/Kl/W0Exm6
WHGeugYZg+6FAkYDLyMUzHlWS3u28Etnd3tzg6oOLPbrdDOAt+PBvPAXqW8O4Ej1
w/DrjxTL3SV84EQ9uJ9gLzdkUx3rFtzk0KcTkHSgm/NtD6P5Qsvv9/JEZyRrt1os
EzXc8IUF0kccXUEmCiB24yt0JeAQfOtuKyhXp1JLOOrh1KO9k5vPKuNCB8wcDhIz
cKnoOLzGzDYfI7GPqfIO3lTv0UconKrr6RXNnGK8kFJ4G8JAgw7l/nV1yLMlr6OK
rve3wHlu1Mmmw4xFOdqU9ljsyxBaEGhGTdeAFj4HMbsWTsIHIR/scJ6dM/XyrzC1
tatk26rMYKTzwaWr16VHSJZur0dye6+u7VLrmKd47u32wm2cgLF0ZBAf2/8wbwlJ
lXeRWq1WpKKVS40N8HNSzronPOJJfjalHvVJ+38gvDeLOo0tNuUmVw0Y3h1D76Wt
tFtGISDACiXrxM6ijx6yE4AMQdnA13D8AYW8xV0LMhbIATd36BrnvBW6PpEJZWbx
CLl8U6P27Aocog9Xykc3VTG+yIbwQbaO5yCzZ8/rUVyPOQpvCWkts89j4ce8FG98
di/6NfQ/Wpp2ZhFt97lMLvrXlZYGWZg7eMVSM1twzFDztRjWKewrJkMf3z4M/mff
J/MmsRSR3MoILJCGAvVZLaNodsqfubI5VVc8LuNYtpRk727XvmLvH6mkM2wCJJ1u
5dHPTPeExyoW0kLfHcv7xqQz8YGrL24MF2cseNjzYSM9jCcGTdOlc43c+D2b2HuH
bFm11r1dMmxbkrwDsEze9bNlNvokYgjvdiWejJa2cQFs+IjL5ExV336li7IpZ5Km
vVoFBdtuh0nJ6biCf5Mf0+NtscAhmF5ZZ72z4CpSdQLYb6Vl/JpmYerzBj2/WNMr
ngUI5VhdrK0g7y2j/Tzw1AoN/rhUiY2mtF6YXmXVf4Lee5Vb0ZMG9KBs/RHCaF99
Jj7anVAHty/tZIEzfFl4HIc/vHNbn985oD7ThY+62lgavMWD4+hgHGwZ03p4YAOL
wJk7v/Iy8aSGf3PXa6sZOZXXscUwpIt12+cUprSWLRLnmNozxpDJ59wJoje1zBD6
bpaO/Dlysm2ox7eLiw69/8YSOvgjJqPKt6U/Ou70YwAPvhl/A3YS2GYF+wMN8eEe
VsQdKXKnYRleCWdqUaIscHB2bMA1t4XBVsnK8rxG/w6urVidSZT5tuxAEHA85YK2
0DYt8X4rJnnc+QlsHgQlw/6uWMFTqdPfKbj0n5Pt09hFG1aXE0xkYDb3RhE68qfY
ItjVabL/WqgLgiePlnvTQoKYjG6YJF3g8l8voeQ8Ct4TXFtzovQxQV8REH/LFQFG
zK6Jd6x+1zXRfD7kfyh0GbDldEGW6mJxfN6qBRf5cbwA96ekMEg9gL3+iTwijktj
iUhoTas9zeezMcj2glyP14pWudDI4bz5nE1sIr2+YRFp1GCZ7QZXQ2N/7QCpXOGr
VVvESr9aCehu4Sy7iUavNvLIlqB7LONSQVUjCdWaT/LYXtYpRmQJqyGKsJeDaRNg
mNi9r75WXETZyVNyBdX0xBG7At0rFbxnFi234BmFLtNVWsUMRckLILuK5/j9OE7y
XCBJ7zQgBt7iMaVafYLxqOyKAONqCPLzApBEbCtZZpdhg6KMecM2XTiyeI/0EjdM
v+B5C47Cu3oTCxw3ust9wN9ssRQhW7pSbYQ9AbiP3JTTuwWVBNI0weNTR+JO70F7
gii/YukNPmxrejh8FpcFKLZ01/HwTqaE0ojIYvibZ7xqwNNUaGmSvl2AQc4yTWGO
kjcSSATF6pw+Y+tJPjOQneVHJ/SyjhoqY+L2Nx9VXnCvXYkOxcNfrBAb8Hx8m+pF
x9peNnuIl7YL3PKv6YGzSyOI/tx4F1Huao81NvRz9zMdmQqDhnoGMRC4b8jE3+3G
0MTKSZOfpX9diqZMGaFzK5OgTBE2LdOmtDmUVHZ/LMv8SVvqbYyI/OmBQ04kKVlG
TzkQT/vmyv95N+xp5/qnA7bof7Uk1r8B9IhnW+WscC6vvTGeprEbpNQCGQOwExkb
LZJbHa1EeBpQmfjUxmHzJ5PyIssRmUdXRKiRSsCOGKD6szqsV02g6vTdcTnVjXey
8FqKFQ3ZUeYP5aG5JnCOyPpsLZmhrsnew89u1M6CjL5kJ/RZ/fesgxdMzy+1dfjA
yMjK9LWu102yyTt/+9w2xF3wjNQ7Jm+wjqjo2nqoUzOdTbnt9w0yR/Njdek4cD1s
8Exn75R72yI/cagjTBW8Hxw20C92wm6a5JYB9KY7e792VR+jU6gYl+rpBYK6YdQm
PJkHwCR173pEbxlT0CeIrMhCpiL9puDNq1RkfSJdsXlqdfY+DqznPmV4DE82Sx9+
PPR5NPftSRmQ4t27SfDA3RU1Mm2CxWyQ5R73fF1zneEvfcCa0u7dMTpaGaJMMNQM
rvwTQLZMsSeGWisPyHK5UI/3aFJ7LrvBDaKyVN1CJ3OL7bi6jyI31CUGIfpDFp2/
bIXiuiDr2TnKVWqu/PiFmWjdb5HDvofmC4XZRNBUE/1jjhNgHMdEQ3IjdmVrA0e5
0Y4qidiglfGj5wXRdggAu7v3Q4clkIOIjhQT/ussaI2cnghqxe4RpN2wStsB9mKu
ItLHRwKXM0fetyx5I3OQh3OMMjwW7nT1z+b9hoY4gIHy3BmbLlbBGBboJuRXmm1I
QCueibNQ2BqcEL20i2C/RyyA5HzKOdQ057Icbs36tW8cufuuiojxIY6XhI+IJxK0
tS7AdsenYIF29fYJcuX/sSywqkQ/XeFOkHq69CgLY9FlddGEcHjiuJnhbGUaJa+N
+/dWvdcmLEwcQZNPA8UCOr4sSW/mvspAe5ErKZLQYf1HQdUsrXD5pwenvPQlvKhh
1ZNlluEMDYkNvzBQh6xDBOKb1Wwh8SJACwxXzgYxNpBmtuFxG3TY7WNXZ0fHGH/T
YPVeS/Wq2cbNKzTn77fPXKj0k6tDi+Eg0wgXN/7ESaghXyCi4+brPHxxPdRATYQX
Z13+hMRNiZXT/k3Zpijw3ZvV0sfW/PSY/C4MAG4wpOByXUXWRGAUZrCzLvVoeRtS
U0wxVk0Q/gtoL12mFN+IW7oJTa+MvEcq+PL0Zw6xxrvwHrSIG6znCzVPFIiMxJCL
yb15HBAtrbOn1hEvA4uODceke9TMsKN+RRZBrHjkd3jVTV6Un3InEhZRJSIy2EzH
Hf8wdiqGgdq3y+XFtBJ1McG+5w8gDBLJyXXJX5JntxpKsMGJnNA1c6sLtcrdggLZ
rGUp64FPKhjtpwv0MZKsuNQamO82OU71wRMsWsb6j7XFNaC/prLRPO3dfYt54zl3
ywlzsTZHXFBSNsYlQfoHmPeW0ubWoJhTIPJDauNB+nxMto4fy7BfxUQwYfxtLyFN
kzrvT7Fu7Mq6TUCYV0OPdXaqD8Wsj7kfHS+Nthu+K2gbyixh5OrxZIJnX/GhUp+6
9XT+GQVGeB+BbNpANhF7CHFsm1mlJCEdPfM9Zkp4sIIAoXOXQOaFdK7f7ayd9vJm
iM/DlfKM47b93+yVhBDjKvuaa7Dyrm8e3RBS6TkpPfMhVZNfotmQtoC3cAoaSZMZ
rmHBBW7VfJrs0PQuGsptRwVBM2A62PDDAbg4FXG3Txon6d/We+q00xSgC3gl9x+v
EJcYoKrAxCzIy+3gQ8jP41+YUU2zybh1Rm4vTUhoIgtuzRcrSF/i97iU49LJTwHW
zXc5EKb4iMVv0lAPWuKtFy6iMivRaoVggcipKB3GWpsyKjWmMQyi3YOj09ZRJDFE
aTc5R35nEwREw4/w3BBcX4D5HRjiXdB94RcO7Vqp34tJnDv/Ncj+81wqJSyj/Y2p
aD98yBY1gFKgAaVd5jtegpxmBqRIzvfMUXsP7F81FwbJzmymoicPr61t5uevSV8t
BOznhtGJV5d9LosZgSMb0mWUoSFurdwTKOBLEMRIIl1MRKfIRsBlV5ayXSXgxzKP
2Nn8mwP13bwP8cxGXPtvLuywEAaDsCgLmdrQHFLqCKeMP7jRLOwSW5q/kz0Qou/C
VnKC5d4SjcyLy/qP+/M91OwhbAmEZOuqjX3tNnRlcuXkcs7hFaA4BqIsTfRL5wXa
6BNWNm3ErYiZxtz4a/EHAT01pu4olRJKHp3rgkXr6N8wjb9tjwX5us0AISOZGvkB
GHZugfcQkIlJXpiEhUhB9f27PPQqoXbF98ba7j8mNMQney2iIkseAJ//Gnqh/5qG
ybBnm4QzlHm9prdnuF5PHHIVsN4khUclnau8/3OfsFgZF3RJy/U/UcmCQbgeNb2C
LVdaMwvCftTTLNY4Th58drFJwQxFGOM7G4TCc45FIPthsr6OaiV1F14uYpDFGpZb
NpAjr5cylAB/kr/YcEGvyBKchWnMEc+wH2nn4P74/ULQSLq26/NC6+Np5zVxHVc2
8j/MeoiyaR+RDyYypbi6RdWoXtuj7Kq8FbdVR1VuAGGukyPdVA4Qq4asufcyXgBC
8GqQpAVfF4yUuO8EnHZ8OvxrZ8JfunlSAakIAJM5fPZQb9OfCxJfVsm9p2z+QaeB
bG1M2mC3leAktJ5A5cW2LDbk7AiSOtTYNENd9M4k1HQfZPEUeTStSoK7KwGk3U4b
KbCOKM/yNcFjzvG0hY+MY8V+MkoqIAPwZ5eW/OevcpaQopO6L77QbwubkE73eyQZ
moW8Vf6itkWAKMrrsYdONg258DpiWlRZQqnKhS2n+VKicRGNNWdbFHJzpwHGycmm
C+UAF3zF1Z9vX0nMgwV6Q8r9xAz69uUZjD20ytp5W3YjfBG+BOtZp2ii2bs2PQS7
CutPARVBBHx7UdlIfkmo5IYGRmq/2yu797DjRx2WC3ORc68h6nRV36gtFV+qCt6r
6MpoQvdSfH61roh9boWrODGMpjDeT21iZSCTvtEt2fk+NPbl4v62T9dcwHA22Wdv
dy1s81fS4vw5v/5ubq9zrC9kBvG4yVYCuFoKZhGo1ohQonUMFy7LVOawRpzxMa+T
S15Wvq90vwVjnd8IZIjYD7TyxMjYwECIC0Mnj9CPKCUEdTwBROFDjgINlIDWWRMH
0rneSPFgjNRlejFOgoDq0/xiveOCvrSteKJMQB+A3vxKxRuEKISv7G+/pbuIAy7C
ieDv8bQ0jhmN4VBkQ4qz/QCsUeO5VNeGw3qsx9sYamugP1DUlQCQ5lUr2TrFJPfe
gQG61ZhYsDKBxHdb0w4TPRIHg3QFMxcYcHilCmatFvRclNPM8EebTAKSEmV9I5si
0bmLGwA+6nw68fQ+lzOJSgtPz5VHuvtWHCnyD7Edty1kmVJwWPY207GMaCThVaFp
Yo8YFuIcXeOCR/046IzuWR6y7ykyfes9xxwubTHL5d25CsqJD94PO3MWNKskVc/p
GHbgkX+ZrldnZgV+8k06936PDI4zUGzWB7yoV7anjICe4k400kwShSkf1sOi8Ze3
8oQxwJqN20Xpilgp4yhrnKRvKKE3YGd00lUiciH95wbR2TNUTbV6g5syMigigcAy
TUDqXwc6wi52LAx9h+gAbtIt67tP1MAyHdoaHSqRoTb2rOd128jePpNH/AVOOFMk
BYwtGYwPXDQtsXSpOsvN8uQZuv8f+BjRSUiXSY7szHZWXYDmxtqRuLY9xivgDd7O
dbL0mdsQ7+79DDY0KzR/B1CsqS7+u2hU8dfnRSq1JVFZ3umoHe4zBgcFgUMIN0a0
Ja3rcjFIyVUiphGbRAk9iZbrxJBmy/F/HcVXtTO4YDk2AiBMYLP07GCF5eqR72Nb
8Ny6GVrgG9UaErAFqp+pT7+boYm+TrPHC0/oTTRP/AhXy7xTkS2vjCIao8OUObLW
tQIkGFq51JrIJ82DwIkQNlGI0SvcbJrXUTpVFB8+j7eAJOGerr6unKEinJqrZxeO
CRS3Atiptcnppk5oAiU14gohekiNqBQ3jX/+aabT2O8nj6r+E2d38gPeK6+IYacm
9D8jOXaZwlARTcpBToa9SRBvLkaNwL821bl4QLvlXa7MrLF535VSm9IGo2NdtuLd
qeRYPHYRT/f35JyXppq4KMdc/lzO7nxOo/ekeeb4UxCENM9cogX4DFw7icJfaJZG
UYIGNWZHwJw3van3Uysv59XYiAWuWqOGGyvx4y5mMdkg9lxinRmS2gtS3S5G1AS/
C5OLjQGyCn2+8NXeSrebVmdyG12vk8MQdlcW+xV/UUiJjHs/9f4DJ2BHrZ5e3D0K
wuLPY9cyjYkhhw/fgMmmF8Eg+9bSMKZeU+Wl2SwznjIcaWZuemUHtNaROfWa7DDa
FpK1qnHO1RB6Gp6PcpXFXRUQyfUG5RvO5iOBE9Za520N/cejWoENyXTFpPxNrYv3
gV4xNweO/oa6DoJA0gtF9529BR7fp6eeINuzwpEbBiydxtpmLqdcUWWuX8pTc6Ub
VwP9AWUh+fayVi3ds2O/4wCmBAjidtkS5m8DqEneqMbjwrXBHh/ioUbcjUErc/fr
QHG3E39QWlDbGCok/9YZU3Sq9QQdfK1fYUsxIA3QyeC1V4YrS3JM0Mr0bE0biB6J
T+w3mlQWLxEe60s/I/u54f6/7yHDcgIbbCrkv1vlhffi0Lei2zzMdkosFLwZs9In
FTNgcBVBx37ydIK8dfqIzzlKB8eUhxchEZHuqgYN/NihfRPYslREmG41E7s6GM1I
ZH6+HOH3OXZXSWeFrrAZT/8TdpcDIg/ASB9KUp14bSR8ogwGAHOpkvsi5AmL5ELe
PraL/9ZZLWm5xW+YatUoLdby6L9xj2FvEnHGQWKA8prlfJ9bz4zkEaxtf2xUf+8r
7jtB8nN6gmQ0vEvJ8N/+IpVawgeyGHLoNzqnOyQthbhfGKaTYf/xANxCEpD6cPzI
MKa1NnFKAO5qubaCVdZ2GZl3FMMlypaYKPm7GN/z4hpoabKtTmz+Wphi9WNJYz9n
O7oC1T2Df55VGoDZF4NZLMzwFQdEASDN/YVCvOFyX1XkXGRM1WRB49+pM8ah5B/D
kTYuvizS0a3NLs7Z6Gm6uHLVSl05JSmNaK4IZvb0k4J59A9IMcsdsCb8kiHY3JZN
u9gWNJZRecyey+5Ie9xFH/T2ErrPs2ccWex6fnwZxctuUAzAV9WXxxvy4J0lGLZA
tNDPQni2yKI7CkMDngnrapDQUgbkw6tfNBiZbclPud8JFNkvJFrfvXiC1o7YvaBm
9Gnl7Uc1nRmv8n5SzDil8phJwRSkyJmySto6g/3SMv6WvacIF5iCjL4cY/h5UrKu
EJSGaVwNPHp53xAub6FTC7qp9u0rTHesOofOTNwMNyredxWyg8eTIkL7lZySFddk
jQHBt8rxwKHjCx8RWTHK/Q5OxETaZd7A4ZBviz1OVA514zIEWxqgcjEewZd+LScD
9qEX/is9m/64Ckah5i6yuDX+AuJF6L+FRUiwcoKAAhJMLD081OzXkkX+ElpUdpRd
HVgNTZZ0+kQJud38WcwFgpkLY8XbLQUYYV1kk2B3YjG5aJqB6zUt4BAEqmOpuzoA
NilWC8uAxdaitglzkagRwT5imxAEumSC4bMlQDuv1Ttl9yX88y9bXwKsVGAGgrdu
/CclWHXplZcKe2WwyVZlbNtQ+zlMkmQkarRe2flkYYtdZ7Th9BwIvNpqqZyJgS7p
yEKq/RKpee+RPDgzl2buQWVkXpXQIagQ9+DMJwgBa3lF7oA3n/BuVUaLuTxa5o9j
mrUqNjNe7oTw5hMfyPNjTOmhtZTNy91iDCUNfEnjj3v6CF7eExn16LB5D28L9n6n
OUm5ix95e/C8PheSj71oab0Ly3xdh36V8ZlVJX9IOdEptSfoIr/uLe563jXEOd6j
UIRccG9MsBYSWWnUCyl20ZEI+6QiTvzuOlA97YFIQ4MXVptvEgeBiytlNHiCIbEE
cVBu9S/o8h7RQX1Giyft5mz5CmUg3jbGpSObwezBIF3gqUISZGrDHx1fAtYPEzfZ
QACTRDfeYazL5mnkpjnbyDhH3HXZf+G8qpH3ONhl4w/zb1UqGLqHYjz82pC9eJFG
j0yaDbXimysLfzM/bZR7QtoGxbXNDkVhqn0JJ1LPANKmor0lYhlQYRu8a8Nqe9il
gA75wpfh5t6fsBq/1MK35KeN3phaQVDfat+U2al9O+ZXIzAWi7+n2CtUUUALIXQV
3Pi324F3Of9Wu4lqDVKq3G+3MPer4DSSCAr1JKwxt+6OgHnVTiZnwbx5cEnGTt/t
79k2FkTW8SgiMNsk7h/rF7DMGLo5tC0Tr2Tqq+vjx+WKj7gfx5/wsXsPnJhPdU4T
dS9G3O9YHwrFvs1adthUUFEHX45pPP5lqWgIdxImCffcu3r9jFH54kactg74aG6p
mJ4vTcmfBzVtYhUeDnjvs1uJwS0muvyfUg3+0PuHbYoX//wUB7nhMI5p9lI6cVhK
rC7LmhGfK6DeSnHoU8BMSVCq7ch3xZa3TFYi09i34+Lzh4vsp+NxFiuNwrCuAF/t
s0+nQbSeqq1APnmsXvMtBWuc80lsgUL8L8uWaKbVIgk96u2gQwBVy8ba+kB7OL8r
QoeB7XTXjaUxhey1WzdZJ0YXj8LBylaVIAkVRysGQ6eJEwJ6ZPl9qWPNP1BfBzB3
IsDvUxfMiWTFLBug9f5dsxk9GJ8qJiMthZIT3VPCMh57Jmvdq/yKlcubspXcHIfD
h9HL3EMirathVly9+YM6QJNYwki4HN1t9LwYiUwVI8SuCKQVk9w278PLISyUxDPy
NK8c/E8/bOMrQONmxcyFLUK7cTVtE4gVYxAvkT4X7a9nbwArQvrBlweexGQdbavV
mesEW8HefegorxozheMTb1fb2gWCfhjjyUbgmlsPfBpd5V8nC+/epxknT8J5oZBs
1/94hxEy4mMh7/iK1gE/Ssd53bHFt5kFtMqu5VWnoEiNLylWOPwpZL10mn8VI2+n
jVFL8xer0dQUk+DzFq0fotZO231DRgc9NJk3eIfrgs0rrYQ3XR4u7zvNMjE8jXu3
7gDxHKYRjGwX8kzUKjmudiXdxZteuV4UWCUH20qW+2fwuAQn1ljjBZYumwaoWz7s
Zr1aXwAlktxPcL88AiIe+LT+8XmArL6UulIgswpu6BtnTdold/K/zseeegA+2kYt
Y0/gZpTXeKEv8Z34RdM8/Va/223hjnvKLHRoRvyO0Z4JN3JX5uzS0uJYBWOJEmql
1+JIirakaBvxluKVlX1ajGCJ1jTkIe0y9hbzTdRFNCKmIbfdNwbXwkflLGYIunzF
T3pjQXHOF2mJzwZaftlCqBlykId+QzSG2MWveCO7LvTiMvitSLI2+UdR+saSPZjW
Pm7+2qzKAi99tqnwgyFoHyv5p6g+XJMIBcDyZ6ZlyEEhMTPqjnV7EFiTeM5gWLj5
TBfNBiuDN2YcksFnNh6b37+XvsKXGpKbOLW1c6nSb8Lk90dbkNbP33HxaoQC2rZX
sVic/vIs/wddiLwCKK6kIN41Do/plt7KVsaPtCXRysYUtFOgU+uXFcIT+2DIafWZ
6jTqB8dBlPWAY0KOCfOnPyelwhB0lgjSxdO3GwivgvKzUVf0Vt3Bn9ktCSqsZQcX
8IpUevULQHnpFyDnm34gICav3LEQ2ztqOS2MrZC/ve3oIpmkzMZ5tQ+XGxVSvbuP
9i0bnp+7CzfTFhQWVdHh+erv1v7tNaZtgpSEbYQQVJoH+vUUh5rikxZ+GtrYrR/7
IEdcKAjsAJs2IjaTK0Y92bwjJav/YSxRwNscgtNhNPFivDtiTVkMU1mYjKi7tFW3
LYH5YyHmEmySEWR5ZATB3ySdYDfxsA2gvXu4v4ruGhkc2w3hye4T2yncmf7iTe5i
Svac2kSICz/5UkA/cfpDAfk+Fom3AZ4/8oSI9VY6ylj3Aq22tqmqRn0VZ9M49QRE
I6Pa92ShXA6e4J38ZWgowIbxardNuF1c9oalH24SVCTp/7/e4VQZ8cdaPiyNgjb9
jfOFycTxig1x3LBskaB4eNCpXfCJrGtYUEBLGlkOsay+FQ9EFAKT29ADuYlAdi5M
EY+lrwj2LYyk6JBJ6RErkH+ztfT2+YHfKo3JSBF19JRyQogRD5z2s2J0ZbheQc1J
ow+RasXquqmlZT/fX2tokopIaHVM7aVrlFNPtGv8rpg47Itl+6Oqdk2NfM0nEtjn
lVWnutxZRQbn+aok6fAoyWgZjSRrJW9FLE8JGssKq55EVxiswiKWX5kZBWMORYDm
2cuqLEHkM3/waOQippspH5ItRMI4fNnjvyJGQ4dGT/HcO/weYEjtJvPfcic88LXN
qrQN2CTgChTrH2RVhpBcwoJBrsJ3fW9bH7b5o3f8HoaFusk5YdQQ5KB+KUe4jonp
5dv+4o23f4rMNNpXNiwp9Udw46W+Mdl92bB96cGhIkOmZoXbp9zjtm+YQQegukZW
v6XwqqBSADU3f0yX6t0qpKgFwOdNvsw904Up7aYplmzdWYxryEqkCosZyPXJbV+U
9P37j5pPPeVsW9DCQnMaDAUuAreSBqEi4XPZ/9kfaT0f2RtwmL6ytNEY/XoEh0gx
k7lkm6i6zxnBeWOV1OB46iI1Pc+6WVf9BaZrlsz8+lR46BhMmsis/3IjZWo2RIGy
ZZBPhiI63E0eU9bVw+BmVBoX5Oh74Syz2UVwIPbE8nDoWTHKYtcl+DzGFvSyHQ7x
KMfXhl6pIAac93N47tJp7fuOnh4NKrRAm6/0iFtYkX+yIHk0YaIFUiZZw2RLXqCa
1pAtUeuaaK3F0m+mOpagczMDr3gcnH0Ksf+XOuDKc9AhKv2rUgZ8T/X02uYFyi/u
YvhrXir7rhd/sPHuNEoA+5+UT4OUY9GDXv2rxYfcrEqkd+adCXsOPUliOpCH/LTj
W7HojvFa+twc3BZz/bbQHmts/W+AgjwJ1GqW5qOd5z9XodWMn7BQ5yo5kzWtDiUV
u8Mfn0CIDI1BmMHyiSX5a3GbT04sq8sdDbwnGQVO2rAAo6EutRvDTzvsYq3oGqle
03KG6vX5e3ZiYldhF65ObZ8rDpAPc+oC9LpxmzKae2m6BdfQ66qCnJBzJr4YysKN
Z+aGvono78RQFr2QPSkWxAo7LAuqguUtu0SIMUqXf6S0D9Qkr6nW0+jElO5sJJmR
TuzVuOsvqTVuqq4SqZfyN3Vmaj7LeR5NM0Cqe9GbYJshllIxJLgSDi41/fDcUDkR
kBwY00hXP1G+Qx7rJRuJHk3TzhjdvA+5fyzcqItgwCHUutYoLWEVg8PBQJop5JUg
oSpL5bLvTbIlBDpN/x23oFYsGG+Lt660x37W5zpXKks3KDw0qton6jmoQMCMx2hc
E0WccSO1yWjcuKcIPImYn913cz6H1Jb+X94dBm9hiD3uBXQCCtwbTnQjJB2ZcAi9
guiENVFl7FVca1mDZtdbeTMfz00Q2jBZEoA43/Ycp5ab0oomK1qG7dWsVvGYSUTx
WkcvTgMkoX0MEmvLewxQ4NIUQrN0Hf9RpZK2ADJRvvK/lRRFUAPHNi0bFlOaHyx1
MI0eDdM+n0CdV1Xxdrwq+7ZFi5/FrNLJ1T5/Xc1mloeeuZIGMBxUnmmTQhtgjbMG
XpITjPZhx5Asz0E+WM6FyNyVKgnRu+/maXOHVbvZv4qkrV8NT90EyPhYUVt7C1rp
3hytpuda58QcFFFz13UOGgpTzKHPFrLzW99J2SQ5W160H1NyaFKss5w3pIBAr4OA
n0fzWc+VkVcjN6XyizMqxMGi4QnHKNKllFnGhhKa9LJ6T+ViS5zwMpU4yoL1jtJ0
RQhtnbG5UgK9CnZ7R9aNCC9dbkoLx9qVHWDPqn19fA2qWAfoo5Ukx0BoCbQ+2pSu
ocPBz8nq7ooaXRWD6RZINCq5B/h4bD5T534bePT8dBbp8YI6KfBhWOhEeBhRwicg
ft/g8iGWSeAyBn1zzmHRZAmhcPv/+CI+hesdVs0EwT1N76e6DI5i7SmtUAbWpZPk
hYsuhJv8pMpi12yeZWLWlT89qwHo5wjbnGAPefU6w0mpf61TInPFUYcWt6I7N8GD
iWW17AEtF6UktUGDgeqEWp+EieqTSsm4MZduirPyAikgV49+TJKKUdtxdCGY68BY
OKFwJ/YrU+6P7jxibNTCRbz9kHKuDKCxXuSq9M/zgmObZjpUhZVpFQHaitBZ/ej1
TeMX9crHt3aujQewHdZkJPKHj64FFcdI60XAxaTYVAGP+Xir56SVwQqfPao5eXHE
XA0rLFjMhXNdzDOuutppekcaUHa2wi5aPsbvISrcRbV7RIZPE2qyb9/tkb5S+AFR
KcgwXzusVgkogYLn6rFUtBpFTbLAx1e2D5XZty+WD3mNBUExFi/jOm7sE8wZ0xIE
FiDFrdEsiAUPZi5fd9J4wGe7lXxJiOKVmqkzvr/cU7Eimmz3ZvTtAmwU/CwcGf2L
4oM8nZU0QneS1z0qyzQfj/xHYko9w8Hqh0ouAWu+LXI3VA3gq3KigCzsIE2FVGtB
pT00hrrwPH2GedAMqrAYg+McFqjVz3beI4mg8ysBiPsqZcxoAub7hBDyQxxceUHi
Hoc7ESrS5BrYgzSNPvW8tj133APjTPqyVsYkCh1799olM5KyVBTyCxxlKvtiZyPH
0j+SywGMYNAeE4GDcmvlMcs9YHcSjKNSzrD/o8MA+87ED3QXVU8BGZ7K5CHcwsdg
FA9NNjVuQ7dUWAq3SqHrQWZk5yGUoS1PPOWy1XT/X9MCEUG6UeYs8RasE1beUIXm
F/MCP6ti6d2I6dsYrDgS/7r56KJkD0zNiGtO/OZOsIHSrgRIhc6ZmThhOlT7+yxS
LC989qOSl06aM/b+t/FX74fNSwk1YLmjSvSWsTsYINaQQRhn3ohGDSZrnryP8jAD
/6RCKbK7lW6fo9BElYlod2womik4VPHfxlw/Rn2NciG1iyNQU5DOK82SH3iYNzZe
hVKa5fr1zHAZsKQkPxpdzUS6h+hmvFLM2TIfI7tp+QfzugHRUj4q4Wg3BPpBc7A0
Gtj5YMMbU6Z+XyYAiMJEpnAgCFdRfUuKgjJqclWgD1KleqayCft+3ElP6IPkRWSD
+pITY9TrV0Rk8Ti3fgJYrc9eSE5zegBE4EK7AmEQefKlo5VY7f/7s0udg3D/n38K
6O/W5cel8HUhcVbm3YJ0Iwz8Bp039p6YIyRHo3bLaHEqFRq1TQeekTnOWgZiZ2rj
Jc/K/Gi0n6Yt9aSQAMI+u4uajV90ExYObIeuupxRyw8JDRKuEPHHMR+y8LaQZJvc
TtHorPamDAHXJTHhl2ECw8SUE/egswSqCxpyU30WWxhYrGb400wDNu4a4i+/PrnL
x3ReAoZPs6BNjA0C/mLMoWbUxlvs6CAJGbsMEpvA2YntCmBPwyjyIf+H4InBWnl1
oGzkfqytqXqHjwLr8PKMU74zllbGSIJquQpPJGuFqe7X5UTVHvUmCtuLiNhQy1oW
EpAUpZ7tv8wSch7wThXnfcNKs83DxfLhms3Muu3ZElx7ZCSzIISF3fiUruQ7m84p
JYYpMIqYF+mg5bAziT4T2nomgPDBK0lBMj3lmCEGMhFq8QEnGkWSxiuxWxj+qfKN
3utqrDrljg+byqxrqByqBSNp/kSEmoeYZkVA3mCPS2O6Z2YSmZcEeZtRQGNgNLhp
hUkl+4b1pVOxzAgn4Dj1GCNgKDmGsoYZ6ffrH8LIqo0fY9jLLuZk7TDNQ3S1b51k
4ejmhhPxsosJ0T5uOWTd+4xIyCeSIq413Xn5waLA50XZQJvpHieiacWL/N8dlPwW
TBCZ2TdQgRno3xS3vlJBwfgLV7p/UZQBn0QsHH7OK0IT/BVsOoFPs9br05WDB6ZY
8PwU7i1GK6R6IzwvpbAEV2W/bmLyfmGOAchosuNc0xEsKt1tbcjum4whIYuweb7m
RkNKwv+9OI+DLwzxZusX6zuDCsxAkA9O+/Yivepp6HzOVgXZ+qOdcenaYCFNTBsJ
y/pqRi7vJLFAGfj+AP+NBVYUu0gLdTAkPqrqproV4Q+j8bNas7czKJMyrYkByvIc
irPaKZ3nPurElNXruL0mcET0d/w5kAgJJneIp8hkFZlUc6Is36zk3CziZYG9FfZj
5pQy4HADMX/xg9wYFCIqgj1AeqVR86Xm8e0vPyCCkBsjN2gLcvY/a6VBKOIxgPax
eFN78HWXWmzIF86T5mWlCLCjdLpzBJ46OTI3LQ+nYLNaCikxyFiUeZN4vv/Wdvzt
oaVBBK1o+krYJbH5HBRl1bV1V3rcvl/gmnhYnu9HW3oAumu90cbMcUVpWDoDevCn
IyLdlL7Gwlj9nbabHhnDgHm6gwx2t8akXd/deXSUjGL/rKqdvM6LQVsyTZ+OFwTJ
YqXC/UAiFB1O9eBUd0oA0OTOtHTQVbivhdYHwq1IUAkO1e9VhTsZazhd5fLHc+6C
BBKpyn2cqH6s+AVFPDQuxTxXg40xaflElVbGnN9DvcEaLsnTE2yoSw2dWXyzBgAV
kwoio7DyyGlVTsuLw+dH0v+HXToBxbrxkx/6YXcc+QfdbhKrEwqPElGt5MYg8909
7PunQH/P588JtpgmTjnNaoA7PsSNhnv9RVi6G6GCgDIjOPh0dZ5jjeHTebTyLQkX
piFBNQKRDScvUhnNQi15HywGp522v+4qWqbTE/J/i7upUYGSRkX8JEnLjr9gtzJC
rJ5ANF5CHUD2UCYmca3eyRd7vUV5N4DNt3SX0Kjg/KcGOn928kedosDrUuMuzNaT
gYFJwTzilH2yZcupK1K/VHI4+iwelFAkVvRhz2VZFYhEyHEv768DZ7GWZfIXIR7V
C/o4yNL4lsQIiJm+PmkKEjhE6RZBFzxj6mt242s4jH/aEney9x8+9ik/09zJtEro
ZjgilVwGQ3z9jYY0/DXDpmvX9kihE8m5FiE84gFq/uq9wyL1vwHw/fH68RYtB8OL
x4VpEyFRRn/99EOBVkWkyZ1VODUrJtrHy28gzJAwnoBJhOw7oZ5WDBkjMAkNjjjX
U5AMQq+HaOEyL4vrY8542YlBiGMMNeX9tdcRcLhh4c65n7l4fq2bk6DDsFegT+3z
eOWMwGA5HSRj72GiisEtn27lE5g1ZiC0/VD4Vg4X9Ecpe4OkhiwXB+EJw9VKU205
fRb686pP4HXGIEi0adZO0MnroqMcw1ymowSzjHKojZfXdvT4XorohIqqPz4088ZJ
MTVgkZhfvle8tvEC6RtKeXRP3eCK6R1KYhtIT5FBtiVoaQjYVRudJHUCe1rEy4YM
CLkzaEc2drwY3yKkZneUBTmRDqYLUF9gm+7g8Fvv4DhqHketfjOhxnjSm2OLa2Qb
7mqs1pAC6/8diwKiWh7MN1xTgF7ypTkpaVuxXTUyZ74N8hub5qo331b1IACllcAx
sBFAsFdbm3OXR2JyiP84KNxt6qQADegWQu0svw5Tjc8lZWKfaOT8O6js3yDiYD3m
QnL2SpSvxUo6qgxHHdRaVbExXMlyyRQUK6AfWl7s4yuCGsaIR56VgLdVrU2joo88
uzdTJwjpQ4s+7hP+TS+0VhvijYsiNWBnP6zDlTmOg7OlZudGLZF1vv2bBULrclkK
8FXTsigKgbzWlWf4eYHbJbuWqR5bHBzrUwBRaRzUG1Sy7dkKkGMa3vzhIYr6Mf0v
ngtGyu62GmlaASRP/AMlxBUnHGUGVbtiQM5cfIxq3hp/nmP1mF8JZNYlxc5zdyCp
4uncXmOYCA6SnjQEt1JQpM0wEvLiGzXLuYluqWHPHr0T+3y0gv2NXAShKNSyO9h1
+lEWfF00q3Qv6WLOKWNdbo2gJbV6vWhGGO+3g1Wb52OkfUwUSbAJ7yQ4tznufazh
AuZ8JJRO3g0CMSedz5gcphrsmoud+fs5IW1HVrFhXD/ZHYj/Fq9XoB2Ysiugec0y
RViSxVEimQBrDyztSJLcKuaNZbiFPZf3jBKKmGhxS1+ZYFeAFIBKttFS6E4E4anH
fPckrw8lb6HKdg2HBV0ysktSRaa7zjxfnITUjTLHf/Rxm0Ep2e7R3nOCMCisb5Mf
Hoh0USJEd3GEIkCTZPva2AunZN4axPScFQk9gxzafb/2Y6hGm3BMub5Vly2lXceo
oUNCcYiTMNKLwNe8HkcDBfodXnNkHpyxOCRrptSbjKNqRNTvmr3+27fsKmfr004E
iEyPpBKEhFmMRGIWazlbZHzUvAMVRTpx3NfNL0s+lfjDRIoQgBYeIhOUcAoxA4Ja
AzawWHKno+cCUrB27S7zxuRCDO3327Hrp7QW6+ydOfxwbNRtb2CRvFzv2Juzv3qm
6nEYn5sP0MMDsC8VWouVtAn0yP2jzSTy0VCIA2SH1fz94HxBe5Zcq7B9k3v3okm+
uaI12+vTW/aZySDBv0hWpchf5dDyHXLHOwSamR3jfZSsPm60RSffJh71EyEtI6RN
0iIsTcpjKJzQIx/+7ZWCH86wujviL/ECWachhqXASyBDczobGmcSqWjcDNpbHZqI
fZlIM8qXg9vndAhl7ZPNmFuqG9AMg7dHHqPwc+diAq8nkfYpTRjab1P+u7HqN11V
LYe5+QWZnjTxE2xgnsIyq7wcmn2UrKA1y1bmiZNUzw6jH+opv/l5G6Ox07M9+mMK
Gl9JT+Lyxc2tJFMJIOQQ+WXmYcEDQJVvUekbR3Sctj8uzslYlkcd2bbtKX3yzeYn
7korn7R+8rXqpGguR3j3rdlvKOs5rcunx+ZW2EINW8xqNLRC1HwPT75e/CKq4l4N
IuKXpCTx116ontR9W+azmknLyNH+p0F57eMLoHa23vfjyjRRFPdcaU3oZcAq0+UA
3N727hJJf4UglHF0xRKD2Zd4lQOknAnJWlUPNpQewnMWwkuETJhxkjK5C+Fd8jFg
yNi0So67FFsC1cN/seM73y4YEwBORKyKP6JnCXkfr0Jm469yIYw1aWIw3f9JQP1g
BNqs/do58t7k/MKPXlVCBga3/0Du1zDM9s18V8N0d8427fn867qY+iGWlicw288N
Bp56oYbC9IF8l/1C0364Za1kXAKhR5xam1brBQfgiXrpqumcGvEtfIkTbHDkuSyf
nQIXmj/uWqWI2TNnRZOz77Fhcaf46UhInYU9FzY/vGtTQgqz/kYMvLo09ciMYn43
UPasQpiBMkraF+Uo/MWQQgz9kfsX1OFVO5fb6SZqGfuqnNL0PZyFfpE4gnC6N6k3
2iyGDK5V7FQ3ywqiTh/yUQFQR+u8wTjM7oLLJLX9mpJq/xz8IlmSKdb+uzNS5MhL
hThwjIgcI+Kqhy60eDxrI1DTh+vsC0c+mq9OvpIf/QXQMrNGCyeJ0oRlhgJQpcDt
3Q65q0R02W0NYtJH1bE6wnltqB47iO/nyrzhoVG5j41I79Z6ooBiDga9xYGk5hxQ
n2rmhgtSucetic0AdhI9DkvRdpgPcY3csJV06WVahLz4zRjdx+3Ut3bOXj9UeJXn
gYI3IqJxLCPIzrSdk6siI6OJ1Y4XofhQBkReCfpZxTRfTSpKbqAzaFobWk55pgj1
SbiXCq7lvnhh15bIN09mDEq/MVpvm8JNMIJ+gTGZSoIO+HSLKoDeeWZyMmAwNgT1
7m9wgY+QQ0+Bhxc/vHO8taqYBYNct0FXQcgyaS4BEMvXZeG6Xsq5fFQIO+2AMqj5
Yj80WYJDB3dEw3qxncjsqJnHLpbI0h9/0V1xv2pxjB9zayulMaeDXat4x9ppxaTn
IKUfDSQkuiaDwY9mr8jrZvgVQcJwVBZeDUk0r2TStNWhySK1iXjmnANjIaFYdVMr
8L8POCOLDauFRLsulI8gDEl2syS0Z5kck2v673wI9NWbQkZZMWV/wEsebJJlJgIa
oUtk7Ly2k8RsXhk+5VpaShb8jkyJ/b3NYblBEqGPEsHckLI3ikG0c+2UYxaxPlUV
shTdnanYcOJawT4a8eFdRb6k6PG2bumMd4mZLHq794KRFXacmKTnBB7BxdmHwp/p
kJEzpsKX+KtyKIRvJ0yjKtRPKMD4VzLI5IED74nSkOtXGuuEGyir6Q4L5aEp12wk
FP+4qsolhueLtygegb3i5ICqKLZnpmq8bMbuITNuUQKzqZJ29zlUvGU0HL9ue2HR
Bf0LivhNUFzyk/VbTmen8Ah3ypCAR8XmPkPUQ7PSC8eBoqn9fE7yrnvSMAk0k04B
Em9oHelsTri7l6ihdvoDLs+lAF0VM0RD7Qo+OJ0urTodaGmQN2p5/VuZDCPoZoDS
7HIAgErh6J7WYvRCbk4xvZwaq2gGDIl8xmC0gpnNiVk2BiShXWUKXC3tN2qcBMqn
VX0lZrs6CDvhoLuR0MWzgcMhIG1VeSwwKQGwsU+xMvUDLFQLvoA259WWrefjeWkt
m/hUvTOkjLU3HVOtFZmeIB1+q4YQPq8yQeF6LYGUdScLFZM2a36Mex3tZohAQ7uU
fuHZH1V20y7YvkHjUNSAqOmuZZOmhDtEWh+si09WuVRVXmXXZSa1dn5G7Kyp2Vn/
1GF8QesH2xABu3/tpIUjxXCjYriOTXktFKGlAzt4PjyLsxPQZNlgFtCOwRImgvRj
n+GOBYfZQUCUy0/n2P0d1qIsfoa2sVgNzNDpmrYSNgnCZ+lYuS+YVSHFTe2uDLnr
ocXuoMDoI7HHP+ZvryCxkDFAoSgYXeRxquMaHGtIE5fCXyDzPCjC7rQY9q5QNcCN
UH/Z+Y/kBtPXEz0v1q5DqlknuTPt36fL1UWeUcZO5j+yIvVRSpJfhBemZ7hMpyaZ
aCAG7Me8oQyXRiJs+jiu0XwL40bfhajG2UgKIAZ5DDYppLmGr/RuwwwIV0bDlnGz
i+JIxhZ5wcbR4HjQy3ZP+nZB/r5WpXW3eIi0NRs1wUqZRTLDe35/JAuiapT1+qoQ
/M93c65Lsn3v2g6gJ9DqJHnrF2kL6aobaSIZN+ByXDEU7BWF5IZK8ZheWO6HIPiO
i4+BTgoUlMbZRTrRUYX2sNwvE63kWs9/O2Dr9C7PbY3kR/eJkyv+XaqyHOmq7bfL
f+PhqmykRt38djZRTbXz87JaMYbLBLDcHDhBAht4wmz7QrDlhE/3n80RIq3AgBOr
pqT2v9n1WWqpMxa1Gv4nevpPHmNLIQ/fINWgzR3bgtIQugRhYX576WNm1wtjMqwl
7SRAggRBtmM4rwHd+C8Pz0TVRWX45mn9QvZVT1xEH+plhOPxbYwo6vBt1VceWGW+
pgSv9TGYfZS0jxv+J102GKOgChIMACkYE6wGDROwjXVo95JjbEG4USMQo78cfH4v
BGBxQnImYobuiT7Ef+b+zx9WSCRmGKFtuaHjYSWVjMqNiwp6maup8uQLEVg3ol6Y
K2Wa7OSjrbDBn439quGdKOKV10RB6s5BBeitPJMpWqWKQGhI0TSS7NkxbaXm0K4G
07v/vfeBxfkcXkWFkWOgiQsLf0d1c5qonDRURS8Ltp0iCt3eCjQjtyI55loHzqa/
wY21ihw5C1+FmtpqE6YaK7OkNj7ownA87lgwIy1Snm0WbuXqn9KHh+N1TzRWLD/Q
vZMMBNhg/mFRXJPlgYTyMDgqvLdX4Ba2sQgv5KXWMyti/k62EFHcJY9Yp8U8f3bH
lJ4RJmglrQ9kdpFLaWumgbx2lQ01UlBJIEEVNQWUUvsScM9D5B/iEwtFGDp3/EAl
7vmliOX4mRCNgsb1HArhKxYgN+WZ9IpdlL5t15eX8rloaLrjBFu9mkWbpjm25UMU
dqmmbcAbNuKVpCf24jPJYIklmmryzFttKyeGfpMSg1HW2z2B2VrpKgX0VmcjgaAa
z4GOrDoTTQOIuWSjarDstnoZ18h8xEosPOHYy9VKLjvRAWWxt6xW9I3vzg0fKPxL
ur+YGMz/2RmVVLDqJg9rfBl3ATKHdZO/z+a5dAx1vs4gwheewbBbLTQgz9DkmcV/
/Zge6EbPq3lHczi871WnKkdK7DvcvbPrmPPlPLyYqCpjCmxyAqiZP9pLH9niTJOy
WCdVdswSdtC8hsU/+tQxhwC6hwsFLh+XeuLmH4N6xQd1VUhuXJvsk9awUzj2EENv
G9Q4Ap2TmmTC7pOEkdiRWqXoTsuU2SQakJVS+PNkZDgfRegMXeGUtfy6UC6ofHgo
p4zBBKotgLa/JAxnkQh/UStoYezMGdVxlUGD7jbN2oIwmnoBfKhNLCie6T6jLq2D
OzZZLY/LtgoJcaEXa8FSTUoguoqL1FpicEFG/YFjBjckaKiWHTXceywBs22Dp20v
Tq5ajn13mOV5NvZlup9thd60KVXazLlbhmplvdtQ8r/6tZ1poQNjXiQJ+RWUytr9
IURSh6SEJrVcpmjolRxhS8GvIc1GwYmibuiQ96QZWq7ES4VOsnqvA5l/6e2izErw
aX4J0ZGuh8VOPHVJgiths9ccI90XjcjJFUVba62Yc6F7mUejZgkzb4B2uy+mwBa1
lA0m44UFiwKm7hVEccvSWIoTWffFOywt33rEG6aECZZA77E3pnI7Qpc7M1RfearJ
5KZlFQPuEQwmLBboCKgZL5cDNOcVqfMB7wOpCEcN4OIpxJfcp7CNp6hutJ7aBv7m
rEs+6sSUMnUxIVn9mjURuENecDep2GydImx2RZupa0fclGYjM2YE2Q2PppUpowM7
nxd2eFrdtM282QlMN6O84HG54qTwy3fLSTs1hR0xsTHUzT1nOuoK0hHLVqu4F4Lt
LwKs9kh+vf+76Ko1Y4X5esGDD/lDc7Jj96bAx4DFe83IMjFyx1uXHAUGVpYkOIz0
zPr1l/nhwzaXFmKx81OLWMYQnlIzxNJDNwS31drA6XH2bbIrOWxKuGYcTSqOdNPC
fHY0xoOuHUqTahXwoPsO94pL08uFfZ0Uw3c4PRgHMlk8G4bh47pP9qD6qqA3QviP
tSrIDahyx3mqMEm9aII68EG45a+IpxZ9RpUmX4L2nUSso6ogGANmyakbvIxwfF0n
WoFwyQsRSfoSZEBPoVOazywjLrxtZIxQbB5+BI9+1dxvTuk/lrJoDei7AACFn7Cu
Tse+37BnWAjX/IrAHdJ9Z31qu3BcN9nebIAQEZ3sndv/FF6HyKg6qD00QjoSKD0N
YDwnO0LbuIrTfW2PfldlV5P83FQR56lcMswYP3JHPdzK1ROwJY/W/iEAyiDpaS/Z
zw/M8705NxsqMIJ/PLohZZSKspBOtPQMHzbX/LM3A4/1rfpHqI55/WTjI8ZOXyMx
vpzuELbdTsQEq36kdzWm57F8jTsjpT320+GfFiHQRaw+Kcr81G3gOggR17HjYz/Y
B3M8SI9+EI5XQ9fJ9miyRVny5a0kVwSZOB2Mo+GoGcBX7ZaDWvrd3udvc/IdOFGG
6lZ8/HDrfq2DVL2SCQF+GAhEGunnDKGEqQq7GIS5ua5tb1cOeUKf45tAJJQ3sBn/
OuOSUvfifGYmVadl4RsMXTkZUGZi1CoryHf/NLZ1nAi4Dd+NK5BqeKrsuapUk/Vv
Iun5VhTZZ3X49cAWQYC8jyNG6unW6ek0a1jBr565DyDVHftaJH3+JDhdV1iYXEcG
NciZYPbveVTCetVrwyZ8qOIOm6Rhq6YAq0AsGDVP4aslnQWtoJvR+9M2tlci09M/
a7SCKr88q8CMscBYrGv3uQi8+jBlPhmv3XzEsVtLNHDePJMdi+I/gAoipmEEpJrG
ycNdSS73eCO5Dd7yGOghumhUFBWkMbWNEAPe/r+0pPLl577YTVWKB69tc/iZuK7G
QfSGgYF5i5rhXpGdmybXwCjeiHYjUkR+crf1MWnVx8rnnwZkwGkrtCclMle7e764
Mc+FO9/pieCUr1lFuCo6eBckgjPdLX88xTuc4muWm2PsoAOzPZPUuazUwo0bB24k
tQk1vMuITp+lZWN+D6nCk0yJ/SSukAeJaVh4sSZ6L9ejVbk9Q0VMr+X17L95AGh8
eaWUBj4xw6ll4Z4DzCzI3tdoGf4pDvMm9CSjhTlcft8wYfcH3cmMI6FWT6jnCPI4
ufjHspq3VnQjqbzP4cC93kroeeSeZ5QzI6BoPQix5vt8x5EaytVgqhyGbRc+spfD
3yfyG1mP7kFarYybLWV27d8bTk/SSCzYyiRRua8bssfDmsMs5bKcr6zV9sFcfn6H
722WQyYhNhZk5PLMVZF9uVJ4Ovyl+9Z6kcBLqZ9FOHVrsG55mW7wELri9G5lFRzN
lamFGEB1C8cvZSQRNmAgr2KCzBapc9aIVB46kDr4vtLYcU6eSWtyZ6QMNcVbA3RZ
HL3c6vkEX56cCMlLeFQX65XUttpdCkEOjRQ4BYTmqXm8i6tPJT5AVYrNjPrlKqR8
p/+aBf6nKN1OhSdvz2uz6V8qMkIGVy/qBSWvGQxzUzrCAA+oaY1PhgpPyYPjFBlY
zRaH1mqPyG32GgF8mZ30YkAmC+haAa2qZt7DACRVrMuATHywPGAmgpEoGJFY19wo
V6kDS246Csvp7mvABGDBkhQyRyq/6+Eq5XbrVYnUePzgO3qJh/FmxTU6MuW/I+vE
oavUActRZLj0LTqWWMoAHIQ6U5+PwwR5NSTS3wPs5XZ4s3fdzX3pGflXP10wMDxH
X9Qx/gUGKIIFcOpA1N5yOtU5nfbBl/DXpuarlhbNGWd5BF/+WyEHTbN7Y/9ERIk9
832KZnzISNzjiHL+bMrgYgu+ljYrpk2v2Sm8uPkW6sXP6tkrkLLnxRxzwvATzVuA
yUOoL9kL8JqnsfnIaMgAz2fysK2XTKxuWrAQQ2IDD+oCOQclRAZA4g1e9fe9MGC6
icNtYh/mQVKLNc65WsBiaFUpzKg1ccd3gs2j+RWw/CStFTEUT6+ZK3LNkYCnIOv6
ZO43vpqVry7PHakaFGVdFqznylrX0pYiRyAiA4TrgnmXlOQLVX6TPMwnpTaVkqYG
6GidGn6QHcvnkdqQerWqPvPSGw+CTasJcvpuAKA3Enzd/BeFms78I9JITZb4KvQw
XBLH4q1jFh0aL7ivPLzktwSjmRkrmE8FZ4KBYlrCAK0wEKe/fIBcsjmt9eLA23BY
o/0rm//bk77vyhfL4mdpkZqDGIk1bgXzVvAnpWGFqPfrhA+Xjdrxsh/mlBQ7WP1h
LaRYDSE6EJvm6ZZoiZFjt6QN9WMxkHFugtnNS05ObuA+tkRup8s2ER1GWC0qwLWz
+8OlyI5mebPzSJufSwDjO6lDOu27ey5ykQwOURAQK0ePQlV8yosTzk7AL3Q4Nlh6
lkZrah6CryrZ413HCNzKQPonAondL+LqNa3qvPB0deQvecCzXAz2ijuBgpGMD+dv
VoVOCMd/HYbB9BJ/ponW8JHbiq2CTUwu1ff830jmXbhVxYoiBIwmZ7bQk+Q6381D
4iO9xYAVYWLD/XWoabDI4V35YiN9FVDz4Tl/yFa3lorKZvMdy799vW3tg5VdYIXc
uCrzUPwV9Em2qGixIGHKnoVyzU2+S30TL5YpdzIbqi+fgdxBJMNxpZ6iqQwquz7A
wn0bw/plQcRVG20Zblr67sJ/vyJL5vej9I1aB2lYijXOAurINX354upxtHn05cM3
YGLB15VwMA6GeIoa6oBXWEErBt9W3M6LcEljm3zZaDPrcOIwXoQUsORh1LtSNb5i
rsDjMqS3qUI+yR7CMyyjhY8L7ybWIFyK4ujLQjnfHiq/S4D4oK9vn87I/ZDkZEBy
dpYDjHUky9rRmZjDFudaVSYcsIuEAjqPdwK7g7bdkuCyPTWaSfvcPzdtORGt0Zig
vvT976lUOdtvUH52YPsmT9V6oxZYAbKHyX+yvT/RxSBKvnVtGsxRGKt9UK9FvxU4
URyN9MFIR4rnseNyySUb4c5V0zRASUgbKF9cvZRMq5mLeQvb5o8ExEzXWNA8Ad9I
AtmHNwJ+1zM0oXX34/1BQ9g2Z+/BLFXl2rdXBnJdVydGQVGT0/6nykAmEiIFjnxQ
4J93WnF6Bc+EaF2AXNBk78SmJ4VSkXdK1PtoSA3QMPKDQVJa4jM2sfRu9nN5ibPw
OG7REhscd1ulKnnvd3yEkHK8TkbgaEmWSIVY0qYJ7lFHHNb0IHVTwR5KLuGOg1U9
Z4kVwiwiD3D135X/djekijVW5NAadtsma1Z86ThlkIVKoX1TaXgqy9b0VaDTDO87
pUMTQXz+3BkoUyA4W19kWcbguDTcMaOvP017mzKJsWSUnk3Did1nRnupZxtKN9Rw
n0DcRvQ1yYiZJXDV2iTH58dT1vboWYin1+p4fS4rmjeFHP7RkHsu9f4xnXNBWrkr
A+SsGo+n8+H7Wq1fwlMRGMbeuq9N4f2jmV3WUX5V/+2Vq82X0EkBl8NmN/vQoY+t
KGTKEAm8hbFkDYESOzXLBjRE6oBV/TzHZptUq1oHzfbueHzSGir+VWEsX0z8OadY
9IImYhfeBoD3CNLBusSe6FHCpXrUN4KBP4dh/wiCw4BFem0JkSZUHcgIbilh4dnC
HrHfwk3vJCE3a0WPDQKWoPAqzsrGYlpghOz3TBpDZitD25SZkNuGvhbBnZCb0lrU
rlNdZAG/2l6L6HnDbLI9PYIKjN7KmyZHq4Garo0tBif3NaxFvnbtuG4Bmdjc2jXl
Eb6fYMSuG5DBLLcRFV/DkZQoAyGaWNQwiE9+w2PP8kDFU9yPd/Z2/Iu129o05ZrO
typbtFhujKEuJRHPRc0pHB0EtyGLaX3C3Gk+ltzMrUgJoic7KRGMHDyK4052Hlu0
sS4ihCO6PlVOGF0eMILi566jRZnBf0xyRdLDMzzOW5sA/1tMXG62mY0ypMYNtL6T
WWKIEVyoKy903PXZ9UPeMDikGskBAVGHmKd7Qu+/FMRd2zfYRG3defUhttyFhnTV
ZKOjoUj4/G9Y6GuGk+ssPo8oSL6pw6UFbvtbILQ7zPYPWb81F9AlwVEB71M5MbSC
Wjew8qIs/uZKaV8anERwwzL4GYe7lekb/WsD77yDVfPKh9+1zqvtfr3pNw4KpP4h
sUzXbqMQq052TDzgQ+Hens9DHKpxEC5hE2ZmLVE7XhSyyjbh7N+kgt9ZPq9X+YCl
QxBNoOMQolUEfqLTkbAvDVxSVjTr9A8u4xjto+ebVqGH/x9/3CVqJ932gx/6lzyJ
br0a5sEgMy859yJkWJqbtvZg3QJvsFJ/jlA12LJ9mAMagsj/muwTeEulyu11cvLN
Eit371Do5sQO4QGTd2YhRG10BWm+lMb+Q+K1PpsLKMLUB8JuQppLZfIIQUmR8eem
McLh3DJa5V34A+gjDrGyqfiqtMoTcj6l7CkY9tHBbQ6bqmGgiOKsEmBEB7BBXMSE
YCS05/IvG3qHgJ+5Rceul7N1B9LO+wygdCZ2L1ssOxRQ98x2rifC5wI3QPyGuPVp
TxWODx7ewsssmT0NMtKrrL3MiENbh/8kMd7UAIF+Zua2Ub9NBiR8jkn9Q5pX/Kob
3Fwu3v+dUPXl0UUCDS78MDOMDOsEpblWrYMkeKqg8fks3A/qR8Tf+dcn5PJIyhin
sfnFN8z7VkGiI+D9aTzM+q8spKxWS8QkZOGVX9tmPy0KIMX7HfRaNVtRxIZy3lRi
epe471yDQrR6FEYR3w642JCn/QF64zmJ4a9ZfOdNC2JHJizc4EwmIb0Nwt000ILH
MYAAT2AeytUa6rvUFXJJp29q2N7AZN8WMCVGkLgD2GsPds/+i586pxBpUKBc2KEs
Mrt6mS7ynvxQ9bedi7AOgggJaR1dsnEosfTUQ+/vSKwK7jIiNXAc9S7rm1+hWdjn
FzFLQdLXmiuHDhH03x0vzJOJ9Y61YP0nXZXtGQ9MM21pljGDnIAnloLaO7T32G12
2J8PZkcLdkKqCThrKmR/kRYMO7S7wxjVRIc54fgPNNqL53fTkHBxwqZT2kO3Pa6t
hH03GKV2SLFn+68yOxpvE3iSaIYWiNOuE7/9Etl4fbgZue3M3AOhwIqCN8pLhMnP
NswL3i1yfvLwWjrL5R3UBpO/i4gb0NtL4fR3gk8Gzb9V6Y/eA6bi2k0HmHBjzGuQ
I0rxZrTByGFUCxUPuwDrQ5zs3+t0rQmJ3gIGEAtXoWTyJlrLiSVtTVY+2b81G1+8
bu+9pzRRkA7F/cu2VEr/O+V4fRlRD7TDbsxpg8H+kYL3UxR/YmuvCCYyRnHHfayW
B/KWPt1fB0Krp47fM2cE/g6m07iGYVpry/9vpyJ7OwL7qjjReQbqhu/FYYJWjd5P
WPYNx7Vprl3vNNrktsqYPoJ29kVdrsyAdYH5FzdFbdgY0K9xRkJLZKXgxzOshy8R
NGp7BU/dqwWT9/ie1D/aYV64BZBrjWUFUkpG+RWNHND+th3zqGijL05yAgUJaELJ
AeCUmblbej6okHYm4J6Cy6xdUdo/DgigmkiBelFaRU2j7M7Ug/hN90lvs3ecGvMP
QRBBNYcqvZ8Z89W33DxJiCerlbD0Oia4HzzZPf2SvFM0OUHyA3qppON+ZFFIKeXE
nxHLdlSsZuGDVA8/5MFquT4xK34EZ3Lcc+4o1IGPJKisWdL65R29l6Jb1rHCdvKK
9n0pq2nk+PlbsTPiEGFre+jZ0ofbecxtdNbKlK+HhoUFaQJC8Bt3ODpMU1Lpzphe
YOQ3U48iCLNtd2s5qsISTSWSKlHb9Be2mtjMBqPetDQFTkUjyoCgZ9K0d+2I0gDi
lwqfELDiiLftPbnc3mb9IGaYZS/IGGWZtdaEFEARBwXDKA9fE8kXnUNGVQicwBxN
w7LpYr5qp6CyJRzPuCQmkGC0V31/qak3tp+vaxlbzVJugvw5uksOMh1kcmENmlqS
Z0cU3boGX6g8abCl/bSWKQc/FdEx4r/pXolosW1NGAfkGdOJfBM9D90cDE6EAwjm
Q4uBwM80Udrpense3QLboccltFccEQuUY5y3rFlbTo3zx7zoZoJ6YSI3CmE6+NYE
44jpes0HL383oOXaod2S2vnG5eZD/xyBV996yGCvY6L0+9DU2qjhHtPz4XjG1oYa
uIaWcRFekxAXhhmMEsjDoP0LEq+qufZPCLJwEiw/zLOx4iSVh3f7Y1bkJdLYjhG1
fU+d3eLt7+JMqWrX6rB3K3sxoMEYG+rr4HpqBZTlgYsKCtQMd0ARfyl2NLpSxU/X
OveW8WYgUBGjiIWt3cruTAWMSE1mbnRtDT7hwzFOhBoWcXydRdkhVPy1AxTXc9Za
PudH9R7cCpBPlgJrEe15JY6GuariCJqlI2Lm2UcFTRSb+SjFEbwueDYTxzU+0bDb
O7AJIjUKfi5ZnZWzJumIlMhKNOWm6KECIfYoBdc+VF2SEgaj6f9hLJKBgQ/Nx6Mx
F3+6I2AxIszA1OCKBgwpIjSGKnyOR9u9mixM0S0a5lMME4JmK9OJy4qdMwOhmwAh
cWTjwNm2D0uYYMmcYtvUwXK9cSiqm4j+ZPSYmPuqgqpZTuZsNCNUrqZsb8hzotK0
7bua7qG8vEsd0fqMh4UdTHRpX69OKsIUWlsiRi4k2NfBOben0nDTaTENe/NxD2c2
ReaFshVSnR0IzIvtfKvWIgJvzBNeiY5d4i45nuQJkd75dbyKDXGilEiAQIgyuxzQ
dik69FBtYlK/7x5d1RO0L+c/S2hoh2A6DboL702l99OB+R/5jnvr3USUZW/XyRrK
65axUFTcG/kge3U7Z/ZpqErxdQE4u+lbVYIiGsANrS7lbzQjeRuP+OB32ex8G1K6
LyhBzsK1GVUscvLWp1U4BjdKLQitHCZqHO40Se6nL8DwUGWJiupGHeold/Y21fyg
nYH1LTzIQ1sToxki60Iyl+AU5mcdV7zx1RjbFdLdDkETlqgrwyYXpcnw+7OGZcR7
qXTp0JuO32DS1ZQ3lN6K+fxspO2+3rkTMQPG8usSZCmaV7el/xRKWxvddRAHhFJc
G6o7zIsswxTZ5dbR6zYoEiGY9AHFhoAo0MbMjjmGOriWqgjcU+XzvYL3fM+oTYCP
eDzz8+ERfkUbli6jv3JBnYtA+b6GyUA4TD7bQ/2XmL41KaNKQPnMYZmcJINZYpBn
91XEdE8my8U22ah8Ar97xGZRPY83KKNS5PdKxppz3gYejGnp4GfjObwaUaDKytSB
/yWDQjD5TF4q0O3ojo2PR/akQ3u+H+xTeD2AACKbbT4gHxc9uMICEvPK+zQ+3uxy
tEiFbktDWEF+PYodFelj6r4fR2ecSO4tA0afbFQYBZBNr0zYuyudDewnwkkI4quw
KlspTESxhEUvdq/xmLpxjSGDwJEDOqc8UydBRRsOVnedxnrFzFmadjXDjuWH4taC
rQxhDzt5hbRvHu8d8UiGbuOmgyrWgBo9s9jxEBc93YTE4Goh3zaPUEI3HOUIi7bx
Kog80T+oR11ibvDWx7F6AYo3RkcICvW/ZUScDtQFVoMBynySdcVpdFd7UoLAqhrx
XXjMf3uoyTmUOoT1DNYftPdheoceROuRfggCJB4OM85jSnRGevX0Jy6h7h4XBb8x
LSLrwZdCHx4yU7/QL2Vd212ry7UQU3PnuGDbK/QXW61xmDTO9pwYPVq6eKwzRaYB
ED+CVAVYS1Xl/483fCZuuj1l+p1qiKJ0e1Mz1s2MARyyyiKxMYQ3eY9gbaiS2NiV
yhOKBhnwQcyyahk41OqZd84trZoiYDCZwVKmJe46OufT2eRum9l6wR43d3iSmUf5
in59V8D1iQyU+FPKf7YCQ9IwDAQIX4IEXf++FN8yT7TMQkms/O4cRO9Gb2ZyPvHL
koKE7JgEDR+XSsHVciFIMxkPshmi29m8MkV6UoD5/K0OhaBtBdARB259mPNSLJsS
8mwUEFo7q8huuJsGYwZhl8+VkrQakwLo1VHdKJc1wzNsjtUIACEGZHD9QwWvSQBK
HTnHeSDroe5b+DGXD1bnxwa6xAhUd1KGx3sOshEFboobBPuonPgmVGH9huAU7dDU
NHAMD+T/7lMPCbNU/bXePvsHwlqCUCTSEquRaTAjfLZ1wPLkMqNKQ2UIlNvibNuX
wF+ej+qWcz7DNJIDZ7OyE0J1AeloGBNqpreKRKWtACABI2yQmb+JBnD7KEyTTYgc
pZJ7L6LPjZYrr8f9Lj9Ra6rRWJZBbPJkn4y5d9wJ3PnN85b/UOfezuy1iC1DwcBj
EdzX1S4VlCgG4En6jtvPhxj+8FPsdW1aOwivScNeg/6NXq1KxwXqkdLnxVMN3mYx
5s9IjKzSo7MQb/RMvooDvjVh742gBG4u8lQIYhkJsiNq4GvOVZZT2l2vtHftbmsc
SMqDROWKFzoExEdfaiQGQAI9+FtVFD0rPwdDI9359c26SLF2etcl6Nf/BeZqp0qG
EqbvPeBzwCLHV5T1Z1vYg4Tb1foQSk65NR9EHpviByltwfYCf797QN6pdA15PDiH
CVTqnWWXOZDmzpTcoRDKpYvGhBkXyzF3zcgMsOjlHtmqU08uns4wwG3V+6Oo0Wij
d9tPOz1M7ved6cS95hv9LU68gjJV5UlF3RecPTNLESTESWu+ln3Cnbvz5OeWNMvd
TWXA2armVmbbpgzwy4QgQR+sn3V9posPDjXXfxSeg5NC8B5gerQLJQzhWWDJnu6z
uNUekWYFvGOxG/WSJ7Vb6y5HoOeV1iZ1WPG1h9dX6QTTu5csVgeSOt7STO3lwcBB
H87n2/eSzVfDvfxqif8sGHphZnhsuutTxIdFc+Ey/PI7JjiP9rp0bZ7ZmtjTAsQX
qKnRwK4TSp3BTbcJi5Ba798aiN3OTzk0cd+vdMat/Fegrsn3b3H7rNVyy8yQhm1v
wnmraSzaIbnPWSprNE/Rf+9rxf4Bu65J/ZdbJnbO5lMi0E3VuHVA69m0pnvSaqS5
SWfLzq01gXqU2OsAAaDhvX2aKAY3MtQ3IrUKor0dfLk/qi5LJBo1+CvbUT9yWr8Z
V5gt88hc3gQiQnluyGIP5kFO/vpiBsiCTyFNvAsaLgkHVqcZy8nlsGLPrTZSDaxu
VW8EwXx1mbRQ3/D9wkXQsmJLWgi3yHYmzmK0tWGCrbpsoQj7pF7OftMM8ZoEIwhG
t9AlWID+vMjEe7503SJdXgJGv8V+hUzaskwvlgogSTDvT96J0fgIbRC+fxroMxm7
7+chVrKz3+S+4sNfVn6BylkEjmw4e6SCrqqbbg88QZRsvX2JnHhRY/L6o5qLF78v
QVSM9I95i4NRlG82Lm6w1+0qHX2QwwpOP0ZFKcEySnrfIkSkpO5Zp1eRHn+5A+Ze
yZYYI6crgZB582lOysYB7POsFnHrj59CjEZYcDeEttgyRTjyD+C3pY0WbO1PWi04
PFI79vc1dyQiRvAovMn9hbcyKzZZLRV98F33iIE+Gqi62CDUx521Ur+Rf1JAtgUT
EF/rnfgnU1mUYunKTdEr0AqkQVk6AQPGUXofAB8DQVCu9JG/mc80rYRZgchLg0nB
pX6ngSo8kGXtVwpNYuOX1mtDZ+DlF3xzop0pfwTZiW1PdCYs2h7KoP/eN9qXcLZc
7kYSUa2l8gNXBlV69imKxUeifYM4HleyGYrclHdXXfTHTh+pEGKqYVHWQP3e0m+I
pCbFYmDove9y751R4/EQf13mxMbGTMKri8pRsx32DjODiO9m7+qKXUPf5/LMMH2t
xgT8ESp7mqKLo/nvZ6NGEJNpSi+ip0v9gxIOfxIStXQWWb8gyOdZSI0qXAgYQcJb
I/p9vXaIMRbauNokjIrM9iiLAOY3JEXqKu+9w1vvP59BV8+L91E4fZ5gTuwicF1p
b1DakIX0u3hOloNC8YedCATP4xSKGw227Rr3cQt5CafTkdQiHKowqfxzMPUKpll8
jTJ0Ikmd4QTvd7KN8GAP/y0PY4tQu47IOR5LCBuXvK5ix2nRHqBpJPX9OPrpeBpa
HWl2r2h13+u8x6nXkpIhvt/XZvBP7sP8NnqFSEwmL2jbpJWmiQc9f/xA24vhBYU0
lcsO+SKQJFBsviwwFruUma1gsy8TXgoWB3dvd0JuzkMju5SQOF2hq0zpNfNcxXg9
baHLb8zizXqZYDSfnAww+PGAhv5Ovkg15FXR49igvarcoVIuSq2ZP5p5zxNNklqW
n/VB3TuRvd6GQHy8RfxeIkFFcD/cL7RR5lZWGadLBs6ZPbY6OvrKwXc2w+lFEg8C
ygeUDNB2L+0LCSsMmUm4laSDJfsSaxmmm3O+06LPhiXI30u7bs/Ae7/axfY3IEIa
UMegj7WtB+H3MoP/LGmqS/hiGS7uwklhi4r78ib6O5jchMH5em93Jq3V1S6FN0eE
zZw6ablkzQscy6ijJnmtTrWHwZyKwBTzjBFapIvn2MPeRaSMjAf33gQp0TPIU7l+
fHRTMtUAx+O/gyzVd1Y871TPFgV7BXVHY2yTMFU5NvrMRw19ycDBjiPCdx7w8Nf8
/0Pvd/ebcxUsezfWYNm+tgh/LaB3RbNSQvaR6LKKgXbq77nfrVOTqZHjsIpT0NQw
/PPNtp1wkQUXJvDXlakokG1dvrhsy+ubsaHnu9urhZ31yT2Z3m9HvLv9gNi2yb+W
U/OtO2BH+IYP2VASbrRBtzAEdKCSuxUQCXK9RYSzO2NTqyzWc9zMbsEgP54WqMSw
EMAPLAnzMzkMWvH33A24uJoofYfljLjefFGxIyhxvAeZQwG2qF/M6S2c9nWHndVC
D2x0UaumYvG0+2GHGVpmcbBG3Gajhq8L5Izar75s0e3k6Ux24c+svlI3VCC1/+B0
wuW+dlvJW2+gMLm/IftTxg5oqILKfd+ytULmjUW67nYPoOAaTViGTZ2ih5Zraa6b
mHqMYRjCxeT+7w+oSsJY9d2GccDGI0jAjhfeQOTq5SU+iK4NRR0SQHOGsCI2LUDw
0RsVzO23XGn51sKHRKW98AXxlQJ88KMSiXh9p2Swg5JklueqUHgME/HpjSvLwEzK
+0/4B3zoN/GF1+Yea1o372WTBpgloObkcKTTHXj2QF3pG2bOU/Xo3l+dR9fLSCy/
UMcxJv+P5Atlz12PqfzGenbSa2sxwgQuEkqoS3u835YjerY24mv/2N4i4K87JheM
X+ZNwSUZXsCOaX/i1bud6SuHLsTquMPE8geoYExOFFmjlYK3nOAF7paOsEm719Cg
MwHftxu1/jHAECl36pZfhJRbYZr+uc63UReLGrsH6dE9z7hokGIoMjB9E0JAglc8
mbxGSzfHhRLSqsHj53YaqJQXXQ/WSMyXh4hTOHD6C8A1O+CjuonA0CkkovqcpFGC
LhYhHjdaCgPDz0p9BDYlNM9sBmXeq9Y/W6m+1fKiBALXImPcGtLAVF7/Bp7lSCtC
AjbF1/sCgBGAiRHRO0ygJwEjub7PZilHDybz1LBVIyP1HGTcBVskbGgi5crBV1/1
Yh6QZU/GV4fEfXmRJEfOwTHOXnkgM4SsqE0RI/0XjLFZwhYIZl5WsTsWHOHcNj3h
ZOeOF1EoTJRunpRDzxKjJpKm19MRX03dWReow3+AY4LGHlgYi8KqFRF8GzH7LIdV
KlwDwKQDZU9lPOPwtAcZNHnOH5DoK/9sLdjzwcG0qN6EaflQ64V07z/ePeaiT+9g
7jMAxknp3y80v37d/KVGx0BAJfswhYQbsEz1RLy6cmsCnzayeJ/hrJ+Cmf/1NnQJ
Buf74jGvwkXfHR7fdK7RnNDokEiu5QDC7TN/uTLm9gJhmI5EiC4kY8K8xIaN/qI3
H4QInKtHoHko0UbsOW5gV5GUq0011EnXx3v+yp2vmc/hTZmUfRxgsNTg3fq3vfBq
0vxhEbNsdInogGm0iVyeBYGHIWpYGIyuJNlK6Za1fvRqT3AOAWdl4Ll6IqkrIMAq
+NQEOby3aVA5GAg5EmaxbqdEB3Hayi7kUWp1X6Ev7jjN24CLNO2G333l71AROSDT
6Hk40bNVvID7WTlJHLb1x3NmsRMgQC89nt0D4IYe5RxSxtgBoOTiRilaHnF6LLew
U6famKyrBongvTwO3BzL4YH7p7UoxPrfP+QdkJ9BLi2Zb5ZfskvTYeak63qwIOw6
6FRZ3KSUhlqcONA1G6uh60C86aOO785u4gmfdQQeLLfYQJ7kJQUb6RgJZAweDrWP
J1MGvyECgKZbvhoXJ6CmmfuwdUTG1/RVSgOrCOqR3UoPn/E3yMCW5Y9ompjUkYUg
qadFn3ozhBjOBBdtucL1elSV0qKo9bbHhVnbcI2sRPYx9maXmEyJEr+jKgBo57RB
u77NvlVmR8jPyF/jqTJZyZY/1WCP8aFFRAB9z6SgGrDS+FkD0OapD+EiWAAgoUvE
XHOO0YpYp+c1W3OAynM0IZqmlQfOU8txPnEs0GRx82Y/e81T6tb04nvN5Edyw/KY
xykgGv6vFG7c1o4z0dDMMOgqij3KI9W7gaaIliO5g71VmJh3vFcDM83fYaEajiTR
tRQ351zuo/kib+Fn8ziPDUstp0u5AS0vsGIf5LcW5leZZ1gwa1d1AK/eJ5YI/Z/h
x8zTRyB6j3/z0NkM+OJxVvC38Rjy1v+QW+0e0ngDzwVFagCEYJ23+1/IRiQYgJM6
6c6Idqp47WASUqNxBOXmPnkjYap1cQzl2nfXW4EuK5QVn21ZJVc4OBvy9FbOT61o
u4Ap17xCDdG1i5Zvboa90vhBjZOlXMYJbFi0Y0vZiSdgS8yWuJKhyUxJS3HEfjQW
XHQenir+uM/kXnINOWqiBMfsXw4oyGYmOpg8fmtAQ7pA+dLUzvkK5ydMJW/EtTZe
33aTbg+MI0WdV7oO2yEx0R478z+sBnHhQxcxdIVqbehVIOVg9CQR5rSQMHq13Fcz
WorazHYlDDydCGdNMK7ysLa8GNT8N3XJ2wr1TXLMwnOAnAWB8YcjNfXX0SAXz69p
2DCg5VSOYG2fNqYfuESfDf7CEjPR/1KgJc5UiPlrgKXjKKJ900oAHFPrIiP3tDs4
5rRFGn3Z4Mw7pXYEAjGnogIEbs7xlJB4KAVxOrNxUMkkQxNwvQJ5ijNm86Xv930/
ctubj51QHfC0noXlet5p00hHPH+tfXLvgPJK8jGwg6Vtqb2645ZlqNl/sBgK8LAZ
0y0J1z1sub4X7h1w+yWMRzy6fR5+J4xu9WEiHYFz6x/wBipurBZdT80NiB4mYthT
SjUffsv4B8S/dWAO4Hqo4aiFxGVFHgoY8vltDj5I1p844bHNCx6mtbPXqyXuhErg
c5no/gn9AQXGSVdfiVNlNnSAKFmV2aMED9s76P+e+xK8JTNyU/seah+9PlUaLA3f
o2R1su2Bbaz41/4CRA4DJ1U1gqUeF0GJ187pPiZ0AWS3t6n/mLQg8g8OYTXP+5QR
aVthRgy3pJNLNhLe6uRiQCyYyLG5nYdFezWM1qCGM1p2dxnHgRP2AGjL4PN+BiZy
UwtLEUH8kYBBkr+mG5B6rgGetUDOqAEwYd+7uA+U6sFoQMRQntJs9KYZ+kc5ZNBR
2n8XKoX3YwAjLkhVEYUjBOCrM7NkMfsg6y4JQmCQ7T1ThDRMS9XDw8/FCQlThhQY
qbPKGr94tAzRWbSigtXJyq2nhwONVNII94iAP0WPucDbELp/+acbUTsbyEZdm0gI
VzQjDzZ7gBLOK4we2fcgLdycN/KIckzyE9mSF7KxVNlyb30FzJ5G5PTNhAGfOz1z
02AbeAwrVnK8w7pENXzlJ9A+b9bWAiABhbRYwQEEcm12PKPzQOxfI+EutLQz1jIM
clgHGiP2jv5vAz3gWQunq9DHdomG56fdsrpP399khy1tHvipU2No+p5kHCioMmBv
EHgppeMIOEOSPQup8MkdZZZ9pR5sbjs1jAuuczT3AI3yj1vmn3++JnVImd4J/yZa
pbDzMcW+ysDILJSkG8N/Y2iJfd8QCgw/a/PjWy8rWiMBMlLAEURuuWnrEglt/TQ0
WXDjnTlwWu70UMsAOA7x0HLtKeVi5ZU7NGpYTxAJfNTnTog/Kcu+LIcXX7Zifcb6
EG4p9juyv3bjMRE+ELIkUa8agSLfeVIiO6oADTNV1aHxRvE9aovklevP7LFQmyIH
xksWj00ZCjCKIJ+4Qe+94P+MPhL6lzpPCigcqB5yX1xnnyJiYTe8uX7pZ1VwEfNx
i/2pHuznzt6uoPNElyfFcLijoSUW4AbrkWGhLM3v7ncx523qXsRBknUHEmRXAtX2
NtJOCR3ruS86kmtFAn5Y4E2Lv21w/grlGwO+M4AfBmeYzkHgqYq4Qx/C1MX9tNgY
H0Tz+Vue+Ds/GSG+JO8u3fymwRGOaxKoFaplochCWEAcqDxHdNun1riOf3kHkuDT
uCPRiZmsI/GFWuUtQ1AC05MXn/KVWyRnKew1aY2854gyxPBuIB8StngnWg82p3v8
LJN1IXXZW8Fb0c1+6PeQ0yo5qlydFjNHludipQIJrBbthW6Mp2h3vXWjuHCh7awJ
tx0FrNaJwMLlDDrrv/aAQhx/dnExuE7bDp7GP33xxbMZqq0BwIfSx+nzv5kFdfDo
nQPuR2/u4R/z/LFmd578EPS5gbiMRUCDSch14wximyGe8i4n3+RKM5t8DzXWK3CH
C+bbogkPupZMZhkPTW7YOsKvbDsngeacbesxSsXA/WlIPLPAkgdfdkKPa3dZ7UiS
9XcCKzSJWkE2DIoYdd3Z18ACuySkGSD97JH5whUK8NuNlRx5Hf4cfDZaBb66anf7
6HmZAV/aw/L/VE4JYjy96a3rx59tuE8tfj/ApiY7XAXX6LoB/XiNx6PabMO1QJHY
vDoR37nil5CE0jKvtiCGun06aK8Hd6XK8CZyvH13Fv95FR5laF+mbyPf/PCCDU3D
91ZHV4DHatVk3m92QDiy6GnI1d0fwRhsTp5RU+RRHapOPbe5a3JuRHGnZTlEK9pI
tGTuOj5qFaSnel2FnUp2PEyiN/hboaFK3PCThd4IoiH9qUYWgOJmSsk8GT17jHLJ
Idw09nCHo3T7bMsiUCl6Lfhv/mwGWQt52YU7oxNgscxTbiL4SBycxMDBy/qZx+4M
l2QpkuKQs4Is0JkICfbODG5/HKgUO6XxJWph7M9eHA0pLldPP50KcEHuebdik9HB
SOe4Ik5xavWC7t4fcuqxBZdWzLa3Ytag0BmmNujVCTjVXxgfUylUh8QLA4qBZpcI
se1xlv7w2GZXee1dBGeFTXlyvO4CN5A4HLQMbYSM2n6IjViOf4iGj4DoJqYyO3Mx
Cys+A/1jK9L0mGpCOFQpXkHtOlJl7HoBPYA1ydc3pGYi3JUzgx/r3b7E2fFIOb4S
hNHydjzXCPClHxBSN/ou3bppO/O/rz19DcuaqrBf8XSCfm4CGVw5MwlL6CvsgnyM
jmpktCcYGXCHSGKNv7leQWC8v1zSMP1ZNbWBa0Hjfpprvo/ke5MfdiC+VOVczGVh
zl7gY8FkJ1MHBtOCVGUM7cs5/iJlQEwmZX7g7auuQ3iXE9P0W3mMBFE19afkhdPV
qnENF5VqYdiGs3lOTBLenHN/nsuTfTIi8JSNmwJtMPYwN8YLZBN21CIZoHbam1Oj
oFWWgkSb7v06siwJyYz+ESUz2DNCITLjDxfe5KCLlGYmQYdqYxiZxU58zwYysqmr
57LP2tajOLErHOi/TIj3HUMpZvs/kbrj84ReL2D+ywoaG95latxGaM9g5togQE4N
B2n+hSsiWOrUG/U2hYywUDQ9FuRQwcWzhezFL5+nK8Nx/w5oP5/+VdP8Fr+2YoSH
GfPuadU2N27hfqbNX/gaqMTuRC/dLku9QZkeS7pkBbgw528ieiFtsb1FWkTaD7rB
CxzTF7uGCN/VmduI4MicDPRqsBXDWKI5E6Dp78QxajdyVHOiEi+zT61XcjwXOSn2
ROqTlVGf3VDQvesQRegfReQlft0a27o/ZaBqG4a8o1ukWMR0uTCWTdpz3xi8zZRi
BlmH55LT4RzjILEBBz9dMN0Iqz7zzXEd+eX11HafwCVfedqz1mLxNUrNTbRE/HUU
ghX35P6VMSP7tLmOuNIV/0rYSxWWvWvQnvt0MkO7qyPhWtwRVPLUelyTEteYNJnT
cY2OJnjp06P0s2FgF2DxWe6khTRwJe3YquBufVCMcGHJb8t80COXfg+qZTLZGsD/
6zYEvEcwhUYSARs9cALm0czOGC6wBDZWTlpMgAIwOaUvuwNOnI9aRgorHxEqhpih
wJ3vVZLSTOFJa/yFlH2YVDxHjUKKDll9HglLdHYFz437D9BEtQZ9I0gLlVEPgKpm
fqr0KKFpk7V/L49z/A1fgIa8BodevJbYJeRl9WT3tdpdHptHTFQePepRINFd85Am
sQduQW6fCuSXcdf/GBwu1AD1GFJBVaWNXy4TQiyDOLgtyVJurFkvh+BSoG4FF00j
LhcaVBUl0S49OEBF9mIWQ7BFInH134LMWzs9eo3hEZXSEeBzBb4VmMzttU2E1m0V
hkSusFTPouAHHUy1bfwDtLYmuTwtRjVOuvqwXvOBh4DwMtHNLaDPeV84AAJjtY14
tySYuynU1KCrUFUVuCkW62eZ8ZyutDUH/KmAiLZsqODT4RqdOZ/ZpcQGt4KT4CZR
rP6UoitYZB6Abt8RfLVAiW2cR/It3wc0QyVBS1CceRfc23dbhSK87aBmGx9ZCwwD
VVl0NCbdrOkcsEP3YmgyrvzzfmzX/UtNR7vh7XhQpGHYe25KIHWDgqW+ImzD7UVT
Ofs2qlBeoiNElGQ0QZttW/WeQlxuAtR7DMCX+LHs/SzCr69BnF4kNrGegug8tcP+
SLUql6GzUZgc84TgQ8LsNMfdP6ADApLJIHTRc4eneCbPzM1pTpSMlYVjW2GsIq3q
Rlm3ZVvrFyRUJC3C6SY/pxBs0Ceaf/8lkMfcX52qAYIRR9O7j3RslLnY1frE7Vlc
MzYWXKXBL8t4gZbva2ovF20IVv6xQx5HybbLW2O3BOH69QC0rRKCafQUEbV04q9C
f1suH/U/EOptv443ykAx4yymcrcLwGBPMgimPPUdMcMTQJUMMtsWHSNx4ue/H7Kh
u595Nj9xVhXPpAGcpgGq9KwGjwdwbPjeayKUa+7hBA3PArXUD9Q46uXvDTKLRaoc
ombsgrETWADI/SYTS8pCHmIf9kNIlkbN0mscJwAOEsB/h14CRrSMZztEd45aG0xP
+6v/uAsorq1cQGZxKogvCECZUY52YQ1NStcPFM3/1VVF9aMg5356I6UOb+oukbuV
0MkLIFFqXvR82aOQ/opyLu8Y8Pb0AqwbSShyq2TQBkTctFf+KpkRMXZADfV8sEV3
612IE8aP8t9MULYGYsMeuGP7GTvjOnKCCYIGR2UcvfQA/okiMv4HgubIxsipYtVY
OOVUpE1B0AFOoJaByUBS5CDL/QnXe37gb44DtgE547NfBlLjty02zDxNpJRthRpD
sx+lHmumnE2zX6XeJML3RPwVOGLLfQoM+Es8TnaOJtRiziNMD/ql+O1WjjTKtT0e
ScrNT8lQk3A3PmdMYrOfSUgArCyD5Vif16Yy4ZoS+/z4q0sguLufby43kF1Sh6Ls
KFGmGsjwURaGdkd+3jqgJqJB4+2mNuTafLfBC/+QavZrf7GvrMjLYwnfXk1oyTEG
XiOfej0cU95YKLtFJakhD/7WiNsgnR7Dl2hgOKMHRg16PDJDFHs7kAvHSMRbd26N
Y05P9DfGIn/hUihVYpxm30jusz++gNhLMBsuTe+3eDHWxcrbX0/W40a+JirpMS9R
arw1QDEJX9GibvRiDBzfQopBGnNDC5sRiUEY8QRRIme2IOqsbB+oaEBWvPSOUgy5
WZs3C2YAlKnCmmCJNXBn/QUePVaSStUwaR8dHOtFGS36aHz2UEMkKYPdu+dmmPD7
OheiItR791HmOrQWiJVWa2GQmoNMVbumLiJIWccyTkJz1eAdxTEfFLWzIN8PjJM1
46kP2mStBLCfhY0wjlfcGzqG/CaqCrYw9eb0FFuh5wUhYV3sapVLldnkyV3NA0Sv
GjParyAlwaSV/rxtWNp31nv2d75nd2hmnTE5Alwa3FXseezTZWfNumRI4hQT4M9I
SfVO40XtdmHQ1WOsHo5JQHBHG+NPfNwj+K6QeauULJ7qUjol6/7OIkqC++tfoppD
9hT2SanMwN5KROamQc3G8Z6q0Im2/r0IxfftBzl7lWYOXMkI68ahWK53Qtkln/q8
3O67fky4lRoOAenuDsZOcgwGbgioA6TMQClIoKa52VQziScsZDdIfEFtCbocpDBP
zSp97S19QcFcOlvD1NUbHKTy2C8/KpQs31v8P5Cbp80a96FdDiuH3dGEcNtXGZLM
TY5PM+SAfphfwKpXTH1GR/btkk3xMSYxAlQ6PM2+6Xqp9YI4fyHxazvqxQUxFKmW
9JjuD6WIIm5kXPgM8XfZPPaUxoxt6/yVAar54Njm9AjdaGyWADPDVwdd3IqnNXy9
D8rAMAm6zgfaP2B47VVS4BPAWKmFWyAsjuiH1gy/a7USgWhXdy4ItM+li6hBSIj4
imwC641sGVSYsgYbckgoe3zO8aMcgq5W74iPKrTG2/BquKwK+m80v2j2XH1LcCpX
qTgnTwysGUdxrT2uD/ffySslW+BeXRBYYLiii0XZXSdZWLWHVpUkKiul+x2FwxuC
5+LLYebW6C2/2DzDLV1ZXPhHbUQQ8VTrQH3tay1GKDVQ7pRUTbSQ7L2MCUFtqUhE
HK2fivJ/NvWS6XO1uKicDfmx/U1BYDxV3FAzQ/E7qfCMmTrTn6AjKIL+xqMcp88m
vbCBi8jy3/1FaULQ+r+AGh5Yb5IABAGEIBo2UiyEPbM5Pvg5ld/F2t5LxLoDumgD
6ckcadEOkJL7MRbbHSKML1hC/NBJ6n3sbs9MJRk92SFWSIbjDaPYvMuAgCmyEkxj
zdVYDmj/S6DthGOdUywqoO5mIcmIHoyjhSLjM+6PuAeuSYNiKuMaHxjrtRR9Mh+w
mM75TDNjb9kRjFFFmIvwawD8W8yTfspfeE9FvrDRUCjkiz+JvAtdN6ee8+qJG2Vx
5/u+Fq/nfRzXW4J5Fk8aqzM8b2/Km5iWxc8pLphoB2lA846YJjElL0IMs2OCVq49
Rb+DQk/FuRAN4S8dSL4nyidxBk2kmC7/3har+QiR5HeVwo+ObZMSgEs6azofJp6I
VUtbP/opL0abKUhqnnoli96uBfvHOCQev0o0Gvebkt8bbNTdU65Fi42vu5gmbzKY
dzoAVF/1qyLhKJGQXFPN2abU5Hi1txefi71+zNZgAs+dyXhoTGtXo5HYrYqHWPYk
RiMd2ryZO7r4+lcjFlRw7gwmkbwaIVvUKCSn/uEV9k6Ir5uGnWpIfT9KEKeRfZrr
V19hbm5VmN0F/PQRcW55/k9gZZOL67tj86Evsuuz/hrsE7iarEIhJwpW41tSIFmw
jc0g0JM7/RsdNB61Pk25xaQ1jLG25CVsHs8e4R8JB8lGpsExQtBsr8nri1VFXN/n
6r+z7RIM5qeIjy65vRuIovIgeNi7YwlXDnT2SyEpW1rn9MiI+s1nqPP3jKlzQHos
ZRcIFx5ROmvXiCpFhCMiPEIQvTrGR8/we2J0hBGsBo+CJ+7phsLaCjMe7ypz8xju
3b1anRUJF7JQHGel2Eqie1Jap1fsd/6UnTL9ZU5QW1PbzpprrXH6O0eoengxO1SB
22uYn1DZ2NeuGwua8f0JtF1Dbe6ppExKczKR73/oXomiQprEzt9n1FLbkCnYBE+7
vRto71UD8dMm69M1gKXrdwQLctMpHol0cE/rHa7pIPQ0ZjDh5zaURYIAp5/lu5e5
bKwbrz2eE0oLf4Ola1nCvzSbWOMB7dPHMJdjWQLXQyh1l1GoJdr5zFrdJQMsBkz3
WFv1zM1wMMJLOmaiJV/t1TA9UaIPIbMNw72zKuCS1YnpOethm4UuAoV9m2/yV4/L
J0n2eYkUqIO1rs5DgO7JOs8F6rVXuFZLAbVTERkimvmPGVCFp0Fb+JilQH3MtoMp
KnJk3Il3G9MORwpuOuxpf1apScd6TOxdNH3qUXyw5bftz4HC20biyVaPoLif+2NK
pwS7U86UpgLbnlXXaOZSi39sBba5kvwbonjfombSo/o1fb/qO7Rhv1sN82Cr9Wrp
x36bXHccq6Q00olDO7EYQhqSqi07kCPtHvEfobUyvW5ctvLVeRNUrBvKN4UuNNkH
mY/2S9WbJFXUFyPqmHmTRmn3dj4wp0Z7hD9udbTswVWUpR4BvRBVQUaw9gTvacip
sc5mzn5IKphee7vJeW4+hKhGkXaXu2OoE22kilqcbPkLPPqbmJJA0XrRqU5EtfIP
WTUJ8Tlt6AE2P5FqevRM8rGfCgLkoaabsY56256/pntsttTQwzIbJ3apF4frkhMu
Ks2e2vL5JkyNZHkusDql0VGCZOW+i6CtTCATsrQIlsxeJ0cXlI8bAT4P/wJgbUUP
IjfKMU7s3iuLUQi/GJr2rn6uST41d7063tm+vFP8dz7Vn2Dp0XoG7Vi0TI3QlpTs
FKCfU6XNVRAEEJtIPSj+JZSfjM8WixpdGhr7biLT57yI/8FVW96jVifGZ8sCbDjT
6/ADDqm6/6ITT6fF3jyV9qQPU+OHL5deicgk5CxSrCWMwifsi8+WxjcHJjfOx0n+
2K3csWwOrc/O1LfdMbjmfEI5bckPkpZH4fssnY5oHOa9Fc/1nTYzngreYLJv19eK
36GZHCoJnxn4JvIa3mkAQ5gXJwrnMYdMnPA2/Tw1EoW1Vvo4oia/DpDFpSKgD4KQ
DbIrDlqK9jV128mny3McHWlCYrHAVyHxEWWTTZajfzUfhxQ6r6wyFZHnTrIEevDN
kSPodNSKRKjTBA2wxAdbtecXMxpyfkWqGYTXqt67Jxmc5rFQpR2GCFKP32Jvrv64
u2I7474c3gnD8nSflI8DhU8kXF/SPTNajI0S5CVypujDASeSLXROQHQKE8y1WZ3p
9tl0HTmlH+mWSx7+J94BiVZirEmLST0RerFZ+R0nm4TDW3fRhSoiV6OzuUZaLc6i
axOHVHOO91hp46JEuLqTV4aGzds1q3l5gHfmXGIcLLIZp1qOBYtIYhWTq9dx5YWG
SijM+i0Fx5Ht8obXp9nBlCclqp3fzUbuWJ9+BqvceFVoX7ANEDrAM41uK7NmbFnd
oqgFoFgdjUvRsAoTPaMSxZCgJYv25OXPesk+PiGXV6uBsaFKnXblqrL2sagInAFY
sDx5j4c9R1IPpaUlZSvP10np1XL80hjpzKIyJE9sLaBCr6TiYhE9bouzlKk9Ze7H
4GMOiSIOORCLaiPaFa25ELT98pRd2ctL8UITCNHrGjNTo8hvckVImCnzLIN41gNo
RvfhV294Sh3SIKci8FtgEY7qBSELFwWH0fUqT5xz3d45Ar1N3z8T1hRNQRDSHHnm
y/qP9Br6anWttVM0rPecYvYqSRgobtHrSM8QTUuCfHhORnmmRVy4MFgauVRqnSDv
b7CC0Vc3T5aLAoHe3SCqxmwAVnLaRUwH2F3JfA0VLzVva3/abq9hiKDWSgyTHZ/V
qPMq46RNbLFc1zH061ROwruxXnSSCRbRa25ZwubphKI/mLcQbmJnZ8etg2X86IJR
CGxn4ty65QJIqxPW8KKPJ0GYxJWfBTRQsP3h8n28W20IPnJenhqEHO7vA7YfULMD
dxFrT7fid5mnGXEOgnhbjUjSS2ANTf1yX0b0stxkNLnXZiulwyyeqAAOH10fNLGc
E0ISqD5uioJDypOPwtFdxNRt93Uckf6SLCFLvpwhcHA9FFukYopmSbuiwnHhi6Uz
i8mu9RAvdr5uxguhguYaaYPDZNyT8d3WiYe6pE4mx3Jbx6oXP60QOJCgk9FLO60e
t+7j5DTiUMGW8f+WaDvHfiMW36A9F8PingOAUZRx6yJ65LR7AuMYLoIN5CvwN3jz
9cvnKYs6jaxj6lOvsSoSLdXiARhOXn98eePDR3KX8FmmqkMNRgOq0Ij+y7C5P0Pj
P6zaOTeWxnbxZlSbL9zhznOVxjuuyIy+rkGpXRKFJRZQSJBdSIS4bsmkc0LIr8lZ
EOCxdDUeMSscuWSokkv0yoyLb0kkXjHz8+wJObEc9sj1DiPzc/9ptvHrQQ7RNTX0
MS31MGZ8u874atKjnJgsrfHyZ72G+BFwfaTPqHn7cBnXselfVDk/jMrma5fljXH4
0aCE687rkvJG8b382EhcWjnh+6MAvllX2tjrj889HObk/J3lLP/sKyAZDsFpQhAk
jpWVoC3D/8jt/DGFk/t68Qegh9d8CnSFVjOAXjS7E4TNK5h4PrNWW8X8mfRl4dd6
KxJi7zVbmu7Ohpl8B/BlalpEuvT//k4iKR+WSYs19vjJwilDpuKeN2PmDxNK9D1M
TbkzgnTp5RYEuXoWCF/qXmHPrrJpk6vZ9GKy8jLYIuQu30WDy507UxANts54+MBd
Df596HxocVbm3XHZLP2x/M3DIIrkptgKB2hNvgqVTsaL3Y1OkiLDnT7LTycTu57X
LRnGhiVkYdDwiV1vbIae3VjsJe5Y2tboKGnoJaM/i8ms4Sp3fQUzHAp1rZM0lC23
qnn86imZBhcfKIfUnGAcRvlY2jFM9opXBBLvXcc8H8W2UgDeai5ZwKY8BK/Ld78g
rpN1dlE2VJdtlVQb7/i+AsCWRj4LLOPDryt9FeTeHYJSkWiG0gNfIrJ7nSDmHGdu
cke6/uVh82OFRfal1NUp1trsCFG02VnAyBQPttJDjGb5BgrwECc+CnFtyZjc3T1A
WaI8MAtjTTkmTLh90vt6bmYosHlKLE0RrVlZANuS0wOdSTiJV4zxxJqtgwMlTlFs
yEYBtp8xJyFzQGWbMpkFTRzL74ZwDey6atcRnPKAHDspNDy/HQ37Ui92uPukzlSn
kWVwk/op/0FGCeOx6JfJebl1mBIPCsBJJ7elsyTzmUd3nyJfAyaSg0hm5fuyCz97
WhWxFDXGHr8/6tvCzzP+DqE0frHxYPRLN8x05eBjG+t80jDE1zGwDHDsUoTvXyEX
IElnIZlv0P1XS8x6AM0rPWl7HfSoqeBBsJCpX7AuubTV9jv1T2CG2wzVpQxDx1fg
31ev0NZN4BE/Ds7fJudyKGUOrWbVaDO2AyFEdUNE/9BjhYExWbmxam9CYHGtZjqL
K3Ic+qJxHWrLBgrn8E96xSYj2XTeHNJrJET/ZnJgA9vphACPFwodE930q7Vp4zfp
4YCVqp1IKsZtsPGmmNCJ+rxQ3vSGAVJ+MXoZr8MvnN2gcpipogJnDcQGcfdjh6lS
yNekG5RMcXVqKXxGBVwEZIAQTT122ngqEdyekN06/0n9Y7Ue1MDUvfCxnldbdKYT
K3fFS34XNZgVpwZHW1rKIkStMhODbpSEjPIX1UGl0GImkkJ2EunBH6nKHbXNwwXg
k3u1bnIM/4f1Wi8kstj//gA/IO8/4Hklo0GEbnapturV0NX1XJJxQLXZYzFlNcGN
oDhFCV5cy8g683CdNA1Bgu94HZO/Zbp8qOZExS5ybR9WVqdvDJOZ7UmUb3LXeKok
jGP8PcYRAI8F7qCvRCoQH6OdvgJm1GiD5m1m74jMzZBPnQReMvtnSocGDPU+Tj07
S2F9UrtXiQF8R/U9MgHzDDgr4f1nKxk1a+Slue/qSqUMV7n7U6kB1cOhG3g9szPc
LNu1AJrnnfu4TWFHVue3RB78x3LBSkEPOMig1ap1qKDzqi3UTjjGJ03dgPx8w5bZ
eHYXsajH9MYWwKGy71gLXlQL97ztL2C0bt4pEH9KV3r0/y4w+IhWN2qbZHHvDJDS
GzXrDq4ScnJp33KS8lHdAD7Hi/0cmPiKpNshU7AivVgP4iNwbuSjH4IuwrBqL+HE
ps/ti2JfI7lH0QDT/wR1Ees1m/IgAxE+J+rfz8Y9rELLAvx1sldpR7FLXrK304G+
iCZKgoShWqJj2wZf67XQMYfL0BO+SQgerkNjZgdNQ1FfYiJrLyJ/TNwGufiytXfx
4EAUXUx+pb76ou0M0YJdR9m0rOoTvyktLNwznE+66kNti92KGPy9aeLHRTJXeBEg
WDPT5ssa70sMITmYsQJjDfEGkWNdwQVjAG6njByHQd+PjDqCigReZo2996GbxS55
pFKEhxucj/ny1n5WHasysIPGebvNNevzvu6qGhPQvRtKWG2+9Z5JUx6GLFRXf1Oh
Cj06+TNA5u8EyoxGrxO/SgKpn7d1Tbi2IDM6h75VPkFmnmkt9JJ/rBFc0aIkaSSD
Uedtzw+desnJ2ImxPgPqu8R9v8gSzn5r2N35hYT72bl5aDnthnRGFE1ZOM35PbBB
5LODHyOi7Hddd/iXWMgC0jCUJwiThiXDp7xuCe0lmfc/pI/H8fdq22iWuMc/8IMI
jBCB89cK1A07r6CKocI61WJKS9AB3fj3WWZvylmM2E03tzYuc9wicY+r5Oh7+qrL
27dyBaUsX1n/NhPt/biiXmOKWeIvLdiQaH571a6u/YvwGDDknVusckH1fkn2UbzK
jy3XSYNmhtX/Y8QZ3Kb1IXWRf+MZ0VwL4qcRXfiWi6cJJYz+dqwRuwZYzrb824I8
/+6NTy+1UQJM71Cnqgexa5PSnMBGssRvoHcxt1MxTqhDi7W1LhWOAQFcQhhUsolo
FJkQ3e4w1VYCh0645CsWN4xuvC1TP9kLPkb29+IMHVsFwGPPhiAZG3lnRZjg7I23
xN1dkBlTNk5CJEP7KE1eig1UOKXOJxHicN0Nq0FZzs+2S4XnAwwZsvJoAFY28ANI
UKBY210D1rjOtk9A++tSBv+WP7hcaKm2Pgg3Vktk9xUkKHps/W4KkJl/0TOUBMT7
/2dDvyOJthnv72bh3NeZHySAwQ7wIbHofoJZx7PVgNurnWgF0UdVKr66oW0RAQ9/
4RDWSky5EOr1wUpG/h+vubBmjXumo37UmJgthPzByQa3R9MaSsAmWbqQEtJ9Yxx+
Ky/uOTNx2N4IWJ4/WM1rEm8eA0FCkBnHwBLCeNwScyK1LEbZD79QW9ktFyO5gMLk
xjfAo0S+S896Ka4gSVGfyMKUxWY4TKHb32mzhbLk/qdnnkbbuajl05umDKgM0W/p
+zg0D5jdLgeLDnjzImbOhbjlFVsBKvVzYNXQmf0LalrJBFtVPkaUvTWVIoPEakze
sn6lhkM9i59R5d6wdLfDuWnOX4w9G26pGzRkpxxfxz0zQBKZlfzoLlVxPXbLSAym
o5wCQdIdJXbfdEIAjI/qja8QANImLTDszsmbQ8iEqlddU7L8bcffmK5m7k8ohqFo
TXwA+iHfFCAc9k9KalXG9rCDztdnpjvvQ0D2IeUqDwSbZ9UX1XZoeeIQOklnAvdc
sOJskQMbHcqkKFXtp5XJPaHQjAJjMNFra0K36EYKoRUbXOPZSRRh/kl9nRO6B28n
6PKs0n2S3JMVitSGJ5Gsksx9e5HjOlqdyJ6mjct7gh7NirYjieFkXUJANXsHDG6y
Lw91N8+lPov5/K6OQUE+wFDouirKUmDtx6dcdp4kdm1ZKnYg9QL3WrXOu4wRSvLO
aS2xTLMdFmG7BYi3hZLZHuJQQjWN60W4eGs5M641LeY3ZCOuGxJ9aq6KOOih1aFe
/Q/TJ15CydfXQf4/7dCc2SAC2g8ykufAVLNw6QuszLriwmCJmUUCjT8sPFn6PDxQ
dEy7utlWk44+Z5j+YIeC8naHRJlj7VdH+z8p8T/LChq3IKGIbWpn/CcLWjRvncgU
JKCew8EZuV7oYLQgE44wjwpbIfsg8baQAzzkTJ/Sn7uq2H8fuyW4jBk6RlZa77oz
wM50Diq2ilcYCY+WT+/wcpijqRUSWNzQScDP1NoPN4EicmqlUwNQKC3CiapTWNkF
DVQYHvDZ+6TNeAk+5boWP2SqfSd5Yp4J6G9Icfb+Y90vdtwmbBUe0pePlTtJPeEX
bC41eNBV2www2G+A0KG+g9aihMmhIyordPrDCKGXRPRf8GWl6WuXZrv4ss7IKvIl
k9zxCqgNwU3gOktwd2GNWkmp8jZNK92T2F/2V+s1flh4HLNXwJhdkrXw3pvhs78l
PCTJRKq1g7Hi0m6I8f4k3Bk8ES9rpB7Q4bY6HIMq1OsSSpbyNIjtnOrLF3dR73Zm
+Dm6Tpo6Pxj5iXr/M2uMVsAZQMxL0lDsG6ZBaDYOJUkilN6wp+3Ruvv4O3myDq/T
I/zwIbQNB+5dD3GOvkEqWMpDx0f+EdZjq+7X6VS1NlU5FZoNKLkSVtKVmzqhb0Xn
NzbTdB90/Aey1F8isiNEwxST137B0FGcpQp2Sh7sDhRro7TdlFFzl00yjm9p3lJ2
3WWz4RSbTtRAeE4u6qwB9DRGKnNVBGWCudOOuuUaXbOlfZ81V+Wx96kx7smhNSXc
LOvc2C6f8Q/vC6BVeZIdHxy/Gq8G5O3YtnPbTQYwcydPzvOAQseCI/wQ/dI3tDQE
KIn/OjQuvb3BXsO3s+5PpflvQqAMxG26IxcJyLHeRcOHx6SQR4jyJ3J4jxppAP67
j3329Vb1l9PycM3f5OzYbZW03sD5p9wxXtSI4OQlHLuVHTkqYENZmznRfLzDokjd
DQV1Q6wBCw3FL1jRekcJGgCn6Oe3y8IDKjp/icYoSqBFOswJf0/sSmZvhizKB36a
pfyZcOarokO6RhDR7Wcpo/ZtKLEdoKqmAlblQjTLury9/cTNpoJLk0P2zsojarlE
lkaf7lVap4c+OZYFHd+QMkdqxfhxs+6GmP33arWp7liwtAU7YS2Fc0JODhZ0pTLh
dIHBMgBQ68qqEftPabOmq3ALHGk0SXEw7v8XXyN3zgBVmslD+kt2Mferoxydv2CP
N5wcqCn6AkZCbFPECHoB80bxbAYYYR06Vr1r/o0IOeQKhyl1dKx7IbNbMK4ytuyJ
akYMF3QngeLXjK6vcJcMme/b/ObZURwgOQN3XUjtBX8kUAe3bymMnA6M8XxJz1j7
W8vlBjEqN4xVWoYBB6a3KfQVRNcgB/l3qPIskhRcRe6JWA5xBa/7M224FZfCCfDk
Jmxi1OxPFje/iuIkryBcQ+bYti2IVpe1ImQvI4Wf7zn10sa5Fz0sWQ6pFlBdGGDd
7qrWGWE7UWPMsmvQmuwZZ7++cNBwwXmBWnR3NVGRjK0xyILomVRn9amHSUGnbfM3
Wq0Yu3PE20NjlOBuE2r0EXEPq2dnlvp6L6h97pRnsipCZWAFBg73Pojko3nhkfJx
cY4TG4xj82uMRtzqQv37Q3bX+V3Ppx0AKrfPrs7Cirb+XG1y+x+wGC89IqdLCqko
tXSlgEn5qSKTqKWeBZmmW/h/8CtpcsErpPUtBXfI4/tV7YXtpTuw16FxEHCuU5+F
MBoRk3c8Sl2C1vdfxcB0uuNtx2AE449ujJUiQVH5JjkKDyTGL5xlklVCZcpE15Kk
rsoHfcOtjOK7rKyXG3VzE3YACUWyANkwpQjxrnuGhSHcdlKwk/qQxCu1B/6BYKdR
DTY4Q+WqVKnwNbfjX6PjFR41QC5/gp9ibNuC0396OKzRiFyDkOB5O2ZzHcD8lfgT
xO/80vqgX1sCdYOe56pqUNpdLQpeY4MXsLXxYAo5tltzVcJ2+f/+kDeIdY5vzE/k
iwpnXjf55+JsrGCYy1K0XUeXjO0MVuxkFCIwjuB77QbxRmO6IOlsm+NOigtsAfyq
xm5yP8+GLTvh/5qlY2qbkkZhoM2nCpZup+qC4t0Ri3/F4/rvIb7b+Bgppz+U3PwC
jWWrL5qcKJJ24HK2xvRsxzIQX0iXUkCcmS/eUjDOs4lgcaHMLi6ze1RDVhTjYPsa
yzKNs4+JFjI7BfXk1BTo4477Hsh/KFMLrVyHRlkQu0bCaWWO35Z32yichU6OTgyw
H0tgxCbXkf75e2p+tfDY/D8bcLnhnatCZn0I6bjTPpjDcicTmLOEgCOeoAhbgYfT
Ulj3P9YlZ0pjaP3+cyPuI5fBrXuf9/g4nJAWGOPfO0qU+EAbTsPQXI0KpvUdkpdz
v8u8TAk2kJmI95ck14pU4vqHrMp3/elpY/xF9i+qrhn1it2w6gBeSAATBaFpp/pq
giDSTHU/W+CNcELMvgK3XEw7Qw2PV3NFpHANE0rXMuca3O4L1iXQinhauBeP7YS9
nwMs687vSghXetKtA+FjujaNYVuuc3uQW2hkYdYPem7qEexqD3sir9XbMl+CfO2R
EptVerXex6WsiIGC9ps55J0GwlNWenp7Y2kAllLaYdVxFOv2idh7qO/br3eqGUWS
6ZdAgrwN99hCwUQvuVQ4IbQhZqo6BfuqnPRoGx9fT7GL1cKl9G68fpEyIqRxhk0S
S3rUQ3+lPOQj76jUp/R0F0ZiB0vMtO3WNHF6DM5JCwdH1o7jsXSOvN1RpB9slNr3
z8/3iQLio/f26tw3xIT9FBN2uyeHeJa/soqLzED1ceb+JAevCEO/25M0diyMgLQR
h1yNCOoPvUplY0rhU52VU2B2YEYczKlw94RMVylg5YEIRvYSLXoHXtbrUZadkYFv
WOqYJD53ka5MqBYENB1K72NnypO6kOkLA8bV4aAgxiD3BPLMyc53WKwY5meWAVGC
jXosaJTBkdGzAtuDgDHic+EvPMvqyykgSBL2gXH865+31eAcrAGRRFoXI3D7x76l
xZmu0q/AnebW8A5p6wr8oGmsKOY5lNjfqI0JxAQg87Wnk4Qb1icUla63pMGgVW4n
GoSVHcfzZ0Q6IeWL4HyeUQTncZFzpnvixu28Nec9uJBGjDhNDWF4E12zYivk+/+v
Sbq2LBOHDbQiHaDG4n4s4BuCV3fNqE9ohzZp0g6+eR+mEOgmGvdm+xxq75DbPFnc
gRilJnaLa8n1HvVyAWcScFUb+INxvGFVUPjlI1tQT3Kagnzctu9t8zz7biqFwqsR
6Xis7N9/rYzJWZTcJl3r2a1i6AfiJwYFyrv4mc2iMoJHqpeU2xlAD8fiybLQqB6L
906Q+pxgN+kdBuvyhksQh2L6He/Mb2SLieLEfMGae8554+iLqLlF/+Iv1lXcCzvH
9irzG8c97fQE3gJMRPdxi+2CELeA0ZmE7XsTZgdYBlNVd2CH/ihI1NX9JTXh6MDb
9jC5Ob6GJILr4nGs0YEhQqXC41pzlW6EV3U8Wz3qaWsZeKCyfz83BeZg3DQkIz93
AOZWLBuPd9Pyp1VVJhY9OstJsmampjGJPPfA3JHx65QzREbJmdaXq0nNNrHA31QN
sqOU0g9+NOX8fSWrM7g8VY1x8m3xMgW1vNU71GvR2vkMaWvYQVnlKy7lOeOZ7tfC
KJni/dCVe6kFjD7ijT6RXEule6S9Zr0NQLujNqG8/nm8slXUTL74FBrm1G2WlPl2
KnOWtt6WbhVckRBS36GsFgPQ9AVvOHSDefDp2sZlCYJVoIUmAwZH3c21NDTu0KX4
PPdfQk5Bc0CMxdJQuBES9bdJKUygAcpm+kfosgM+T0QcCzz6FaGCPLqLq/unGyBd
xsyiSmIRZqizNeu7uonNU/2F/HfIRv5dUgnNhTAAggXvKJgIms+W6FlrzjKFswVZ
WrQhsJRAOM4C6BnPfubhkc+FReV6mWcCk/3YZi0mlEr5HnN0/7jqG/Xt4mkGAZ8c
MMVAQimqNR3SvhL4nhrDt4epQbZChiIC1w3ctSUpRXVoGr51gC0gfaIfcy88Gi00
2D6DZjpals1hw0jBxNXSATRMBPhhhkgjyK8UnvsBvlTNTKbjUlbqEAK6nyO78luM
fjFkxA1GhQ6nM/7qEYQC3LcdIMqng0XKbzxCHrn0DXfMQMF45wM1Ge9OpNfmyYV8
iJP2DVHYpOEEqvl7JvW/obs2hs4PYiP5FhcPjyyUb8mzy2qoMa7vJAyug6JDUZWn
2QIBjDNa8Z67kiTZptk4yzskavWNGjkkc8IwC4lFTnCnctYWpHH7gplK1L19MtlN
dQ1pkI6YKBv883eQswzge5l/S7QOjtGpnAwBAj9O/ylaYiU9LN0RklCKUcwHvTBo
Db8HhB2jcED2L8deVk6n7VcgnNqCf+APHgrEHgeKF6K508uefIou5ESE36mURKjf
jv068L1/UodSyiiB7uzX19VgrmbijaUNrS1or70+xKBvxi11cxEZuVBPC90Ic2ni
RDfyeL3PPdalTa4UAwUxUiSUh1MSH1BRfEfIq4Do1mvjNZxzZKU7EMcvCgn25J6l
r+r6oA/6qO06lyVxGTGflWpIBwhBsm53+c+CcB1qsvAf3jplqoLdmujpkXjRNWAE
eKVqrT2/p9MNDBvVtuETnoe0HHBDZuxufNmKZGklywXWVLQjakKheiFN/+opWDQf
9P5l9JFDgKP0s3/txA3FBDo0BvOobyo6NaRuTG1hvRnvf2aqM07ZPi3p6l3g3TqI
ynFGeowfGrP3wxojdAwOcmp9yM7e1CN5wdTgxLN6qsyXI5YiCYRDW5Wx9gJifwfj
rRSdzcanHNMEvhuMI/7RegFAdC+a15PoUyzh11pXFC48lJwRk0IEfmyNvkytQlCb
NJRhXH0UQNb60jXxWIqfc8Q0A4d/UQikFigPhTEJv3wthEg5yhLGsJ3S9vgk1NGX
FSMOkprvLo+PMn1eGpLzuEGEM0BUTCvt63Vziy6xnXLyYHxIlxRTMgzkWyyXcpiO
+byB2tYhAgd4wP5aLTB7MO0sNukBexRbnQBR4Rfqe1wp3D2UvLEfYY/d+nW/cm0L
hKoIRe8DzCFeaYCteZ+PZZFVxtZk2sF+GJpukv7RaJzPFfvejVAaJdmbXm6xBacl
7FJN+QV8qKjTsY1uzrB8MeXRs8QU5xZLAsQ+1QyXWblOBRwE7SILBxtjFCQgnzR/
W7+SbycgYaK9TYw0imaqKJqSyZouJ7FQa8oEfOvcaW3JIJ8EVKkSrmpIx4ekK03p
YKDAd+JbO9gm2j4yGuN92oYypErtQwM0D9rY8uVkSMbeda3Wfdu3KmlhjyUmlOUs
vGpY2pKV34kzBffqZueZuzDIz4+vm3X4SvOnOTFpfMYqsIEEF21Q5ATgwzc8V9r7
tuDHA3Qn0fii2ELbJloZJ3watB4KMmGXehy6D6VkZDX4UrkTeuKlQwD+T8vTjanp
0cWRutHQ01KdvePhevNVUbnhFoZq02xmM8oJbXYYwp+Kqg0U8VTsWQcR6OMSuUNI
JSVxA1OXOzaHItoFPo++iTtzNcc4039fmKV9OUc42xfGPMwdyyY7eBsA2CxwoisK
KHu4UxZkBPbSgNb3b/N3Ysg9RvY5RnCHILwBJSxJ6YqmkXI/89O1IL9dB5z+xxUr
MTGn3BUCatEOVoZz+HaWELxORnbK9wnH65mWlSjE3CXlVnXa2gt1YB+EPPWBk8ha
/QByMGVV8IFE3YSyvi6O1eECvvhH0Zg6gqDNu/GhcClyjgH1Q2ok6ntbJc1Z5675
UBSrKeRg5+DPAh133+Kl6raSwiZsfl/xKRRd0oA8FwtPYEdY1Y4wjDVOgxM5evk1
kthBgAIGXQMDSPXRNeQ8DJI3biHnWkbZj1HUNg9hU14g53lGS6fxADIDtJFozLMZ
Z9JzbeQXXqqBcJT2jB8EiXYnfARGxLyIUKq0GlZvGaTHbbyC42HVTt3r8FuVws88
1b2f56nPGoDd5KhmIqkb186KGfLwGYeutg3/tVfAI9EsGKx2yCAZMLcHFOZJqOkt
ztCS6fgQS3QzFjuqCCyYXPQbDo9MbyQTV0h8+3gllW9qvqjZ+ohMzfR2aCCRn6/T
osvgRAiiSq9YdwEIIaYVLCIZ9qvt2aEiKd1SPnpjb3f2cu3lLQ0JJDUTPj9kys1d
XR9K06PLrrBjxj+KJEiFIuIw6+y1dgwQw1Dr2pbGFGcOI8QOGOheV9sj45GDDF4C
+jbxxsTDCAXTkUIcWafdpmNz61Pr1jI4TIgkFGjUOx30OTVj6Q7KhKOZSqKgW7dW
jve7w/8NUVaXi0RQirU9gcHI7Pkg9mXoXFxMaKm2o9819ct+sBUaZvo5E4Vsuqzu
uTGfa+UtCTuSbAejwL/2H/adM6s4UvNpd7jzSttWTBM990uYC1szXytECxC711qb
RfpBoZp3x2ZPdGFZjNyaerE5/EphclK33Rbi16yVJE/wd7h5l73yXr15hzqmDu9W
+Ox6glZJt46qVZLzaK9aLJBTMRSNUjQj2+iBhwhhDYo0MXl6tsoQ0cxTjrjojEbl
C83iAv6+rBQ4JKI2vMZW/vIhAwtWTDTgp0BkpyjJqAFIKBg+kFTkLX0IRYis8yZG
SHeb86d0RzxjwepbHBIBVKoGJMnTEPzgWrA2Uyx68j7v9LXkIKXJzYYxHFjGiXg4
W2CYZ8eXiNXyQrYbK2wsw94wCGafp6KoAcAtFD0gO06LfyXR26LqnjXYUw8/tCB9
op8wJFTbYTkx3oMkZMxLLsPJgqZ+arpxboE/iQNx7IBuYW6lj1DaRzC/6nj4CLQz
JZaklVB4X+KlhDbyz6VIViEk+VN/bYH9soGdbndUdqFDjJKoRZh1nQb5t+rKfvhX
XhPgqIswwjB/XOvIynTpqP0SxpGJOE/78UhlZA21yWUL9LNkGW8R1rpAooasoggn
MIlVi0w5ZWWIr1ED2bs35UklYcP0O3oEBd2SWFPuuTJMiVj3jp+GP6h5fMIi+Zku
QIYdkPgQpp5EnEfLkGe0B2wsnvNLe3tWzd+L3lTOV2lHGBLVlVDbOS+/ein3TJll
CDP5MWKdjkSzkDcNcmSUmU65hNHwFhs/J1aW1DV4kpYITY0k6gBs/1moEUE4jvF5
te6zMY+UbFabl7RW5aNl++el73FPC8LEZ3JJHOFijYqZFIq40pG631wV1gTuM6Mm
wI20tHF9xedZiJfmDd0OmKD0yRGp+sYCajmWEFshxKWtyEyLI6QVEkS058BY01XU
4fisEcPtMuOqqqTE3r55iOMdJ85OS3o7fttNcv4RfVivdhUtkWG4QB7Gpo8/TZM2
//SRF7Rplvvt6Jn7u6q3SqcE/pHbJmUpcExMagYvevZxQnMx+kkMJbmNpVSdvhL4
ZKrZeVaR/WUFDmzmX8mmE15NbOsx4LfAGaXVtIlJkJePciE1Vdeq1GmHFUUSCigs
PwLpcICXf8xmgRq/Yuufcc/ueTHOw3LU8hq00gkBRp8KBTRS5hKMeHyUWEizq69z
iLM6UyM0n6jZcUy3sBrITeIVHz2f8sA1GH/oHJY9xRBcy9RC27w6t2WiHeyKcSot
hklS+YWCQdH5bGWeFH1XfpJFZkV9+8y1SPtpUXPu5RM4DAtarN0dgTkmenuJvvyg
FGUPBYunv9VteBjfAaMpixf4ezsHHg1+lAABctO3bAHGtPkGMunWQPjtGeVa4kga
SZWcEY10PeKqc8s39X/+niu+sWdj8xweV7sG3wCCM0B3DIKI5Oy9tInN+1E0nl1C
+Em2xU/PadQPjyQk9tb3rjdPir+jZZ/fqa7HmBAeJBG7kwAj0tK+IvDvZoV580OE
ibdUTgt8Zzp+rpLzMj3CWqMK24MbE+yxX7ojFHObWz7hkjzoZY4H983IoVQoC7Oz
hGo1njQVnKlY1iH/yaRV2OSbyt6gfUHkD4aknKuhInf8ORNDoQRcuKBwNjs79MOM
6x7W2rEc8Tv6Rh4xPYEo6uEpxkPOeTIeujxiJYCbk0GthdXa5G4SL0KFTouGCL8O
VKCsmAm4mBlriuD5/gZw6EGloX2HTu6LA2vmwhI/lCvIAiERSkyFxKCOrdgNpLsH
m1hxnVA+gAGErtKl/EdZDgsRFxNR7objdODFZ9OZuPnSecgU5n5ze2RWB+IHfaJ0
WzCpjJX0mDyKO3JeOzKxsFJwPVOyQ+/yrV0tU/0jFS/9skXjaIJ1c+azcOHXJGkT
oRmJEvr80SU+T+wiYRSzezDnbGY08501WE2djTiKCZXvfcim/zHsOH5vlSDmCAGd
2ukoSXSyhPEmpVoD2SNzY2zkpGCiL4CNLImY5fBtwANNm4UNNWtTLoyFqa4JjIFN
eJq2lhE4Vo/ws7vPj8UzxpUynWAH7VYHLvX5kQDQOccP9ijID3emX50lb6Sbp8We
B1+1onSZc7j1w7zhpPbKHxWDC+xzMHj+2t8WKfD1B6Er1o1GWhwjzlyA0lessh/b
HRia21GvafUSQA58jFJcXo1chcv3yL5NlAoL46oAatDLgYDe5x+yrDgs3yg7zOTX
yXivzISdr2l5enoGL8+CHEKwvcnuGUwcJP2in+lGxZwbqvM7OEzdlg5bi0plNjLq
pFeK/2C/xmvAdZrjcIiria0U/d1toJy2RN+r+nudnC3nCDDNiqo9f4OpOmZ4tJxM
S5R250jzTbNuf7H2KVe02XVVIqh7UbnGOe6ah6NFWmiTHVpn/EPC0gsLc0eZvhnh
KOU4S9cZGv7MKcJaiYI63dKlcuc3TPHBKF6LnhXxKj9Pq/W6jqI0tw4yU0r/4/fO
3Es9Ea+OCn04zcFi2u1Ud42V+nFwmRKaDleXLEgjzVz0Qj7Jj6Oon7mm9MizJOyE
sHgw+J5AYnzA9+AyT4qLBRPM/FC7zsWD0Rf7wdNX/txATXDZxeuzn5s9RBdKitEF
C5Y6gahQ8IjaWlQpXBtmJ1dm40TzzirpxAKjKuFwXRBeT5zlXVgGWlIikwW2Zuvx
e5mMmqK4dp1QxD1KG1RysouMcIe3eiZZWHvynWpidxAUe12DEZo/wf/CwadghdVj
AcrK8JnlvM8Cwx+vY9/FSVrOkQ1G35okOaoV+uN54UPn93kDZtBAmFXiaOzj8AwH
ctGLOYinr6MkNRYKjuBqtw9SAoEc+A+OUlt2u4/2iUk0RnTTY0abHYsiCjQJPmq9
yGcXasIwWXh2d3Hzw6ZeLR8BMgGm0UFECyfGs4/fQOsFY2+iaP2Q2HGpdmuSTeF3
REVub6pcTbc9BDq7HbvF4NIbkgzeHp6GlEQeTwy3/UeEDV+ygr3u/85Akd0jVi2e
c8krR/41kt6bqJ3a3d9hf39uG9vx5qlNUBNt/lWXI+93bhOvMV88087NkO6WxU//
J2PdE4j8ZWLbYFEpcEWjBMbvbWoG7AGkP4XPilknbI4ESZZ7S4jPbxOrOuHwd1Bl
gEMAlpuhUucIw1L7Jv+Qn7WJywUEycpm9TRdvL+y3IqQpNHOWJbLIptTVrqBcZyj
fWIGAN7oM0bnoSXpYa0t9ecAiy7NtFaOKPT7fJHCayy5fC5N+AYbNRmrV2k9oNQo
8o1SUDjOCimtxxuHIhQil3cJ78A/03ZWp4oFND0QDomXw2x9v/8WBrM8VbK8i/Jz
TrCFQgI2qp1DhkkochxOZM3gtKhJY2uKHKKJiV+sPvfQa9Ps03/Ey0+YrWCo44hI
4L2QlDNHNvNvRKUdBv8Uxtx+FQX1/jzkOluA0XGPkspgmURz624jKUyn7NGtmpCE
/bXgCSB+p5Nx6zKJjdwhRfk/YO6iG8schD0xtvC3b6ztO1qaVc2AQQGpsR8ffyeV
6a1wtZ7CCALe3nO8XsCC6ZslzK8A7fbPO6FG5rfGrxeTKaf9u2dHUlqEsxVr9MYh
nsE/x7589Z5K6e/PHyoJ291Bg3lDNj29stoBLLh+1oIcROuZ0sCms8K/IDcjtWdI
J36PBkbG0n1IA+Q6jM6NkAzWII4F/lUlEpJReDwyJzr++uhYc+tuIoTzEGKk3qT4
NODw7vkoW5zJz1e1w5vN88e8oozk/gphHvaE3WkrNbqDbWwri4fjvkIoKbavj/3d
3aN3H5eey4AENsN5coNlSldK1e0frgHpfprFdeWdgVSmOOmnQ3pdi+3R0lE+X9Dq
hCrIKfa/IGZUP7dUMhVj3HkN0BcBlM0zQCs30ffSi5T5gdtJpc4kSafoBI2+B29q
GS05zsoLBqiVkEuH//AcRTc7CoFqNOsz6k8gaE3gj6lbyZf9qmezy1qGbOYUgxdR
6laVXUDSP3Bq/TxLf/4fu1xeaTdWc8jficJRg5IJYMhp+KeGare2Hc+PYSGnltb5
J4QJaLEgHP+xRpJDyM0VfMTmMqieB44Wb8C1TbkXeWimMB2xB+eVpNUFhsx/BWNk
+o+BkXWiwSE6tkZhf0Zi25RaKxHwrU2Uxnf5cZjSUnkz7O7Ijja0gI/q/kZto5o0
rFzZ3qhXIEqTgROPnHjmeoPOyOQCXuSUUb4MhvtwU/kHB4bKGg9heGignLmrsC4p
5XDwv567xeTmW/wsky0UEAnKHK6s5GfOg975nPYqAYSTZrV4FcKDTUg2yZMfbsfB
IMmbctZIDm2jLcdgQhjkABqxrjrqwSEPBoqM6LL2vQHbgZmLxPhkyILq4aLDeHTL
2IuyIkFWiisEGl621nSF1umwVsdNO8fyL1qdgHzMG6IRFUPMz++c7oFfg2s58oIj
/EqDjW+933NRCGlssmyWwo4STlRuiDDb8BeENxHz5SKY8P93WqRoRLP8C5ZM++lA
1bQ1QLRbZILqg4lcCu4+Dn1QXpxoXeFOTvIA+mfLEsR8NZUpgxGboKa8DkndsaDp
mbvZlkXVZrrETo4V7i6u+wlMtdrkPQfeE/pVZfrc7QiS2GjZ4h5mMv4gzgmRmgEY
FwRFvZ1B1aNQP5kKcsywNLrIo+6b3jnTDYmL74dpcuJDMLj4f3GUh5pcXJfL8Xr/
SrLWiFR5qaJzgTc96sICt0FB/QCIQujxtNjZ6PFFotYqABJhKx+VwexTd88baztP
rQ4lc/H1i9Lo2uHLui8/3+/rJSNPXbhYvj2t/khpaWVVXxOaNNvOruyYVwPZSRaG
WgffKaev7OguTB3vM4ETvpku/FDii2g4pXWvLXOSIGWYv71z4FjzU0XOoemcYgAg
8QR9FfQXY8o+ehifPAE36PaQaAeznHPtShfoSIbKxtprHYLTYv+4eNdlvaDZpQa9
ZjkxbDq7/DMd7Nq670R0ttq06uzg/+ZzrHLRAh+OniVuvqKFARgg7KWZ7//znpLC
zYRuR4WJy52ln5Gt1+u2aBeqV9ciqAlILgttdTcEZafuG8nXlpb2/pBLLuiGN+12
luHSDEGuPqioCcNqjtCGA0kJzGS5J9V+0sLGPUAmXfro69gduvf5zH9r+rMZPxuB
TuPZdM7QWb+x9/nqH2Nb+E1Q0xcsZDn8Y6PbDePckjEEHrIKy0EGLwRdmIFaWrHZ
X5RzLKnpBilKEt5lEFJ+NaWLFHe+qvqowFkZnef22pguk320/LoXvz7LbM7dpLi9
RMXBePCM0bfBDQBQWITxuqqZYjbJq7DgxeTN2DSG6mTM8zS3QmRXPU1OufBPtbv/
h6q+NpsrQzPcf5bXBVFWCiFg1ej0vuSTIZELkyLM66fKsunT8X8cx6s0t+cIG+KH
JoZArTaVfwV6h8q3YC9Y6OGrLkIH//xLh/CJa3P++fzn7Z3xBnXoFzF9j5uw/qOv
bLGznD1EjIMl9h4oZ1w4V4IuYDF7xVagPFP8oZuVtRzLyLs/3rvyqj4etpXWHNQM
MSwzy2/pSZCpsa7lYsvYnJv9DsIzMdfrZwAXMHPgrcbSbiNMarCeyl+35xzlx34r
hE16bSu3/STgsku911IOHCEIZya2ghDi6fSm+22Yj9ZmfRjEHY0fXpcqKzjOxVI1
nnP/kmzmca1uoTsZ0CA9TFTykxfh2YMIUGfwNgN2DrYNU/e5o4PsIkUYixgVCY6X
wzMvnWVJSkhEGId5raLPxUIGaBuhao5VeEFEfDoNM6om02O1KNSvhkDTl03XGD8H
hpswQQ3Nc7P3n0UGNB4822OdL8Jm68A+Ao70IMOk3UsakqOg7PuGF8Bv81UqmU1l
aB1/NccXz7PujvfiVE2kIksIek02HXr+0MT0IO6YgTBIZ9C4S1zG2KjDY+tiXfhs
BXp0KwYdxFqsCjgIg9oMEDqjT8OHasetSn7S/Sd4Ao8qHEI5SlXmE+uxqGhIUFxM
VfTtXSVnBcSf7IjarBm7gh/y+ebJGbf/8+aFnZZRAqXFqw7ABnHoXqY8xHX7CrF2
TSiQ/iNJNWdu/f8sOSWEGHJQHcucUN7j+nbPb/YLqd456ZUQY+5U4gHiEF1lc8EU
v+Q8TOGuNA7lVOMs4XJPf5CQ/LEF/RTuSjTmmMK5i04w8qXqOyVwcObmfmda46jP
wqlh5VcJHQ13/+PZ4cPrZoXc3otYUw0Dkgb+/B8XWovlZjNgBf1nxPv2vQYuQvUl
V8fJIdpIyldvev1tFS3tjjUDWbYYuVG1y2RAga1GxNQI8THdSz+Fn5kwuXwBV5zY
sJFQB/3GqcXPJhvRpd4Cl9yN8/5i12uSdNb/o/JQVqXquRAYKY3h6QLR0Pru6VzI
Y/hqDZWTER+SRcZkObfLRzlD+DyusT9Zv01h1UI9tE1zuqMoeXerfF8VvJtiCIQU
3Uojxwblj46/y1Za26rXy21yMq1CkSMudWHTXJ9I1ItZIT36VeUodnNd82cSc4Zi
z20fN2Pqajr024XqxQzB0f8IdnPFeT2TAl8N2nrlM4FC94nSc6QaT/RtZayMfs9n
n47NE3yxRX9zSVOBasETgUkP0Zu5XEArZGHUbigbVO+kZT7rbNhkjnAWpIlhrJzR
QixRsYy5ukSr+6DKdU4791M5qhc+pob8B/xBYdYDzsq3P9PBfMmcvZGb8rkTYhax
iMGasb7cN3WhpZrZZV2hlR+QQOzcYm51dd/Gl6xzjSnqzrsHsnGEDGwzMVAuyEcy
SahR/4v02YPf5UNY988xqVee1vBEG43YIuiotHlLXHfwf665KLgx6hqq5w1ENGcI
PDDL53ndJ7kub7MdF5j2n1f0aWlPIKObifu9uw310AcQIVZRRnZjRx6U6UNRwtq9
98qbc7hCjLkO/KEZDaxrSnw4hobGTzHGu/HAll6xAHWppdgMepkTL2xgtDUkvvrv
MXVR92ED3JwLCJVWwJ2r7ERT4ilhDNHsfk5mgqCKKEFP+9duixhXq1QeWb5PL2SS
9Qz2/KfrT2VxvSXgiP+qo8AbkgoLs/jCloPJPOSE5koZVUtsqS34wxIiBTZq11hb
jbWC22VxSWZ9nGZATkUggnlRqUGvOYo7gMsrzx4KQwb5aq7mB9ZOs1hVAkU2Uov4
7hML6jnNG9N7hMxL9Y374qMX0J3MfsHRnPvDFOJ2zeHXMF0KKpGL0A64fqnSZvP0
GoPgwUC4hgtVZpnUptv85lsfcmNYsaBeSOz5sjGucx+bOgByv2nUMGF+bbfPHG3A
dbANuakir2CRuzvhR0CD8J5P8AUtzV0eIcgOHj4IepK3hWHfhvQCm35uEMdG7zQG
q4LikYybr6DZ8K827o8hOBtq9p9Chu7f5xLNSQ9oEZIyhKVWomp/aMl/ZqDXtYOy
6DiZ480/f7UiX3hVzPo+xl1Qwz7EK88/E21KczB622YUfrqtqZjtW7R0oy07fMPk
f/lq+gmootK2SQmWKrNuhp7LcMGRRslN1rVpQgxDKRfVsClEmJpbLVE0afZeeemD
DVQkLzO7rFeUUTmllwo8XIHevPWTq1cB4+n23HPQkCDenvJC78fG3B6NrsS6i78a
SOqkJe1BcBzMBs/WRq1jfI9yrgCR32NtSRT8ZezwqIU67G0ulTfPkytr16x7k8v0
FFeHeE2VkVZJPIHhNrxog8xxODdQMuVPfvBda8Br5EtZ5bMh1Di1+aUdmnpcgNCA
tiUQDIotfyD7Y1uVwnq7z+S0h2ErPUCHZck9uKOF93dblGgcL6yRgzqGoYOqfuCz
YduTyYSM33oyeffoK8huN0r7XrnArUW8+yKPAlDQWWr77rHbZKwEUdQaCFZ0mjJC
56D29Nr0Q5MyaGXl1eFm0UctHOPRVPsOQl9TMwwli8OCHum0uRMoO9JEhazrcJSC
E6uS+19Pecx7iQMc/insL7I4qXQgKS3+8pj1f/dudJ5S+VlAR0JImMxwWO/Iw6ar
V0kwa8+E10Uju34Boaa3WhCL5pXvm11gwjlx896Vxv60c7IUMv5fYyQxEo4OSchy
I0vUrSDMnOAClD8NhKd1tfCoSwPP5Uz57Qyd9B+IRdObyghwXIuICjYpyJ5Oqjs+
rDuwskdUgKgdWt/PRm7SOuhvsbPFPAPYWLWfDGMJ9tkpoAfoWzU9/6e9DpEwqgam
HUaTuzZQzadqRi1QADtx6cuDh7FWaymUvuPcK/mXJuIhNnPJwk9mT+RzVhCjtZL9
5+PMlr0cOd0/N07/0czcTUxhZdo7BIz1zLCHc616w8clsxhAa9PeDAbyt/6OFG7p
Pb/Ct8kF1LAaGmyY3R64fofeSj1UBSREpcKaQWnuJSqawWFu98r1NXmU9WrmBNmT
U/9F0wm8UvfEb0p38rfUc6KfT+JWsuQeMWhIOBSQaCW1PDB8wjUnaqTACMBJ2udA
JaxI844ChZqqnroU4jVQ3la2/U9Qt53N4nKWf8RIVQhdmqEoXmd2nD4sOUV4lEQO
AGyCwbflRExa7G8AyPS7mFjwEupKfFRRuMtuk6u+j41LKqqeTqVLEGZzCjWIEyUO
OiFvd0TsoQChLzSJtKYrsNkiQKhKpD5LEaiSgcPkAMPwtC4bfbaAvHzRGeTvmiNx
UOGaIb9mlOHzuqQvQu5b7PVCEha9WBZi/Skw0Dnf2aZ7b3VXrGbBZ55FJo79DU1L
mSVAvh/yF0GHT/B1fckoT1pBVGuR6MGCEl9WCBShcwf89qYvnUQpWdd4hIGZZ7G/
v3JzmM698yqw380o04Zfeap16Z01O9rn8fw7zEQMXMxsBsj0smhBX7Vs6H9IMLT7
hRtocuWb5ShIkfhfyF1ntx+VdMyLUYKgjHHDcaRdwgo2Rku0xeTSpI8uVY9zQJ3Q
NBn99f7k8zBXtcXA4+Xo6r8U2GvwafB0ku8JYlbrDspeNvWBwO2ykKM2YHRyfhNQ
o1LClXL+2Co177B9QzPrypWsfG7dFIRGhVi//pKupBjjFjM1Ac1mM6VgnNR6v4vw
HHFmvMP5Ux0c1Gl6FZn+DStgFd0Jp67zR1UOt/MTur5Tpt2YYVEH0FdROqmMe+6q
UGCngCyNIfxoOw6Q7SJ1xhQNQUKr44GS+qcarNQPxn+JfIZ4r2wkZPxauvZCsnEP
ADt3zNkhaauYe/L1ZZj5PXyLp+Lzl8SMWnhIg2MQMFapxncm/170nxtDQtK8yJpE
wJhvVQBj4R8hilx6MGwx3OeRJID5hdKL8SSom/Qcl960TaeTBqbp/6gU5JzGkoig
PqMC7tMch7oLco3Le6nKZ82Xxp03UUH+GWVmZUpoQnLGw/mH2Y2Bsk/IwGU0/As8
SlowVroFoEKJuMvl1/7CwpgRSd3qlfL1XjTVK/Wp5gQ5a0Xct5qGkWAGdTI22n7E
elfojarU36ZCdHEI89B9upPSNf007t85UWIoa/WJYn9uFmLIEfvfFCQg/BsoxsUw
3jYWNNfY/9oh7Qk9ELnHhLh2a4THoqY0ddhXqleGAGqM5ia4ipIChle14zhc6ja8
wwYdEo23JvANaPZLLQa3fPel67py6thti7QJDN86ii/fP7y0OYgZZ1m1QQgQnLcG
YrnuBYXXo6BJ80jWOgGyUimwhoCnRdvFLRe7pW/FmzRFSJTvhipTb8Jdpo7qtsap
4i23tX+okHN3ARQD+ZAfs7P1AnuARmJyGscaXj4JRSinwUZ7sMUOd1xD0ve11UL5
or1hcxuGl/lE6f0T/Zmx5kDj4EuA74nXmxam46EPIpO/Yxnyw3ppnzFN/ukoIvZO
e1zVR/oGd1tXisJsZYLq0B6ccrkimbv98/bETJMWISpGSJAq6tyvcxP2fj4BerFl
9u+WNrS4OEggt0VNhd7H2E/gFu+JZCMgxKw4nQHASL6tws/NVg1m1PSkrYBvQD25
JdtBNkk6nfgUkp7LTmZ5xwNEwv0YeriubUOgb/q3394JXSZU81neV35/x2yJy1Un
X0JAuVaoHhWaxXalzr0QTtPfzpY/Mrn//qOuLv9xpIs762AWq7QnMG/gS1wFuKtC
cdXFkzQRTRhombtw9fIBBd6u7wvO4sY1ME/Wh1EETgoSnIGwh9TAuQR921Z3YcQ5
5lEbOIdQSdPjzmkC+KP/4sbRh4VR7zoDLcBhsJSu+dayVGoSmIThtA+X+az74Qlh
aQV0zsRgMbJIf44X/LnpC7TMkcoEp1plBauGCd5qSUPoWPjOx87vbVJffLNmyInt
dvmFUqQmwBuxuc70j4oC8eXHc5KFMfj0UyG0k09BdcV/WKRf6Cg393g29elg5XgH
WXPFScg/1NNIwVkon2Pd5Sdk4OoFxMDgdhnuqc9ojAIrhFE/on8/8/18P15EdNdE
8ud4T1p/c1vyjBv23J3iRXMsEUw934e9vGlCoJFxmoCMA+htQ6Lb9Jcm1Xge4hEs
V6yjki6uuN1rAsI6InB9vt5/eWUJIv5a0YxJIbgtiYe1mpzqb+l02jG3n9AEKwQq
JeY8nKXfyMPmDmam/iRau7E/bzSNO6xwcTGo1P4Z0fm9tBmeK8Udogv9RJTAP5ee
pmqrwC97FP6BLkoWoFn4qc7VENPMzgNkrm4VxIjkgNuaC++6aOxKbslFvaUWsFhm
EeUmlguLcq3xaAARqdZ9XC77C6KRnZrSluNS2oSdc4sw3PO20LDGWTb2yZrvUWzz
PK6fF1PjSefpFcN+6MoW3Eh5JquIaQk8vYTvo56QL0l7V2RaBAhoM9TRH9zqut7X
E5keVhCpFy9nzAGGvXlVeqEpPrDajpA6PCmSQyoMzpQibIqRr7OySnliTvbwRCbD
TBCIJQsYCc7IZup/8ZtXMcf7OeIxBLYa58x/4DTxIpao9oScvH537pQ4UlZu7RwO
eFcqw85FxNKOOxi9J89mkTAJQwKMpVTeKM2cR/g6RhS2pTnGM64gBb9a96GmiF6Y
egYRDvtahmixt5ppxAP1mk9ZjgLWSYKJQJU0NDbSRoC0EZ4MGHsClSkf8Q1i5jd1
Mh+NazsEvjqJJVwO/DPrKq5VAUqR6PT8ORe0Z5BHtRatkCZFIRXKuoXr/JpRWZoC
1VApt22aJRmTUNhuP45zTrDhJxb1jwsZWV2RPYEvkMkm7doZOU8Gq9TOlj2WA4jI
sQb1EVSnWafsZBjQWhRrCPJgNxsy3lv3AraWoqi6THIzykJ2JAE11aSmhzvxLi8v
WlpIzus0DedsGXiLnB2G9TgGsh7yPssCltboGrTGI/T7hcFZxZpDhcmCN8ZWUdPy
Wt/g5ZTc1D+V9nrX0Oo1vOgMzeLmF82uT+UclJJKBokYXbjWgIobO0K1pY1uqYUI
0z+sYjaCWeRHfne3igWYVbPkOd8sPmdm4pKbSUBAG9O0szoPlSoeIeD9nY9snIlr
ZOz/jwHR2frv2JTArwohCbOv+SZZaARPK2kR+sw+auSrsdE72CnMsMrnJ0uLvuow
4QCt2FKgkK1orWAbts1MD7sQQG+u9U5qpbxGk5uSAL651BtmCuNjJpMxrU7OmSCA
3MuV5V/QdA922icoOrCQw7vW+b1YMBHMf5xts7PO7ri6OK7p1EdSQM0JPqP7rdwI
04/9/gddYbVsLf1Xv2TudBVkSfqKs5YxySi4Hf5/sCIj8v08Z1ypRi8oCsfj7WSZ
lcQ85fRd1o0jbv6bQVHCsUL+Dy7Znib/oDNj4LR0MwwMONWz+oQmR/OzwIpNG/Al
iP7O010IEPMT1+pvFA+KY58tzzZyk04J2i1J0pyL+lnJaGjyrcKT6c3Qo9cpoy8L
mEyJLXnw7o4BO4a/atskK8hNWa13t7xO4Xmg0kEpLiEe2PdC5C5afYxD1ZAsvRIk
E76UGmgJZ4avj9gA8UBOcpSeA+H2sKDp7s5o+2P+/FrVTnSNokbTD0p75iBZftjZ
5czkHL9dmDJuU9U1aGGfK86RCd2GP70QzO/8grTXSo8lTWA19wNMlwMvP0V7BWSP
1sJ6iW5vN3QQjxTbtO1SvbDmBqf5ue0CywLNRrR0YCvunbIEW64z0Tyr5MgLd0OT
pA6DeFbBSKqGzf5cIlI/E/PIfxB58on6GkEAe7DtE3c5tPi042SmZc1Qo/NCZLMW
SEMG57rF/xxk6PAqcZVOj9zgVebnoQxEKwGaxG4b9cInLljTdReUlLEWzWtfdPW+
z2TlH5dUgANRAfhsH3gzC8LfIECHfyGzTzit30kJQNJxq+Jctx43YouJsGrMyp8H
slyOkHWTBEUs8/J8wIKMU+uxqto2rrW5Nf2zmDSXv7wpQ6FFfagifQx0sc0av2n4
aesy/YMdTzw/5Hp4aWrLnCjZeY27bxFmcxPliw1cenaPjXJ8W8Gg0M8Q3h28F3FU
3nsO7KYmVIVW+M2NeQGwfxC6Au7fVgR8+TwB3qoQieG6XAXWvyhSQQxLxbfdylHW
4FGg6aYHOSkbGvQ7hW3ttrd8c3hoZHAjQ2nmfguBa+NvPeAQPv+ic6KQYyY11kyD
Yg68TmbSYFLNsWn9DlFJobJrZhcjYY4OD/5NBaaq8w6GsX0yfhfQlyyvGrjE29O0
EzR3lhbz/YxzfElbxpj1RXDGyxW1TQz1pAjNlKr2fJCc2avoOeqSiTM0PVRUG3jC
SikP2jy+03vvYjfG6ZWKkvcazM3tIgMhoYiA9/l7vHRn1A8SkwQ9J2g3AyALGOPr
zVtPZViGDzKWDJOaC7A5QyslZMPFCAxWj36ULaMuIm09aQ65xn9PdkgzmqzBLvFG
6dK7etlVo5E0ArcL+HQSIyigJYaUsHdt83GJTcsxVdUn8Y6Vj6nJCgt/G2lkRahy
v1EElGwI310APPk7kQiWz84E5/VrORbpmIvAG0dKk4bkNHuD1YMLbfMxMsuF++/u
2SgB4BWg1y63955XVgf4+SxXg3RmZLOmCk5R6cYZZJdXLOY4I6XwfG3Dm6PD3Cq2
i+9PTsSCYFPOlNx7GvJKpDENUnMe3DimrOt/0eutq4N59pMh3lHpxa5oB54G1VqK
qHtfpruuq7X+hvdHLity/myc1uv3Cf2VVRC/J4+2fH6+z7Uf1stv92zFMccOXJXZ
oBOgyAd1ubISMO7JqAMCQ5vHxeNc+qSFEItZj7vHO38bOB3XshZ6RJMF+3/ufwue
x6MaVSf+UMGx+H3SRN6gObxqMIkwK7vW9OweyvSLX9lorP53wMr8ZLhjVHbzKCJk
ohdN/Uq7sBzwb1DcPVdbBchDWItMsRA1/aiuQ95IZlhPlVgM9hUgk8tAWY3AogkC
nfxlFKQRuyQ6bEQZ5OXLQJ8d37LyA/qIzmB18VzQacQYQFJ8VzcKrNNVP+LdifaJ
rIFiOHQOuPgOqt4GWs8C2wAIAatdUWkvvYuI3I9e5NBSKD84TQA1FuRHx8B23ZOa
iQzGq4hr44nH2SzeDl2CtBCeth+JBGoOJYAkFt3wYo+1jYI1G9fTVbXjivbdoJgW
2e6kX4H/c6BHmd6BbbKIIsKbQh+4Z1wtniZw27+F15NKo42GzCNTSdaXb7m88TpK
irHKuVLkrh4UDQSznMPnnJ1NMhC+gDCEZulS27jNpjH3hEdFsFwvIu1luSgiJfLE
fHolq+WaLpaYvwDKOxJM+hur17OY7Q54dqDxCsZRR8x8Tx6yTu5PqUxF8gzheHpY
HsN5OVDp0KU+jEuftpLR+Ulmm+MVz0liJFXUHDwSxaAAoClF+OGjXyl0IR7bOZ7U
CkPaDtR8U1oAIRmr1S+gEfSjkY7+H0UzsVHdmR++Z2p3FRTebBocoARSGgvOoZW7
m9hBybH1cjTNBHS1TF8DwtJjfCX7FhZvp64dOOBynq+yXHvkSNawk5xSguqHv94o
PCHK5UArFWVxe/Y14lGhvQETXaPngmJRxMeQPCgN+vGm6fngDbYyibRcA3CcRH3g
cFj1ubDD99ZmLOhH1msmO+oSbh4YgWHWKPsPpWoJyYj4yCukB+Hp9WZRpkA/9Gxf
FHZUR8suYH/YCs2Ygf1W6SumG0FG0dM3K7PaQ0MIHYP0glolKwOWMv7tGoFyViYR
UIb6I0G5pzKxMQNm28a5lMBCOtW+szrwL0CiGuf66bfkcpAuOtv657/GG2DkbjB0
4+NzMg5AneeTEsk/v4A5BFcllilDj831siMrnT0Y/9vGXE6i3MSzlbTkSDdWj8do
fckMCijhuXGpm70F0H34CSM8cVrP6VYgeDbMbi0m5odBpICggbG/QCJQKQcB1+DR
2uF+M8Gy3k6FsnbqhZO2VZ2AOogGWerXU4xxwxk+5VzPknIa3tKtK9A7rZiZQKht
tVQVF6u9yjO+MYFVrafnrYAZPfozNYUzOCheC4U1RZlmEPvGhY43yKbLuPsZKCc/
sQaWEmgqstvUZ03FtMqJfIypO5yiWoj43qH+DC5tJ23C8Eeosd98f8oX2CdcmuNk
Mc/qJ18f7bFVeUyFfL/Kqi8l/kBuGefH9peHoUrCINYAde0dFCLceES2NQCEacBa
XS8cQrmxAdQBjOgwk3LUCUvqLBUYiDR+l7B2LXavArvr0uhZEkxRng57XivVlCDZ
ytIwAgUo5BLOOQJ8RkqXcNHeEqFN4jYM4cYQIapAXqowzun5+0j3lc0Gq9cKIbAE
eg5Og88i7Lab8Ll+riyzXrZUCiAQWVszCuzBvVwMybN3CwAftdliTH78YMy8l1mA
xo+KyBMF3SjlL1wAZw01qkGX90lQDcD1rrpDQt8OisD9dkK8sJS953XyPHAVkS6z
nuvxMic1XWka9D2Oei/0BNhVvrUn72cA086lFYgI5fj7HhwIQRgb0bf2YkwNyDKb
h35gxRZPVbQdfEL1SFk+H0VsnnUpCChQKzdGtTIWU1msLhMuIB+zXh5R+H4A/Cjj
BaByuJrKxPJTdFaDWbEAjs9IWMhEAm1Tg1VVrw1Z78eu7hVqkj+5NbbsRvfW5UFI
GxoNT0G94GsIiV/2T4CXn0WGEJ47GQAeK43flHPehe/KLVcCxv8PvWr1nQGAbzsc
hCQ1ZtjXgFFfBKtvhEZbK4CkqAvmsNcubikDSM5EdDBDL0cMqABHS8uAckhQoiZw
dddVSOgtJDjFcjRSHRljHbDXfWjKhL4Qs8hHDHgc4mhivl1TI9WuEi2YHE1bC5Uu
8AUWkpttKtvHAIrDwJRABRVtjDvRwwSbUFpVRMccw+7QBG8Ug9C8LYKgVGHlvcuj
LIleyabOom8PPJwcHtdRnulFjW8sAqJbmVK6rV2bToZN6pTakonONjcF9rWDElmJ
cXr9cemKJxa8XmP6HpRyXJvz57vV5JCWkR9StJC0QGyhp8qBqA/tR86L6jX67yKM
OCEomqqF4EHFALWaDGBXKWs5tard2A0eNDMmenCq8TVKfZ0MNHlN1T+k4+N+r09t
ggdmWoLLxRuzluX9kpYaY5lCsJlS/bgiQFUyNFhSDbCi9sPL+a2RUuJGe1Gx/zoR
Ys3BYg9NQ+C6nhQTg+uXbPPd+0Yo1kohIH/zF/gKPTqZzFnHhGiEiyf/f10ndWV8
G05yZ9W3hcXibUEMZedoA7H4I2EoIHjj7aH4y7aVt5YNBwaKMOl3ynxOx5rNiWbP
daMBO/FOpqN45fyj84J1d+m+qM9sQcrfZFBPHGv5ldoXYL5U2Yt7gLo8NRKQmpQz
zfVoo2bQlldYSWiM8wp07Sh0u8K7OwB74trJkSRxfaLG9ukcJrEc7A6W9g6ze0K6
ZTg0aZPiEU4Ydr2LYn+Dm4LyaXQfE7uWpehRBXU+sUeUwoILObkgJiFRz9x6trKS
7VAXKkXYE7pULHzJBWrNOcaXQDSGxUhhqL1ZCVlYWoX/lptKgusUBLvlLaGGKwIi
W/Ebvssy2CoeNgaAFfJQwJu2GqSvbq96pTeh+n0skzphtlI6QM+iwzaWChw2PKmB
YJKJlnYkjtpPM47OmKDEoN4VQWz65aGZo87gzst3fKT1jW0w09sFlrqmAgxYa8we
JtoBoO/bbksCqr1an/0tPJhaX10DxAMRHfamkMYmTKHdenMM49KGsDToVqIG+fHi
KovLiDyjcaKPvEzNZ0a/AmJz1v+LZVt1s5WDcMmMPeuRr3qhfquW2d1ERJNy1mhG
mGlG2J6E6sSGvNs9IjIVlmNM6SCENdNk98igVl+mobOdVr3DnQMEYTw2HKHzaE5h
Uh42VaAnItbLIFAOLpf3+gxGmfzhHrLoUmnOtcKmadfudjCPYaYW9/IMQvoBiFGp
LXsKGwG20AaSa+Vz5lS7CQGmeDT1BwvcFh+WpqcKPH8NbMtt52LauvZou/urkHo2
2dKv1IF7KvtS/KWfBkjmxeczibDP1bMSSMU79IOEKCOj7iVOuHsQ9R3YQpKNno7k
kcWKZiucJyRYqzS7ebXFcqLbpiJBWBlQKljCg+pDPQlXjMU0FquDXMHe8MHM5zSd
Veo7hUJhO+Cxn2a1Um/yFMtsJSbtZuF2xmTIfdVjow9y1IfmA+gSPRwFo60ur4vq
Q/auBBuAa/GXnLnUwQhJnskGPHXGseDHAnT0lc3l1wu4WDVr4ZRsr1dlVxiHzYik
1Wqkf4pkh22NiarkeELLplPoyQmZ9Mu0fkJ4YSvtlv1p4Yu47z1AL4P4t20Py+ML
prVlAOql2NOmHo7IDKfPYNZyG3rmuhNqmR1HDRVQ7qdQgZXQjZhPxaAXu9APZfjq
LIvbr58/41t8pgfiP23DE1Kc7BZWmGiNVAbnzdFBjwyX4iWXk3JHFTqcMhh0hReo
H7b5I0DsE+Y8Gw8gl/7YdRqNB2jNmpignfJuLvxZzTt+ijvAdIWOk/H6lhi94mRF
TVl6JHjHgcrIAh+yFbg9SAjgzk/oW0Q6ooze3HT6aCV/nLvh5JMjvuY14AzY+6UE
HEdnh+2EdfzEuUgO78jHwAcewH/qylLzNFOsyyeSPSE0g7LrOX0nFxmj+Z1aq0Pg
vbR2YS1xZpjCDdzI8fywW3GIbWo8N0vdm6v14KhZMzctaGZWqytkqs7pILsN0G8G
H//NR5cuBSZwYaqNnMm2+RNGck7zruvjR7ma+yHxAh+XqlwHaI5uQt6FbTf1qilH
By3EGqXm9ZLgMmeRaMb/MxKZdW+M41B4bFKKibv4pOe1MLDqawxp5/BuVa0atJVf
x/1DtCUACDCZ5E+FHbKlesd1ImleHoKNbIfMANBUeqgP0Rhmh/LkCgZ15ww/0tL/
8jqw0/yTqPyocVs0NSneS0TOyl6eJCa9V2Cw6vwmov5GF6cOE4smM1j2nrCrlGZo
07BXjhivXhXyJGk7Fd+PmHfOSPkmocaMesH3nZ5L10584V6lfPXA7s1ehogDox7L
r4QrpmO187/e5VZyRiZkDQ7UL9QjS2HQ/dVJreYZITVTqPsTcW5Ayj+rs1E3gFX9
eDzX09+BakvFokDvvV6nvOXjEO1Svlip+x6j5foPA0p3jW7ZPoiNobn7BePEFGYU
vgCDRBCp14kWIBySvL8tknUAywDi86t6VT6Z56UXOZKnQ7ABgmToik4QhTLYZ5HA
ICIn8DI7Yu7G5lT2tS8Fg+1q+oAbYcOfeflMeK8tvEzpVji6eF+qM0MdqUL6FB/s
TF69ao2s2pnUVkzbJxTbEfdRTEvge1LI9sYqAtaYEhJEYTvnNiX5OttpB7W/1QND
gOCU0cMKKUef+XVpFUnury9xJoJXCb9x354BKjw0muOrzCqYecuycsTDSLp4lSdN
7ZoNIqopgJsJl20jN53nmWdwuD8WCfkCG1nLfwc6krKMutbm3Co8PQiXE5IUthl3
oqHkXqD2CF0mGPcbli7FWpxX/xKYgZfL2vZYa/OT1UPfGQWlpjB+8B9xEb6TF1PI
c3XCym48sjdqBlTysVf6FxaIpmNEwByrSZXC/4YwbBXzbcPlBgiyySdOz1+RoZB3
v/nmDZ1yE2MIuBx241Smt8zElVWohyTENOYru9dnZ4clKZ3z0S54MAaDPyeca8Hg
PHV8d/pANJEuiAXAOYH9qQIzHU6IEk+7mQvsdBBmio3Uk2Qsm70rNcTP+qx+9BTm
CKEzpZ0rZ+u5BHpPkTqWRuyxxGo0iCJzV/11BXMYR3YsIpgPEdhCUnp2Jj/+PuUS
PftYcUp9Ga2xgjNJ65NoIL9y+zLca6A4F+ILedQOljrrxPmjh+KUrZ+AOuykjg+t
PSMpBk7eLtPMCnQhSmL2Ydb93HsqQjZeVqgIWLzfLl8PaKv+zve8eEsoT463pL6v
ysFRUiwWhdTaILInvFRDAKHjcR0sMmM0ZOj/v/q7E9DnpD/IcbxsrqTCK69QkD3t
7p2peLl4eNOHcVYUnWaMYddyYRiQ9WljwvaIAAlDW1T8dZHza7nSRMzASXlfCkpv
NAsWUN3xxkQx71H0HZfLHrnTL7Cka4UhksMHlnhVmVwQP7/UuvPxiidAzksF1XjR
UMVV56uk4gpfAJaH0t5SzCd9JfG8D3IBbmm9SSt1yBZIEsAWwnIJ0ILfBXWRmVbb
3SQs4ThhqfnACkBMtwDxNQcTNPf+W3ouo7EL4DeNlYsqDTMhfd9DbgRyXnH5WVt7
5up4PAjjTc0qUjLLNo07T9lZWXsXrv9GU9CIgT/Sw7/T1r3azQ3reUkyKSkxxWox
dbzSJXpGaAKIVPMgvd794Gmw2gOB9bp5s8k7kQFHtUcwQrJeuwXCFmKBUIUKRfCS
QNCo8vFhuoj95NGHTSYrRRLj/y60zJ1Wh/GKHRg/NKhDdPWSXPz3HDnJpgrgRY+d
44cX3kqrpagcj6nLkoA+DfoyC4ieOLTH8Yx3b1se7GIv3lNGQLJybY6XHiInDt28
89S05fIbYib1fcDmbYF4MgMtSsv3lWCVApatpQOk1mkztEHiYl4HjkZGRPFMn1gV
JbpkaTdeYhJr6IuyPRp/DYAv+58xTUUggvGJjvWUlPEXVaoE1K9r4gO0zE88ET59
yVBcBWh0+GhTgwy7kdPwmd0P7CSU1XNw6tGMy+NLRhyHKjOkYoqPSTL8o0Oj7Cvh
G9CfYPPIwHJktjgR+kWVVAAS3h2M7TzQiZnEP4/QHbbMCArcSWh5m6BM5IiY02Ti
O75LmHF4hLsoDq432p2jujJj/fJ/IewQg7NlTyHd5b/mS3VSr4Z7hKEoDFtDOzpA
jh12xCr1oOlXAUaC+Zs8laWWXQsjJKZB9GzTbLffW6kEtJByMgZBHrKJE/IlRxtW
YxQVOhw08SfEGuQMoGX3ZoQA/SOA6/sQwkiBm2yQwVtjOEhbWGHPnEaV+eGh/87v
bLnZn4DMLpXFpLPibOxNLqkOUGPntDFHtHWz3QjKiy6biyQ2kmhoxedZVWifWJXF
AjpMORn6yfM+74TmL+zuitaIYNpnDzq/OjdrGu17WEbOav8YEp4/P5B4Ay8A3nfH
zLXYGJLwEZefd6dtB/QIutQw6QFoMn4Dp6X+Xk0/ppiQSvYsZ8g5oWC27z5UnGD6
AVCdzlm/M9lhUVHKq09Aiaa1MhAsNQc0LYlNPyQCAoOMJS7dHPKlzD5E251dyRu4
FlqBaGPUnNdL2cP7voVcrLU8XIK23ZRzNx8NCAuNhv5/AgK8wjRbvCeC+Ft5MIki
YB28FibBTcDSGKzEgvGf1wFYXCA8SVVg92SSkUwiWbmlvREe5QSsFIgwYwdQzKaA
Czb4C5y2mICJohK5xnGgYebv/UyaZxInJ9zItrajHWmw+C6arXU8BlGeB2FxUjF0
eEZmUk3Xp/sgRRBfJE9yy1hPhNI+Z8ehEfgODxx0N1A9yiOQ/D2hTm0yJnKiEjVh
mB81cSRkYDAGDtAYvG1WAcxAcy8VltwaTTkkVbocCg+NFBHQqSszaY53l0DhUPjh
1tn0+xH2kcwMygwo27HPWJoX/1eth9BOzK6S/hH9IyaRhaJ7CRv3DFc5VvQNjjT5
tJH+P5SHq4uMPSN5PJqoJx0t17lb488AB8/UVemWV83bNwcwGL3tkCrMlGzBr6fA
713KtUzmSRB822aXXOd4INwSpMjlZgMl4TiSFEESNu60isXpAIQoWnNzWy+LIaoE
PYeZjWr4co413K8C8RlyqLy+T04ky2amW3dykym5wJus7IDIE3CgttqI3H2Z2jtQ
uNNUL2ZV/UOQqT00e9IaoHCcjYoIdUYmdjR3PdbTXqkgfGpiZO739/esIS4txC3z
K6nswT8Rkc+M3/ki8jmDcZUJR5iFSdes6LumofxY7Ex0L3dE9MtM8dm4GGiu9mDK
l4owSDOLag+xtVKkZHHPjFZ7nXiZslQhT76avJMeB53eNPatN7Mek4hIjMgux08n
NtOxKh83N/FMmfPUVNxbH+8zq7QXuv17Hdx7tBXbWJCFNw+cUyqPKjNcCKvkwDLW
GDLw1Y2kHeCxSqq8aXJi9yjvYzINar8wE/cYrtaZvII9m0iWzT8ITybFP4P3vAFV
ZB7WOAOiyPk5Z3L8VRMs2GvI4Hy9z9Z75vwOOLq0RP+2TXx+0JGJ7WgayT5Q7BRt
byD4RtdkLd5Er1UF/KXDCfmqu382Ie3jpHtarNUfOBFkBo3cJOoZwe11vNXPMNXH
R0wcrPTO/LoMHd3OrbQqXOVntK5VSle7XaCZBd9aiowu49Yr6Lvp9awFKiNzs0Lm
00xeBnJdhFXQCwHenmHL/yrNK32vWU2CfAE3bvhRCYVomjMU5XwKMQPnx6Vaye2O
v2ED3Z5gfVCu9OPq84Gz9qUkmwdN90jLYg1ZX2ba6THE3B5OBFk1Ud9zx9vEFzgo
lYbrtZleSuJnCqwYJzXtYVz1+J6BLQZzLxLPqt5bi0vZr+jrmxmkgT7/AhxHY6Gj
7pWPcbldLghjdTJLwg6VaMgAr7XsXV90QYZtudtzdu5qUYzkrbLa/ljUzTXXYDhV
rNJtS0iuML2QbraMVBKRM1E1/5/au8qAMATemU8MP/2RV5CpxrLYeemVUSOlJXye
NkeGMKfHvo7XrJYlPWQF6m97Qu0Mo1jCMpTIgA5nqZ++q+++cuy10V9eGTBz70A2
TO/TYBrIZcQFmRIwpcd5b47vamD0rgygK0sF8s1N3B6xO1RBLCslYOWVYVNEWkey
nC30vYQADYgBrA5gjDX9X2GFRgshcC06BbxzOQGaF5mvRqCY4+Ji4OCf0BNOIxur
N/p3PJZ32GEEVOuxWurZEoDGOcP9il5a2RjSpYVI84oj3g7ggCY9az/vr7El4rQe
YL4KQEStNe82lEw5McyZhn3HMbP2rwtTdPDjvNDLu3fd/e9j5otVeXVVjyy2UM2c
AwIn4/EpIAFJsXJaeSzc+11Qkd1x7rnHwdvpHi6XDVod94UnczhK4nfljPxmqyXC
DkAsFEjen8ClycER9Q3JPpQHnIz1KSw27MuWdY0opfQu6NLy9DajCZ38NRy4AXRx
Mu+OqwLyZmQKs9fyZFSagZ20ExSbHtHVFF4BJE8ROl5R15Ys+LaCW+4xpEKG/t+m
j3ItUPIO0XtP8xTso+cBBRll1ectVtyOQVh8PXsP9lnPfmOLY3raPcBkNtojReNZ
zDH4lUw3qa+vzRWDkLMIVPAemv0idS9z8u24OketWbCYfJ0+0udDdSYzFb50/kJ4
cJNYId8KUUWBSnqH3BOJZMwg2GLVRpxrlARb/d/LZXUbSlgdyYKCH+8+pQH9uNia
rcOzd9k+kU3mIE5DO7CMr5oc+CMIhajhX3akN4BmWX7OFLfnML4+nr6+5EDcP9Cs
hbaQwX4LJEKh2lp0tn53HF2UPvvCli7rMd/VSZbIZvKYCscioVY4bnZy+piTWVf3
8MjTxgOAskyJ1ypR5ORXph6M89MtZNoPYEK5xGZruFRuRqK3O7UcXlghqD0aAQbi
ZbHKoM8X9moIa/2RWfMcT+idscocbxplR9Z/u5JsfnrdxsxHvLIFZ2prD9u6OU+W
zEUNntOjzQ6mWFNbN3vNhkfNnDcui74w0pHKYEbdDmieDp/kH5BHZmsUJ0V4WVwA
Mnkc3JwjWJiiAIBTlngENp65QYCGA67YKtDLLI10CWva6cY2YNSrQ1ypUzfvrd7T
+n+Cpr/5tPBwzNinBFbBiXiPWVBQLOC7kpPpN5OiYBPsybCLAptfjyN+h2UxgRau
sons4AiDRAno+jk5VDm35iIoxWzfz6T8b4HZ67wpJfaavIzQj2LJqdkRdtWVvms8
7rP0haqwgfZA7gdNAqkZsNUQuurGTiDV572Z7olW1vwLDsTcxVaHcwA8Tepe5Iow
5kyoQB7GfjUZ/YpuZTi4breypE/izak9gKms3xkZ5YsMKX/iA2uFTDf0mdFZUyWf
fMoGLV/NKvhOPiTqCqQax/JZvg/cmAfnG/jmBPSDnS5hJEIYobdJaVzBj4SMSY52
OH46Wi3gP6fLCEzJLIhSUaMcu/pL0wJaQSIV3+kKdIm4xaYSxoy/5T13TTn30u6Z
j7WoyUiWrDHldfBfAs27oKSuzcZU3u1smJeL6Y9XByxAv7xAgBxku/npAL7dvBAM
k+UD7JXiXOEVob4FywLKb0Uq0I+/iyU/F9bFyKxxPxgNyOdGYhAlQbcjsZiM1ORV
kqbBPfWaMJyHoURoZMOm5HpGhMnfQ5TkuSldl119Q0lV7BLBOWnzGb46GQqnZOxP
GWaBPRVVQWMzt422bOn/ufOYGs4qCPhVwGI4IetYyLF/FD4kducJA+iABQH+OJXH
6nO1hEOYeW/4kaXHPAHxgFLkjFyrwIlJKhlfcIXcAS0Bp4IIONFUONtkULv2SUpu
2ARqmdIExGkM4BwMiY+2PK1BwmRdfwapNU0jcgv1EZIiTVslbWdMJc9TJoV+ukPs
XQWeUDhSgAgaB+ODtS26ow+T19ySS4PoRzd7CbkvhEJQHKZfZqv6N6T/vnsA7Mus
1nkVD/CUYYzWyOiCuA1/Xt6Se0omG+Mg/BJ99qU7aKCJNWtIperI3+XmVltQu/Rr
LS1JyzdfNZ0S85BH0somDG6X45CtGWaMGzB/IfmTwoe3Zy6uiSe33BxNXHnReXzO
mLLnuVKSlPw3kgmxIT/Vt738iIF8LHtfGm1c5RjSXEVwkWFGdUCaA5pv3lccIWM6
4VBlLZmJ5XntjZIGX3k/+RVbOcnhg7hZKYMMOGc7rM7JjZunlHjTNjxrfZ4a3MQG
hun14xTmMMhtjhayIaENMu0J1ooRitPzHCdABt40HdBWqiyV8ANoVSvqnkJxx7zk
QZaunnLEmMJ8HMAyh6T7AIs2BTTAvBTEA5ASfkFvYd392jTKxgPcjh5Sw5UJI/z0
kxpXNsxuQ7eRS5cymdD0jXsTbAkA0YJ542o7BKqTaVm4GHmzpCRdZBfPpj1RsHVo
1v804/TxX1+TcjUE6JBwysYhSwFPPJUjvRrMhasgUdu2UfM+RagcLCaKiJ1CH9mD
yUPWlTtXHBLasVOTgGOeuZNg4MqZ2sNJKXe4HlLlh1nQPLfLvVau4pp/Yx64y4ng
LEXHDUviLcw1vbkyu44sUOu0mV9P38pXEgzyfaSU+OPUN4obYYCLrGjUQxaq7dl+
+hfgOJNhZZiDRY0UPom3rFPJDvv+ciZVli3n6DRNZtR5czX+3cx8FdvItR80Dt+9
vFyJ8wV4eQ84KNRRKe+dfnn9+Sdq311BbSiRkmJsWAWZxY4ZBAyDC09UDqNSmhGt
amfqGKGJ8oKCmwiQ3S5XF4x7U/jrIvha5l9huDnfl9Y89E/gIMV4FVUdwI0AaNFk
91GdAHN2whFhsHCakRNJ+WlrKpwW//Za7InyiR9T0hw8e/ooQ4Iabq+0T+w5KBCG
K8XPu/kXtiyF6FES+I74lir4Xxn3z6XOJjSpuEv+2jfj8F557xsoIb0HOQtjDWMl
CSkhZWsDjCzWwFQnu3YVPBmQFtVrVrAQaIINZCG7+Ij7IwoJoJwjq58mOSzqlGDi
+1004ubTHfCCmjDKlIK3XimSzpyVBmfAFPvoGDcNvKdUKkKk7JhOfmCbeKyKttiR
uJOQr4pH9zvgfc9g5fE/l+UHtj4l5bV1slnZ7iVNYonu+ArDmdXGA18NcOSmaGu3
xb2cAtdIavZY38ZwbZkzqUiUMOpx3eU8CHIEu/FHRQ2YOtqobYALoQrELPOzWy9i
+YEUld7VCxcx4fSJLMne1AhtH04W/kYEDFoq9irNyqHJhvTot742dBXhEZ5y7jVw
soCooS1pnVrJpd8yXjXOS8F0EU0fdDFMxWB4SvOIAH7tTI5UZbKafXEAkQ0k9bQH
PVfGuglHPe+QUv0bOtLuchdRNEESq7+vz6YTUhHJyBzYnS/G5cHUfQQc0E8PtQdU
ZIXC0o8shd0elP9rrXEL1KAjgj5HjLD1JCWZYe1Di4pZ1qrzn26NsBvVYeF6qUap
vhT1dR2v8U3dNLPl30wXSlHqPTC1CVI+o3Ul4beeZ2rbHiy+KopsFfxhMs3qCg5V
sM8FZzBo5bXBSUkNkCd4+HnYXb1OlS5aztnXF+1N35EhTGjzTRiRFACGmCUxBykg
Aw2YVdPmyJzq461VfkhLKq/ITGsFsJKhsld19uZ6DupCnLbUnLeDkNixbEIA7dcr
sE8Ue0iaa9MmmEexOHUCi7jTYa9tnB9XuMtMwC9uKAyNvnkffu7aIU2dlgEa7AQx
ou+F+coOiRGbAGvJxf+jtOJql5YKVN2QqpbbDbdHrsc9oxw9BvJJJI565sgmqwdJ
mVrcPvRD0CPEhPO37kwN49Kmt/3TMmbWPCYUMgYSd9LE+0dvTbDp0T7lRjzsMb3X
I/wADOy4dVwOCxVgxvjaMqFxqd9VBkLLndVVxf327to0XZS2tHc/kTke4YgdKx+W
R4X2B7bNN60KGdUVS3sa8jtnpUXyuQ6WidwVbcRrh7hSCBEezTqv/a9x4TEL+2mw
DDI8knpAdsRc9ihnrA2QFBCv5o6iA2n1xfEJGdyCgTnkIUgWZswLU8GXL8VBmbhm
7knkOGg7eFIibWpBK0nPKkbyLTRjs3koErFS9iLrf1agWSme1TpSiDtTcbzlomvM
HT9aGeuJh6ejwMh0uA2YbwgRZQryEeYx3wD45jSVbtv0rBXocuo2ALbTTYK8V66G
WO4o2XcpzFrjvzY1SyGqSYOl3sYO+Et7azCSHUNPsHUgPJ4rmyFfq0rGQ+GgyWbw
V5wGfTuxFL2VynhCAwqkJZrr4ynjUVQIEwNyST5v1lxM0RgP+oGLGNOIOK5b8h57
+MDWjCQ3elz5XMCk6OFHLdk/qAaG2aNJhiThpWFO8psKSIthxeVITlzbae5Fr4Hi
McuKO0UjSts+neE86TWeGNw5Sg9kLFNFJ6/zPDOH/Raka3zidljCJtwvg4Hka0Js
a9ySphgreX6atV+mdqv3XyRt/ggiji6O/Q6kvt8JJgF5BgfpbkD1aLDcaZnL6R74
rrumQvVRXml/VK8zFLaITyORyb6ivVyKgEv38krTISD+WZMGJXVGb8EXBpkIcUEu
RZ9fVZSXwGj2G5EfoKtwCTdDuGdt/MgoPQAWAbNX5tnfT2wFxFybseytL2oFH8IY
7H6ywKWGZh7T+g1/gYj10MkJ2qnp1A4Yqi0kE2pd7T88u4X+XZ24f6Jm8nxqVZGk
p7lH/Gll0xK2yBmsH6ZgUbusGjZvXsZuuob+3miEC/fUSLZr82WqKEkr96XnUPhS
w5bHvRACyPfIytIjDZExpeqRqHhd8Mj6YldB7keIa+dNf1OB+49BVe2OfSUpbm61
uJJj/a7hTt3JXrKtvyN+1P0tYTOavPmlc5aS0jxqS4TyXX7zCc9Vm/8m0AJfqcLx
Q3pALi7Sw6Gim78OYTuasGLfAlxLE9XFLMNBXlLqZ5xg5jjFyyAWi8slkLg75HHl
GQ0i3T51axSK9ja2efrzc6pUW4BkiVt1R+o6Cxsp7KsMpB7BZYElvsgBT5fn0CBR
yTYHZfqyst1vwzg4XNIp0Mv68t0hwojpTIc2CnhlhcaiMlsVTXIrjbQY4X2nv1Qu
zrAxtXQaVAjXBbLOxJkWe63h0rZ6JfOTUVETdXSwgHeTWdQVxRGVCNcGDl7P0wkL
5FbFlKGnlk083sSErhSP43wbEW3ByO53lq9JOYmgmppKjEo1UPn6TMO0XA1EGjFy
XHY1J830nCauxt5P0XSKYPsYJLHjoLN1WhYLZhQsclodQxH9gD1XMSLBtZMmUjMI
zI73nTNa3Dd9Qp5JppY8hV+U39dWdTS8COinFiuJ69/2yl18qG45LAEWCqO/s2xK
YDOgkVNUuyjUGS8/gVC9zZkeNYAd+s582CZDmjbQnbfUnxrCoa9YTviyT6HFx6g4
j1ypiqt5dZ3Jlf/NtQtTUgeWLrgM0vX0DOohmlvDnuU7bC/DAFMfYvjcUtH7OPtO
H+dfJx+XW+cEYSqbzJdadbMoD7D7ToFFz49lU7zZcOvJHuS2t+UP72O/THqASah0
DrKKNMjR3GCS1fAf8U1QN2TqSflgteP5sVs5jpvMmKkfuPAvVGIs1qvqRREcQMUI
UmcA3hP3LiLz/Tey91Q/55d99WADT+4f8Jz6l53HHa34zxwmAIqHUH5JVhecqnVh
6iOi/GYCXWAY/TncWcU4VUeCkJyhbMVRvkXUd/uRfb4H3mjNAcl8J+5tW5Ev+GMy
nZfCgnTkpgLxrsqjCw5UD9KwimoSMRedrIDwxIaquWjzWYTlLh4hQIB08ng0y5zg
7JoQN/7A/9XcPh4EqCSyVDirDxQxvSp37TlKPcm/z0PQP1ZdnaoUvocjxVV8YPKU
UA5SOZ0dLcRLJDyPq7he3no/JPCG99RyrAjXi4UAZrt8xLresc+6zpNWoHYUjRMG
XbRfKWFg62Q8KwEpayq6hHRDz+0FaLWQSHtK4Q25sSb8C/MS959RqYmLapF77kic
ZpgoeN2sDqI93A4sLUanc3H2Ym8xk3hWjcoYtYE1zX8QmZkF9mBYZQ7XyECEo27e
5eyyTXQLHJJeyxFU1fw1W3uG4pRsmDkjie6teRIG8R/AxVXEdYhHpaJ0WNXJ/Lb2
ypgrLmqmY3AbbuaSkZL+BEp13faY5obZlp8bMKqXyRvhuX8jv1DOUvY0/YLoktAU
wv+litwkhKRFwFWKSWDrqrHrTBaVLAW0tqf8veDJvm5I3KVT046IsFijNU/zbcML
OHEqMPzdoHyjt5xsvr8P9Dmn9zqtYU+4peR4BUZ8v4Bkv8yDaU8fez/l0AjA/xWr
6ZgPGxCnrd+3BrdGbNNvK4N/fLN7lD8dGQExlGjKt1pfAy57eAF545mzGikSqRP6
k4To3lqgFmz2/qIz9IHlQun7rTVIBYDvjpPxX4gU+jzx9f8WBXuXSfkQ3jbaKGdo
IwyEuVmpiC55rXC/n69FkLEWs+iTqHFmhtUBLz+L6RQv1zhJKDmq7WpE5tmEGpa/
ee5tA7kZSMRAeP3ChgVTgxYfJxND1YBtYuNKIHg73pPMiOlEwxHcwrSJcvUlLzQ8
885gEtuaq3NmLAKerFHzSGBBItSYEQZUAkf2m6GPfi7BY+MWiJUUwnJ+qJyzxik7
0DQ2G0eBCMnXh4IQKNrEHnYXwCw3aCvgtlRX7wi0MfoM0bYheWMXMUWD/hhAnYUP
0kUw99QMKX0S18eseOrMz9C53hTxTOMEVEpax+/+7jbjsYt88EUE4bm5u/kjAlR+
hGqecl3Lh/zvrN5kdA3TVPwzpHmSkHHbhwT9xWNN7wQo7gWw7r5iDSwXCedXiyjz
XbnGbi2CqEYNC0fcSaCrED4T+yP+/t/UMZZAZQ8fOFkeHv4BvwNwXH8roqdOoYFv
6uEaqeF1hKfGXtBuFZfTnJLz5J/ADvq4lsbR0Z7F9U+FrTHf9pa0v1BXF06XiuhC
bq74+ybvpQvZQJiMrnYlkCcTFBsjfl+u4WQIEPLx2XD6PuYGQg07dp+mcsiKROli
QeOiXR38IUW8WTDkWRfSjU5OFybRRQhnNS4Y+UQmP5+fpVTun/dVPu+SqcvRC1N8
Mr3yhpG61aE5QAhy94OdGLWRjMIHB+Qymm5whzO1B1+Jl1X4QCE8h7sRq+kQr2xS
Tv+vSi5SGSWGLXwhs0alxB2HjmDbkgb1xm6W5xr42EH+hutbAfD/8RxKGZ+ZQYor
IUqeYIT7xJb5meodmWzinlPkkOW2p9fnweR43GDrmObrrSfg7APOdzOTqFdXWB4v
rZaJ6l8XVWj0zi1/o6YQxVTKJ4oQfgTogZm+aGHYEPbTwFMACqHSL2KydN7znLEk
JARZDP5Pedsrx5IcpMUm7i38UqZ/+svqH/FpnlpWMT48lvlgCrJH6/x4oJKls8dZ
nedxh1DhP+rXzRI1cc2YfvALf3vnbWKslz0iy8+fZCDzW5TV4BIJ45bFQ2RDwUhy
lk0qh9uaO9V82edyog0YlYkVTbXauHrKogd8BYyf8rTyfc+wogeRCtfhiyKGR1F4
nvzpRCRZcGCxN727j5GBnhd9wn+g2WE5r7KMZRr3QgGEP+3tOw5mUCyFM6MXSWvj
HiiFDsFmzW4UBBK3mva+XGCX/74ZQmltjjNLr1OdNdctwFRbvu8Q0IEYKWleFKxo
IuoekRzbO2SP+Y17wmLq5iPW3TbjbJKbNhiB0vzdasrislkkUqrtGT7eVIvk36bN
D6hzf9Vu5qoKKzA8HlqDoCkX+LzqU/n3ztXeWmsUZSxsUESHhvV6983EwDkwjktW
75TW/kZZ1BYjjgq3OMiOyiGblwG6llN+9T9HaHijHlWHG1cig7n02FFwKuPI67j8
5G/OdLbgogsQe/kO936b43gSpwk7q51mI/GidGaAqz5F+O5vjJbBNOIwgC2aWo5A
d9Wtx4dvgGKQ13p/t/wch+Wk4mOvMJ/AOpXgV26bKUuWceDPVxmcSewrkEZAl3L+
mvWrSAgqpXQyyeM00ecL1XXWKO6N6Yoo819Oh5D+3dYWY/LrL8FRNE53ITMl07U+
ol4/hzvye2RwY4OlPnegxjQloPAOPS3g0FLZCctis++UkT9SY/olMLDxzIOVr3Os
M6f8cSXr7qaSJjIgeMSGX+SWGB1NKEHqhBnFkq5tfw+aI/ZCbWfifusmZCy2T8sD
Z0tKWFCkpp0iZQ864FjaQdzr7FjG+WLHSYYfwzFdxa+JV2nKPjqYdY48cHVH59CZ
vb8MBlKJo+hC4I0pGJJ75FthwBTWM1hF1cCW+2IOw00f5ZkWMufs19xIOFMbAkWa
l3EBDBVpIeOQwy1FrdUt55hO4hh4yxYV+fj7xX+cYfctA57UEe7MKPQqtbSaaKYa
wQOThxSnnoLd6IsRJSn5YQ3s+Am5cD92TYJRF7HZDJQNdAST7ewfh0Oni78l4YYB
SGIUHtbLA5G3GcTKiF1BmWroBnIiGbaWzM4eh82s9cKKwPqHVWHjEXuckG478gyO
y33GGY3Zc5LQnSvuAWs851GChASiEYxLF9LTVSyiGacUfIC8vmLdd7n7Uz17W33N
UexmooapXXNOX9dkqvIclTAsaF81B8JvpO/m905qydyHNT0Fe6BPu33iCE3aGbKa
aTiwxfSpz3FIoZU2MWRASTOeEbZLvkHeBhKe/jXGQrnZPRk4LgxTAfIAe/hdisjA
HTAitlzE4LIaHo6ceOr83pkalHDtZitSN7uMafvGzPMw7VAtnE7vyAydcKlhnpJO
yrwrVAWBwwG6Tg9l8iQrGVvHkKoORo/iiPgm0QcYy54XfTpYNo6nFFUeaLjr6v4g
g1RUu8f5/awYqOpfxb+hhyTwLGDbF1xohjYTLcdigpPAg5uV+rZH8G54i3tcmABu
zlOHS49re4jyNo4FB7loXRtICtJwdUrwnwZE1wkMHDQQUE5YboYXNQqxWh3KqmbF
DFquUIEWTqpX+LyNCyw//Aa6D5CONJPj1uo37yK1ERgsKpvZgkQmuMJn1Fwxz9AW
z9XH5g7c6lO7rVf8PchYvwS3RcaR9NSAoBNLuUb+0ycteNY0V4JaV65mqJiUqEvR
Kz1hCXB07UasPD0VAMNRpBgk1XNbGOsDcWWEIMVhiakfm8ANpwoc+n8PiYTX0C+9
ygn+pyVVvbGas9EI5dmhICSh1L7g8uSJ/XdTCe1zgJJlYQS+eJCtnSZYIGhfrpZq
8LBA5a1ngSfeQ/tsSSDcPSUvvrW/iyogMaa7n+3PiTlEL78iCEeEEKLlzw6aQ1Fq
wqC9CeJiOl0JFSHHQl469/WZNTYyELrzEx+ke4cfr11hy/hjnG19k1FSHK8jaa37
mTB30Hel5OtzKoPfg82JRPur7Dipib+yfp/nEKEdov7xkbtz/wYc6lnnUk3o6Q2t
Egmwy7eSxfP32r66pi5y5yIObKPPM+f5pq2GJ3ArHYsyZJjYn0cD0EKOEmz66bGl
D+peUp6998ZsIONPH4xWdO792qemOYpaJYYd41aBXU4UK4alL8UiRn2WT9nOc+qp
dLNdAnB7u9Kc++TIm3D2+cGjEj+dMpnnV775eJpQbJnlot8r9vmaisPgj1aTqISl
NN2xFX8UocS9ZeG0dhnRo0Cd/MpAaBpISAn+nz2se+paisizHbO6Q+y+OrOygs/x
mqiJT0BoznmngYxu7LaAeihbuQNWTXUzYlyjmOs9j6OPDKh6rBoFBwckJX4IxYJo
Wf9B6tGWPtBy6aJ6M4bQ4tHCwFrOKsA0SfcQsrhbG1RCk8lc572H9nUaNfdGn0py
ximhBWLX/D5jWYXAGDXJ3yugAxnMFFmboMF8edBqHvWhJQJ1ccuwOTnBin/mhpPK
OOZ/GBv6DkGT3ujdviEsEtK4uXR0YLF6v2U/KUnRtn0Gx0vKiFGbcsMdHg4zB4oO
+Y3/v+h06/BPve75dk8Ej7xUVMF6g7JVftK3FP02yTCe5dqeg5/oH7C9HWuyihVD
Rp5znbsD9OkU5EcfaFzw00tOu4Yr1Zz30jcQIU/N81vU5BI5EOW0dlU6aLrKmANp
rD87M4FYRnYve1GPr0ACq5hVEfTyqd7PBnq7QB4RNr5pJDmNmcSU2dv68oKvzwIN
Togb+Jas/i2QB3WUkBhe6/l3hJsmwsExmmkU2FuUkqQllNieUKCt2n2OPjSDPD1O
Z4PAEYpmX9puZm3k9O5PE7H9P0X6RMPZ6vcxOpIM/nRI+Ah0znc+5MQBdn96JgcE
x5OUhzE26IfjZlfinRdH7VQCX7M+hI+RuMTm8x8/HCjxg6xMcu7rggDlFl8gw5TF
doXJmnPpm0hWVeZPBN8HKOnqgf5vI0ziZXE+B88xQGzA3TejE+5YuVrsFjha05s+
uXrQUN3L+o9164z2e6KTqHZJFNfkmEq0HK+29wHnA8O7Us7P+5+59v2Unzw32pdn
NCZqfHS2CX2JErhZM/Qd7hfP7nF7hGJEvAfqrkv8In8oBTg18YZYQz4P3eXiYZtU
GA3VcHTeMZegmGRX0MxbhZtog6ACo9+HKGrU29WSYwEjzvHjwkZ1RXUbSfdPUw6w
lpU5KD2jKnPxG/UD+/LFc8AGXlNdkeCuhCVZoCsnExCmffSxMmxshOHbyZIzJ/Wr
seMxPUenZH91A2Uk4UiPBu0GglRYDwsGbbK9SqFUBFZUorzBfoisYZc05uS6Vzx5
6MV7xmG3/1l/RkMAA9bNbOB8mz6uiHOU+QW+BCxGELb5ha33t2gwvsVOxSHwi2zG
76D8MVZO+pzojHRHFaeWVK0iB/FaOn2T4yBHqEPsyz6I76J/k9MIC7xfVfUw+JiD
l6ESuavnXYtJz8mTUSJwxnuGv++Wh4Y6Df/XJrGy3JOpQuCxQJw+TequlUtQxOgz
xuero74lXm6H/eqCZbUjK3vId5dMqgcoY4r2uanEQjWBAEVAxDPXZX5wF7EgfPku
GS/hH+lVCPCnFve+XA2oEpgM0x5Dq4apd7OIj9mIHXua1x+JMpHkES7PxboiGGf3
ZrBka6FhD6VjnWJ7vgXTsPWmW0uRbB9CA8JpvcaBTXMhWxqRVcIJN7b5lyNZar0l
fMHpICm0LcmSDTemlvbrFmqfG177XPr6mlwYjhYp1VTm/POa4jBTQ8g4fx6Kho/u
/2VUZzdSkTDNU07PNHbuNC+zpZqQZCAQNc7aQ1fwHHiwvZLgjsTA0K/5ZzokRgZM
a79N18Z/Fc8bR93pK5cW4HWrqPcs/oJLrh7fI37Pj58ME4zkb5xqgokJUXvnemtG
eQSsSLeueK1NHS3JGgXBAAnN9PBt+SybjREJ9woGKvNt6xgdaC5ibWoAVJoRJREn
inTwcfwNC+Y2aFnR7d46o+eVh2e4jelwiJrWeAMI+IOKF1VFs7CHJ5Pm6XEgZQQb
AaM57mOMIeaXmYogGDyF5qG81XgTVFjNHaqSkiQtn80mnLp/d4wRizCCAMYt1cmb
KeTzaz04J6o5TJ64JW8PLrde65S779g3n7mO9FKcFWrpVKp0bEOyHA7hm1w23QvC
2n78Nmkz3qJad0B9J9O7GbsoynGXghXJPPM0NxAYsrtDJIeCZ+nU0TIP1o15EBl3
DBf28sNQAWbrS9PaRJCG41QxerEu6HT92msSU9ee7ZH6N4g0gh9FbVd7P67IzH+2
2G5wqm/bWV4OlN53kGN5aEH81IjlaPs+Q/9B7YMZnPEoi4P/Bes828iWHymgW1Qj
kIeHo+/gmmBR4UnBMP2TLei8CMDaIU/V555jCKxpvBKEjgBxxzlPuJ5UFJEd5+hR
xGGwFbZMFGs8YsnqkU/Zn9nqtIKLgA7iju3mplLGl4afKMnvvHqgBEM/wnK7QFs4
Rsy6/vV0zDDuHJz9WyEHFLmTHCMrQfmtfAhkbuqzLbpJ3csqTJwFmzxW2EObCGhw
sFmV01pV4OIHamQwMHS7/SChfXsz4/miLZPt15/guLcZ/HADWw1gMGGRtAL9MQTD
XvO8rUtRihQ7AAwM23HSfptqvYScJjyfXld7a3iULHkIE2efVykJjqkMueqK77FD
ORlfNJwATLrHsi7QHHndOYoG7hhJItD29NgsVl/9nHHN2mMb3JwUQUtMgBlWzl2Y
Vf8GgZAkgfpInmVIEhF08uiTcna0vccSALyoSlCWRBFb4LLc064vNCwX+h4KczP/
q3mScbpfC6lS4tb2cmd596lvlbRlLQQzuNjxgAuoaoH3fwEcjOYtTA1cYRvQeg4f
KzDZaArLOZZQHsZUMpc/o9NCT8vwx+I5rE5LB4sjSsY7MXbOD91OKeocHPqCNM+I
Q+4+Uk7v49yH0GCW58P5N4+MVFLsL+RlUBvqmF5jDDAcWAKtJWKxvJx2BK9hxGp9
YLIGFshJQ+7cnfy/SvyXMOHS+st7wEdhY8LZpap4tvF67Uc2x9lf85ZuB2q+RDCt
SfAE5IVteJP/a9S02+jjytApkcCyRoK8QEc3bm5c78k/D4mOu+N9h5EpHhFui/Py
EvUkLwKbQkYOSl30GpaNTlZSG7KACzlhno9cI9Ba5K87cMOnfRSxoGrjL140n7xh
ScVa1848iOjL1E3JEdKRRaMxQIrpHekxj5vgUAJMJDQMVbUa+fVHDpL77351jn69
roQlOcSGli3F0QmEnhycdXLPWq2b0dVEegWs7M50zIO9nKd6DMZOyTaX7k/khz75
rchz1TNvQE8kChRb81Gi8hMr1bGXM4LSIz4LULyWnz6Y28DTX717YwbojC8EkbBo
BW/8vsac1DK2WXCyhiGWOcLc1pAU6sU+PF7KiRdIh4DbrKZOxfHfGR42oBNiHn98
d5KLAumkeEjWAhVYVxuIcXQ7uQMy5JjpDldH5jbq1+tJG26ssDpF3/J0fE2xQXyA
lUiFfnDK06WLFhoTGPpZciH4uJAS3NUysfTfHnDv4QvmJHaBYwcCU8Dntd74ihqa
L2tjs+9hygdXOWx9N0Z9TZWoQGsblzj6PCBZsETsXkF0w1LF3N6tZXbe5uw5AQWq
CvQVHisz8tEKlkFEVGMoksUKE5Z/xs0IVUzzAJaj3Misb+5yvX1DpLDiAhvOZcyq
g1L93gDTBS8HOJiiApcbLEKMcCCy2UOKx6vtBA5vClhEyJIiV14KFnrRN3Nc74dg
OgNlloqpS1o4LOvxKrRp0X2KR1T8TU+bd1lf0mVXAodg2QPXC5MrR5pgnddCjn37
0N4GS7Hg4FqZ/mmZVyZfE5+vSSSoQK0HJHn1mjjfJxoft9RhE61F0U8hdgPO2rxB
4tuQn/+1MtSftYWwW33EyjTEf+tL8YDYMZbvQOIqElzYJzdU3dm7nuJF/7VR+XOh
sBiohDiTWwZ3S33ov+Ld0zHLveUGOagm5MUxd26y4dSq9unBi1v80z9ERReOqn4f
AcMuOij/9LqvqSDUa4LwMgFuhpacA6CSFFhcCm72ozqWrScuSXtqH+KKnrIP/L+5
jh16uEi9hh//HHJKrlRgqfGQASRxTni/gn9nmBmxEE48lAwEqS/VhUnIF49IVBu9
CUApqD/XZiEd6duBiw+9Qm0knx3pP9zjwNKGzK6+Hy0UleS9nFHI7Lh6GD2pDIA9
wR60wQI8LTlVmraYXfP8FtqvScDQX5Zf84iBRY/EOVmwlgaJLJ+IYcJ2fQvylXYn
Jf+vrRJyryLF9I6jGJgofxwdykpCZvgb90ehOb9kqPzIAOFsBkVC7QT2hJvcSkP5
D7L8Y2j23S6thHc42VOGWZC61jyhEyIM12XowgJepYARlwDnGkgeenemuzyAbwbT
nVo7iDWTzD5ASDUi0meY5MrU/LgH/ehQvSyoKy6YRJs7KAST+2uCZxi7Y2zuLYsC
NqbA301jbZRmoDc5jgVMMHO0ZSBB9cH7tuwpSOjGXGnqtutzpanQz+WlQPn/Q6KS
c+8PiAQfZYDCiPPdDp3tDJGFxgzcIMFO7nOAgLmQQ8KB5yxBsmBjhuY+8auPIgWn
DixZNfziN9run6gF/xnB0VeJADJ8A2lDLa988ks7JzyCVrIj77uOn/l5M2HTi95y
Zd9Aelsdmmk6blJXDEAh+Ejb6+LujN1V1QnwF/shQk8z926ILuQQR/1IA8DSrAfp
2rfOVh1fQ4JQktlmVbLaMqZVrCGNV8FgC7eoEH1rVCW44S1iRTScCOqPWUp2/B7W
QV/K2McM0s1eugL5FniHEer9YHEX87otoTFcA+64btiraX6kN/OxVZ7wbYb/7tuf
pkzlVpUNOiwuotTF5heSSZrwTO9j6LluJRziJmGiIv7iOGHV9Rzym2106abcXFjt
zXAYSoB11lUX39SIVgsl+3WCj2bVQcAVKlJM2bko0vosjmfiLFeeylh4sSi8g5hA
WcCHjbv0QER6IdTas4vYzIgG2fv51IzXGjrkpTlP0xshbpiGSkV8yZovoqhk8Wd1
s04Y1rNR7EyP7zZANQ6ExTA8q9zoQ9uAd0jGfD8DdkefymPFTjNxFcixF7eVo9G4
57TTQ4QWr2U8KetWJo9qVNoPnT9zhQbNPu1advZcWwkaFd4Bozsbp4zkgj1mNVJN
l9f4L455YnwG235hNus9OTJO26T/Im2N1iMW1hTe9iw0/q5b3SMmeiDc2WlUuMjc
TUUHdJR3gjzwDWIi0UcL5i4e8K8RfZPPB3f90q4JXQXnA3MpjErP3Sdos3l2v0pk
5aBp9YO9rxzWwXL0nHii7LLKPv3SxUNqJP0yQGfLQmgVXwnLbcSG0UEPGdTsj2Zx
QR9+zyjF51ReQWF3VxRUlosfxMrx5UVq91mUF64SiKn+ZW6sjcklM3DLyZj7yEff
Vc3pNvYrcXGTvD1XDur80sJFc6VJAWvvAndyIsaQv5x6VP5HrC2md+HdJVELG5mC
Knpqk3jWT2wX5T73koAW+q05Ltuq6TBng6k/vlPMbYN99CV0cCBVfgVJD2jz9ITU
/1EbUj+9B2wI3Wg4vKw0RPO0x882hB/Js0XJtDOh9PH04YM3DDANuirsCLvi39d2
Xz16kIBq7xdtNLuVkDz3yrtFPpBH8b3GFLEwgXX1q61VunxRL8pP0IBi8vzIagab
UBlcNj2MnwEqukt5EMo5kWhH3aBSdCPniDtmk8fOP9+TdZs7I9k0ua439z3f84uN
gKuPW4fAKONoReMKfve7p9zmevW6DXQMkrVp/GXhdhwQKUQNZpmGzTZSdPgFGw2B
Pak/hjOjgQa4JVGM1vNWikI6hFL2pbPe6U49O1AZkExAPXc7ypRf/c6CcaV2exvP
aFefK21QD289UnQv9nYaRujOyHBIe0m9u/1t8a+zLz0ZdBZZzcJlfDz26/CtghR8
fb5/prKhACc5Qbg7B4Kq3TZH42epc5XbSnrg2pD1JtCYWMnIXr+uMqVCWTeACHdm
wcfO+mZ33EiG2bc97hx5v66eKk3x57gWkg/hPqSJSgEpo75rcx628Tl9eP5JqHnd
e4UDEOOsirQU4e9bANfU9SyhZfa53/xTUm+ZMn7aPv7dw2BZcz2ADtW54rb1YP/N
Ai8dIQvTqcOpYqD6OVL8rt+uNQlKRWM130k1C07mXmkYRR85l4QlfXoDjbE6LedQ
LSIfyT/TtXxaZmjFjvBKBGSypdDGOAqyUeKROI7Q70xQhBAg9JVFSNfpTtv6DYQg
nSXRrbkLcF29d88YssPXZSkiFIh14S0o+rKG4dltraPgBSbFaejMFuR+IYDNmPof
MRlIwbXs3huyxh8Ky8s9QcTvWpGL4UxDqPsHGvaGc6kklVwrQKUeKoLJ/mjIWoXm
awkV7vpI+rOJBdoGCPXK+QU0Ki288qrlxyPpVuhc9oqSV7ptSzFrPMrzs7zKz0WI
ntMqSgk8GPYR2siyxUfVFbJpM4TJObA+EMfqg7yY5aSK0R1aYA19LeqHkJuEHuu3
gFzbWGfEpFbQCRBMOc0aIk70DvMY8ZOv80LnFa0zqlZxL52l9FQq3W6lSUHUquAN
rErEdHRVEFh7O8E0WYM1oYU3U74oj3EzIKQcVpOvK52dbh9r2xMCpoU8eRQtYu4W
Oj8uWKZV6vb1563WLA4oSaiEt4gzKoKeA4Le8U99HvSx7CBhvK7PzoA7qc/2svgu
/UI7tT2W3H6Ly0If1ziceY560RweES5477r61mxSp0adgbFhr+/P1nHPr6sUeg1b
hT3zPA6KIFaHKBj/k6B9iERS3KBFEnOjp/nJHr4T4XPetkpCzLMhWPOKetb/0cml
o3jBvebPjbfzhYC8cShOhPY0KLToN9cP+RRSxCwritWU/qh3mpWeHYHRh8JfCMli
1AcT2vdI0Wu/59ijjrj0RzeSPpoLKeW2A85ebvkzdt7qhhG6amxw/2TZwlXCtaS0
avMg07tCE8kzn+nOsLFhN/x3UOaLFt7oQuyQKfqg3yP7H77Y0XukZIfa8dvEF2Zh
6VsZ6AuERVbUBZi6W7zLshejM0yLAjHPYeB2zYh8CH0V1c7MQwHjB3qgYRYmcwjm
K8KYz9bY8t4wrucN0jn0L29AA5uAnnQpT2vvY52xH6AjCtHOYTCbTRdfC6s5hk+v
5n6RogG/ZXit/QXddeWkWK7mGiHxwhyYs4bJly5u1Bx74bX4llVm6gLaFqsqE0sg
m1j1wou4tUOtGZXMYWbaKCOBcxMTyvrhS80P7WAeGMFaxsu/Nk2lUg/7lIXy8lYx
TOYjMFdCKwEm5nah35m3shNE3N/MERLwKpVlpk767Huzmo0P92GlsVHX3CKneiE/
cHgMN/388WICHOokbvAAUwmsbsigXXc7JWSRGnjvETn9+MIUIfkjNcGlEKKZqF4z
vRPPvIyRDuImTWf8kVhrCjYF37s1MFwWojF9OGklSmxXzvEOmdck6DhaD4WnJF8L
D9+glhH8G7a86yBAchW5eEgRAl3UMorkXSabDjNLj/gW9qB2xchPLQ5bGCZ1JcwW
LKR7pxQxVhon8ObQhjC1YejyDKe6RI57wVVL+9IxpSw1eMCIYEMJ/ZZ6GWE3GrYG
/+ix1uwsZEErRws8KTj8IIz3l7sH3ewRYiPZkqnPtYB+KjC4OiPF+yZRdNR9sacJ
Kl2MGlzAv63pEB6fGh91CsX3HTMrsLdgEZyfnOKOyC3euHd/Ee6w1di2LmrspLI3
mYoQTBKmiyDmEp3lS/T4lptohWVq/em62K4eNu9fe5ToPRmXUHE4SiWDCeGcSq4L
hA8KdkDGBoC+K5OQJ6hON0dEASRy830x7PUL2X3oBgz74UhzKjzwjpefbW87TWiq
3F52N/b2088eQW6YT/9xhoWaXzWYGYnY1kNlUaiK0tyn2fSsN62PaPNgZJKvS+Me
YAaZHMEwBigV3VvSzuUgk2INhqloW5d+D2yDZgiclCI7uTqPFlTiQ8H6L/DqTBAG
UV5vY/Rvuayle2uAVs+0DwlwlhfU/xwiSo2DtLU1SySfwDznWHKQ+zcTQHFYnLUA
c4H2lk9skETVWX+ICZK2bbACo+WU1rxqj0XJn4kZvsH1dEeD14NNgTsXZUp46go1
xkSHWzpdUfQfdJG8QlklihJ5b5kroyV4wRQ+6c8XG6HBTsFOJipo65d74/YRpTOA
PC3AURiluB9mQyFsYpya651YO/7tGsMJGRUiShvqaXpD30pokssMDZtIO6irBD9+
SXn1JSoHm7HvYuqh/N1M4fOYfpZwst2YOw2wer0mcGZgdp6mFtPuzv6YKb8Wmw/N
pwm4+umbvJHotzvZXq1mkbRvvR77hqC35ApjU6hZ9rx67NbwgOBFh/2YIrYYNMMW
CB87LitXo57EW+ntAQsHIeJJwMQ1rvMgW1Fy/zuy9Io2toBn6NMn4TBAnSvH0fg8
F9vJTbsdzjIzQBibK9lzHwwh3iYP8m6EFNMoC2f7lMyB7wimtlgP1A8ET3Li96fY
FdVI/czoxp5AzZjMOpsFuKh3SCAbu9F3ormCvgd/dYbVWG0oPVpAIokwGmzu4Rxy
FpjFQHPvwOp6U2GNakZwC6z/n5YzlVIQrqVKLTeZrL1BN+gpoqFv9qtFEVYcEvKa
E2EXMhkyk/46dQ7WW8JDea1DGyxpy9qEQaRH38+vhdjJZUNy6yi4jXpA4ou4jxAu
nhPHlw2IrC7OhV4/zSUoqZmZcaZsokCaXEbgcvGFk/sUmWvUsVhFYqJRfQhPgYcj
eHqljCJBw3IZMJxT3JLtuV+W6gcir1ViwyI4sgBj1O9VHUV4XXu8DeiDymATSPgY
7B7pDrMjaXS7FoRVKD+Z5dL3dge6acBWXYDkFqJOHEEdC5GsOgbsiappUCmrx8lO
Uvz26kn0urKC4GUwFzgv5RX+ep2JuCnYECQlAzDmjMdK4TiOMlh1eIB8Pki8ajnh
P8hJ1VL9pUbrEE2D8RFQyX33ZxikiAoiGETGcGDvSMwFvTgMV6ZVNiY7l4cCrEui
v5EXEmWjMHXiCV01CqbzYJOgkX8Zpkt1Ld5Dm2mdBEkbLK1eObqLdW4rx2Qk0Gsc
nFNk00MN/ex8sOs+4wn/T0meZXz9oTwCanBTvhDr0rvE92e4KVpGO8jq28n0HO4F
f3Bd8Jcgkorim4YZN/s3azCZJQZs7IY5i/BzLKViuonaYk2SyEAYdVso/LgvsWA4
CSX+BEu1Er4IVzCfcQiZbD/79e5LqegWYsRAPNrY4csx/cYQR9hts7XRDLGku/1R
E0B4e9QipzFaAdZmyCZY7XYv8NDkjKT+ED9AaCRusurgEYG0buI24YAsDZBhYg4k
qA4QM2qQpxoP/V66j6fk/uuq9XgRgzdR6y7rMWlZr6AlK8cI0O+kW10myLmf8qYU
PjJkwqWyNH8/z5zfhKnCZLb+zu/PD4UbwM16q49YY/2VlU0KG63rPP9iCJ+Rtq9Z
xgssi0zqgtgf1YxdRS2RkO+gr9LyDiN1cIt7ZK2zrJTLoHyNx/ZyTMRqpADasu6h
YiaeU2A32DvioeN6cMLIAN9DOtSnrzqYmLNsiwk8+pdH9GzHClZ6j/C+PoHaJ9E5
d1/lhwgmziZIFmLBYIt8XRSXOVkM8VwNcElhmUKHePUrzF2xvGy+Vvge6vQHZiEv
Z62DmHlMpVDPhLtVYcMFNVbt1b61pHr2VcZE4F8TqpCObVu1TUDHVYURS+XIDpd9
2zEqrICYGk98m3zZ/6N+7nyHvVAHg+09dh5h1gsZnyUuvVBsdhJKE7izSGu2rln3
/l+ylrHh2oqbRY9E5/gdBRUYVQoxGFewBiyB5a0mnz16vgH8Nekzw71jGt6dEHWG
97hlc6Km4aBclD9K+4blImVrd7MSOXHLKoUu0ybCroK7aXHjD7FTS3Y50mSRBOmP
IdSaVWO/aegG/gdEtW7OTDChaEwAP6QbTLljTYLxCKvOKm7+xgkdcWmq4A5AVwlU
AV/dtJE297Ak++SUkx8wRZQXfZfX356+ZO4hgQZBKSbmJy0NUVkzE1PdiKgW629M
LccOO2QCyh1Cxce4w8uzxrIXsYxnAiapRY2D/9CZ8qn7hfq+VBcgOImc3U3UN1wy
VhpiKG6Bs5BAXbmQmSKSMIGequSpNxEiTF6aKnYbebNNx589V05nwYENgXsTh+g3
MSmLaV8n1ts9hZfV6gqixzrPMSjdzkK0UTIIKSe6WxYPXg/f9p2MOu1USYjQ51Et
uo2pvYAfKEBxNYX1XMsfesQQxntxmFAHLVgSZadQHY5la9smhjT+92WUknqh7flx
8pbXySJvRvIy0lo16omyU1AJPENvGSWfQOR0TYGg8x5XPQmva564nMqKlOsNVhNw
h/XWmGVY1eiKN+k/CNT8ACmqdeWiOPM0S82cmZKCWXVLPVxTjdVtiv3BV3JD+vtQ
eVitGEF6zHID8kwYa218kvC8SXEyhPIyOhdcLY1sKcf0HgmLzivdB4ZYYvVYWkp6
dH6YNO8AJCTZFyj7WefMg6n8L8yfYbiA7IK4C/pryM6wGPwrzqU+9KNJ4QtCPuFI
6PeWpHzT2cpENWAj3YEVLhEBTovZbXWBCs+zwzpOOCtwfiJnoi7iJUNVsvtoJ2Ko
UBmD9I1oxzOLTytXF5X8suQFvQIKV/UvT1phqZkNwcQzDrYSuC4egE0xvRN3GnHf
QE0u+HTfKum142442WshKmvJC2BEF89py2+R4FrZ94/Xk6qY/zG8To8oGczaVHRG
aYbNkDpQdvgMBmwxeU+Jm/DsBrJ+eQ5lCEBiw7/4TsCw2NWI5sHdwDTe0YVw+CYP
rV3fwTNfSiY5pOIP6/Sx2Bj3nqbIwyhcbruudkVkgQujpSPNdtp30HcdtgTegTGq
dIG5j1gIrNufjgHYsL2+fsStjsd6LeQ3sdWemnoklvyyXbSNsMu1nGqPpVwMWxkN
CDfLNp0ct0h5+kVUGheHqPQFj/XeWFch6FBdWsL8MCHGe9CUqgqe8unCQJZdfRDw
NYKe7G4JWyGv42m6LReQNEy6JX4u/qFZlXMn+Zwgw6d/tGxCLRPXOBQwTgLoXNQE
WsuqOd6fbAb5XI4/uWvFBruuiiUr/aUrAalqbbDs7r2IEnDQGG4VLHBY4YuJMKGp
5htUrTjR5Iv8Rk1BnF7iLsyet0Lw7AE+VUA5+IRVW3rmgn9+Lyvlo8GaqltW635w
OvgEr5X+9/hWm7Tw3VgZ/CWB8gByyaPjd5J8XutPG8hs6vffqWaIdNUAZJiSZx9q
/ddSlhmGiaWGPNtZK9FY2ECQovlXR8/Z5ldg5TDYg0qchE8B+lgl0nUveuJ5erew
/czxJ4WS8Dt3T6xtEjsLm4Qh1dOtjGSetP7wB+La0UCOKGSRceOPG6ALCHzdRG9e
VAr4KYuoJTMt4oEkE5pBokIiH/DMZkD+M1rotHKi66SO91hBWOB5/01T55YvO/01
kdPWDwrHLfoRSGRBLeQplj0Q8WY+9qfQKMbm9gkF7oczVwAc8rO2ADxPQ/VwTx/q
DkyWzN5FngwLz67rL+tMYXMd7R8aEKNQClMAI6WgwxZsKxcj2Grew11nZtgi6fRk
j27ntLrJlkYowfFQMWNMepUHM/sBNsZXPFuGyakr7bt4T8lKuilt0FeNggNjV2ZF
UaAxxGMDVgLT3NeL2BKq1xS7fgVeBpaCSUVE7aMI/3F9yh4ay1ExSf7AFgMIRkQ3
mCGni1ZJhEUUyH28BI3K+H125yALLjyWCY9vchN7yUcpKUnJMkPh+uFiZhQdkUFD
d379JS+2ema4ih3PWSOZpGeFkOyBUm9w8KFOL429J1NMutMH33bbj3UAlxuc9kGb
9v38wuUS6aBWHDIEXX+O0b0CCCS7faEbO6fmd+TGuqcEyYRl+qOwDxuD/HbbGb1Y
dksPblDBfOOfXL+MYk7asCkx4i5fpxY+ojcK02jd3J7UWh3EqvaVd1DMJr1GKCGn
dyHrxv5UlZCCZBaayeVTwXHjF5S6kS0xPEdpMltp6vwX48yTKcvRRgViXcq+drSI
dOx4IMzFgSM4SH6NMRzRcuzo38CwyFcIFnIvFkFwUB/P6s4TqIdg8D9suje+400x
sFMkK9w6MogsWjqAUyh0u7sfFqL11iXErXR9k5GMMcPn9fZxAU/Qlv9bUoVYyD5s
krIZMBKlPtLkxR2aGnahOnzm2+4kJCpB1WnaGD5dy/X399286LZsSS+ZmEQjgFO0
i0k9fol/cUAobSICbX8nCTR+juvQW56f5z6tprSg0ECh7G+g3VHQLkOJ7rgEaOba
HpRCQyRkwlJ9ElSZMp8UGmREkfBDNMsgZ66+6Iqb1bQkUqKjL37gFmEXg32MLhbd
6W6BDdUgVPVbq1liZuGL+CDjuKeD6PdQn4RzAn4r6vdBlQiKT7Gzi338YLfpRxBl
wmtcrhcwWJlYqegtFJoISQdLoKPmq0MAJORXYvBYEIYnDJ95IEUnQZjQNXlOWOs6
3ALTuSnk77/C5Y7IS6gLcWIJxjv5jvPzKrtmzBa5cjQl4gt0x103U/2snYMc8M3o
Uc5q17muMlS702mT8x0YFGe15EH+gNVNeCNCxqRWoShKPrDoViJeUke5kAyrKOa7
eoIMSJBmhRDUZjMdHFBC1sKaJNL744kdAwD4KVX/Guelyb3q2Mb0y/L0ZjlxJoDP
Z0+nE26q4wEPQCtdYHm8Sy+8c9Es3BXEIqSrorTt5540OltDHtLytoYGdbF184yA
tpTWsRCAirWSl5hQhAdhDDRqlmBiEPtlNEo5wKN0n0PbH20Zdwvq4eflDtkgpAqH
/lsKkt6CkE08s3L/ufunC8Xhhq8ZLr1CdGUdUGK39JmWwY7DEKogHMkKvX0qI5l7
+avIE2wNYB48q3E53dCCLTyiyp8lTubb5Wj/fCfrnUxZ8/P6nXOuigRlWbait51M
YorQFY/rxeoZMuquMZmNg3DLwDOU2KO/UrzmfHitwGUnLIb/nHnrs+QVh+FenICJ
iqit9x1Ja2d1LKz7gZRGVucPcTLlCPYLgFgWxVZ5o9g1QzZWmC94s33G13azsdrB
uYetBqGfk4KFktyqfaHnMaif6xVGZhkhCh0eTBWgdZYWOZliPr0Ed3Zt3rv78mVe
aExa8aUVuE4KnsD5jG4JkWPpWi5nXq+05lG7qvYyzKnxMT5nnE8eYkNdRC9wgQMF
ZKLrHlgGhuOcnhPi4hVbJAEykuKs4ZA0e5PAcQlxQV+PjuEVUtLtFgJi7ClORnv1
E7/WfnWuAQdQQrF+aBRWVbGofULXUoxfeKKsIXHthYJQRGxuCSChDAjzNYUUUKY1
msKSL6g2SR8lZ6Wy0FF9lr2gNeyUXcvMOTnV7olnpAmuYOUqoV5YI4k5XsRp4/Us
3eQhJjj0dMk9MXZnRqbjzyXW2Jdu5kGrVfUmm56URYtdrpaPk7zPrjGR44tJSWq6
1LVLiNhnYEgDN2D6cE2xkp7KQKep4PqXvqrfmg45MTSLBVJnTuDYC01NEeHin5Ei
84AOSr6kCKOLCp11s9fGyHFBIMbJuUcxYAjESvioDNkjFSIwBT6szOchGvbLb094
PMP4lb/ysS19u4xs82HEs6WhzlPmO3QNSVu4Zpu8ojI9x1RsVWjEeCodzWhLKjuT
nwPdUHObY6xB2CNWKo8W1SSmGiS6/2njhjfHdcRvl6ZImKMucakEcOKdv6PwscKs
gMDhGz4Cmr5391U9lhXNodzpBDJh9oN+xuGhI0pWxE0Wit/bM1TwWVkUzM0+BF+J
FUuzdw15fHxkmqAXHlPhdzYjuWrVvFiLyQ6SFrXXTuy/BXILWH6Qa+8QEBoVzFmZ
a2Aolhok1DZL2nQBw/GBK2aun2g4gRxqq43Wn/9NqIYWee62+5f+YR+2bSNz4UkQ
a7THM2PApvJ3w9gZ+SKcJkuQBRtl8vnnHjvBRQsL9gOwH+8sLsE5/qZq1llpew1c
IArWQN3VbZX0POi3GbgOtX11F/FF8cFV/swWGFStsdTOE/NiNnE4VngcURvaEsmZ
fzp7ff3CJeaj/P/SDVlXY7vaK02FlzfjflllDPr+YbZHj/QpTwt7f2cScr12E+92
XWPuConelQFKiOT2rD10BzKREfs41j0OKc18//t4kEHRAUz9yYTcq2A9Ix1VvO9B
ZLFitp0gIksY+Mx0Im+6deQYoE6PmUdprcidYOYDd5TMcyCuYAJtQTnWlyh2acuD
rH0701hHZRSXTIjVVl9zSwqP6tAFI/RtMDSA2LS+yNH/AWtImMEfkocjmt9mUlGR
N38fuFqCqjrlHL+U0DAuoSWehNUOT5hibb53wNFkspn6NsYfdmgrYy2H1WxqQV+0
2tuMIn8Ai87p66t0QU/5kT49rfxyRC62A9ub/xBkXrgU2hV+95vS+EtNXRfKAjfc
jZYWyxP43gkZ/5JLwOMuh5tGv0stsxXBJXkmDD8djhiE6vDAcAs65wIQ2aaMOH7e
K4KwSsZiT0yVbmG7B4CiL9F0PlcOFH5YT3hoT/lmVGhDEKh3Oe/UkZAawE76ua4X
hLjuxoPD/13R7ldn7ZaO76o0cAk/cYkQEMol3vT+Bkv4qNxLOpIsg6y0aXv6HLzL
bHU4pnEWpVItm9t641sXI+CfDbY+M5+IjyMXDXWiEfyVHVNLGWl48uHYrjczRQXg
ZVgLnOdWxHmuA4Z2qW5CXcZeQzBzVIHfCSQAyOm5Q7obVqosvX4FHuzswK1emEmC
hRQh/AskyqeHBwS80LP/DEYyBylbicFpbT2EFqWUofrB2dg2q+440KJPFQVvRj1z
4s7utF7Ru7KUWQS7yND0dbfF7MHQDq329jkPfeZ78BNcIMccJabiXYTY1BfTvMWE
LPBiehI7X7qfKT4Zxx3w/DW8Fdy8tMp5Ho0m1qc1nOJkDhdd4bRubgUAziqYoBHw
OAPH2wGhvVkuTFnY5KsH2qVP7gA1YWuTCP2HgNgu/khnB0vl+uJbxmL79XaN67OY
BnzE0wiHVbzrmgG8KNnVdJ/2N09+HRSHwK631ur/+YKt3P49MfdE0Asso2A/q+ye
30udSo96VvIrVDlAi2Sf/fLH//tJSUX+sXMTBDmwBwpfPo/pt4APKR/4/aF2gWVN
0X9bpmUtQPCk7I09p602uphFER6WPbZ+A+9UG1IrRhCaApFkMGsawv2MZxKO3nAp
OM5Q3AKlUGiaCPEfBQefI8f/E+i05wUHcRy6h+ARcLyBfGZotZsJHBzf1io8qGuV
6GCGXWjDeaWOqo1VsQnJTR5oYmkxP+Vq9T2F6kk2xVAwwwba1kFWvxo2xgtlXhxw
iu+GAfrnApA01Gilcq8sBUq0oSbMhwf2QMdNbUYI1R3LbfvBAfsudy+N8L3xwyu3
F7sxR6gwPj6zNMUaL6mP7T9T94myUs9lSfQGkfB3Etg+ZY0U/TqrtqpR1RsuWtmQ
EzwUccCBRQSYVaUjTlf1LcTQp5kCV84v9K+I6SVJvd2yk66lD/CBczgIZ6K4a9QN
ZjcvI8vPNL2wAIBpCOB+eQPKhbZM8oqFS/HyB4a+m4W5Bq/XPNNRQHdHD8XJUOsa
0X3H4ZxXOWreOQG00HqKkCykbibEQgOfqNAU+3VBtlrpHNQkKEC/b7D4b4qRGVf0
2eqA7v8yN2YO6ZL+L9Wp4+6goX4erDutnwObb0YNmZDoVBkY0vl6HRrTq9mNF2n8
mB/YlHTaP9rrSSuAulEDxR9iTYmn7Rko31WrsaWvlL4kmsaDm2f1G+r3wES12Dyu
SH9vPA/YeE2gZVYGdML6r6wnX0PNR1cyM7XRzwek7rlguDK8mk0v+vyxax/CtvGp
jUUAWxavb0NRFczDWwYxnymVZ7PmaHWwbwfm2a6jvbzvBfevS1TI0GLcwJAFKjA2
WAsxpsjJZHu3OtZyII4TBuhwcCiHRJq8nu/lJlyn7hg9Rzs97T+MwJwlv7QsYm+R
WbtVOOV4D2xd84FYNIMcqJnaipW19G4s417u840NO6yR0K8b7xKtXk4MW1v42in+
hlOqlo/wANjkw4jNs8El92axUTbPU8YkttRRhvgMUNaFWC/8P2nAGPvu2x7UBS25
ubCoLSipzg3W69EexYD+LLQTPYuiADuxBAFr2agGHGSWk8prbi5gAh1qVmfl9XQE
UtwqLnpojGZhiwpsyxDcLkIRoUHLt/bpfpAwWKg/v5JCdKtf6jdFkGdXxMn8DW5C
I4B86BqvJeGK5/Z0NdbdDKJmthLnRQb6QiXAz1Dg28pRw1TQQOe3qy9s0x1pqIMA
Sf97DxOx5iR5rV7OSzbbke+UAtSBrdTMr5px2mDHJrnKR0g8CU+hpYe+naYnpkmC
/f2P6zTgZcheaBNIIDLVHxlA+ik78GogQudDjnMWpBXKVKRmIaa8g7Mnj/6uSm+V
i+H4feRsp7U9LMvsKqRwGQyd/HXicGk2vHW0SAS0i9hcaHzzsnv0CV7vvRLAuVoe
zn1z6W29n1/A3Zv0HziGbHHzQpULbcP0OtXt4Pbifuko7wLMn3A0E5EhIVMCU+hp
FKw1tYoV6UH40kfS7bTJgT9aHwa9f/bDELYRkYDFreBEvmjybBYeVofRLSwcOHhw
lrCVFB/jh7f46gg4GI0PQqy6IlG//yfyeOZZztLbEHh76R8JttqtsyvAN3+Xoee4
iUHwUkpXyZaf0p+BU6qgES/NbisqqDdhN1Sxvykg2lda5hucEOe2YVuxWnN65oPC
3P5dP/+upkyQLgGGTb+zzBfuW1MJdwivvbM9cd6u19gv+ufAHsZtwfVKCncw9U8F
Ez4KsNTmSJyLxeVHrT5tUTxymhcGQ4GkAmo+AcMubpge4AfhDHZNQMV+fQpfIEwj
suewoc32m8o9rrwXPb24i0LCs89i/eJs51DEgIoOWHXi9CF+fD3ooe89T0ZsNC+I
fNTviKf/zE4iF+3n2Y1XQE0R2mSMMSXBgtwZEmHfMpzqyt/MkjcpmcEDh7d3uWKT
le64/AzKQPMzIZ4rRWNON+MkAI+CsMW/pV6XuxgOsYnjr5hZNLcsFLU3UnJaFgok
3tVHLa+fXVCY25ultLAKkNDoYKXfjLyxX7G7CFj89UC2g9Pc2pU0tJYO9R+CBGGw
TBzsGTwYhOGapO8isDEE6SsfVNVuMNulGh+zF/Um5xdk6akCm1tELbtHUpLtoEvu
SiId6Ts07DZJ2yWoZvTqpsYp/VcMIKH5+85UqYe48eHFZ8GEMFA5WFBgSyYoqfaR
X5gKNJRou4eI+F1I84ykLBdKFOHrx8hydxj8tnDN945HVdfhjjurn1DCpBODW4Z0
fEKrWImhJnY8rPQ/jibL9VCdZWA79esHEjlSMInMO0/FVZ+Do5Ay1pMtMfopu4RP
L6PtWWW0ia1EvhilRiArjkoapRWxDyI1muzorGuARiXeSuUClDWBJNI4FVx3f/7a
b4zIxkTsBIuLkD5ARmEqlfo5ydkJnvmEyM5ivz/NbcIn/0up7aDYe+po6ZiL1MUC
VWe3W8Gv9/8fSscAgKNO+MwA0RD3caMYR3EzpU+Z5bI5/qcDTuEGm2DJUOCzfdnb
POzbunGyxeQx2ti+0fTnSL222ngFzftvk9B5wwfUnx0zeo6d2YsHC2uiuAEb1/X0
49qdG83l4z97jgfqpQX1zb4S4aYTZC5sGClLasXAtm/lq37AdIqdICYLLtmd91FA
DOZel7bzmp5qLSqeUnktyto0yYVnK4hvuOfJOIef02ILZQOPuaANkJGqkrAVbgAW
xnCeAHbIp5RgWZZCsCYDK8/ZMEzFIv3cYsPqKC1d/w479Agdjf8yrUAxbp6n58Jz
Q4j8wpyNTSgHZJqNuvSzxGOjsUZPnNO9OC34Wlj7CBOhuXj/dx5M+magTg8nIHny
r+T43X1Cntz1ZfCdN1zCKbK6Y67eVt/2+4zK8Gv9kZIsGpTgpT6nYEmTTKjyq4vb
XPpzhsOL7SKHPf1XPZS737i64jPiSbjO/UOu2OPcSujVDE2ky39WWuz0fLD8JdRn
IB8Y6/cxDl3xPrj57NHEXIU6qNvBjIjouuzItefeL+Qs4PSeBWoZJK5RlvW18vEr
19Pp1qvdXK4eNvOC+NWDbVincNg687HlMgR0lhkeQ3H3u+4uPkUHrBFfyDr2GKdS
SRGEFrJdsISqNchnFZrlzvp+jWt8vMz1dR3O7ZjBgFPp5zh/dO5xJc4BFs6jQ21T
jrOsVL5W4qoRz9GQep6kwFavWkY06DgG8J9DO/2b/ekkRdFob34e+XWeGUF1HOTc
Ztnshz1QBP/bNrd6QjcYyN9OiZs4PN6mfQS/AahQdiqqTEsl4Sph+LptNhWytN0U
cxasQxbKxwcORRlBxPHwtGXckMSxdfb8ttOyeLRVnB8TJyLzK2aHg5KEl8MI5TUC
nD3EqrJlzTq6bSCm01nH2TO8rYtOU84AjuUImnIH/Zvf62O7gDHaHAefuNEL9xdo
EJ1k2KSHnvBYRHjDzcwRC2yt4kDe3fzmDim68fgbSgvVZXGu3hfdRRGMQcMpiIEz
fXSjtRQaw8ApRDNdt/LyILzQQ5JK4ZNOiJYYWm6C8lUNYlDWEJtJVTP8OYkgU+ef
ea+GzQKfSoJFlqw1G9wv188kxahjh0sKodoELE15vm7i1wKsAjMrxSKyF//2MY6V
jmudHaNUFz0vEdmUV7ent3ueRCLdbyJOtCvqG+/eZ9lBgIehCCcejzRSfMAF8DIZ
fykXvJVet5Drofjcro6vrz32o4Ol1F0JNuRzYQhBeVNeyTZtUdfTQWXyB2++DKGJ
CHAFLgoBifO/RJlFv9iS2XOERR3ySj/f6xe+pTTnoD3w50rJ0r48HYE2Cod9EzQb
XGtoiqx1n0QCYNCFJHoaEMZwHID0/gKFQtl+HeFFIIe+DpH7/rUaDy+yMHFOONwh
/te6NQLnx2Qetza5thrANcyhhm/0kk0tVYTouJYQ8tMPZtwyXSprk09lVEhfHZhv
5JuIA/8fwDtgAEC1eOZ/UkZATmtyPY9xftIUGAloR+y64Q3bGtYuYzcAiENCXeVK
NunomI5L2HgDP5Dg47gUkawXU7BGkXHOd1RAIsrhYC6WcsivcJsz9iKxK8azpoSd
zyx3JQ0ve5v+5MrNu29kIUBdtP/anpKcgLSvp5xzt1yaxnwQRDEEWuy58kxICvgx
gbnu3luo7wCEGZObaLPxMss9ghXNs2InIxeAJGeE6Wjd1oy+B40pRVG6nJupGvHM
rU6phzpU7k16UTQdaTjgu+52pk9V+nejSQX28ujJUWXuGVAxr98m03wvW5VnlbDd
GhLSX4b36Ia9rshD2I90e7Q+nRujvvoT+u1gtSc7Lhpc73VPzWteTS/9hZmr3NQH
MO9/4uhY0e9mv4bcAKz2993iB3as9iGptL9UiS3dhVYSkIdiLPzMot1kSs8RJ5y0
1E8RMqEBLzQfmYwQ4EVsbR4hOoZ9s0EU8w//DRM+X92X+79lv34WpQ3s1EK86AAk
QpsoVj03CFrayPE4a+pIS50a9vAQVzkOE7R4FBmSQnxRx1DkjBXPfEQp9DhstVt+
hljpP4qavEsNijVHRCxxW2UuRDhdA03621qqcVgi0/dPC58yXNNiA/g8MN3IUJyS
w+1OtJ0J4Bs0ynZy1AyKuTYwvgfwXRO4twgNmyZOlgP+6kQBTw7XEza0GtLZCiwm
us+1iEMJKm3NZuiG7yCWi6UbrE+UolvLSQM+3VExii+tBaTfSmP6pCyRF9sUQvwo
TI7pQ9H5jcAuwRdiWQAjP9x3erImjZ8JeBRnCzy6Mjm7ziaO51qkinQKhDKt/QYt
yYJe8hu1HKj6DjrW4iq+MF4iiHGSSbJAmQpCf26YbHZ2cisX2seXl8hHJjKp6WJ9
quliXuDvpsoXsTdzd/yTlEfwCw7hJEUdpif+CQ3porN/4i4an8nlEn+IQGZUYG7+
CdbTVnoC8cYBSMJtZ9j37Q+lzTFDIC607vT1hRW22/ZMR9WNhE+niLS2mA2J7Rd2
UPIDUH3BBvfCPQT0HUkgXSwvMLF8jP20VMXuE+J62RtWxoJKvIt8MWRxjVxVM3f4
4ZjdB8XBZZLzMEYRhAv7PIMdJuRXoxhlTI0riOTX8NG/BNimYzutIjTMZG7RuJOa
XQz7EYxHnNtefSF8ted7kdZyc1oaxnPOaqYKJKZRSYtfUKU7gFUHC/tP9dMCbOyp
trYfQtYInFaiaNmAaym6Oy6WLaOGa85KbEtncWq4kgpJ39h2nOWebB2Lqey0AMr5
5vSWjm+6CS52eQUbFnPaheBGDqaYtdAStxWisexdTYI2zM2LGYzyMWoaORqHkty4
uTgyvhabpbOT5gq7uOUAkPCJjNGOyz8HpYEjNmeQpA/+q/2hJ+e6CtisfQnn90e4
M+nPAp4t9VKKNSHCWdpuBBv1XS3vGZ/GN7nn19AYcA3EoLXanAnZnzBB3xtsk7B0
YD7tdrQiIhXgBlzrD7UPiOYT+69w7tOIbco1mP+XTsil7i9dDTngJFLiXF7uY+LJ
VNmruTvSwZPipBt+D+eJt1HYTaoryOoxcnUhiEuYOYNSuYI/mREgfJxdaec4flUE
vrCXiGZzUy46ZVECwN6N6bWtDRtge4oXec+6v43Rq5QaK1RsIERTrwU2/3QG2QW4
uVTIrbFmFvxciwuR2w3iRFh19u8na6FKFPxDbraTpNUTCV7zku4C1l/L4a7JXC6G
aQDtCogj1QZ7786gavhvtzsZM0N3P+jlKUR9yZXhiZI1HmkueoCVCVH3QzJeJYbj
8fIZH0TYmX5NcFvHnjWHmFwA5EezNT5ucgdPJPLaWnHc47wfcBjNnx7dfhTgE995
dc3gaQ+k30L1AaS3Wsn6V9kxD0xD7W6fp8zIH0BS4QWc8XM7hPjCODD+zt3A9tFA
qN3moWbWsSrEKzBlSoQt6Y1tcytWA6rhimx4PZ7xU4WHT+oZdDyx7xcpuq4Efqs4
Sr0MedvFhZGDcqvdPqUH7dBl3kCMC5Zs2tk/iIWihN5PO0wYHRrqtBW+tN5iki+k
dcAF6IQsvj+gwXKOhZ+6csLy73ZCzXhtr2rC2Rq5PdeY+y9b1Y+jPS1aqrCXBrS6
1p1KeIMnxDv8MGXImNmbJo71c5//FAxmv8SqvG8j532/n1CVHxgElMLldZtkj9ZU
8r4mVhx+VdKIDL31+iXLPcCntLeRBRgwXOYALeUfKD+to+g6xB8uoeLIecVj6v0Z
cf+4Bu7ch9yVNvtiGDrmgf4R4Ri79kp9seI0V9YArFdcqjY8cuapdLMwUHgwX26L
y4ivqEi+7jAJ01eH0akSuOihn7wmRmbK6ttiCoG2o85pK0tZ9h1ZapO4BhfOBGy9
HiLJwWYkxpgOSPby48jDsdhPdp4rIso8YJ5VGhaB3WPZhlQflWsSESVHeGvrS7Kt
ZHaKh/gl9NWM9GSkZWBAsqjPKA8GKv3x5VSkHEuzbVHZVytJvR3zDDDHsayKL4yZ
Rzt64a9BqnO7P/sQ27zKdOm1z0PhmqO3Td43HjjmN5bjfIoHY73X1/yA5JOZp4LG
680ZBbDcxIWDd5o78hO+Fcpd+0nQ5HDvLj9g0UEHR+MC3jPetkU5dWoB+RGSG8F+
R7WyBXqq0rD1rwykHWX0kKNycGQIlSMfYkc7+z/A6hjnhnwRCr32ZHqhxXu1jVud
ERaavpM1r049V6IKjq+d7wc3gt4RlqgF1lCLnzv76Sjyg2TVqShR4m9fz3hBqUFb
smCdGgGL86qdhF8sH7FzSPzvzklvYbs8hXidDN8602gFiOKKxMLVaXk7I/KCLrp4
dZFeqiiIZkqooAly0CyRABNGCt7gUI3RRgdZNKrsYIveLW1l+A+W/pp48MBM1VtK
qk509q6gJHOTlm5642cV6bXL5sHeqHr7JQEQJI/bGckynlc9lWoRIShTuPn2CpWr
Vu3BsNY4zMypK5YIlSl5SYTUmOfT7IRWF1UtG0Em9zHOGkZGTbEpYo7pZ21gv09O
YlvBFJOfkSP6zkRDux1uU2VBuvkm9ba5CqeUIcvhOOJYJVI/w4EQTVSR7qON1CNg
vza5CgMi0ls33g1mQn70Y82HXKnCGqAzD/eXBeGc4fKCyvrEOuBA2xvTH/fIFTPm
qv43hfRWzNXIE5uBE6Xv+y2IY0TajhMuLdFem3IDRWvKVygh5X9Xgoy3QJ4/m2ZJ
qna8eU1rknQ3sPx3KxrqlOudaQDyS+LHZdxst72Qi/KE26vlTIc8KtepD5D4PSgc
GlhYikLJgM6PDWhAIAYMflpK/TX5NJWJdVmk7znv0U+Pd8HnyUNd6PboaGxw610W
pUmnaQu8VCr72tq7VQQzec02x0uhQutzDdccHoSsA1KZkv0Ml57yyl20vzfgBlzM
khWt9+Ab1ZLesUlXqJTkjl6LGbYesw0VjtfBV1ccfRF4URnYBcDc6QW0c7zDd2Od
TkkcMMOibVw6QOzNQ8rFgB5cskvQb0cG0dHY/Ove6fT7S/W72hBzaOYHebMef7ju
8KMWXUOtzOgzOT9wxQeDKO9TXN8e7VOHlzyiq1scw8yAGIj/sqkWaHVCkIsB37wH
eY42IQzZSZc44Hh1Wsit004cmqUEo/Qbp1+FiaA/YbMnQlVPeb2bmm4htxxB3idk
AUGMk8TvnywlkFqe0xXn9gV108O4dZYqU2ql0SjwcRXcLtZZNBIDecz4dB9Hf4On
i27RgXb85TwdEHJHBgMGEpJEWTUC0Pja76HW92iuZ6ktSS1eyNYmHojE7rW1yqqu
m+gMhD62vViLaIMPbAVtGLNLPg5/N5OTTMb5f3MHXju7qHJGZXX6sIha2VHYj5nS
Gz5AwZBis1E8JOc1Hp+dAJM5RXlf0abgRWsfXK/BVcLg8nJALttsc6mwXffc83Sy
zLxYYQs5wgtp8CRRVIEYcTpG26MR0LxPfOlpAFbiZH86m1PlTi2GkJzSebOW0Yuv
ciGRbNX2JJZ2I3mXpuBPY0YXUmEOTbvshiv39Zo2DfqRzXE6jfmKrRFMZd1HziSe
sRagbux8iiLNRYhnd+wDPy0m/+O9587B18R25D7Qkp+cjyzLi/MuB9EoelC9a1Rt
QJu4n3NJEdflBSQrrbGUbSVSJYtQOa3mjNhrv4VTdQXy3oNjpPbsT2wwMt3JYT9x
bSi60YtPuq3TJhYbREJS6G9kw2Zjd3Z4JUuOOzVz6HKlhjbwd9J5PpPRGJXX7sKE
7F6+7oThdpyPH+hdKEVB6jWHO2+TCOTCfn89ZO4r9ezxO5wEqtJelDgL1kVog5IY
T36oeqPn6aE49xnxBJ2y/I258bP3i3x1nBgg21p+R29agm7HxQWBRgZ4lcdtuMJk
RLGebcVdWTzYf0eei3X7b444FO+ZwhGp2ReZBFZlEap8wtdC8SMt12irVagT6NyG
tqgR22iYwoOPIIMD2yL6Vm6aXvnpC9weV1amMzFDIF7YpqeAbShfzuG7Mzx2SIKe
6aR5iZP8ymbolP6prZ8bIOedTy9UruJaUjTnS9yB0TkOPvMDhLH30eli8e9S/cwi
/raz+/dTarCT40tEi+YIJqFesvsvnjFiKUJV/ZrF26yKl/gKmWBpohyA4Ui5oQV1
g8KtA48iU3UHHHAZTTyAYlg4pFQsT3Oh2e704Ess+D8Ex/GZYFtfgqmqv0mkvO1Z
XWafCTjBgB8tDFiXTjeemPsu71bp0r+RkmoT4QoPVwvy8U0jJCX/ygQQWz0RsY2L
XJurUzG29nMcDdOf6h4SIQVZY9kO0A+D+g/kVm6DhSEpsp2gczY3Hke53IS5TZIM
CGLdVuqbKhhO1MGlunqLyf80t9c9JBl82OPKh7s2Lr0OojXd3vOJVUYqC87qmmnj
Kq56CSuPeB/IriA9CQKvFyF9Ij5qcu2ErKIHfVYZFiQtATppHkHSz35NZZ7W7zjE
lPdbTthptBXkof8rJ4OWkvFNGies72MdKr6HTGVaF+5+2oUynvy8RP5lGTkwIMtr
DMPopaiMON4O10oK/xrdCaoXm+iRhS8X5xEjJ5K/EAWXJzPFXcee0ervxFfZz5Of
9lw6csOXIRJUUviZwvTZtDCLVa6wLEmTIpeJyTU1FqB5fqUbUQPRfZhEg+ufI64w
j/QJmpg/BeW3vXqM2QZrbc8gU5J8A7+JZuZlxSWEPZ4YBgZcZuE0wEIB9K1su02x
C13D/6RpG/6AsSHVbFdYQYbKyJa4TAkl00PN3rFSB01OLBJbEpQXDlauMJiQSS5u
7LN1JUksuIdxp+6zBqsnlxvEUDJm69DvsT38ODY1DQR+oXCD4UZ3cU3IlESzz86q
2Vrfd4tMUNdNn0NGeIGxKux5YaXnVj3m5g9+ELXQ8vJW6ZstF49KUIOlHgxXaPfk
uayHhMs0ShaQZNsfDkqWnwaVygiyWBxnez4C9kT9jsEmVxM/251VXX0AJvPDcOAP
Tjq1pVaN6xG4u3wZJZWnVvHWwv0LmwBCLt+CizaAx4iOQwbtIRJfnhRkrzsHqCsW
xyij6xoR3USofn3fI26uxwDync95+sjELA3FnRCHAO1M/ZMoFjcRGhmmaeAnJmoh
fn0C5E+uRorol9MQMLAOYZcNsk2T8rWGLqr9jmxsS6sAbj+PPzfb5DxDIQ6glwMa
dSuf5QOjmO81nsyiyIl5HNh3PUopRxIHA2DR6pMOrCCSwowSpd/uyyOnKGwqOnA8
n0F26faqHJjWGj+XGaY6FNFtslVBkjgHlxj8dY2wLpO0DQyWK+5mhVJK2AN4f80+
eNHirIEbhzgRbFt1/K0ufqSxLtrhvHZXjHw5rUevYZx17apZ72TrIXnPlcDGfDkU
NGyc+gNziK6q7Y3SNofUvYVCfMDCX/3gkRgw9tUVpGylf+QSj34db1tIHSD9QayE
BaEVViPTauNlNW/OLTTo5n/tBKoX3OCvHSWQZ4QsyDOsIuOZvNbVUht9hWk3asTe
9juIBigqy58kvdomhoOhzbpn34Wa9pDgvB2R6QoaMQdprTqioMpzFu8Fe5pZPcvb
bPv9LWhGk6aP130LwQETAYXywiEbYktAWUDx2XFA5wNm0gVZvCFmX2DMMxoGESTd
xqJBqyMvuL0N2K2D/U7++Z59oGUbpYr4sKRI9CqUKa2bhBfFLCr6vJHbvbIdnby2
6pcjaruJneESrwoRpi+h5Bf1wXpYxUCoPghZFnsMRTqq/Gvo7ItGYLZLBJm9hX7G
CvEpC5NxBBXwRY8su9I+Sjn0zplm44SoCYXxd01kSGkkOoh7L/UhbZPQEE3QNMWc
AD4L3bYXDCa1Ni1h0zOfKtJyUnf2mG+YqRCOoq2aab/G/1nBN183WiOHT6i29KzL
7J2Xv04+9GO5YTPm4IQXbJONUSaKnl9qHEZ497NSVtpgPqX1pXcRqKy6R4JDKgsB
JgA53Ode0F4ekoOKHV2lTvfTtnOoD8WnokkeKukX3KXhlW5PnQDKXEO0XS0LH6l2
oN06U+uwueL1hjynMrXu66gTc9iF4O+oeLHqtUpIj7OhaCzEiYKKMKUcWtF4SOrY
Dw4gyx+fz84N5x4ZCYu4nEzGqDJJRDp2ZRBTSBe6QjZ+qcfYSrAwuOYjcGjDp0J0
HDuxmzpwBhltwj/OQfKav8NdY0r2tKAeExE/w+GDVhemOlCWNeACYU/T99h/jcqr
rHZue3x2MpT8AGtUwQ/IXCjtoLfVXvxhVmDgdnp1YUMmHw7Jasm9tTaGYz8ptKrO
dIpMjflUWpldZH9rYQ72juDnBf39xtHdE/6pDObK/zRd4WS6p7PZsqflBFtlrQe2
owh91ZvoC4CoMyTKQm0kHc1HVEWYMpft+ByuGl/Yy9xCLv0SONys1IAVqP/6XiB3
D9fUr5uY88ZCrcIsoklMNKx74lruGz/TNQPro6RMT96hKUwiKpDBPoBez0aeeRqb
0PeFZGtGU9c8FrSL62GFyRmEfgMAO82KgXSZnBEn+odeHN4zjP3M7OIB90KkYViM
kH5vva4qgo0cCIO9nBuKq8pT5z+TnPGmnp7E718WRLuMqqPO2+g0cgA5mzE5l8Ip
+4R2wPbuP0msoG6PqQkpxDYveJ3UH9g5N36fiDe2uZSUJgcKimSixVS+yPxNCvfM
NUMpVBSR5fFZ7DhtDZoKtlk5sPJV4tuKZN8hnKw42LBIkkSy9H+0p/mGVi2D1qDA
dbRI3O+pP+yqUJVGO9VlbL/0y/Ojx5ra+QoJMtdqP0eoVpP/ty3TEje8Jdtpndp3
K5yJpDH2worcEl9P2t1LkZk4cW+7qLrnVaLfW6ZC4mI1lzXCGfwd6dPju1D5pcXq
qZEBzkZ6wkJCw9gssbRboEMVGPyKCdcmZg32ydVs11MpHSDY6HiftbjVonBoBiLd
a+HoW/qfT0wBsiAA8f4BlN4yBtSV46wy7jvVlZ6y5K3xIhZWLIaouzlGIXTmbFBg
D83aBMdRDNga0kULknicHmRrhrhDQey0TR9r7P4ztPUIFkreLBo+Xny2R/46qMiZ
L1A4EHflwyI483mVMxVZQN6k+yAbmtwl/FGWbHn+DiYel106CIGvm3xCSMCQObhg
hVJT/Wf1B4ybcr9DDs7k9ZmehJVfgfXj1kXsknibEDLXa8Ta6RiE2eL8cxf0YQQq
xRJ3L/dv6/UX93bKUyuaZkFplv34F4Q+p9Ly9k4yLOjw8Pn3fBrC3uAk+9FzwcXa
P6RuaY2xfeeX/FoeyWmapgD86rQxVm7xNiWxvwEPpL9HRfFGRDHM2Mongz7scLUG
CnGLpfDXg120n2Vz6VNVxcYx4zItNWgTzGFxyVR8AWpG9WOfru0e6LCeJ6uCxKbO
c3xw0j9IBif8fHCySozxTL9xel+gm+MWouDlxUox3VUHbPrL/r9w2Vgi1MHzR+Jz
Lqk2BS6xHUnVGMa8SZWUuO9XxDEQguMwWCqxrSBKzWTK/KS+KyJhUM8qlF+FPMf1
VwTujDijCTg0wrBnN1rIofid4rvGa8fACmgOsxn+XjSts/xVRhUEa1g5ZsZKGOzi
r3so8DyxeSVfs7mhFcuXCm/+svRVlZbI8VO1SzE9DvPhO8TmAkTjR+NwylAgRg2b
XXRnBhpE+pM35I3qVd0ElaHQBkWX1VajdvsHmhSe3JQ5DdgdGDACDyjq5JCBJhIV
8v46a2/yZWLdVqWkAciK5hRtFQVKsofmJCufne5LHQ6/Nwi1ZGlQgI5Ae1KEXe5l
DlSaxQE2Ik75X3x0ZfHVCq5wgWCM+jOJ7HnSkDaxnczsFezkGkBA69dczjzbU7ju
Mll7pxEExs3wgkZSPCftaSIUpQ3RvdkgcnnZJ5R/+k87oac2oAW4P0Go4P73KaVA
iGgLhOzdXbpoOaZOvCaqvNTQR2qyNOKuSct8Pm+BPwnTUNi384ZRtEvPm1UNv2DJ
RKztpG2G57UMhjwPQ1L8MQ75lXyZKSYVG0BoVkCHb8Q6g4G8WM0om6b47RoDoPpb
GJB6AYijjTu3+oUVCKmbHSM6EbEZuYFEVpimd7GQbKecqZD38/hn+JN2T/Ce244L
6rO0mGhZdupGd1lpsW+ubXiJEsoBIl+32GCpgXyFHqcuQIp/5PWoJrHki7bAifkf
35H0hW0mXKF1jTm1I2WYyhuFza4awgYjikDWQ68stf8IeQMPPhJ4IZgncJWwDrJO
nxfcxo60gwbo6EE+TvyedANF3E3d6GBR0qmpcBi+gprLZX7uaetYaNdxrow4l+mG
K4KGCQZCu2i7XvtJEjGtR0OMJ0EmNlED2Mdel3ojkbLZGMgTPUQROuOfkoE3HbUj
WRRPWtxH26eKRAaSF6paVgdRmJaMGYsSlDp7f5m8YmCMPpScWu94mRz939DVx1Ob
kt00qg/TD/S3s4cP4Jdyl9y3rQetSO9mGKi1cQZ6pMXH7o28ZF761U0LCcsNqduO
9z5hZXYhjcewQssuPJgKbPe2ODGVqqEPnBn1m8tvpRJId7vmVdH9fI+r1ZWWfXAL
mTvrUguoG4clPyhkg79dFuT6122raU6xoIswD/SeVxFFd9IepUUkZ7lY7Jh/8IBo
3w2JYMhicJ4WMiYQiv7n0sehsU05C1HEqMc30xoZStiU5emYKNx9bXjyKwdIUJPI
tZIsLZ5W2tqihAfjLxUwyqFhjD9mzhz6Yayey8KTO2Fb00hGUYMYo4uX8r2xleHf
L8+hVSJvCxQJs23zJr96glB4bAlBfPoFaN5y65gBKo5RPo68khNeVPz33qrFUkDi
9HInaQsbdSqIEQhl+rrReWW1bV/iz4q66VVviE6LkOgJi3EucuTlk0G3ZtIijFDr
PtgWCM2HQKzkJ5P4+Eyw1Lf8Cwj8lf1AjtgQKf7oHa20pINS/Icvl3ZgALUt0VXV
MAS7rCq4CrtLhQyeoHr1Vz+tlV10vp27yRdeZHI3E0LqeSU2L3cV8hmyrQFxwD1y
6n9tXQdusppQ3eH/6nG3O3qH7FplIX+ovbNi0fRc/+odrpvv7t9+c2tRb8JE0zmS
VBCRSyDxz2rAkwroJd9sOrnw5oPVLqFdNCpvrto0P/mMjqIjrqsLZoFB/BcK33x/
DEVebglCYqJHf7QKAM71Sz2PbMYKsbQ5vlbYXFeX1x/8DC7UleTLcGrj15vqtAdc
k0tz0pzajY42zV2cRcrqwm/z/ST2SDyF0aP3aX0198WwcB8EE6OhIR9fmNGNkae+
VwpCEOE/bBZkHjNxFfhvasU28UAuluXaBAR7AUArCxWVH2ByW+dHH1/QKCA7+1Lh
FZpaLBeUimolBqv9A02qPtNHRPnrbAkZhXkGAC03+xV4lC5Jr18m6pSMHbJgQa1H
uaEoFrvhLJXTzLmqLRQXQbqlKU5tO6xkkB1038mosMOl5XgAjWyk8ee5AYBfm7Jl
BkIdDt2elXKpZT6+QQLlqP3CBZivHE1k7jryL6mGh5hCqk88kHvBz+M3QcSHaPLt
vbB4QsuR+iPsvtOZrWV/I/qtgYpTyO+xy+yiuv7/Uo2gl8bDbKbQMFDEe+CJRXoA
i0jL8tGMk4Ka8NGV1uAKUQrZjWIYAPvzgwvotWRhg6voFKgbLMhPGyVQiosfv9Rm
NIe/cg8r+gJUhGlu/TtGaDIM3vdAqIkYwapVlGwTPzfmUqPO1WOfWyckXwUDJ6XO
uNJPiF7SzCSqI/hH2l9ySvDb+xEufcFmHbOna/tufD2QmkPp5wak0EGexDyeLCpw
E7puxF+SMudP85wK6ONp0fhAXkCoOVoSqlyJaw33JQhAQKOPApWxzBGNSQod9d3N
DtEfzDHh40Mg/0EjBxvXghuwH1xSeWqSronUIQZxi2q37wjRrgHkY2Ictnbi+iAI
GQiIa/pHfrz7fTbHgx6BCqB5hPMBlQfXSwgAZuzd0NHB8faO7dSxuaAPa+GLGtW+
odCz853O7Sy3w3WrLZERS5Aeuca9zt38Q/d9ZqUXtY+5j01KK4vQu+cM+cKhkJ4D
Vk92VT8jIq0f7lH385qmfmscUoIXBlkpsgQcECj8qFZu5nVEGPnSlHIWcNoQ/cqy
gGrLPqlFDRJm0jwr7g1x1wW6N6fc3FhOLsD5tbT/IUaGrWjpi3mr38FbfVQJhgTp
RdXdioMR32BOCbPeoFkYGO4mHf5M3oggrw/Q4tyh/r6cYBpkfKRvucuPX5aLELHP
Fts1NVGB87S2T+VXgZBJYDhXY0859Zh6QIy3jIVBMXs+NX9dvkWAwZWJMmE3X7Pn
UHIXqSXGGjJoAGTTRc2SbNO4yFKPzoOTVsjFN9HUQ15YWZTS1gSNDgtAd/pIfryO
+FBlAg+XGcxZuDwpUB54uq7s7PNEuSeIfL6rXc1zTGjuMcqrunwoj3QBfDBaX4Uq
+rqibLV6oczlylTXUZLOOSGimbSs9hImU7neK1JbVLDqa215x7AmFFeJ8pHU6pqn
YGnQbsH4Z3gxHmOLcws6Zh1LdfkDtgosvBlgm2dBpK6IXd8LJtZXEPMaojmNgVsr
Kpj+XpmUFbPsNqpNkJWHKdYHRp5KCyVbyWgfSdwRPPs5gfktPe+BKxss0w5NDjX7
tL2V5o1b0K9ee4ipwbLzhHtgfrabtuDxoTLFfmZ5KY56f0GjVt/tICdx9JOaOa0d
AMZoGJcYzc8AGsWESJIJxrHK8VBLgqcCcaT+1PszjjR3olA4DVJeRm+9DQ1E5ndr
cfR6MiRF94vT4WbqgCFbA6HMFcutBrNQVZVMkvawS51w22r2YHhP0j6WkfpdvXVs
gXeqqHWmHUkTdW2EU4ircgOkFYqyYSVQnWwir2ZRob8MluZpqt2Hlz+vQP7/b1UU
g/FQ8/3CQmKHr5za+jNPsyYtgiVUaJbLa0wwv0WGNWt36Zb+p7Jijfhg1CKEhfpC
zQR7Qthfe5pM1WcfRZQT9XF8Zz3QAoh/dWScq7wfCgci+39ODJk5VNK1VXgfE7Yy
HxOkrUB95Tmo2J1Z1eOcG5MFPnA8J7luFFqG8ZK4UnY+uRU0AblMTEUON0AWuCvP
Czwvx+bR9TxeGvjmuufx0ScdBriALPe80G+eIG8IZflZEPMeWdmRgkxCvXa4mV9+
wcj6WCrIpytXRBhY/Zb3nGuxgB5E+s5JT5dh8136Gq/5lYdi7JimMfQQapkuz4wM
CVyIGvqeoVQ+1Xpc9P6J8LtQ2XwrBsx7qxLAhp7URzd9qLFdmmlHZs+KS4CJdPOb
hgaBUJc4DqtAQmgsXv6kDDnZ/d+lCTzlDKREvI5VnD19PTKjOSnjfPSMikkW5C5H
rhouoAJup74FtcxEBijshki9rsSsJjib8FrGDxsI3eyv/TAJr0lUMuTKKLiHnY/I
RWmrq7tek3txmytEwKH2XmRqkqdVBA+Ah8l9VaC+dNOuqdTvvHMGxAOlMb+i8/r5
weKcdgnbG8gTwLUi7KyXjdi/wGP/AyUbH3IM6qeLiq0tk8KRcTGNnkmB3Ag9kt+7
k3XSdGRcrztstKTmmUcZOHLOz3mftv3mr6mkiMWzc/hX2F48by984GbxNRcqSuvy
RPpTMYhMQZ2spiw+2Ho9m1tdyx7DZZ5ECxzGNDM13K4b4WbbLcyRFwV7eV2aThPx
x6muHrQPHJPSJkgzoZGSSR0VNIJ5FWFn5a4I18FlE743AB5cPg8f4+H6nbKNTrSg
vpai/67oA0KBi3x0x48WNdwfJoM+p7mZm1optLa55RJeNbr6W0QxpfdvoXiWjG4G
n0i+NbtffcGFBpFWX63xIPC8MdQQiRsmI3ff+G8Ez8GErlvqp547VpPmu6Y9WbIn
x2NZ5egaS6xLoQ5kzoWP68VdXJ4wybgLgFw6wz2gX5ac8mT/d4Pt/NfiM+RMLw1o
ywsAAvpMXX6SvuFITLnNJRgW46jv0LGBI51ewXWgk59imlTiNLE5GCIFupxYJpM5
VVjyY36NAbYmDUt++bxgsZfmr1vfFsK3lwrG+H3+BbBn9mBYGpCjOvoNeLB6wKbM
K5Q58Onr3WiH9KNGKkvWTSM7pgjs489Zm3pVoSMWOC1dMqehXcXcnJxVonB1zLQK
wjBMNpzIqfKU1UfI9JoH2EVfBKPXJ0YGSxDT6Bq6Sd+eeOB3Myx5HhcHRtMuWi/o
q/9ZVfgOlI0MBQbOUKjmFcXhZeX0By26Wm37LL41+CdIVEG3q4wK5nnTWaTYLHeF
7b0fclJG/f7yg7d1bp6vieq6SFiXaUqT70woqmTfW7f/b7RonLCPUsqCuxoeIT9k
Tcw8mDDorlLPgU8WtQzOFBqNuxUmEYnrF24l2ULLUKKATp1I7VY8yLWvfzIt4y/M
lEjoJEYAWvG5hj8i1p/Un8kiCzbM0FgN43HaH0YGfbbO5VbQDV7fiDF9k8GJ5od2
TiT5j0hlZVsVvGoF7TqPF2na4vBXu7YSBEwcOGLYuTohnXgGgMbDMWQFKJS3DBGQ
3KJGnzdVopzyp9s857eUEq0Krmsgtr8wu9pgcko73EEFc65p9IuFXJh8FaRiA+JE
7qG3RqcQfEI4IFjZm898OHV/9oaZOfaHq2Sk+2zieq3rLEbDjYsWVLCp1i4t09hs
6cYXtoODE6quC5yd3uxjEu6nwZG5LHSc3AzYH4vFuBTxagTpHsOxaFEm13JxBywT
a60aJiEKVZ7joXngj24uAOnscG1pF/7dZedOe33fBKJP1I1pCdnRe3AmUe8sSCAy
5bYllRDyD3b2D3nE08E19uLRNnOovvhad6I503Z71KO4Z42KJcyXQydPG/E5525Y
sjM6pM5f6GfLhV/Z/BbebU2X1KtsQ4n8dtuAtGRv77KWUdJtXL5jPjiiWfAFhFsm
MdJBkqOtgOf3vFL7LWQB/5+UsF8ADZdPzwNOEfGWo/TfAlbIpmHf1zy8IEP85xMB
Ga4mfJ6gJjmagRHVgW4uU3cA194R2qcRFnJwYOmGWqwkbB0wJop3Wk3nPhD4/QBl
t7mK7IqD+tekN7wcJK1apk4FjzefkWUBZR1m0YoHUOgjbd6makt39g5owTPHqqC0
VNygWE35QndzWecoMT86qOGzgh4bk0JdQC+ApihesnhPjWql2OyPDAQKmpbaEUTV
C9U9Dz/hAp3K+Rhe61cEEwl5ikoHjuEy45Ym0tRZq7KDBOTUygVyIY43mMXUl2oh
Izdw3qDeWkfWcp0Xvw+DGAMxHP60SSuniCjGXsXulml+negIxTq+/4sVy13ZbLhU
hpD/CeiBp5D7pgiG9kOHziNRDdpto2XnlK1AT2be2OgYGwoms9M3+1SXfBw9EqV4
AsM2g8FrBbO/QKJQFMc0muZc/mlV4mWC59ODGbq6GUlirvUpaetoRT6vbI692L6v
17NjBEmHHeh0w8rH9FvdOXeR8jv1LcbvD7TPtwYyDbvfctpfXZbt9tvfsF/uBIFv
SxrAE7MphZNt8TUlSgT4k/Rq7fvzChAF6arggyvSXBpcDp5Bcgfb9JHLbQJWn/+p
QZBwhE2krLOnSQnibVSRGsQpt1SxHPY5UXPG/I26HK6ny7fsMy2G/I2DYS7xv3hq
9Hf/YJ5uy1frF4GrnU2RALampwBlmTWtVrZNdIyGradpTiZonCGuH9k6AAbJAe9z
f4bhEBfSspVUG2lPqKhWG9iydyymu1vJ13prsi3s/vEaRDpamb61nQLLX+XusvQL
Gckk1GDZFXvruNlxzcyZAhFgg3GE1nC5eu0XeNiEHi7j7YfNuqmK9Gy9t3G968DR
pHawHFhp6werSeGJLgb1m8K5KF5ZOvLI7gMSqFVCfybsu/TjoeQMKpuzI5dNUcmx
qyOrKqr9QcnB9s9rXa2NIimLiYmN1NCGHtC8nGmdh4l2gBKIpt5DeETUFgYnkFy3
bTcJSj6vJ8H15IR3fuatB4/SILJaKSuNmnQATMxwpG6q8O1Gg41Ata+k+nHypT41
N0q73wM4lf96Py+YJY5YWBHudhc5+iyNA7aH0AYlPnr0ZDVveBXhoFUVaHPIoWpC
4uHz0s8dI7I7o1s643VmVPmFi9rflDniNC/x8uVb5Ouar7uByH41LOXDfs8juVc4
ZzQ3UjppXqrsAM3V9ZlSqiur737caRN4qDtBeobpnLAowhRTcRIc5Ty32Yp4F0p1
av/u0TOEomGQlhcIgxaktBsYcRl/2cvEcIgOLz5c/WWYp4oayDxRY69VeF5U2TjR
duAch1Eu4yhkK9q/iOBKNheNQUGT+RKVidzroXYAabFmirswhK6XDRGbJZ/RBpFJ
voU+5egJdVkCfJJSDf/BruPLKAvVe6Wk6RoaxUFnvo6GcENl+/Do4PE+3NMJSwbu
GXSo4lNL+ya1PFqmdh7HFsyqMNjQbcJi0CyKsK87DjPhJh7PkqYaossKYhXakw1u
rM/+hSIyU8kWLNhhYUgqIhfQ2UabeMnpfF18L9kJvRI/LuZ4flRVTUjwNRQjvDGB
EUsj7j6hkfXKOKtnm0zQU460hTjffki9h7hSsoJI5RNgRFZbJQpj+4/oDVjJE4Np
3FgE5cp7IBt1YoR18ivMODjfIekyhJHbfvQvKlNnYdQPZ66krcWrMiE0nVBpiHj0
nVt/63hfDCZOdxyHxQ0EnaePyPW9GrnMbCaRni/ltH9eTOQtV/EEzr0F60ALLzgn
KAzURXzWREXGJiGgIBEFztGOV6Hcqs5WTnfs3148DhiZnDtDwGTkU/mNdweqwW2K
Z09i90IF44X9tSPwfwUFCNY75hOE+rEO7qTceZ81Jw6itvINo4sbhrzDNn5xny1b
9BMqtaBEG8hqLxWV4HqLknJdtq4IdO3UTLT2O4+s/hCAj3MpuElI8nVeHCHDpunD
oFtvpUAYZcD6c1KrB3DMSmNq/hB38K0nx+LQc8XsVevWIUeoe1E8hDrVcc4rk5Sn
bPafl1hlD1QGk5EKA6O8dCHe5oUuypjGmIbNDgED1+ikxyhVWnbQAq6xLuES/C4M
1FNGs6qx6ceVdQCqdNomvy/PqwemCkF5moHNExdhhxm3mETPjHJZPA78N8DGkd99
BZyL3Z9a+2RcKiKf74BYG2F4JHXNBFE19FiEjB7ysoirJY46R6a0Mm40y0EmWpdc
sr3ncO3bHpQ1iscB+wSiM58Y2Q4AOOumCpQD5CYYYxzyIyb+UTiBkE0+uw/2we6x
ZmHwaQITpbYxU7+XcCxfCXl5kYEDGy3lWgOh9CLgGAP99pcTvkgPEuJ03fkHbfSV
KGkEvopSAjORBjaZmNEZ7YhM447ZQScs9W9Rzzk1gBiC6hS9iEazk1Vz4Fz/M/nw
zAbIe27BaZMAWvbGfJxuZyIInGB9rW6OY68ZomZLdmhbF91mBYHdDz8WmTcYm3S5
8wQlqajgKPNK9G1Ub4YAFZpGwsYR4wVvQiikgy18KnRHSecA8gJnC27The3mMr4s
50iqr6xV3A1geiirtv3YXcggn2uYgJpGULarR74zx5+3Hevyen7iP4r8Qa0bjD/w
yKOkXKV8QOTh7+295tq3y8nKml9gXfv3m76bGTE5E4uEoQFY6+EmXkqIuGuPiAcE
RSxLY3dtVIA3gdfY53IHQ3+1v3KdWFrb/1EA+qaU0rS+1YjpG/GkjexBJ3jNmSCT
O91u7STLRAN6nZqPYZYNt8xX57JIBQxYGH8IiCQNN9fW7Bm9SWTjfwywj3jKoGwe
Faa8NvOoRyOqHG2S8N9nZTyWtL/yeCAYRfKlyxQbdrBFxcfYx3jFdbvpiGr7EWeo
5+OCD4B0Gfeadz7TyGCTQW/zu1vqOENXx0dcRj01+pyf94CucZBa0GmiGkoCg18G
JBg3uyhq/kzlTgbZah1SxJarBGiBvMjB860IeccBXvMp2CfCdKJiC8XSlruT4zTE
S9BgFL80uuctToSX14KDGw2jRIn8x24dEm/003OyNyS6av2dC/YAeSss2EBo4yKX
GZb4a1aWTzVoztGNEbqUwoAvjDjLJak3lFBIKwxqrOGMuGgBn2PjqoLrgtHfiEWt
LJwB62Lj6R8iLqJm3SFmL9CP3xkHUSHVkIZ366QzJMySIFz/CDK7Z0jYCSAMP2ea
vKSMrICQRcA8CWSxU+LiqnxRz0/mbzCqqxDvb2V9678GE7DlHhZIJtg7Fyp/1Sfz
H1cRmU7HtosBVNarPE6JwoPn2udXAaHCKnrvuWHZFtiZjXt2SWO00UOsrIzMvJIH
ZDBYbO4+DBE/Eprsv2YlkfGjmfEnf/s08pZ6OnWfBUg4SWBK90mbDTt3GzmQKXLq
HPBCC8Tdet8j8qCOXOhCoqzh+qNpQAx5ZOqXk7alOK71hokt5O0rIDY/QYvL1gCB
uqD2F+ostSzplV/BGmtpKaoYt25+8UhlxMtDgVXXqO7thWSWeNn3PipKuxmm9tZQ
KnDBXvlVxrYuU/Gbz7CaQ469v5vrbuLbnLmHza10HEZXv8F7Or4QKXn6dVLAEsfR
cufArQbCvTVHquWXitZki0zhxuRU/6+E44UFJWK9QpEOuHCGfgPFwLd1Frf7+tNR
AzgTXcTiqy0upd+JxUWUbda8dpn6lbZYlIToGMGSX1o7PlR+BhIF4dEyG6nUCdSD
tARrFno9W1JH1ogv3TptP+1uxT9Y8XlDPHvcug4BPopE8A63HbCHwRHit/+coM5G
iBQCent2kYnpqrTgIzdCEaCluImJyxjuq94Ue5JpJYg40TDygP8kQLlybzHZmLGX
DB0cuHBY2UmKK05nv4VfiU1mbLVkPisXj2C9LmqlYV7OGNXuaKl1kaGZxBHoehiN
7Y/Z5H4VmWfoXBBE6MgfqQDg6skd4HBU5YIpFYvqe+FEd3oFktPEIXtHImk320Ok
I03xX/2wPWpa3NHl07G+UQPZsqBye7LmJ2vhMd4ixOB+mfKcqSr6QXeIsCFFX+9G
nnkd02eq2+o+IHhcDC5zZ5pX7AEYSrZJpv9RwL1dzG44vkpsSpRDpirt+gfy7EFd
jzvFHeeDl0Gwjn5Ndji23HGX/GbgeSQYl0qckwkV7NC2DN/VCitkdnCgSzm06eEv
ErwT8Iae9tgYaB2sdi434aaDFAoyyz6+rqP1f38cLevFVU3sHh8kQYx8LdLyEEJF
GR8S78/JrjI+9n/TQDsX+6TN9h6bTWmEdwomcb1jddYqOpmZeu/3avM9/Hs6/1wM
AkO2xVmYzeHSI0AcHkqOwYw15CQNsLte8sn5zw0aoYemWqh3g91NkSMleaY2/r6K
acK2rEJop0Vwy17JW57sTHfqZJfcI+evRJJmWXIfsoNLF7odVvFQm7JzX/ywedGn
PycI2MiuNGGhdH8wRd6M3HoBh/eOjDpdF7jyxggeizHvDA4/Wu6YvEx8gg0rkbkN
keCwsNdri/BvZdVj0KKyRzxM8z0O1H6JPJlSVv8zb/Ua213vPXgUIB4obH/H3r5p
t9K0M3BZM8bAbbtxFAPVE5+kiC1Lgcc5toX8pWmCikh5KJ1kcpkpyrwaXdBRImtz
tDw2HR1w5+r2gInYl7P2A+F8P+83fHRu3wis0Y0QPWMYGy9bjduBRUAySvvDJ+bX
IaTmB/Ua4ELs3ofahQssaBYEpOvz9ltgHLdVzdUdVQMmSX522361dUsZvm6RCojd
kFwadvp64XXb6oRVphD4HdC1jpc9MzjLrJoHM6ldK7R7LVvDz14odrKDEezVniYS
aGNS2Wu5p/2h3jBoT869C44Q8qemCfZ2VnmFqtqyZxTT31QfedBg6MZsPoKrvbRG
nXEWIOq/mVhzWTK2qJRh8qhIAUvKqVFGYd2fHlST6KwsOU7Pfcf8om8qAVKMFH8y
ydCwcgmKHUiCMLDVVKugyvwZKiPmL4SAcf5P19ZZFxc8OJ4n+IYKqD1vsYwXrS4J
Psup9bgOJqdNsPuzDTUCq9HD7e8INrCYSJWXOOBvLcDnbbb27So0C+zlKwKhD4fh
mWeR7Bb/FOIcSxZ4WcotbV8zcY/PDd3WR1g7TLt+LV5fDw8b7Mj+sFLJXnXwLjYy
pt5ZdXvBlSbDsr4QNoi971eRv4asF3aekGrAsPFuujyuajWQORy4RVgP3CJmBbjd
qsc3njPfQwDLO9Jw6EyR6PEIUGkq4ahLrQJOxYe+Ap452ZzpFymj/LmMEHAA7Tes
MGALs/HexHvEibaegOBwWcBgvumog5X+ggDwKd1iltILbTsbu678QIkrNHYkZXpr
mzGmzhCf7jlU2OlYtKEQwXr05/b76p6/T4v16lNDsKWoHwjWyO4K6sZx/ziAa9C7
cIVLVB/+ue2FuRVk2eIbmKjMsqf8khhH/CaUaBttnUQ4Owl7oDBLmXrf8VmljFp+
9NQWv1oAfJWMXmwbK4cNIYrFiCRpB21Rd8ZDULMb+cFHys8CzEEpI4gjyOa0NIJJ
HKOJCpMRzZCt818V2kAQU0kXTZ7PNUUQoW4KW43lUzpu3uBpDtE1nD+pxgQIPBZJ
gd9TI6HzlY2lXRN+m/32ooMYPFcr973XXviuJR/FJDq17UC25nijV32MNU5ayNmY
DBYywuhjfFQzMeX6KF+cojPDxGPVteL+pVudauq4TMgpyqzkfvI00ebh1kB+DvOk
wtbRwIU7FcHngO3itihwflwXOq0SR+dvNeLzzttt2QA9MKfI0cN4Pe4qX0g2dMp+
LB76SgBPHQXSxfFABiJNYwNJ6Vo3ZqmuSuZsoSVc7nMaWyapv6u9CqXgHM9Yv2y6
utnhG/FAGmB/KpUlkPhZZ9D8OhrccWota87dSZj/PEJSD66vN1jmMJh9Fyxw3UDR
Ff4J5V3j/RIo+JOTp45piwD+V8xSeFEgCR5GWaguD800J7yGw+XQ26g3xYsQhwpu
ot7TlwR9oRwzSanSVuILHGdeEOwJLsN1mWfD6N8/SuT6cj+bLJGPecjvUWUJvAyt
5aJ4Hh26+EACvEDEp8b5toQUYZUQKDygApGQDdRMbCzV6pYhzcjq5VtCX6udYA/X
Pw1BEP4c5IVN72sjI01pNNBcYaZfSGYNS8GhrTJ49SX3SxGo4N9FqHc9Fd5YDU42
S0Zl4Pvc1dBWLVgTO1FcZJ0Wbb4vrXn4qYWTPRf8/wbZd1D95hcsMaQYCRmcfQCn
gkLwveIyMaWEU51JdfxVN7+80iDrv9jIxhPoLH3YSAq19MVV51JYSy7e3kk9+t3X
mv0/wlFUbs6E54T+4BFkkpe/V2gom0A9OKmKiBadnY2N6/9W4iBN20rT2LyUZfZO
pL79TeZdiZsFrYxbffOhXen4CH+725zDRBFmtJK+VcscQpRjYexF81VmoG0pswGl
D2Bup7meqF7GpN6V8s0w5fcGq7RgkP5Kq7IrSyfe8RYBOch908doFvsYPC1kbvFp
Azqig2ZIjiHQL1fML0S9ViOtNyFSstL+cCPheD6u7GuD48l2UIuiGQJ6zlROTUiY
i/saQsx4vZqPA8ImtQcjMlKXpi1FUvUWctCWsLjRAon8p05KAcSJvl3QZ817FbnQ
UMyBt7TU5DLZ7ZPMovPazp2WZKJqqaEvZTsHPqHfH7KUjv8uaZZgodDifqoFN85j
/4f3rJafzsUfdBqevIDYkdQEhKzc/TB6svejFgOFJkP1Z5NlO/JlYnNRpfhYOSGV
qbqAg6dk7V7F14DniAL/xROw+mQjJm8rium/hxN4wZR5/wGy/75JSmtQIT3Thuwl
Wck8pBEDWqDmQncMdhdAQUlswhxU1i2197V7xFKt2EbNrVyJPJ+gKn15cV5zyCms
vlDi8mGLeEbIJqJXpmP8GjLIekIJ92bSaPz+ENm0NQPC1ffpr2tgR8ecL5bH5lg2
HimaPC07SoNtB/30kjP4wbV+yBDFLZE1hq3Pd+jv29regmHFc7NYg5G+tLGn4skA
EuJRmfA00CUI/CxO5UzWstb+HSn0hYAFF3wTKzFwAMqzJ+EWHv06FeIyhAyFT6nS
0RCULDgLeTNCt52gkZRpRX6tkzwxIKv5IYgWejdx0aprN8TAxqurR6w24J7FWx4R
fHZQf039aPH7XF+b5k9d8zf6Pz6Exw9fOlNeTjlIwnY5RtJDw75UnptCZe+13nwr
bj5KvRYkCts7lNyWjRg1DhiihFoV8As3sa8Q957bBDR9fotnZnzFuZNVIgt+Y92Z
TvA1TP0B76WRHUMlZtIUEypWzkUjX02MzWKyGhJ1HAd2Z9pQhnldHYlnAuayceWf
IJnj7PdPSYtBd+TKa4gXnEGvo43SuUOmZp3ARwalxobZMLb9GVhW4kJFhY4DetCL
qVsoZP/j2PJ1UhNXmsnFoiq/oKHwxriNXaUmQMZeYC2gJRDD7O2lYFdQ/ONBlzzZ
5tjOI5HtSWzIZYmrZy5DLZBmjZVJeUlNcxmKzTHck2KCa6zgGieu87ApgHDkw+jU
vbS9Pe442Eg/5s6IeDVwltOajY+1GBShbbMaNXlif/BxSUMXTMsqMLyo7y5YHSu9
UWsjtZ+ZyZ2NX/zNKBc5rHtsWHM4fYW9Tw7p5GDZtJWGKgdQ5wxhHoJYXal9wny1
9x+jfXZ9zq8z6Xx/ZCz9zNZkxi1VfrHLg9XWRyuHIIghfnLcwUrGSvNVTGU154GB
WGFFib3DhLUsguUGvYoJ7uptMR6PF5SYpJx2ExihqjqGXl4a30AZZjzZjHJ+gZ4O
H/FnzSRA1AJFK2oLR5lyv5MzvZj+8gN+899+++2pjuD1ucTUS/EnQdxSoAmyjfky
I4WsR9JE3E2lkWqzrSFYLw9fIey62EBbk93N6nMUvvaUuL9wajTsiT6WOehjC4Wk
yfn3+OOpRYF1ZIk3hwuoJuVLZuKK5nhDcczYHvPTKyBpf1V3yvAyQXijmHSWbVsy
R2O9uPi8pTDXBQlQ5BdK8omYgUTOsL3hEpFVr7OkmEilQlYqqedWFjVjiSrgmOYq
p4HcN4u2JivmRDvbTf4c8G/nofCp92d0HK5X6uzUp+kfljNSRkGh1dJ32Ww0SmZR
a8EZdxK0SUtWM+VToaJOy0aW/YgwqLGNbf+93bCkwV4inG3VzivO0OUm8l9xzGsM
bg6o0QDqbzv55WFkQfv+a7whmK1y/k3TwXhU7nN437T3smONcnWfMDLjtHQ7LQou
XhpmCsDs+0S8cQn2ZRh+jkuJwruMJnc/VuWi7GPS2DWWNiGE6Lyc8Y34aR/vI0bq
zMNEoTdXiDh69zvB9+9JwO/hD9i5aY1DvvFF65P4AFUfhvzsKuTFr3NNNE+l7I+k
K54ynS29uisROAEsDYPCcnFP1r6bX4IaPEO57T6gChthgDdxr47ve3uTHA0UdcU/
B4lSFI5JhuPWeL35gtt24jUGMJXHXuXqp/IQLN6La55ppwT07iGgC6PmASy9WKi/
hWXwZRwtjYfU9Gd4FgWPTY7UbCgXpF1PDJVzPTdg4yr60xsr0gcRmLao/9MEBK3B
sQECf0dQ2KG5yx7ZStlvcWVo1noPSRtSJrZGiRLD5DhbwgkgfoBK0T4Q0c8mOQXM
PC3RfAJjDlv695tXQJqkeAFs3oIhxWH7fTXHJExv46rW/jjQinoT1Fy2U/mfvrO+
TZzxGmNfacNCMFtZiIGBdni7HHzrMF9s5sBHprWOcr1TlUEDpXQOQlJ+VN2awfWc
bDxWs0ocT5FnDNbog7KMAXepov6tm8mB0bf8tQHqAO6BbtG/XZiywa4YCi+i8+5h
IOXjP/eNkPLrmQIEbOyb9FHmFaiRZJPiwIbp5IwgWp9gWfLPDe3gyFD3/Eyrq/Ie
INFeAOHdi9+Gc38K5bgwzYNqg/+pMgg5nLrPovZxvaJvG+hHlxQi9NCOCu69+LC2
QUd5wy+QsTDz9Tf5ZxYq63KvY25kxeHSKX09yPceGw96LHNJVriliKWVUckN0wg8
Uik+oSmFu73FaA6sjWf6UmhyPIzoQSCjlwddvRiBoj65poXu3OBRSYLWm6EIQeGx
5kcfsHNURigFRDepOtGavu7hKt/W9rAGBydhDZLIkD+CuVFIGyNlxgBBNZhzHwKK
NiQRo/+B/K6gQJ3Mezh6+tuiLBXm3xCkASeQ0nKCcsWfralgfR3tEWE44IVN+9LD
XZUkiGL0EtnvsyLLw99lPUgXz+VTOwiOA9sUPMoX2rFnTuVVx0iPPy9cbymEG0Tm
PKIsMuEK7nWWEN6e8jO1pKF7K3lOe36+0iKQ2aSk+F30GUzrHKPHSYl7u9abYzOn
16Bm5mhc9CTinVRu89Xbo+cuvBDjnT3H0ZWtEPc4AlWdvxb7dp0U9H0ahkhLBUhT
dWklWDj0lQ1Ry2fkSf+81r3xbsF/iAIwbCd6pPOgt1kuCA2IM6amDepfimmvqECJ
j+yhJzvdoWls+MnnBml7ylPAjsQTPiJEgZIGCmCATJbBd4c0UL/kHFO5VuB4MFyR
+BRwP/n8rBqVDBNhCG2r2fmp5kcfp7yK87rc66lAGbzJnXJ5hfp66cv7Cgn76aJz
mYM/zS5ZKABn9mozPI25j7m/Bfo2mR1LdTfOu/y1B33ARH8j6Kab3qayIE0yJK9/
gJY1DN4Jk9kaPkRxX0531kVTAL/Y8t3DMYdKqegc+hcOwERObaCj0hGPxhbLnnJo
tNd7HjuWSoQsJrWr8CeJqO1u/YDHUu58zAUSklnsdG2BMKX163l0eG87KLx89OnD
VQXOkPyp/CdXU3zhR4X0jKEveYTl2AVFgNRqt5oQCEP1dokz3p2/DhaHs4QG10kd
FYIr0XYIiSyRwj6TKH5+c7Jp6RF419DAqYWjiU/Y722aG5eFWLYLSq9DYxNOFFqk
pWO1JlHcJ3luSVz9d5Q9pux1Esz+ar1/1QlVUsgcEW8bjICs2MaLrZ/pRnpSCjqi
rBOBNzRSKIOhy2JwyIEWqU+WbCzB07XO2vMNCNwDjOOGxMT1ewyqwq1ls1wp3SZV
8N1HAi5RYzv50756kURbwacfhfj419imrc6rXEs3I8wAR4vlWx0YyStMYbeUP6ku
jh8ihuyFVExCextfX62XbZRISbnkQEm3CBaE8AQ03vFz+tGk3qXx6RXPHvuMSkNy
D0sVk3mJ2zBdlXttyWte3PwRQt/Js4mSFaXJRCQhb0eSoiLRBVWDci/43qIZIj2S
daqYkrc1A1tONKKctq7i+vY8jJT1+MumI0QHNoZTmltGIADIldst6ADkYDy5abgp
M2DTfyvl8ktNARVwE9OC7jR223YwzKSE20OSGeizfKRgoDqy6+t8WFwn05zSzdMg
aC4y84cwNURfA4HllVq52A4iSfkTbgrAbLw9H8Ac3ADkxKKX657eXVlZYCEOwhqr
2JOzHYcn5QJEM7Qfo8G9SUV0fx+aKthl4NLakPZ2m5LUpSjG2cM2tUh1120M08wV
rxB34jcCLtqtmsj37CmqUu4fdqQuKpVfpRLzybRsGiRyB8X/fcFLk0rgABtwDe8o
tYExq16pSEUVliPTQniS5aKwHtldOCF/UFUn88G0cn49VjPYkrRSoo2wr1O5rD4D
7HUB6hTE6boC3nCKcLcW4lJpB6eG0Zka12T3YOHjuMlDqCavM+rTRH2K971ctvxh
0SUjLM2S2aD9jr3d2cRKXPk8+qd7rxUtAtwIxij6/gwmjvUZA759HmAN4/U2Alzu
TgpR9kqwRae49yM6XXVKTxdD/RKiLeGFkh76QH2AKPSMLTD/mEaN7h/ymcxSXTkH
sXxjSjr4Wk8PKKrQErwPoYDoAx0WSngpip4jj+zWJLUpxZN/SDMWW4uuxjasIJ+3
eS6DzcI16fnb5LoK/KBq/j32u+3fngqfkpsZlkrjBheEEPbVPui2Qlf4d/6zAbzK
Lk3WP/UN4IQQVm1qr+ezLwYwuoM40M90hMSlQzUL33UPrvuLeuDfcosYQPNZjkwr
mHIa7k+M9nssvFL63yG1yi31ZKSps9DaB9AWuoPYRQOPIM53BY4vITeTrVcJT9y5
r8RoldefycmmzUlOGab4HaTJcKEplsk5+Zbgvkiw2nn+uXuzhZbfdyOnzsPrJ9Uo
rRQnkrrnCPiHrbxEziQ80FZf3O7vCiKQzShnYxFmRR49zy8NsDq53w8WIaQT9UQV
SvhF06qM7s9GetgmKavipXhGGHUJYD8cC4IKCtXJXTiraHyJsd0M4Y7Btbbj3tot
Thj/K4hedpNCsxvc4Gd4tkOTiDlpEfSdookghiwFlIE9Qvnh5Rwr2nVdbophDoVg
l8DIxsU8m1/VbuvDhkSsglxWHSDeNWym6JhvxoiGaJ0qrGNt24Q/CiB923hD3djE
JU82O1G+vtSKFqki5KKyPyZnBqOS9j5nxKIt6HNGKsRZ4SAjSm459NQSb/whvKte
Fk2U/M4D2t0d3WQ7fb4JdCgV/1DI4VKG6e3LH2cQ+Zdz4CuOy4J4dDyRfv48bSBC
1070/zHASMD2on5yXZVWXibrmYeNg5taQYCLe0VRmk9yZSrjwdLbnhtJ820XsCZj
Dal2+21GkbNrGkD+5n3kEA1ge83/kp8qzfXoSKbw6CaovcnYu2AGoUZsivFwTihK
WJ5gs5HCT/K+aX8PgVL1zubovD1k9U5X1JBnNIxeR464WNtoWtSwsWvR4G7ukmTS
0W42pF+NZne0UjooPZ9gMTBRY2pLfMOfgQlbvcUMCaG+6aEepvl4XygpRJ6FQGX0
uoKCXWi8+51g1txmdpkaJ6CGXdLZqgYVtp4Mrj3/MM40e7LfM9D9+raQToK1Vop6
t08YASqIjUe9daAgLLJprpiUVs7bWtKcuQ8oAwuVO+91yrfvmQrq9l31CHGc8gyl
FDpSMBLHOTCBJWdeOwWmKhtYZd49dEi4LpRlEdAVfx2ND2DV7i/Dv0Sns5pRsgou
ITzZ/rEdhf1X3oNfdpWJC9D7s6XRijRdhnQ/3tyktWvjHuGudjSP4Gn0m2jWHGyu
wog9NAnzGnskUmROBsq1d5ZQw4W7Hwg5Ci4XbD3c20aMj74yqJyQFv1rR51wxR1R
bjCd6tquGm3IRge+2T3ePMZYrk//BFLvZVSB4J3vq9J0OT/KVxHAjeZQBmIt1UT/
c8BpFNqSqWuksKFquvWkgvkGTWwyUyRNXUJ4te1O3UUVeea85sD6VAk/hzX/2hNQ
owhOuF4558M4WRQbpYoKMjgpoUOGIPVM2VQ18El8JrUIPWOKygIoQfSWs3VfO0yE
CtqRPf/gNtLdagx0Ybs+ffguomtPKGo5376OAvbIMPLrVia76W64EwJyGuVTeCnO
IM7rVls+qasVtQ2KdJqqZqfxYCRwrsKC1jMaIxRwdcj9g84kgCEx2UEfbD+SLb5+
SCAFrA/qwQeHXFnfLBk89UnGhfKWYP8sTmNw3ytUQKQRSBOsCKPFCKuXtc0j2THy
3LDAyz6wKUCoP5BHXl75et4tr6b4CTXc16/31I0nsVipUFYtXvkw0fP4wG8oQ8ne
9xFz0cRLFqd/bEnKP88+mx2U4k06i4KtyFlxBAsR4Q8OrTmsttbFDawi7vVWEdty
NFlfh7aTuWflQsn0NNFQfztV+60Y4dEIyYCvaCAfQL8OvtruLl/uXCETB0AMCMeO
K4y26HowrqvvYpyxXpf5ih5SrkaQmYx10m4YTWUZtr0rioICpD21t22QMP2lz/XI
EeBqPG1x6lhixMw/1G6GzyEcN+WCRe2gWWVtPctIp+ezY4IBeq3z/MvkSbj/l22x
rH9vrxCI5gPdWILk4hwVtCcTlqAnrV3XzGMdPAGEHq22Xbfcv05aJu752gcuOdh9
YDEI0AzmFjSMqq0GQNcSMTKf7e9x/sYFtkaNMY7KKxYvNZ+/bLLqfn+az1ZymsX4
c2cK2QY/cH54l3oH/vQ4OYh2SnVAAnChI1OfVV5IoHsRdRGkGH1JuHx5l/iH7otE
kf2SuFxF+s6PAxA469HXDQoLs96gEnH+PHvpQqivXV9QK4PPW+QEbfdNKF+06F4j
mcIeldxDs/F6SukACv+XJc2jE6g2ZXA9yGOAPBPtYIhApHpNsBIKFdbOu/d3tKX1
SrN66x35VaCdOGVnqhzA9zmVQe/6JKN++MMDmhhHoLs4EsDbpXwpp8Ff38tThH92
NQvxcFJgMxQatFwKKE9PD90tyN30SEWaeeA2Z8LAVir2vaCCqTNkQ+iGpLNtXrno
t/o2GDLVrSROhKF7NP1h7nL/JQFAq2g72nZl7a/7ggRdRXjdpyKlulESrnlLrFD1
JOzGXPTLparK7uQz7Dz9Bycb5FINPIMIvmSH64VDf5S7NUI1R79F2vujk4sr4HMp
+f6llOWo8IcyW/wuCRyoHLAg4JMHoURu0RreN/AbmVpIgbqZLfrz2YDCztIdnh1R
yvAtnFLJtdPOsYbrnMH44gS2g1sYpSpwqsi6/zq0nNu4qJOYadawGbXaPsO1J7Ii
gNYWXz9jqeUv/VYVUOzxmGLsQAdPRRCkY8prR5r7rCxYG2Y0VlSJAUjk/4nC2rNA
7M4glrdrqBD5TNluaSDU7q73QhZnjZ/C8shKzWAHs71ymDOTZMEw4wkMj39UwbQ5
Y6voprQgQB+jUX2yo2iXGht5YQXOTh5LmOVQZIvc7wsOtJ4Sp7VSG0D70BcoLw0j
ZjgICx0INVD9XgeJoOy17POz9JlrXd8DAOCVfdDyWnynceQnQtHiCQaTSJNg8cqQ
OYp9r56J2XHfcSrvNa/t7GUOAS0kJ+N6ZzYFq6l9yNyhj7OwQ/Te3oqxKSipmbXY
UBUX0lfoI+XUrmEM4bUiK29vxh07oGwAo2dB7ExGJg1auXMRtqo4J/svgp22VrP+
Ji3oxYlW/e22jo9XLhqqiDHHOcnfUFk1WODUIf2akVi8mGB3QzzasxRZ1lz1PgOS
dk3d+cOVJsPsxIZ6oNrKdZL6wqCOrRWIkOEZLCnRDOGvrnxhAmdHGEeamUFVnXy6
c0gV+EW+nHqLnLsHz1Xp0+4CVwY0cnM2R+t0OeYWiTi95SnFxjRcjebmWI1BruAS
bmNbQpRgZ2VHk1+AIIyDLXHuOK6Vvkwo7kXzXmRk4wW7d99mLySB2vjwC4MFYw46
9BJt3JdrYr//LESnwr01LhRC5RtTnc1tL3fAtHpGQ7Qt39Mk0HWjJ4NtsuKRoGmS
5synSTorGwLsLF/IX9R7Cb3WjAR20rzPaC8Nt9W9jhEMr6I1JOVVGxs6R55b8XC3
zRvrRSUXeNW8mjoAByvbjP4oqszTO+Kpzlo04h94lbkz69HT8K4PzcRrw8zxnCOF
8MKF+9V/uM3nGkKsno1DcrOLFr8lFbZJ6HJSbuZgVGxe94+qdeAcp/Zsklon2Te4
hxWY7jCq0kSgIB9WYTrVtUatcQw/DEIOnYzU260liN4DQQgx2WfYyF98dUUjN7gd
Vj+buwV3KsejUVqSU3RlLlREN+5c8OXYkDmuB5v8ZmGbe4DuXmCrRyyAgjUSdgXO
VndV6zP6qZmHJVDaR6Hk/25qNFLxI5pwwYDcV39tg08UFmVeVbq5q9UZS6Bl7vd3
BnITIKrNFBrCicQf1o2nYNMBB42fIyshS6NA57wFESncFs+4Y5ljqLKAKNSc/mEM
mZMNg2lwRjgV8SjWL26vua9I/JVD07voyigu4csM2b9067FbwgyuF7b4t2mHL3dc
tO/bWZgKOjL+vReRUv7DeJAj9RUwI1NVOHDEtHSHAJNGq11GXXLIPMM83/9UML7Q
7wvpn14IgNHm8oYBa288BO+7st6pFoFt1sV7hNqqufXQXYACMtqSyt2eluFqKrq1
jle7edgIdYu2QSA9dJF2CLkMgDnRg0FwUKnWybk+QI3Tlv44AQk4a7GY7BrV5goK
7NGJ8PSx5PRW5OZD9pGmJm3zkFZt57eZemE48SqIl4OA6zhM/gF/qviAB5FcZShX
SSheHM1y8pzizmq9gDSfK2Ffebf7SuaFWm+9u2bpn3InQWV7xDoYGkKxRBKfm3VK
eKVz7C3YtSxw3kjVkWGuBYPBTEkqTZuEO02hNXpjhR9MKDtW0lhJdcAYxGz0YpKI
EhavzcEEV6rRNCGotCOgsB0Sp8x8Ir6hAEmgIF7L4DJzMajY9Yf5uRF6LOjzOtMj
N0RQJtcDPsKO/V/31fOXcB9Rj+mHpH8A/r5MRBPhNLFquOhVtuzngxzLC3kSiGEu
DOKgp8rzfLNhDC9GrHk7Xu0eRuw5huXsH7oKorHPqA2V78IqkK4f0xCCS7OpKaRU
O+j3uhQy4iQuR6jom/6zDVd1iFPqx2Jg6Rrqf9Vh3rtOKR3vmO/Row0QRLnFVmvh
4OvZx+kfmFoY6ZK46I+vCISsGnKhpr4uAiq75kBvTTwH9MvDKU5oq+h0YNMCApba
sheVSVn55FAZpOSswfRQBxSGxqiqnCsb7vtJaiAQp2k4Q6W+PLM+rY48NwsQAt+1
pgpAIzkDUZaZ0DNC2vpWp4uCgNRs+lSrGSsGlFE618rnSrA6JNkEeDuZv9mAGuHd
DXzwrR9M62rlXFQuE/5B7RxgaAeEuCijTGA6arN/FKuGajYGBgdjRTz/Dkl3/sV+
zETc4Ki6v7p+QxSmKRw+VFiFne0NChaLcws0OHp+emtNekLpAz5D3pC6ztL9Yugn
PLqfBDhEjQr+fEKqnsMtzMNdvh+Q4GYb2tgUoQC0Jy1b6lO2j4n0Q4h4kPYRRvga
s4UCy4Eo1/Tec5E9IlECORlQ7KEfd4TAerO8yr7MdXIrF4ecA03vABmD2FwLWahe
lBsHGMbryytLEshDPgMsY2cvouUqoGubbd4ZI7Q6DdEYoUfRL+/JbULTuV4Mk4oG
5yDPqc9/LEcSCtkRbkaMSz0/pRexGw7h5ok3+WhtLN2Yjb2ulYzm7i9n9N1NhiTP
Frng3DLJU4HuIYgvUEQWhFXI2V3GbCVvOIJYi+x/Td2d935qXN3QIqGxE0OcvMDV
HacrXSPOCHpGG9faBsIfJD/OASao133e98farQDTPYJBF22VYwMS0vW2tFFbR+la
slt1ftzpbLdbaV3ybemHwSgsl4+7eJryz/OZdsKGrDy+T7kSiuTT7lXRph2uGvl9
GTdGgw9PWpxEg6IW7f5rhkmRds13TPBXIV8mx18K6zoYf0DiQqmwISMMmhsRt31u
Rb0J3Idhqv8xkKFASLi+ICN8nxTZqaUxXtKuOGHUdRIhVMQIYLAGP8MMCbqs2PnH
iPHRFMJKqwC4SQ7uixno8ySYycT4MeSIXdKdYodNEwRwpa6VTpj8zsDJf6eNw9PU
NldtrVeVIXNjBbDoeKmCwNoOm4ziFGJVKvd6n9zbZSbq0kICFGNZdZa/zJmLkfeP
2j76Z0jGwu5txU4bdTMo+qV8vAg7AmqoYT65h/98OOCefUTrJspZGCrxDJ5jAzYl
vYX1/7nuLlsGXsB3ASARSGGuwuxEbJj11jEaEht1YSTrLHEc9M3nm4LonVpGBbZ0
wMhM2RI+6RfE9gzixQihV0UQ7DIpi3Pl5XidLmvc4F6GJYhqdrfB+Wod+bXHVr+m
dcIRN5efPaUPftx7fHylA21QMtViJIbEHDdX0IpMTIpr64oGOhK8LkNVqZevJb1K
Mi86+oozXWLC0wucOO7eRD3I3YqvCv9dlvp2KuFkYJhzNqLmNIIrTn5u8/ZWQUJD
3iYrl6lh4tYoWIHg2W03hN7JTWNL/7jvmqJXGtin+i9mhOO6mJWj9eHFi+AZ6a72
RMd7jS+Y6tgnjWu05IAAzqORjrSDUUTWLc07qxprTNhLFZTXnyUJbJtzweQZKD8d
suhIgy3m1tGXTZP8AbJXEHaJ94SGp10/G2I9UkLsCJHNLlfzA7DDh39e2/hCR176
t4Hm/BemiFEsuxCCwVMlj9QFEMT6mf8Fa11g7MRA/zxCMIU7r0hEvwuFCjtXBW5o
QeVT1tbvhfVMu2bgsqUTaxQka8k548Hl67WFjPKxui/1N6Fbx0hpg83JUMdIl9wm
1SqEI6feApVviMf0Akg5Br2tz2gEluFXq4t9T9kDQClyh2NsrYcpv+33TYqVplDa
m2Wfto5qxMSktwtaZaiQtqTLdr0QP5EyoEzomV1jt2jY+zL7SiET7JecU0qgemCd
sev8F1u8UTFZ3Ofjpjn256HylW6Ye4A2Qq6ukWEaGnI51UUaB0zF5ekf06Lj5dBj
rhdf6ehgJzKCwrElxAbb+q5m7FMHlulvTSs1W5+SkxHQgsseK0Lda8pUEYDy+sEe
QAZgwvi83ZySFeV1dlLEffNP1gtrLzZWF+VtRjSXLYEIziOT0k1itLtW784L1N6k
FpZgYmq2j8F60/MD3l35YFQWFRRN2MRIP7tb7eQ3jZRg/DtNBx9+PJiYPfZMDgjX
niPqU1Wqzkp8k+NYGUtBvG1KyLTmkL+N03P50fy3SmjyD2p5s8Yheq07G9dnuY7G
MMK/7ZNCngX9f/rbFPVpGMERu+sLMfqta97+buhrIz2P8evKShw93cH5J2sVvutI
66LGj24Rwg9LEsuY8AR+TcOql8INAExJI00dN+0h3ltn/eGeIjW2qYvtw+yQ/+gx
rn+GjqQ+CSyKzEhhkcwSDVDvoMVwlTMUWuZu2tx1a9f7DeMeH/5tPVZzZHe2JyGe
7fHE9o5NNCur9fJD7FhNpw3GVQgSL84aEKC3N1mPmS/9ocACdEsVah/SSqXcvXU5
1wQfGoTvc+VAC09ddQ5185YUkhv3qWe+zx4dM5e3ARFs+lwTI4UFycXgRTOtkr/q
MI96eDdSofBrg3HMa/kjGz9/BWWk5WVQwMmiIrlUcubmk5BfU6kNLel9Doixgi0Z
QdBgMpdSoxm7Lc5wusEXZvqwkoNjfz6R5r4ktQxRl4Wyivumn0E1Tz39RQPWCQ9B
kwuJOm4fjdurTGURU99Ocf5e60OAN5biH77x/4xSB8xuwOdLTkKXdyXjUE5r3piV
bC+X7N/YwileF61LprRET1o3VDwmuPEMB03pBwYXBHs7Q7aPC66aR+YK+LkOTdDq
OGSJMeB9C4vwnrjTLcsi9kNBrSQEk8x+bINUTLv5ueVlXVHDbj465SvZoyr2bah1
YLKHKyRaNoqbAW7V8beXF0t82YcMG9nBwbhUyJbSJPrFHaTTT9ZSPzwuOLeYuniG
9hr43DILyV3UHRXvqhKKM6ado8kKO+417SkGGywhPpxEdzuvwcUNL3R0BpJFjHak
8Fq9Vvp2F9NYu75MrwSZEtuhCpS/hzv5EcthyYOq00OrJcXeUfuIei6j0s9T7E7Z
RGU+d+P3bw1TM6t0MCTKasYM46/YIlNz8iZtCB4lMbDnyRmdi04hcHWnZxm4Bszt
Y+VMcMbLXDZ2oy/L9tn+u3kAsv5g9J+L6CSS8AIOGIV8G/GQeNWMmRLiW3XicJ6h
TQRv5WE2tYaDWS3zl4K0vKI9bVHPIWGGL2ljacCsX3H7rG1j6iCExCmR9vSP/T/J
UlIRSFvBRVgjol27J/wEmBWdVrOnCKMdKPHiPNvFDKEKQf9iJTCmJZ19bGDfelNn
JO5T/zqjh9isDY6RUrltNjiPx1F1C4YQDHIkBOdxzDXv4hjpVzcUUOC/BO095htv
aikVBBdSv5p5ljHKvfpoyA0B3EiSBw1LH+fTI3Ik7Cu+Tv3zQkdb8fJzBIQ3WXow
fj1UQgTseGUgeUvTPQr0UYUAfl8igM9b+rz4B+TAeahzZtq4wDYtWkuCvF/Crkty
8moDn60v5V0LrVfaUr51x0eW1cV5tpOIP1NigpVJTcr6ezzpJ7545qeXUQAxRfwK
A63H+wrkPbUFngGSoYc7BX90GHuqMF1fIgdamSHw/gZNjyNKmQzY+yRJUl9eNTN8
bPAykMAGe7rMM0bPJMJ+limqTmcxcrjwIi9HW3N0FXCHbrbNmrql1wqEwYOkHVkq
an5vzDr8Gv5QGqmkyAysNyC7jpg8rYBE6GzKmrGyFOwVogebVqPR8i0BszBx4kal
K6vrMUV9Mq+Ch8KBkCjXSRU0dSOIYTNWDxj+oethg+N+IbFYImVmb5XJ/iJm+2UF
ZIoXStEYU36um1JE2Qvm4WYvftQVyCt3DLFesEF0IdFjBNehO0+y9qJKW7BnKPjW
dqomQhU/7W2tpZrqA+tCDEWbM0jfAIjB6R7rkGTKbh/Dc/luSbeVV8bkzsloPgI+
0bSopEJZDFS38oujDl0bt0Ok1j1DPiApQyiOV+ObR35jGjpyU0Dwbd2O3zwsK0A9
pw6kSPplBiG9P1NChvM61EImwkqMb0uM6kXJhxbsw4ZcEhobsfpUey6voQP8cIMN
wDPLU9dOFn7bOi49Q4VF5F0Vjs8wXlan21eKeFiSWWF5nt3uXrU42X7RnhAqs27C
blGzSl/m8+lL4tu83zAinOhB9OxRCCEawie1n4gRx7dtTqkR2Eyt2Yq4vL+/Er0R
o3S72w1gD1q5gmJzfq8t4Qp+oXo/mVbuplfOvky6uPn3T5PuQod321mGxDohlEAv
UPcwC2xlrek9i0D0A2az11EiOQmyEOHjXJsoifqUXoV/E8pm8qQGW2yqIRrVqSpQ
t1BjxOLWUkkWh5YgZHYyFWjFWfYjpxHLpTqgvcSNtQLzM0otgMcbHH//4ui0owcg
IDqPd9pct+hyTeCDAbkXucUhtBJUbAj3zs55LJrcgw+2UdR7bJ3yCpPNOda6b9H0
xbHY9GO0efSBbHpYvKRtmdbpqQ0UnHkhDlfScnQYXa5jgGe0uJI/w3VlNj9gJfja
25+p+wKuKMmYWgxMVUr3MWxYH5ciN0RGSbrl+f+Md+f/sjiovbqkhNHlfgLniW51
6qRCxk3PfYjAWmKvy2SfjjdZ7zx6vZS+UMIt8w380ax5ypcXeNOfaQvkObaeJ+66
fTq3CQgO4gCbp3f/UcnKWUlp3KwQoK/q0IBO1YdJZr7FGggVet50fkzL+jyZpEZe
A+7XXPu7lNyELEHzRaP91oOwAYJ+EepHcs0hc7eFm8T2DhxCJyz6eMuJBF4eEdj/
pXEXtAc4GbMaihr89ABEojr9ZYK8RyEFC3rvyuR3SXaE7h0HwjXJnUXmgvTuZT+N
f4sq0hkw8Fl1ehkfczdk4FnvehCte2MQnybic4TlRAIBE4FduhWRPjhBNDpT+KGp
/Fg3HemmiUHLTDPFpv5vKkqCA+vjEPMRfPatyLVERhQJX7ge3w1wUw6VZYKXc87x
vIrqmTAOZVkPYxZdKUL8UnQB/0xAzT79MvMiFjmbU7BUeKxwbLYUSX+j5VwEDU67
Zfy0znDTvB2fidTqed5XW/2Lq3KOA+0+RX2ymMb8Yh4/jAHSTf+136aaMZZG10du
xVlzo508CJ4rTS5cZMX/3ailGPiZ9LvbLPChx4mWTM73qejKIEhkSSMbVfJTT9Oa
rfonTQ+vWa17BNiz0aqybizYJ6f5MLBc4RRrLD2mVHHxLDxcrz30iHh8YhFNS7r8
ufTqQ2MFbF6BbbscCmKnyl28/cyeTp6Hy6U+WeBQyXNwRVdejsxogqvbJ2Ud2Upc
kLbDTjpa9GPkP2DrVzi2PiQURJUlFs1q56kHuZTC++/4D31Pg0qJefWoxyEtrFIi
se6PbR3eTSJE8I2YfkhPjQO8fVmKU9NNGrQ7UlbQFQwypmSLVNHYqox2AnlMBHQV
G+qkrQFD6fTkEiEVHY383iUmyKn35XzsnHuikCUYnMjP485IP/xJG7DCnOC4zc9r
XRS14Z6QNU20qYTTS3FdJy9PhsEvAEKQW+BXOc+Ok5SqLeMOUsSaWw320DV78cxQ
hewHvwKA4QnWeDCtn4vjBwySPdXIzAKqPWzxkJzDCUcyRwjHiORZcfgqPftEdwXw
zTRc57BnIWLoGNS9y5vnTK7oA8L/erjjMwd/JXi++vOWg2OozEDaW/90VeL4VOOm
il+qBATDP/k5phcLuXXqQ2KGCtWeZ8V1Npfa9fD/SahFdTCncKYevq3x4QCfnhmC
sbO1eWbJq7WExJXy1xBdT9OqXvtoYBNU3m50B4+2f8tw4uKa5JICZ9A6hnP+Aufh
4PGQ7FfMUtqUpuFqNFQiQSRy87E+pEn4kQSaFhfAnMR5bWtzEV2yA4wZVm0pOftc
jKHJD08njx2hgOPmtpa0of3O9CGHDH5XXL5EyEtmvuYPn1WujltNAukSmVK1O6bS
L0CPTPvpygY8PIXd9aTVW9YGIEiL+nIxYqvvLcvwrtky/pwIe8L04SYIxd3eYSJl
6iWkyB3AFgYYI2kV76ashYJ518q2rDuDno38Ug0UBueolKO/CFyy4jEIKLHv1QA0
80lWcnAEj6ybd0ymq/esVPnJrhEoUSPFv2bcFZPzzjzVpy1vWxThL49XaQBtoR+W
Mqhgprjv3bj5ynOK4OUnELr9rbkvwH5h2s+Ds8zMLe9zSQJNUVevoo8q5QMKLEQh
GonVEupbUsOlGgYGoYhmlmVBzk0CksALhDvrd+5YPdeb1s4+4HBbqWObSIhYR4aA
228IIuCHJ4d8WOcfkIazGuvwxkVF3bgF0IEu4MT7efXURg7Vh/0krovQqrkEHLtu
FLxvQqct1rfgvbIFoVVGqbtNQwxAnwPiwoEXMDYkU0uD/HBT+JocxIyItSfR436i
0N2Tce8gXchf+M9eOx1o96cfOzuCbydGifOMu25ECsOffO2IF+KqoLjXFEmu2l2z
FhgEZQzNG0glZDWbTApcJve7jk4Izof8n4Inxwb021RX19uzhjoAObaVMU/sBPOU
hrgocmLOmrs6khyVun75ISk5HLqLaxCENg7fa6wFk+buevM39nbfAhGwk+OwYY4c
XLDvpzUNEERv1c0/UGUwpYfmnahI4YFcCW4rxH6YcHCYzgquQy5FSPzIAndVWiNR
rUJYBpif0ZOc53LsIWrl5rv+AWnsfuemgy76XNZFZZzwctOHnzs36WTP//ESWadN
a0LicTmEHAfJLVAcl5vCNJ8iTpdPs7HacuF1AEVVKjdtsta7LT2NRK3Zd4fZLZw+
tQT/ZCGMTTmcyCHKL/mq3AVGKKJwJ6etgafqnA6/nkEVpuINqswvfK9ZjjJCRkKq
xYGRX0t8X/kIyRF0cT9T6af/AFOHZ3ixfmRf9GjXn7o/zwF+BRBG+aMEhNZw3UeH
55D6w2Yii//s0+RIx+UUA7z/YLi2mVr/yx20x4DbWjUkacnhh3Gu90GL1oGSR57q
uz2DyWjHBptOTIRij4/hlVqZgUfZJWbeqDR4XZWMWtASGribZce5CHpFWfXjxqaA
GGtFD5t9ODPLEXWQNBQEsByhcGKRipzKD584OKr2smjSJ7OEYwM7NlWoE7mWuxkk
patRzvXZLaHCOVkbOZkzdAec3KEVGQJdN1WtMmHbQ07SYlP/nutkrjjbspCq3vMm
XFftWzfkUWHxRtpTumS+gCtJS7kfLrXHDL3s7nRkdfKjurgY9xAcP5dB93ZmLHYE
Uv6c79S5v74gqliGFv9v0Ll842mTstuCGmYDOO91oku0pspJ4rDr080G34vEmHVP
jPB4YKYb8lq6JohkCI7zS4QnKgRjIQ9ExPbg80B6nkTiB2rMmeOACFxLiu59KcSj
HnGvwLbESjSy5q750AQ5rsrbSpJn8pfNDmU9Dwfvi4sUmhJxlJulnYAKYyEtad7w
aLYjI2f32srSIg/udBXd4fMb10ptV3Z43OmIiYgIsaIKVhVFNV9WEV1T7z9Xv1Ic
lYgQ00lPHNw7MzjYOlDUr2Xjx5WT+q8eujJmrsGDUf1EXSzAoqKgasZbM9o7CIoh
FNqdj+SrSOT1aV+qhAIZ3oV9q0hVLyN+rEsMWlc/3xAOMF1VPj6Lb0UH9mes0dkW
sQw12n+PJTU8SGYBXdwxJzTIQPFYM0CjOtMoRLDCWinutucbEEw62Kxb33mYhl33
j6Hpt4A0dgHMT0+TjbId4bB8AwC/lGtQDuVJOrtzX3+JSdLBB63XYXN2YA7w/CFZ
N2qP9t8/iIBrX5Q8ueHtPG6LFQO0cnqq/VYTPYGRsAvzsd6CLfyDj1JvynTsxkK+
RRglW1qbcPlwDuRykeza+AHVDM9E3j7XzsyHxkNQU4XMKEYxL6R8i06lQzxx/ES6
vphaO358lQSFK6oKDa+1dr6g+4tpEvho1pq37eEtuXlM25EpnX8yRT9bg5fkWH9l
tm0BTh2y/IFf9XUQcH1Gz8ZO3HrmtZ72kIg2V51H7knRSAPRURoBAB3WgFVpDjFK
hLT5z3p0L8isnF2i55Jj3NZ1rElHGROQYrjayatfRd9mrssnm/2GhSCvY/NtiPMR
eKooHRINtVME08c12sW/3op9MYcK7N2zHOBNdRPJQFyvNZxXucyh9JzIqfPw8sdu
LNV2dUSkhuazyDgZUUvS3ogDLz0f/qWcei7RpzRseTqB4wLNqyKdSBbqNDP3X09q
uAmGF5DQ8YoQnsUvdDiJ8yPuC+hH2uh36m9bB57LqRhyZCcNjxlff6KTq8/S5BdD
/O97M3/b5V7QN5E1ylHnlh2+pqdQIx+94tRAxEybctw2wF3ggkHwJp4pXhSSUayF
zh1f+AM8vaPSld+/EROtXIq5Yzg+uPHuYEbsL+ciiIb3TKfrDIftN1QgMleozQc6
CRn/rM14D5dXKN9kQ4w1xlSaJmc1AnsLFRagcsAX0cxMMxtNOXW0uU/FbWunmFU3
ETj1Ut2aEYREwfw+ipYIkxJE7XPW40wPCc/S94I7lNmBa96n4IGrfnL1qwa3W4oc
xevKhp70XhIVnm6rN8R9s03WfhGXHQgTosLL/6v0FzZrIWDjGvv1oxKqKSSZHNHO
AgFQVrvLqJpY9uoGBAZ06BIYMPncre4dEvpP5ZLgd0TbuRbJ8tWL9I+KG2V8YeZW
5DqA1Nq6eiXcseHMDOgICZBeCSzK3Wd+iim1m1Ut7DU+QItK20PII3y1z/+ctzJ0
Dt4h5VOxFAy/GZ6QX1aww99F2VsdyZx8IWKZNv6jmVfOZXqgh2vuRzNyzKNwoMKN
M542U6wX1XPYgVlqW+6KOG188Nqorm7rULuDwvIveOfEmzFB6Kixhdu6iAzVX2Wz
cIkYWUMZn13zjee4HPjWFTERGhKtwKMrJerEjWBVUH2Khcmvr+vX3Oi9F4NJkW2U
wt7oooPZJbG31MaWpkJfn3iL7Wqc8+PZ3Ubuq3M1z8IvXY6nQQo7bxgyVuMaaqWf
I/bG9Dh/49G2QUexGGG3fK8BhX736C2BE1q5U2yvk/l0gQR5PrCNapqVqiNPc/qN
0JuaeZcmq0VCqXfqVSocNQ0TLElbWnWcR6YMOlvBx6nrJr4Z0y0W1FvkmoUrlIs1
DylWe8PFeXql3i7gtmRUM6+NDkV3945LvK+zPzH8dePeL6VSmAxeHBOSeVIh0Mjh
vRxyeTwwyrMFy6EIQ4ZIzwt4lTq/VAJe89wJN5aAit/dBS4M9FrDO20J7QuFESjo
dIT34cOfYwr/H1zHbdYH4EiMKWd1tc7gpjw9vVNcLQux/VfLW2cGxPtuBkRMnZIb
p3P4CKKKSj/R0Qahc+u5L4QGIbaaq+i3ZPNF4WpUaptbh7bLogPrj87ECkisq1Oa
dbuKSZCQ4KslUzdKuSaPEksDsGq2QiEExKwozlQxvd3jZF+Aft88Q5ukGn+/PiKO
+FEwQRcP0KxUDjBIEge91+jFMgh/NgNRDx3CRf/sddznbz2L8cM16ZWQDRaa71Lc
FJguW6HBV/D7d6vRKOfbj5jW/qyhU77ZuiF2T2vNhinw4EGTxG8tWn4dPna9B/V6
2akaSedLMYj2bdaxJMmbLE4eQYbmYmci0+BWPpd5hpwbXUAJC8gKWB9vAEnwUiX1
VhFme233tR8hNQX811GrFFHN0U5hMwvJ67eeOY0+kpDi0KX3X+BokOf3Khi4GjVs
uZ1lcbHFS0bLYt/zrnzUVWV1f4ltW28YnZRXG8SxfYufqaKuejxZ3QFWo3I2HCIN
QjYp/XUdQQzREVxJM6dB3KbgbGYobQdfFvLZnHOiRWZzOBF8Lf0BPaN3YZd/APpT
WdQFJKipjSNzXOSNyX3xwrRnq+p+Q1eO1jzc9+xAx8j9oKoDgjTcd6jLzet/SVaD
BlmguHWC2y+BH4zou37CNW8sUe4Ka4MQjsbnDagRTV/YjSqDN7lq+fMkyZ95wXyi
jhCDTPOv0D41i3X+nhF2p8er4qALfh8O+2u99CX4Gwy6lHFYIbmvBYCCDzAaMeqW
3h86jACrqjlWbFsKkZowqfA5U8YAm687xdcuSuF+sDOr4OquhNDlTh5tmDBWcLpa
iSQVZ98cTa1Sa1anjfVChEJ/04mEnj5Yq31s0rUjaCo9EF4RPjuF7nIxvzBvIgzU
C1uM2N1oWU7u7iCbN9Hiznc07IhXz3p/Htdpg2MxEU282fkVN9DPubwscW4/o+IA
mNAvUWZ+6wkNwQxYuvQStRz91fQOFucEnemZKzTfo+lfSMA/k9P9CCMBrUgPdAfV
oMG7rFlyz1V0uoPV6ezV7LUlj5dqxqd4IpVHE4X0WxwF6Hc39+EfhdJ3wT/u2a5s
WqcP5FIfhhXMOatlhoUIL6VzCPRpDsLLNIxZQ2n0H0/DXEgS6lkFskWrg1lx/LHG
xXxBCsiWwdKnaQbVNspzS3v+mLHzKfTdAF04ktg+XwM0bMfVlNWMyhbJW9PlVKEi
ERO3EuUsnQGyfbqy+tQ8DAx+WEqTNXOI/ZhoGh1mwGcsCUTb/M7/CzsA4PBWYSHT
hpuwtusPQpSJkT6DgaZLrPD04iJIW7Z7P+SS0g38nGzbPQo50CQXKvsU3tTw51mJ
bhFdRn1etASg6Y3cIDMQTCv0tdaiTqWSLftCpFaaAd72fTEv89bHWUMhLhnKCbGV
J6Oi4o0Zzh+Rd8bGp3KE701dHgFkIdD4/yfsl9wm2/J/kB0uLHudrErkH6SHWKe4
bVD6ja7u90INVvieuK8WUg8NXc7h7yqlMNomMF0fcjgPz7ElyCB493PdjT7kA8Tx
qTQeEFBHZtVZejTePrhyIX3y5pHyVl30zumFAo4CcGp5sa6/G/fb7Ab4Pq2qekpv
wl3o/FfpSv6wdW8JIEPcNlQ74hU9TYZBUwnWlNmukon1nHbSZ5rLg+SvJMWDXFoU
lz37Rcdx133uMe81Uw0Mj45XG1oADUUa51dTryPyNb6PuSkGJX5tXABZebAQYomi
3cxHFMJaS9/yYvt/geRU5u/q8mmkr5262VaEbXNcUYvIEgWWDFEenD0GHzXyHupJ
AYXqh3jxNpbnlQo4Alf0+eHlDnDdkU+ceSeg7Iq5vvEhraemOo5qQpzvYShTjMGA
3/IOwk7uGDJgajAL92Jc2S0mmrs4jl3dT7Y3RIWSJZFlpcHfxbHNWts9UnJL5IjE
TCUkSdZn+0TCfl2zLTUTDW46gspnzrEvT/lLJ40EWa/rtf/hrl7Q7XB7s5i7Du8f
oeT1OimR/64H/kMWjVdpjC9wwfmFxH/u3EW4k9nESjC28YrmHiLS/5fbcfA4EsWi
ufUc86VRc270ly850pIv7LfUXgEARz0SN1clybRpZgkn9QhGFCSrX3jmtilt+25n
zz9+n2EeMVCI3pg6tEVCIXb75DbKTfgb8b/empa4rFCDdXlG00HZw3yVLQpB+wO6
DZ9Bd2PDgNYz05UyHJN4rlbGrDlXAldkzjUrxraf/3/YR2TIpyN8PTcrLlJfejgw
1R7iZVjoBzBsAEyEvEeDlFrn4CzEF2GX9ATjLiWQlngrFaAbbHerXNZkOEmqX2Qz
WPBoa53gKj1yL1s+kruUpVMquIeuPgeZDQYSHH1xSMmBpVSqRh2mSYFj4JZ3uqMD
Kmv/QofiRNMQnp8eEHIxUak3yvUPwT5SAdFa7U3nnv3bLB9dvWgZRbyYZKVhSPcR
z5Wf+JTmyu3FOoft8oZ5Q24M8YCpWvWoZoNHf1UFtUGqbOfPDAPPZB807p8yLnyh
iHUbY3nZ3Hwp2dqvmvsfdbwqTHqnX8bqaGDx2esnHRwb/EFH+AKwBHJL8RGr7dtX
QjDnogcEERA7ixP2OVgCcNBNoVH4KxXEcDwshEI2zwGTCCEDHAAU4Lgp6kGwwyGL
cK0L9Ryhx2AuNAL2cPmntzrAgBkGss8RQEhEXhPgH6U/x6pu23jadZNYNXIfgG1D
13Zw4u1ZRbFlHbMSjkBVtp8ILCgt7h7p7EyseTf6jNBA+uSB+t101uj8yTbed8fh
8I0Hv8ICsz20pXY4AXJmGddKcyoguf6ooxvt879luth/PwxuAXlr8xZklpg7jcqH
Ff+zFe2vAxfpupswhvh3Pzjn4F2DHNWjTKQJVcNOIlOaKzJ8K8PJgtxkAGNw15ri
MT6wbFAQ6XM9YUxhaw9URglOjdUdR64sksISbqc5gro1aLwwTehLG6hNcYSiYT/W
LvA+4kWmnPEVlIcsJLCbsbLPeSo5XiPOsFOHRZO1Wi88P6WYZIoknla79hlXbdr8
itIjNC6Toxo26rcZGe46PfNco0osSEhFT18+T34S2zaxo9AwtEh/G/v3h13icI3j
IPELocM5HPVK1CLMPlsmKP3onNQl9Tx2uGEQ7WHqjtky4YBcPxgwJjz5c8c6K0HC
hdUGcTmLoZbm4mvf3YonivtcUXiZrzUIhZZQXFwi1kWtKYXOcVIpBoFukh8tZnM4
CxqQ3YF9jjMahknBY+4SKd86+C9ZqJQVMZ8Uw3SWhkXUQ6eHBlOlCOzmzg5uEajE
ytV0xwU8e8xQYC2IP9FvWvFsla+OzMg8hXQSKpvQmG2hJEmrUhlTtn4EaHtwd+WE
GV4WA61hSXFKpjKpMADit3U+gsJ+rf3GlysUbFmEzyo+ARnUI239iEFrGmGWClAy
vLqqbPlO2gJ/lsmVFwGcWe3uNC/Gg9YqkXRjH+xD/Z4BinPsSK5sEaEQeWjkCcck
GovIiwZILX//sz0EEc/BL92GmLuhZQvo+H2xVrzlg8hz2mxy7MQw+n8biaxeWg2R
+Ypis0kSzRNQ5Pnn9340JA28szRA7Iw8egfJwSJU44ZE6FdkOqz7CXchw5fSehuk
ZNAvLrOZb+6hgoKZOPDHzlXgZ/w+1RmUce9H6uqX1FpRyFOlLirgjcJxDNI5L2Ur
pVnGxOULBhEPMYyWD36md+vIc0J5YxjovPTfe48pTRGUQdp72B0xl7qjvo1WfzzT
7+reKL7VljbrDkxUiHHM4Ut0q4ZzHbV76c5MEBwapsjvpg48WLyQoin0VBrP8dtn
u01EL2scmExVw02/MFFi10FwHbpD49p1FlkDduEHuW44wnNOOi1MRCeCFpXAyTEl
d1QdEIvAzMI46cbQsAxPQmWv7sWL/dyRJEmdaN+vuIgn/tEsGMFdY+JHV5xBCkK6
0InTUeRA+eK60TLFUujJKucNPuklnsuU9zeqVSzC+6h7ruzexDw24jCUaTFHPCVt
ZdJTx4yRTPEdHRfHFTFFNKy9Kzegrgmu6F6hBW7g42YMZlR0NJxYj8K40dHMFkzK
30Qcal89KOx2azr84bnL5ymsYnlU2KZhdIupBeJsJUOpCH5R+KXWCzrm9iKLNquq
xkh4cqBlAxesnwDLFimafBaKqb1xek8PWMUKbp3qlHpDjf/Tq+NJZtNcJEyYK87C
vdKVRvxADhzIRS1/AoZxoLbaV1oPVqka9F7RSjJWcl17VzL4PrjxcnMkWlBHq4tK
ZPACgYqGBbaC2i0TujCnZ++mLFycOf6NUjJQdYN2VWFZjLhTVivvZMZbW4rUEhRh
fHnUcB1OQRtm9TUYc6YlSUEKLJrnVZdPXyngVOTF3ZoecNRxL4rqau+Pwh/+nJdz
0PFvqEuGPFw/ylN8cuD51bsW3OEU0bF/5hiGONopGOJ2x6oC7y6+le+ydGL2AI4Y
bdDS7ux0WgA26NWMUtI5ofpL3Up3xjy11DREAja7H0RNHZsVVYaJmFex96+El3rq
S61NEeiASgTgqTc1GFGRceb6UXObQXNcgq3Wu3X4gV+sszsYGGPolyFgWZLgWVl0
6Dv7U90aTnpNMCz46A4rxn0ImJF0tee+n9IvF7vQvjwzhsGTqPO9nXcoJBjL2SBl
IzDgNwuVlfq4Sq28gsyDJZgNds7qbpMsPKn579rr8lddE9hn28PLu5Ev4sJqF14/
/VBgR2rA5Paqi87WEDhjxfstHoSE9GDNLkdFjUUTvp0ERB28ERLLoMRLdHVlKINC
99zecHCrd8lGRr16XpfgDOmxRADlehVrDJV521925P7jWpHnlSPjQub9Wo/9B4G9
4YCSNcX6e4UZuuR+9x8WFPmMlAa4yslqfH4i38/XrZ+zWchO3nB2euLiLvkS23tQ
os3s9eMwMAm1Sd3fToLrNQiNn0zIB1rGqHxQ1YHXNgP6hWFz2BGgbi+drjeS7hcA
eFc/IPTe0xCKOlTrlJ3Xo6XXqEiEX8gmBsmzXCdnA1XIfS0goMtOpZsguer9dk7Z
CFfm1auv89Usw/9LgARCzXYXWCa7Q1fY68sZCAR9z/B0Rq+gHdOHpA6JQzqBual3
0HmmPLaYEqBiUnyGezchdDxDo/dkbbDTnR726QFKAV1BTy2im/GXo2a9uGVqR72t
VW5s3ZGYR1S+UCAhE3xQyrnXWw5wfNxiZW9KbKWhmLsJOBw7sNvjvA90b8UUnY/Y
K3okbHskD8UDj7ifGs5oUjns0hcElbnd7GgMXxMZ0cjT9UCxGHhqun1Q7daoGsvO
U17Q2Qq+qgHckJew/RWQrwenQPX6qfDbueN7/5EZJ+ipztFoOi0lqBh/Ii4Tc13U
m+QdQDkgAY/U2uQoNQDpNM8U8DAx26Dri+ZA47Frtvrr4VRNkV0i0sgRopDqtHF+
gathRwELkhnCVjgHhKiOdnmYvakcg82QNsv+wTpCbEf4aAsI152ecfxUc4Qy8nY+
cOOSC9LAtRsJVfqT29kH0HA14hsrQg7U/K0a2ig+sBNQOLwE2hiqUWK1uEX4h6nd
Y+KaZUDfPwyjfHBb86Ql2VjyNy4XgClNeM2bbAYw9cvdXcoIddz7aH1oDtYrOi2U
KipXo9+8SMOX8b/LLq91PvZwrR5poWCUdPFqhkjUkSYW1Tf14TZqFiM4BS1E8dEI
8IxabBvylWKpe3mf57LvMlbBjixWl/C69Fb5Az5uNpAZ7eiTEaF3xpxPfDIgyAXO
x6kE8FknmPVVxc4fOD1QzkDY/uHiTCkku1xuNyJYnK84aGXHxUpZOt/bIee24tHw
WwY9NPY9yrHRTSbeDYDqP5nHKS/uq2JMKLKTCgcLpwOX24eVSQWGhvNv9QV1ScVT
lZRmf41r7TVnomqyqlAuHqqDo5VxBAZ+izKbiuU8IJzHhNl8937uRxy/8QHgWYyD
CbAmmvtFp7WoBTbH40RMXySpRDQF62rqhtC1cT8myQt7uX1E3Fg06B/7f2avcO1D
4AumQ5XgHYxs8OrpxB7mHuFTuul4qICzIZR2EpKfmkxnKl9zIRq/MrwryfEfwNvN
Zx0c6AeiCou7MY1iYSAcNYQcgqpIXIK5VHEN5Jfc8Bdact683TxOMRhdnksd7lsB
U7y6jsYIQhBBxCLcyuTz1Lov5WXfd1sba9/IRrF1GVpL7VKi+wi0BVGVblQSBafa
FtQiDBT5atZENzsQa513PT8nVUzfW/3gppJpghGylWeEjXxci/4huLPZJA6VG3cJ
AqZRl/gadkK9MN87po+fuf1Tf/cCC+StXKOXGFilIXG4mg47YeKVjs/O8rbAT8JI
00atAmxnWnpgldmMfkm+hbftsp/HnnikWBJDhBfsvVC+Gkjl62Z7IYibenOF5ObP
xGPQECUFZO/u0fRGnG+ueTPgAk/1NEgjIbVOaENiZmS42iCVu8F/awicJx2X6Z5V
eVDiGDn61sKCqdiw6+bGSPFiVDmvJ2xHLONZ7hw18niWc2GxVeigSxBvL7wOFi2l
ZivVx/BgR9jgvSEbc66ZM1XumM8bByfR4KNXE8KmZ8DV6ypPLGmcC+0KJhVBg1CJ
gvXh6DJ8X1pM7gJwKqX1xlna1Yl0WKyE1ZT6VlaZEVjBaiQlOesipWUzmnErks1K
37VAg6OuuTvRNda7YoLeCyzKXlmL6XX2iJNYeWdxntXNIw2PZ3OC388OJXgcIWiS
oVsdayOWoexuCklIgjQSsfYlF9gK+5NM9ULraPClxf0RRh9/SvUpT04JrqS+XKBK
/EsmI31g9yildTK+VW66+V5Q67vuddrnA8HTJXvIBMX7zv2S6wWhGxwy0gL+o/TI
NafotZnY/tBGGK95aeTwV2ux6LBBtfuMbf0mSwPU5zq3BJVnB19OnfuNd+cQh6IB
vcXyAmCWXHRHjxoPM9OvyqUaWgjYtgjQA3wWqR5eynCHM/UzvaYXb8UXsfi0bQyN
FzTt7B4hlfC1TW6qK8o4ydb0ImhV4LUOLojXhLHu7uAS21mWtcW0J1Ve5QQQHhPe
2etjGhPFM7qNLLWR2ZTfqyFG2mAs8n4knyGtOpEzG8+Fdfy8/3BsjfOqK7JhDWDb
Xn9I6dqryEChl0paeQT6qOUPD1CFLXLvLgR5g6HzDYx6ul+6IYOVT5XBfRGNVmS2
BLhV/7J7ELQNizdgA7efQafKWSJhY6kRW+tkb4zXYX18bQlQOOEOYRbD0HKpWYMV
QnJz07HW1iZM7mhUMRfJzMImxYUcJuCWzW9DA4/M1H6GccCqU2yXdJp0leLxdNJb
Drf3Ps8EM8SbPEc2WpoX8vI1TISYSYgPzH7FjT5TimetUD1YbAtuUcWj5LNig+9O
2vVdkBlkpTQx1X4Z1jO/vBNXvPlDV5grBO7kh4GT/bu6Djc+gE5iT+I+c71VYjlc
AunyB0gAH3ESgyxN1ci2YmcgooAHvSoGIJL2RHCV32nK/xIftdov24s9+C44xc5U
z/UTEzQkmBtcqkn8rF6NXePcq/QFPdTEgXJD/FS70hFS5sVm5rUlinIDziJgxtK7
gEBaJd7TUUzeSMra1knmqkxVbw3Tn9s75Neuk1hsURBberuikbqNYyfEfaK5udDK
gK2cT+iq3SUlcHM9SWLAgz+6axUlErPpVTZ/kGmQq2FNEzRjgaL6xNok509H4ccs
p8bIn1wuC2nwU2Yq+QS9DPn4e1z6grq7wsBmnt4FOp5x1ICOelEVkM+Ii4RjUmLp
HWk8ttnjVelmlWV5R+2T5YsjMOfU0IkOhlFId6+SIqjzt5Y+zfiN1l6lKWLImIE6
A4ohe0G90SQMvSq+yNP9M2nvlPRcuodziMe41aADCRlCiACkI7xAKRVTNoyFQvFD
p8sKOTVUk4wB7UtARiwgXj1sGbgoKS0ji5VbP8I9O8Etpj/EYIhQhZXGrLLJS+IZ
y5HaltRoiqE06ivEzWlirQNEFOYvR82d3Xo76qgJioALJJHlJHBfjs8p36BmZnfN
x68palWzd0p2aDHXnxkxCjSacyWNjkQRIHxkEiYiTD7JwNRpX9S4mFtkbDUO3uaI
XNqMMoHpK7/YYNrTkumOOfqGM1Pizxmm8/jiCdDDAhadILsVMGonQ+wI9NEn4/0I
wiabQz7M6jBCdOfckeVfkvFi1f4vIlIx3jjrvpR5Naj9tTDmHNexzM6O6goTK6sH
AR4rSsYK8BzgQpG3wyYW2cgEcGQJB80rPXYgVXxAHNNz5vjtTsNwW2QhI7yGyofR
/pzZ7a2kMiD4awiLZZiRNuSpl+kVxyARHw0UBGkYhKrNwTqsi+7WJQm15vyAhDuA
HSrA1VPE7rFY/Hk7doBKPYQyQ4vAMD+z4W5+HCHV9YYVeX5zVVzsxLurvFQaHjlt
VY39nxpMDzN1WPVFO86j2GEtWyLl11e3nKbIitFKKsP4Mk4ZsM27siEhw54Ix8Jk
utp6taJXcUcXuz9Gk8G0r/vlP+owSXxFzU6TBEni2mvcYxOiaKNL5y1wpN4b9RMu
w0rE7zpSHMwVj/QiaF29jWWUCo4AMfDRkzJkOeOHlNGw8Ip2JRsFVFnMAzkSBIwV
mxTSwMrsz47gDXO/Jqri30+MKYO1EVeWEZLmX6V9wzibmavX06+9e97wurYBFJvj
UiAIkSlABQ3ePlWLrXGV+5PysxZ3bdcEhFk6RXzaLqrjPYkCW/pas3F59JxVlTI6
rlxoFdeCANG//y34k50L5Vnkqar7MiCweErY8ZhmhpmcV71LjZMb19JKmpOtTCzw
+laNHeJpyrusZq6VPEEprrQXmsEcqh3pgy7JybdfD2Ah2VREz7V05rMCzzsvWN7+
iepbQusvkszPKcpYWscnErHmf4BxtMDvTd+UJjDUOG7maG8YAy67dN67Xt3iM5xj
FwfT47GTWt0ZD9/SFWxaxB+zZZXsUuZVIuMExisoWO2sUdUyfsTAq6dHIiOoKFEk
RaXftjZLuRow35B0Y2VPuS/209wlDon3VEihuXfA079P6Jgv6nHGjOtF5qmdievp
DXMx1A239BGnZ34OxdfWeT3rQaup7svvgzyFs9H0rcXEFHtoMAzl5+X4naaFZKq3
JvaZmAFYKOW1GaxMnjj/p/5idZyYJ9PN6KqsCr+8RRNpHhllBOcJ4IxO6iluQGxA
Sqmy2GMP/WcQQ9IlddFZwx0ZlzAmU155Pw9T3jQSwDmEyiqd4NEUOAJrzI5jiwUq
eUzEFgjABHeeT2KsVOa96erhpjMD3lGC4XURxflaxFMhChGSUF5GoA9ZOuqoKIb9
qIy2z8TdxkJQtnQHqXhCzWVdKe9DclzXuiSsFS7iDtfA705WA4u/usrCIprYOmfZ
sATsx7cg5zsZizDfCqxoQheNxbo0jnF6mBwbHX5R1/HWXgm0ktjnOJ3/8VzK9urB
iCOG6mwHKVr4A/kkeGN9bvkBytjq1uJC0ittSmbojPtP1+vdtsIt7eAv77Tk3coI
HGr1FkCL91PLHbUz9doI6f8uUB+fo1k6wGcJoo8U3bEyfwG1JtbCg+Qcxlf4qV8O
7mO1Fl6QiPo2dGg+DzjaD/xOxVPI2Q6HyaRknweubPcdr3nPNjEbQ/S8ityX7Zy/
Vn9Z4jOLct6MnmtAqsd+Jit+rcllfA+ihW9y11SwRE080W641n4AeLGwNVoSAmg6
tylZttZpYXcG6oQP/pbAYsE30+kOAno1r8/FMqTEQJENI1aTpaAxoGSmKR9h05p/
DWCG1gTRpONTn0SMFfjQy41/umLwb1PyY2PZQzCLWiOes/3iYpYhga81SUVcucwc
zvJKo57sIpiJmo0ILZAmzvyOHPqYsdKnvQtA9+7VLmVkA7B/ejygTWfYYPe/9RTZ
a5s5FPBku6/8B1Qjj4S/Bq8lwRsR1LiPr257a/bqlKLivIY/8l2ASfaW72NRBtJW
jW9Z3SQ/J6Oc2VddlMe/1x0Xv2gmBUFHAVFip8fqHpmkUkKZzegdOWFHWgt3M2M8
mlIDrSO0W9pfoq9xm0qFRJWx013o3V0gCpOiquOyHxVLhkhOxkWPDqT5Wb7lTov9
LloK+fM/RYd6PajvbAnu4boeHucyVgsLvMX//zm29hHLPZQRwCJOwjtF9N71lS7e
XIhLqsh020Ix5HmclAUzXO2YXoSQjPI4F2U60x6HFE8PyCzWsGBZ3F6Oj8nSlNn7
ZNlPRBTIh6teUq75k1Cov1leoUdC+Hf/PUlxT1qclvI+T4sbbgnep/GZUOklOItH
FEBf1RX5eF2EOXtgvnTiCh04H87Nlre99TFyU0vEg0I7HGq+kqGakB63ap/Vlb6q
wFYoHD/793Z4juWH9Pr2+BK7/tTCikQfKnFtG8DSZT9qpJHsqBrpn8Qc1Kr05Ak+
b8wgjzrJYjNK32iMb6fy2/mr8FF6I5Mqw4C0+unUrNOLoTot6wYRDzHZOcqZ7SC/
dB06EiZpKW8xIRErWA2mD7Gl6DPK1jvxHBIWyh0A/QXNsLuoLgq64keNMu9ILKaK
8r3ahHLOxjSlWw3EAlDBuqRi7h9u+aiwu6yJrxGfYC6CHz/57c5torgnHNOPVgnJ
ZVqU1Y1/c6f2pghXP8I+er54A1WAiw0YYIQOwfAcfOeOh5Y0SHSwpY7Xp+edS603
UW4BRamVmx0hunz/AnQbI2Xraxud0hLDHb/7HkMT9cjXSBpjqcvb2eQHE0Ci+lzF
nlqsi9TOBbypMu9LyWw8i2NMwnJP4GHUdd3o6EEzkF0wvvQi0jnfjx77SXw9w/kP
fNwaHIBigs12l8gl9aNnI7jbG1OIvmeYWphBdpXs+ub18EPCOWn8xuRsQgSTpmaZ
ofJvRuMYXtNdpiwCbtLlrKvdHVO9K5IWmPlUyAhp7mghp1aDfNuCO0J6ZuE+3xvv
Yo6mbqyJV7hfAr8qRGZCE40AJKHt4nF8y1hrbES84LwykD6sWi+dTey3fkTTa4yO
iFbJxjAjpW0Vrfq1Zjswx8QV8Z/dMW+PqxebccON6FfLxTFoyh3D7+/r0cJFKDtT
jBkAs7xGtxfJCiVwGHmNL7PYccplUonUhriBjOypM+XFm7psSVDgF8QnoEf6HTBx
zcyfhAgeQB4PpsFNB07juxGkl3fadjaVm4NXusPD7VRvva+4Nur0DCyHCZ7B2Z2T
UoRy6OIpOMylPBIpXV7D4MxG75BGxAeC5e+vC0CLE4jQUt0aUsjuD/+cefwXX4N5
U1ct9Pw2n6OrZOqdfYkeIROzHYabKQYTrB3WVmlnlittrRVCZmAvCt20Sir2RpdM
tQBMgQE+OfPoMJYlmXOrm9sjsCeBGS2X7iy3Ypds0PYm42NJGH7C/a7JhG8my/af
L/Ty226qzNLBtMnBZ+p+Y5NkwNXI2mrIWyT5Z+3wjrRRp9dsJLUlvhQGQ0hRDhKr
Sv8XsY2satP0U0C3OPY3O+kOSzUPd+iUZQ1NvtR9EpFFatP7uMeWv/GjcLOdIsQ6
iQPL6vj7UPwW9rN9IU3nm+mcqXUpMDt3/RRwk0/L0UjvOiUtB1KO1vZ7QIblM75K
bXEn+BhO8pYnY7lXSvNNaI5/nPDurj5ORo3lG8ZY6U9+Rj8ShLDGOYkvi5Lu6qLF
/Fek1RXCJf8D5aMXiQnzEXpqY4TWA7bPuv6V4FtGrjjXlVnY4Z1Tkq4a4wWPzd9z
gz0adIF+FnFUl/GFoVFsrLuIjTmPBlryadwFThRszj/smMossPcMYh40/aNrzZBu
izoK4GjWy3jpGMK5e0EgPjEWd1kIQFQRds/uWcLKYjd9o5C3zHkMIGEfUYAZINF+
/Kv28lKi5PbzDTm12sDm1ooiT+GK0ifpsoF/TPWt6rAZXz7YcbBxBTa/muGvFqZj
nsXcG4aIvhC+7T6AX8L1Jwk/qu5o542+QuV/pp4UYoKJYwU5nSM58fdzrHlDrKzx
pM+MjHWqGlmxsHEz/fhI4SHoHsqBYnxi+V7OdNuQqt+5VS0s3oBMVcg6gXF+mxrQ
eSEKug/zORnMNmt95f7DhBYeTwJmFUnyzE0GISXVxevB/PFOZtyHyzSVxTjX5Ska
fDqpp94d6UeqdfQHN9lz07zP9EI9e+8tN06Qs5OwSna8e7EqeGby9OueTfxhoKR1
e/RHfvuy68Wiph+3LjnkVu/epuxnqzAfnN5GjA0FG2pOKAtMCr7KqIKL6dMcTNw/
MTwYFeVp6lIRRvlXcOIWwYAXkyazbwx/A9j91y7bGkYpqVIDTnf545bnN9N9N/Oz
Xqvml7oV0tSdgJ+fMt/cXVwdd9/k5TCaQo1MpgzE7GeaFAtvT3AScmjbsL8ywO8E
9eeO1PI6YtLtirIgsp7xmU0Zd96JLXmbwGeLluoXi6BhKZCycf35T5vHddyu7P0m
vy1oSdDDBzi9qorSq2uMx+BJn+yf9d9SjvcJ1XiqNT1R6aEqoIksph/AwfjqNZFN
5bXxY4hlfCIFw0CxlDoB1ahVU5sFpag94AKD4LVlN/OZwngLq+NevYez7HME7Wzu
AGzgfuC64XNEjQSIBhh1jpw4peh2gp2HVCWX3DDzwQ2joILjRwaOHPSyTdO0L6Dh
XRQzJwNTMGJK2GPam2LVxjY7l3GIKhBU/1IVBd2YvMhLAR3xAAuYiOyRu4/BA6xm
3ZCaW6t7MGROYdQqKLFf9w88827XRo/7NKVdtsCZw6GtgtqqBw3NsX+qQdIru6m9
0sd14zuWmhbsAHVBZsu7AESBfLEbDqRoF4j/Yad/0fAuhtiLF7CbfLS4Ql0cvJvZ
s0/5i8C19vuxZKrtgHLWucfCbGfc+DwUagX7mTPJi5fpOgpPwPq88cCXYfEnoAmc
AjbX3zD9eXtHwAqwOkJgLKbQXZQrHJp+V8lRqoRO2kIGVlfDOVjbshWYhQwks266
WvjmRLO1vKhVCaTI/OUC3wwi4TSGCBYHXI5hMQJ9VINrYY8204XlaNj+aYK2TUyl
Smy0ffeslLplb20m1RdehrgqtWWZnUyhSV1Q1JwiHz3mftl1nzFEGssc+wD2FZi7
QvmTlSsjAMUlCFrHzXA4OFW1nejSvL1SvWS7IWBiEndFqGUyAtzmdAl2hw6vlsZY
9dtNL2wtl7FFax4BeGKedWc9MCFJ8IKlGTGR6mPvxvHQO5YKcfE91shb4c1lZwkn
LD7yAv0oh5nK89fFM5ZuKazQizQBqaClZ2gTV34r8J+tQvxhHlrukMWxXLbrH9Ng
vbGrWanWiXFnGJaBjBLwgg8tS9mH3oszoVwSC4NkPjuAXnd9HVZfyOc+qKrOozTa
va2FXxFHCHGhbgSyLxuZvDr1Du2AeILLTZH/14qluPF8m1Cj7r9TKpRnDSxWrlhY
/Asj+KmGbQ3zYVCVs54seZzN57ESVTxJbxWlC95hTdOk2jP+CoVb2PvxDo5phP0+
XtBAUsUETKBY07o0uONHolCKtn/zcbRRUbYQdt6hQSFlzHChQ6uTdoTgKbguwEB/
uOGKvCDP5qQjpnICZJ2ozFI6FsCROgHH8zwtsH1W6Md3pbdDgdBjW13BVZz/i/z+
Z8Oq/2lsUu39haVjL/8TiencLityXpW7BPw/9aGso8oOh+eWtFT8XJDTCVYd/yOf
oXdCzA+7S7L5DnqMnlyoFdWgY9jAOdWiU9ayN67JqFNPzLexBfC+4g16kqKXXA0I
Dd1qARDtkMDlxBj8v+tHLIJboWUJs2kqS0zkZ3TZGbOPoW5BrZSUFASaE1ogFW50
1d0TIoHlLzlNT4EZa3nMxSOn9dS1mh4xoh5263EftaWvyrh2WqU61tTwueVzI25S
joDSt0tgA6tJndmXQjZhFSq2kvKi27tkz/7/pV9+WswW0HGOEtuoxPLjI53qvdWa
hoPfVufxFk5PMyb3rvwOym8facqiVyoB6KkQM2929rvE/dVOZMfEvVgDTqN5oUTh
q+zvmM/svddojcYBmvDqwltMCfZMYmRRX1TdmXZoYMPJfMCpgALX4JBb5XqxpqVK
AJBMyUmO/3Ahe8jhcCsBko84fDadUVTd7Kp8RBhIaurn4WwNoZeJyc9chJB76pNo
m9AepA5Htz8mYGnEtpedr36DuzJ1YxOwzqw8Qjl7wn00jIuk87K+YmsaFBYZEnJq
T//4GU+Xse9aACYTChyf5BrGYcCk+PvI+2hwhsvV4dWSCJFuTAeOzcZDcVs91cdK
3JAVUYpr2bmdt2WDq2DlKc05LXXPVAXJ7xUlm6Df8dHsz+we4twAnrTBJ0d0wKYN
rr8jqsJJaTRyfxYeLc6OG8AaDWF7Zx9I3dsgdhcTLK43AbL7PQ4dl+XOCUHO0WW/
L7lhFQdRmAeOdAx76lbVsBYMCdN8DSYSjCOe6lzCnH7hFQyqkm3mnu5HRSqTSwUS
Hp/+FmL0iHEesRJqo71WsBazSxjyc/idPvOae9eYiE6ZAlI0wwNHgAM01VSEscm8
OQLQpQMq+71FSW2oDojv22Td5UbdjwWJS1jkXMa/Uf04uaxOifrvRMGj2P8z8XKV
GJq7peqbw1j2k7nxcYI7/AyzBQht+EMKlAvRZKqZv8AVDDZ/q1P3/uzXLpc8svTw
unD7eaCCipi61Hq8pfWFoC5ijoz7wI/TckuA8qfhaP/UxUmQnBpkX9ctZ94ZFVIY
0Hj7lIMt9Ts9MNPwsIJkz1APchff01/6ZPMVsM5hKZ+Y1zgERy5Hd2YkkKZ96FnY
V2YEfIpQfU2uzAoHN5bTrKEsA+axasFf+8gUXRQHqSxYTogEZFbHcVVjDH0TxPFX
/DnhjKDtPiKU+d9QP75+9nPMhuHrq94GzLB5lqgW+xA/nMqZyuYn1aS8QL8Pd99S
JEXJYObdoTQxzoZ5GH1oejIhgF+M/bQSucDcjXu2i3AA2XbEBomG8fiOLt3G6GKb
D0JgrCqToOjmrXcDJWWbWGtHIVpsrJxwOl8sLHnOWbwFfvVsTPjNDc6zAteOP6ol
pp4YFsYJF9rrmpkGR4qwupugbKxg3cIq5CkU+G3LkyRlQx9jJLcgWIdf0m6tktWm
W14i1M/rPrCGfcixtRSa1AMra3pPero+L1S1UrJSVobbv5yVgBcC2TizvJq81HZU
4CkckU+stzSX2Q2sq5r6tAENz+Mm0UDwdVn86LSs/zl+FJqlDTgCMPAcJZs+WiPo
/3W038RRaYdCO0QcmlmtQYekzpVjuRrouU2Nbe3wFFgROV6TNVOujd4hu7pAHjGR
5xORs9RgkXfpsB5vkfijm36b6eVoC4UEX7YmWgqY0poiRgYJYeZquIvPz8iIFFDJ
oG+vZqQJ9SefOb2jRKKvfza9byL1kTPVTnNESTZgpCnBOQEF54IVu16+9vaVEUEB
mzVgsBTWmslbKQ39mMOOLZroEmbdYkeuVU5T73o5HIbEp0FgEwIYfIMNhovqdz1g
UdytKjDBfhHVwfa7HHDTc0+sDF+4rntDDQ/LRDX7df6yfBTrKigKBrRVfsCIR1r5
g6PXOR5Chgr1GwuQw2jqnwrLX4nqckws1xb3+aSJuCk6GKNtbED2DD6mJ6jWU7Sc
wCMbbp0HLrWW5Ch4uryFuQbrmChyrb2sL5aGNgWC1duO/QFBgDkYegU34aAYi/wr
FSYMEcmmtJ78Fl+aGjzh5qI203NAnG3UJVlQDpyCjLJE79Eg89LfIUnV/l4NqEEN
K3v0mBsQg0jPTZoFDloU5dgQz6ezeJrB6rj/upAf+iBBHEO+qsbD1T+Fs/7ha2KP
QWkfUxkLwfDhkJ7eltrWW1nDEhyoDKO6w9XRUF3fdhkxynlF19R3f0EHgydQfMXv
Z67V99NL7PfpHB+9om0mPRqw3CHQiy2zSdSEzGv014P+BOAQm/q+6vEXKoIZ2+Zk
R1qLySBCBatLNtPI3hrdVbqypQqZlIGivD+imGafD113KKsrctvMSKdpw+1ozQ5N
RPx2VKu3CxyccTN5sDA2F88UnQipewyx3XFdFhbD1TVN2HpCAZ1uIb63ouvmkvQ2
uPnmz9cZgNVR7oKm20I+zzvSc071YFoRgFdbMOOkNB0q7MFu/dQ4l8+tHdBpVLPu
UReCi4Mmtb0gvahjZJrFqInuUsKUpWewGV8qinxdbWARs6nJ8/lO8bRJpGpYiiUi
r0Ax5G2IWz8HcnFvSTyMWmkHu4NUYB8b+aQHTR42Yiw4L4ZGqSCvFqmUma1hOhA6
UPSQQOZbL1uQE/6PchkEFoiheYD1hAZ4SfK6yz3++izIyinXzO2B5wsRNQk//hlR
nWl6Oqo5kBxy/Jc4Ya77U7HTFGHdUbm9R/DN8yTzMqDPF1aJpryv1BjEW5GbFUFA
zIcI/IwVcU3U+7nhSYNdh5oyQUu5717Lh55DOVLtcn8Iwdq6afPwkW2+Z8iZCNnB
B93bfl6wBvnj5TzGp+7xGsE/R3o/RgpjeLkUTPEj087vpXe4glnkVvu2HOJdWpLQ
SDjzINo+Ljy+jrr4Di9HYLP7uBYmffM5S/MI1teKirCMqxedvrbE7GZ688+Fxyjt
bJ5zQvD0QdnAhcMhycfyD1gsWokXR2Tik0PRVC14nMTTyLjo1HtISODHyUK0IaZS
oYGDaUUtTj71ka+IIT3302ZjerS0cbgUnnwivsXWD80d7BHOqDM1celXrmvBlz5L
QeKWKzDWldHFBVy6HAWidhk/+lRd1Pizs53P097eyEKc7bY31HWxjDJOUB6Dkd+g
UfpA0TBggqLSO+ET0zMbgMFaxWArdW2zoNapWhWZXkbmsBsU1bXMPwWHdulpbx7W
j4/tQmFwZZsqiv06ZXS4DXrd4VWR7tDVWZfPIrO9oOYH1Skog5+YDB0PWog2pYUn
4gJy/hM5Vq8Ueyo967f0ub6e8D9ldNQuzxizKh7FDZ6Xy8J6PnncX0GBxrwU9i8i
pOCbc9OK8DRWmJK7SAR6LmCkWOZcIM+Gc/jS0FfjJjoCjDLOcSrY/A8yqTy17qh/
MHu6Bfv8bA1uMY5Jag8Eb2ma504QBrt+3I3Jxl/7MLJk+9Igm30gtl74+rvtuGR5
v7RTawuABOHl/lpm2j1YEKwaRdjdG5mV7RgY2p2P66SrvoxU85vfkkKH1Aan7cfB
fEz45HdoB5S4p1eOEH3NCDejtcvsNo+HQkc9B53wSBrzobb76hv9a8K0LD7I+O+k
hkIVXbCu/ulVA1ijLzj7zQBb85It/ORxy+FlsMTMtUYclZ3kpmW+ux6d2ieRBjep
xhIY/xm0XzRxfZ/AvtYAuOFn/OORFrM5i+8fb5Z+bu8WRkRpyZGuE3VCNUeeKTQx
rZV5UxNbOqMrbPm6qhEnk8kR/4EeXxdczdB3DOjxiZzhUNRLbtU4pGMTqyuovdvD
pu7oRofNuuhF67QLmPKBg+etp7oZM08Fb0sTf+iGXdwNQzq+Tdu9HRibkaf7w/mk
NzkqJEQYXLvhbzbW8B9833u6JhLjHVvqqecNzoTQwHIA/YzsrDTCzu/AiJ2GfWfk
cTHdpa8ejpzfegnHxiYsBBpcTP2j0/xkiSE97rU5gWe1LfUgPl9+qujs4goQ8ckB
FN3hn/1VSYp0t3Z5Pzt3Zufy3xzylAxezSdNM7dhs3CAnYlqtrZdmxc4T8UQbJGP
5ipErOX93bCKYL82/C88K2GYhB8thYOL0Hh7D4Idnu5oH/jPB9qJBYvwFcScYwmA
fdXhZHsMaeAw2MtkfWTJNJKu21tOpNykPiLlfzaqqKdMvMbuuS7HnWoqvkKI+1ZI
noJ2qnMn8MUm22Z9Iue5SqNTyZvzl+VaO3mxYcxsZm7jIkIcXq11RYPPQm58iafU
rP0+Dh8SebSrWnwSt5L0EZGoGlUu4oEnTVSO9w1zFeN+zzjwp1j3EmISHO2iYvkd
4neD/cSjQBo2UHF26FkbH4LJLXXNla8e8r92jbUrKwH1MsFYeK34YDsfeihAZSi2
3dPZS8ugluE/xvVAAurP1vzW0FpGu98UmY+mbMoL+yKWOjoj1sZllSK2aOiIxYnC
CD106WRLYcg0y9V58GPTi2OYbGHSqvFJQUIdkFxiscoOmi90Ec1j05t4Lse+qDbj
gDqP+n0GLq1vAMPDWXDqfbX/eeR/VNv5o/qRbKRkQW6923wTmda4gbdi0KHs0DdS
IjiqZ0aI1Vo76HeiHbdSSA4F9+MXPcAPekUt0Q8S8Cp3Qp+0n2jLZ3q3ekoHYbBJ
9a3Xqd0n1HKgRP/yNdKSWSycbbHf7Ptg/pzo/meNVCuJ66fdTqDjFOOfV4YF2lYw
wXGeyrZ4dK2EwXrXgWgw0qdid5Jp+0hQ4RvZdlVk0ODiQuKkAqFKk1YN3QWELd4Z
Z0OG+k+6ODC/rNxeEz/DCfV7Vrd0GkhgvrvkNeHobNg86cxtATGhIRJTZDmEq4HK
4AE8xceDuKc1UN0XbHj7zNelvQYHINIBbn1a9ONN8Qdl6ivNVGm3E25DU2zhy+xh
c3HRvBSVkY5GRaTbyVUdEBSZ4o6fhst4D+zLQfCgzWFNK+J5Ce0xU8ZF+2SG57UQ
D4K4nw82BXbiGTMlFaIINVLov9wZOfHda2DlC7pfyuPDBR/JPMJeffc+PE0VWB2Q
rVARDAl07az9yOAo6jck0KKNzm4LeCQgoH5PeiTCYoVR7/QZW+eaU58fdNbyhXYO
emToKFkJp/V7GfOhlqwMaT/7eWO/ryDodzOagkCyf9h5G+LgZ/FpLujacg5rjMs4
Np8miJuwPRvXuhPgIC6WqyWPgTJdsaw3eQ1VAS6kBYZGS0nPPbaeRHz36kfwVrPm
nBdT7t+2iQRiwV7s/AFtQqWrsYZTAbn5mdnOg1+E4obRMLWXgnTrFSzd7wlOQe2G
RHZtqnWbV938e26EYaGwHJqmUu55op+EQ9Rp0b4DvE/Ow0jEZfqOCwBeWXM7Gjuy
b8b3/ggmFg4u4F96wQItRpR7zMBMfMDFqWxs3jzmR8b4t9NMsdxgt6yw5DErMM2K
mfGqNg86CwAqigp5s8KWXwOda5q6uEr+8PBG0MMMD6V6vKsR7Uqf34l2KB1pCMsz
XgvdBfNx/nzchHvOFy4SqyOZDsdyfvB8teT0L9lqRcJ7ZpBpUpN7PMPu1mCEkxSB
c4pqgcisci91Fq3CaLH5/6JbvbN4XjgrO4vaEI5FbWnCQExqzkwbqzZ1Pq3CR7Sb
9+GNj/ZpLEM+NZp6cORUHIconR53fbY/8/b8KpTpW/fldcx2zSNtVpwPvqVRD+nB
Y6w2wHr+WGnvIecb4d2KMfjYL3PJFcRrXlYewI3Wt9GpeovA4LHB5xoaBfym+r3j
SFD/4l7SpM1eIXVouTk3IxF/T28ALpayGxiQePeC6QnDfIiUH62DFZAqrRt0xjVv
zUle21IaBaa7l3h1wBq8+5rI6kppoZd1PdaAoFzG/q1JGvoF4gaVm8mXxNf5prSa
C6sIrcf6QdgVrqSD9o0CCuFRR4Ob0CyjqnsIDtqd87E+L+99/HFv/dUumXPxN1Db
ROSkuKMvL4J4B9sXMuwLokqEl2xnTi1/FvAwTd2W8yVA3NkWDLg4sWH5KVI7n/FZ
33Dum46SrqIWALtV8WxkLssyWv29CgoZbvoReqvR96wEGaQLCvDkiwX07vm0rPod
LZzI2Rdk95Hv2B2J7YHrJ5Wq/wm3KP+eb3CnAy7q7RJo4E66q6YTpfwgs/dtcrHd
WmsSW/uk1IEiazqkH6Asrd4wvqO+gtlttolEQaLwbLEB35EdrKRnT578T6ZQ1qnk
lmjoaEwdYSJwYbhReQDbf47oWWKFQgJt83NtJTnPjq3ZdGrP3EbU0yxrfWpQ4LiD
0I8EVqNS0II0WOPPSMcPqsHwitdKyVDqkjzmIaqON74/ZmoiIvzv15pkjkWlsuaF
66epjDCEwhzfdd0P5u/Kh4BEuP2Mp8uxP76MvBov1QH2DqbwevipZ3NtQ8akb4+I
bpdhbqqy8vG9bGuC9bywvbWSAMR20goUz2XWfaf1sfrAwXyfIzGqTfPuPS/Ki3Cp
aHYyhBV8b/YWUGK3l1ekmhqI/9jGmNhtfCbXEI0hfp+K47SHG7kQyftWN3n5zlHG
unXs2WeynrcBzBBaazsgfw0/b9PP5r4Gq8tTDW0coDVYs8qvWvLAea+HGOEvfHsq
NsFn9GBUI3dS8JnWO3rT9skqg4ADtxHIjDc52aBa9l7wvRgyRn/sMnDtD77xSDVq
42lHyV4ZjKMY+j+uixvOc5EO3iKu1K75R5oh9j/s150Zx372SYg4bDI3klOhBiew
oyobrjpVKfwqKmtnu3fTlbvjoeZE4NViGIrjEyVdfLx7XIvjosyM2m9jMQvfs1AI
z+Wo+cCeAXhDIRlFkWaSgkTXWfYSz4TozoWZEr4fBCx3mbSohOruYrMyVhAmhSmF
Hh1Z/D2/wNM5A0KFuv1U+NYExa0RF9+ru4TbhFAjiy35BjT/swRCC+DgwJNyoxW5
1b4jOpRW/HvpUfK3rSIRk/NHs9bpRLdXQyZ4fJ62eL2ZiHtKhZlJkJQgXqfYhaw6
l1KmiwWICLbhvN+gzQcdXH3eJCsnCKTaKDsHl+i2Hvk+2F/GmCHk+AZlLnnlsjXD
reaBhJ4SH4Vl+0+dTIG9Okw+jlQ9OvJ+uDUlP1AexjiW2SAoPuQjExVc0QRRh7k9
MgowRReNPAbUQZ9P0Ufd2LZtKx7wW5ZAyJq91rnGajgsuLyWAhQbYdQqlWBy94ja
fJdDvTg0vYsqnfk3zRCofp4ZS079QMU+7iiDnW22eBSsruxgassvE1Te+vJ75Pu8
vIQJhKDYHkJ7gYxdRFC21PDsF+v8NLapVtFzxhs7GxNViCmfvt7py6n82/lPPFHc
5PjaK19eAeM6LG/IOYdovgTKyXnhM0Iybg7UcvjRwe1W+k0pi37ltZ+IAh/m7qWX
4+9LZRu5hVfLxbW5BcRhceO7HkbQugKBRsEFdWgudZ7LUpm8RyALhA0lL+Jar/2e
8Y7G8UOHSrLfUC1ZlGOPys4gtmGwSJ88jXXhxVLvLlcuVn2TxZuHmHmtIvSl5rlU
uFVOz96YfD0qFXY2YxNq7UBU5to9nyL5im5A1V1OBDIPM8mtpStSHZ8bEp55TSh8
GyLYYm14H5BiX8HZED2NjEflQYean+VCmwLeo/PNAJx3eipsARoKviiqrmvo2o7t
V/dYOe70uEinhd5Ne9I3eWl5gwzSIM0Z8hf8P0yjk5UJqQNN8W+Y6o/VqvgphokX
ldHW1CO6GyefBtztoE/TNtn9ypjaTmP9aDwsX9n+Ai9aFTkHtUJzhEMWy3ebB+Uk
ctKTFcwOevXWSahpCJWo8D5Edjgd7hKcUftC9f4vSgAOSTz/rAU+gCDYy7X4iAtu
3evbvzN4xt1laHcExtu1AhlKdl/u72YIToaAqU3Z2LYcGMdQzkNEXnzgfVZ4NFtf
4E+PVL8ls3497LdywSzbPGbEFVMB9JNKqtMarK7ilX6JgOcYwJHKztSe0peqYEUq
+oPDogj52s+EqCVOitBkk8dHFj2003vmdiwVwLiAaW9AzRtiDvnHN5W1PQbnWPuF
tro0vG8TpeZAz80pcxXE91nICZ4f0XxUxbDHC8laThVKuKSTzCN2sYHrHWRUfVym
HtsdBasT3wAdfaTmitsmOjNriBYTnpi6WSspcKhaBvXX+vLgHlU4VGzOyiMiTUZ9
dYhdRGxnTklI1F5kV8fbqwFirkQ/jOYWyx7FurttBrJlBWcQLi036Piml7BO3Fhu
OZXHi4+KeQhcK79GOiybF1d2E423RfFy0ZAoPk8ErFwYReXFRmaV9QGM4BJArj3I
fJRfX2T+JvUlytfZGKdJS83Wi+uKxEZzihfdGnMDf5BiGonRmmTuxoNYqlwm4Tds
BRR1eFxbuKfYok9tDx/1RWV6smhFvdEM8vpT8yWMZllHn5Ax1c9J03fgcSEVrxF1
S+Oo232ECrLneGrUwREEzs6vIgQfeV7iV/zEl1EogIgK9Wu7Y5Mx2s1uPebpyx0H
QdwkOmjbVfQC5Gx0YheOA7SgD8MnChXUSVXnkRdth4uYk59UkTLJzDmFkCcKGOgX
YWhJMoZcX3gb3LvA/a/cYCnu5gGaqmVaeFMSnzPVJABXwWgFO42ek0TcS/DjveAy
Q8DZWuQTxrze9vawEL9G+wMvhZOzJJ71f0Ru+g/N6bO6TvGwxA2eSfV8kZiGk/9R
sKGCa/76xkc4fFdHIVTEFQwz3VY1OfISL9QOgOWDxFnb2whO/ZlhJ5q4D0W/Y+6W
0jGktsr9j0GGV2EDLTn1xDWcuOtLS7rQ33HClPN2WBgHxc4evsIdoXp0M7hxPxp/
s36xjLmoYc164avdsGGhecyxNilzNNs3HxrMBp2eJMXnvVg+iQNWw7FiylFJP4cm
ei4uwDsZJzBtaQsxt5+FsF3UMuagpyHMSyKCVQCUmM/1mzWn/CP8w5b82/VU0PYY
YDvM9PnrNzUikso1YLSoIduHu6+OoSi8N30QP16zXeSD209tw9q/0zuMi+6gNGmv
sgsWeNOgYPqCmo1XXOJwmpsb0SP3Q5qZn0RfHth9QMxb8cS2RvO/BnqUB3gmIe4a
NjJm3Wp1sxJjf08K+RRTtFio34oN4xdiRVwwUJjDjfcLx9bTnLYR5wZOMf3HjVdg
qCWS2i8FXbczmqNHKi/Lqp1UuZiHKhfOmg7kzuxTvPJiMgPZzeJa0D5+Tp2nalOB
RzWn5jM8ibKyaty7+FFMa0vVQkEqPBm9k8flK5wFis4ka5az4ySZqecvVbqLfBzt
aol+d3E83iz25TGm1iWM6Tjjgm7PML8cM3JH/bpQQtK2pZt+2LJwai/TguJGJTRJ
baga8wmQJut0kDlDZ5FJl9e4vDMOCXQHXMMOXyqL9Cu4p6WzkbT8/p/iOcUi9h8E
eDyz0oqfjEz504xGo1OLXwmSLw9ldXGqD5P3Iim8G944u+b153mOUmS6Z+yHBEjG
YKgWknSnOllEeJU1t9IuxAvcf3jpAqdzxHg1f/O41je1DblfHMTY6npee+KWp+OE
62couKL5GONy5m4lEIEoEjHYVcmc8QpZ/l3yqcpYMPscavy6l0LGeTTBs8nlW3Tv
gSL4WpWuL/FSA2QLht4G5nOhf+2V5/+QFzFoEIPFqSej0AdLhy0dHPbbOQ2DZNK5
kRHsiDr0fbr5HIWENQH59cF64UI7eIJihkjdy94Nzj3imJMF4jr5HJ1M9xVOVCu7
2Eg4hX75BbT/Ih7Mn3XAqLUS09nUUXw7C/g4/xQZ0RF0MRAYXp8mVUy5xBJqlJHC
ebmmZnOppdzHmArJqmpOE1eBmiQZ8chuA+YFJpJKVmO1O6vQLW9U9vYL4PF06maQ
OGUtWYDMktPA2QEsLlpW0fIuoQ1Zf7p3O5q4XBV4tNYwt03c93A/1qSEghaXBuNa
2RoMHAUc/8XhRegYAiDBLJjg7D3YmR5rHY9NxGQV7GmYZpI0cAMQYiD5anafp1fn
uDGp7TDMD7RKDbK4SDp0cu1LleB74uKNb5qA9gDKPOlqPMj69YA1J3l/fGwS76Y0
ElDxYcTrDHG+hVN15GhO9/dbgQUiGzX2IwHvCMbgmQG9f/CnWltf0cxL6r7Ol97m
X1HebcUrm46fsq9VcFjwtMOwpN34qlFD5pgSqyzynsqkmiIZajSXLK4/GzTY5bnr
CJI1H/sRGcw0CD3YgB5DZdJIYHs+mwch5rcauXfEMaYwKbM5a5C6Z1d4+GCtNw1F
4SKRCDfyv6ovADDFXV1ujSkz+3WX/gbmrZMI7n43F0KRSSxvQnf46SNS2Hbx2ci/
BkOtkf9XE8ge78Aa2ZrXR+wTwZTlcvlbZ2z27LADie8RgJWAr4vrsCBqtFYYRKd5
mNfLTW++sRSffseqrf+IBciU2PwvQ3lnCKoM8qw1YeNHtw7VDAvpqGwjMCsYUaeZ
8g9fu/ZBkv1lbjf3wrObX0bpRNo4O3zM/ikHt8CTwbH5S+GG7Zo5rYIZ6rFDmS9l
AHgxZkepFgSg/RrDuDLgK5u9aDpsfwpr6UB0xuGqcwPpAyPZg2yH4DOfjQD/8zkx
ShCS264ePlanUu5j+CmA1+t2JllubV+6mSKEoRLefegsalX8ZhspsvNfccvGhDWm
sxUlmzOhTKH/yVHON/cIoYIyU+9AFpTvuO5Ha+k1wWaOV5YW/QWH+/pxL2NMVRfp
IAXMQ4R9AUrXEmzSONluyowe4KlDliJN7TEgrBxc4oK2kpl1DHdcXl8EFKCQTD3M
6yslYZwVi4F4Kcq6gT3YDYqcJwZXcPVBB53GCKF+jLTBjDDROGC44IZedZSjAEdo
D2XpdpU7eDfp0e3XGK44tJVaPoidzwFiLIDe6sfwd+m0KhJzLxDaZTbqEuGxGOzB
pvUoV3NPAZCvVgo/q60x+l5dEJaKi5i+UZqifXcRFD72s0hZC1niW4k8hD3I6Kdd
+Arx4iMrJkZwrzO+9zfQccjrwB1QubuGIpNuU+DGKFXXz84I5fhBkbUqLdwOqCjC
R2mBk/ioCR5ffrGvFEOmJfdZIWhOAZql3nIViV8zXPNaRJQndPwHfAKGs9ny74Yb
wRglOA/91Uw661zvhJ7lzCl/i3fnlko1MEr/GE/M5fbd2wet0DTRVUE/3pLTAXki
raZErkH2D0cek9E0KiA5qJVeGqsWDoa9KCHzlJzBe0QKTuusU5C8y1oCJmbB7tGF
p5YeZCtgU5I9y3gQiKbPXL0a76fshCSLwtRnyQeSka5UWZP7Ud4URoU99SD+5E+g
xj6/03yC4nF28h99C1Mjov8QTY1t8AggGLF/WPFwJc+jfa5rwb3waUyaxTjpP2rk
2JPO2iqA86oMM06Z3DaseDM7sQclrh8kkKXQbt5pi3LAxMLIyKHwHjYvXKYEBy+e
QgBJnK5avT35U4DNpL74Ft0jp/DxCmIW5vM4w99Ef671ObINXDC28IVEwVPZhcLh
xDoEbQ0hLEjkPiHiVZcIJpvOERHb9xoHIxQ3bGL6uKIxc5sDn6Mi9gaMHwIltkug
a2j2cXJuef/Rce1Xs7A6KmbloW7pxk7ZlonyEFU9trtECvSX25sKc+yhe9MQyFsO
Rk74dbVkcjoB4K2qHBJvuWfwJhQp4fPNyaN8ziACuLIJuk7Vi5ahG7/uHcXfebRW
v9cpNbbkzyQ2E5qk3Pq2ByKvhhzDg4sL6GxWPCWpqxWuhU6ngi9hYlMgDigEFQb4
sTbWN4UwwmLhAA8INqOnevoIKmKrqxRy5f3OxxEBW8q62YU54qnd57tWx+DRwstc
VPmoN6Bdc89AcFkbpX6n0xLHUWDPYQpAyHX09FPnGHO4vp2g9FJ3FJBxKBB+n6Pz
V9yu0V8626iD64ji5HkbKwlLGIiNPe6Bx8Xmf+19Z9Rfl3TerkoUrO7RCxBvzYRt
1aaIWMA2Mk1DWPFXVGRA2Y699H2/jDN9y6p1+mdX0XIvCV3wtFEzGWQ4GCTGzEXc
3ppJh13fb4HnMMIIciUhNSlMRkdSsiJ7knARXJLC3Qr8vGm2djCaAKVGk7SPGCW+
WKoeY0oXVYmNKVbUciiFqhhYx0yVN91cZYspD7OdHFIsceVpv9LFyUiYm1GdPiIe
dVyMGPsG0gFqRfZdHiPeVnrr7L08mRV5DFkp+6MUkPpbkwNFl/kOXT4t5ksq0FkI
X65nH1eagGVOyHNejBkwkHzJ8qL8WYTnj9fn4dtbqZA2kmv6O4OaJw73PIQCp0pm
ZTHyrczAeOi+NDGcowYIeAOHFmSYOe5woWUAmCmwg0oOZgHl3Qxbm+k72uNLRX+T
qlcDMr2QZNpjHvGX6mk1V6Gs0bljCgVwYRz9lSqDmt0sr/y3OTfZuCWdVyQTaNLI
+PGT4BxfmjXuFMn4E3iIAfWZmjCS1HvGmYS5Ag450TtgetDUEw2YZrkiKewhUNVA
fSJN1mlj38kzQsLnvx0ZxIQFv07fAFf98crCArBtq3ZnqnFn3mcZDezf3ImTylM2
QQfHuv/1vDVJg9WSJtuEZ0/DjTfshLsnzGg4qQHQp/rBrE5Fh/WJhtxrV+e6uwKK
MGotjfOEQy4ba02BW3DL70SJkMYOEShOoZTvwsNSECdAmuRz6JXg7SSB6tAW5gI+
AEjFJAbTCapbaj4tO7Zpc0B27Ec5t+bSXD+uqgYmDZYQG7rNtStHPcLIUVzTPxHy
sDfEa0Aez4HDuyCzsJpKYazYDJm74scUBIM1tzl6mXRhEEgEXMq+IvdXtqjohriC
8FEWcoEe6kBdeNvy5hwoPXyueIgSxiy7i3AzZYU1QRfOPenqd9RmJhJuNAqy6qNp
D3JGRPl0VNBSwaOKqdb7n5s9zhRmXf7WMkqnBI6j5mpiULVs9z1anQfKM6mwD8dA
RjXFHsfikJtG13Rj2vMFzN5mSwrxT39GWzYsdm/lrKikdUg0vaq9HHDQoXjDlf0W
zrSvrFFDGkIdC5Y8WbNq4tC3nDMHOPDy9/sR3quCfYqFvEHtWbm77rL0nE18kGvQ
Mln/o+9e/s/gUZStMXE+eaCMczWNc7xvz9pxNep3iiMZOnezpYn7W1j4NvLmhEVd
eH6ERSU2ZtukCvz4GQ9qZRIcVm7DIjMGq2zEPVBJ/haGqvCYTNsLZ1qLfE0g2gvg
N9EPUVcHMniOaYUY0jKPAOohWJR1sQvE35vYubRJ58/GqUZFLMYRbBRx+gQnxH/E
1B6nswk/NL+dfKIXl/UVmok0Gr+3ktiQL3zDp+cVokEw6Z2JV3dhiI+Nh+pRQO1Y
io1E1QZqCAeVs8G1zb9lN35+59LIxvsfkJ7HSkYxDV301yCvCoULpFVQzp0/vEev
nOHB8hGldLPqWHhEfJgM5ZPnbFLhQhNlT5EOIpTjV826n1gxszSKgKBls1fzejTJ
mGA+wGQDFfgjxcSS7307YAE8YdrFZ44f7rXKAmKOT5lGANdhYgXzEs7t/pEjhPOQ
JTHF7XJCWM2mL3geYmnE3CgbXKEyq90p42BeM3vtHW33nYtl1Q5jIPaa1ZpovuDR
vJ0u3RvRA1bexb5JshWNSH393F1/5xhBkGoOMhc9sVirYEwngS9vmid1wlpm1rN2
VgPCvnhCK5IrLnkImAKP1fBVM+bICwrG0T+DLyTzDZv98LUwT8jZ5+pJTy+n1isW
mZEukIwqm49ZsmS7shN916wcBLlE/rQCF1llKjZ98pqhdl/O2aIoNjilsyh9ZsqE
IcXTQio+Pn+HoT746qzmzY3bE5rNHXEFCbao3Nvb94LQZUMO4f6fCZ6KqJNwr2Df
RxcZG1OiSS1cF892i56m8cyzNmaH5RQaJEP0RZbqx9rqKTJt4AcN2YHqLpedJ1Ph
LJSS02GnFWTK/50Rs2z92SIbVhhklC68duDTlXDwtxWew7lsNXCfzBfkA+Aqj2Uo
qRJjPOv+IwOvUGFWXkCC06T1xbLYHg3fppWHbTQgmhaiQsofJdz5FYwkUUcvTx18
YdlUjelbUwHp8bKFMRn8uTgaz9ZsuBhjVf1QF8WXYIBAsQcWGtMMVbv9pThSVqUy
p8PnHHXGfyzu+A68IlqG/5IroY6Ya9eHFQYau37LixpGiOyR4kK4rvtQfSwvkOet
dS+wqAgJv/nbu8CqZyvm0zQSDuj9hv1TwF5MH07eDB+8N0BTNmS9fANkuwKnxCEV
os91uF8Vx0QCJXPfWgOpfRDZBKtSz5XsAkWZPr8Gz5nWwwtAx38bYfvrF7odaiZd
/qv8LblkcYH9tSBo131+jmx92k1UhMdDbBpN/bUwSwsZphDtIUFQNHu9IOxfFDrY
FywAm0fWDMKBv+sZOKzlVz0/T/OkBi8E/fSnMq82ZdcshYj9iXbvsJxKjTyGYG8Z
GY5B0CdN9HG7eik6AQbT/f5YJpz78Od08asfsFLFU/FEiXjAHnEYLmCRtLyMvjos
iXigLPsgC2dmyegRPMJHjOrhhzPO8swiJPKXFWiJJI8Pwy/f3u6whBpmfIGumZxf
4PhhWstGwHCh40i6l43JeALGT4fqwdpwPujuf+fg1N/qEdpWoxMAq3kfs5ftMOQx
eOxS/A+OoX6qvxOERma/+8oSzmUU+yHx7+deFm5q/Pqm0V6tMhUeRtzPGw0708Og
0yge0F1XZn9LJiiC9pROOnSJkN3Zymh1WNKtZAAOuBgnw2xDorM64APlOBveoncU
7Y7evyEA3gBR/xT5pq/7KpJnDx5IQv+GT8fw2WBWqrjeBFIWlDkky4cjtqmEBe81
6Vbchq7CHGgBpw/v3CE3d+Ttw3fsKnnabL2zsNpUkEVYbaOMfBpit24Q1Ry+ua7+
otlVdhkys8NOqpeuhTs619wZY0OjVrCtMTDv8ANF276YS5mO2QfiV4r/Oy8OdJZ4
3nlVdNLqWb8+96FSNnRt1/N25Cg+oUYObxhTasJWE91Oq9GyJYIx6TQQKcpc9JpE
Pll8IkjonmWCnsa/6wjhMyhzk6tXajcPIJY1/kqeanneLDtyus5BBkJQLr6oys8j
HnLp0TLPIm7bu25IT8L7u1xg8BvbBdy4usPbzknD/OH7R3z1/4oArrYx7bQpF1Rk
I1VjAetv57zDLVgWGveQmWe1u8qx1FMoV3Txi0KSgwAHY68f+rAlYmYHuaYV5bYy
uFccrI2oO27PKx3C1OLhGDHWmTebywh8ARJDtMorBB9DoC18g3Vx6SyvCV6ZNw3r
0FhU7eNusgvVxRe+AOl5Rr0/jIE/uXwrDf65UFMKhssekn3OUzUgDKxoQiJ82F9Y
r8grHfNxh0chnjYWyutETfXkS6dfv4wb1OME75mK9Zci7/voV+Tyu9ocV8T/SPO6
U7NLcZ4ytX+d+nq/r+4TBQimlnZCLtZRrSVOMYVm/32a0cYgK5sAd98SlFF59G9A
dz7qCdB536RRy7+2z1xHC1vRky4c8RlHihsxff9EMIcFSH1PRNJeyVAMANxqKWJU
KljwDOfxzqSKOkuBQpawAPPGpb1lwLBqnXKN8cNVkcma4ukZ+bFYrS4PUQmNG6VC
uJEvT2jGcUX5u1gj4cIhEwYRMi4GSt4q9Sn/MAjm0hMNjDe1Jva9NuTygunJ7bMG
XMfcmF0/3mNcwvVhJ+cWwq0dmfGVKBcZy8lMOvXUI9QyB3p2hbnWDbTr/h8Y0r34
YCHiSxkJDL08DlH00KWWQsQHGhfwLrdQwzclw5aaT44bIteGk8MSUTuu6wX6ePMB
mySJkv3gbyPusV755DGXtl1RTsF7wHiwrkJp/4mcGlorRbym1oEYc5v8LUyfBrKX
qwZuwshwcK+inWk9leLtTDuDtqvQWBpztiAod/0OAXkiJwYgllUsNYzYq490TI8/
D3J5bY5s6xuLxpNIFugdcpHjOTkm/0NrI1UDQNPK6nYVIofYy0sl6GrgLnvl1yWU
sxghtkAYhpWFd9GU9ghZbG2K8vwEm8TPYRsRNFkyB4iBBe4HvEsouH3jJL98KOUu
rDMObtsX4O0mVdeFJX6qxssg5loZUIRhOI7LWxvALAeNgbKNJufcCmCEqaT8a9ce
d5nQqpdBywedIf266DBR9tPewpRBlWnwc8Dnphypg2tOPvoVvTR7U1lt11nKMraA
ue5qUVyLARprDO3nt5pj3TZy/kKXrmA6HVoFB8Gtsm2DaMZfXl8tqU+rfUUHINNv
0H87aYEkyJ+2I7jZ966j4697giszc3USjMCvEcn5CeIynRm7zk1mCIx6KC+11Y61
qU9PXdbbodeUcETV3fsYc10mt3KCQxGJdCNF5kn+JzHlcXNNVXgMoQ7wwsAQKAkm
ZHjb0etIgcTHvaa2nGzrziM6eNpANJLBJoaJP+IINN63PV6IRYl6ckyTYBp36glY
OUzyGa8bbBPvC8qRRzT0tXOWlPZGy/9cLwux0jWtKRG1H8DdpGEfP+/sjX/6k5eL
C0tVDykUeii4ERXm8XkuUr1m6gLx4PAhZblx6IWnhEUkYK5/xBpTWOc32VHWhetD
xyEISFusYfn3p+LAXTKFDdwI79kfa9IhUF6Jmxw6oU6Q8+wWpzKBRio2R781Q1IY
2bFCuMas7LOq3WO5mZzcGyD78fNk5KifFYQ2t3c0IXk3OrDVVelpQFsA/BeNm0ma
gQfXGCyygxEO08dbM0RxuwlRNCMmUdl3sHKCEMT6vWNccS9Dg8Omqcd7MhYJmAX9
urZduDR4P/GVpZK7WCF137d0jQmaavVfA199asI8PcOA54dnq0l4064koLaY5V1e
8XT/T597gO3prWkEACKI50TeKUwycS77AND3mvsJh5UyDzF7MQGhbcc/CgEqDg4m
iB3bM6MiA7fOROhqZfQmNiR7YU82VvSoPyesDtpc9j5tyajYkFMLlQtpi7eeQAXq
hdoyJ1TC2sIMzMLtxW1K1cWU/P/ujo0L0B8C+VtwGZd386anaNCt/4tY3L8nOnrt
/kkpbAIuH06BpMqJu2W5eSQAHK5Zkg6BR+rJP8iJ4/AInkCS0IfSN8Z3T+FkiMSJ
2bd8+/DbMO8FY89Wg08lB7lQr3Gwu/9Ookg6YFqBD1JtIkiZzRzsko3Vk6wXVaVj
TH1coKJIYv1Gnr+Zv2ZkGaB9oxjY3aPF2w9AP26jkrfmpZHS11VsWIugsGiuxNgs
BfEtaaT/EFeQNZlXHmwZ+JN70hfIStBXH/Xh5hztovA3ti8E7Um7lmQlmNdVfRmm
7AaWcjQ45BBhG2JSE7jZw4BuRrHv/DAWjifZDvdS6OSOI5NSmgJ1CKL5eu0bdcH7
QZKIQ9SnrLCzy2dNbq8Jn87KN00wl4Mv+SgVDNXlPWCGlS41bJLXgAOxxBdnaXbf
0KEbvZigxJFIGPyAsfK7M+QD0VXtrfMEf1MriPD8W03VWS25KCIKNgdkm0dDTLBj
MVkC3Xzqg6PB62SwI2BMRGbqgzDMOVyFS8YSl8tkQOBBOxgQKYMzAP3pze1+YfXm
O9cpbB9Idn3HdaOfLF49jSCyZLYBlWbn5BcG1c3W6H80O344yQSCEbjwGPg7xI7P
Iy2/3/chg9sIbF2I2LVezthDXuJUvrsmc4FOAIlchUFgXiNMd0IGpisDUiwqKjFe
Ixkxi6c/JOGEKAHy5Gw/lNCB66bW/uhpDUg7gWDnv3B4NrbZyo/fnLyemdvxVG7S
26FxDNkRNoerueAzZuuT1xWVHSspQrxmABWgRhzs9b/fFPEcNYILxAEy4WRwvDuV
JS4nLicNf7hCTzGXNXZfoz0cZwcUR8ofn5rVaAH+XNbWta/R6jwNwUjlK56vPvAd
47vlIOYwf1qCJiQyiSFRe8JPj6YwfIb76p7c0VPYka+aYhPxurynDXmmeN7v2EJ2
PBR2ppB6a6aq4SM6r4aHRmuVVUtlPnUc+/6BXErBWKjdGZztfOYVUiwrAMGvayrw
P3ILS3QGfzY9ZNOWelz8TxHJAS76Njuwq0vUjrDYGAGqwnMFXk8GAhNHr3KW16eR
l36oX6MjcLgA7kv2AQre3qN8CA8UMV6LpTA6jTNP53ldDGDk0l6n2GnrQ9ABA0AZ
j/XXN9wI1JwyN8QvXnqKU0i3AQ0e3fSG3c9tfYyl1oD/EpaSwe4sqAQ5qbF2rIwP
P5RBfyVXcGAbmeVdwbXH7LVPYIBC4++Tu/qeSJG7cPAkm8f7YGFgXjRe2U6a97Zb
XYK6BSQoA6qbffwC7Js0/uqpT4pg3z0aeCJ7WBqJvhV+GLaGHOaOQzttJvKXy9e7
NIh5wO8+BH7XaidrxQvYQXM05jBdZ70E8oVs52AUOpN8588eaOd1DZDpioCLnjz4
AbfsFZrMW1JdrXgs9AxQhZ2CBJO9fTf90cpOnUEHy+cIqOVH61p6mrjkD1r0dBny
wmllU3w4O0FVcbRlGzdpZkTduT3AUPHN/QKRomIQG001SX4QOIJ7COgd7TMkIg4+
V8KC9qKapHyasdb3JxMGsaTMCmFqkiGcZ3DTY/H9sMSsrab/d8UAIWo5BoXP1tfx
971BJwFjogOUh6nc21Ay7UbUC2ac7EyIddDhPk7EwsS6tG76eJ6NPGjgengVuIj2
g4Z0+/GC9UFexFhU9Q/7W+JGN8Sb4vZSpybQLn6yuopR+4fkazfTZhv5+l4yQMvN
95SRrf7Rt2yAmaNReSmztfZZa8hpfGEGXIEqo9t6ciGte1lPA/Pb1DdATsIFndpM
O5M0Uaso28tZ0l5sdG7CRNATIm9GHAHoDXxwS59F8/8w8Qez/2AtbI1uDPpdoQe0
cDR4IjMwQRq6xccd7PRae7nCqplRwwdcqdtVcM4IgNv5y0CP7991U0gf0MnlWr7Z
YzKZlpEDbuFBjdIyNF8OzBMxVE5fwPZmix4B9I9ZtMVnSDbr5BTMGMwVQ9t1Rrvu
+dNT4KEmX5ARKpQmhO/wABVnj/HrXuQbWGkK4Xp5fZBGTEYjmVqyNJBN8YePB1/R
ZcSzvdjVisoEJgEpQCJl4B+YIzsIRDo0dtKrmmZFAA9z+WKtzGfZnLCWBY3eYs6z
GPBDje+leOjiCimk8ursKR4VToB/U4ZrEpgheUgHhHSVW8ylKB8XmQCF/ybcv8OT
LAZrMaYHr8qM4pphJ4VuBdQaUTtqWp6v7IBdrRJviTf/rb39x52piFpGQCpcZBSS
weyMT46rpARC2cqLHPk1tW2X2iXct7Re8mh0+wd5QdDl4S6Vk+QvJ2wzt27hUpkL
FccnDRg5JJTHEXZcNdDEJPK+ofFxilkivcDBEQdlQ3zYdSHc4Jtt1J3IKt6K6eUX
gJafHL4aVjfIO4jy+LapPzC5F1HWU7oQ4tvsQ6zRbRW55WQEJ8NwvenE2DHaNR33
jM8fMdTOIuNMyzz8oQFY9HamEBzbcx6udXTHv8578GZbKr5PgAla0BNitdhPmM1V
yvwJVT++9R6BbJCP7lefR9lwlkYXqnHfuC9Kf8gkOJV+uUOhJMJOtWmuM8qtRR1s
Dp6Fy48HnNFqQL7ANOO059JEFW+ODozTllgFAxl65hhDV0ZlON+snhuaXThDznZY
yX/amPh0aXdTQnsnL+nrlFV43QL78+J4fK6kawQB4EGH9yZwhO7uNs1zStCbd+Hr
0HpSd+UBDLMyo11Bh2oenfvcVQRxfAlPX+n1DfB67ZOIvGZ/Mh9F7pu05cu6P2xC
0KTw/ZeblE/aVXXisbh2Him+oqt7BUxe0pdZ07OmKdkj06a0TXE56Mg/jOp0GedU
3oFzlwpYibijNS2AoN2qCE8Rg+fq8n6oJ4QzigW+nfQoT77U1MG1eNkXRAmXtpNL
slZK2q+eiosglBF18zm3VoHStffv82Je4M9se2d/NlZZfR/KRqdGBzPK2FvFC0ET
JpmH8rPzORnzC3Fbu3O2tC5w01W7ziWizF2xahU02MKQPbxKdtQgeudfCB0TDxCc
+M4riSPGkCNfelyqfDr0493en1K2CrVQlXiAyDvCdAr8rp7Pwgs0cOIrOqkhsa1B
mnUFVGSMMpyhs+TJXjmhmlJk1s9FdJ+a1+Zwx8pUexas6f5qM42vmdoiJKvhNPIl
3c05wn+7zJwwOewtMsIP8evuXofNUpox/9GNNohJ84Ljbv5oU5Od35xxoMizeDQG
eJLnwZGCmXRrWgt8enx0YxajoeD2XVc8x97p5Cv6i7nR6LbKBsiAxym7gmlClvsh
W5kRbjVeREtkwKZqA9q2sok7nyUOVfeLoPRLAQDTpndR6ISclVjoW36ehKW02IFC
eJI4xacuj4vbULytvP+e552BACAHEcPZdufMnbdOMolvWpvv2q7NaS5vHTo44nzg
0CLpQI/u3uTmkXLZSFix3f/bTZxNMyMkX/iI/Ga5jFOIvdECg35Y3RDDFD0semdf
rdAMPiWIDm3TI4x7XDVf1FaIRIxYPS6Ul/E8xHt7pmJIKxU3NzweovkEOiojqKpq
HYGJUyTASwfLuUD5TcFwwXn/+N+1u8BRco2ySYAIQ4GcLzZkMcTTYur913cpc0MQ
f1JqZnxtUv9Fz09lXJlEaMG8G5SKwFEnTD7vfoa0moTgyjDoZwC5ufGtDz51FvFP
bJyEi6pG8wnlQP2wRsLE/qSPkSRRneGWwFzkpRGI/ijbmXSYkZ15101w8A/SnlLj
Tdf3N0h53p1yIYoBQcqEDIAugfGt/HbH/i49A+qvchpSP2q92kbH3DFp7RWWlHsV
9DLu6FQXbNT8oDmE9Aydk4cgbfkKPrCXxRYjA6jr248o9kslz/hNtcuSYRBhSdc+
Mwlgaj+UGKLBk9s+0uZ5/31S7OODobgSf0DOKUkgy8mPAzheX8OZYCbdxQZJ6/ML
2K9Sk/1LuFFCsBMiXsTvRHPWgdjPZQDvDg90z/gpe6D++xdUB8Huhg7e85zfUZTK
ObelMWTzFzEoT8X75QdkE6XRDh2/j4eRtJ4j4bcv2LSbXZ1zHsHvmgtFMBp4FV3x
SjRgIaGi5gCz4LPJpM5d0FWnRA4zglyGt6d8v7hLULx35ObkTQkHaC6lbelElB+L
zZW0a6QasSNcnMMHw/V8i1ZNaPQH/mDYkaPdycVmAtielB62h+2EAHswkYNVPMDn
SDcHmC2U2cY4C5wda5wpDAb2LY0ceKXUhhUVverjrLOLxpIeFC3i/q2JOSuOGqyy
kV3b0amF2K+2BqIF5pK8Xlo42fj054/3W1wAj3iAlt5nmDvJbW+Zr+6LSiuHy/Vx
hjV07VOm7szlRdAhoP75NdyskKTaLBzg/jtnSdD1Dtx5KgVzywVqxPulxboeGikd
jMdst/wM9UX0Pk582tFApaHP3cxB5Fi/mC+RZ4hg62bQvZW9DHtnu1NB/DHzET9d
9f4rwOLMVx6yGk/D/FzNNjdJPFSaUwMApR0Bu0Yl/4XDUP0rzUJfLXmMqnPioVA7
Io/qNhbo2sX92QoYemVvTDpbiXQRSjzOV7Y0dcAUE7V8qJ3cq40+AWezP1tUx5/I
sSZDcxnK8KJ4QGARigtSMWE9a7ULsJgWfFD9WZGd9ctxUxee993jVkr7WmaJKWJg
T5g0aq9DEOg+In4jhGTtYZYEsH4euE11reI8bO3lJwy9H1iEuvh5QYnND0WYBjxv
YX/94DRLRhM2+PF44CThMfab7bz3m5QOkDFR0WEXkzKcg1T6DnyzWZS2f1jMUC0w
/73Lf+M1E1L6CfdoycAP5yvzkCRJEvaSq4imeiV4a4tL0oESbF44fybdu8uzsJr9
0c8iC6G6WqUBuTTa5D2+qJWEqRbVQzkHYg+Fu9HfYU28DHI0e3wa5bZ9MvvXFW+3
hXzW9c57PKEg9Lx8B2hdudWcryubqITdBDS0hJpUKBoSDQ6g77dId9aO2SRFNxsU
7t4EmorPrHrjTp7e6OKEI7fkPBmaWMHdVpOrXq9QV4CEoiyEbpWUFIC6lvDuOoa0
PTGagybI/ki0nXqjRUxC+mprfeWL9oQo4KhmdLEr0CUS7rUiggeYcsV5Bt7pOhW5
ewKNY/vQ8npC1ouEYMFALmilnOZpVybD3Ph57WsG7JwTBXbEQ4fJyLPoG1ZSSoKG
Ibr9bD5+unFZdxIRz/n8IjN+RbIsiAHlpKniT0S7bnAMguI6WvMNMBFAEPWXWWTw
v20sz94avTNe2e81Q2XwqbLPJ7EcAG+uiu/aKlIuZ5hioWwRGWS6yEM5ZMOcA01F
HfymJ0Hb5th+eg9SAyVo4iAD+BKPgfHsyUZGIhIp1jBqcEbN7BlOLV/NWTy9yPAH
dSWHOxpCdyF7z0u4cAB5prbP7UWzYYd9ASdLocGYFKY24igfgtXiUglxZelwAy5+
+2N97vFhOmur6IRahtcFFDdSlpbrZUyuE1K6mHf8oZUFX3egfZx1KbimrdaNFLR2
BEoTMtXyCI5x2Zsd6ck+KAo6WjAsChBRK4vo2+bYaRRifwWtvWUBgI6MB16muFo2
51vWSc2yCI691PT7VE+v2m0l79fs9D3N3viQm1Jn9v8WQR5Dv4SCwgPMwyeIFWRg
bhrrkRjz50pvB8stuFxSEQZ/ARWi2sgT9XGWePllhe4JZXpCz75CVeCrHbjXsDwQ
bsq6vKW6FFcTdm3dnsfNK/L/8DQ8cX9/6YtNWOGZwzcw/D3t0moN7mUUm4ZEal3n
M7NDvZd3/PaVHqc1SEXwHbXyJxTts19qoXsiSwEmZPXdAvdsUjnwg6xLQVHtWzkS
ulYF4yYPlclqs2hkiAqNvzcuuffjWSy+evMTfBJoEhfZLb1XAZmvthgfNihb3d83
aEA4mvtEvt7uPMoCX95GIDbnzmWU6OG9v5G3pBKLrwFyj5z/MCYnI4sTLlDjw41W
U8Oawmb6X6TYjvLwmpkVQu0yZj1pLnlNsuFxSOQf0dCXBdKuw6Wg48Ygx7VP9RA/
zVUk6Ct8hNOt7q2pZAs6hiheKxW5YYOCXx0ja7ZUO7aAjA6dX+1IbEoWZfw5Ruik
w8oLdcQZkR3+nmluprmBsTYvn9MXvJJGhh96rYyWfonWNBgb1miCztezH2KJmWxj
MrdsKwgXLLTtYGd8cWORPQDiJLzTXNZoKBUs5i6LroWxxwcoCGN8An5FntAd1XC9
J9oJbh/7JYgNaPgHUHnVUeDGDWFHxtdfoh4203DkWGWpHTMNg8VX9xsTKsQhVzEv
G4DeHjd0yMMRui2YbSt4ZvFGWYJgKfcj0zaTMDPHWAu+XAtdM1vabm1TDYMK6qy8
e8J4YG/xmDTTs/K//sO7LUxs0eV/z9WTEoaJFNw2uMD/SsW9uyPE6eeiRFF+u+Dd
unfz6AGrgEZBjrGIGG36vxuZYU91NxnFfg5y8/hCZ6SCoQS5uruGknC6MR17TQP/
oxjSeeMAhGRBVtHIhNlYB6swYvlIoyzYyIXOIxN0pqTayBgKbf+aoy0T3VGxsstc
zRwn2rkgw7hYqW15AfQ+hD2wz9A94PEt44JT4C4K7BAdjzvNeluVo56HIm2V5cbf
RK2+EXumfvFaMmoIlOJUBouHhPnJLyBYfAu0X8rVJ2yFWhj3ThylgPPPWikl7sdW
rBRKuycp1PjD1qDn0Xgfsfk0bXw4z6wvCbx28nYQxhXQuFXWzAXgtHYSiMxEdb3d
H7iXWiwwvrkXeAMYT3eRwpwwkBhZfIiYBMJuvRvxb/hF2W1Jcwx3b5v51ZSCI+kG
vxfjUvbFnCNXMTiR1o4FHXFhl7rwdJKoKRiOQIPXAGihTgmThpdVgOguQzFBorBG
e46AqK23d3/1k8PnD7bsxJZ7/WfEQybZ5qteyX51I4IEb11B0XgDmxyHStJyKGrP
isYgeBTsUm61VzvPRykOD6frSTUKBBgAmSZe5T397aDnU35m+rAglY0f3ImcCW9+
1TUcTf2OnusQqu8NBwt/pyPhIiK8R1P5o0hcU1C7Q0GKy1xjJULm15nKyX+Nw83V
rOmH7T/6nEW1tkIoHMZGYstn1VcI62HmS0Y7jusGx0nILKldz+EqXLX0udZrdujF
ThL7KyaCo5az2D2VROHMKO+FM9hRT9tzuwqnejN4lN5rVGJqrhuGKuIGPwVMtxeA
uZF0Zm67UUKa0+zgJHQ4n2D7H4jCOitF7OWP+5DQt5aNbgNWVAMIV4dM/EwFsCyv
dteDX/jyKsDmDsSa4ZZBdI5feOJWhtjg2BfyMC1UklpyY/OXLcz7vCetHvSk8T+I
7WdJhwmyklont0chwW7wVMi2oRm4tdyWq4PoTbCoTSpwEbjjuzE7Av/n9loQIfYh
F5f9ekKqZjb2mxYnsacF23WEK2oBhh1K3p/HpNLd398VDRBGfxXOJMt1dhTUoOLV
ey4SWHWsfIUX59nPeLvF90s3y+fjfBGHOkaCwEQSeojJVvOTm4NTvILLrxq2CRq/
ZcJ8aBrG5VyJRDqM5Y+WART6LToPVHR2px18TaWjurG0QkYk3GGWUk3rd9yJXPLp
K4A7KhxVLGa05RrkeWWr/D7D/3t+ZAbAZVHsVBNWN9ALfvMbUOVufWRgdTc1GJh2
TxvZy5re08jAWsvr9pb2YRHAga7wYGksngJqjPkkPi1CdFsQG08hKoDBZby8+/K8
bX4CTd4Yv1aGawmnbvbU9l3YP3UbJvF6BX3eWee5K+T3hX/tW/4N7/4x/1LW5U7X
F1GbxuRLiL+3Vr0T0+p/Vpgs1Q7g9MiOqjitbLC5j5sRG6V9mXwQigXNB2ZVl/6G
UoIk9ETm6/8M8iUbemWeUd+FQeq1Lrc+jWDivv3CIAH2y1khlAtBC+sHhCOm7QGt
5sNhP4E4t3+ObkAcD6DG/N6CMp1qsArHClK5Wr3+pRf5fvD+sh5UniAu9T6PSsgx
Kglz4ijNB8X4y2YhEqr5Jygk2HZ31OZ5mBqBNG2JaWsRF3eA1VDZ9GZxF5DvwKEc
QDHw1de8gGj3qAv8J58wyE0pLO3AMisXWTbcB82M5XAZ0OXrxbDSRIqw8mdvy3Yy
eAPFwfgIbo1OdUA7pcJFo0vsbR1ZFx2wHkUFdAfe3ql/DZP7ewNWoqZUVgej7peg
JflxlhNvPju3jE4ch9dAlt02YD769n6DHlf65LbPAA1F/U07U9ok8al7psMhAaI6
o0fkAEjjDXzLxipoqn2ZNRZLWMPlMa+irXb5nqYxRRCiJc81hwqUihGaVSkEf0Ok
IR/KZjsxh19moXGcbjWiJVilUPZVXhQi7ckW+IOiVBVESF6Y0W7q6pqlGDR1iLKV
cNsubizM09Tnb2HJd/BJcnjpMMbghatWYet0D/bLF0q+a/7DKjgnwpo9uI1olZAn
jYYjeLB/NKPlAV4KqHTmn/k/NduIK8iZIPDblvvehIkdiZtyzbT8ZdJSko9015ib
iin+wWxVlycEfZPipQODqcNmcF5y6QgjLUeKmNLa9leF0fMkyM0Q1WgEyfY4IGA2
pEhQdk2AXWhtNQsyNQXpgSGfOvBUIzzrwuS60y/LGSFveyWZrpsoKASLgA4QOBrF
rwzDbgizk+zJ5TZO2YqZctudpnDs3kRCjz+6g8UNtzlZ5jbRkkL/uEznr5R/GpWF
QwFtL+UEcCZ1qyxOtI/Q+k/WRtj9+ueqGEifw7b4nyIKBsc4poUip/0Oz+Jvfsav
qTZWwItLmoXrnvCmMWyJipJubYSS9FrE+LApjVKbWGXEJarzketCnbF8qlbaBtZ8
GenX7/eTDI5XJMdcQciTy8BHgPsGCcNUwZFIcA2b+OeZkR9eFFuaGZXOw+2eAOck
956LnUV5beh3Gz9u8vMh81qPagD/R/aHxsBinxmJ7qej3yDPzAVc5cJ/dLb/m0GI
CqtwzN35089GHws9p5s6EskYckq2cnXARVkEL91bD5jJpb6nyRrDIaT9QJl7Mtta
2LldgddLY7X6FXD5uAxYUTf3jitkwb80GloqNAsEKxNKXepHKu7FHouWAjDN31sG
r4PidLBNmty/e6S60aBAqUBpUHhfsGHtItfLhw5x4Zod5ennXPnbGs1XI0Zj3jAq
u9jimvvCgfzfi7D1CXn9csj4/U9PKOBJOTLdLGMDUNNPoSvOiisWoDqWajq0YT/o
/VFfYS806Wp28YfmDBkh9QCW3AWxbO8ZN10CrnmeSmuCyYFi+NvW2BO/G3mnnysT
0lxlogw4SeZqfQeXJ7AbQd1ZH8PxgSAvL5tJRCZ5LMrHlkModZnCg2DFFdjdRq+v
64M9esYr8PYnAgUlv7WcAt8ysQCjeqY+vDd6B3vC+l3BRAEUWGo2lm4lb4/X1+9a
RWgQ1vZwjZR/67BL+o95xSmGXsZhQyhefC8hUMEVJQWYXRQM+Qz/Ug/KYqQ2aZs8
Jl+ZNLdDQup/9sxA8ogbEW5jQOTKeL8q/UIbLpMgljDDxwxmDDEqBwibP7gYgekk
6lh/OzWW/02fOX60NaQzYXUChDHf/hJeKi/Pw5ydk8tsOEJPA4lpUIWOUYLPks7x
16OrsucagbLhnK/CaLzi3/eIVV4lAYcCRlqhm/4DMRq+T8lqxl9GkkgmsfRocF+S
x5Tq0RCQbqvplHmuExTBq1SOwrKHEBFRkVLz9UwULWKFAc5RoM8iebKRiqZM83cG
NtV8rYLVgCxcn6VykB/bE7IOja/Sx6qFUOejSk3QKuO4M8Y24b3X0PXDspw2333d
k/LFnPnC7A1lxTkvY4+fnqkReW3HVXU37USmM5uNmCPDYInuPqiAgRI2M0Wu93PJ
G7r5ASqSdPUeOwiXdkbNJykd34T1vGNqxN21q7RkNdcC+rLnF7DnV4pw9xmxntPy
NyRZnpDD7q04AaFBveCBBtII2JVlYYB5yB6O821cB32vda9Lp7Rg/8QPuRwDOz5M
ApvFMw6wx6lgCPliCl9xLF1gI8K1V7fcFSA+jpemSjP5bcgh971gyAMHP10DkbdS
LLf36gODDGZGfbNmfZOwS5upboWfLGbH/dyaUqesqNj0ADcXNE05L4FDMCMWW8hc
yrq8rrIjPrUQw57MyAHQRFCR6FiUMvYPSYHxMidJouFAG8lFMGxFGdiQQ4X0aVpm
QODR7/od4gcqLoJ4sR3AatnY8mZo3TGRUF6mODU+Y7uAfjlxaKx/+vjRjF6yru1b
bw0mdg+Wy345xtctz1kDGIrs7Sb7tF9NDnKFi3k4blJA/Rc7u82HGoXvKoUrn6Z7
8E0ID1Eeb7/OkUozfrWXu0541I3/ej+plhmXvcT4LT07bIhBFgBzDKASZxO99NVD
XnHRsYt050SvcgLOwEZpml+AMChSW0WSupYEsDW7vpHTEUpGTUWS1w4PoR6QJH4O
E7s24wdNaDQyCNIszG+1YALTEdW4srswiU2ij485S/kQ5pvp6c3z9PPTZ6MKpyKP
UC7LP+teh1NOE2l3rb/1gI/LJflHf+yaa8+5vkSdL7OcD3vNziKf66NQJWj71wjr
njyVfnj3G5UH39VgxQil/ncxQP6cPB3aYvSXN3XWoUxqGjCTFSr1wJZkpvZBIQfw
0x8Sje7N+GQy3GaxHmIX8s2JlqO4gkAsUQCBhNg9jG9xECkx5h4GEbUeePbo3tzk
8YpbIlXpzOtJTzz58nJReQVtZU+rStRPqzKt0Pgo+e68/TZVMwKmcu6bBrMyKlDF
UXh3ro2A4hCdVWE5O/ZEpu61kVWy2eU0w4WlGoEYdk9zE/8Y+Z/ZF0M/4a9sTyzc
luGPPeYDBe/sOOSoE8DUM+vZ380ctJQHP9cEe8GTHRTc3ImfyPi/RSqE+LMWuZkA
ClyQ6e6L8ccsIjoav6NBLQSp/u3tzBfohYy4QsriXvSdvquF+04O5eFRB6YwshNU
nDvSJBCG0e1+wMa3tqd6s1UAzM951KCDeL42Dy+DIcvSWyh6Lp4OzG3TCjL52qhR
rUq0TzPQCEbky/XSLoLu44q9ItmI6dC3Hg/5YXjPIlRE+GsVpb3RxfbOTKzFzKJ6
j/y7lx/Hbt2SvvAlYLKc5U3bE2rJ/oJ0wgwL4g3tnNlc8EqFwzx9NacO+M055LmJ
JU90TgdqlPtu2L90WPsC+DevWuUVRTP375TZjiqjbgICwIXdIFrvZAbyUnkv1QuK
/ja7IdiWVq96+mnxjW9Yo/l1/xkB++gnIpiIxBePJXUW1FxK6bS+mkByxO4GeyvE
U+dIDmq4v52W8DsufMsbkuigJzfSltUZDXc1tGnQAAi98VXwomxbLxmQtKm15/HI
kNYlmq5p9N0cszxBQD5HxNGaHMOKyi5Neu4q4/QDS5rnzDB/KVyhqPC8aqWtV3mD
CHngzsdQMyr+joaJtxxtd7jBXO87kLSclkjrybcwdB4bu5F0r2KjAy4h3Kx0TeBf
OAUAHad/DraPg1V5izu+EClKwq4J3XBNqa0f2DHfa6Q0ZZfCKxQP4mDUUG/YSF1g
rXKSGNlUuVfvn9m5FrfAUSuOw1eorCIz43nxMkTVsv7zKKbQYbwB1s5tI+uWo/mF
bixmfj6i7nBx0BylaLdoJ97nglQe27lSKk7hy/C0vh4zzAPKww4ZbihOwmfJBtlN
CXFOnPWG+3DS6zS6+N3QEkUpAYD8+nRdnI/sEeyB41FCQtPris287lZ8qOW9BFYD
+JfmwCIu+4lCMgLFe+pEeX8KrbExf0kV2sJxdsMIYdf33yDtIkXOrBBNn1+rC//v
tYYhdFu1Q4YuML5rP1cf6HQGgpdBdsPiSvRvobaJLvMXS38THoenSY4XlmnBx1hi
/rooa0sYeLgkxS+DQg+TlbyPHpmjbl+hYbbvecpqkwR1oUupXLMvqM4APOQrgdmm
2zf4SeLwGYy9hiW7eRFdnRRBVlR/eGVyaIrVIpwf27abE14ier5kNdyZKMljHmIc
W6oki9G4FnN25DEhzspP8zkcGIyyXnL107u2pVcxTrSlHifIVIxUxM5Kqcma+KA+
OIpb0lL9k2ibWHcCF1SmnyqLk5Zove3oS7VEtyRyVG6ujAR7SJiQgb8LZlnxSHMb
uXT4U41tFrW2K7UdLuzUzwwCRhrCKxNOA38Q77mTRPWWiLoPqc8+WF2dB1XSlKBO
0DmoTKkwBMM+bN9b3+H4qaJd+bZF+TemfOhFEVFcGUZbMj4ezfTa74czPVO/SHPn
Zl/tDm6YSumFsyXotb4P7OOw3DjZ5G0z5iJWIoOTNKa9uc107N7yNyvtfZUa9LwW
zCqb78SH2PjpXHrGkC5xVPuVsdbjYMYPiVwPGW1UudPiFMJAeI26Wy3GFye7amL9
zAwWJ+aGtmS4iEkxJ4IQFJVoajQez6LPpCRzO4NLqMkN85ORkaGq31/i2yenPGmQ
zcUkQ4K7SUwhetxN5udTHVnlZSUPBtJqwzQ2Nl9JWw3662pp2Fck6xHDU+Kpj3sA
SOoEKwKhOmJhc4aBcMT77WxDbzpp49DeSJiuPhjAin5TCDkZR+SQe9r04SQiar7v
oJnx33ZLETX5tDZmA+5jtP29WHBM0rGPe7FMZ5wfmeLS3E19lRo6KthSgVMxkPqs
SwQe02Q4baVkrkYofhu/7vI5T1LYykzMz7FnRFgYubH7oMer2JXVqzSc96DF7zB4
xP2OQm/IBF1CuJ6Rj75FMJfylTqMPSKyqtCkh3P44hX37qnS+qImgKiz/TwH9mbr
R8HbtY4XxzSD+kwwHZP4DqefbyMs7HZa8H2r65Nuir8eFJ3pSJEWFW1NiAvCpSwX
G0wGpFHAXBMd+V+JFE37ZNf1uIzp/vHZYz/WvyaHhyeYZpvYrwBBgTe4ALylYHl8
kSfjMeA5+qzkedGUpaVXSQmmoxdS+gZ9FwyBmjlIxSRNTQRO5gyis6XmlabOikfE
zBGeVjzvNgBSrlL5y2sIaqrxb+lLrdkiD4+aA3/Fix5cEPmwNY39j8CnB9GazHsx
gJDbpklbsVg1hI6zeuA5vkjfeO+t1ns0bx6gAt8odS9JEKoX3175Am3E7Nlq7uBu
JFF7exZynAGzJu/h36i1b99Pfg+bpU4VXYULhManWwIESjzO4GHklSGZBt/Y9z/E
eb5gUvDSBnivH8weKmLpAnk3dTBBZArdk3KSCm3dDwd8mvJJydJI/Eb7PsSC7BOf
O3ArOuW4rz30DWx/aYyaLhNesCSamY3S2PvXUUptkR/TpwVve2t5nX8GVrnP/vrx
wi4f+uf8LyLW6v385xinKGCcavQIQu7Gsedw1c8/LKz2ua+eMu0JPhj/fJjQqPJZ
YqqJpLQzDx3ehbv4dqVjza4nJkoM27KzwxBWbpPiC67C/5KL+Ib3pJHAK1Lpuqzc
WyTFUOm/h7x/qUf7vA0TjB8C8aAp//g7+XH2thj5tQlumiRpbePCN2DGjr2tMmRj
8A/+3/jVo1p9DjGYM2OH5d63/e8U4a7M2DenOc60PEPEcVFi3g2HROmX/zlxCtr6
kh2fx1JmNL1+i5uBkt/rCB9MQqRnVDZwpxsYz5ZC0UDBpBPIIMilpjHKbh46uN1+
sdsuQ+7LA3j6+/KRxzcesZkNBSP1qQtF56f1RiwmoRbK1fiY39EBeCM4iww8Palk
NjVzb1MQgizHsVgC4+GwM7uhGLqwhcp4w5GOMfXolGp8tg8d9maMxhdYGKWNCLmy
jZzLvlmMsc0GFzxkKhfN8T3g8aZiQVt9ujEYesU5sWJHZsV3YmnDlSikHiRlnrE7
eFKjuztMrft+1E9uuOzdPNer/lYQs0Vye3hzqnE9Ckw332dxtLNcL/bd34+LrY8Q
FGnQb+HXLA7BSJdRLOtFXx8zQhhccIPvEdiY5ABFv2V422k38je7ySjRzSbfHBQK
zEJy8BTTxv19pzskz4+ou5grp0PtRCVfua0HFUWtjcnu659C1L2imTZKLA/oe9Ia
Qm4a1kJdn62gvxFK1m22YlP0rFh4Uf3yBArJYF5yRU0TXzIF+PXuorp3jCtE+JyS
xWAZ0XzSSBPdMSRBcv/by0sFVNHZWkQBSUeJFNx+aVQZQVjLtEfmWGAm/BAwcYA7
Gs9TXrWnDkX5Sfa9lgN7JqWN3luA+Xvylt60GMUDrGo3emh64aI8A2B6yNoThcRO
s1CZafBsKKQ4jk2tdbG8CFjZQtxjc8UNp29VTsdCpadZ9HvCw5hmA9LSDmLPtfnm
mVhzlsPuxtlrITKipOlnte41nzqUgE97fZMUy9TClRynjxYJ5jT4d2UxX1RSl3x5
YaR/qtiJA56NPORLlKxzetbFHb07tQHOtnnaSvDEVWRZ3jc+RR73qzYcRSdoYVgZ
rpSXMFFO+94MvynIGZXSx1g7CaXx0J7w7L0SohGxDHbgoNmCc/DZg637YdRBZQOc
aAFl7S+eR+BDM8um/tZPfyTTpIubY3xiF4myJN3NIETxZVy34+9yabpXNnVVKzlA
uqqE363HZ1I3hM1MkLRmPJpP8dw8LBvaYI+8Kbdvl6/bPR8o4LB16jJWeXDNxMj5
oInHiRJnKmk4lYPvJOVnPW0HAUEm0OH3Q+MdGniV4Yqif0sQskY2Y5p0GNViWPxs
VWr2vPL7xDxyzSExWEkAMJ+donBPIk+mIwRpfHwATqaMczA8Ycww4rPpNP1uxipW
il8rozOlUM2EF/g8mYB9lpuZSfnYVRSeo/RScnzB+hKyrqjjGV0kD6MejXB7SyyR
JOOpXtUIeXCK7LYsepfrMJUpU8NlJOce4QwdNJSGiuRdWZrlNWznwDXSCRJvDZUZ
q7kSwSv0iQGHcckpY+zyrXukv+9FXQXAYu8k2Wt+ovAJB3IhVC03+/3wLoQMoXJu
lM/2KmzK4RmVYtl9aSHAjGCzdMzWXZxoJn2N7x0vGSEusiQowOFyZ6gYwRYvkR6W
Iwzsom0tB4IdhvVKyrc3cIR0yQ2GbW9d9DYmTFzKm9cTzIL7gh65LkxWiVmjoZOj
2Yunidg1ydcmC9po2eNNetdv8FWb4W/bVBXTQ8NXwxKZwts/bR96zsHkXa4Tp7HX
yMVwnx/60i9iZJAzEEOV2UZxknm4V+qCztYzDm1bdhpiHoxT6eL8cORcDiRi7CKa
5FhvQjGqx0ySbXQy/KNOzFenzYEqb5D5F8u39HPyulZ0N+HU56EVw2Q9HTPCJBQj
E/1jdUyP6LdxrAEN1M4DWw6GhopG0Ei7ZWItotwn+ESqcEvY4QlVv4C1myr+JcpX
r5512TBm5mvV7ISmQ4AG9L5G0Te3zZNbrdsypz2b4kncHYoILNaUPTcf1GKYVsrI
sJR0jto+yHP+TTEh8VexGqUS56mOjcoMJx5/RLAue5C13BuKAu9C/y5bT/5KSVXd
h1UVvjnFfX0S30pKPPrgolhwVx4lY9YLfcg1RtTIJIGGX7OZC5RpPp18eUMM0VPE
6UIvetXEtI6RQIcPlcdvkVl3isy8j/SzYBpFK+Li7tO0trDreX4lDwRytfzBT/Vd
bx9CEWazHpznyV/OqpUZvjX/2IchNQMMdDV4zUcCkhPTjeTTm1CBPkxBf2b2L7xg
RwTLX6snLx7b0DJjBukl+91Pr3veNHF/Iq2z/uBB0d5HUE8H4Gl0x4Y37Qs/am1V
EuZwgonsLmqyYYCZIgYCNnDWElUyicmroAR8iBlw2LLX38xz44JJjCiPRVVY5kJ2
5ZMaZrybDAjRuzsQ1YFmSY4ECh0W9abFX0wUU/VaaajGAayWvS9ICFyUagvrHrOD
R5thyF7Tv42BG5B/I3tk6AmRlMM12d5VTWVU+0uwOfvunz2UbvLgZzWVKOIHmvMj
dm9DlEOOk+itl9HIWT1iqY8g8IcQss6ZoCdFfNssyhcYpZ/eywkhSkSHZeE/oqSA
QVDQAay/oHPAnLjKj4YiqGEgvwy8hhNWA8I36z//9lwsVICrseGgjxH0S0eYIxlY
azZj8mgyd3mOazNgo3tQAQjOyX2fAhJbp1YO3RqBkj1FHo/1tARv7Muudenf4CtS
VcwdqNxz4HEtzZl7PjgEY0/mCLY6TvJb38fmCYEbqc4sNwu+cOUN9r3f1Vgk0WR/
CvZVLNJj2c9+DRIHyd+kbqfyrVqNa9iEsM6IIaT4A5zENoRVhIJt83pMYSyVAdJh
47de1jqPOyIod/ATpcp1qAWKGsL8wx9R4SgEsFrTUBq/amIw8PSwhlU7GBid54J1
5C/nj77V/xBPv6YpCfRsyWi4PdWZMYgI4tDADI2KVSFuz/burPxNNCiFTBKyUfpG
UA+j72My8WyonBSNOtJYVxvBHzs+oa68tOnCVH0yIQQ+xAUemOZZF/P87b1zpyD2
H09lAroW/DsmOlj1IR3x4k8dIKJB0ww9LJRH2PJWll/Jyi28wDYGg3ti3Mu7D2sT
NYZ0wlFCIW6sg78sUWz7a8J4pP7EzKmX5Yi8zDZ5DQM/FPF00lVvSJa+3JPOML+Q
r2AWJHfagQj5AV3Im/mBcTENGRZXLN/74jVQDP2pFbRT1absFBwKHROlT7Z/t/Nd
5ocOkvS9PvDb10yHWbz8pKe208+gm58khZIvpnRCE1MvTGPFpmynFJbiKdrIUsKC
MJsw9wGjcroHPUnBpegZ4PYz10WWqQ2LF595UbTYZII0Fc0vk6rGfF/Hj9TqvEYw
uIJPkJ5eXmBCvm/Wd/Wfc4CuhtCXkTp9BOZ5z8sic24XUbZBIf/jQrbcUsvyC4wb
dl8cVONdQxTQiaUoH0LbrO2Ve+sMT20tEoA+5GQKdJt+GrFMYQXZGQ6GhLTWoBNr
DgC1VI1YCXlTSlNeIuT742XOCEigQbJHeM0vfmUjNx6W4FQhf6YCwa1N1nEcj5lC
iYKGWhDkYPyMeoIdLjQB4TQOmSIKlGm4CHSwht8Ah2ekod+Pa0XAOU2AQuR+UgPs
yAw4Wo+aUsiSGOLOhDJQSdPBlnp7/6S5Huy+z9v97UO+znzZw+Dx1N/pdcroi2bQ
lkVXpRQRyufdQXMz7ZGmLtYH4GRTa68lMGrlAEqNpX65d5fH9X/WuQMgtwImy9nm
O1CN8VvVoJcouMKgWoLeTnBjm8ZoMyhUaETO02rs34/0jq7qoeX/rK/01gwtNhKN
VGcltj9jAz66IkAWZBMBZhgOCUcR8zP+ss+zefPG6rTQuH3J2AOcPcfgYJ7S/bVS
Np5G4z1yFtMuuVF6ABslikzwwyNDlNZDki0nklkkkZqG7mh3NPgfNXyoBluC56Ld
Xt1CfWzoId4l+Eu9nAY756iltrNcXC0TAP1GvdkMXtALkj2tx3OgkN1uw9FjH6Tp
d/vfSnKbroJzvvjMJ3NEDT8IWsQ+2vJMlZzU+pUackra0P5Q/7KCZoHy6bDbHriA
ZTmGE6wITZ6EW95fAS60D1APJ5fd2UQ3V8HTq95WmKnPJuKaz5jzkVCP9qknuNBi
qvaprjoIjqixX8aUCFQnNYvty22EURgpAMwbFLQHemD2CV16V+/4DEZFbjnjHTlF
eeAFxLRzsv+V6SbesTtKmJx98BKIdPi8a2PKDfs4mVpo+OQciFjouWEkC5UIrQR4
9kC3L42WqsTeoSP10smuqLwH1oRmWQVD7tT/oE2TM8+oDYa8rmbdM8RonD7BEHhz
9QOAA1qxgDuZ/4+3aJgg6Lc28+r8AI1pm+Tu/O33U8kBRRGztMeM3LjT6kTu43EE
+vqJfi2Q5a9lrkqEN1Z4sRQAcOacoo9AKtQRoxgsrrEJLzxES7rIpX4DkFGx3hwI
taPFx4xz2z8TPeyA9KTh+m3T1L6yTshK7jNN9dUfxBsN5++Z0U6LzN4HpHHrVn9m
E0qr3rmeSYdNIK2MMH/afuliqsDyqAQpYvuxBOQFnP2DAicDDRbHSo1u2KoA2ajL
Z86EJA+aEkaFTqIM7Fb2Edeej8qP4ZhZsQ542RFHDdMD23o9ygJeZGdH2wmV9Qp3
+vO2DIa2k0U8GAm7bhqDGU7iL3rSgFaWpSbCkcAII/g+f1i5G5WI0QqxWCJ0yf4C
fuapcLbZrHicROGA3byK3HTZCDJ3cW3HpaTEWkfuj1c8PdiRkvA1craembuXkJiE
eEgek/GlrSlBxhl3j2vng4I174GHPJtXV82qICjch0H6GtzJ2ymDcmB5OZqPT5e4
WABMerPfnXgAVFnncFyHIYbNMOOq8HCaFJOKlOYFI+LR1Cg9yHA8OYkGzdZyIiL9
cT42QQH5CUnn04LZLfTIFamgSkSXwqOfe7QKFJj0aRsnMgNu/UI5byu8uXbQOM0I
wy2alQ6eM4zoXhRzWVy5lGf0zEM/uX2ib/VHeJ6msRqmkT0cUk2I1js/zLQ+D/6M
0QwDDmC4pqGVuljhF81G1BfxJ7b90NCvVlQiOwXP8dqc1i9ScIuJ/oMAY6SVSiHY
paClURTgYFBB7uSAovrH6W11WrupxgepoJD3DXAl5H6jXyEi1FNgwb/Dj2dCmKch
rO5fj+22UTC+5ZKwRGToa41Z7JhgSZqrWCFWLTGSDmyQHNx2ShPN5jtGsSKQ5pzD
pCQ21vqAmU8Sx2fz5aJPSDhC7kRTzM8R2Mk3XfYas8UYp9cWGYniRbYMFyj7f8Ry
wx0Bo+f7rm0bDrAsD79UaK2c4/N+y7TvbQnqP0+oiuk4zEDAHgBi+8ig2Rs5zclq
wG5JknRrBNtE695Six8caKnHnRT2IlX7z9Umz3hkdt3rbiqpMcgtDwGIVARU+J83
SMrrk2qWezeM/4/pc3OUfUIl2ANd1D9IEe3fqRZ4HOq+Tu/Y7qyW9kiLIIk30vXE
CVKsuob+R2X35Jdc3E3UU/DgMMnAYNJilgoQK4lkOzylxRH8KXRxus+C1N8Du9TS
pa2X2/ISNNA0cvpfCdbLrztZ4ZwdwF5BwNG25p7cTKyXommfr8Bjn5X5ZWoLONCu
C2vMjZ6bDkZZK1r0pTK6m/1+hsnpxa0crhpDbMTwMPHT9OBTH0CR53fBHQlCV1Rd
irObrm2Jax6Je8O1NrCZPKAB4s7GZ5doxBFxTrE47EyCaNwLLQDNhx/E8duSdn53
kEELPJlSfbzs651pKb/e7ISdttbhK43jnayldT+E7MjLvsbfDjyLSW+R/vfBlvF1
18qSzWWN++dtF29ra2Rn8VygoUK0/zq1zWrVT3T6kmdXG8z73Vvp2K0SeGKtIzyc
UCF6v1Ptezc3BRvj5oy7ZXIiSpb/KIfqaI9lwux5eP9pApRCP4bqHZs4ut0sB+wT
S4LxyrL+qnO//NY57A7++VKF83YvO44Rpu+j9S/Ko5IUnu3pC79D5XKiZIkbCMr8
437pTS3DhCJLPImOylXot1mReQrTV25YD1AJdFifjQhzPC89z51Cx1kRsFwXYZr0
fBPZ63XA3Xy97tasen6bqRl6gXAi6aUKY46qsYTDrT5SFiFpVFMWXqBLs9F2ET6E
TeIwWtWP1MjWDBDJKmbYgz3i8/2+RO98GNGU75A72BE/qUbyVdpUiLUZue3MtGsZ
cJKIY3XWXe0P9CSOu18TH8Zho74kqpRlwszv7aIu2n5onBygBFRi0vCUMqOcvkJ0
rAumnMJ7l+Qbq2hOtq0QBROBotvB6vUy+zyzIIK2BJ5e24gJEUjtT0ukx58BggQM
qMlZ/9bUCupCNg4iG6ZYz1mbooIdkExWoV8rCDvjLidMyYo4McKyBRQhIfyFIwf6
egwpEVv3c1NbbVkD83eAse7/sRdpHz4YLrhCZ+ckzVdI8Qe+tBBdaJ0U6w7YNXxJ
ZyBxKxctzuJK5TL9euJ/OVckHIGHCF2kzUq/4sH5aQrZf6IZzyssur8zdvPPRJ6d
CrYWECmsaoi1XYyAEDkky2ic73ci983BjiuvRXvPRaEmDNWrAgtcmvbip5vDpR5l
NTZUNACHDtNPiTeqonF61YzR9vg/L3/yA0Aw8iizFo/tQ6zEtY1vhmHRRTdn8n5+
pY//UDGVgVCAAjRJVNiSf4mLfr3dQYuEGgbJ9icfig/0Fq96cr80rUNpE301VPkr
XbIv0wU0hu09hnEo2apO+ID5BgvCnr2X+xZTNSwo2cz5X2JYu28U9ACYu8buiyv2
2k7iS26EiugTwPu1HNx9U71XP9W2PY/r9mBi9vzdFFsu2ewomtYPkZHDGo02LWZu
ziBKyMgkqQM9MpfQhFJmoA9oHMtOYbBllKUPbJogZf8abDLCVkvMeI1IXMivFG3H
YzgLlNhKjx23Z43zm71ztrXEcfgWCDHqiXfHhuhNlbYK3j9i2oRxc1x8BDqAOWf9
SjwCHmFDrCqZZdnqJvaVxBfZav8BU2fklqwkihX1+ImNXwp1/1lEnruQUbwe5bGc
UTI36X2STjlh/WE6IKpbBnjOnLY7IixLTJL+LE3GAZaNkllFm+FNrHFhsmhSH1rJ
vBMSWoChg/w0iaHbAWaEooLujxqxy7Mr3HdCkRFOkAOoCwIiKu8YiVmP9U/8Wf6s
doml7qyLtD40WwLvmiCTx4GZMiLOtGhsfMU0Bj4dGmF50Q1W1XlrPfDawbgdybXW
7GgHdd4jkpq1LWbk019ZH2yyeSmxq9r1KCF2EMZ/6DzhtIA5P5TOH5sA3PT3UAPX
de4f328JuIB5SWUwn6C0oTDeyIINcIuUI3M2RqEdc1SqY/lYdFt4AbkobF8Ptyma
1QOEzwut4Tx2VhwsexHvOjjUp8oP1PJBFepK17ZgT8ndlKJ9aDKD0PQNCLCSXPQr
8qHHCKaIRTMpzcgCpY7L7zbJXm2eytXeb89EY7FDwU2ZYBUB4RbZZgywaVxjnU4B
yaCuXoorhBl0mLzD3HEiTo+mznUvooBcEQDLfnBvh/DLncWtfRZI9YB08rOJykjy
5EU5REtj1EhuOtOv3lQn98HpKTAWu7sT/2rvUH5FtRcDUI1AC1dBWVPD9Ek4laJt
LZwVh/J6B5Ut8JDI79NJtwkU5cQaFw93XDpmpgiMw1oh/m50fYcpjp3tcO3nkkna
QZYxHzVhLO0Fo5tXVINHJ2hbZo2dbUc1QR9Ao1XQe400DxmzaCPp3AgFWjuin3tj
/6EiYvbw3sfSaLSyBVsBN6fLK+ZSTgKjRbYdy/bumx38onLDqFw2XcFHzXsgfFYT
Ao3xN4J+B7Iy/7bqlIe9+zt3REoLMWQK90ZI2+cWz/ywl+gxPalnOTFIEAu0uhaW
XIZB4cN+K2HH9thN6YumIgui9PzsQnZceC0puVVe7bKDx/GIeYuTL9iFDZfF+Mki
qlcTx0N7IvAz+zeajS1REp6nzuciOrVKbu7/+QtEGuezQj+46BsxD6H6+Ra32BuL
QueciO9G6MbzyEgVPvi2LRI6JY8E87nrNUOubbH6DkXEuM1iuIAwa3oE7PfKMgUe
ExlNFk0Ne0vq65/P+8k102OQtF76lSAy0DUL6kfJMVEkscrW6vujJwf1kv9ev4mX
VfmwdzKVL83cA1ZonkmEqIjaOzJu4VYK3/iQTFVU/QZqhkgm4W6JE/CPLnkYBwSf
hdZ6GjL/DIeZC0/H6lOa2434zxa+36X7much82VLIAlbLT6rcz81Dk/P93KM1Wwi
SkCozhT77o/+VNVE1m+u0ubROzZeXGxku/Insi7QNWTMYx32EK0PmjWWz5iq+Mia
O6MuA3+wc8t4nwz6Pem58WB9tLDTwzXsYYqj2DW2/iI3uVxiuEHBEWsJxn2NM2if
A2TDyAiJln6FEo6vlrm4b8s40cK+o9Dsp5OaNWDyZu48qFvmWR7v74+MOPryyjSf
VKRqcp9KF2e0XLXtMGQ0kJmnc7u0CB+yGVqKEPeqLkLvWky0VlmEDaxST4sKrbp9
tMMuA+235WvgH/MXGbVl+st/ltRwFSqoog3ic2GzzgFAbEckbQqeVx4cZCoHU/zQ
WJ+jtagxI994/amotVtnEf6QOoL0V+RsiE9Ym0UUkjYzNhUVWsfNuUDNrnJt0mFN
iC7O/Ycw58bsWdRBqmPP3bPp5e6H5WRg+kpZps9eFRCtqUvIjzHVvoGRXbsRO5Eo
z5WhC4YXIEDPoaezxYII3mc5ugDuWVpcUn0gFzORp/Jy2Iz5eBnjz+JTUcua/V4q
dZSkwMHWPIo/gnwmBdqEq/loACn+NwF25nNEY79Hsj0hX87Jq0K7WYK6RblGIFWY
q0QdYGqDv7QlOvwFzVxpplsaFJhiEqtwAx8mKKjy0Mv/pkV8rlIHYuiuTxNOxZqh
QH/yAc+VYjcNjl6jcvDQYxSxRNu+IAK74OiGkU6L0jHskm7kGur5MOfjyLBiIcJG
k9VpOW2an69vhIYNJzAVGdIvptvDJMDVGuhFgsyhbT0rU5V9Kq3a46g8KEiLNv9Y
fzsV808scwkeAlbMu+2sybWlQ+pFMCLFP26UbynzSs0jsmATvmXk2PumPXxrc98M
iyP8U+GJbLGBikqhd3cPnFIXP1BWBPgM3f0zY5K/iG4twv2Z8WwnA8dgiZGQyDqG
Xlm55UIm/GTPX1Uwpbv1DsbDPJqZ2pCxqh1B3C6rtKQmxUFx6pyxMjmYWOp6BniN
+f5eDCKNi7P8KUUe5Gwy0Z5DaVngtU4BpQ7XR3m2aoDBcjXKVLE31nK6gmVT8Onl
DFDEMcKIS2psAM+V38ZyI1ITShgoB/02bGU0CgZtQwc4nmk9gAfsaX5e8fWPbE9V
JDcn2s0B7cjYSgl4lzX+9YezVLvVhUFIwVyLpA86qNMghcQtXMyTIA84tIi54Cgl
Yh/9UgdLXc7EfwVnxSsN8ji9GWuNg4fOYmB76qgvwe6eQalZZC3Y8xP6ajaB5OeT
P1F5JNyb7BrJXkt7cIrnwIF1uSZlSIhyiRtsZRfmjxCX7nxsNjpxGt+gvlzLLUVZ
zkg5zpnmflLHvVWv37uRrCReO9W7Mm+fZMs/5MR+LhM2REjWvLr48iOZ50z9ZGQO
9P2L0Efyg9uUD1MLMXgjlHHLFbbiHJdEADIC0Fpocf4nxKRj/w8W/YbQqfubVQah
gbSqWVJJSICwlxkqiKtGfst6eaKwhSosYIxl3+uHU2Zgpg/vJStNO01mtXy7UCAz
5dwcwhOWeJrVYjH42fLbEE/skFSRSZ0uJEe5YYfIZDJ9LGE89epfgCFEwxRufpdY
8l5gs+Jez7C3rdnKD9fgroZ/nvxqOHEvMVTuu4k4Ot6fHqt+4mRJ8S9OlqUfBfZg
KSnlZVbzmffMfZnmuA0wvOKHD5wsJ4QmIygydCIQPeUpwC3dh60g+zTYIApgIUXe
sUWRF+lDLplcB+1jaRTa+Ur4A9NDdOe39e3HZl4+2n9CL8DkCD6WsiL0/nHEmgw2
mAVvp+auifpiNfdfUKjDSinU+CJKn9U56Z29AcqORCZAUKjGiwVtTK4kkImSLDql
Nfuq/vLI7tpEpsYRR5yZRZUuLhP2umD8cCNQFl79uWSNkZju7VFt3FAwEdcksE53
G/ujE6sBu9YzsDl9iOXilH4zsNjZ+pOI/ql8quknYPNrrkSrVn4HCt1w81Smompg
B4OhJZk8vMvs5iu5SUMvPWGo9AW0xIGm7Fnlis/UYuCZ8o5Q9EoJ4FAskFIz6SZM
BjGfj/agGmcco3VKlA9hogjldEaUjU0BpdpmWJWZ+QLymHl0byiVXTLrq/chMJmw
Xak3+DQkwTjrVE+c/MEZ9Brb43kzJgIZp8j/RP4TL5n9nxHj8Hk1MxlEHuLzXs1w
vlQu8IZGpRgJA3w5w32ijfIs/Zukwe5714mZQfkw2/myFugIO7r4m6C9Dc/GMGNU
qgKmB6dBY1m22y9XDm+bJOgHWMMsCcp0mTm0H/WeFh65sgRC+FQHyMWOVfGXpa50
GsepbLVDhd5CSOM/D7O2L6qp2jyiRRs90UsB+FQZd/lxQW+tvLfmGn9rKLAa2PIL
dNTM01t5v5l8I6u0axgnE55OqbLu1b3pz1q7x7XQh5E55QzG05zRsAtJ6LKhEnJF
r6ltzTkmz8Y5UFVKJqQh/+nfP/gnbqvPi5oQgvZA3OO50bbnSoP4J2X06YKdzxDr
u2C2IAAB2RMJ9+Igu93Pt3a8OQKB7YqJRWRPEljcCkNYXvdQVkfiB39xcDGmHhPx
TfejUxJQ7PRglY6Ze0DAC5Dmqj4s7bTpch6kaqRB5Fwr9kVVEpmtPQzCVMOG6Dzs
sI8dqBZK81z0RQaQmJJGPEThUuP9ptInk3GeQSVexNc/rL+bE5C9sgOwLGBR/f/d
kRt8t0nOj6QJ6//kXzLLBNQtJD6ACahKbcV8JSwFV+3xMqmE3NaeOfr2JUcMfQCj
kx0m91Q4z5x18dg5B/EsqNSHqsB518g42m3j6zD12AaBd/guVVvRiqKb7JFfRx1F
bisD0on+7/XVNqKGI5inS+4QWW5w5sZQ8+/IgltlCB+O78QBROY7z/vepDwerMPg
uTt4lBzPlS0YOV7eNb62IjYT/IHPEBub+536hSjrCTJhK5dFfX900ejcneMgladQ
9oDilWWyZK1KFNrQha+nhxVjxYt+qvXCZlIyXvEG6C2NQL97/1tEt1wLNJEyRwDq
PFL3wh4kklmj+IUOOPRk3LgS1YKqYLQ5H8F1ggQ9nEUBni8BVd/c/XtiZYeJeQ5s
dWSWWDTza3opOuGHE/PfO5tPdayGNXOKgfbKmt1yHyCkUaizV7PpgxlG/EfQN++u
zfmFKRP/xmsJUAb0I5fZCP8feZd90ntn91MJYpA0a1WtXZ00IJphhjxTQdtDOeO0
k7N7HNwERUZZrdetex6tSg5sAFAHI5sCc/U9BgC2QXIzeSk1/7A5gWxtd1MWJgwr
8L9YiIF2PCJMK75FCGTjgEadT9Edbgf9UURRj2PZGifdu3lE2bNLXteDOQSc69oq
B8oS6+3TjJriRmBheaVwgVk8zLbR0uAlHZ/CHM6oI69rf9+bcASokF5XaLxSR2eA
Cue8wA90yQItnR/8cPGeXQL/thkb32EBAf6XplLTO7EUpVl1Cw+SS+M+bZvvgYGy
VUkrDR+7lZ7SDV1yjZtnzRodmup+p8TBSWY4/ihn4ak9dQvDan7ZeCTfo6i6aj/6
P0uXPlM+nvjS/Aq+tOe+FpCJk2NsOHjWBB89BB8xg6zBBFkMRSzzj6EjFl6f1ufS
SDL7wKaEgyJaVIlMcVsmQ7HgOfx2vgAy7PvFBol/Xk7kNrzBq65FSYzFDmAGhGcP
sg6UK/Wel4MVNNmjoM0iENG0nHjT3HdNCYDGC2PsSdQC4Q6tI5F6sUBBkbBKP0eT
7jMTXIIfZX4jKxgx5gVrNdH20Ejm83699mNaLQqmNKeZIUyAAdsUDV280A8U6xyy
jeqT+q3QH2vz1NweyM9S7ELuLUsJPwcNCyyFSaN3o3sZwN66qHZURnzukq3CL6N+
mQTbstYRAsqVG/KXAU/iu1S9kugmt5Ix1LRJOaNX4DWNGNE691B6lk9TB3H+Y/U2
QL4tFYTJ7SDML0NIUPp43Y2fYurgu2TeXMnjsD/A1S5hTeJ69MxERCQc5D06Sy3f
Zvg1VGhFfkavmmMarUF0KicAfklS8L2+HkIKAN8BHidjQ6frq8EtU4Fb+1IRDxgR
ntdg82dTDryyFW9iIL6ZG66CIURcrXImfMAvgwX91ciUwvVE8uNe7BKdGILBbH+v
Nqx5kyIrFth5sT1qqXU/OFHIDx02wKgDmh3wxOBEBheBNgclKKaKnPyAM3Ntz/8e
SS2oU8H2YM++KrtkSm5VqAJS2sSYODu9mBh13r3WmXd7SHXNyp0+J/v3VIPhb15h
BgTYo6MvGzpjiBW4Vy1qzsBFTZr07dHeLqeZAm5TxwrWGuo7RSwt3QTASLxk9wPR
NaKYYwy+KpaJO0N/f49nsCogPseVNiqVArcrAHOJpaZK4P+MSS5tcb0VmBan6GKB
j9OoGDDaiEx2IvQwPnFd9kw0veXuKhiTryK7zIf1B68sS205AYrZgYoeQyJprzPy
T0sM8qa6scmPT/BRF8wKxS28NUFyfCxaqqORs3Zco4ur+twCXc0ONXWQ432SaIZj
TS2WvF5AAvONmsO2ekAQpBhk8cDnm+femmOECIWyKPqfB1pkixnbwrlsQBnzkqqP
hSljGhtUFqyJi7NwX7zPhGjE0x2kB6NIGw6qi7VCH677lTV1sBgADHoUtd1jsB8O
LEhsVVSjEL5sz9fWVfj/tsNuKmwhT4QjkOYsF0xcnWjFnfe5Lm1uX8OtHdN71V3i
eK0bwY33KLgdTWUTvkrRayZgWgtyVOZXeSiuoVnXjuKguAziXDF3+GkIla0qyh3c
VI7VDEqVQ0WjgL/A/trPBxS2GUZkVQ6Lm3+Pqc0KvIKl0jhuSQpN36REXrYcYM4O
68wia6bI1zuaCHN5ewHpX7Ns50c7Fqo+ObcuAINcjBhDJ+5vDL6xkhotneuKjFaK
uWM/4PAMc1raqNTMPapiBXnaz1a0+sxVV0EMwdMBS8R1EIielLfU3fpYCOJXZsEA
OKvgGobTTjRiS2MB5DnGHPUrH4YvRL+cDVnfRQH4NhYtCyEhmUbc39YMQlKDXyD9
CJ17c5OKRYrpwHWaVSuEeLRX2borDKJL3ljHVEA/c7I/pOhpvZ7G1RB275Mpr64x
pr+iwGzBM7Ki1ZwDdRkDagXNTN827uiEelNvkDJ4oWeQMR6Bwjyuv9iXwV2uy8uM
xKJYzPmt3+czAYEwXkGqGIw4thviRJj8zIoCPuaXG/UIvmDVGhO822zKLvdRvAk4
fBSWVeWD+vHKlEQKGjVXMqtKE93lCUm7jVRl9phAbJXS0Cq6XAR9r9x/AwC6ltO8
YoSR9Ls+m4PluQNwsk3TKYuY/5pMMETPBarEQrHZz9IElN6SRCd/CXIN4lxuRTFM
iYbmcx5wq8SNE9a4tru3jTLEF1bCuXvj8xhAbOMVArgffc6iFR7Y9coq66hxXiGg
ka6Qe79JbZ4f3EiChSTg+EHxjnbzvOfR9ixBR2W+h5FvFbH3EskTKI1tQwAuGh/v
A5du6RxenT6iqOdoOAtX9i7FWXnmCTuSk3Btvot9smf9CZxVZ6SaMQJoB0r148vg
HnoCVmTyipb8HyXnkLZgLEHDIIPgtMRzKDxlnonribGMZ77Z1QqfnJ9P9i+ivb5Y
SJrTsxy+oL15rx73kD7q6i57xgX3X/QAfCKfUQptl4MPFqKitywrctb27YOUMVe0
UYwWypMbDl8oZFzI4JAhxPzvTeLHEypuv2bCUxwV74ArSFgpDy++q0XBwpOfM0bA
YaGNKqE1Y456PafHXzKsvmDaxWxzWTBH+fvA53QMtqxJMks4ZRFGGgaWrWr1MPUK
j0Vwh0qzcWNEHgTKS0CK8Tn85GXtH0ErDgwi/LcmCbNfQbDwwvbFUfap0uk3dVxS
D+twZ3n/QwFWxthctvQ4mzRDyyacy0o0BpHHTXAgeZtoj6pbwIuQzVH/IFWLTj+Z
kKhMgfC6wZRx+yxv/AyOdogNbj/cBtmemdWcmT3UPmeAVyF/b1SztQvn6GpKhGif
5yoIu2xrtNRDCex1GnsYtMKTuZZgglodoWUOdebnabMkzhuUBHeCZ9NzQJddovgz
a9bIy+i8rNC3Kv9LrjZCBVVNjaZwVnlq4BwQ9Vy/Z4qhdtFRgeYvx+rXs98FzwkN
u/phdt7UuIwZxJaT2Fz9pJCHTL8ZP5eVv+vanY0f2g94ymPVNwwFCWYalOdPdmBO
MvyvxGGcQ7PMIu+tkdOVHwBUUKxYo3NMo8veCBcQbOWJ8bXq3KxcebJ0wdrUiixJ
qILKTagZbCPGdGzDDAJLyKJWakglRmdpL1n7AT3k+n46ypW16L/sxAk23u++y5/9
vk2oycmvpY+rmERyLkC0y2z0a49Xa7nx/tPutWKJfVZ90oSeoE+k6nWvUlZgUPgp
KGY3py4KgHtXt5Fh1IETNJK+ovicn12K50Yyiz5wZyVnzPg27BZbHN3oLru5SJAd
PbH5EsQ8TnpOZuKEmQuZ3pt405g0Z/37Jee7+NdjEVViIxY5vCIGPHKfO6lwb58U
IzAC6M9ugm7eoYX8I63eqBEkdXarvLWCd+hIuoo2x+/Re6ce4ZD3eRTfKL3vgWi8
VwSKn/Sk3D8UJrl58YzTatG+adjGsG82gygdc85ML44zWIzfhSHTHuv1//kG7Iky
CZxd1hX/5Mru+nMfrsTQ9WheqqapKkFNBpvn29dDbb6J7h3iMAHCZGjVo4+e7oBq
eksH9pYG2DopF4og0K0wMQSf3brsd39wt94gmXF2mHpRzQO7Q0ZcRd1DOVvMm2sU
b3swT11Mhxsy19rDr/Cd+pUINZwJuGGKyyMbxrAyCpmdUb8wF0argQi8GTfoILua
ti5FKuM9m3+rarmjCuoQO8CSy2lVrzDXpQJPz4WUrw9L+1n8Yg0WRv2H3uvRLWvW
eISlUVlPFbXBV7lW3BZsgnCPhPaEmO93IfAbcDONhY1YAymzIIqZpMN1qhsrEahC
S/eJoYNjeVA/k6+gjQ7yB7jkcohknNsInvTNgxVHHt7wT2p2/7m9vXma1hDCPmQb
JirmjoaXD1qmW5h/y0R6AHF3oK7qHjWUdMBwHev3XIZUzGBrlsgCB12BSMvs2upj
50zel+3xZpocr2rmqFr9unPz1HyCQK1FasDJvwCaICdtP+CTJLH5qfVF7AwhMJ0q
vXm3bQrbsK72zrFV8iNLyfEx4+LxnfKnf1OmWknfyGMb/Y2NeRLxwqmpO7zSXmLH
1YAbPBVL2O59Rj6MZCUfcDHORD792fboIczaBdhc2SSApuJFkHb2X5TNVTDj8PCN
Hxa7qdIb8wF3Oy7dcVCHSxLcZAuHL3GeefUt/c4VsbvRaXbBLlUCo9mb++c7Kcy3
gWeFrZWxYEfKPd39cgCo6CnE6S2GUZCy9VsmN0TrBihJQM6dAm/uHCFXYsmCDuGt
vrSAr/QFp3f/CYpUeH8QZcF3r7MiDnZfFY9GIYU0ytvsb0sKDwtdpeQmNUeakVUX
S0oKKyZ0fV2nRlLfHVcmI8RB1MZA7xWk0SZKulnRJ9O22tQBd+NAobLxFHHLfb1H
EqcGhp3Cx4iJA3SuTXxdDBvFw1UFFZKpCVDJtMStzLwXOHqNgFoYVVGhjKY+BA+7
vcpdNR9ks7uPHTaccugaJVJYxtgMspFt88bZujPOZUAp94RcKekH+TnouJMoKQBK
hCiSBk41IeIOQhgHscd0mpRB4Pu/hohMa48ejW7mqglZ/OsX37r1x63EMBgSvPzv
if4RWHi/KYuNL3Oo9QX0AIErXal4nkHd86Mf7jDK1laZNWkhSoK5ANPgtS5SIJXX
H14AMc32PgaEKIuI7oFeu3s9ZCJWbkvFzePV5izM7xhCjzbwp9vQaiNgpW7zcuJJ
C7Cw6utD2QYFPgtET1ywKYs6sPEeRvSERhlCubi2Jx/genzPd0rQi885tdC6srMk
F6DSwDKrju3WnUgM8tADhRKuhje5XiQMwlpMN1ZqNPYj+kzCAsJ4zjulRQfUqjcQ
7HuPwpHE4TuZue3r8oJIpOcar/3JqhhT0tBX//9Sx9ayYySgdmUY0g+mlltmh6sf
XGsvM4BUo293soL7jX3VwbVKfFmPuhLbQwyFsAfWCCz+/EXkwJP7W1a6PECxiECZ
fAFME3qBFl3JDBOM9zBDr1z8+m+NqA/DKQaIb6b3kgOS39wD9iCyBuLN+UUbZWZX
Uuab2nSGZBElLUn/3UbQnauD95NL+6cNTVysCVf53Jt4cm+7er8s09fuWNA/+Te5
9LN95JNgfSOkgFU9MkwEFTBA/kH4A+6HtuOJmh9Jfck2lhEI0w+YItnkM7Qgzd+L
MRKbDwhPOAuxPNVX/fwD6qTLKjYmOif4k45w0eANugbCyQSn+z8i8Zb5qoG7Skj+
DzcibkIICdYSlgcHgXw7nJFKaYKjba8S/0f3Z2Iyf6ZNydn3jUT9YS7vl01A0miR
d8QiKZ48YtHMv7UOYCLUEqBT4LtAM6Ag8qmcNwGJ4PRmHtqvPGhUR7o0AFdJ2LN1
KXTWq8TR1ztnYxNsWkpW71hsJln8rXZfBtdG3mJsjo525mRywB3x5Xy+2oAOiKIZ
3awXPW678BUgWOyqt96xiE+2bERy/J1Q0HuG5IUljmy6ISKPrEc2PWnrPjbaNeq5
HI7/5PnYHCxymgqbiPzDhc6CFUmuG7czKxBnnMQ+b7wpFJ5BkgjJ6Ky2t8YvHxGm
9AUCKwnEj3FGKj28Py/P5HwKHclbfJweS6+GYW/TsnM+lo3LLCbAeqyDs/A+Ym3B
VT3YQcUk6pM+ZiHykwEcIqw8v/vxZdHaj1a1Q1H4WlV5bahGFsJDSrQXcifsomuT
npDnaQEPVvDZBwhY1iBV2+tpYwMNsNpZzM4mxK/4fo7bFpBGXa1zGRTw6OAEBMgp
JjoWLk9lkjdTjRD5LjjyxPuENCFOivVM0E8YqcnhhfCQ8jRqrOC+HleEsUpIb4VM
nS0xJsVjPIgmaqvLlADQWkqoQywEy2PSrn+IIbADOB6lmQbElRXsMrwKNwPZNus9
cho2UIrbRQMfkX97GONHB31TP99F1w1T5xmNlh0ueD5G5nE+nQfFz0wjzWl8jTXn
0kJzXuKh6e8PFdAk0VBiNHpRo74v4xfaNjqc44vOp2zbTI0l+SLbmBNcRDf74447
lacxaMr2KN9PmjhO+ZzDKZvkLTmJYehVv5ezSgxqGM0eYol0jvWWz84yCEVXPOZo
0iTea9/mB9Qdy2wykR4AlhlD5CwFniTSDjklWCDQ+bJegunprnxy9ecAonpxn02l
7yBwWSsQPdahgMlE0rZ1HbJbQqBbo6qG4BHLCgPlfzpvh9fR4NIlvJQEpqwo3ixx
jDOZ8XJAxbZv3JoWLA8BrSQFJT/C3JaCsYIgMYy2fAzmI+/onEX3RA8Ugdlac7zO
GmBzfo6VzPe4ZIFizEPxy1SDnv1WQDntyt/X6RC7N6Kla8iCxbzj+4GqlNXCyhOV
pUhjnjBwHP1tA1qZE39vIDBCPTxj+E4UBDF0c5KEM2vVKnJVDSWLUP87B2oUE9wm
Ls6g8mhog0UZ72x/uZR2L2VUIpXcT5TmaND6XpjSVgLsdLzlkLruuJ5qrrx5EaK9
FHHO2/UgC/e9g0U+jjcFwD2Q0EjG/ZOuCkQtEyrIVABgaVUtmob3K8ErrbrdXR+3
sVfReVSo3eDJ2/lchHPgB61V0Cs9p14fJVkthWTB7mKLaNkwZ6I5F2nMdZyr0vqO
8ew6IhnvLo8Sen0FGkheyK0DHLw+GWAasySghdh78C+6bVewDJHUOcLnJJwfMKy9
rVQiKQi11HAWXjdyN2e4fmfSKFeM15aoL7bNo5CmVGWPMKJ1SJGwCoyiEvpaYapH
fmKq4sGQRP4ESYIT6+RNBXSS7lbZvE83liSp6aPKEbyU3asEEtQyB6G6nAX6FksB
u6uOT1wqEJ95p6S6KuIeaukyKtU9xcJS1hB7Xc4s8vwE7yeJNhaH8/bs2yXSscKN
Kwo3tQBOgSfTvfiNB08z4jxSc1hdSMX069NsoCEvExG+yuHm3M/ZxFvKj5Eu1Jst
50AM0Mzlzk3nbPkyZ4Qld3JJYTdAVaJ1Hnd5c/GrLmVNlUsbNHDvAiYqHrZzS+3b
/MKb9mnxJRW2L0f0xUScOmWmITVH1q5U3eebu5JsoGrDN/T17DSlXtQ4rVHad2K2
Eo0tdhK2XeL1WcgbsbxNN9sfmjA7bvbd3iseKiS4E+T7cNZlCEmr1eo2R07qalVS
VEJVL40c0xdqld5fu1DOgZL8J11SzFF4U8ovJRAmKTe4h9F1uZgC92ZNWp3Pi4IK
rDk9IVyMSgKrmANwBCnbVkbyc2Nt/8bOfqTfAnJSzkBtrBAvijjoORC7YKqnPULV
o4GWMY/Xy5XdOhxoKwmtc15kSbc1gV0x9DBkA8qJHk1bsCNgqIAUACALFfsQPke2
5h/QVmvW08fLjxko0NJRFSC5EqN5ZIYeS8dCBDq7qaCEd2/6Bs95eOZnUN97zinL
H62V7P8p/mpcbayedCpmI/gwMUqehf355pvF3gVv6EJIwwrF89NRCenZfa7qf8dx
KwbQ3E2bRno4ERVcyOPWExCDjG5qXntjgF0rKYNhMzCn8lKuLtKFIZRfXViRmGUV
NmoszdAXXa7rPj9TbDv0eJY/samvQuHxXlzhk02VDe854BS5AH5XoKNZDW2PST+P
W5J3kbOHfnzfTulMySrraU5iuP2a1nK17GjP8bKT3mpA4YI/MuruN9rnE0ZT9f8k
mI+5APE88WU8ehrVIOgOIxADHAmb3RY1GPsuywZCRO/RBzlLjqOayklpcKlWBsl4
XyBgjc0w741s16Q8VCxDOBzg3rK8zn5jb9NQhK9bso5tD/oB2+0dJh2Tkv96G8si
95UHCzj1nxIwCUQQm5rNU/RcHd78BFQiYYRMm/ArsVHpgP7b6JJ4VUytdF54PDWj
Nzx73VOXHbKNndIWw5AJUD5bVxQzBqot69bhkwCjdNc5XaQfxju1i+3XN9A97//8
7jUoZgw/o6mcg7liVrWaApWqHKlFQJA3zEyHeINF89QDDyWfoUqGL4G+Z/5l8aNb
tO0Qf94ymzRHyIQR9EsE9EhkIMMPgqpjDkbGBSqdyFmd8fP8ROgm1TR0fxxoVJNc
miIzy8cGQNRjrVtycc1a+ebNUiQ6I1Opo8XA7zTDTNRL3FQVPgpiHnuw/gW1AMIY
kzXSZ30AR/xxzkaVxUVzd5YamcUqJrUpxWSDbKsZPrs4FVz7WLT53m/YsBa4shQ1
xs+IQjsrcYErxHvwSYp1RPb1sXwneWkxG4yi84ucqpBY/xAhzovXZb2W7kGwkqae
eaNqeGz8uq+3390VseGMvFqqolUCgJD8cIPzxEQAXHLnu4tRN55O7oW4IBOGJK4W
fFN8Vh+haNzE4yHqLKa5fSPeatgsA5PfhzJhc9DtQkcQREbBQmFidawz4bReZT08
QyUIIBimLNpE6rQCbAE9UiTujDfa5saf8hGeknXRzLLcw1S4Vl2DC3CP3eJXOuXw
O+p4MLwDRPWbxN8ePj755KQogYUASJqv+tDwkNzUqbZwVupxvngS9s+allRzh+D0
5wGFYOjBG4ZNDb7Nt3k7X9sKsgbnIYaUhvTqNldNnWZZOeDR0K6jnNp6QHn7uv6O
2Wnp9EfpKIuJD0FzXblThxVA5nGu2mAVI6X06b2EmOPcn51lY9w7h4Obm08MSNqF
bAoBOWxClkJo/u6fUvUDAnbvCuu2SM1BtWxHHN4ZEDtb3NE8EL9PadqtBLwUI8cG
l1fa4MXtHpDzl2D75WjRNw99LQx8y6HX85uzCiy0k7DF2JNum+7XYLPXkh18C6gT
HEAK3ttTRvzar++iHF/o/LJOmkAzLLyOV10JiOAsqWgxkZ52XRp51BDwOC+ylvcT
EbKNOkz7A7BKL97HvZ2tyRxrEKI8mAzAOc8dOxe4vPrhu7O7pW6vWEPaJejdKdk6
hA31nvbh8pPtENjA+B0hyjbJzhoOH3qPyRStM75wKGY59+iKLWGfUUAxcWGGquEk
xiPbTFZrL3RYONWVgFfOgBhKFA0qBKcWJGaNAtlnqyI+EOE8FmySf5vvBDXHqDRR
Xtv/1Iz8gK/2yMmCb2vKeJUuO991+LAzf0DEDWXZWgTQdNVKL2yQ7H3Ktk9mgWH6
byZrb83nXoXj/TBeRnyCMQUcHVWdGTGNTAzN/NLyQAgluvnDweIZYneYkLizZK0M
iXBCKarRnEnxyFvx/Z8qAZ2Zx4TrHPu6KcLwQK9OnYENktDf5/uUtEOvx3SqH2Gz
9gvwdZexMiVOjNQRmZrdWIdwFULMu4RFkwWXp04Yv84SjTa94MnBVAo7AldvKdBu
uA0UY0f7EhE7sn9aRaDKVZj1tnNbeomNcz3i4V6KJ/VQv1MLXHEtNTqFUjA3P2fF
tKfQXOqFylaRTu2VyPgNIR6c2AejcIdBGoXXJdIapSCT97SYayBebtv9PxuPj03w
JR/oee+CDGaOtiQd3mzI0gBNsnmurIozUs9NWDNg9JNf+NFy9U10teyhhjkkYY0P
X1hpZ8fA+WDgGvxya3XhqHXpc5DWhczVEyKZa14iURuu0ozCrqsvCVpRl1nX2B8t
i4iKpMjTzJsYiJop/zsmfO4a7pEPMaYx/xaHVFHbbxcLfS96MakfUl4HwV7DDMyv
11uefNaFJN5HY12cFtEZbKuxUIwjOJgg9LTQQY3GR9XgYlCP+qGrBpuSCM3LKCgM
6GwSXP/uvP56VECoxGBCIgHRYv6Bhe/qo4H/9U3g8WJoQyRVPc6cSLQaVequdjez
WIm4yePRotEUjLkCJ5mexeDOKX5UI+gJxyjHWGpTQmMZAxMC5OyDOblM3hSJzTXC
87YX2UfcKtPjPCy+rsH2wR0Yt0yd2+ljUTiXWVEwIuJ/WBuei+ebKsVXy2eM+H25
yVnIzBvA4iM1zcvupBM1eWdXyXVvzXvSoSUpJSMBpkuPJLlpDMLSDKC4Iddg0lhl
L93U7K7NzntXrXa4KEPVXWHXkjC3RvlJiXKONty49/FIvtCohlsZvy7cIUfGL3hq
QOzLEki5X/jW1KKEVzwq2yiYhNgnwTYzd+8n1gOHrKbIeq1Rqxi7K1oWvUo8q0CO
WYMmBLU1yip+k71wERD+s6HhvzkbIUiM1tsqGizIMYiZ04HklRI/wAXvr3xicflg
ae2qSwgA1BiSozVOP72sDDGg6kctpHG8FtKizp6UTBIQ8NPjaG2RLGYaNPcFBFMR
UgDc/m/A5L5qjE05Os+dwIMFTljkopayxURxMmgygaOdEnhGZBFiBdFGXKdJwq0D
j6HPYT6cVGRQfzIIrAzCChEHpw2A2xNntovgmzj23mfkSchZ/8Jtw/mGI/cRfvA/
VSgd7O9NW9HtdIfYtTwRS5WHIHq3rCLSAQvWHkl60JNdKQb+XQZpa4M+0iTqsFFM
9/FeNL8vOdBjwh2eraZoBXAO4ChI/S2X3zzHq/ZfgPmkdm9LNZSYA3EsNI/L+0Gy
D3SNwztMIJJOe0WS0OQITnzxzfRtmGPKFvUdvrJHsHYwm6t3dmo+KEpw8TzbHYd/
yGr6idkp27UxmwWCFd0zDe1Gu/1Pr6QzqzEJIUvKQGcFr1+wEgvxj/Z4+58fcsCu
Pjp7+7dgkDI7eHc/fL4JNVaMRyI4g4uZfCNDLyW4Id0pV01KtVTYCzxut2f+eE65
6y1s/zkA1N+yGZlVVbc1k3HKspsTuwBo6ZysrZmDG97w8UL5e7thHUh4ndgFAiHx
i1keGJkdVKto6mkhHU4L9+kItQOYD9CBNNlOmvpCIqXMzyX+eFc+Rl2qKM/RS32L
B4cpIL0PPffmxfTy3ZJArYbS23aLaGLVHGZE46GmNWZXtFf5Kw8BtZL+5iJn/YU5
OfKZWUo5C0lVXOGxHwxbZAjhkdPJVE5MrhztV7u/ZVgqJSi9860D+P100sGI47A9
cOujfQ6IDe5twpOc4ls9oNWtxPVYMH8N6fGce6/t85N7EXk0w/hh2GnD5z3uDAFn
2jK0Qj+iF/6m/VcGRfvEEFSPenKPwlkQyo9KXW3cw4kxlnSjx5ilXDGADdQ86zyL
wirZB/srdVVeE7JFOjl0O/hVpkUqpZucSeMAjd6LKURUobFCDnqiLPzUa+UMXuOR
W2epPtgYvvXvUq0PCxs5Z3hP4mxMk/iAwxQuzAqL5WKmoZX3PQzuARFgwSBKZ1cc
15/0ikS+QpNUF3jbAE+m9ga0LYQevOfbIAp56+RdKOQG3nAS+xBXRW9GiFKeig1X
97tJ2Ue2MdrnjMqZUBCNCZWJjM8U/Rf/5fpqcyFWV5LFtA3II7HqsOGHTgI4LHHe
SvwtSIdhdk3ugdNvLblL0iVytRKQYt+kZf75mvsL/nRNZnq7n35i8h+CxDcpT1E0
OECOsOyZYqwATwZvGaVv7o2Qy7QO9NxRmmrbD8YZp7zYHbanrqeLDH3V1Z0XLWdE
fjc8cof8LSW5TEZmgnp/qekOuvv7mjCyB0H2iSQi+IXxMX5nwrZ2HZXftnly0H9t
T5h3aWkpVQ9MGwCEZSIkb2G/zOwFegbUCO7F/Y+8eRo2bQeCPPz6Vo23PbAHeWGf
juR2tOSDnbV/3Fkp40L31OvFrNHGkifVwgZna/1tc/AcAz3T3Jp5uPiC96/kDMOV
m2CXqi+UbwAz5kSHELT744WFZVsIZEFyf4GkyP+S9v1sFFJHzUAA8xjzpSu4sIyj
ztor2CvycZUczAEyrnGSvqjyykT+NQKnYgRAuygmImVA8M6nh/H2pAENoNW5pg1q
C4/kKroxxDKLjjSe42T+H1vUVcYLw4xYIDTcsRwj6uSAe8LYxz/xQlOoLt5tH74/
uiWvasC26lPSNk73FmOnJUSfeE/vqInfCYq2rHVgRVJT0+KAHRnmdhQ3HXqBjzpy
QKs+IkhOemuGEjvXEUfv6+gt1tw35UstqTwFx9VjSGZN1AckBr0CO9E/GVmdgx2z
N2WZtnc8naHsmNdUyW7P1cwU3lbZ+8VfKKUTnG11ACDPRdt5z4NaETOGZXhhMET9
LTYRxqmpyX5Utp3deAxp/lcQuGkbQ1+N33IpBPrrXfT3c2zUC9M2tSQTGipCoEY8
407+w4laVrHYip+en6/L4TkMKadT+oYdSlrqYifMt5dZrRPiKPq1o7UdyJRr9EaH
ecTedI5DM5RgzewPxv5rF16479rnJIA11H0lRcfKopPimi4sZ3PGgjY6ZA3bbxvX
KMAeAo+ODsl5k7bw15VvVd4xEMm/2jNfiijgTqI0WGyPZm48mgbvFxPZU2YZZ7BT
xhjEUZVxoa6VXNR7C2z0E7slAl0YtyujX0D+hOULiEMUIG1EtrwZOFqpFxAuwB4b
TPhSp1p9p7en+9Uo1Acazsz2FsE82cQ5jxenEeVBlZQFa8OBKS+JIRnaUCMzE6HD
SurUnAU/opJNCCeI6dEgHSEP3BRflIDfBu/3oDgf81usqyO0dspuM97G6msKUlvT
S8lnzDrihBIye8XTme+RRI2T5arrI1K2M/Sis6mGRAAG/soEz/KyKzJ/3mGIncnc
GlHwdHyEl1Qj+EfGgCzKJZBQMYpsnUPoF8bOLEdDIXfotj5o4un5I7Vcs6h7NHU1
zy2uPV1coPu7C1Y6Uxl1QMQicRMns/sF+wsrEF46gbHTMAzObtC4eE/5h0dHCReN
uer8vLEdeC/uy54c0inOhGRy+RhG8J/uN9lOfLxLFV9EovQIhIxWuhrK76sBj5j8
AwsVdqOV5tEziiwYFfm39Nl4BUhYDoXrhnb/Ow6eGZLJh64VzX0Ci18a3A/8eQZu
26rpO3qK6nxjDZSe5mbaQ7lKfU7Jx8cyKaQcSZosSLrZ/nsvoiOIwBufO3eJVh3E
MVALyOh9WWE10Ao7y7Qy213aI/P6XP/LjiGHMG/D54LTgCoUu1dFxhdTRnzgjzcW
2M5JyrnV1zY9euvyUy6yl2xx61SOWdqk20paFaGXbUgW7v/DH9MBsd1NW3m2a6b6
5EBk1vVZwn4L0pD/w1ZmJ2erJXi1h+1OGMc6ts5yI+K453gdv8UDODYllk1tIcsa
cio/PoK6zbjY+ALyfHQ8a+6mwNd+TCDWEKgpcXShssUOnal+/n5iMVbF+mhmgmS3
JHfcSvDHjsiEwfrh64qOd1jzcCs3m19adWpj1JKsean/DEIXCJfb7h0/0jiba4Mw
N8WXirvTmx1m9XAH9piYsUPEeQ6ZJB75YV9+fVnSo2NgqIlInzh5dcGgtJhIjqYp
boLnRdy9brAqn1U+KmgXN3as6e62csCQSU29FfSrgM2x1ztYVRyVGm8PheHP5a4J
6at0y39RPF4F8ZDz01wHCraO2ArD5htV9tsKtKiVoa5/0wUnzxky5bC/MM4OZPGM
usc+KQHBKkeHTQB5gMkAKrWxP7rkyyLJIADBD+er+5Rfs1HMZPTJcUmgkj3cP2PU
zyBhNvJAqeDG48CZGCK8QD3cDi2T5rdRu0GIEJHwHFis9yh2NNvsCf1P+O27TA7f
BzmficxIckagIe3KvwyEgbeoIlxXQQkuozkg2Y4xmFSu+didblnoAeaafhF6Rs6l
Ad10njfhlxjlKxNvRLTfBz22r1D6aW4d7lwAeu2etyLH2lOI6lIEesolkQMCVYqD
2Mr7OLg18FA7Ev+w4VplDVmLJ4stYqniVIM4S7VM4EjtAFcfSmZa9pbCMq7Mq41Q
RGWHifNDZPaTCPo5ENvvvtnemIVXXJTPzAmCwhjUWRIXvpPdRt+6/m4MkMznyEog
2nP3ZgvNi7u1Fn+r3X/JJKNGP8sAKDM0nyCyNkDqbfnJl9IViyTCv3MkPMCdf3X4
o+VsSFAy+JlhZt1g19mSwhBBgtziulrT+/8SKGItCRmPC+FzsXneVsqU3agmRhMB
/tCYyn+TeGRzqk5nOvxjZHXmUsBysDIDgFX2yNC1Bj76tbxsL+lg725riupdHl/2
E2zGYU+yGbrzdUkFtC/bJ/39Q6JJl001WXruud8AWBGRdNLNK3/mcHTSVbO01nhF
oa+oEL+Ae9kPHw5kkct60KTaSqLAbzfZKQUW7H6Gf3+WT0IZsIC5M39qdgK2GXNE
NIjE4rIU0i94TT8HXVCYNNDV6/SVXSkTrHaeop+USVXLvTq5gCj1VpjVSe3Lk0Cw
ewatkz5l1rxyZD6FiMkvn4P2ZvfPv02RbFs9Gr9jw5OuLbGq1r2/OYXIQT7jA+Sc
uTwTEFhpyPu0XPuY1LpUwLM0ldfzzDDQDkxV2Y73JviaxAcISRKjpAh39FTsv8l+
0TrzT0tNyXObiJ1QIALH4eGsKTheM4UddpyUrcfi38zeAbGnLW1DvNf+nQNx9IL0
w6Gy9Oyl6tNgjSDU4mcsElb2fkj6s/6jQKzycxJWts49BIw5GKwQ2s2zhtqDPbVx
7iS2ZcomVtmXLs6+UsAwLryLNVw80yoYYvZutdwn+h0KBIMEYSAkB0fMTX7WLwmz
pfTSRs0aey3hBpy55XcOKgUMw+KVmrVEaRlI5QQWvjS1CETcdlwKMq2a/uoyIoxd
F1IO8YGX9awlvnS7L4q7+WOShbiBSyJ916tYw2QGxskCDe0HZeSn3ix56ExEXgRY
HVVmYOFvU5t2ZSPaXwlu/tv57Mu5w2rJReuJFQvWtHGNhTc1ezxS6ijEAERv3LSR
+xfiMo3tefaAm+1AwDLTFIvLXAyA7acKzZGvWY4Ud81fMV9lALyHcKGWqTWqm5LC
CUo/XS4cqIRR0jUXXvtBKQ+9qaUHKTx9RZwUWLu4lzj4n014A3J45tYvTW6tFekC
qlU76nPE2k3Tv2zj/4RFHWNuFTZqQi97B/zdfcpZwrbrBfJrUkPoYALZIQYoo2ZI
fEKH1hk+kgFr3aRG8o16i6x1l13p7jmL9MUfH01N+LEPLZiLcA89fVWWtluYdn13
GdMxVZHk90QGRu6Sn2RD2NStNkkt2vcWJGQz2iZz5Ul9gnnUdsPwpf0rzTz9+PUn
qlPO77dGnD3TgnxjK9LJlGcl+5HiOHqGlbdHtME6JSY4NeWjoxpFHYioYp9xhijs
9661hX9bY8I/Ctvxu9c7i0wMP2S5Cx3HxnnuKKCCA1zUreQ7ky+EoOzLnCsXa69B
ZhM66HN36KAt1eJhlsNkRebxiZMY8o15/gxWs1drHGKlRCS2pzzicSswWEO2Nnsq
j8vfTrsAhbtFlhC0K+pKRPfDx+Iq/4RSJEaOJ9eNlTCPiAwwoyO0tHYUEmI5z1eb
+MyLmcUa7tla9XSA6NFbWZDrr1f3wOM0ftlZFG4GAk17ydfdb7npnTiXnb0BEInG
6FmwR3tbnGuaGAVT6Px6t9FoMQtf3wprsVnf9pP1xyjEKUb30yuXPHdNMV7sdfkX
XG3dkKBJh+vCY+Y9t3+8nMQzhd3IjGhhSLZFJ21qNyOTGcI59OZMu59EeyfvIbVN
q+738xpvHThOajV5PouUkG3EnLrhrlB4r1x5KjmeEMo0QaovlgiAj1TiNp1E7MYD
Sx1bW9/sNtSPLO4R54p5BBLisL7/xuqU03NhWXItpASWlBUdfnKb6gTKftMLfpv1
9PP/zw/H7JBohnZwNTESxjcPDWP+wvAS9v9RINIL3lKKMsq8W3y3Bki+4SQrOJkX
O2VlfWKXerdGELuB/dKOABlRatX+dTyXnl5IfLB+BBOzIqmXUDLg+h4u4HysBA/r
/wRWaWFmeQtYxUjDUoUDISFxfiUqMPHPh+1eY36kev24d7s2WNOrvAO0a2zSLLQo
pR2ptfyvfFa5kvRZcdu8evbI8J7oaJKl3mc0TaZDgGrABEZNtZ4Rb7OvWJBVuAjE
jDgmM02Pz6p9CxFZ06wCDeS4FNUSaQ/fWFQGBUwq3U/7XCKWs2ASUom/dgTPGxBI
CoToRWvnLJ9ceDmyDgKsKBiZlmLD6u+0r+qPlAV1uzsz7eVhxKQsBuF9XRM1u/ec
jFW827T0LCbkZwDqtWqWE8rYP1JAV3bciTq0H5Htlif4XCUlLR04ZGdn2epbFeaN
V+16QEN9bChW9wTaF28Ow387gL2oMKQ5fQECbY/dV9AAwNOdLMAsjV5nf5WB2WIO
8PovYzhtNhAJPzj/qffIXayEuDDiP0x++dEHOeKohT2IQwE0dAz4pNUI+hlPMa/3
lEEwKtbkb1tDfoeAdOM7T7ODKRn4G2yMpW6TNDdgYh5IAvmVTlQKoKVFhlaw/ema
tjXPVR9Sj7pMH8inuWGSiJfL5WZcHuUjQ0xgGpQpvkatGSAALUhEUQp++2Gh+Ub2
2lnPKAXXoT8bKZBXbep3wvDTg+apame1tjDpOHRzDNJKdRPxMWDaTVJeHFuwTiRj
5LF2uRtfjtfbwcfuLThcRKJxwRGidrIwKkr0bKosCWkN1HCpSBn3DZHg+8BmCGIA
9LSJXZEla2kxiOIAuBz6XXBIvp/zXJz/z9hORCX1R39XAZ5YkMSFmOe5yEDgCWXs
jtsDkkze+Uj2S8amxn+OTgfZTQAvVP5XoQYC48d52UpWqPHg0rN2s5q8FwOx066r
v821a+fuam+zjMzSvt+GY/RPj/i5fw6y7HFQlYSFEi2hgpxgW1fb8IdGuhT2leZu
kKerK+EBLvNBinkRVo7NfGB8pH1RMeSXwluEBYiiRKz1A0yQoPOPjX5Ss5tuIlaR
Yh7Ks7GIoRtN2bcoml6sov/Ffva4wkkWSRqPLU04UuqBSw/VD0tcEX0L7jbaIOcf
191dv09wO6Sc14nLaVLcrtJD1W7eNRzA80gq7oo3RvV+NoqlVU6KFMtGm2tvRXOL
nO9ruH+3Lpvps5UV4u4TM76VvyZOL+1TaGu3WLEpmS+Fk1ru8bcKcVl06qXZTALd
t6nsaajlmgbkAuM6u1Iq5EyMopVvTn3lhiha4gkGvLlZpzkKORZEx2rbfVQEcKtj
6k6KwFhlUQOqaoklcHi1qTOSvE1SfHLE+1Ozw87KQKLjJQlLMkXZ14Ap0M2SOqAQ
RwVEQI7BKrQRNBq9MuJXExxd2ViKwyoBlFoH5AbVe65fHxFZeaejGhu+X/rY+JuC
e+QtazHqb5kebuHXkrnpTJLuXTKUSsrdNp9sroDmRZlD5sYh1lzrKplUCi2QM8M2
8EzLgbO+46ejrwTwlvnSgSMYcGkf1gsNXLsbfC8doI2wfsOP/Is79zkdLACtxmsa
jKbIzuoL1u5mjKBY2CH9kqZblOoKqix/PhHwlpZlsxjZRfLiuu8r85TRLnbmmySf
umVKNilAiBgkOG+5GXjBgzfZ2bR092K9tUVKx9TnnE5AizLsYDhx8VwrrhTqMzgE
/0dajHXXTtYkvrkr9VuyLEnvFY6EmrtkgS4DjJ1uKxVrBGzfu+UP+zDjgyXd2K6x
GqftEqjSyVfcL6YE5lKVjTGcsg6gIsXwewgmlv/N16TmAytt9VojLtBVznkI0JHR
0mXe530mZyNWKiA2oqEuAwojCJxC++zAlmy2Ab4JkP8hVv51QmtZlAH5BDQJemys
JIPqaBHXLl3vE0QGh6TS/XQ97JUm7QnZZiHGBZRVpJKzs4PdXnig7+PLLIi03ooq
U3+B5OzvrcT9RVblrHKT8dENaMA26Va0gzx1pqTrDyfLQYWRxIgUPaMVL1b2rLdr
j0pAUGWpieqM/BBKqAua4pgzdiv0duKetgqRAzqAAIZ8zqqV9SF8wcXZpBoqzmEQ
2SKlx4jAWiei1CJ4s5TuouBwBOGEabTZ2/zL3pV8glWRISX2wd6+qnZIMPrAnMEY
wj6bjKAStK9wywwM1kzPHJ8Qjhtlptn/m6MCy8pLxNg2eK1/guziJ2GNf9FEGVWk
8qLV7DI9vGAkHnQzgxq3lJ2b837IzjUS8lDJZFVv/pqLjDsPTmB7Ip+mi4ugnreg
sMviTM2k233DGdS/t4onCjdnVmPw7MTTUDb+BdbkHZRWUKSd6Zxl6vz9Cb1+Vycq
UvPZtaVnasv6s/h/MBbTAWQEyZy8lvV/0U6SMtV0j3dfPc4uI4y2Z4dH/iUFm/If
zifVIjxe0uB/lwCZyzacugbwSudI8xMFUpetr4K67t5hXubj+lqQwSdpOfU910is
Gg7n46/lLcPLKnwYK15qqgFvkiWzAMZECAygY4IFzM8EaM6iXZU35uv500My34Te
IggIkD5vYAJ2h/aYfjAT6k6gG81ihkOrA9tL2VLBFlCiH0TvB6zFEAiE9QHYpVJy
7+mceVzbUBqn8Sh8jtcHBHvDzXHvcnxCIiK/c1zkazW0b3qglO1y7qLIz6FNm4Ad
a9JzDw8GxacW4sUa0Twx32onEpk3uq2+Ju912hQoYxJkvo8qdo1d2TPdW7lMazOR
Cm37OYpXbDEf1UFYsRPreaDOfyIquorRTM4dJdpl45dlxxvZgS+N+mu/A1fndwtl
XAtH4kKneWDtFfd027PtQbjAcMNn3WoLIuZZd2T1D/oSWRR58cKxmvIQtY4zGH2j
4g3v/Pl+nXnmrbJEym6vsglK2oks2TpJPmzILlS4tAa0RoJfXwPSOkoxArqkb4U2
KhNxIwPoWZBIOGlEdQHneSqSWwtP8LtclyhtHZyyuF/aOtaKGS9Lq4jcOuFnjGhF
93uCZwZpeXod46iFGLdjdItaLcmqhwabLIBKSSU3qnVNgMPBOczvSAukZAlPNtk+
oembHNeZMP6YZiSjUgdpWpgbj1OGBOqS/o4YJFZPXiR4oxcdRElZ/kn2xaHyyl+k
a3t9mtwhF/UeWlWQetW/cSHOcQR6tVnAVaVQYFYkoILnYfLJgs63V4J+JaI6ekjF
xhqB8cnaL/X77Zmueduo/7C0SdJgC/OazNS6PxXN1KZiUKiPA++EnIBLB25nmElS
qC32JrszNFGYtcBatojXQ73b3HKnD6AVEBejutLLMqzj9auiagLgeAjPry0CIs7L
1Q8QZggVnbtpjWwIKkfFO4GnVEqN7RQ+QKjWFlBVDbcCVY7ZDKnVjoNftjEfxD1t
v5KIoKdYNYnuJKyeQ2OGottnomRD+3WUjrx2WNiWdAPpjhyM0fMtcFtT6L9oTkY+
q51tAWAZ1TtEeYF5ktImN8j5Yo7DOW7QQEko0TI6gr/L8OsATUzYSV2C3P81zt2W
ZxG2fd/bJEpzVe6tyrkg5zXfVbzEfC5Tn+XFO1ZBntpYK9oHa97bbw/QqjHLAaic
KD0QecmWD0tfKWHjsqTvo2h3AT5qp7U5ChPCNz1Ftq//iuuyvP/LBw9OesCPu50d
IqblBKA2I5M84EAdj4KhZ+uHrvDQ1IFmblWHlA5kExmhxdmKooCa0wOkvBLJeOGJ
HUbPzKtcu2YOoKqij0qYCCV/GZ0sYxHRSjvp2vul6VUzo6g0A9XjNvJGjLju7qzn
TkUAg8rpOIJ+lphD1K+lUAWDiKu3LroRLL0YPdjRJCX3ZyvnkpIv1kITzFzvAfUG
FSqirHYuXmLadVyU5LTdOBQMnK9EAU9P+E69iP10NdQcx35JzcHZj3MeHfzNdXoa
h5hX4I9kZEuv9T8mBCJxjkcaszpYfbWSmMUHuRPbEbiGEoFuqzckiDB+Up+LIUvE
TK9uHl5xHNlaQ3CNQyhUTsvc/uhO4jNZ6o+QjKRBJvkbiwExlUmj4khq3NlqbyWM
+Fp8k/kpN+i4eUtIjv9kRY6CEkQY/lUorzXzRL81+Xi1aC1v3cVTENuVcsr0VpIx
uE+7VW7BudxGyWUIoaHUNDoU5KuAGjv9NbVq5x70NNVPjSrSBZsLpHqVih12DJP+
BGN8M1O7iuUocyWso9+Bf906ESJRRJwWkUfoaKjYwJHiTjLYXPsxpgPdaVLx5JZh
lGHdcHTYjp/GFSlE3iAtuw3nEKpfRGW58L4Rm9adq5raNIpCZBEdcozwUs7/E9/z
rAuLzxyFF/Frr0hAenHZLueBymLay1Q4myTJ4WwGwm3gtdMl2Z+2LRadEgBfB3mS
pLDlrcjQcaGvrXfdUSzqgEkdKXqb7+vmcx40EkapgYAczi2GEmrYZjYgmcjtW9kb
Lskx2D/vJrnC3RFaGfk5JF25BsouTaLqZRhqfiDcjnRex+AObbvHfWrsc3g5puEM
cpiOkFEcwigkfVldwWkAZhiQOZx8dII4Wz006t1/SKzyr0DiYW+fjcJ3vEQXmin6
cEtiHZCwVsZt9bJpMBlUHxIh82HrHg/3uLZ7ejRQ3RIUItzitAqDssFtYKMy7p8M
GPN8iZ/UgSe5bB5eScEVXRI9fJ/RiMre74Y2RyUC5sa0DFSpRy/fODyXudkvNsIp
g6jXvxfF/Qrsld9vZeOX8Zo1ewk3Ks2u4Wb3p35H0CepG2uPuS/FJCisfp36ewxG
zHBiyAIHYla2Vw/jSIvvYc48CHQpIPyyuzwlch9CWlKEV/6v11QHXupVnophMRTE
8ieDH5L/ZAmHhX8kfOo/Fsc08tEOh80qRr5kq+C/DcjaFBrIDN5hCK6zBrr1R/2Q
tttDKAQUA0pCPB5IQXzTHygdf2uBwa1uQkopQ3ossWRJo+3rtMF4TL5Cf2fwB0GG
7eswJNTNOZ1QrfDM4P7ArNDWc6Y9uaK2/9yCLeB7jOFwwFGdz2M+wuW4paKQDpNY
axc2TTdeUmb6Q3F+ZqYcUILahqKo5mLk6cTSt8Dvkt5mSYvrAn1gXBYH7MgMDdIE
fElPriEy5U16le+c04zNNAdUvzg7FONNckV6izHF9tekBFNIVVfidJxSzGcNu3qf
7E2zdmsjwnyRY1yeiawdQusNF4feHOSFglmfm16HldtzmUj3IQ9Vh/1A/f1P4XhT
VVEotwz0+RnY3/DLBL8LI7DVq5CDwMF44A/ikEZ+0ztvAqxzWKcbHM2CzF72IyUy
JOG/gLc/scucQacC3QFxCmtXUCENb7SKZzN687kNTMtCZ8xf78C19L0Y2plQ2hW8
8AW4lD6RIVaNlr9cFPwYj2fupPPeyfMtofcAWgGQJu09Pu5rPNRLS9Aw+utmH0Kg
kodsf1MLKTV3z27au2sv1jJwkAMPdflsxiDkeuab5vrClVT+f2cFb72az9SWHMyZ
1UqKcFYuSvhtgXTozY8HuUyvj2bptJ0PfypJoWm6kOqmHHohLXdjlxJHuyDf8ejU
ExGZIySVYTk34SrIy2kP9pCuYiVJi17cZCQ80I/iUtVauXFS3jqcQhzmzsDMqI6b
J/WfhZuOpT2fL4taqM19cCKSbkhEYYQBj1KXAJuh0KDIswLXWlRricPPpnHJXQEQ
/YrmRTYrcwDqjfBpQQYx6mfCzy/bKfw3ajFDjSxjfPj5Lpm21TdkuYqnS1hUQexz
qtbX2vBF9/GYYj114Rz6lg6N0TdDZZAU1wp7A0NtNst24n3Tf9ASqGVDFNHLGjTf
1c/6UKakqpaiPbR7qarPjmK6GR+H6G5NUFMUFoM27cvTiDU8n3+Tigeny2tuUkeR
8e7L7MD3axag4rI1U92xpsXlztr0tZfxXg0I7gHf6o13zlOt4kLIffp2ADi4aBSg
9/ayzjekHqC9Y0pB0kbBoTRqjZzUzkj5naZLVFIjiH2NJ4wNiP278rv0wzbdKZc7
wBE0xUfCraZIYUnKR0+iB+aj7wCDyma9EFcLFN7D2e3WSdlGaQzxhA8XyWM9XWaa
XOflwhjDxpxWYv+xPIZy1KrzsduisuqVYKfL5qpTrTti2D3qwrukAwWH7npjCP3a
ZfY1pHflGE/L/zMjV85xj95pfCufSDNsp2ZelqzE3zS+tAEv0Sjiibd3ULDq26yE
Z0J/R9bryP4WcGBNMO70Cc5kIzeXRhXXlUL3tqF82OUjr1mQDSOXW7PJPp+mEmjM
GByvgv+l66/FcnFMpepJplyXT1HN4AXbNOXxXvg5XDre26JVzKg+QfK8XzaCntHY
vnQuPsgr/BITRceJKoJrCErgSIgbx/LygZCC8rOiqTTX7vuto/nWZupAIq1EMdUE
zw2E3Hi8/AD2jMYsfCOrJvpYLAN9lo+w8cVwNZaeUxAwT3bWHxZJEx/qNNZc8VRJ
qwMRpL8swNz6hnZDQbeYNx3vk2hQCbcO9V49O4Dac0Nev1OSN/buBlqSLmtWR7JB
oXaXFHnLHL2b20ctxEhRDVXwCZozHe6h7kBdbqgIkb8ZHKxSnfcWNxtpCYcCZZZ4
yEidGiu3DrIw2vIl+oVXdO9GViUHSOxemW0iIoS6GwAGvlpgIoVyylUC4bsDcvr1
UIrDKeTQhbR1zWUskuhlaUWBOveE9fTYkNyuG9WwkpZ0sI11HP0Z1CvUcCBioCvm
8Gm3Qu4iSoT0+FZ49yKog0OyPnLdroYWaD06o8bRqw2t+ZvewOeCAe+UyjDYBtqf
eoZR7RxfrGocfXMc6lPEm0M+ZijKDDIiWewu3QfimqVq4bMgpLbXsjISU8KXaZ/h
BRpDI/Jr77SPSQfeTJFmhByD+ugelYHS5m9Iu/nYMuz3ipFZ0nxIkkHhSbrIZz0F
blRjp1XgERa4F8wV9ewEJ7L/1A0zutyY7eWKXnzgHdnW9g5eE956IDo6Nstl6d60
3SjomELi/xtiAdTgAjkseEsyoY8iNvLJcGBOE7rHPnrug9LuzJu3HPfjx82g0H1U
mynoxdm37Sp34GeQ3iNeix9hNtfRYC9FsMdK1sTCqhcPgmVmyWoQQvD032RKMIvz
csYvDbR2MnG/YJAZ80LcRyV7HaKx+4apaGCqMoz1jzk4Vnbuw7DTniBedliJfyhn
8NSpxsijzR/MRv2YMQlQ0mSf58iFlW9pnBJVOHN14JPmBkpLd0HxkmzX1loVildA
F7ebP3hHPoC1ovU1JKd0qNxn6WWEA8pBpWi6SD0jL/vFh2cVrUIZpSJYjDyR04rp
ag+MsPZxPW+rbftFkNKkZ9j+NiE+doTOt+y/0V8CSirlgCn0qMqK9dKYJ0Rr6etj
3//Kyf7DySordXSh2A0XuB1pS8U+AsqYLoMRJOmduTwiQmKn5pyL477e15FEB6jC
J/NG2cOfbYu2fFTUYqkYdWIezz694mwc2rrGlLmzN5Fz5ruwpDmgnpNhRwg+XxPb
Kzcf8GXty9P5S0F3q61zgpAQXDPs7GWa/eT0pE1ldPxY4vChaGm3C4XcBQNrsM81
jEoKk78Ov/3Y/3VeUbZiVjFlsXsim2a6old701VBuSB+rqF2d8pDrf3p7IUm+oE9
Q7JQcyxb+YGCyEgPpBpWxoAJ8dz7F8iJ7IVGpdEg5Od33VpXKRYL44fPY9Ep16T5
nHveyqfKw9LixenivfN5DllK1HHjs4UOg2QtUIwq358XZedD5d5yNispc1e4JvGu
MDQ9WzGiMajAXn65lEjv7gh6DLOSrQ8gupT2VxYjSYWTcTM79+OFqQtcP5qRgKzW
+mJtXT5m6CEgu3WVVmkKbsfqNc43aM10cDSToGplmYDFwPbA3VUjyokaWPfHK8tU
b0jEYqbjw8l7dqnqdARr+JBWOlrJ3+bM23cjF7LD9ECQmXbD2jUEWP5WD2Q2ghsl
pm8R7r7N9dDl5k6ApOTdr7wwIKVKYVIKEFnjBEkTcr16Uc0SXrCVtMn0fDc+EhQX
1cMzliLqN19HBPBmiRocEJmnf6ovxcGYRxLrakouA7jiaXMOkyRnNf2sxMhLdY5h
5cROWEhU9an4C85OU70PjLViGhIT2/faJ+nh6PzfyIMBX95bmXoV7cyloIA+iLtC
R1H8TGHytEaRRauZyLy6LQaBVPoN9I05fOUJ2Ez+fI+EW8Ljzi65D4/rHXHLnfGs
okdVWj5L81xzfGKV65hKea5j+9cIw2Iv3gU5nonmjzLEIor/ew/weKBrCC8cMk2h
6yO9JSdgLnYrCfSFvMcBWUumUxEfUPOuN3fmVhVgZsScgty0DtLb/M+s7g99H9e/
qcwg8LPu1py+zt3sQ33/ZpoplGSMJsmS+8m8LxHqpRO1n42X49Fq3TZEipuyJ8aj
f/3F9jXBz9H37J378O8JUKym/veTjTZ0fkZTHCcdFOQuZiCuUULe7l2AfQvP5X5k
bD8StSzzPDcIGNv0+3rAsi5eC5+2EKrKzZq0q4pVm+keFoewERDJhMNSAAlwwNh5
G6FXhmtO1AIXCc3AwYL+r/MiSYHRwARYFRba2NYD4iFDte08mpbk+qQyHUw/VVFe
dp9OHwNGz/IVKMYjKIHJvyRVF3Ud89bW+g5D3B2qLBVUKDrqPNpb63b9coJ1PfXn
KJNmT/w0vJFGHvZ29oDKUNxuLgyqNCjaxAqAt9d/pYcHa7G93Dl3LXUQg1x+yJuX
jpApaIKJYt+Ol/guPyv12MEkJFJwmSI82JSMTiOnoyPkXnGEJYilP3weZCkEn+p+
/IvUzk/k4sArMV0xwXDQaRoOzpyQ0qDwmFz5vB++TPqYoHYIIB0V+aG8zwhJBlmH
ABYgz5qU2U3f3s8lYdVJq7bW2pB2YNI2Vh5ju30n7MZtuocVHtckgS0II78nWy/5
cWPMRVB8y2UjYCyOard2zEY08uJWrR5yxT0fC1doKL3ZG0GB06/d/raycOpgOy6A
AX5kV4H63tKw9wB1OvaG/WKjbTcf/JJxg0FeTy/JvNcPYCpkC0warEoXuhAAPVXZ
1d9uFy+2jHvxN7dmZT9s5Pe4hnMGVO8SZGR7O+pDbuCM4la8JT0Rej7GnT6jejhK
7Sb4/RiFTAGPTL9m6IZiJXSNXG9f2OTwzLGQ/OAnF5sAzBRSt8g0HZ+RWtMbmFx4
1EjeojZpOCW2F4rOV4x0T8NgTB/cWWgGZAmIPk0ygUiey5m8inMTL4pentNvby+k
KzjN3E5o51St2qVc75k62+hHaosuazOZvMTss0csVgz8zLKlK5WxwWBto3DNfToC
9nxOWQEe0kNDtE2LadlEX1OGlpnxIe0njVr4CuzafmC7lRHdzFoCc8WiTPXoVmhy
BOKL7yFNn2MBRorc8o3DWXPDKDqOe+cJg9io/jf6rG1jM0DI3+5Xh+1yOID9fanv
rkyhjt5DgQ30fzJ8+Vth6aWKzXlKgTkDlu+bTWs9wvVSUQzPb5FLfBcN5J6z8Jme
yZhSHgMkSWJhIRDddi5MkHCIgPVtqaIQy2CJWRaTA7vJIkLDrKk+urafW+njfiLP
ezG/2SBv4qAnKjibfXCNFoqaZcwkvTbf3qkt8veon05mjhMSKpuw/crmYm0GR7Ir
tzmiZHuEBxt+scLr28yeuvEZ2lU14hlW00sgU4dVF6QehhMnllyobYAICNx45Px5
GZWoyfAdXPIjv4NT/hMV8ctt/QQRvippYyh5MyW8DL5pXGjMirDfrLU0E9v9r+me
EcpZKXaUs+J6sSmnktNRAUyqyozUw2ZDoRW7uFStu7RB52y0HoOCcwhs1EQ7hhrb
SPGCz9AR5HJLYqGfHhb0mg3cJQUdJtwU0JmRWKPx2rMvu2vhs7x6luND9UHeNe0t
Pm8Ebmm5gF/XcZfbzRjIJJGyEEWKWEqq24oSRqquMaNSdH9EyM4LQYO9hvS9IGi8
uAREbPoxg92WtnNJfK0LLX8TrYl7PLFDN2jdMjb82nJgE2BR3d6iJrwgwVsNKQlO
Spb06g4vXEvsEXY92Q2YwBRt2lYU5OwJyyz3vdFGa0hvTzuKbvOzRzKg22b0aHjg
JVlc7LxcfrVy1YDfj77NSCVfo/jsAhiJX55PodwOhZ/9w56Lsntmn6XSRaKCmzkS
/oG/gyl3VedSA/i6MIc/suwn/C7Roh6En1KENYBpW5gMBzpLI+fFTB28qOE9RGBd
S77OegMTeQ5PZlIfA222urozbLnOdAHvFO+TRQpr2LsFyAFFPry75Dt5jdfosHZG
bAephroXRT3CDhIW9khkxEeHnAMxLcOXFy3Ys3ur25ea2XO8e4w0AsvXUXdK3uep
NdOWqI6TWXm+Yj9Zm1oHggs18KxMoihCOHTf7cJO3UedC7+JCyPkuEMkIpxcbMlH
2oaALX49ulROz+kmZj1gfK27xqtwlFpd8PPwoMK2owB1y5AJv/OWs4OoB7jZjHeQ
Mv6ToTMYUSAO3u2aTbZyHfHaIlC0Sb1cp7A7yJp5fzRl6i+X6zmlWizhFOu+mdBg
Rj3e3o/Ln6z7TZr9FtTvopi0bKa5wAF7c8Wp/4SkLO1IUFH3/Fgb+QZPk3E8pfyc
uiu4Lhpis5A+M6XLOjoy4gRqj++47QesLDig6k+OvMjVIzZ61nayLdEOrpSvY652
ZkKET8jC6P55RCCb08s3hADW70sZMORyUTSOHMOPzfPm5v58BrQURL4YhA/9twer
FEt0BMjNqv2HheDQBQLTE3nlbxlqcIrfew96awB4XRvP9dMmCvJXDr+GDh0XwapT
jZMqtUWM0O0ZH6yjW1GrrIS4hRadeZCgnwwlehb3Vr9RyY3vR5uYEIgVRFbWv2Sq
MLx4Ib2vVeqOmXcqLKjMLmMe3ZLd51KGEu8r3i0x+RPl1SStXQj7qXgrvTVhRBbl
sseAhL+d9jz0RECx1QeTX5cm9/HgoZlIJ27NIjnLNdXm5PMdSFp9uBQrgBWfKN3n
+KoO9kE/5jdVoR0RYayK6o7RHPYiVHy7MzDeg964Jrl46v2CnQlUnjX4FKtKhb7H
za4Ly9ZjWwHNgYF5cAonCLIROlwySXg69ERdFVW3xcZbBU19S7nSx2yjXpd0eRbj
7RsaaG6ntuozO6/YRZWe5yok+oGh60thXwlU0Hgcy+xCgxyrMgNdvdjYlMuej7I2
Zg4PG97O6C+eiVv6dlKsFl9Rl9mG36FB3oY7cawuy1s/qrwJkdDfZIyzUtpaYF8P
KfFVlu4xe9hLmsQsYwF2PNDbBuv3HxZ3gRUXMYDiKxCNoeQvUnQadd+ytOPidRsb
6cw7lfZtQ6N389VbHf301S6pcOvFoiH6F8nuvQXxQ3lEOio/g+aDbffkGcvBumMt
xXuiCzCrY8Awtsb52i8CYdMEDFYE3Go+erB+wTqbrwUOg0Dkwfa6K1lV/fj8CfSm
YG35D2K0qx/60q+4l2jOly9dawJeia+vZBC7XREhPjrGNGX5T8WrHjaNO7K2FY24
2EFOtKwp+KmJzHYzoDzo7W6nVr+8T4GjamJj6SlHiTyXDSzq9aGRQV2xV9dUEyf7
ROKnsm3gYFwS0pSHQUPbO3mVRvoYT+2BFoJak60aHEoVp3VDoaUGTrdzPpZcrYOt
llvKHa0G1t63qQfvhqNR10NzSTwfNcg7KoEui2lbMVmzAd0pwQ9ysIId+9m+jb99
NT3q/OQTnP17Xbbztdbwr0brAqwddxQb8iLKq1wWwhzFHXCdP+pI+Yk8lqNPhq7L
To/VT1l0b8DLyrM2vQNvrQq/Dgy6GzHBb8fN2SvPHpw7W47ewUNzSViqJExwzZ1s
EioJHHlVL2A2tX5bQ5Xi3aPm4WVveYGKzTH4qYa6P9uvLo4uvR2SYQKo0u/jo9J6
+lCwLftIMcKsazB+vQx5OfyASVj/9OQVP3UZdhzEHvpT55xfFkpxyZaJRFoHC2M/
sQptPZLrCZ5WD6Bur+tClYEPksWadorw/lRjlmb5YPDunDGB1XdlVnfjxmKDJTaw
Nic/X9Z1z6z+IjfFBFqeYoOWkaP+potY82ShHa91e5dcgB61nRdL+8f1NLiDQ1gu
TlL1bk12PSn5g/Sj68fCzMjoqFUWZCcyHBvfhLhOLYVsnY1CgdJbbHWaYuqQaL0K
Kej+nrl8yjv25mHhjoPGmPYw6nYdtIHDfjKMUlzY6t5/kiZcOG7x3aChoVfon1wK
QYv6LljvVi0/Vp3S/hP11TPQyzite/K6vWv5a9q4Qg2b30GzQ9Hq6bHqsScOLIk2
hoeQwO0daWUL19VSE1GyXl2cTMoNy98bSyDqmJQ/xHTuFdvyBnLDuVjWcXHkhhCe
YFnarCVAHK6tdCo1XeAdRHIkSsGCt4hXMFBwRE3KfolxBB+QCuhAQEm9LRHKl0im
Oi1ej7b7xRee0bL09rhRI/Y9vodEZfFdLQd7Jb6zCQfmGvjPWr7s1ekFj/YPDXvG
WJEH7JDjhqPd0H27dyRxaCOuy2sXwWyulCdRSFAJztCz+TtZadF/sBic3bNE1v91
YGRS49a3bO0iNCjN2Qsx2X6/vcSYtvuwDrt/Ukjq9K4izvC6mHCFS742VanGAw1F
WXROFqxNi+AT7vV7rKvsAEukVtVDUMK8+lWwjtjtxcGCwM7j/hi9h9ETviqGBXrM
DeQeiroDD5PxsLaEQu16x/pKEWZvNwIqd5tDs4GYbCPpkw9O39X3IRpUQf9DG50Z
FqlkPX0QduzYeFml+Irnd+tdbllltByxitSCllrKI7hSEH1gV8gpYFniuXT3/H3N
rve9XHBpCMx72IBladji4wgk1PhrKc8rNl9WJDJnnPK68SbbS0OhBLsUQ6rS0/M0
O2DuafTJS45YxJ+hLx0n/RMza2itAX0MiiFGwL87pkNIeSbsbNWKAMlxU9yE+lLx
hzGn/wTJuv38Z9XGUZ1+Bv/3eC8NhNQGYzJxQJ4h6ejPFKGv5Fp5tZQKMePEkBj5
1Comf5JvYdIY99M0rw8Wqw9yd4Al2hewBh7WmsyZuZCfetspK8IHA8X6m9KUiC0L
h58PN+TRpxXooJlzHZArEZwrhJgXOFm8rbYpFAolUWKes/MDg+EQsMuPi+5k68F0
Wom7tLP8+VZQPP0POLIoBrmPEW7AmkcpPs/S4jn7YR7vI0bT5E98CTAVgQUProZ0
v3NdFJoU5fuxykB6TKCFlh7mUCMyB2ogXRYuZkyAmoMJtBH1qege7JLa7L+9OPmJ
UcerMCzpP8fJtgIDX+qN3jY4ws7Cjnuw+SYRZhrCdW4orDKnJphSFENyuOsWAxTD
ItzpoehOSoK8ViERe2bHoSIJwbXeErL3tAhy85mmNSlbNYxAHAyD/D3pLX6oAcbW
tTTnTQNjTvwSGBN9EWrM2MyaiHToFy7ge9OJ2sQOIk3Mq+dRa1pbj3s71pB9rzXR
ln/clNqKeGcAMMe8gr6cFVjbdfMvAoAK1KxRDvDR+9K/57q/AsM2yQXkK5ewrQ8P
Y14R+h4Q8l8am5BJA36CMuyqRhxaTFKawXd/76wJrBDibcL2IeYDLOZAEia92MTA
5uPyjnssy9H09OVY0bkBi8NqawtrVo4nn2lPUjztGbjgAgiaUfukZf1MHZaBlZ+N
gL1wCEUntl6tALfj/Rb6zCw4Gz9ecdjfSwhzc8rLz3DTpFA0aZWB7gU8RGU9j0Jn
HVvn9Rr97/DB/IIp1gZEgs8cTs7/Z9Qey0GfL09uASCNN3H7avZOn/LBa/PCcN8/
FyOZFSHnwimWYRckV9YyxeHRoloPPJgLgLjCsJSd37zeRHXWCEpES7rjo3KxDN3f
NdJS1ZrYy0QCdVxE/r3ZKB1VZbIFnscVjZ33bno3D8RbeRK5fFAxg/0pD8tNi40j
3DzC8HYKv0TcuHcel/FenjMmnMw1KhhKKTbPIERn5eMZpD+hsuhqIK6JyPwInAwi
9IY0+qvdcvOSz6/hpxtQr752W2W2L+zllGyGkzHEb0kkCN2k6j1QUUgru/LIp6jx
Gglc0BAqbW/TNUODtmzQf/5ihGsSY2RxKmTlCczMjG1H0EHT83ixqifTUNO7mglC
V8qS6J8xfd6I6MDe2RnvPrnT+a/b7qCD81wVWealyPyrgF4brp3rKBOYbsFy2ugB
VOmMw+LnvDEIonqV8fRAg+3VTrpmDEN00hEf5f1N9VkOPhp2nH+Ll0LHxIaAeE6j
DnOl0dvXNRh5cmZTr3AtI/uqvXOthCfwt8WZSVU8FhWFcrW69oo4lvEhDTWmotWW
QwpoLhrqWEzsrLrIlsLuHxHuF+tJ5HkUMlQZZHl68GzmZ4AWlwbVkKROk//M6YRS
pYdNBZtGwu4/Ywudyc98Be8WJ6svM8VNjDyuhVy+fY5gE3PFiTjDVxppuFdIyFiz
+lExVtpSBH2mm3ZF0B1ztBNJUqFu4/ZwSl/RMHC48kDEq/fhdXiqHWckKQHkEQgv
4vjvCKqnCPr2Kvq4KFG/RHPOUB9BLsdLExxvhFMUTc9vprdmc1/YgN3Jpll3mCNu
tNyrlehMqbDVdTFqmiiZScqPyUePWgiDu6FcLl8kr4STEF7pXfMmIjNwqkYWRrrl
PlHVaNOMMITS4vaHl3QW1fb9vFihhToR9i4iMGonk+ER1WsecJ5J4WlKSTZ9CIWC
Rzh98IqzPKhychtmEt07M3yzPjP8ubKi2gvaR/1JMVR2Ysy/FGYv5KgkDGNR1+29
XWTPoU7WmOofdzlJwfXQKj+yH9DYm7qNatLEgO/MWyjKXlqQQbXhMU8F8L70/UII
aYxLaNlxQ6A7/D95/uJnQvOj4oDHth01BNcyeqcv65sIZEPZuwIzhfradcYEf75g
/+eNfZuOs/OvWxHj/RQuv8gj/lmw+K2w4d2ZCjWsd+1QOWA6DXR7e7wyf/M5m/QK
mSm0T5n7vHVZu76BqX25NkKLnnd4x3AJLluLm+I1WkxlDlkMY5htG7PKufG/c1Mm
sEVh+gPShS05q/MVQwK2ge+mu+qT/dkMHCK04gzPNCtTjXCFXm0P58YFKn3Hl9YP
1RD/1XC/ANGwawm8ulSKIphnhCdJ2VUTgM0mw3OfSxr9fSix+M5P053kDDZYIeCS
8tpZytukBFj2lPm1gQwRia0jSmESEvI3WVIJjNTp0EgEoqXrWsfNqzyTQxVVbfs+
Kgv6xn/L1+zKtI+ytI+kcyLk8mzHF7Ix59ksx0+utuI7GpqNAQS/Jk5N9PdTXbVF
RFVE5nhfCXkAsrmdaljLaag8fVSLEtAgWkGLSToOOWODztCW+PzSYpFkv/tFFCcX
/h4EUNaHj9EvtLiTQfta39hitWxG4Y8Hm+8JG3jrSbOjOfzOWnNEL+iBL3xwC0o+
wsBVcWTiaxkd3K5AIvphOiRCPbfOm4x1OPYhLm6i6cFzXB0Ffs0amJ4PbNpS3D6y
PX519nONMmCe+Ko0otbAkXqj3TuyRreza3PyqW70XkjyDdDEZVrKHrilKLriTyUk
Qrw2y9uwscsR71hQtSjdXh9AEFnSDkpmxvtswonv1NnEiK+LCLnlXJJGWU+OasEB
V2Dn4zmbyOkuOZSA33yHX+rGiEFX04fUPsYBg77AfPv942YspRi/YNoadrKuOxbC
F3bntcB5MjYA7YtKv1Je6zRCr/YoTMMKuZCuKhN9MRzHIxhDAPyiHW9RbL6k15fu
CKZEPiE21mC/WufJt7OadOf9XqFWFR82oLWGQhEAjf9E+sp0zlpZCjqjOWQlWVMI
owHGf2urSSuGvPCNlrhuSnyhbplhVPXzsBfKDxi+/u/9zW0NQ4fIY6Z/aCiikUAI
ls50D3WQWUNs7F1fj0zQkX60ewAn4VwgTuhCy0sU8kkS5t+1InJq6e/Er2Cnjowh
jQxCvlmU+T46NyqbL/URUb7555qS2Ntho7XVbu2k/o0XuRIJlM0bhgoYxis97Vo9
05/KrA6fVmPorzxfelK64eMMuxmxqa71KcKdpkCeQ7G/2EFJnLCha1Cf4+jakH0g
/shqwTU9vvNf2lUGXhlF0REJEH8DLw1f2oDOsx+RCV8gpXmRfhkrhuFgqNbLdC1R
uyg2Rg6z5mvNyZ0uA+XEfxa6ImbnzUVSuB/c9M9OhiUkaKjweQcYGSUV86G6zdMK
A4suCrxfdcdVISzf0LbZO0rRPdByHsRbVXx/nzx6lmPuKJo5wbAhd9QEEzEcO0D5
1WW/iMe+dp9m+U1zaoL+HnOnm2heQ/sStpEh/zDfzn2CkvqDB+ckq3JuTsCNRgJV
gV95E1LauJ8YJsWR/f2QIDH6Vesn3mMy5B23lZDk2q9CDjshdr7EzGZKsaFS3x37
eimE0873TUd0vIloWMEGzGidsXlw14267S34D/yGYnNpbx0A8qoGd1OesmXCf1f4
qY2IWDck4RtVEJablZX6ayS/7xmMypOIoU5PoluCBPW8NdqvdT/oDAOTFEs4Z7gq
EHPHAgNikxnMTlhSU2V12eAc2hZSZOzmsiiRjWhndoCM6hGtvOp9DMzfyBkfQUBM
IvH+b4kVI5iqvmXkMRtowqTCYlm0QpVL9bl8bqU62WInIEjRIlWE3PHzCinuoCLY
mjz+EUOMR2D6u+ZHqqC39yW2aqOUubuP1SqeBKEz0832xr2pafixkB/LYuvEboxd
wvi8vQ4TAmNX0DofaB4WB/D++TaMQYPvbPv/j59d3ItgI66g0zLD+n6wmpHWKk97
J6G2Cp32RuAT+4fY+mSYJg07BD3smPln9wyq2o3Z8BnvJ1UPbBnqL16pmArWzzow
9NpHcoNMzuGeByBJ6YiFgsGKoEbiA+EH0Wl/bO6lPs1cOA1GT7T4Qgm5eqxZFbv2
cbXW3oHxF5Ky1RN0/ieEuuN+GomZXu+i8NuNRXS3IfgVQIHLzwo5KDKfUdEJ8bID
0syjhWMc6QkCdOTUlGfULsasLrrurMyuV/db4ZClZVMEc5DbBTs+IQwqaQSQXjWB
iV9DmHoSMBJBsZu9ccO7bNm0+DcbFWecX1GZjWHkoCL3Flf3oUK/WgyyWbO5umxC
py6dmRA+6A3Xoao1PoELzfNjrwHU8kJOYnXbWd9UYRM/K14ldCY3FSEsnmk9QTG6
9LEp0FBEi3eMx2JM6WGIfRCObOy9nvHfln0drrijTCZAUBjbtQJNaq1ZAozLgWKg
dHi2j10gX0JfGbnpMEHv30wpzLUQQcU+ut0SaxMbuCfo6ZRexHIys0mcLE+TOyK/
C3PSfhwPDkFGOvEoAamU2GwcMXQ5sTrlh9+fyoPmq8M4gzKgAjKYlWq/rrhxBn79
3bc2chycW0ggdmHm0IWDvku1eb6EfVtwssV4i+ONCpM5hbBVzde3BRbpGAz5jxVg
TutfSdgaCv0mKj/681bT9MkiMhBQVa9SWk29YXvQrmPKuWczpWxYsDa4pCqzgthu
EFCyb9K4UqWx5qwfQXpB3Io8Zd1aHBqrCEdpotbMe/NIok0yeDx2YwFY6DkFEeLO
jpJ9nnGhgRXAfO+j6WqGuKLdOIBzj2HEduEZ6JE6SZKr4EUfHQtfYmTC9n4LjWLH
0fvw2YuXPcB5eazoWn+/MEjy7pV+EIlpMGZ+dtyI2b/+teofrZ6hq/KpGoPK2pCZ
Y/YDHeSPBr3Gg/YTwvSw5wS+yS9GJbLMrCNcnyV4dSMXjunlx13cbnoJbvCVNVQr
OcIpByxH20SbE6Xv4OVrMadSGUdmlm61HROzd9eTahAt02RHcCCdV2iH12ciAxhi
pVi2Y4NHF5n/bczYML6BWOWOQkrRBYoZhWWxSHm/lZbbZnuIhIJsX0C7YNn9VR/U
BATJRiOy6gmHElYiVXTFnyekrmJ4oYp9qStTKYl5WGXdr6bBs4va6kc+ziWELZ+7
Wnf6kEF8ccK1mvdMAFmUESBhgeowRbmKqTwuddBAqAxb+G/FPEqfew951mtIu2NS
nWObnGBDRM305v8JFdQQrItrQ3MLMbuKqAWEe41OQ3vrjBBCFQSa7ltfCFUdbCdz
y42EqDXaQ68Cgv55ic6MvhRoejPRP67fWVBuKrzHMqFuUcsvf0CrRBwljYOP5W3z
VRfWPpzZ0VPPsuxGjZLS8hDjugsnQ/HDWktPewC73Z/mmIx/DWS/PYG8Ne5Dg47v
Eelbz+lMLz5bLXEnggzx1l0oY0mvpSeXApjfX9SopcGHTGqv5KtBUowCdh04fz9P
AalZJnY3MTtudx0DARqAjKLZa9MR9WtQVL2SevmkZR6g2Yccthvrdn2sLZ6O2NJw
awGPH3mABWsr2zftffiEdjtu8Udsk0VzsMCE6D9P3hhOJn8CiC97J7h13CkSJE3J
h1VBxvbttRgKy3KbXLcRz80JPuXbRjBePO6ubZkvUy+iI3SMruw/+jQ7QafCXS8i
D+JDQquXlWsrqUZwL1mxhAFFz09/s95O9Pa3mNULTkSGXpGtVucDo7giC+saefI0
gFDPrWPYbaNVzT0hgYW4qtbEd/A8ZGJSH9YhmpXzyXNh77SljuN033zNZ4NNvID2
6rtEGsA+2x/4nvktjTYL/B22xVsJxXZUADQVG8pE9oqneRyxEOpJR5OLKeqYHtSS
Jpdtneq4j75EGxm0oJdGLOcsRBn4FkJQb94itdWQtDGCkEwJgFOl29v713OdGzfO
dii3uwvdQmPW4Kx/2LAbAUczO/415F1nnGuxjTxjqWlRkUy0wNz7iyiDd+6X6pdO
3WgLR9JC3ODLCot5edWweweqHvBDd1pd5Gy2CHnNaUg2Fup+dxkNK0raS4negZny
P2LlNXzDQi2r0mSAWnFC0nldgLknNJ2SjR2r6XIQeE1HO1/n32MmFWYLt6nmN3jg
ttVzcR4QaVZPreyP6pXmTdXZg8ned8O+P00Hc44aPGYEBeI1Us5tbxdN70EJXoY6
SMg+OZbwMGLdEVr41NM4QNwlMZzOXPBWGP9V4Jr8qXazAA+JXHbNDLhCnPicPqqi
sz2Z39typaWGwb2U+J2BhUJQmz/l7E0jFP0kD2P3uuOXb9xY+g0Ghl6fZMYrYVP4
FDTwdwtoEyf1Bq/xBm55M4WrXY4E9Eb/tG63RcU1ERtNCswvksVyHPoLB7XPTaYK
gQIarTLIQ5Q9xTp7lcCpQhbmM9TKCBsiB3VTduHFREk+YCHQdC54BPKPJ3aqd+ya
pmm1S/GGwuAL57yUwpqIqzleTkPORP2c2TwrSWlJ7l5e6Xg8B7220S+zsXWR8WQ+
ek86UkykdQWTCnoAo5+N5n466yd27npwsiBRFagFTXIBvkeoZYPNv2tCmtkVcIX0
2A3HHJ4BaaHYBUUcAYX4StRAtwb3gjtTuVvMPldY0bnB3LUXzLfg9qEGySHRsquw
Z2mv6fR5bO+QL33XP5/YlKvuSI9kXp/A7735fg5gwnAwuzSlcE9K0iM9YSG+592M
h1buPqU/YMyDxwgfMWgFRhARodNeHecxDSjX3oQ/QutiaHDByVVNxWWdbLOJggwF
Fvp7H9138Joj3ihabgoIenuccXiZEM9gfm4PJvTYSRSLidJvtf5pIy/uh/k7WVid
NTETVXV0uy1d9wKraEDLuxOt0560k1v/73oROlzPZ17nFFXNVtwzCWNEF6U9HOJC
JOBCdmF2qIzmgV/IdfqQGmS/yRYp9mXeiCWeSHqH7GE5Gxvu8lDayyiQvBXiLGHQ
8xKywRZJCHZdw0jPzynyVggJWMgSQ3siL4u/mrR+6TD95IbGWy/3laButVYaNB+1
kbqi78KnOr6OZzgD2vCW7+UJlxG1IeN4U1N6eS35JxTfbrj3YJcAeMXmpZSQxnND
5hcFC7sXKKk4pcKI4dD9m0sTTgTlAlWZsctTSBlIY/H0Pa80sz0mKiJjL02Yubam
sNPD7ix7+Pll8h5sCYq6Kvsysvjpx+YL80GnrQtBm1y+waIPWyDTMl2Ma5w/8L5M
tVbJfnpa2MbBRzAbXD0GN3YNcgq6GLH/czqWy7HztlP27c7kmrPF65BseRz1krGO
wjhmbZBUQOmTaG5JwwsX86e7R3TYJpgRW/IWbpIt04Ygr2KeTeZ3YnHhvutJBsfq
g/WYpN8LWeBsPLkrvQL07RdAwKUfi234YnVgMpbL81Ex7zZD0DBYpOF0daPa8WoO
RwPuXLkoBJmlAUvgXMXxONw5Ebn0iokSaiiTRGxtDxGwnB0qD3xyYPZwggORIqRF
U1PW98C7j6ATkkhj3MmHVvJTQIgvFLg2YK4yowdQZVt1UoJnvZzzDDHYtLW3VMkZ
r51kKwC5dox6Xnp2vbtCw6rYYjysQTt2iUB+36EiLmNugO+KtBckYQl+BEHs1b4H
V7Bc761eq6asIzUzLk2MhDAKe32Y6FWCZihRufrccteSD0SCPqAxaBu640cHmzTR
7Kv8ypzpdljBvA2uLKkYc6Qc4mWs+7LeN9qz9SdqmjfjjPpaOB2yRF9cPXZH12nS
7b3KefC0m+2Awq0ErXTvegj0yJCA/+jD39fZdT1AtJ5FEp6k9Mnvewo2otvU1znL
TUThn6HvBWPQWQGCxyZlHI1VvsGWAzSnbV9JDMLE7kz+EvMsAtTy4qyrWlDD8lpT
5HnqKAyZr7bRG+lJ9J4/W2k0ImaWTIKSRM15Arc+8I+AXQKv8gyYZrd60r1BbFe+
0xZkXjTRHcJwjyI/tOSW6J43uR62oOWSM+lojCO8A10bkKAgVpTqNRvfYfv8THjc
Ep/Oh6l332glodCyjnMMFO94HgsQn2R3tRjsMMP+kCkaphV3rmqlddwNLa9jFY7U
xAFaKJ3ntQGerZFGg5ZhR7hFlY2rk8PRchtq//CYiPbzxwhvSCo2FH89sw0f3c0D
1OqHhulRCWIwRLU6/P71kNOEdPZGcF5H0k+HmTqnEDznbz7wBcUHBonqDG9c4+21
enW4Qc1dhK8aYAWqg8C6j9zbcLe9fvf195xUsyzvna9b27wRRTekBb2jJ/24usL0
EPsWuqRLCLonPXDwfDrAZNWIE/z/XNh4xq2S3E1jh63CRvEiirS9NL5tSZCECLen
rLCKsctpcnK6Zmrs6J7VvP7e2nu+irjMwGGYLTQgm/klGCJIZDCH7MvKB/Pys5g6
1f1HzKJvLFohFoK651nXZvivWLsk2lRifH2ulZUw7dStkOcubqWjcGZ/2Ygzti6c
f3lSKOI5im4YNw9U6iahyzqNsGTWz1YxPZgiyr/GByVl65+42Wjgo7eiJSZDLpD6
jak4gmbV+EiTS6q9hHBtgYsrcBBD3DYrDP+pSJw/y2i4MPwQWQ5liRKMPejQjsU1
hH+NsvfMvXm9STKEi/YUy6vwmEqR5f1Lg6mSTp1+8bHFKWY8T7VUUMnhO56ZdVv1
MZGCNiEmmVFAFBpFbB5AomnqwH9NvMd8q08K+y0oCMG/HsVNMXUSeDD5xUFDKSfc
0UQyaAR04M9qx3Rjxm6epTG8w6GR40jsRa7xN4Lr//bQakWoHPU6gbsbh0BgVYsk
eHwnIKOtKoYCollJmvi9aG7XSQiez83/Cyf8RTkbwdWOyBV0t3DCjZj7lPulcClw
YWUDn4cDkkkpyD0VeeH+/XlcLCl395c6JZnHBChI7sXaO9q0kkm6aAhpYQ0eeiIv
lMeF5ocC93DeC3ApTaNkz/nBeHjn+vA+mGCq7lF9m7P7lqnereik3Ck9Y2IfniNF
r5sKFFrXDemsh7r9RHdWKKbY1kg6P/2X/2u5Jqm6f2rpU27Mhhgk+iuofRWeuibI
XtySWReedNhy6Q5DOvm8AxMoQ/LfW+NSDEB7XhlGdAAEZWcBHYqNqmAv5PfJNhmw
g+jSe57TfZS5pJW25OfZFkLVGqjjc+ecLsU5eih4XjQS5lLNaZ/1/j/TzCmsCQQc
1drVTQdL9u8la9qUBxVywpvQHm66RcA9aR3my0req9sx3w5hOvsH6iK2fQI6JrV4
F2zgc14b2jYDu1EYAtR4K2vhAnSYOiMAtTE4RAm0+wfgLfu8KFxapceEE9qBlB/Y
cEfOZ4MZHef6jGVxhRqTrnD2a3j2b2M1tfg9lCfNO0pM6gs/GuUpwlNvuSLPlZ41
061mO/Z3qxieVAVytl8YPBudlvSQXDOwv++SCedGgsAtcdx/fbC/9J4qb7HesM4Z
ABfV6DQZh7R5aB2BQces+6T5AdHK7XunFfRnXSs1cuJaItR1a1kAT+QFzwuA1pzK
fuGKjMi8duNYGf0y1RZhwBBWXztDjL2WJRJcugejz/giEBg2qSa+SKKDcNrsa0oL
MF2h6cYO0VuNC0H8Da/U8+1eXa0TdAn5tIRVCOrVFbZZuwJwV4TjS4iyWY7JpCpn
bYschywf5QTGpXFCUcA14LcAn4htxBwF7ta2F1+F+ni7x7ac/tZUt9+KnX5BHIF9
ZvobWYXDb/yNvtJK89FZvDJfIzBjXRviwiYcxF6LhtpeqaHPIiVCfoOIbEkxlri7
OQkconX7y4fhrIOpQDDw1iOzsDhUfPJyUkft04199kbI41DwWjr24vK3Jt9/AnyI
vHG7a4ZHrRsPbFNGqQxN1PLtz1cqzYYbnlcVHn/qTrpXs+n7hqh6YVq8GkhZzqt0
JwAsCGuyS/u0Fl09b30B6OFF7E9FI9zAHyrXQlmWyW095ZiL+H3Q6GP8LTgQWUxW
0yBvbcyxejqB+Xzmj8qx8o8LDkXWJpV8nDfvO04VHN5NrQ/y4xOaXKr3LWukCD7n
mJai9KNgIWmh6yTzhZ8izeUgaZcLTmAP+B351LVm3ndyk7dBo8YgU4gePQaQaAm1
BvxoFcAZEHcDX0byR0uTCpEwM2BRCd6f9Tp0dcyejxC9R8qFTeWJYri+zM8Ytma8
uVboDNBAi8BENlmxJ1vhlhzFbtCzWcKNLmPIAX9qKorKWGBcSjky3voHMp8zGlxz
ZQ9Qn7vCv0zyIRrtFAwx1Clh787/TxuF3Y681SUE8/qQAvZ0/+Wmvg5t3rJvJv/F
J4aRlDwqD0246gXYwbPfzRsJGhEFy8S5MydiVBOkAlB2TlFN6PZq7EtoP7lY0AMj
Qv7lAka+0oNTwBYizNBhPQEGPrb5uF6xrCqUQ4/p3Era8XFJNJ+NNG17HYsWhnEQ
iZ5fGY0vfoTL/3M3weuvw18gHuemSrP35tYUv+x1W17hrsFDz5xeZaSRqaq5RpjY
ICqVw7wq+Aq1nFkimyeKifbQSoM3tjWaC9rG6sky+35sLcF2eqch1XytkxrLTd0K
8l2VqV0Wiv0VC/N/fSsuqAJI+yQpJ3vwFcL13lD/9wvrt9k88xsf+xDlkybaNXLY
cz+nEMJawgDQ58ZaEjVGEqL9rvtiQXUv++Q1BEM/JVEid6pAZ+UYY20EBX4mp8le
c7yycjWGtufMBoe+EjOEWVyaKKXfqKzX13MokUL8b/qN2WbzI8r39oSHEM5Ww565
s6QMM6m9VJq524Ez8pKHTgmLmq2KF6Zg3lkn93LsZtq2Ws6Iy4E5KJDN0+jfsvLz
2LNW1O7AinTO1hU5wKIUwNPJF9fpp4d8cskqp8NnnwcFSaPi0WU4CEbC11tv1VCj
1JfABXAoxM4JX9+EX382x055haQOSgkqwLzNNEvO5WbUe8CHi3KKFX8+KAoJyIy8
nUGhKR1D8Y9uKWxmTjlxP+boSGSE9lLkTGxXwaXI90hdzKWKBACKzw2XW3E8CxBo
/fmodE6pX/utKnZyFY4SeUT3MlKqNrHMuustcNhIuVQvQGbKbFIWY/cbkJvnxpuN
Fj/ggeBr2uHYygvy9UUxj3k+YK247NQFbeudhHLrleib33i2XkXy+eoG1ZHiTDhj
CTXBJtBgoVe1dOM853md80B7Y1Errd/JW9rda7BUzzOdMoIBggR7U14+UQ6JJmiu
A4NjoiUtlJbkcrYRA89uMQR1qlx/DjZyZXC0XgUqwrPjcbAaJUz/9hzBSJLpcrPV
Gb/O+XzhOLtWNrnj6Im6Cyd3/qRtdrUC73m0oXMjk1dcLngnwu/ONW2SLfgZyWSo
US3nAH8s+t0nWQucdoxpQmM2sx3l2NxRaWH6HU/8ZjnBXYhdhTSUlQZVXilMkhRK
+qLOGpq7WK1CEhu/mZ6UE4GWcC9s6/yrwG0/Yh17xDlWmmuaZoYmX89tD5ZhTt7D
EOAdUfg3NPLINdzyGul9vV7qfn6pKY1nwQ5W5hnIB/jbV3xZDK/S25ts16P5doXI
J6qxHAoSBm7cy3fq0mXMqkKgoZ7CYN/kjd9l2fgX+32UQJYCmGki+aoouNbV5Ybs
yeB6+fsrrLr43hzY5p9iOeF1TJnJPf56TBAopcdIE75BTuf15CgB1Fun/mYv23If
RG/KEfh6sX4qQldryMvaX1JyGG3lJGIHpRByAyLpobm9+zEXNOzTHxCqbWflRzmO
A2iSaD3dJM9T5yXAbewOn5KfEo2qb2QxPj0C8UFEg+nUMRvimWqBmM8fjzowSqzN
eBjKHMeK2cXY8jYZbT584UFqfhy/mnsMTE+5125HAGV7MjQdvSP8NGwcpctrD5i8
xTRXFyvpUmDBJIjB5kbjUsk/iDO2I0Sxdoy9NrG036RhCrGwnYYPRQV0IORWPuuA
JSDT/pcMSHq/+6N+bhpgkXBfpVQs5i45qP/Z54M7meeapfMFon/X/tDCYfRC/o2o
1bKyiFWerUS/8u0gQMzTrOQ0xI/ub8Vzpk9Cu5fNt6cV8kI1l5o3sqyBKi0Zeon3
EbjEjTKnX0n3jEDxuXaQqKmHWLrA+/upr5isNzzvs5ZatXnXolUzr+DPtzTr9JwF
GtoE2vk2lCo4OPj1l5afwUh6VybUP7z3fkm6MT6K0FGG2fDATX7WoZPiBwbMMT8z
6k3yKo5w/wwZi1HhMYZ/DmSi22/KQbcQJgcRgbGTXYwO4NWIVfsiBh264181DjHF
MbHBCnHW29BgFrsj+3uYT/YrJSDdUF54py90I4cFinwP7QRpDy/QdXY/0r+umdOm
Sbi54rIySY9TUl8zGeIHNVMQvPBwmBtSYNq89+e/MWdpOYmnDC0mzEIgLZH/xoBF
xYVT5T1SGIdbKCijYAMMpFB1HfhpoZwZ61ILsHXZ4F5NiU4560ySYEIqMuNUggpv
SVOzniBEb7J73aND+0f+gIX1D4iM7ocpqWyw6bnyNaqtNp61XKxk4lsslJyitVWX
2rKhn5IGIjkWQnSTO7bRq/a24Zo9THxnMDseUGEF+6VAFZWfaQ/kMMdqrNGO02bM
WvYZdm68WhDjL31UMRJnEbuJo0cGEyRCLKcWP5BoWHy6gDz0n7s4qLeKkNAheu7k
Oksjc8JyDjMU6oklO7OlIAGku/ohvhn/cAlfSO7XtSogoHbNbumFTKIaf2uWwW2U
havDcyOXfni/1jnFe4grvkbCSje5infcfCL94lBGUvr6OjU5vogt28qaOk/vPrjM
vPj3hE0/GyC0KXqvB/5zlEZoGt1n4oNDcqTBDjOTlZWQJsant9MiuE3S6JFUgH+I
fImRc1aFnPjncFklAu3LnPDTkD+Y3WtEy15EN/5IH0gVu70kgZAWeOpT/suydP7n
INvSWM0gxJPJQCIR8Ai+/x/738A5c4CP3vNmp4HHXa5QJoN9pqnx8m9VoEv2veFb
e2xgBixFFBh5AHDXR+ucgJ4c/hHmUyUxtJRy3a/eKZWXZ31YpdD/o+dkA5GD7DrX
p7GRY5gI++liOn8ExN46wESRO2w6ei8tXRW0DG2/4KUBw5SrDrNwCNUqFgJfnbzk
TfDubdSUD1ANaEY8+uPOCbaKCw48tf21z56syr2SQ+8SR8AJqiLvOhurh2WxeX9x
tEAJmEiFTad5OSPuPBknaezQGVkaZen2eTvh+TED9bEy4ik0amDPrHD8OlLdPyi6
QYlzkP1R7VJRARnWHzEnoA/Axql+FchcFEigAD8LIisAfptMIvxtvSLpmDOjHzgY
WDeA1QnCtIpTUGJes8OtXYvLhUOZzZj5yOIkOxhJ0YUWqO7TJXdV1eBwtss+0xKR
FQ2g5+u5OTFXJRVoIeKq7EhAx+OBxqrUEoj1Id7CzGfyTdSDGUDq7fJTAoWWyDrv
Od/rtT/9BFQqPUwk3PozVxi1yhxJf0XD0Hj+Y9MujiHyXMAm5vTVCVsbq5p+K0mn
6dg8NmIUEI0Ip8CugztePTlWVFJ/ILVYiPr+MDwVcpBjmyj5RphFDpI0qhLIFEAg
pBd3Egbc7gt1xwtFhPkYGV7RZTxMa2oisM7ht1Y69tlFRG3H7zbWWJ+t8cSTCQ5T
LJQmpNti6KCVMHqT8Qa9qrbrG5GsXl2HsE7I0eqHQdfuGSRPOx0rq9cPx40KF8I+
FeOJhvjPc752ohAcv8WritTLAzL+MkpOjUE+5EqJ0aBBcF4vPdDbNhyDA3eBmpU4
nBlnitGYbsBFojsJeFokPHIvZFOfs/etTCscUb/Dw+KWyPrkFlZtHiMyql8bmE0F
y9nb4vML6tYinhNFFoP2hAw/4Ah6RX4L0WdjRGKwAKI87oekHiG8AhGRNoX8JR11
459eUTDGBjbi4rueZHfoDs/2jfvS2+rkGt0RM79mP0L9qKq7r2n84YgCtN5hyfzL
if4xl2pFf9e6Jj8cns97Ss+1D17w7LYXWqoXHbIzIEOtQg7Z39czbaSWb4PPb1p2
ViVpaw18LTjmfP0+uszanjo8RXp+ehqNE/67ibl+KvO6dtY35wYtmq9PxBcdeueA
80fjJGHPQZCQPLLlHGTOjazPBrJDnbCq5HqwnXvXePAxdbRGf5kGB1oTqMlK2SD9
84sPIk8uqjAps+fu3PUHOtXRITzNYjvGS6ct1HRtYG141EVzgPRdv4X9gQq5VBDr
O0vpSdW/jSFZr0tLVtSa27iax1gH+lpJk980qCa45EO4vqdFmyA8wXml51MguCrr
2tolP7Ckuk9cEYvea16ptYFLPbl3UMV4vXYOfE5uCuaC9LDr30UZKG5RHedGLaj2
UcX65Yybq6+IM6/JwNxSlUYr+EW9L0mkeHWVXog9rYYcFKmt/uBhLoJ7fWBvny1f
w9ujNS2ggBYZkU3SOFWL2GiLB8DU60EaGGcRqvOy2OG/6PZtQNv0sLuXea+xhq/a
wYYin6aGXKnHyHfIKB3hhIJlHHNmFqOx0vZ/yTvDxtGOIDhBovk6Y0xZz1GuBerV
XwmwvThNWcGEF3O1Xz+N13XiXrgeyDblNZf491H5gm8QEOcIZnckWNvIe4Hfn9LX
5plHzHdbHei1ocMaOCbO8RZfYD/Ch4HXD0izo7hYWW0v0EvMBIDepxu4ejfm+3ZL
QammhFv89jnJfppJ+FhwFWLyofjHpt7PP8Zwm7hQ06oQDbnnf1vpWHmWkkCZsOPm
KF0s8RBRryBWSu+H+IHOTdb5i303SF6UZRy3hdRjkO9S/xOW6v2mKZxFQJQvLN5R
3Y6Hi4WoTuI0JMP3gj6G3ZQOvCnPMXVYrNYRSYSnqDQnAVO6D8pLTzdcqs3euTrj
s0QtWdz7OXQNcGeyXDIeeRcVfU8lVn6MURd7PzkSQjuHfz+xNp+L8jXu3bIKC+c6
C9xXAVJSrN94aMY5QB1G4KwDMF22MWohDemsnT+FIo+c4soHd3GHYZV9ZF8BlIPE
oR49HxhIPpryHi+vkcv1FBg49lzNClpq6kITSxcewAWoPrNgWx91VNuBXRezXuMn
Lv1gjG3thBh+aexBk7CSOVNDvWk+phlpBzEMlhBXVD/csgy7p9zuneD/TVSZNKaq
9EPOoUb/6RI+2//n+BPHOKlGe1CwfdH9ii8JWQrm9jB2UWICwiVtUp4NcyiXPowC
feIdkgklTMDjWlfnbL1vxa3TIrBZ7gAQQkuo8gdoT5eAFHgHxPUBBtNIP4jgFW8r
LEuJXCxXY3/37Qqdus4CghwfMy3cv6tjbgJfnsoUqG9Pl1ac5WxPcXXtGFn436a5
yXKYv1ELRZGjCDWU7o/PH2God+9wIVCV3zzt+JlUr9vALkFCfEX0paSg2NxOcq0t
6h2qU2dQn4xzjqouFcJOklQZNvrVvwYvUCVVxaScvYQu2emGXtV0Ux8Ncbn9ca01
yneZatCklQd0uG/D5IZY1EO2eXNHobnNt4ecpN6ZOhFxC39azSsYYAhaK0HLJFTe
h+rPCaqCz7RzD640L2wcf6/QwhQNLvpfcOPF1vtRRXHD+SIyUZ7pn2RmkX4oFbrf
e7VOl1jBAZk/crfFAA8yPAWJGNfQqrqrvOIdVywdMRMoykws5Dnt4DO6xNaHLhap
aAycL+JuyZUno8TcMTbA2JrYazSH60K1kDq5To3JIsd8yHWxSGPAIo6msnnv/8jM
8e+AiAObmizBTB31IYdc7G2fnmsxHoa7m2zj2zI0jvMlanqGXwBR9aRqBu3NFMWy
+zyh0yQs3M9IydhvI3BIyvD/5GgEOH0wtqX7ZbLzSBgse8EDwjAGUAv4kSef4QEu
k2tw4UMlVsP9VqvDB/7xM8ziz/oxknR/BmwLIjPTmclS8OqQp7j+w287BJIiZH5z
Fyb12MfoX9gclUHoMjhZ5/DfSftUXo7vDq9ZygvubBdg7i4BA0RHP6MnV/JQsDGD
PS8ro0j+arSHQDHWwoF8ZUrWg9NMhqtLatDT44lh79VwrUys/K4z2olBulNeeBjL
F9158X/mijNJrWouYB/v67MLxoG7dU3ZYbDHzKEFlH10ClcJ9D9heRi+Y7c/JW7r
qfswn5u4sRPVrcsLJqiMZoEJT3aP8kA5R069+jmxzlWKHXT785KMTxcTyaXNaNdZ
y+TUaw6GyrUZJBm7sHDQbuwhzAjqc39jj+c06H2TZYMm70OFordfkOFui/AIptnE
TWSgK+gWgi6IkT4wTbV0L83QV5YsEL096/FT3Y/Y9xQI6+Wq1hvURBlA6lUuaY2Q
5VRGJ9SmBbpUf+O1fVXLg4gBTL+6y9vDz8Tu54j4apIjDq7qgCyUf662i6QIINF8
r/JbhNtRqbINniInq2mJfMGasIWriVWOxoUGybX749SyCFAsBiodFO+BMAhM9uhY
7K+SqXS7C0PbNzZv9U+pajfN5P+tm+FSHmSpnkfh/q/zUQ2g6pKBgpBPHJMU+Ycm
6+CjtF4yXcrufxv1j7u3M1ZeNRbp7t+rPmoXyAbQ35x1hQi/uC2cMtWvxtRnhIE4
7uXoRFdAz9Ol8TsQTP0KcmP9G2QYyFMtIAHr5b7JEd66G+mSiCruWb0Qf+ecvBsO
9TwzzaEVkvKvjXczOiEc0gborrpBEVm0ile11kZ8GE25kk9816GlSUeqV/H2RHba
7/waCn281zJP96B/GtyccvamT7Vdu8lTewueUxzze2EeDMl89OXmdLW3HT71ISaa
THCa1ht43ehgXutPljp0JDxLRpYhP9irdDj95hXjYTXjL/bAcEUgRNlvfYpMBP5J
gwmJbt0ZFKC78BAk+l/mfnEBdT18848MssGg68K/B6k8SsyCF9FaqhMvfLeQADHP
XjU2DpHn15aBDPRkanZhAKHyYO83vwEMCRFnyRK1W5MD1RrBLlYoAQkAb+8NC/6/
ogpj8/1aGFiX65MxWnPJIM/MtI6HBqSjd+UNZvUBZ8iGxBtbcRm/veRcjpwf8GuZ
cqWdCJROZOZWvPntnd0bh0TbIdQEuuXPGL/tDgsJsqvzp7dVh3ARBRgGwMV2HrC8
/Gr0MBMigNHTPIdDIVvpISwvvSWnI5QIsdkIVgv9p3HaOMQ5McRMyaoGp3505DH5
b20kzFxzP04kHm2iRXBXdqnS1NCN9ig0PC71LeS3DLazBqS7h5TrtlGUQXQQoJho
qnUBVv2mtGhWMQRVhohsgUsK4RFhfr3JNO70yojNSoehDZchgPIXvP2Z/VgYymMI
Uyf8lmfgNcya9XH0BQk2HuxFihi/JykzOC25L7NrENSjMWavAHme6afLIaBtW1HF
z9TK432SAkjtreq4aTlYqmD66yNqsGXFeSZENTI9uNQMnDg/q+9CtlFqv+92aSOj
c84sepogchdwjcVhXXSxjOE3CatBiy7vCcz6JvRg6hfiwURHsplb/6Yc0I7FAr/1
g9cWZihLxqflYP0JvQuAFeR3CJYLLXuJ7DfKP5f1lvY/VYcKMWLq0GTUcVldP7Cw
x3eALiU1Xs8BEChzvaPgQb9w1BwGmpklRpsfsUvvfz3nm8YzQQ9qaqHoGQ2lMyPN
YnrCZEvALNMKsxZDIm+n4lVgrPoGt4Fyrcw1fQCRrNknrjIvQXotwjN+iaij+IQk
WjuPhUQKHjbQRhFajD3tmXcjKRgJiQOqocvYR03pkDbfHk+c6UelDoKBNggU5cO9
WsGF3fVpWPcr4vfXz6Loy+BqMbc4VnBeVKdCnKn1PWue/Qr409X9BfOta8Xai313
PiPdPiQbbOg8hKHF1+QMiLCPmEWTNE2NcHQsTQQwUMMoOsPjdlRdDii3OeSvLXLc
lUAiHWD+cFvpn3sMblcd2iHEhz2m8rVYjaCBnSBwh3dcuW7N9GbckDJwdUA2h5Kg
HjQzfFkS+pg9FLa9ROXYDrhy/EOHO1ClDgyePSbc90PSMXrDjSsL8RGXoulJFRo8
UcZF97UJOY+Mg+/FKW16se/8bTFa3pdfE8MCY/AC578aft5OvVDIQzZ3jCzygyOg
AEpPlgFuT9FWEMKvab3k7s6qjNFSs0s6UPMQzVz34HzP5COuZ8W50kGeyUCtUSSY
iSqqnqhouJXGzR5zwLb5C2fTDfsZcyTqNH2/PPs7GOHar2k4EL5wQvIb6CWDoxId
B/R5/DI3PVmvLdRuTDVlxgSWNp+wVPLUGC2KTCd65JFH/D0O1h8vvShf/6IUqtJa
c95XzJUvpKrXVeGxdkSM2QySwsA3L7lD6kewHkgU6QcNhsc9CVmmCYYUc/vgy0NM
ZLW5403mQvFNMVF9uF+O+gLe/RLdVq6MQvM9idV4MfR9G4GLHnoNqvSmEMjERY/+
NOQ1+64kyP6WA0b2sUWBQmFbUhSWC1cb/9vILNl+MFdcD0400cGg9Gt3XuWa/XUs
q8qZbhOkkic8c89H9oupwqvPUoKvx1cPA3JIguk7ZsidC0TXP053q9w6QEE7jkgI
Id0PrpOCxqICMjILzx9rakgR6n3q26x4wIcb0Z6iRct/L6dDhYL+p82zwnoGarwq
60qmiJ9uXiAyOAY19BycInVebFhMftLineMbqr0iUbKbX/VnYOgJmkQUgo1tfJ0d
J2k61vVnVhtXoHeJkjOk4oPcPUYfcrX4o/6G96cN5u2pv8FJ7D1VretA6CTr5Nn0
CQg8j6akoZ4DX9n6zsguKTHtzShv5ckecsKsPn1dkdOBesXlXho7zyvwwiQDRDx+
8eMSbQCMeiIwzLKC1vhbkfFf0s7N10TeqUhESr7GyqCJc8kiRw9dzLpp79Sno3rU
3G9kLNJZcqzPxOV2fQ1n61PJjudGDSC/nx9Dafeiw0DbqzH5GuVqk9rKAwPUfmJi
N03wirUZ3RfKg8yicojFHVoXXl+rN0tJSL6UcAjwdbywFm3JgYJe0zorBwPJtmS/
pcY+B4eKDL33XhQDL/zZZ2FS/xb7lzjYTsTBkcshUsSVuytQgFKtynozejqpishI
iybS3/fZnfSB6/wcksiI1DWNUgGhqdh06HnYUmqdVvA7LJOPSCyS+imNGokvQGuY
DTAJXK55UWjCR1kWSX11bV6yd7kUrcSa3rEMLgLyvUrOGuii1g2jkLpfIJdvzxuk
mV90IyCNHiIBYlgF+rjiSAityknLejdD2t2uwuj9Y9hXSZJU7+MW+wdbMIiaYLM8
4K/KXmUsiASlTt4yOmfz8nRdq1ZKLzPsNi/N9Vv/jldDU1Yzz8u2yD53qWe0dBPv
F0zmNQctiYNfxLui/BNOB3wrQ7ptnf7jihu+DgKKgSh4zqM89OlpGJyLcoylsqJo
jZkFM7zCrTTUWaUQ37DGDVmpfCGfZOey7ULA+av3m75mF6kkEi5GlpHt2SqK0zIs
mS293qKuLndR0PQWSVUiA/od0SsNclvXiobfEfAS7JvE1ip2P95pkiVge5+UjFeQ
JvYPLxzHckfaxvR4knFSD2Ka1dr3deFepPkmdz/p3jTN6+BUQ2briKn5yr2RP8tc
RNcxuIoYllsVZs2ytY+SxMeKhiP/tou0pf7kDclvZ8eQykAWrCnW86n8QnnnvqT+
+QUe23KKGcWrVAp6VHP3jP+xvsxhMEdxgxc/B976oGxDlr7UUJSmbmSrLKzSbngA
+OlqOnRSxBKERRU0Lcx1Nkz8uQuOn2sXQqYxtlBdGiWSdTuTEVZO1mFZ0mmdv8Gs
2v/HZQwxBfBR94Uk+uPvfYmTW7KPyCJdHDgzH3d2M6MmaOVHiAXuS1LNZZIokSOU
xg5LL20lfrSofgCgqWjJ1dMozwHomX8Z+FgpYLgRKbcFU7nW+Mx6iKMqd2jYglWk
AFffjbKsClMPhBp/nRh/O3ETenWWPOCg7upUwwGU5KliLUnVUFBcftcQF9Cgsfyz
e5lqVT5lN3NZa9gBX9X59AW0XkGVoq/ySTnywPf0F00O7WJIj9ey/llHRiQ4GQTv
96MdUsgFj96yrap7hszBhYA++6YYxz9lINFOHAo8h93Yav7ebc+pYVMx1DBk5exK
szu6ZkLeMDk95+Ru+INTlHi1HdnvrmuQj2X8rMssStBdCorQBFs1jfYNJCgCcUS+
LENaAPOxwmzOcxSwfpIYU2LByr5FLo7MPjJzEmXfUUerTdUgl9+UjYoQcDySXnBk
35NhkQSOULWfg/FoApGbmjQYM8taTBR8VTuDZ19qXnl1120RyzBydPkuFgoLHGfB
h+U8HQpWwhTcU3rs+w2TD+XRM1ojzWIgO7J6zKnV1KALI0LdDuXOsVAOdM29esMe
1M/7nI4p5MNj0d0ZOn0r05VxGuzx/SXmf71Y46IQCG5sdV/27tltXwRElf4di7m1
hbBjXISgOeAouUVsh9yt0DN4OYu008H91zoEKqao1/u4lX58F+8DPDxwAa95gAQx
vWzS4GzB72u2ABFmoe3vYKibTtp5LSZmFaqLzyuABiOh+MH2C83z9OEV2JUjx7W2
O0Qz6TvjFEvqRGeDwX80XX8iP+r7hpuwjusav2Uzvzcy5lV4neDWP1zkpy9Jlr7u
8tIikpJ9sHEygBbOU0ljiAeKzbTryhUS3mEQhWXb0kHAg2PgyWLUgbWDcy4Sugic
9XMEAMCLZrVtFw7QtV3PBpDUF/N+wPwwifT3pA1qCleatZ8KrR/nHHolJDE/OvxX
XCdFlMQvw9i2GDD7f6sPtDb74rW4Td8USU9xtmf3zQlbSyzXj2lrXss9YLt1xu8O
hjxRtTxQ/Ei80gFwDT7RRmVJY3Fi6/u9OSbrHUkgWdT6aHrmsddYvRtlciorUCJ4
r7K4ofEwns9IQ+eFghV3RzgUKlC6jME0wZuOEUtIYteyNpCC6t67WwiMMYhDzexv
9fWJtnlI4rq8RU5UbGvu5m20CpIUgZ2JZ+Gff6wlELEjdw2sz1y14Hw2+VQJnFmP
0ipFSEcXN4cOA4agLrwe7AfXj8gpAQvprB01SYk09uac+DJkR4ez1BY0JObxthH5
izWqI/29975gxjvK/tksaLgTV1i55PaoUURdJlnB8n+fzs8fqrsOI1xXKcgOJlpv
DAgxAydBAd1ucEj3Nb5MttQwFrJ1N5GlXCuGS1s5C0cPB+e1wlopgyDhHcZeet1j
PeqjFaBoV3YiAwCy5Z5Cccuxdkxuvpaq4ZzJie3dkThKvdbmA1j3IBoutHfsYBxr
LmO+VQc6+XPOBk44e3rXY89gap1qFJkqB2np+aK7u/N4gGTdpL5BaH4ZE7qrzMYu
nB3kvpZYuyqaGVQvTJjkGDxBfs6gJ4cfUByWiNT3JPWPDCQ53OZwscTY46cnsI1k
6O8unTqGsuVZbJoZGOR/5JzWtU3BtyHXmKPKoK5jwW/ryvOzsEJsR+OYyxUZdBTy
8hNiSbozrsk/3RAwrNhEXrRNhy9ofMxoaL0U8Z8SexrbJT6ry+xcG+9DrE58wSbI
/Oqj9E6q3Kj5xYkd6yV6NkNjtFH9sGga+d+NU3vgwnIkt5Gpbo5qTtQhtFdSkumn
qZEy23xaRAsjylco9hp00mI5M2Ml13IYM2feQVvd22g12gX2/cEVYs98cU43wxUU
zF+fKYjPNmRaMUpYWhKln9bhk5WJg5pd9DtspWbUzPm1Y64v0ztkVgis0aCjm4P8
iDEXdtYPKM5CKdfA7HNg5zjurgk5i1yNC5NTurgSmOT3IVgSwAjpztf/4UL2Lxvt
1l38J0f7SjVNrfo+C5fVk/sAxuRQ0b0veL68ix5r6UWiY41Tf/duBqyhZMlUNLQx
4kLBvFCb/6ejhR2rgswZsrWFQgtp+6tAev2CGM+Bu0IdF1Emak1+ARwMJf47FLN7
qNjThRpHhoEsAGBVGxPgNjgACOGQsSxlQpSBjtExn6mYMlD1QPIOYn8r9LB45oHL
Ic/sSN4z2//79a6WboKfaBAVwFF+xLt34Z5EiU4Py2uq7Ojslk7kZ86U0M2AbRe9
elZrAZuD1BL5VD7ySCOE5rzLOZUN3DMuHSFVQxh52pVQpBsQum1ZydL5sNFiZ21T
vAzEYNnt1vXOauZ74RjZI7JUxKfmj6YKj6F9ixjo3HZD2JxW5XhETw1R0a4BFgQl
qqGHy1oI9Nx83DUzR0FGBmy1x29diDFsu8uaGcDjgrKmL3DW1aOSNftdR3LzfpJo
iHcH8EVpNtCX8sTwPL0Hqv3E9rmWQIHH6z7vcDsI/+uwq9glmID+3QR7ObPUmX7Z
dHYk8qVuTAoOI+pMWSG8V3cnDSRijwbjLIbl7K8E6gv0BotXbMNibhGq9hhxhYAg
42/aJ1xEjFA5uZpX/5q5kWCGJ5QKMVSpfraPnUl0exGwdym0KKImAfsisKWGQ8yP
V9h1VsmVTQX4zpu7IyWpG0HiAInCtliZsA76E1m23CsAyLtUqJpOVcAv7tToImkr
TLTU5PpptWQGGkiVMcPj6aYhRKEctLDA/Fs6BpyrVSVOb+lRdeT84ALwGwW/PYQe
M//Tv7ZPYVpOOt+HPF5wbr3KTR2tUD9ALcn3zykUc0d8IJmvGd5XqPIGIfHEbB44
vBiFE2gKD2iVdqXUDES9dkjHPtQ0yF1Tv1bnbi+oovnRKCNlrMLlPml5x/KQp+8e
C/GyPq9EJjSKiK9jO85Cbe9v4io3rgu97onJ1U1TvBGZg6HXRVRq7s8wvPQBJySs
O2iQOjJ0C/YdfbqiO7MzAPr+CnKVOJbDvQstLCcQ+FXpv4i9IVUgbDQFawdlARtS
QKuKft6Qx9MUf7O75SJ+0lbsfCVSToC3KnHgy/6+1zu9p502Fah5OIdFYkgW18TJ
acBIfoSVjH0WMM41B7jimtp+kXJLpvGRZF/J60jAtftuAWkxwsCd/zpKpLDknIBX
toE6IYf9AhzUq7HkBGKQW3tdBfaLA7NtYFuqIRI57gXoiUCla4P8Ntyry5ERPIP6
1FglXT5g5RZSfnkAw2TlLB7xDxVQbtLnpCN/nKfzUKBpkz4H0LKc0azYentZokZ9
cF+1ooklAyUeMbQi/gm42VTIW8EljXbK3ydXhsoWhIoei16HlX5hwxXPOoSTvjtP
c/T1QQxek8Q6f20IWAvNPNj39bRZZI6o0B6l+/vDp5gmE4RbSBk6UP5C5xRfDtn0
RRldoZvk+jW29lPyVn7I+4AGUo7HSdZMulxdnvDcmHgJsbs7yc3M3yZMIpEzv8gG
/N7jDkFMr2s/CB5tM2AHmrIuwIyO609ucbH7B1OFqOjB0MZPXvwk5gOZ6YfzFyqf
eRvITmltA9yvNH/W88v7mfR+KKpjMK5N/aivBqIxl1elGsEFnWtTx5fv2BeZlO6H
3Wf3IgpjGjMhkOkQWKflD1D98FyEteCGuAbokwXSzmwXMYKJA9+4rBfGy/irNtvg
sau7LgEfn5wSpY0PoGiP1jSYGDlIXwTbOYVef3g0AirhONbr2+HMzqsxeXSAsBen
qq5TVlA+QrMakzRIdvNA47jWeCJCITRb2xL5FJ6WV5bzd3MbyRQE/EiqDHH8h/Mv
xd88X39j66d50kxuWt/s9QzmH8uXDo9qmOf4kP2FlRrdAjrJGlbmS15+LacNutNv
0AeAhwVEQcXPXIsgDBBfDC/6yYZI7TfF8I3xoW61nLyBGWa+zcFpIgoZSr1XygGV
+JkXFqUk83ygafa3gUz1mKgjgtUMrsUW8XRHbDmZCx6cb/47URc3vZtWy/egejXL
80P2M1SrNpG30ayp5zQWBpaM01XqD7PskTwNgG2C74ojm6lQRBtRZ7Ca8h9y5IfX
xc+X1ZCMpuQdC/Osp7iiWsZ7OFDLXuW4DpfRtVnYUGJzcgpuOvJoJ2D4c127TOxB
E8hsxET0EqQVHfbuoS6ofd7Q96HLLVZM+Fi+FDPjyRA0KjdYypaK1vvEepBBuHxf
nmScopEZX+YZqd5kAP/S/EgSRwO8Hk3rJtSzB+EqsROAap8FUOgfbayHmZFkH833
BCjrFJymXhaOtmMvVQGc9T4zBvDKsr+00HM7wY0iuFQj4mlzIVKmZrshQiEVTfRh
jbCYwq9V0LoUIGHoESIH/dpVcTltMJE1uKOwFK7YYCzdRyIj2d97yOKn240WFdh9
2R4EbYX3ofc9k9q9hPTt/NGkBZ+wiLTTp+Rq7vMYDwMnlNzcGIYfznfGssyBoV7Z
cRCDKE6dCJ11ByvDLHgoSvDvMElifmlvP/Pcsxtd87thk9Yw8/vvg9Drd5mMDKh4
nToF2zmA+c0QmW6om/sHIkZQ57QL6ov4ZsirAPzMkjU1j0ZstimPd9uPcWFhtLjx
8SJGlAOdpAjKnxrkFpsgChhXsrVUG2yg/SSUfRIMKuRrUjNNeN7JvAC4HKjAPC85
3JIg/7UDwdfQiELuQfn9YGZ47vkMKeXFX6gvxFKyB1QSHzkLYzN0iiX2iHqtRFXD
klyF8MfO8ED0oZYXcwRqTqOB6tZMK9WjMsAmVx3w+6yKQ21m4gnrHtl5mLP3F8PQ
o9jcKxib1nWH0KCYt1vBv5aYGbq2Cy+u2Ypo/KVpeyJwnVaNeciJ/vwaZ99KHgpY
1qcR/N95gPI4ra2qud++tp26ukPQTLOOF4XhM+y0vXjvjdME2urinjdNlEkAjL8h
K/OLozezRuRrKQGm44inFewLl+R392hsqLtO0QJASab8S0DEYroUmT/GyvNBRW9x
9UBTxGaU1Xe597m9siJiU9mday5XmR615voFS4HJ8rwAq00lJo9fxXUVHuybrfaC
zEW7fuTIcTnzJvVNyI70IwK1PEufHKvR2TAwtMEmqbmi5KxY4RjtyJKJEtShKs/1
Pv6KuDB5AB7xTlwGg0j5crVkrCQToiwjJp8jzEW0AbjnMrcWmLMbR2m3E8TWvYDq
T5X6O52bFepCZRFu37v3wcXWuACzziEceInQqa4NIOA1Sa0L+DNgTxeCfyK8YCZi
S+k6jptD7kpG4LcVN2JKxg0fnjwhfwH+REc5W3hvwvQOTtIZoVb50LKPElyRjRvb
6C/Y3NunOND+mf3DaGHDtBCUIbhFFfh4XwBKlXb2CK4UJtlXB0gW3XC9mrDKjCqj
yjAs40CJSgQG/AXYzAv1Y5TIesM3xiw/MvKuZVuZ8YpDlKF4Ds7ccLZaurKe5gw5
aVqsAvCA7eKfVMMzN8T9f6HA+THvTXSExIwYNMiazNAqI+rEC7lQA6ettBF10cFR
m5dDp/arK3XePA9+UmWODcj/DYv5ndwS3zqhhKW59D85nwsBcm/0NQSBG8QWwTMw
PSXpijhBTrY7gcxojhQo+QsKyJW8Hkq9Rrw3n3ymzOH3bKUe6SiNmQvaZ75Y4Vx9
Z9Xvju6pX1xhzlVlmTm1oaXJaccwrVtHOhHAdrj2I/7XBzajzsR4gfIWNG1ZftDY
T1tMk7yeEHITRS94e5te0ES5ylLfw8veqII/jdwaWAZEABdAiMe1NejxG5NvzKDj
oNnJjNWtahfxq0N+k1YpomlpqqJ0XnhBJHR/lo7sGBYUjyvFRxMb0krFN02uzV/d
271SCYoI+Oll1xeEq/RXDyp5oqSfUP4YAbhwmS1Tm02Li3HcGFwgWeJzQKt3D5As
N7LZXCMEwQ5AwAscRH9hT7NEFpBhNciBfd46yPodchj5EuWdXRVuYcIYieG31Yog
qV69iquFISPswA0bSxhaFxQQ6Y6s090YB6eLJ9qmIqf3uiQJ58HwUvCWyQj7wdMy
J+SwUxg7jt7UoztN/Hqv+rQsyQsfC70ryJ/qGHxeWUWag6HuRz7XPEkzZizWfnFj
96omTvfjLrvNbz9KHsBs1UIx9UvSD5Q+BVBhrkIROOvP+zKhfDDQSKzD7SH1wyzP
mfdXLRs6Rjt8YuhlKv6+aknYV5EPvifUIEDE0JJnY0zQY5+Fh6ODzoJP94S927l7
j3DJGWRd8OW+87YtSohn+6+ATjY4YrV7RuvT6PuoEvIGQtNTZtl0dimZjvBJVwX+
YWT39zMQO7dOUKN/dA6C4oC7fkB+vkBXLInGfTz+++/iERAsdX+idDvKoikU4gbj
YO3AUHmRVRC79M7T7oVK+B51lQBVLfDjFkxuq6bTpMLLZ8otqpmUT6vbrTngohLX
8T7tn7E52s080lr1vrc1hekRYU6+frir1avTeft8iGKllm8x4lXPAU2/+lR2Hnjf
5jh+zVT5Mn8Reg4bgyCI09WERAM9rA4QLD3lmqNLnv1Hr8aTsaytRwk+q2fwcKLv
HfZn4gMwDiiMMGpjjm+AQgHlBcIckqtauhe/XfO6/pBoOP2AM87VzHKzEf9i64Bh
+GPCLwMUelh3ijTzOmDHtgfV8mmiEx0bF0YpC0imTGno46JvETb35GVvS/Xtscd/
X1hfNSV6tGCQP2iDkiZZWd5JfzbwyJIzsK3n0w7RXK4bHBo32rMhtRPWVw8Ndx92
NJ/c4IRch7n4EuPpdQRqw5NLinvqph+xJdSOIgno31Hk0G9ECag3eCorIUQmGs8L
URKxfapc649JAaeDYl+CC8SUx/uzmTNN13eFIZ5EdzSbEbulnh8OtnKtQVdJ3C6P
KJJ1EErqEsN1QYk5IkDR1JwLJi+mS+slGvST63guIemvot10mUB/ZIe+wz/Xo62W
iB9TAjuxzpwNNMJEay0Bk0DANxdlQRKv3FxeCHm7F2SeKCUZJPltM7PICpBRiHAf
fpLrlbV6IsQm+9reDZ4oJAhIQo/TVdUd7w+0g/n69eBHXDboGM6M4ZsZumiXMhMR
75LLMCnrMx6YrIo97Me3ajucUplY3GqrjMJYr9sM1pJ7+J5oudVEl/dWGvE9YYqN
85V6DgTLijqdS6MeuZVwNEQbyxu8s4qqzJzZVg2lo3Hf4bCAkPUGVwGuqMFqCgxV
K91WNwKp/kAW3eLbU60cvqen7mjTFcakPcZW/fQIoe9EpLmd/8Y79RjF5EbARaUN
b88U37PqkFiYvHAutRjvKPVSlIo0y1SCXLE/wYtcipKLsJgiMXDAr7NOTPMakTFy
nuS/aQCqxbkfM8wKi9Wjhwei7VCYGwow1/M6/Tn45XIHz+icmHY8+zNDS17jW85+
5sc0y4CoruPhE9GR086or+PCV5Qteavue6g8HjrDbWahtGAl987T9FFEEFZBszpQ
PO11rCT4PJtgW2H30gD94B3fAb4+Lc6JcsirUqff2uzlNaOSeKNkPTOFHYtcyCMR
+XwqyGdurB4Y3fEBgLy5ZOdJeBi9a5EzuouLrDd7eyHArf4oaFZhOmKjTMWHqVOh
zErbn0gvK/wypvqw6mo5YoHEOwBMSU2XIjuyLmOp1/04DqbAW1LWQPxAax/ksyP+
6xlII79TeZzTLseE/mhx203ZSEhoLZmsBhr+A3tVZGqvB0lYMgFXtyV/nKjjKGNJ
s/M08uYGwOONBowvsjtQxTzu9uCxQyTdcmRGf2U2DDD4A0SteAciKx8P4DeZKviw
73xrhRJk9Hq7d0pzJtkHhucfY981IQxl5BebDSxmiZRFGkNHxR7Dwi2M+MJTpVZ2
TY5R40QfXG4WiCFokGESFh8KDU8sskI+KBM5zEKRHf7f0/yJmv/qeRdmYc+70UMn
m5Ez07jwMQAQLfr2IPYbZTENmxLc00RErtYWpl+O+ubo3HrF3WmbinyTn7TGtVOv
TMJi+QfSkHlkxA43tU1/jD7wlPVKcglFx/NrDrHU2NVm+usNljtyxJC0TG1EuZDQ
CvCJq0opdpTA9tz05gu/S7+mvVNrAKdGcM6T7alGU2nkO57mUD8UfVru66l8TT7p
5THk0DG0mIwQPOxic1l6Y0RFsvKPs9+PyLXUo1IBO2eO6cCA/x/+QHCyHoCvxp4E
X7vUyZC5e1DVtPfoe3fpe25vSQsIf625GKVEjXzjJg8Je0siWV/6QkSo/Ysx1wkf
aDK/OHdFqcIKzekDvz8IwKxJ8AwVQZYwXRU3Mj0fokawXZsfXfYsRrQBT+dX4X5S
I6l+V//yto1h5IkHhP4ebY6gM8zxhUeJzK1x6Lp0zEXAxI15/dVkkPR+gl7FhCZr
5JEjgHkgm9KmlyNSoWx0EADBrlxoZlDwq2LE1D/0mnnD/KHlzyqzeCcZAkn/j1Uj
+wEgZB3V3V+JLKQdna6e3TJwWzPxDF7q4BahZ/zIOoAFNzB8KGlbyVH5aUvQHcPq
GfhfPYR7SsRIsom/M2S1IWRWrmfvYpg5qXgQUdh/gCileYzsHBywntJlVHdRgHSu
UFIshJOPau5aude9Ou6+7Ft6C+9tI7Il/mw1laRT09bwiqx4JUvtlCq03Cghr272
WKr0iZVMGlfdkfH+zXij2jCiBXdHfyLttzxUKlrn83rqfR2fxYzX/rGugcmAo2o1
stCM+OxiVuAMANQitD9zRWfKNgEL1OqMX2Yxatxlck5hkaVYAZrhkW52TdlQFTox
YCK3sEEAUiap9opHKGO6gAqrBzlauMnPWn4kAH+4Me0aPYyjtCWEDgGXbFKNbvUh
FWP1eGfpX4TXuEE7CZTK03B6bdSL4BEiEk3/wvBbrUWa9nkee7E/q+jCDHLzYMTF
MugVAqcpLlSOZZjCb8CphYSdnWyXmVOvmG4jQi6aOgC1/cggg8DNylbgJUgpEO4V
u41+cttnxYvrJiSCeKPDlSyYoDhC1Ifd/IY1JC6mGnwB0DxeIQo18w4zNxX9ZnIh
FqUJuXD66VU3PKKHTBpWX6fzzjzZyAqi1stYpaP0hm3+sr5yW1derXE+fi6wy/Hy
IXU2hpb4SBdTQmUv9aoFSpQfEZlaSZ+TKwjI+vUgw1VUtswSuTlNl/jEF4EQRWYb
K8m2CCRpeVBIh/Dk9PLjMtEetDXmYFjqU270wcg5WNeCQdYInfM2pjAthuzPE1l5
nsiQVqpLBwm8aZL/EkKeDkIhvZm3eEC5YEmMfTtVgsLko7DJD/EHIt/EKjmPeUFh
p6Gr3Lldk9H3xkmE91AegWG+tr3wDTeSt+HsMdJgCdDBCGGJijMsypYTmHHRp6kP
FRLH0f++OATRiS5ouyqqrm0SrvpvkvYbJq2E/7bmPXXNlD8hrUm54Cm7qE1V2y27
MRBQH3mA9x6ADVxVF8EBRfjzwoB+dSuoz10tCvtbYVDrEhXcvoYbCJGIuV6YBuAz
9N+MwnXcmbqdSA3se7cRVWUENyom9V3N44cW/SCoz1P44s7aUHcnTRr61zT5PAnH
571culK0qLB6oeP1IOz3N6QcYY6pP9TRGfE2hgFI3FIboAisuSz9ccah1Lg7RDmb
WY8kLdWQJnNYySkaeviS4NJHM5IcaB1KRNKH+BAeRiVsjwtzEBp+hV8s8aGMQPG7
peWE0YHnHIlQK7v4GI2MYkJzY1EOqICq9+H60PxD4khY3KmF1wt0b0buh9kp2S7E
UxxjPkgU4YbElR2hcHMGXeIapQG2JLjd0oIpYaDyeHk9oPEm+Vaumf6I2jrb4hwy
ivWZVo9kcGb+g1wgWiItcdNm15LsvlDw/ZLWsoItrUDKYfcSVktNYLe+VqWwePU1
K+CxK/JMf2rCf/bfu+EyC+YJjNOoovT3itaYHZ7pF/Tyx8HyN0kCwzskrg+Jqmbh
4eDk60cN35gf19fb0QSQQE+wcnPXbi5Pq+FytPgRx+tJfpzCyoohLWmxZ/qCk5rP
nvOjVTNOnIwxclubQ+mDqLM2iwIGU2s0qW2c7NBOMKtNOqptWaZT5BbhuG96dEfi
VuemFUoNIbGMh5Hz+gDNZDhw0juxm1rbXKcFkpsT8umA3+bOqf/ACiuK206YeAkD
Biz8iXDKgoYhxVrtXaTLBribyzBT2kSDTJ2j+cvLaKjCQRvhPN2o4aCUnKxywJrp
d4BGcX6EvD0UOEm9qHyVKEUsSLOCn8RUyC/4NPLKfCODJ7yh5lJMSZ1vzlPIRs7U
x/T5H9aAj2E7B2TzgNsSewPsclrcMK2m7muz/5W523gAq7vvausJ9Y5KobsXfBiV
yxxr1axfDd6iV5LlPOwdpdzTTEjID6vzisqUKO7qwi/sRxnR8xRGh6kLH1RZ0ekx
6B6iFPquHoV8/66JW9Q1/4tdQGKX+lXKIl3mxW06i3VtqklG0ELZ5K49GA6l/zmB
sV+WLq1DVGasycVz1bn4hDva2I/j8NshnUi7caQokcB+D6JqGaFgoMG6rpoJoUE4
OOvenOy7yOCIWNURtIVCsN+YJaksUVnvCVdnOXYUdZC121y1QIPL/ZRV9BoEoIsz
9yL3o48e2YuohrxIgtTW2xy+/JssbLK5dsirF3WYp9GpRjBVVG6XZPqj1D0KTDDa
njt7IfMtBuV/xHz1oU28PRJnygUVt3HChCbJhA8bO53d2udbuCkL6SjYblowjYoy
VXCbECyV8pU+wMwZNaLSwAPM/BhpnLpLz6nx/OctGXAnjutnsZ5NoQxKqT5bQvcz
uhiz/d7kpm+NfqEvfy7V4YXtS9jXryUPDlkYG5B870bh2JHhnopUUs4znfg04E3P
i0fKeKgnMBl7iDVXc5f9/C3+65DdXlQWG9k7mi3MnZ8WgCrTlMT38qG/WzAfPO2F
obIbnkMtvCtDMJzdgiSFFgewMVwfdsZoJAEzDG8moK0uCfsGpKhA/CTAlEmYzDSl
HLMIWMfwKEJLjRokNQ2Iq6wHhllqIJzObBtKkSBh90NJr8oT8Is7IP4c7BrnR8AP
OFWQOvI8M16avEFCR3Lcrc59mrlqnYUuNjci4aqx0Ho72x/tcfl6LUXAEcWhDSPO
NG4qDYoe/sjuuoCyy3GYMqgEwia7+zzgnp8x7Jmd4c2dr7Wxg4fnhRRSWzUpDO20
+M1aKcZCWhw9vWYf1zugdOAKR/ZUwHYerCRIUNHwZoSph8rZxs47ETYNavGHhuCr
B+RAxm5hnmltHExAG73hjDIeoYC4KvW5Pv8ZAprqkfJpEN4KkLlcgrGBloQkui6v
6dNQOXZzpT5DcYrFu+LtG5iAD7tTV9SrLG4nMDAYElayY5EQw/o0J/oaR1wQrqy0
9M+rC7ziCewTbJkczeKac9kxB1cT6Vc4BnhH20YDBN9u3GG8hKx8LUgtJ6s1NJCu
MhWMbP6qPwJrxgRV38vTDAsykOXpKxL2IBZdr70XupA1mqcnEqN5G/cjYnRXD95o
Id7ESUandBqriaVDOQjEx3vfYSUMmSpf/FU2Za8KgSzmsez7CwVj0uxDNIt31nFJ
ga/fbkZedoQfvpuwDXzczKsTiaQ5eee7I6aueKVgxmliVk2rzmpWA4OfDeqmiR42
50+LpT1WigU/uYlxdmaMhC/PGeaAxTe5r3iuzir2PUQWGVs2HNDYC+9g0tuL8Zmp
cTFWopT6NQTVi1pzTo6Dxu9AEQ3k49shPyk9iWA1fSBndlziDYu6CBlYqCNwVaUV
MNxuLVg/bs4ynB5pn0MMgHIVG4nNO/OqdaDmO8ttTX8xUUC6SSjiKGatbXnF5hib
3QWqxCy/jAuKLyf+Wp+UUE6RXObvexafU+Y8Gv/t6gd5I2ePJorn7qENFtcMfopP
Ij9t6oQGRXEzcL47qV4rTkNGn2y9e4W3PKmxZvHZMpaiMad81aVViRuavHNSckte
uHQ3rOx3czFAF7m9Kb5uPqVh9LwSqe4BT+HJAimRRqzK32TNwKiT1xlkqJVHXHAQ
NRFuatkGT2MWYuj+EyQ8OfhouNssHVJ2Yv72egBmJvKbBMySSFMFUrH+mnprR3p9
QOvSpL/UyCHTrSIDh9mFusayUW8u9Z3YVY44BT8aUjLH78I6U8TXbUNVPgMzHu3A
b3MwoS1tiz73qMXsU2FwfM/FOjlb/D5I09bA2+kSzuvszwA6nilszG/tkCUJK9w2
uJp5HfxnMI8P1P1Xrc4JSDssHLrUBCyNhRs9WGuYImG/69jyk+Z2yMe7h5L29mge
btXZh92uxDDiXDy1agsHlYNZVH/j1DJzc+kYvLXCbVxMa+6gvlUh76xXQ+u/c0fi
YAJAZs4lytYs73qMogN8Nd0rC09huLlKzQnaRat+33wrbBeUYCgJgHjNIS3eYRFE
6g5e0UMmbsG7/xXwT0dVjYywycW5L1IoLlsnizwTXNSq0AFL6MNRfLhZo9CUoGMS
lSIIkYMBivylT91OWIwLQoqlYYPE+q8cfwGzWFc3ktaP1XaLZ139lPUn3/gJ83aN
dwgU5FeSo4idAM885MTw5CXf10NmrDEk6W1NWDbWWO/X4ic1IuzzpL6rkHMcWZ5B
c98SbkyCXVTUc9aAuCR9gefadgtu6yal+4MBfgN0yObYbpBx+XhpGbPwNB2f8a5k
jj/OxYUvR0fMfd9lIRl5Ato88p23KuiYEf2+f0QF9aARv81c27IKwjx8bFEaKBAr
/KgpNkHACTOnEcXd5zUy9O8kASNINCquQ9t0flKowAu1YCa354b4TJhwhNv3KU8z
k76I+jjIU4XWvdEqzOqfK8HKVIzDpQVTAGQodDQcxA1eC8lWiw8AwFC0GlSxBTNc
Saa+29UaJq0LRGALwDPZcDAHN88Xr38lS4/tjoF0EPLDEQ/RLWvwrWyj+aGKeku6
BWp+ueBSCRrz2+Y5lRNH1+enyNI7RoX7Aonn/VPkQ8/B8FyC2vMlVI2dkI7oc4FV
DDhJNTD/WO62o8VgOtyrTyLyiRJlti9Y236MGM7VgkTl/nQNF79YLluQAbQTqNsY
Hy/TsamUiJvz1NQyU1J0cq1DxQvFXJlnMlvt7as4jJy3ytevqNat+OoMv68Bk3no
hD8n3H5A8VFwG/jATRtpSAN5dW8obmIEd5kzUSJzOEIaorOZvMo8+xgbW2+/tOWV
GvoR4zLFspj0UFwc5Lfxgx63zNOUjSxm4tlL8286ix0Qag5RyQlU4rt+16BMXb6t
ec8HIsCnAGZnZpym8X08MY1dAG2BZIlScnaUnfmPYSeNPCPpI5RiCtgl6pxc/HT3
YlXf5aUnq40m6qavJinplSroo+bDojp5TIxB2SKE4oZLlai91htx9afj39pgE9eT
iKTrYGyw3ZY6EZ6RHTNSuhbGojJTFOyzm8wrOf1cAbzIO8s7NdCwsMqAJYpXtNuM
DT0QS9oE7QKlZG1v73tSNy1N1BLfKU7L4Z/sBLVTJuYJu871qZgAYML3H37ORyGr
hNc222BjAUzWTMmzwbjQlbE29SYj2UIWyP6EWOISE/gDnno3NO+y0UlxZfn31HVJ
RoylUTEx5YPh7fxplSsA9NHcxGqnpaAp/G4Apr02CH30Yjo0FN/8praX752bBjQ/
LUFW7I61/La51wiSeF7gE3W3i8NNv+Z16OeYHDFOyNXpRx4NLvEF1iwx0V5ZS/L2
DuxpNXUpggqxpMAdsbs9DBCsdlOkNXM34822DOkzWaDnvRGAf7B66ax2hHici11H
Mp+asXwqP/uWRp741i32UCYXy496BQbaoehiqvLdr4/UifTPf9DLmJIfI09xIbxH
gPIqFTrn7X3fhDs1Eye6K41htGMNqlcFBVlJvjufqhAHy2lV2FUKW+adfVnA8pvI
FutfzlsCskLoXseVXjPosRnHlD6mBXuSoZqqune8IfrTnkewcOmGm+JPnXCCvl9w
OxYBpeFWpYDLh4TdOmF5AytTMNvAGwYn0VKJ/9XE0Nld7/7wVH+w2tRTigiOuZJl
IvnzKva7iXwXjyBGfIYshDC4DdEu/QTAB1Sm34Xmxvac0owIABVQCFTMUFfnbZkH
B24pbOpfu5jeGR4jnZMSL3WKdEuRCrDtoGYNcDyxoLlv9yqBh9w7I1AM4gMSM3M1
HnSS5dR1coPDw6fyAQUbjirM1odGvjODFJEVAtfipT3iGVrUBrGmrkvoKqjx4ofj
g3yiNvZloKo+wTIMs8l47BpF8v5rLcS0KO33fxqfQ7lJNj/XFucm6M4ua6s5KnBI
CbolMavIyTuTB7bzgWw/SrsIuUDyUzzOL6/6/JC6+KKMV+/k78kLqX+BV0eT/bp7
d+PrpwSeXvRsGKMGyCuS1CwAwdfbjDFdFSVVtIQTcPToWwzT9nV5K3SQKBAHGWvq
KudPOXSH0ThfWQ3uwX+UL7a6A44c50IvgsjkGJNDYn7yvDjI2snttt/luiw6rgAz
dBL02Mcq8BG7kbPoQDd4seUurqQVWbaZTnLML6bY7Cu/2nSGULLds5uBwo7FY6yt
tUxivFjXfrgS7QxwikyZPV6Ndb59J03UptrMMq4sMmesGhfYFduSHCYcxqRYUkCr
qcDzwWRLe9SXnU9Rt4YWgV2mwWLjwggwZCPPqDd+ZHs+x/U/O5BEKOCi6Mez85Sh
WUUVlCGnECzqI9pcjLyV0ufnipgHDAnKa8+G2jexgFjeVS+pKsD9gpkFH1v1i6Ly
SfDHgFr6rjcIL0vaA14zh6UfiCRCMhGRXHu8QJOk7nZghjoeWdRQj3TYnilsiUGI
tuk6YQTQ/uMK/pQQL93kQsBz1O7W3a95WRqUe7dZDdQoS3RkSrPTTD1VMcq+TmH8
469VrEWCu7B/5SeHTeyBgGwLijYeL6oWVGJDe3YH+h7A1AX5vI9dLDKnl7Oqz8/i
rbOMEmmoJl77E5ya2R7GEIVix2Ijx1E0q6+PGFj2k28cLpIZwUOMU63SuQ1MatOd
qhk+qW8A+tCnTBgE2dbjgY3FZghOMQ5ISu3pInvRWHinOOlNTVUqjmsQpy0aQo2N
1C58sV0FCpdUypwl2O9fsTbonjcrhqxTY9d6AlwhTvtNS/O1KBDUjhxH6gFBBvkH
ROWKBAqltHOYQ/nrGnzoWsCtAoYH/cSWi6oMkUZCNZfc9qwwp+ZZMKGWKKNOd4/b
01d4JKh1O6RfLTNhhSGWSdNUmwzB6MomybQxZUimT/2bHK/dkHcxjvuyzux/thvy
LmEFUKWSMVaKH1vXSqcnSZbrrFEsXecSMojh9gj7GedDBYdMCifNcdTPadMl0Rt9
MBsj6kp2vWX5YyL4IF/chXrhu4+IRSV0Tlb+YY46GCdgJzBQJMe5Nn1P+9d64jrF
Q7Bka8eUofvdWZxWBzO79vXdcYt0Rm7GK0VcM6zTbpvSqaopFJ4e9DlBYHhENAsi
Z+7hAhACnd/tWkewWgyjXfOhc/nQBENoO/6xnIlk5r92V43ieeVrp/pAry7UkFuX
PDBuWdRYUdeU2iZDunEX+xqRaTy5+YrSZaEw+cp2R/Bxw1uRcVnAzAOBHq71Q9pp
kMGWqj8vKoPm35bYKk+MsiXmVcTIfEPt1usRjfvPKxSz0UW/CQUe55Hp5c9AEmsc
53wLObUJZgk9xK3wK+6lS5EnX/3XOXZI3hBdRCKV4EukAl01gjSj+xcAK7pC8Mml
+5rQDGX6qkMHdrMMQNS/vIJ3y2zhEysxg6DCuiQmjc5EYP/kAEsCOAYUhPTq2OVV
pxxjJRLohwhXnUgEsZEOmA/6gF4wtbV40KaseqFJhmaqEuu9emJF1X3BvxJb45Et
Dh/SttXoRfZ8tTmUHOV4SF+oSU9HDe/sJI+/Qrn6g9sHFrNxkZ6ymSzLGtpot6wB
7y/tcqsRAgs5p4XLpOcM5ObHsUN4iR1jtk9msp8/rrEJdtBdJFVMymp07zG7azij
bnaXLh1ZaKV07Alki+gZR2wzgHLtOgHJCFtEtSGoZ74v0J2+HYf0D4VUZzoa3o5T
WNeKnKhVhmpD+pi4Vxkjgy2KMtBAxk1eEUcntQcmaGUN3s6eUoGzUsOlDyhdb8M+
BDnrsNrq+GG0Dc7xM5ZtxaO5tqM4TOGttfQ/qO0pjHuRyxurQLvlA4Qil3YPWukm
tVH10qhbwqnJG164koz2AEAJ3PZYMEHNfaLzIKRjlTXrf9EUHC4hTcEt8T+4IVvD
NFH+wf5Ua4xURK2pnLte0u96COvqYG5F3eyDovslVNaSXL1s04lyeztq9iS4EQ5c
M7xYrprQ1cbaiwqc+7PXnoTfhj8JCVqDwBUv+vB0aPfXXbfizegjqUNYANhpuPOI
qbPhgA4sqelcT55B4fQt8qxb8hOqWHXLCohsG91r71C1OgHrPXCm/DzWRD69bddR
kZyxxLhEdjOM2ftav9Tv9s8aJnrOPF2nWUzTgEXNntyznYTvFMq83zPqvRzIyxOe
VctocZX91T/lAEmBdZhsFQy8wYnajXuohpnLSpo2MWXWInKEjSygDXgjFp1uAJ2B
8Uc4MfzR84w4W6cbjTqAY6nHwd8Vc+AKXaIRG5S7FGklpddq8Ea6WJrr+vJaVfRk
79QCZNQRdThpkTHBFV+je5GZP1L8x5ny+fIzM3tiLR7ivlJRPvBrHufq3Lags43S
V+ZVPk7Y1orTcAiEsysphKG4h8rX6o4HgkP5t1Qjs/b2KGEAKoePWNipEyDjBqPV
fbk5zaaUMmfMTQmcA5OPpRgAKnPFoXU8JGCNRCqHLBj72EM1L1cl549Dz6EaW5L1
EIlycw9mPGQqiA+fXtmb3rKAtaLqEZ08nFrkuaqPhiX5H67869RYSr3wb9rMiUfx
D2hAQlSEQv24ugzIxqqtY7gxy5uSiFjfUEWmeWrZG/1ZQoJiClHv+jldKkrc9LFc
VF9rvlNKI9Jc9T4x/NxWNGkbMUfKbsRGg5E/AsfbzIeMv1YOgU/igrWkrZ4ddRYT
zE4J1BnsclU/vcsuv9/AUmda2sclldptCsjCx3UGd/Gm/yK1CU6mES0CX75SK1VB
aQC3c7WPiCgRUvudG35cToWvsH79eJS+rUgg57MXXDH6bUdiyeZxdned/i/4QxOF
TYT8c+cL38kG5otEr7wUaPqvoHDb8xXzH5W8wuhgRSzBkLNbGouF2ZVilP0+9liQ
xVK6vUc5oNGJu8kF8Kr6fvOpvHbe7l+mi76fNp94dbHW9GSLJIYXyE9vNbXCTOqG
tSqoJutwPFwtM/rMTNl9eN+yFtC+anH0tnV+m1lD1rRY1H8+TDiAUfKEPGEet+mP
6bIMkYp3vJWkoIDECQYZyXGIu96vrivtjDvphNJJbo3tGP1D0hU9LoT7vlQtRAk1
UQUdAsxeSNV5Z/K6f4N0E5SPo+4jGaKIP6S5gujl/I/DUlIS/XTnmOGTUy0Is3Ff
Za8EHuYUP7stP2z7eY3oqaujTobAmN7/ipSJadwa4pQEOYxaTxqjywuML4ASrQI9
4d8dinhKWEqXZWLw2QBql8lHBMDPPtrG9ZOdXZigk3Q8YWnrh2OijADx4GuUQFFf
VEYTZeVWJB3Nc5r4Vg0BDOQF+r1CR6J01ElzrGolInb/x0BrGTd+zYMVa9OT+Rdj
DTB3XL8SXqoHXGt1g1h5L4ZMu7hf+/mliy5xPCpmXGB945jKkluBkdARInl5SO0X
SZwYHElkKJiZEAiLLkP42QkZ/uD/x4+bCIr1cfdZ3W2OK31OBd69paz80U69VsM2
kauEW+Sbyl2A+j3zeIJ72CBZPgGyErRtSdXjZq058O2kJ9Klj9TngKtCZjPcSNYo
g+gJS/1PqRdysqmeYVLi6NW+X/I2axzSLnlSGPN+tWZslO3s38/laXCvHgBQPEX5
Ja4b3NtY4BOd8bix+Bgr0+1AzuBlYQGGhA0hEOcZPyN8Cq69B5rT6MWiQIe1eN4x
z3luOeMFJNj7IbYpO3ujGpyhyLV08rXvpALK3+WtnoQ7YhihrFD/1BnvIZSRyGL7
QQYCG0RggDTeL18tm28lN+XbADmRPFrJni51kWh7MWUTg8hgZTqwBG80zFHT0rj4
d1nrlzqcNGt5gsz8+5IXn9I9MVp7Roz0J7ry5FtOo0oVAe6iuBW+//teV5T71EEJ
E5VceOapIjW9ocgLCa1LPgZ1Pypt/TZqqWzBwiJqFjs8p/UW0VAWpJGk/QWuzLHf
czMRlgBfqczi8jum1maPKXIDw5A0dFHroJH1OLXGfpADS7j7M2L0QrM5O6JhXoZ8
SDI43BOhztpPxV+EnJeJk0SywHSKHvFfrkwRlQPIlf+O/X9IjVdFzndl1yWnhuxQ
YS6zQV8JbWkPxEUaNBhTfWMnyQhzJECC5PXwXHeWlfTxcigtjxpOjaNuSeuziVds
sO3KZlVRRMw/9QPxghsJ9DUpes6bxr6e2I1T26XcAj7QLq+dOr0qThHGB9m6cVqi
LlFIUuF6jch4RmzECjQU0a+z/onYfp5IczKsrei0WhloV42VDQ1cIg+CxAH9ddky
WTXMRwd4shfZe4vOzBx+v0EE5U4Jl+EkBXrbea7qhWeem33ECmaSr/uguaBBpF3l
bldV6WMpk/uIvCXS+dyXj4UNvfADzbl0RjeMx+3XJ4dY3MhLXeonJvlAI2OTaTD4
3ao+8fgivp6uXOU8uzq0xzwVWB0KoTarENXQAE/sZLenOT5ddnN0jrREOB8G7abN
G+LQCnh6kj5n8cW4xPpsGmrpZKiyfbVqLCbG/l7LKqeqnmJXxJC7lv1tRTzZ+86R
hPXlxJCjQwOGWY0VmHnIgiRzQHjTc6YrpYW8bro6PK/PQe2NyigGD3gRRouFlF8/
qAebV/2vCoAD7BR3m2FjCi/+oQLhhz2h3DnMUk/BjDOHdcfSo4tskp4uHtba83WT
N4Ni0wE+ZSSZOzdBCmo1e2ODP6Cwl2gIxloKF8QI8oPgSjPkG/7oTNGF9iiOkTtB
uOum9w9WZmzhTm5EAEuk3CzGAgd4Vb4gq/8BFWvfk9a7j3RheXvra1oMGPySX6oI
lwXPv5fmkHI5+n57S3JuYs6EdySArqCV6TdcUBYw7aD4gzzIxpkjE+iemysZvnSY
/ht4+ddvdmG5Jf3imqfDSRgaGk/Zsap45Nd032ae5NMa2a7/SoE5cqcvEqxWgxHh
Ag/yjVenjbvZZDjI19Ko3FzSu6DSl6n8CgiYCcaafl8iOrAX314jcrdQVKkEq9EZ
b64RYgLx4jGIeVz2roYOd84YVPktmCS/aHtyV9MONWQjTWuHko/pXobMB8wxxsSt
/NQAam60Th0xeX1WoRKPzz1dNAMuOzO5yNdsQHP0Ym5wNEWGVdFtrUl+g7Lw/WKS
wtITkZ5tIefgdce51dZm/CO0vpYR1irt8UGBZ0gXv3j5ChOKTjDHUGBFSwk84zoD
Anea0rKVMEaVpsgKLvlPyJADBU9hCzoVH9+1ez4N6770sYAX8ukM5EsJFXu3aMxu
kCndgzA/dj05rJ9sS7KIzbFmSLN8EgoXRKGOhtySvdE49X15ulbXPohJdqKbOXKh
62vbTsFxKkkC3jHzYVx6GOc8scYxSkl4X/8X7sXOj6fqiVARpXw8tb/BipNAkECy
apEZoLE8Esl3mOuKBN4SqkkEeb/hQWKpLRzWkn/+Fa/JYqcXKuuXjMVBYXWBoAEs
4DfdWs/L630qGQJOXFMuSjGlCM4nEbtF8O3qPmnpKytMm9d5v18ySeB1k77/tA13
gHURZt397C6INRhtMbIpvNdeCm0D6gbWj9+g+IBpdLp7Z05GAUN1wTTwzbi+RxtL
GF7wA735Q9uIt0gZ4pFb+2FjyQWyuSg6fFKZVC8Z5fAFeaZO5+JlkCNU3Uh2u4wc
ROiEpPL9fnyShUJSCmQFvFCF4KRzDFOgFJHupEfHVo9TDWCOFn7IK1I+bwhj2oe8
dem9uuDwjiV2XzhUrOV+OgUWzcSMkPKXWtvOnq37JKPZFrm0K86tzOzbwTHk7gAy
yAticsJzeASELPCjZ7nwNQ1v3ExpSWcet4wynG6yHdVuKN80Ije1C/Lf8JeUYXYc
KEgfXpGwdZjFCvv52Mv6PSAfJJNhJENxhVZCCi8QUCJfQJ/fqFZyY9eg1aAbdKoW
PnWIwjJi2g6ohAZqFF1d1DCAUw8bMtKy925FQym2v+UWfGAMSKI3tLJKO9Vpj44y
4KjwyA8+xMxja9wKk3irplkbE69Ct42sIOwkEnS24VBQKVQq+RfER5lbkf1HSm7q
5wwKpPndpywLysinX3w4wdHs0hAVdxKNpDk40XFuIYzT0Bk3N8eyOk5y8UOm0YSH
bT/mV9p5/gCz86uYpUCcDz567i7yQS7XhjR4MVs/wCnq5HMw4mkGEAF27cFxlNco
wUr7cMiJxdhcBfmMCfx8nVr497dwt2+snBTwk/qAbpybUrD0KF4XwViHHlQfEGBj
hQT4PBN7h0MTULOk5xOdMT6FP5WP99JdWS7v9LPpy0JVtkkqduo8+5LOHlftBUEL
oWGt69HYEKmDob647b87c0lmGFksCP069t9HnkVqOvgPfIp/N2ZWQqPoyvwy1NT8
7zibCwbqNWyzlxRX0qLeY/TPoMjwJ7IJHNR1GvxYV3lckyDP135JrI6utuONbcEl
ki3/IG3cWTGLZZqc208qiH2JirXsWXuB4HWmrJBF9jPCoGJXEaeYcOWWcTA5lMLy
yWBZQh/q/1aEThhN+Kk0mb26N4S9UkrenB2QA38eo2dL0AmknxcE5D1ZJjjPrhn4
RWuvZIJW0x/i8q/f4/e+aHysLn+qTLG9Sig8/IcEoR6FMmppKxS/OTqea4aVDifI
lS0ETAk5NHlwjepfQFzxcaDtbCX1xFli3kgIjWJa06rSXGUOw1axSYNGSOxX+jJQ
FRQGOOR2RSMKJZm85bi6ITmMJnlShwspyY/XIA4e2oSiRtgqiYBSsfDrXNiA1+3C
SvkuCORt3kgRRxujq7JbXCAV9p/2J26Mk54+i0eOd0roYZH7mf9TsQFrkwzeOJ8g
XwySIxUQtvAUpdz8SBzUFlwRzufLoz9T1uQgIPasZ1oxXXACqFhgcEZ6xTJBd3CG
LzT211eqgyddj8WMKNh6EqjfNLGsBtshDfVNwRTOB5bpZO1CyopAWHaU7M4R2yFW
25g3aLIvZZkEeZRFyUdr8Hp2AItle2fw0BB07T47yIRa+WVjoN9p1Xl0GxRV/Yn8
+ynxyrK9GPR3YFcL5HqYtp4a+KIkPqlfsEg73aem5BFJprKlGcbJqoJWD5pAnv0m
mnMDpONvH5LcH9KQgXvwpvVKQfEnltoaVChgt6o6KagkPGUumwm0Op3GlW7+xY9a
CsapRDuwZZcXY7HZOGjIwCSy8t9oYU7UkeeyiOyJD52tON577GDHJIuWwPrJpFnG
AzzK/AAFI+qgTRXOEr3bq+jJCMM+HQAvBKYZfugjD6dkjUptSeFHs3bvlF7WGyc4
vbDIVzV6VSZzAiZIfYCnAYVaxVMGjMA0/VqtKr5xOy90je6GxTF3i7DZHIHZmqiE
3RVDZ4tFFYFABt+cpE1prEImBUc034LP7Syr9ZdocGdEvqVpXM+PrDG9mXv087an
nnYCxYqf/V8WW645dRRs+6xKkXuVGrILven+TS0ALKnr3XzsnGHhK5FDCK33/6cZ
ssg7/NTbqpFlhqi0QwYGd7CmigIr3wPn27rCKO79zzs+L5igcFAA9PvR4wdqbwRM
++zhKrGNHQQASTy65D7+z+lzfw/8cOFt74Jqj/T7ETvLzsUQbmn4ts+Y5fY4XlW/
4UdWkJ8ra7BxlSaTvPkOVtJiYbLqAC7ej0AMh64jKfZv48yNL1rQEGTJGUsYoe89
8cmY60SZR8RTVpYCBchrzMjNMx9i3s/SdLgcN1VPTHuiuEBLxsnPK2EaUC1tMC32
14nyPk18x/7zChD2+XNdBUzkW64TQXQ2bNMGs26XinIihm78eim/S0xuiVfEpHkX
0FhLdQ6Ac5/QQgBT2eDKkx/Emll+3i0JJZBA5f8hRXCftnbjVk6qcqpz86nKlYRa
3N3pTS9Nw7bvjhV7qKDUIfqIvIXrv4UvlpXmkzbtg9aWvmJmiBKVuJlkzD+uwC8R
kPDUepSGa6+krfnzTlKWy1CqrMSIJnF2iAwKsVIzQxzfTs9wgWZSvYzSlX271hhE
YpalBz484yRntixqjYXno+f3RtZdGTmSxM1U91foykzGlEwlrLmiCJwvhUVq5J9P
GXcxxOmtQop3ZrGyEK+xhh+W6VxTLqd5yIL91yG5hWrkEHdc9PSJyQ9zig+RA+yK
nYLEo3ly8YtyMS1ys+fUQOWhYu2DwxoLcHfrSJKxWcvcRUC0ddg2gIeqxG2HTnet
VVvCT/3fRqjuE712ThQaiJ4lO+1lgY65N1hivZWRA0d0wtZ6t0F56dkMjrobwd6r
7NoRFV/ZkQMEFJ5RxgcDLLhsDpAaM10SRbamGE9WG3anHoT6f/qiEo5KntkexLo+
n19Ig3cXXxRTB+p7VdILBom4iKT5eewORalrZDYE6IBkLcGhs3/lqFo/9Xx2Feew
LzbAZ7m/0glh1HkqXJGc6cgVP9RJB64j8ZvOwNSucjflARQD5zQHTftMF+VcCSI9
P/G09bIWV/S2+BdJ2ExcdBLJmPHpeXNADlfYgBJ4k4VG7iehEWkJFhfPdFbqXWy3
LH8QbC9mlQk+FhJ1gyNdfEoJTur74D51BGGv/q1J5vlt/uCxAjjj+TBG4S1wbUtS
ZGh8z/FFdKmyfYwrxVL3sK4uYROlhtEj46UaUTq3W/2IV1glB2LyX2nCpbq0KRGD
pKK3DE51EdGt9iML15P6NBNYpfU14y3epwMVUFWpPH2uTfU3MdDzhvNWRxxHLx3n
KU4BdfFHtOc5YCCMq7DlP9FYp8b0A9Qr6vkiOO2PZRgqiTTd7jAK3NLcpnvEh7Wm
3lXYkDkcGPNYu+sPSQBGTz2Adlhf8K/sJqAtNyV0hFZlIxlu2fPFmNwi7Ihe/i6Q
HmSc2pE3E3lsheKU4hZbFcJBu96Gjx165KghnGZFnG6q9F99FTIviH9jontZsT/W
HUHHj2AahIi74TKcYqrTOmeLS4dB4LZwuANCR6IiBHeli0uafjyKVIo9mOnCuTr6
HSU0xJNnOPjDmqUcVzWcCt3nqL9C6aj12CRybJpvRBMeUUnXrSz3/zqN+vO5H3eS
YbwgUWTaT9xsTkrMDI26JMXOc0RptE+4u6QgvP4Im1yBW2++h+FvBR9C5eLaTDL4
2Y3qeG20KdYr/Dzt09UkqlpiDW7g6gA3fSOoEUAUNnzec6RiGaEuHYkyEgHoksRy
IFnIwz5yNv/g/CseE5VYiLdeJVcAW91qqo50aeuDbz0P/0sDT6fR+RZybPqax/LD
vRGHTA+KztlMq96m8VlRNuKx+ed5e8gl3jwFo9zZTIeerhp++WzQqpf55efrOJLd
NlplMa+66n45PfeV2w4tpo0Cg7/gfDQXqPcwZTmUxRnQA6JP8zDGa853tdyfPXhY
JcgfEJLjUzwYGGWMMww/7p9uGM9VHEzIj8nd8qcA8cY8YKwXIuvAoUSP+Fph7FYi
ByFrn6eHv9b12p8D48bIib3vm8RWAO1Vu2p5xyfIxKW/VLy33l+yAewjL6GCv2PU
F7JN2OzANB4MdUh9C1xV+vf8DRB7bWz5bKaKsFG6/41cN+6Uiv+gkjDFdwqWtkxu
YjlxEAkgrW2rEMoYBzVvCX5bhZZAgGX7i3bm6CO9Igzsp88vT4SbALDg4BoeHYTz
SfBjkeQl41SpbWrlsEua6HJI3VdsT4V+Bgo9FSR8qM/fb9A5Ibiv3TTVv1DC4+01
vs4U9XAGGUXfmR6fIHzXJyDqrHHZtFtuQ2i9P79jiMdZx8FIejMQtNf+RAeUKk0R
BDNNvI/YN/eqWLo6Pwh6v/mZC3kpVCaAkpa73cD+HgLPxARudB5hQySSLoEUo5+h
N7Mp9IgTiaZWPbupr93EZ54wnBzee72BG0cIy4s+RZmjRjTXNUL6ucvBugnnp+L2
A78T6o/LjQ+zl9YncmpPhUManLVYZeR86coWMpq3j2bGk/Yhj/yvAx0RhjtDGQJw
8isCY2IrOaTjapye5sUWUPnEKrRLcWj+5Ywf5UhKsrc0CGeqV+8Lzw5Se67vX2nB
qkiEW16Xj22kjhoxzPLfQWNtfN3IHLNmCnhoT6S+3Vxa57avD+uG18ba8p6oJS46
CCMetmc9XKkL7YHsmPOgdKn0tenMJTojqAvRsUG12OfuK7PAKqji878NBVen828E
S+bJQfsDLOA0Hy8OWp3IqcOeYybDcuVaa+o6e56FEhU06qsOSoSwry4SI929DpeS
XYjSbKEjgyH7BD4j2vXLeEv2lFyie9NS/9EEIvgKTzK1KLf5me+QQoSGEfRQ9qcy
HGFacjr/0ro52l6a/Oay2SSG7rP51ogetLOlFPS5ENicS5Kp0OKXdKgBpvCk8/pq
xUJJzhNDwUgcRo5jXnOIo8Ul61asTXRSFfn/59VgrhVKN3fZYHUXeJNfewNZhnMp
pSg/8rezatxSpns2atrOIdzbhIfN4M+K1y/mypiUH8Q/7tqwISxcFWo/g7ldYgA7
1uTgc2J0+/V4ZjJZTRqFtAVKsTCGGrt0aQO8D8zgvsuRm+cnoUtFLR/g3gHCuzYk
H1r/PVsBS56xaUcRj6VvBvf0XkHphTdm9qWQFtRv5lrBdicb9yufbmTMdZv7Dgjt
yM/kN9P82kmnb/+aGdgMegZ/H25JbplT6fIZRCaLmjZYevflvxWyX/cKv5DQO2jO
NngqeQdrjZ5o+3fZUcQMjFQjpcRvALqRPh7z8wSw5eBs5D7Jn2uePJDjLI/SAj5u
tfZSuJ1FJIy4N7Yr4hig05ahdYOqgORslAviPhZDvkEa4BO7b9luXHxOy4kXsGxI
sam0OLF9Ifo5UnS8avlg6Dcb77N0zQvj8dMW/HV041gT3TFS2TeuXTRbiDNVVemI
C0iWeJYRafATA5AUZgHH1tnuDg/ZPzNri/wp20tQEmhi8VC0Gnu5+IVyXbSPgVa8
06Q+lhjE67bpPCBLJdUO3nW9WfiHnM4mZLQMXA6zG+2wPlakYP8QlBY2QhxUD25W
PN+ZDz4cUs4BbJdSZdgW7yc4KgFpcXAnaZ/Qc/ppln/+Bwo2dNhFxgocx/VNnKb0
lns2R45SAC72ACtmUX5xgiYjt6nbzGIWrKs0hjch1mv2VOy5Eqxx6+moGYmlwazn
pxsn9gwDdL4MW1wlHp+WBc3ivuw8R1HmHHFrO4gxV8ZaVWcVyUZdoHkkM4sHs5/G
dIaluMdqBo473Ot47LdTtEHjUAKC5SxKPv2rKX+NMOvLcCfDxZ6hr4cj/hpx2ygz
O61CWMtxlqq32uKHvqD0BVypEKQRgV6pw5xmwOSUjVJ1XzG9BeLWmhmjF/wCguL5
mXFD5Kr2UJLwjVE83LCGu4XEGp4PrzGNT2lJQGgzt/kbdYUBizx9p7+e/tDBMik1
quOHVTLxuAAfjuSkdeBxekXQiukcnQIQ308SXM+imdfBzjgHJB1wci6FLTWTsEWa
Pw1mhVbuUI7m4lKLeVs6rODgfSaLx8JZ0cm4qtFBLYGRMZfpEWblpXEW77iPYefa
t4ZRtbStPVpvX73YlP3QDNO08Zvm69PQpRwS19gZWxpjfWdlTsz6SgM75rGcAfSk
pap4StLavuuL0Esc3it6P3NHrwD/Mb4y0RReY73bUM1hjY7QFGt82shxz+Ioaese
woXRh1ltmy3cTLbb2E3ehmmn5PzN/vj1oH7bLuEqbkEAS/ZyqsQoH7reLhQdcgc1
FHht8s9Ufj47RWDHa7e0s/ktciDL9Ulg/afO+Ey/Q970WMkSFEeQvpyTKK2/8XPP
X6Dh5Akka65DPwIAZoePWAEHlquhq40RZ85ptZFDZ6Zri/spoqq2jMZow2UtPXzE
6foBjPl+1n0nBjebcUZf6sQS5LpRxPJ8QUa9fB8RUIzj9InkhOAt5KAhluKZRpsK
KMWZ9vD+788AJUv3HxI8EAyk2h+Vs/ySQkTeD3+MbQW9NtmcWSD2tpdDDFJWAY71
eskF/1DJSOycxXMJmx1zxGJNuho35SBoiPaKyBx5crPGaR83r6fFIdoh+m601eX5
KWTpmej5tgwS529H9dbbpePmxM1/XH3Lf2PeHC2PhOn/NSLZtqoExc5WtG1LcBOl
jwEDJz6yquVQDZuSZeXDJY3JWjHSHdp6cZ1t9/fPj5f2YbQpBx98fsQtOOvdM2LT
JvHVEeMdGW+CLmYpImhL4qN4colekqv/pXAVOXPbKh1OWwYiAda9bRLJfCzFovYs
SL4QlOGxwezuBP5bF/XkkZKZo6+dnpXZQUjS4qXpy7lq7JXgi8NDcrOCbXCFM+V1
5jqQ3jM4HZyj+90UM5c8nIRGNz0lcW6or061RWj+NANqCPHCHWGlb+ADupKZX712
Ml/B4PAgcppd+RzwxtNeqAr1Eyw0SBJCpFFDGFxGXjBWichhG7iHOvHbs2QSb9kH
8uvESiMQBTviCDJfCmuAjgkDPf9FzTMuCoio5QRePMSaKZXPfhqc9LSxf7NGOwdK
E83CH9JkbcfmiddFdpIGBdKlMqlrzurOpX+SyeD4xIW/Nmbn+6h+8JcJSNFlaB5+
SF6X5OaRklVBOAtoR2wtQKOgDRD3B/d0cmu+/LGj8mC0FLEqaWKWv9+4L+QLVytq
5aTdLA1/5Y52uNVC4UvpC2DvzqGUIlczzsXryVptoLUY6KTMeCbQY5hJrkjyVX0L
2cGA2IhF/a5KxPjWrb4WLUROh0QDr+ocdRydMy+6Ag0zPoUayJT+Z9dwKZsutqJx
qU0Z04kJr6IpuQofMu5jc1fupJwCF2MqKHeuPtsDtPs7ZNbzwq6jTXtTpcAtuZFq
XSm6WZhAZOOLJO2aIl2rfH0NQdRitoFGxlZu4tGi8L5uS2/4i1OAN9QigFlDzwcG
sKKQCqWyeTuLEVCKVyJ9m6d6wlrHYNxZHG1qXaLGtn5+ITG7glZWdW691Fc2ebpY
3+5UU3vXBizj9xYyGXrEq4/sdqSsQzJz7iI4eQatYUTxAtzRhW4yUjfp+wPE5sgP
pfxpYpLdlKZAVlZYtJIQ/1w6NTb5lo+seCgf2LPiRJipi09SaTo6c2W5REPmglb6
HjwEbgzYtBlL3mvJdzHZTEjKwHg31gSG08fIHjgcGvrTQMd0slkh7FfXXRNKNogu
mI/5n09P8zL2nqK5Q9wzYQdVPVLqQ5l7Nur05ygTbVHBsGVji9v8D5LOwoltDs8D
wAERF7xkbZsAI/AgO9xx4G0Tt1MrTYNFKOF8KDf/gKlQNIRhW1BzVmU3igOPxPBb
v4AAjDbJvFIb+9/ykAO7uv7zTT1rnLEM0nPTs3Ep9D+K3J3rSynEv2cwbdpDz9kA
flClfFaKtp9xBiGMbpU/Sg+nfm6iyzXGbNS9uFe2Js+Y/hmWR/VzTypCpHsbwXXe
48wetUwPH4vs/jzkGw/237MOTKt/q7bpzfV13VSJwpen6YrG/HBq4mM9Uii7gt6w
Se5XIBz4C7DZfoMoARmEld2KwCND+pCOVhyTToPtZXWQ+e8k8sFlC587ANr9mIxl
KDp7xGlGrCv36MY0aGQLMB3HdSwp3maVpuEW7sjp8p1wtrfsX+VGTP2DKgI9g+Hc
GwwJg7e43ts/g3AFcPkWjqjzDDhstRteITLd6MKDQxV5gDbCsaduBfcS6cE0vVbp
SCYR/uy0VlvOC0xKD0AGGLt0wKrFRsnUcA2ioCCwR1LMHAwn1ZMcJbrFZU72iZrV
5In6O9qYTbYWFbWW34GGR89EzdlYGjMbcEGq947b9eGbDcfm4QMXhRUmYHnL6ky/
v5pfG1xVNvLrMqy4SLBKmm4+qUqX0Vzr7qgm3i5/uq6Y33eJsfzxrwKpLyvzNODA
MA6o30VrRv4zuJ6VETAfDaxvs8uKGaRyw5Mrt+dbpd/SqFPyw0qduWtRtht6q5XB
65BfZlOJyfMzMm52IdUQLgHZtV1b2fr796cmG1g7Gjf3qNU4C2eEDn1AvRMhl8kM
oPOoD6l6XJ5xTL8qt25WMat9mC7r2PlDQzopjuN4LQzXu09h8ca8HzRjELuYz4lK
0WtRb6wigJR6V9dpVb2gnV5Sf4s8qrkue1hDoxa7ZZ0lqI7mGX+WybOMiYorXZ2a
9DPNVxcsZXicls30IlBC9dtK7PPGiV6MZrMfmvNBqDeKFv3Y0LMwlVdSmQ94HjwY
maSm0QjnqeVlyEVEbC5Vubw5OSpTfOS+fWcDiK93X9rXjKMymrW5BrAMtNCyT9PO
1T/r8e+FGEkjqC7O092FdUchlWs+ulplpGk9Ljr6OSSg/+9ZkuNsES5JfQOkhG/9
WbvvlGFHH1649jQ4M0Kml4x90Jw0iELGq+K9DHAw2lrO3BYdZZ34XlVAvJbDerQM
+YimiZv4KRBBb/EyJ/ihPbwDsAg0oKNCb//t34m+bsvYB76hFKhdqyiXeCYI4Ou8
/RoY6AT8jBvV507NsFokpfoRVOevuBKNjDLVOYS2YC37vwKx7r1gsHFwKOpXN11t
zEXM4+IUzN8SylR666k/x17WZ+bunnkL4RuibHZZMBZ+JMnxF+d4ZzgnH3sEPiT7
nbv/zViBNDf5SXYBM3JhdZ1I/Z/2ww9lrvYVpSYGZD+bI4v5pULFHDwop28YmKLn
cJfGcR341iI+H4LRAe00PUiW0+fgB7YGFVg1chPIIGFdNUiESiOih5XCtngtnIPt
KXa+6wkav1Nnz+OIAsB6pHp6f8u0h3p6nezvB94QU9cBKOsJN/7pcApChOr8zS2D
ZmRUGwcPqoQURDj4acrC8PAYciTAvjYGeK9tfdyilPuKGcyIHhMJtwQxQq/DnOvd
WxLPLUVOlWdUDINV2RIVNMkWTRjAji9ixXerCXaC1a/qdRRE9NX3ae12GMRmuuxQ
h2WwzxmMjCu5QUkv0ljTEaLdc3isDCAzH6U5cs71suqUyGEKSWRRMO05dPsQ1EsA
YeIVl5wKOqsCRfpQpMcqFvKQBRSfFVxN5sKJsKj5EmcXyMim4EdVwvOHyYul5a9p
dD/Eqye2FYb5GshDEpoi7vyWZ8I6NeZ1XCanl9ad/FzxjWI7CPmXxUCw/hTfjke9
zcCIihF3Ny4ZTpXnnXoEo6mk4eyabG2SAKruoM3TQHgaXhGiOw0kg265rJz5giOy
F3os4SkcAsAtFXKdpGkLwEJNKXRo+/bfTsx9rIj0S7iRL6nWjYdh7ZUh0LPJVyaQ
foQ7ipAl3jFHEZw3nldcF1ssgwQewr8JqvNnPC12thwzZcs3lgH+ghAsZ0VPJeXc
keZn0NfXoDnd7Fe9cDlg7aCBK5ywvrIw7Pcn29/Q+7g3tXVXF13Asl/iMCBjxwE7
oQB9HED1ND+1W2PSxt891M+T1bnFKgFFeqGDMiJu+rDR3X+WPHXAxe07jCxgldz1
Kj/rVlnb0PGteUXjLNob6N4WfnBSs31Xs0WCZYvGV/YD6zWm95nbbGbQ+KgLx+9D
wW47tMkoyII0TKYfzV9cir3j+P6IonTuBRPFgwrltN3qLnIAO3zOTVAOJuXalwXM
yzIBL5q8I/ipHFevaF7GxPxOaSfxfTTxGqgdJQm/E4+TEgzWPspvAXrbH/qGQ15E
eYNnfJDhWun50RiSHDS18N2Uknjrg8f6kpi29SMQifyq4RkhOSCG7t2LUGmCiYBp
79PYxxC8rBhwJ1x69/8aVQ3bWdi7s1FxuibWrjtm1ugawIBk/g57Z3up60rdPd1j
Vt7pmv2oGnafvqusA7GTJq1P/1ocypPicUGN7+desnIawNsX3f3kYzq6369r2Lbx
vq3TjGQ339cX5lbAsml3u1gIERsX9sFsEoUhu/HWewKG68r0Ljnvj6gq42e69YdD
XtVauC1iqauQub+ddEofjp4gRJNdsllt1KeZxFS/NYOoj9tVwwL+uZAOrWNc8ZVx
2ApN5+5PGYq2Mul9OT7Pa1/Opd5IS8QtpFnLboR4DuABFblj2VhaLZD8KXppTbYw
5XL0xGlAwbcWxqyFuYL4xFClXFP89KtlYojodM2s12VMBmmTjiS/hhBkDEAa0JMh
G7r3tV3KVGKRMYb+eKN4CD/TcvzAO8ZCR5DzxrZZqr5KumK5r3Xo9623XQFS3wsD
0XZeoMxYQEOWa3u1UgXEuDw2rAW2RFUFJTUg0q9RudmCPClvsr9bhs6XA0mnepcP
qI627zVVWr0ymIKan+i0xrcPhPxbpLHDWR8hYjpeNSNeqm57By7+tukYvcoe/u9Q
L8w7m0gkWlPobOrEn9a5FZ1mtERUIX9zmFv9ss2vQrUZwjK4aPjlLXZgf4LLcn/F
cRr/remU1hVoJqI94fiFatH5zyZ36DZ9SdAFcqwul3YYNXnPDY6BeEELRgkkA6k4
nSSC/coQS7wLm2h7UO25knCwkHOYN5d0roUU+4HMH6ijjKNlDVbK1BmDOB+Wa/N4
3R4jeYaIGxzYc09j2rDstUTT9MKYoKt/uU9/4scvrv9IDk8NfiN/EntHcILhw4FS
TM+nkcasPPnEQY2+JXl9GVfyQiGtv/Mj29jf8tiOb9RIIxu57Lsv3D4YBhmwbGIk
Q1lpwaJ094T7dUVTClATRMDxAPxV9lKP+aBwyyJijB+T53LTgRtxudrS6enwd2DE
yTR+/mJiigDpRfp0n0C2NJ29Nk+XhnavV3irFubIFAoO/VHtmy6ZbfvTpcGHuCF/
YjdVJG5YQoFmuv/Gr0NtDOgR45YqQIk3Cc1tG/9ymk9L6LcHpD8ffR7V5NMTNwi0
XpdQhti1Q1H9+rybPuKVxSiI99kZ6oJDrmxkEnkvWhJ21tU1lO8BWph2QmDKsQeF
n/D9IUY1U4LmZnwv/gqCKLDsJsZQMCEw7IZmwoRv4BBLo8Wn3WPckiQF0cMNiQc+
s04PJIdbEgArfw56DQUDe7xF52BowuxepYrIAohVwriX8kyESGFSu/s4lOXf79z6
cJ1lDitOaU7aol9tZSjyGZtML9Njo7/s7srAv5oIn3eRYbxb1+7qGl3QIQTQerQB
Yj5tb7Cgb4/tOvzWCiPGFDSCZ47jtPlFOP8YTHuJrPTdQ6XmxFKSDytLGfDGVyYM
wciEFEOCBmbdCY9xzAOjAid+GMaheb9anEBgevbGYh6yxPu9Lm2TA1Nb0WqjagbN
4LIZWcJQJOGfhWSWs0kNLFNIZntne14LxJrfrhyzxt0tposqKsqwmds8lKtmQkF4
o9TuxxwJUC8hW2RwG7JYicx3xNv+X+gSM6vVZ16jrqJUJVN1HZc82fC+YS6HS2cX
YdVCiNZtW5CzYt/+n/gGar/xnPbxhKvneVRrJ/dApflbLS7TXHdX1fRLb7hxKUvx
D0pHa/MeEcVlP94vEYKbz6cQlTtj7XAXYYtiYUH/1x7CHR8/SP42jhTSzsicufaI
OqYZGwZum0jMF4j+HYd5FMkFOlsu+Wg3OEO/gBG7IuNaxQFzeK4OCmFaQJ8UESBQ
paMPG7pVJhMTsQ6ybUoaYUVdGhZrvCNRjulGw3wIE+TjqhjEoTO6dXvj+BlXtguK
i3q9QrqVdkMtzRTMspQvWTvSWrCJoOLaSxVHba94JnBlhCKpNMIsNuZ7+uSw3sUM
rlxySyOHY5mK7jKtn0zmhQaci76kQCezJDwE1yePI793eGKQUOR0qsHDH3P5xnbK
vfC6RHP+2h7ie5rafI+3UH6SWIimUpwW+mu4z/xLCjDvbzcdMumJqnPkkq4l5UAy
DgJAV2xRSvAaD9OfLmfExiAP9JbhLPjBwHbMkbzatV55vEAKxgO59wYOsCEvtVqj
oOEph+QHpyI0MWt6GTD7kgB3s8StfqRzArxVi6sIoDEFaIsB+cMddUvogEbBj/nc
TUFdbKCkKp2oDN/8el/P/U47FOPxQ1+krKGlGaFul+DvLN/Ef1ZkBOqilOCF3jXd
3L7EyQurzgan2S59qXJlqi5TcAxDJKZsTGt8EAFN/g23NcbilyOHNV8XXQC/1SQH
oHtxJ4uIA43+ortprnT+80tge66a+TbbOM0KIzIu+HLjSDTtgxY+mSTi3228or2X
IHnFY9/ouf1dwtL4C7Sqzr9MMj+7WOriL9MIZxeSSFSKmGCzYg5pc0KtKsIhQOt4
IY0UMJPLYU2Bcg/Vzad887FBuvVlgxB0Xs2VKyDlwRovyv4Stjkmwj4iMDibbU94
2FVyv9okJBuNxMa2cJ0LTdZgt0DfjdscJnAbBeu/cfTqFdCODZwUZ0rrSORZ3iiU
XAJDP7qvKWrc+LZ0dHNt5GVqI8fQbdTnx/0TrVfyDv9M2oAsIr2TbdBXzIvxjMFN
whmDNpqkEsDrNV13g1FhimquLz9D+jSg+SuuY75IjrgDLveSf6flSyXedV+DwObt
yIkODcE5v64JmKhY41B8vKFIq26pP6QfDYvux6oF3KvZ14aMWDTRoU0wf4yxLtk5
GN5kr1/tXD517/keeyHb8suMP+T7FV0aN9ZewPwbgefawIPTVgJzoBPB79kp9Qjg
9Jj0P25VJF0Ku8P+R+AaX0qP+p3uGQ5tpoStlSBYGmRP6Jqlja6iRhG2PmKewvYB
oqo9NBtL6vO7eFFYw1l1v1ZbSV3sjbWUSd2tqdZ4uky99dvwai6IReqxG6wZoaPF
hausyb/yLim+1J4GdUhUBOTdEX314xxSNtu6Wh1THYjARQijCb9HMg3MVM6e+ioy
AHd/a7UDNIzzxhtf+vfwX4l4QHYXoNLl9ZVgg3clErt7tSsBMuayoVVS4iVD9CBj
94S7YHlP50ffoTQgJOC0vn5arLBZ/ANVf1797R9lrD1R7voz0A7OuD26NTbyIeG/
cw+jVdhf+82lJX9VD9PI+ri7WoWdozZTkazpZCKXxF5PiYqxrU8Miktl0qjIu34J
RwflivdIS5jX0pSkyUAKfYQDx+ZJ19a6eGRKewLlkvCB22+HcBpGr2wcvKsILz5r
xMw24w0edXiGVh4wDG/Lmim7CnvTqMkajmJ8PDo5yHfPtPv3v8vL3Sji5GpR7XGp
Ts4b73VnyC9HaZAqV9ObfSy8xgvItu8TZ6ICCTUQqLnrm1V6jqILOIlJlPZHYTYl
KZJspEcDzK6CXCjCtYjo2NkOpLzA+lsLOJuKGqz+rJTN84LUOeDSSlAzVscd6fgs
TgqDqgn0u/+EPnBWMEXZWu67xsR9c+Lde5aJg5KI2SzU4zqRVesNN9DIsyFBMy58
+vzWySgbHVoNwOVES0MfL7s0eG/iM3JKvoSahdaeIkfcqx00iR5wZa8GF7pVBHP5
RttpH0KnO7FKOprg1gqTuDZGgl/Mwbde/k3cpB9PY18QtlelSngWHA/bQZCtottk
ydVtucI3tPS5jIohvQuLTHtkgmNuQS81oIS7tIi9EIrKaY0ZYsGOTGTLCsVLnjT9
nM9hCMlu2hL8ojK3GJ9cgMf3kVjLTUwsnEFk7+R69CcTRL0F2CrrZN+awWtXqn2K
su9ODI10D1/WnpL76Xgj13hevGcWXq11aVSW2Hs1HhKK6DLbSwSLIbwgCEL+7cq6
sZ+BneoxMqwfPsG27E60Iv1REx0PDqDtf/Hk8ELwmyCBecrrbSxZ6OM4OShlk0gu
WUPOjzj3qLGxiDkFD0INL+FELPQuwrdBC2Lcsqb7cksHOApG4k9QEBVOXbh6jEnJ
OeMpBA5sDd+ewYF7D9MIUYA9eBHmITMWWOwkHghDYMaxhVe6H5NkGmILc7zL3Mkf
Rn4g2X2gmUMjm4COeJHzQpnXsxAE0+PA7+hMVeS0N0zBWbdgvAce5Fx7q2xVCRUt
CNrZFRw38YE8+U4XoGAtsJmuBrUz0Qjp9HVqgPIj81aRT4R7eSxf+PekMsIzhoA7
Gu8QRnprbd9c6hXf8sNWheg+kaIXH3LQonyUWCnllXxK98hhVBLDh0tS+aNlDode
mLOCaETvLyUHqAQfxmG20Sf1m3kip1Cz7canWnwCbVYk22QYAxVSKTA4QQ0NprRj
Wv54OTSHDZZ+78XKHDWr5dmV8zHIWTZfFvBqlI7FnyLdJkSs7RYPSlUxE3pfUgY/
0mV3ESn3oPGjlr0EZ8UsIqobJyY+o4rWlORFjp2rGsOTd/HZ3M78UTV1oDls49WT
Qmyz29rwDR617bXqg9RGigUp/FZLSPXglfy70FmYXTXEaS/w+28q4djqfYW+rwlq
gCVfO5rN9WQauz68Evq2guZAElIvm0OFwsZpvPclFfy7D/OIPheq0HShDf4Go8PO
Q8FFHK/+eIgQLZjCVvvmPBchx2t9AJvLSwTE7CVS6BzlLFwMiVfq55YQ/jJW7vdi
HI3sKvCGxIkiuInhovJFPG6ZLtL7abxPsPphlSkqIi69MipkBaF11gf801qr9pFx
p/inYk2DuLM5k/Awzp40RggDQUqQSwuFgqlkqGwLobQqwvoto2RTZOPJFaXG4qF+
pXAVD0M+B1Q0VFT/vOhqnROGifiWuoDEhFG6frsERcLIwSZtz13NiRz2IeXrJbvx
Z+ixfht79oAxeFr7z9MzuBf68j4ljzKQGIOaafPlIPJpSUah5kMB5n+r4tPeNDV+
NOXl3A8OAbjzQgYJY6awRdWFCZsX8RtTgR52FmXEVT1UsXownp/HmDApigWcBZMa
r2Xwkkm0L+h4ftG9nXdUPAmw+EhZI8jw9ngiIlde74eim86XqPCkTfGqPKWMSKZ3
yCRV1xc4WlrBUULtROgZGmIprjRmiD5QWXPIfWJDSaU0qiv/wR4Q28AXsxWd5UBM
kQcvxJ8q7QtK7/tM+LdCCpOkWG9AkCmDjS2hKe8SY7/KZPMUJlMUx6BKltc99LBq
mKLekiUopvF44wD+qHeEG2oF8ldyGmmmqsDk37fJnxFc9srN9KAdB6D6b2t20UQv
oekIQK7P9V9NT2Qggatu3qebBwR6JClspvPjaOAOrSi3YFzBwt452Lw/+WT5WLnk
dGRQ/apFUmgYx2gp7W8js5moGhKkfoNna86Lm9lpaEiKlZK7Dpvlu7P6ProHExOj
RmgcnUriFQ5HLYPGzvWd9GcRI4mSwYxmmmaPJxmiiEg1i1qvWv+zvTrpJ+ZwQ0cF
NzqBYRBBs5iiC95Yl0WJP9MThmxFX3IyL0A92kcLZ47ee4LchKu6U8aybzoZfWUw
mSn00srcSe0gRLEeDfkFtWdI2ERGHuRTaQZtjpeDPS4i5yAK+lODflactKcsOGh1
C84F1UiTU6TU2kxrx9d5JJIF4CpLR3+cVjbR2kHeFiofo0L98cXhQwBVHEc9ZeeY
XDtcZCr9znrkb4LCBDffEdefrhftvaQslApGhNer9Saty0vDmNfvHH2sI7g8BmpL
zgFxRTYYFVKuOGAltJN+OBzsE0Oa72T6Y9YMSCiWo9P8WDPFIGJ4p8gMaQc8uyUu
ksZdVZgwMo4mff0bnh9S48KR8xACpLq6kAIDyjURnqek3TY7MGrpEKUEHJNyAAAQ
WW025qqtYyjMxQPZVfWfR9B6STumf554QFayf77TRsHfI22mZN8CrB1bffpjPXnS
uDipD2/4s70zaZOy3lvb3SxY3rPD/LxiUhHXbPVPGr3EDxzHcn/Wh5TQYnxNv9Go
PIMZJSnJ3JUQLPrNchuGNU/a4w9HYsWTnWf0o1dmtNu/uGzkyAE3njICJjHqVexN
XZnFpNv4rIje7s+gyfOodI1nxg2gTsUmbKumNDo4KgyrlA+tYTFO6sp2fdHBB0kv
ndKXaWNJIZIsqm1leOr38clRhPSywRH8OqSuxJR90kYIrmbJLTO3yjlinrmbVnBA
4RZ2HoHGKvgHeXS/0hJHXZ9JVIaM9gkI02T/my7Mz3pNnHvCX+MkInIcHm+mWf3r
uBbQF6iaTYldVKpotl87baIo/BsZn0bsikI64tpTRs3zhTOPeOxiNYPS3pVB2+jW
xWfpqr6e18jDkaAdR6Uw/V8l4xUfPDZ2DKpPwwiv715xeIueDuPJ3S0tsV+4a6rJ
kxYVrP+iHENuhZAakJQNLSHV8EZojfkbwaEFsLFxs96kwrf+DPJAPXtyB3tfYJnU
qv9uK2/L82k6zLviKjkJ29ONR03wpgMWuDNXIcKDTI0apPr3TKCYRlNfKulGJBtW
IdY267UP8/zDu4soKjhmD7gWY6sqDIu5GWc10XLwf99bGv/LAw8ipsbV6YtXMk1z
JWu58a+ZE9b5GyGbI5eKWyXlKX4SK2ckh7dbtdjjXN+uEdpNypUCHUmGbmiHHXiK
G4VEOatpdGJbjP/HxHplT0NwxI6xIQUpO4VbwAG86RItkF+b3cpUx55jR+eHJ9VL
kMlljrtHzigXRdyqXlZwJwxscmYaH3H8y/dnGApk/G4Bw7L28IHvb9GPb388dMr0
4+/muVYC9khakdXSB/LOcCrCuBTuJl/LaHnLimpIVzIYVYQ0i0MrPfQtElidO+20
5+Jm7x6oyC5RjxRRcO20jpnFpXoGOowcFs5Swg5ZPtfReBh5LIGvrBa27zKyYVEz
WA8S/BhgyRnRr1fuO+j3uU0mVOWATR/c2rTAVPUOlM35PKAhg/oRnjNgibojee/A
cF5ZtIEkJXLiEjRyh1hLVKVqrrQPn7iplDMuG3VEdt4cwqruyNkf494JWQ5v9b/D
JVLNKI3eHpYJmoy2UtxH1hqc92qgJ09Y7Gt8JERJUunfYqbs/RM1FK6NWtfQYdxv
VGC5DyMT0vJ+1+pRJQWX5wpapju28lAEEsVYWDm3fn4wU74rX77cR2teWZUMJ1f8
TJ/dbsnun0Q9O2DVY3Le3Fn29pOwghMMKccbN0Mcz6BX/lEyDV+41GGYDWDrSfpf
GIkpC00nRFFzH3OgmOTWw8hJK1zw8eqYqhLKeE+QtBz4rilKWd0p/xNW2WBN2yhS
6l78LCogSxU6xeWaiDW0PNeEezjdH78yP5mtiGYwiyjnpOmVMGdOaGtmM+G11Dld
SQt9CwxBzAS7h+/voFDSasnJH9k0pHcyuf+DTQ4ijYBGc1sJ6287wA+Y4SaVvsxw
VeOBEIIKam9f0S7I0ZpX73tDp0KX09DFrhitFN1J3cRUtKt/zSaRiO+X1aO6rtBj
8O5bBzmYp17q3uTWzm2ibyKOHxBC9KE3tsb9IvZKxAYDzeJEtzfLtGmhF7nyj+3j
wfW7eLWE9KGO2NTkcKb/AmwSt7ktPjHp3fp9HAZOf+kuUBRn3yrq616I81zoZ9wd
LXbYL1a/0s7zNea50R0xmEM1j97OhCf+h/ezk1H8Z3/eej7jjFF9GmNwSjLVzeuW
LxHSScrF/e24Awkmsb0Z7v4z37r104lzeQtG8pBTLuM/bQgIDY9os6jIf5Fi4OCj
pJaNkSp5OKbY1dsIJy++DAsIc5wkz1f1n737TNJB0G4ap1nY/B1011W0cYpqCVTw
0t/Ao4VKjAalAtre+TGTAe+epIQDTHdm11uj0YHk1B5eO2BvVv5/2TlErpsLJ1Ll
R2on8gW2GpfEqtVbfn+q9GU4O1/eXKo5bKRk+DVJNy8m2MRly7AVBmMYYs3/exWI
BH6u6XxnnZKkHmHbr3JvQHcEiXKwoZBBtIrSG6sBp2jyT6rAKmMGXktBnds8XmRP
bime3X4bj5HFxzs5OHkJWDSeqM3c9eyVmOrdeHGNNnrnwUoIVsBQJHgcqFUF5pvS
ni8HjhhTXtaNWQCss5qRAKdlciNHj8dOEf2r75AItSJuWfMn3vSLJfs6ZY9bBd2g
KOSZeysTCx4Qavb/sQkgl3yPPkrdu2eR/QG8bLumxkFIc8Ke8F7FhS4e1y3Jh4Qy
eugntSA2XqgkKD/HiZQKviNh7D10aeXXDdU1iyXxwpbkqkI/wWEmVzBoz4veMk8y
OPo18aV2EXiblAiLjaf9vd9mXikL5JriU/BCm00tCvgBIdFwmUytAfyZ2O0FoVif
YSLm9ANElmvj8NAJjBj91CPi7Qyb/MvMeXWmoXsonb9m20p3gIisG+FgcjOJZh87
ntncKCcE/OrqAzObV0KCLdAU2+gf9hNY0pyq+L+VuhHr2xqSNb0G6C8WX3+Afn9/
/Vo6AaWIoeZZg0T7zey28GnXSPmRXheLrCu2ESpYSlhFf1MGj6tSE/UX8f43hdGY
fN5SZkm28fVu2jh4niDZXzkxPwE//T5FqC9VxSIgjgg7fIfPnqh2vTQApHPGRpbN
1yMIBN/wpviy7ArPchro/jFZtsjvJnWIpsGcM4AxhQ0Noo4bhzdJjyp9AKoaWHR/
ZtWN1JeojgH8lZm3zmsJ2GxlgztHZAYK/yoHRLroj/54XmI2jNV6bNeHUEBllo0I
d8EJ7LYa4cYId7eheoP15bwd9Amxq1i1DfD0UYoZgYVHUgItUc4oLlqEl1r+TO74
+49hYQEgZu93fqWN0r2dfWROwt4eVhMbvWbcYaHMMWAfxOIkwdKbj5EFBUcy9OAC
ZPObyCm+//uyWrn9OdK3TBpQg1dCFkf3Q790A6h80ZPmcYVqCPaBy8E9BURIpk04
v3Xa2ImL7YxVXeq5d7Bj0/3Y1d2B+j6ikD/5MdRLdtBNqfJNAC4tTUco3woCkJYT
Vwiol0lkIHDB+EbJdTBKnOQ7Fs6Ahe2a7hV8HthkYOF+BjSOlQJN+hUqSix2FFGC
EPHu9CLRFJFVbSxulfbqh2hH/9hWqzlfGpycGjchKnNZRqWwGNiyfgNBpThuai02
RXkLxjLPiwl2s/vFRgoc9C8KA+fyVyDBwq4idz2EU8ZiIOsJc+1yMJoFm7iwFM3j
Ax85Xin4DhtNoXJDJ0tUgC4Hs+YjITPXqEI/jg5UNCA8eoaKuQIOwO4sSv5Ypd2i
a6B+1ZioZLwO+ICaUqzEmpgqnvRU648cjOmoDC8p2JJSi/gG/PJS5Oqf/2ypo3Vv
qYPgo2Nmkri0K0tveVnMyvM9b61oflglEuDv8PipwyTsoV23d/yF/ZHvyJCGlX3Q
nD0feEiUVJb+tGpjoFTbAYyliYhZ//+QaHKI/Ec7XgE638yeMgwbPZkSBkf9dUCS
fd/DE8nIcdXAs8l5mhCm5Gyxl2uQmzQEgLc4brw7f5tKOUXKJde5HcZw9J54o6NN
IYG1edjv6owJGiJbMyRG3873Kpo7jdAveeVxDFEH3ct/z+/AA5eNQXURRo1XdYP8
8kMAjryIQQTesTKu6M6z0c/CQHbNX2l5N7UlKIz6leRvev1DS2+ILxjHV0OMxUjY
4VB22Z7IoCmN1aIdQ/M/IEMZHPnJFK4dord+9tB8ocpQhWB1IQVfgkbwByl8zlDR
A7aPpAthiEFLEUimJDcaGuUne45xmmT+/2LzZjLidahuMd9qvM8GLp31iJhqsJoW
lS3Zw6kedZ9ob7hpQNSJcXosG192dUUhYZ+Ierxz+FjtPhsNp5mfSq/8VR3z5WTO
dbBvLumcYcGFlXV+umLqjje6maO5RhChzfv+QRKN+uFPGqPDZMAe9yYEqLHN6XJw
CBQssqrAQxHpVW1C/77qn95B239Plos+BH+dSI67IoGLHhcVAoAbzSBU1zaoqXjO
ku7yU/ZuNkMMzGb5nrnFzSkRW7fAD1V0hSejcV2PVLqDlHeUQI7jmFpJ94U/K1Xu
q2OtqLlvlJ2nWC8dM6J9PO/ICml3yOq3sBvYDEEEfTJ/L97iqBw/LLqCWWv7dXyZ
n8pWRZcThd82wrydC2pbqCRnl93llH2dN2MaOSvz3XLUSASzkwsM/t2pihN4CtI3
dI8+uMJ3ljtuYnKuW8nmrn958CQ3649MKgtNfgiDl5I9vZePd3gcYeAMezlQdAoB
95HfkZRJhsSvXaWF4kvsAw8AePItvH1A+Cw7/7iuVHZpYRzHUcG/zNm/kvq2MU0V
kkDvVPuFXExxf/9vX0IMlAid40EGSXeWAb+TOaCZ1FQWXMUCqHzHK1LpKdqYxK+U
0terD5ChO+fFiLYZvexOg9xq7qJHbKRRuL7OqCeomXO1ZyWiRAOYNhF21oXi8CKh
kSq6F5Twx28oYwIVSMEBUwbQZ7urBgX1bY3w68gW5nCV8ZjuDOcU+JZW3f4XTBcU
uZBAOBh0Pcrih7lcxlXEnNUyCNU9OKtYdZPTY/lqil3cv/tBe6K25uPL20gY/hH3
6u5KIloS4NN6L/UPehm4pDAGbmuzUreUAboGkSRLZA8owOHmnfwWKUno4D1wudzP
8FwVOCKfWeFZ9j1UqxdEm0eZy5+lnK8VBGajOIOxH+0VGr1bmxG6XAaWyHsREttN
kKXqX4W/8fy+b89LVVmSqc5cZq8IMS7umhFYgoencSxCsqWTZgPlZyPWy9SeAC0w
0v9M1d009nsvjKSD9tOhShWfHKCdceyr8HGKoE0bI9hFr9intLcuEHO8h93f+o3G
KevZPfU0VyQBulh1N3mkIgQKsn9v7klofntViR5J0rRXaMo7GQR+ydJyzQepiUiO
+eppMLNmpSrHnwRq6tAlnCu9yvmu7Vh9FgpeHf3WQLvBdY/R9k31a7IiPo7JhCuh
blZShWkKfqOsPmctgk75X/9uLMDcxKGfCClvzdzaLg1NLSyuo7BuLJ9RJvXbS0IU
0UZFnSKvDDVvnvrk/Ex/d2a/9Ic8Wep3f90xsKRmUkrfA/bdzBhPOnqiuPtN/xns
rX48SpS4GDbCOz0JYpJ19dEFR2LjkepuBtl1lmsvpVhMfWy3p/RTA0GplD3+mKFf
R4FOmOS/d2yBVwvpdmUQdvRwbBZSsFqDMegBsRW9bzhUqCYLCf7lLEHM4vYiarHD
J9ntE2oZkn0XNnqABW1xCIiLMNm8zdWegWusdEz0SdPdmpnUf5S6RQXguDqFkcqG
0Vj/Ji6E/SWhfznzYvz2FyiP9UfyGDigUAwXExQOL+QeWfIdcGkBrf3wx/lN1uQc
68kUA/FUuATZjemgMwyDR19rc53koCipAISvDP2J7SsAH2UsBTZ9ROkJNQmMFW5h
+ZCse3I5dNPgfiJSWAPCOCODf3J8VJ5WG1MBkneRlt21Eoap77hNS1HftL2ib8V6
fOZdFryY4vY+0VAy02kamGHJfVWpaiOuy4/75Bx+EDPZuQnt9gKCpQAh2UbVHoks
B8B4SBykpyQrk0KWio46anPztqBLWriAXlk37AgEAH2Y1i3kp9khKbGFQ0EGsclf
eD7u+HhPXFmbCRHiNMd7FtYewRMV9nIhlyyBHY5OuLfKtBluU7g/iwPXdcgM22pU
YvzD8yz1tpMUiMI1GLMZPG9ckupS9m984o8ZAgZaRgq11F5W17MwvaKbbkhcYsc0
xFxM4VqgNzbbCRxhFdjve3R3UVJAIcIggyLZG33nFuLwmFxkzXAd4S+xdf3NOuRR
BJRzpeqgb/DdV366Y9Tq1gYmvP9avKdzG493jKU4JsN5PEQdmorkwVT2cwHg6TPS
7BXvncrz4sSHvBpMjVugfpzXGUPAt+HSDy9fZdeEnETnsYTQv+TQ9uJymzLHkS/N
7NRt6YlLNMRRcEXv5BiihEhslOfXb83JAurvhFWoZpBlJzgBvkyX5NLnsKs5Txvl
dJtm4NVbPVfTWwGQoofAWDW2zTVtlVnIjp45ZQRgPewSS7dFQppDLklimCUeTo7Y
POGbfkOH09Up9nHP/cvcUGn68oTwfE3kvcaan/CpJgwXnTU/QbgxWy629Niv2Apc
BNtK+qnnS3EZDFYWyNCbIg4kGTDcVnylv0OGuKjS0NYN5iLJvbslw1GbDKkKx5mX
cUkHSt/vgZ6gbu/xuZ3jh9KtoGOxRRfVuCqqeiWIRwOiTAsbsts9asbmJOPWrguU
e1N8ZkzGup3z5eHAnxmEJAnYHu8m3SY/2YnhVoeHffgKyGcL9xzBQbkEc5tv7uvF
spRfibT+RgYL8NUHnswbckwvkBjEkuR5+8k8KCZpCINdSf32RP2d9a1GSEFOekho
5TcBDG/pmqAiW+nRVVxT4eS88+UHZR25BivqHw4o4H4AqjUG7d5J6vfD9SNgmnCi
Pn5F3vdLbkV6QL5+uUCzt9QTnXyGZnpF6yB+rfa8C6AcmSj/2hob2/+yt6qC/4UJ
rBw/YG9wKufRnOC6Fnt7xl2JGN2nKGdlg5q1x47aBe1B5z3vGax0Wf8QNZZffNed
O3GVdZDY+XGq9kKjewB4j856ENViWyWlfhyBv5Yz5dhme8VMtXxCUnOzNsa41bdB
kCQExuxLDpwjHuicae89ba8vF6fDYkS/mlSvbjRPfu6JTsGhLeqN1WUcLgi4YU5f
B8IwgNWIsUexQ5WE1/7URU/dz2zcYlTuRTMGKMombFUBjf1xAB2pp/ti5tB5kK1t
rtNYl3k1LdQEB6IcRIcKj0EJfdRiZXbaqq1OQeHmxMhvZhv+BlhgsIT2ugfuVVAC
IYptDBr+NnkMWgz9kGbci/Lz9jcL31tElktYbrZBhG81P5uCu11BcoPmYJv7QIzH
vBEF/+/5/jMYlxUsnKeaAfGMMBSLveRJanED2PXfVVLqwTPMjWQgKlwNsRdMd2Xs
GqQ3qyVTWmhsua3FoVNTtRjDbJ/zMRmqki3wWFm4om0DGURlDoh+wPnSJIEvLDcU
qmy7jIzlLrJrsHBlgpo0O7vggb61nbDy9dqqcQdR2wGNq6CST/iG344iGcgVGvvl
H2ukcClc+Xwu/tsUui/0cdU1kWQ6bS6Z+HtWzRdv71dO8I3WYeNH7H6qBdS1Yc0m
fsrUg6sLIol5XEAUBSAdUaA50sqwkGDlWZR/BdChiQxKNvW9qoXSe4IoIipxStoB
nIztJ5YBTv08C4TZpYe6hEYj7vU3fnSu254cxrIZLLyHNzzzlU86EJ4BhlycsGjF
2A+I7uS1PujZ0KrZIPQUsnU59LF+uTQI/1E26uXHQzqMdyBUBsPpdXQQgBQTBDmH
aRf8cUx7QSYmh7oPL8FS6X1loLb/LfMF240bpw6NWLKfinNjlmRD8RqYj9GxqzMs
3xrehbWDlDHJL2kk1zrj2WnOdfKaBC0Q5q+ifIIJY2ux1jMegPnWgdifyoW0fsck
a2mDbTGcbCVemBzcBr7b42srYh+/GLfrH9s+mDfqHu3C7KVDmJg1iOTT+OaP1Frx
5NQ88Wdx9rGimmUJzomj6hSpvXm/H6TbTs0JP73uAvP+cvtzBhY+j4eBrIgV3Zru
Yv3FbEtcSdZTZpJA3gt7ddN3pFOKi+E7M1pSulZWGS8MvauvWTOXcFhCuyjbDwu/
DZGDj5yolcEYwKIxnsQ6qqAEuje8id7R4axTARz/FAEZkgbAoVsIOwPvEKV/j8DT
lwiX1J+6iX3ykx4APP3hz0YrW3faogpBCXufyc1MIbPkXKNJbF8ResG6xz2cIfd0
aYE0y/uJzncatNMwzoltb89YfxWNtg0t+cXFXnivoEPp7+PrsoC0oVqcT/aN4bbA
d+xHj3ryC6GyAv9ueh2C0g49SU0HLIfW8MGgjX5mMSfsMmTUlNwsS8r0GvVoQRZq
L86PypOIzPIRo0600VzdU8+i2PbtokuRnYwg+ZHQPrgDhkWNuEdD6aT9NrhJTe7y
mAFtSlgJYm6EyECRPHqH4dslBVuatCjpo4pR3wzWaqzwmqxGF9XKoPJWAa5p6YWC
lupnTpyW3O7fHEDBEzYI/iWQzfTo5Dt5Y7mSrlPRauOgEGIbvfeFYdOvQaU1RN5n
VeFEFpj8qpub2+vqZPDsiL0pALRZPqOFhEPAmuYdqzPNEy2STV/arnoYwqeYLtoB
SDMdltbonaMVjF1vD/aQw+CzAiaKj01X965pS8ZrWqB+6LT8BnFUXLopgStaNmsu
DARJEGKsP/6jJi1IbNIxg5uPtMVY4Whn/hn9UGjNukdh1/zujgKaddmZLNwsdHRn
YlLHEw7y2WB86vfFGPtS4Cmig74JGbLQgF6wnk1X8xvMcDZkG9Q4MIl7DCA7qPnD
ottxbaUzmjyiMT+ud8P+AlzM39A4mndb482n3ZQq+yzHnZXOUJgo8OTY17tFMIXI
WWDCxWXUtVn8mmTtpcF9Oj1NkbfvVKrDiQk1ZdQ5BNOnunMRooBQ/n2DFw+OmaD+
Q4S2SRzo9L4Duj/rPIeEVq7y+Mmqxz9oQeJmm2WA02c1y4CbyFt99efR1IY5vtPJ
o27BAX9mDzWb3ac7zrxgXhQASTGMxktIWrHzprhCnEn2z4Breijco7u+LU4QlC/z
RfvNWBCdZblHBqpaNvGPdPQu3eefW78ZrhZ3suM4DugRuVGW7NI9UbE5fgMGPDCz
ZB0WH4Z7x10MPzK4zA7A9LHrBiovOtll/26qVS7aHZAwn+dOfUl+gxKr/xoVHq7p
lSIgHdFlL/2oCJDREC3XWkkeLoYs4buJl2XFwGh5/J0jWvwqCeX5nta0eX697x3p
HT54+6Ifc/aiK6aebmWxtuKlPZhlLQTvMAyxtRk5IDk7BSI9stIyMIHOPrCksAHU
9UYLwoSaBg1ZHNlPgvNYO87hGHIwUefdts+po4BosIv1RPUXrerZcJz81q0iOQ8B
p7t7tSMak5oBESashQ2uwiUmW0I0RP7Lj8HtdPLXBBbn9raHXC8C35YrIjJCRiLj
/2n6QB1DveWxo5e9xC/qdXSobVr5S6hOEyfEH2Byw/sPzpAAxvniUxHXvHm7h/vE
Rn/hO3UZpA9b6E7BH5V+58ZPZcsekWvzEQkJ2kVPBNDDRMQnFkhoCHkXuzMLAPUz
CHHx4YhlgoXXm6ryVd0Krl4yIgAngrSjrqnSnWvSLa9gSoLxjab9aAz8YzCBfGA9
DWj0u7WRRGjGK3fw/ruALHQwKpdacMcNJzZpCthTQ4aXlgFIl8Was50GcZDGM2gc
/rbqGrOZ1puT3pFiXZREA60/xeXaJRu/LQisQxj1bFwPR9750WKvrrsSwrlqrIv/
OFCQax8Dp/UWVdKS6sqfH956rmmkGUASSnlY9/b1uB3v86M1MLZFgfwhyKjIAkY/
Df/gAlW6EU0Ilv5lkNIpeuKAnf3UxHb5BP3I5ShL+Q1goiYAZmCK0Y+e29j1ocEv
xSlRpQyw8ymWkZrAEUj++ExxI/gIiO27jSwOnWN8HLJ10VdgPZa3dHio0uxO+liN
2TzSkzMzUMsrsEDFmFnuj++eSO8J9mJW36O9ABQiYffOAHfy2MI+MS3SBFpQBKfC
JaSTYQquSaTHfKS1BwpiuFJ7F9FZeGEAoH4qRZks2s/X2Nq5s5BkXPmIRjlSi5H6
MtFazfuv/MTW9zNpgR8VsiNFl3KjQrgsUsjVwRh1w2ydmc23/6SiYu/WdxoC7rAq
5MSyIeztiJ09tI9CcNypGai0Q1FdE0OepB3AfNR7Xvr3VmR/rYBaP6L7zhpOXA08
SL0pq1+5eJVrWXnuHXfNPSGIMWtqoxH72GiFV8FMJ38/7icieYrtnUYd3U6/wYi8
3H7JLCjkHa89EV3PwNfhXrSeIikdTwWclv3j77hhBCIX+Q8zZXdn/+i1oBdUSi3x
GmK0u+apyy/kahu6qqJV+spFiAeqa6EzHDWcUJLi9uCK9L0jwgIjgvf9VotdHCuF
F3vISk30TxJ75UNBvbdBpVfCfL7Mc3IHaHWmH6GtMw1doxcnXjrVqnenWBU4jGi/
Nl05fXfBhEgdjtwXQOU300ZtlIswdlzutpfDr592Yz8yycR6qlSuOMeYGw7qXVYJ
eAfjKpzsTipOUfB1kPtN1harVg3Bro7dL4x3+HVwEruABoGUQaAPLJB5JJvQvHk8
37OoGresLjHF+rio+FZs8fMmmFFsjhAh4RrKc2FCS9YPfkhIzf8StE8+Pvln01gL
iNecEOv72g844yar5vmKmWNfxz2R32xzadvpiVRS7MHgGLrGhxfiAx7tcsnNHsjx
kxtFpMB/MxgNUMDI+CCMux9K1gN28QNwn3yb4848x/QlkbhP1ZQG1vXWcs9wm3Q2
cELlYhzvDxYSzWi0WTB0S5tUJDP6kcbipy1G6DmUYAG0C+YEqvtj7rjYcnjIGW+k
Pa5fL+wkHLG6/qJv6cxLst4qMVLoG9rUzSuIfoFVDOuEPB2zsAWxmRBDVFOAG3zC
/PlNrCqXuMp2Ug3sa2I1NlbejwHtx2JA0AL0aXZopvPZR+4yen2wb7PfbPsLfVbm
3gWEzRc/L8xUbq660SJkBscNI96cIPemUAGI1n5m2cgA1UKEuEgX1ioeKYqC3c+u
FWUcmpFiHD/JMoItIHUhs9jAanGdEUhTbVisWCd3rC0iRedEg6kXLD67NBppIk/J
u7SxtS20Nd9AMjz+bIzdvi48gOc9gukpgi+4DWFcUC8VGlXzgRG10nZffxSI5DvC
2jlui7/T2FS0hAp4OOjnQ71C+bw43yKYhNpRA6ljv3m4U43BiAEpI4pFDm2z6QTU
Wm6OT2E6lGC3+jPIk1AHKa90/DCyiNleY/Te7tX0Y1bP8j/dA5ohwg5XeFz8uYz8
VFlbkcobNW/yUieC9DLGeaShj67klfdzAbe7piDmreGPlkSEsIh+T3l4nochXknV
hn/Sc9IJ+1XF6mWZIV32d30pi4UmpWO9qneVWX1SWWyazEGPxmW/dstCck5Y9KhY
r9YqZnwsWfAYBaRGXpYuBWUJdr14D4hkhctMe8XeUbCBanIiZvcMKVFDTcf2ewsO
QQAqGOe5LCveXzUhiGApdQ44rHN7TlCueVx3hAF20m+gIfBI2lOdanX4PX4P73mM
27Saj4VX8XCppEUVqd7c6xaL9Pke/UapviU/FS3j+9aTYnLp6gMaAaegxgyi8/8H
LqbpD8VdbbwHHCd+tJQnXNgpyWuFbQbdf4ED8rghlYX6pvHfk4Mm82wcseFTSl2T
lb4vWR6ZArY8Rb+oMmpkrEk3RqDlAdDwqDvhcHum006PHqe2ubVuKRTTPaDt5B0z
7bpy7/VNsEuyu3PFXsjF4yhteNgUPAm0yN14kICYVjt2Vg6eO//i/LnR2uHzo/S0
1uQ/9A6U673P4EIj14Vueumn9vinUgDANyMHYFl5KQyOcjqgz9P1FeyBAZmbRXgf
DNyoAOyACHpxTbJkz/HDUB7dddaeKzo1yyyTA98kFAaIOucbir87KjU8SqdmqCr5
IZst2TCdweK4DxvuLaVFAyREdvXgRgLtTDTq4bZDAAf4Sm420sjnbK9e9HDY0za0
j7VyPTdOBX07/nptwyz7Q/pWkl3EDsv4R/aBvyLWrKS9sVJ97KfOLbiPrMDa274W
4ejQ+9T0P9M8Y5kz/Q+/xbK6XIqkbz6yNBvvMKEvkuGkBUcivBnKs3dwKIaX0DB/
VEf71YqQCPq09cKpTSL1hiAQyv6dNmgQF1HXBMTKSMkJIP2yE9JVhfxPzlvzY2IE
l/uC0vRdyormXPPp2FsxM5CIgXDfeq0/12GOvyLWfYKj+yYq6U3uYxvjPAf31krJ
HtVJSkuwK9V/cSQMwwse8RPyhsYVMgL+oyMpq0drBPmj7burnRAzI4IACAHaohyY
WWZh1PEn/KdfntT3noYkLoqGiYOC5u3svpZ+rdBKlPLqiocKj811xhkzxsjlshxh
yIQbHzmsohALXbIEuvS4Weo6BhZ4B/BrWJLM13TQDU25yyaCEM8sdMJfGRSMvURN
IIHW+4GnDgJDwLGODho5K8wD21MYOx/WJZoMdnUKIPLinJmy2bPaSWdr/G82bBxf
hqdeXRBH75HHNCn9I2K7qHQRxCpm0EFSfkWyIgLWsHc+XeKEswRkxq4uIHlGMXrT
CzYo6MgZ1iQe+G8iin8AobLNamP3UKqKgnpJjjYT/lcYvbqH4YI5IUigOvqlAwxO
FKjU9/BunqgVtZzoVR8d5pBk05ADGYw06vrHLNx1GCQF2T3cFpyqcQjnRFwBVu4m
UbilidlyFeCc5l3nLtCPwPomUENRgvfY8osC9EtNHhi+29UoUusGqw1pxqGoUn2d
4AZDMbgs2kfIjiHZWTxMr0/DAM4w7/2eusyWUlVqO75GQhGDDDJRuNVnKwRuOHom
cEp/0Rrk/JW6J85NN9asJDjo2/uHoCt/N7zyZTJx9z2t3tfuFI+W0NtRGmah2cKI
SZqKXp0sG7LHcemMZjIq5b8j1HScxEqk3+appStTPnVOWghHBqQOK+FdDEK7YAJW
+Fse0+8FytGgqvU5JsLD9QhafFN+BF/1g7w5Vcrwp0GQRQvoq8w2qDYm2GPII/D1
MZaGNenbeNRBdRIjY6WtCOGi44FLv1ijqh2fAx+PRI3Df+gsbcJi0QEcTdUo80XM
g8VLNodcR7RCL1mr7l8EXRoJyR80qJ4/8IIOPeUiWD/H/uba6VryCEceltcTfQ3m
tVHtLUKxeYU2FAIwD1dBQDqfYGQc77Z+CLJ9RGlfTVjDSLiqF31KYO7xR5XgWSgA
ZBZSAvxh3Od7JEUxrVkdNxRY+fNAaPk95w2lkJ2ICSn/HYHUyI77aYlgMOWI4l3Z
92pggwhi4AGRwQWUOykjXzq0wfr+Y0MFMMY0O/tHR5MQIR8MgKAx8GLoySl5qswi
nfO46+6XYIJKbduGn0yhnhnLNe/5J3KQSelV70axbXSKlIIIASYG7KIMc0RmZYUc
QEqBNQkXuRD27ek1SSk4xeo1Zfhr5O8Vl8AMVShZvW1rjTlfudu/VCKSkkjJvpMy
keXX+l6TZx7w6PiEwvQVR0womvf4jRKthVfHr7n2/xDbTrJmkesUWndp7IllCnaE
46iXJyTqhgRL6sm+jvKx01FxtMF4pmSf32kEFy3uqJrKEP62yBRQY3ymnU0b5epx
TRtEyKr6HM5LAIU97X0ztm95fTOlvIz7IMTHCmMhkczpS32UUqz9c7D+dBiuBZGM
XIXSM3v6/E2ciSvAgTMLQ2QdIdBJxcKOIGmIwHHibMebi0BAnop6qw2k8EW1nRPE
uXYi0oKM+XCkpEldLmxtKqimCcOyuN32qpGyEJa2RIE3sGpukQdp9BB6ZR/Sj+aZ
CLSYdwMtswf0JHkBE6kezxlx/UVB8RYGW/kjay23mhC5s93sP7dVosGyAsaB8nHr
yEOqBL9/LvN8L9du7HxEYsXNDA0xGC+5zcO11HNSF4+e2cNcmyO3fZ3YjN6dgfvg
y/8H9m/rrgg9fNPyfO2XpzLbz0ytfEQk/C9UnDSZHXLhDi/1hK9JsmTNUUEVH8VB
DM9s40NokjW7B+Q1iTH8hsfOobq602XdcyxqWxltPfDPUhIBQ1Kwia4SH4aKVN0+
Qf8EhhtNAT7s6/pNMy6OZuJe+C+xR8xf4jThObXVTCfFvV75GRNK5jZMyv1/fV0A
7+TDUxdH5Loku2E/1ysWdM35psZy2vvPOspCNIBFZsJPBFRmXHtYqJ9jrP/TLfaZ
ysnZ6EiGIWbxFuwYOxGAl358qs87aRjZXXVp3t232bR8C+v8TBm6KZ3fOg8PTLpQ
4qLumAUzi7WdKEBSJ8ncNXJR2d/8a2mpADrfAH4rwoLgyaHUGQ3veuNJOxsCirLn
CyuK1jR1+H+7PPppISo7O9qOnhJqtVSn3+bwQAzXzOMWIPd/A0eyRX7AaD5hcV74
MYPbISJlCuGhi+nP2WXTRTJ7kSCsHP7CckLFzQNuvwx4RL1zHITqlw/BUb6vDTyl
cjza0R4ZzaR1LpGIj45UlOzbVpWUtTcjqtS7eL30UevjGPYKGJu+AYMSL2PajyN0
onya0WBLXqiOHlSMcaKVXaFbnVPOjpVyHVE3lQQngbsKMJz0YdxjctYoowVohBpM
Urk0tPA5OS5yEsyBFX5/IslIiwr5plcSzOd9Yrq7PbYwXqWEBcoxy2rxa+pfi2xc
QJynHnQUIB3LtBrraj8zSFo3JV7IA76ufJiNwJgm+zXXrYkLQcCvAUOm42M9ilLu
YuBK1lE4S+jCloQMeWXkJqnMKj6tnZvHyKpQQi82RThTkJRhxpZb4J5j6M+T10jt
PDeNNSmd0ybABMwQiUzoDlDkWx5OkGhh/PPAhyP3qlxSa5KJ+0djss+5PWTWYg2r
evA/quZSmmCG0NRpItQn/odrdNixXJE+P/UoZIx4BdrU+w7cs4/7tN0CXfHNbNN1
dSjWIsME4v62AI7UtJF2NRDMcJIsvLuF8Cqrd9esXTXA2m5ex27Xu+B+gZxVCKvZ
b0kUidiFh7Ge8hYbaKyvNGowyWn7LgEuvJoNdpvfbe2zH/iE4Kr/UNKd9uDbMVvT
x8urm7a0GDr8W/4vA2YFMJYX61WaPCaKcl1/F6YlAmxWBnpLiAxe2VhFMIZGFR4n
CdINE/COnDl3S2fS6+WsFAZdpIhjDa5Xog865KGFJaVlLQ1igjrm9DNgIKx0F9qK
/oK/M1v1g22hQn9JRO/wQHpHMRzYbb+iGjasp+l8UtGbEYSK7BI4p2Uf6lZAKamg
M+loal+p4X/cSpIiJVo9JlZCx581J5/NxbOSz+QiylaLYxgV2v/X1DcwFYXqbeEc
dnsN29JcwiAySRsHHH9G4phNIhpFSa2ieSvvjf0mk2CsH+PC1qoikNIjsYZfAjQC
vHU3uzTZB6FT6QI+CwoLuFjE4ggcTGEB2fMnGG/qGFJcSmB65G77zEcV/aAQ1Rb1
cNdXCRpN1qH6M5Mir/qKQQP6oBjoDZGofZpu7U0RsBJfygli9ZAwwEJ1N4c6bdMc
KdPBGbsM3N8Roo4dvps1VAPBRWnMjacAJqRZOr5yfkMTJgAKLwJoJ4fukUrqIREY
uYUrs0DV+oWvEi3B8OPXfukL2Sq3LhHMadAO7W8tOqV4TXX1CDrRI8TwU+S0TLpJ
vFHnBztBhaUo1PCYsiKxLBZ10yf0lhtxoLcEl5W6lWLl/Un60jByXW+LrD0xfPIK
IhOOjMSWbdQwboRveZvTH27WlKWtOlNsxipw9T9Ybn8knCUC6Mo4NOudxnpQLB2f
eOKrFzWs78Hr7QdF5gSpZHp+ZeyJlW0NTncS/LPU6AeObdPIKT6M07x+OLEyRvmF
o+4j385lyzvWceKcypS5nJj4DmlFi3Yfwz5XNWI+uSmIPah2p6B/B5/eyRR9TF3R
Yybpp+S/kBp4U4Uxk8PwZCSLL6gzfQTMvcvTJe6ki90oHPKRVCBq041u3WWi0TM8
hfdR5VY5NbwuFX6DHka9Xv4UGyzrGAxYcVZu7upRC302+ym3EyIuZopzitsvroSe
uiPD37qfqa954W3UY0pSI8wWD+3YOmwpo1G0VTtKsap91BR/LfxpYMOgxKSqw/Vq
1wIVI/TFn54zkDZJMApefo0n7kVWsGh6TPvAzQyERcvbvd1Z99EWE/ZwRF6WT1rD
U+zst7ywQxOhUUAhHsUFTv2zAH/bWNVFawWELjrdKKVzyLggPR8LGcQ4UU9zllFq
AS0dH3w1J0UwO0XAdktDBM7qjR8UKNINARAkpCLmWLsVFSDMayhwBfC9S/rxWhry
j24OAAQgfpQ0JHucOsqedeF4b+u971i1SZhp3++77tQKtDMuHrl3ztxdk33a8a/y
pQYAZudWOlRdtwX7p1OLgYeeyRaLxJg3RTuNNB523o+qH6iIhHnk238gG3OQskNH
vM/3z6TRJ81QFMJEWqkMuJ/yDorcG+H2Wj/JOHLRqK4E9QLqUIuhNS/GFgYij+k7
csX6NzEirRZAsuJ3UnDNGRXjEPJsqJeGaQYOl7pfd3D+t7KFC4RZ+tkjO3O09eK8
M0aHkumtPU/3obG36m+v3OTNbPQ+LcEgDbooJ7K3kpbMaK0RFhdGpt4wZGAFTNrD
usBYgu+QNQ7rHM0+iLul50+UzJTUt8My+iRL6gIinSTQRinU1iiKiTl206SoNFt3
caPaMoY/CfncQlGHv4jQAVTqnG22aJ98rY8YbhUUcCvmXK97J2Db6eIvxBQmJk+A
4HumqBqtZnINV39Fx7qMomQbUD8/9UK72hmonH0DiD3JuAqw4DwdWo7qcKACaTMQ
uYYQ/H5A+ZlrtnTvgficki069C1o80r1QBZGIoY6zMl2xdJcqNPCx7XgE5n6taBE
2mI0z13n+AVN1ETdxuXZOvTb0yEItgyLSFccAVTMzv4bEO0s/s9ph3WUESCsI7n5
hv7cc3TIBac6VjcDQ8uop8zxPuddCTWWCmIn3FAtoJiCVF45q+Nn99DiFybBzsCN
wjsPN7+3xaPWWaNmUjl3kLFoWoiaRV0TI81zTZUXNOF1E1uzUMUNLQ9EejOC1yLz
DNOOOv2jFCZANGfy5S+OGmpGcPZoZ008zbSMnQONGZU5zIIYWbu5l/tKO/ULmGEr
7CFUwvH6MuW8t1cDzvfo76XPIuO1PdO65zgl/gHyJQiO6lP70MTFdb884iAwhpf3
U16i0zCcaxwKIR5fUV6Z7FZJ2dPYwl2fbyO6iZkPmaX1QXgfb+Hsby+3uBORQAtJ
xIDH2Vbh2MiL9Mz733E7HVY50HBlg/ZEDWwFdVkCHyF7YNf8uMwrG/OpbkMvM0tu
wGHzFnkrlTX3XQWEH8kBCDssvnr6Fil1xNS5EGX3skFOZpUywaZdoKdTLSeX/A9B
C99klZb3A3Zu3SeEIW4LgYtWNlwf+q4avLprAeusPvkvAAfC89rD+phHa4RWvj2R
51D5roAtn343AAcWrG3WdUx/oXKSW8kcelEvMc2RdPV1nt39NcHIlcIOI9H/nZv0
qVSRVqhr68oJOLgz+yhF5Nw+Pngfcq4eyc6kV0WuXHgpdBlLZlrgtm+OuTz9R/xk
WWEx6gQOs5oXgw662a7ynLxYblokniiMjujUN9CWYpi7dnaQVaQJJb6jc0ev8f3Q
ErYyblo/fCPTztdIKN/uJvAlmk9XhR4t7tWpd8UAgje0tLoI/Ch1fZw0sChSYq/b
Hm1J5XmGOccSfFfGhlLkIfGqw0XQZB9RCYc/9X2PicjEyhFPKwaBRNk8HuYVqbaQ
nqDH7KSt6kc9ad0L1PZN53ssG2tblLsYlJj7D+5lPvlZQV8MfRNQBviHW73FU8L6
LW9zrLuAvJ8imsDyroWvu5nDPdWieZbCmZDqE16dbjOSMCC//sgTnYp2mBbdYwSb
P7KX5Ua/y0kX9zJwABrHsGDEF3e/ypR9CpNteHQFQQ/9Mv9zfZ46VjH13PfymZ6B
V/CvVPKpjKRyiDnKdzOGjjMbPA7hqSa77sY7JN7J8jzjXfH5T5p5v2L8ClAyt936
+P2xSK8BPzJ+hpWrCq1HkSw6oxd0sqRMd7i09XhBTEDWWwuuPyRASVWWztVXkbuP
bhzbmVIWeVX2A9p8CLjDMAJE+JwEi1YP+btWQJ1o5z1UDfQi++2l92YG+qQu/gkA
mrPrfXNLGSJ4X5LNfR/uEy8m/qyhSuBSxMoyxTyy+i+N7QccsqqxNwLNtUmmNdZW
bfUz6lCA0pybuId5Z3eOUXXU4mijdaPtao7MU6b05q+CrVlRpip7gbyJ74EevNTd
uBnfwcqVK1gsZhINpoW9NLPgPKricD/Cq0zVdrAe4HAKJx9/uYN+mru7H1fRo1NM
PZ6VDU7QcN4EydjIdH4T81L+CKS4Q801zXQe4EHchagmAOfJdUqcMElNH/rR+LBn
kFOr3lgjvXPpZMOStWYUQqlApY0UPq+006X8E7mkS95ttyh11ORv2cstTSI5NVRT
BajcN6s6jOI5U0FpooVdPwqpM5hJ1qZ5a20Plu6n3Rvup5uBaX+6X3H7v2G+Qzam
RaZKtVxjIJ3x+St9TI4jQCQgpsXIMHuf9nwzamMIsf5OqlL8cmoNu9VH0mbgOO14
QOSZTe21d/pDXhE/gKFhHVLhclwMEYWdwcME2aqbqMFG9OKXwpacqdhdYudTxv04
rydSWWkcYsuSF2QIMJiNgq5uHtKRajOyXqn7PFcmCvljZrMd15bM/Mws9QZwc9z+
fHtYvnohE2PgxqOarXVOOB/Y8wz0Mmm9g/PTFFp4w4FrWzg/Zvn7X/4RnQ+fjgBX
8Wr6U1OeQbi4Ab5gYsbxvMpdueZvFg1XbquzJxjj7wdRSUGBokD4KM4Z5npzwno+
gAicJhDDyg9WOCyaE7LKVIfHmg1Q78jd0whG4cadrzN6g02IQgcFYQxDShgR0Tvb
ZORLzVX+p3qPhinGuvozViXnIhX+034JiavSh5/uxsPTFAOUHvBgBGy3DzMwE5kE
bbTS5GWff8nZswXyUHoLqwrltHX+tAixedpZAb34hxxNVB+RVEYeCYY8ENZZXZe/
DmPIgrJMHiUKKxXwFt2wEGtqLcN4alIJhaWKjEZyVJiIJQ4l921epITKbi7ZV71z
WQ6DZEyRt2eWd8+PUYocYUedQxNERhy8vg6xq3tkuFqoK9Niz35IzfL1tGe14nEX
Xyq1WFGMhz8hH64TXsYKSdcaCi/dNoMZKGYEqJaPRO74ROejMc0ymGuV+ivgYUcp
zrennghwNmlUFqKgaC/iat/exmXUoQXuj+OHe0cFiX9dWgY+jvnsf27/atr0e8sV
wzJdSji02k7TkmQE4imsNTjUaNnGTrg7pf8cQdgU7VmFuDV1PNpxHWr2SyvD/U4T
B1UzxIJeTQmjqJNRL6Jg3b8zHy6B6kTnBIubUTJcjEta9tMZgJG0XaGP7XiLoL0W
c6KYAmApCXT+1dfu1Tk1E0hkM4axZpOLViCrvf8B5Y6jmd185BHI4RMxBJK4Rq7g
m/6FOokJQhCQFRD96tpo4nV2glhhyC7nuBLxAEaTPbrWvPpu8Mte2NV88hyD7S1d
ZxAmsEab3fENAavuVmrcBF1N0T9QjKNSoN8JtkKqEF1Hjh2834QpnqISC61JAsUp
wNY7KtBcA/P0yiHeM9D8nZj1156LxhbyBBnHBLpuEoFCu79WdS7MPxffsJdnxM6Y
4otesSubvcerN6XklcvEvBrWhsEk1OTFoSsiaKiLQYh0Uib2RWVSKN8gMejrLMuu
4QLYJO8tcj5F7yJOwo5e4uEJV/cd1Kzh4Nss1D3H9LNneVc/GY9RGqmsTgcfck/U
6sYmpH2LRtg6OsI/vnKkXHfM8BLTZ8ysxB+rRs+Zkc5DZ48W1aStLrSaM3V/MGDC
GyJ50epbd8gy1qkk8aVmriahYuJpkbjOywLrtDan8S9rSPOAG0nM2MpatLxw3AHV
J0zVR84ybU5yls3WlK5JHiLX56fV+U+gi6pyKSCPiJXNb8Em12CxK29Oc/YN9nY3
6iqaX3Xd+kk8VfwSHT3AdTigvyKwT/XKrljtzPt3KHfmIUDfuTwA9L3F+XtnkUjW
TO2VYjHU/DhT9ywxGB9AMTPpS/2YTsnYkrnohQozPi2jfw2bI3pZC+kgqN2379/N
rfQ7BLYkEm5O3eQx6O7aeDbgTCySj5B6ROfxXnEG8+cRO3M9sKfIhcWTlznYp5a1
CZztJRNa2GCYJ38iCHIyRSun4eX1Jh9TMeDNKKJFDzDPGUP6aXw8T/j0iWzOQJsx
tyW2D1ocfLdv0faecZk5ozJcicKl1Fn8uxDhhz+eALg+fjJkEaT+jR7FT26zAiuK
+wwIfXv20psDlDoDfiLjVICMbSQe0t7Znh7Vlm3Te52p/qOinyiVUlqYDSgPZr1/
ZVAJNBX3oeA1rANzHy8ERpsattCvWVa3EvfQwxVqLo2bmHG9FRZie0Ci1wqmwykn
lT/y+iAht3KkvwzmhsBogNfWhLgKWsMmO0QbOI7timd4HW1xOEoHP3WulRaSYCD0
05Nl9K5JDE93a9RqVAYxL8ixGhyg5OYMG4kwBhZLbH3Va14Mt5nhK8PDoMj2sXYa
2MMSfS7NzOOgaoNiAKhocJmzO5/cl3OSVvFR96scSlagwwWZqH0f6i3BlTtP1SRQ
YFufsNvthkj+tICA2BVNoba5427oAsKMMmqarD4GA0DtClOaif2C3TZToV30H0SF
xfoQPo4mTiXW5Mb1efve+E5NYIk+xflC1D/QOvaflZ3p2KfeiUleNEFTCW+i1qBg
SLkS8GHkh5wZkGv61gml3Wbc3UUFfDggPHAgEfXk260dbO6a/CJIDrgz3zlYhd35
4hxsrP4xpDwQfvUvoxK976lthOhoqpqWd4JQm+uDckpEL1FXP7pg98j7eOGqNqwt
nsnxq3bMGQ8ug7QrPXMDYOhbFspueTX40H12RLTzZdYFYDtlHHlj2oVKaHQjgGbs
Tp9d0N/VhYbbKTYIajLBKk1lg3s7VHUHi5m7kWybiJq7+TrTJbhaR8uCGwmgjq/d
VGSMABAR9f7FdGQAUmskgV00C0aVO0QWf32o5tNbIj0FkDl7EHvSwxik41XrNioz
9eAbsQY9TJGzSTOrAzRYDT31n3uToaDLfif8A+tmn8MaylkI3DII4xeF/X+qOOPs
V2hD9ia+qas4fG0/fa7yCQ75bMoc1IT6CGqB55d/KvZZl0r0APuOrftCK179LD7n
v5FbfexLS2U6cuW29XkYFsB/Peti99wOr7tbUuOcdbm9ah+/BJdGXxghDhC3Uay3
f6o7mHVC7fg95YYrLmZ/4wDhp+BFN6BlvKOu0TEIKMSSTcSPi4bVNDIVuQAAh7hb
V3cUPXcaEXIGtDMymwgN6hahX8++eB84sIStAMSKbPC64SzGVjPa1fQwxai3vu3/
IOrKXmtcvH64iA46OZrxH65sv3Rk471ztOcRn2YcV6W6u9uBqnzJT2PS68KJJ/QP
9GYzpfukco3eLkTMu4ZR7fPMQRdbPZg4eSDV77kqmms5wj5DJAsZ46uNx1o9YDGO
CoDNMT48u79L42bFs5BwUS8hX7sdVn6XZ2H34zqoUQ+YAYWlkq0ehrYXHe/dATxd
meBq8wZBe2X4hs9GST0kHjV6ab8E4tBM4v9etXeTOXl7wFF0FEq5Ouy9Myqwyi4G
3XGo4PBP60EIktXdjEgTu1nsSCv+BT39xQ6006yB5IYBz1jiV6gwTh9KnFkfWSYL
6J2Hp6vFY82AeGdeNRctX6DqNelW3RQUj0e649pWmWNsqdsMOAfc/9x9Pz2VAL5k
pqd92Y1d2YH4VoH5mKLxK8+KBfRrenUSLkesH7SrYpQf3dHrGmab8vQElvBWIBCV
AKoy3HyJl4Isw/+zvQwyRhEiKX05yJXGBK+wyiMlBeYcQW6LlD19RtvZrrW3kLlF
KjgHjLbPgDZPdMcAtUmCz2TapC2TPSCa8FwpMmwI2mDjnJ8w/fGeMcrWY3tUHNI5
WxoiiDZN/btB/s39uTf6lpTKVw9WOVcbgeWGTVfbV1ameLA1mVfOr5gCjrzYvyl7
/E0CEmethrzc2m3P1brKKdkqMM9MTS5ksluVWc0A1I4HvHlkL5QhscKfpyzW8Cc6
OlSaVpIsfqcuovPMygWsRnmsKhv0LRXnxUKhx8SwTWJMrobJ5FyKCWZXsJ5ted6q
FuJY9EjS/fYh61shEJMlOXa68bMSMSmqamW1NwErO3lIwA/+qzCL16ysxu1PjUCa
Umcv6NdWQV0zbOLNzUS2Ws/Gk7uKCU5vRLCxFqg6Fe2yPAkZrA+ryYsh02qxvZ2k
h1JBtH+j5YQvMZgelWKneOom4VxylPqiUQSM5rE5fsp7Bqe1snIs1OyJBuPNwGLq
JA1ez8DuxefTGql2y84cpzVGD1qU80D5nJZG5DjPvXXDwabj1xRMJOdBZiyc6pj4
Qc6idBJkoeARYTkjv1bzEu5ri0c8BIIV/6dYMfjybhjkbU5BTVL+9/aYbWNsFevU
PaoJIJTOAE/xspaselcIGZIaZUSqZiZnVAXxnu2p43a7ypyDDLc5h89b6r1jCdbW
83KjozsKF9MsMkimgaXIld1LgvJEdR7Wj9hTPAk0pzfZHQ3ISfPhzLuH+vRIBek0
Q5Y7forCTMVI5vlWLVOog78791r8/BXpZZFcGxcv21t/vXbLmCNaACFr+ENPPLms
sQKBXL/zuEYwdGzzCs7o7JgT31Wes/o9qNEQx90LjLIfDRzB1OGHiDpwoQLWExOD
auTXuWJiLAbt4X6kSqaRIu/VS9orsTlY7xZs2WzQc+USqNAUh3BPm29t4HBzGIzv
F5iO/9mI7y3tfd5hSG6vGE5+WCbjAVFvb0EWiC0YL9LeCUh8r+sZY2h4v276WN6T
dZ1WjY7xUi7liRLCtXOmYAjGaac6tZscBG297to/LCfjef/QMcHr7uzUS4gE/pZ0
lbLOLTJrlB6HHTMP3tga6zYZzfOvPFTcJMiRuXVpj/sd9HaSd7QDb+rSDITBelMo
yIVAQEGVk6B/PPXRP1FKwPej7hPX7smU85KHA7KszavDpiUmuPifW31ITLG5SKY2
wzEBTC1nHhL/dBQlSt2y9fxCcOjiuhUr5GenqSCieMlhtTHScgdryZi99mtktkzh
aZOJcMr1YWKLYZ6o8k53qyhpCDHGdaYHprBTU4TNxBjgBt2AzkXqnHyzTSMyWjsI
ENCKjVy4s5wljvszQKfSovPR4jfL1gpIwEED+htsKqL1u8s5Dp+8crsYGMUh8zmc
jPh40LsHvU7w6ftM0Eo5cVrogkF67c+haxIDWBZHW0QnJ+fqyVZ5IH26XMfZNtps
/zeEGaWFaRWVoNFSTzjQesUKtMX+A1osONsQmTynbWAFhQt9rOYzNa4ifP0KkFIK
KIJ4MzlyAJIte9SKOUbMIKBfjYxAolwqFHUFM12PjwfCMdrNZOv8chihJmVcX4St
ErYK7+7SfU9FiPRgB7jNbqIv5y/LJgCgz2hVtGiVUzdHapz4dBFFSU68/Kw/7ERc
faZ1AVo5N26Wrl/IFFeviUSsTerM6T9wKedHyucDyj6k+FcoMYcIg8rCMJU+GGh/
VKXGv0hmoX7H6KyJSMP7iTg0DmtjAzbhgNVbro8ApUnZW3I9Itk7/CPq9KI+9CNB
p6GSpSveLc/mXhvayy+KvIDp8uzJ29tURieUYevYvbLdi3bkAuwWexnCAQwdXzRX
CcfSEZ3122uKL+vmA334C30deFz34a0N7YGe6hy8ej1bbkmpWdg/W85hPKSqbH3z
pWXEI8xpOK3cTRoE6wIE4F/FnMZqxK5hGUg/pJHDhjJ3oxZJYxLrzAzOvc7c1Ji5
8vDJ4Shc/NO8h9kiNnc3Z2jRwv1mMWqXwanalfq/kkZKXlJ1aMjxzv/44ZqKoKXl
gBZZekmt1F+AN8dYP+aSJISmVq55n7Qfgiui81XN+8fqsXN0/xjZ4r8IHJ4KgO2x
MZTJWXV7CykgqOS5Y7rB3vMektUUl+ydmj4k+klb3acTUH2vIUjRW+2mwLoaBIOe
9hm2o9hUKcZqhdD1oyRiP5TFd4su3OVJVJ+NtHu4IbOI02l02qDQu8BRZl2iy743
zDOaSWqnyUpuEfL32Qsm4VxBbM4bEOqiX0UBfcYaEMVZ4bmC9N6k9Ux6dQUZHAHi
92wMrA1grXqy5NymCqcZaJS5VpGAiJsw9LLuE90bblPMAypTRRTBr6Ns9cDi9Kg3
ed1+17WAEYmB1XzkZp7DPa6XGKO7APGzGZdBNwb60Rj3Fx+59oc+izeKcFpUmLtd
IQQEud8lslSaZR60iimD6yKNAx1vw6LtBpRtOFvdrAmfMQrPuwyaPiWSI3UCngoY
m00Tx+XksbU6nDZMHortVdYwoV2xUwGcoIxpCT0sZ9NPRE2KZEggS9ubWsVjzyAq
pKVjlG5Au1lLWkMSV2DXqorR2GXYx2KxbRw2A9/IEvCwwlfHuZi/g0s1pgg+QawM
btg5mqZsWA17JlicWGNrZplYgpgwhd5KhZvZb3QyqtiNaYkEv9LhuGthtgu9RsNa
SbhMVBmZG4AIrQOOVxd40klzuZEJp2gHOFv3abWssTz03Pk8ljYjwXXzIWYlBWfx
guKHBzjKp2wKRXNdlrn/aL6zf8DtBiROiiAxREPNb1rcc2Wf8+9lqhmXFppZ6DKM
8bffRyTdbnQUyEDsGVPWxl6i8znGQPiUwOXkkQ++YkSuhgWc6zQ9lAi3pAlkOiJV
vlB4k71J2pfBI83Njuw9PhmTNkogv1EDGk7Q6PChI3TaXpYaqCp4O2BB0s7Z8us0
59bp8u/yaSYSGNf+QfieNR1Tg6B3hz2O7jazfuMesipstXSfq/TKN9iV9hFrpMKU
DYuKpuy3hYtESGfkeJKjMejMcqLsHERTaTlOIGISB6BB/PuLGhiUE+FlBqa0mS0e
E4gECmE18l0sm7oZNeZyQWQuKk3EDUgI0mWlkhpFkzA4jNIryz/0rR5e8I+akEfT
Pk0p/VmjAY86YuyB5YiPKA3twiLn+9orXU7qSCT9PRiybHTY9FaT8taBgkxWUkeN
RT3e7u8nAFMEnqFaDnTI0eBdzjn8g+4rA5ZgVz/zg5a4cgmeVK2AM1ODD+J43P9s
BNuKZ0WJjIOLolKFY452i6DM2nig7sbQ2C+T4Ssn38eR3AaXJaWflyFcSwVAWeZY
bJwOckOzvUA1VBZkcynDhyF8VMrx0iXD8gTvKetkPT79T0+U0mHI3tYUIuOfc47W
M6SF9bf8Wa7y7GAUoUxpxamjdZBmuyctB5bk9pQ2DzG7He67GAyudtnBYTI17Akq
AyZPvUvFzHfL4dhum9JSbuVHlrQJMj0Y1ZEM4FTd9VtrZn0Wy0ldLhPAtDJLvFWL
/EqTCv3fFJSCivp/HvnwLgfkZGMRRiGCFYaMmKRnGWj2wI/SpsxlzkJBTwpPlA44
6wEiN014w4XbD+3APHnH85A2Q7uA79/NyJ2T/vi9QmyAJ07TzBZH1P1w3PwLtMm0
IY/H+ZTxpQj78io8Y/kruhwDu3KmHqivZuoM6N5Ohp3rPD2hwRIs73vuYPXhkdn0
xQa+hND5LgdjV2cdBrPGujL5KrNSntQ8emCh7+cebfbJfgAdj1SJKMRYw5/qXpf7
gaFvU1Fqsq44JwylM/mZT61/ocSe++ud7FNOiPY1IgGq9kNQWS4iVdvYF55a0K63
H9CImPlMrnfVlNRXyahptDp4LCs2DguFokbUYof/+kf5c27uXcHKMG6S200BZmkO
kwrxPDqzRptYQOc2uzhXMHf1SHiqA8LnyyXp6Zh3a938ySTBi1DdRoPDEILCXFbv
QY88kaPf7xN3TTmQNg2hYHiEZ6yZBRt2t7Z1IjH702tgzIs19Z/qDRI+XiPVB01t
FuDbbhf3D6hihaBlYqGCyX+JsjUNhpIbqp8YTEZvzhpFRsvSxk9zqmkOeeZ5c2gv
A8htp3f3NVFoWEX1x6E4KW1c8+JxfmfBicoz8Ga1jMgkJvCsSTT54xPEjV2V7XRi
N3FYz/07/K6IRbn9T/YaWkanCAmnoItUV2rA1DwgmyEMrQVYmaDCZ2zM2F1HgVWg
w3OoBvseGz8f1R4B4u+aS1ZcCBmlt2hjk/cllO2ZLwcEZYfzhxQkg2ceY3shnHrV
zGt75VRPGZmvG6VAJgmG+OfG1WTU3ASH+GiYzqMomR/MzDEMNN5+4P3Q1o2d1917
jMJBi9yQdgCGOnEcLLuNJJ+X5kEJRK2SgKeBJxo/PGYWmXA3YvtwgujnR8g1rNJE
rZnZNkZL1v+u7eZQ9/fEzWHFeX69V94cUemThht88NV8NlNzkS0aWuZVuZjtbs1v
3WUAwbRKvAJ7flaVtZ0vY5yYnPgnuVt91fgkpVczH0lB5r7iPPmtK0uHZWuQJuS+
STAcu8XO0WuuJGz4wKdAvClJTsvc/Mk06vAuQtUqH7ck96kUtNZ5COuMpHBk4wcp
yNq57G1BlUS21vctWxfH6NsqP3Q7DsSziZjbtE/0FJoysjBYIip9loJIJfDpEpoC
kPGtfv8e7WY9b63uEjulPUFLRsc1V9GxiMvqVqP6+cNZXoJAxP0mH4IXlLcGNMee
aXEg18dwRqO4iZFJncKQa91uRH0hMiMaqcxg+FXWmdBYaNZ/xeCRYgW2i6ZitrgY
bSFDylKXoQJaghTyMAbp5qKPn5vn6MvsYZkjfXR0AJgYwpGSj3Lp2b9hqeVmKK3X
qrDv0LAV6OBw15fTfknMCyWUMhq3kVW0kebpL+pB/3jHKRKDmvq8NXv8713rA/+b
cwota8cVqpi4Ha80THOm72BD/n9gZTqXS5cDsTi8GhYqN38OXHqlHxurXjXZhpFh
ke/Jlhr0wAk62kA2zdAEidDz5+hs2R7YDMOyvGvt6KOVF+AXdwv3nN453gL/HNlX
/AajCq/rKH4sXpw2s3836I6v922+PWU4qi5SVThphd2g476Mek0d/kksaR2fn+jY
0EOZRzxxl6zI2x1P3Y7tl2i8wZ0qLkx0mRTBz9w20qhlP2wnOaLrHXeF53RWLaye
g6X3UE4UoQjjqz4gIOX0hQRiE9lWKm4hvzBdRP+mJHJTTfpVzipPG1ozq2LLw1T+
fLwgZ9MF1grT36kS6B012T7dFHC+iPl8le7Cwdpx/cKnQy2U8QzInCZcu95Hb9qI
qydQQPYmp6TcKDEY1zJTFQzNVd1z7kGpjAJClROyrTNAGeySSlCerTEXzxncww9K
oN3Qz4SEl8gj/yI5Wz6XvpdU/TozEL91BHr4V74JGDLcm9lzlei28EeGu8rraBzr
jK+JAd585bTsK8XAHtoj9lKqyXxqHXC08Am32wdLFC4A/rSgXL4fDw2T02H+sRKH
0ogfmMyrsnDVlUa01hR0kItHl0OUXAR1/CdyxbcRD8yhMD2Os7CfW/JQIlA20E+U
kQTQ1uq4VbdZthxPxcYUIVGQ+tP/5D+ZzcVqrJMTWBK3JNYT0wzs8XW64lPJv+Wf
j93ED2ktAKKWdX0ZwgJ6OH3etBiKlxaW1IYmxJuLfGkbVfPQS6A6yeskI7pDJQRg
vsY6GDcpkmeo0LmqjCBWCyBreJgiEZx6LZkY3v9HKn/6tuZTPi/LXbidoFhWtkUP
8vdCUw86LKRWeJlsTtvqQToK3gryPEEBxAYECNePc7Gfu4X1+NoR7d6s6fD1K1gW
rJ9PDDbBdTLj45+RpBcUHzXAKRZ9+/bcGT2+dhWYvPqih4fqKCy3ZvDAddEyjPzV
E9ybKgJeYOYAUSP+D0V0D57RXpR3FYywtPDgY92zBbOR8wjvpufvL2gicpVtlnPr
dhc7bnIZpvKY2yxcETWIx2DRH+UizEWCx30Z92L9Ha/HniXREtQK9WVP7WRs7ls0
doe+qIH1EamL8TvRaeRhfACqFarATM4zxpm23xnki5zN2vDh4XQdHveXBG9Cs92S
kxFrn8IOkbx6zoptL2uc882H5y19MkcelHrQ6og+MSCdEpxMekeIF5hEXdOP11Ai
EX8lUDPLaakNccz+YWdI64tMD7bk2tbYCoMSxGVOSXCtXeBHHnBghzHJCCfEPXxw
FKSSIEmo8wzorSay4cej9UNu5Kchq5mIMh9Rf46rzmNkOlpvtKkIJuh6gegIPVXE
ovUxXkiPtp/CboYxI5BVPLhWwQZqtw1vtaEbzpMe+/bQyDjy8M9g1kpPtaTvtniR
HwshACqpZODQRE7zshOQGVSBqCgcW/4JZ1c1QibTq9iUQ2mX2hLCBB/wPgzhP5mV
RSlQRydlZdmxATK3azI3kYw0J/C2X30/yYyMmsCVB3caVWAZw/wJAfLjPPaWMOaM
/vQ9NAeuhJJHTBOyrP/lHd+hWojnP+xj83QfMgL0YlWHNJq3sAj9nNIy1sdPE1WH
X4AMsi4HZSM7ldIROj1CWdfVwXZJUmeO0Qy3y0p4+8SjED+LfDkIdwzqUnEQO5VE
z6yIJJ4m3r+YG0Y3y3Vpio4l1A47AaaHcN8F+yEWkwkS1CqhscTqBAfgFk9m2ZGk
rwYZ9OjmY2KvDY4u9uNCTXhAVLe2DhBJmudrBrJTIiiHPtHGypTWgOP0cuizVEaN
Wx89nIVUrpBA2mS1vByedKEov7aOfjQx6UiPRRF6xTT3F/AQMoG9DIdYjjADP0xQ
Smdok2AFRibsj4Z1O8AI6LvLAPyXGxS1sQGmYOXXihiE+eRhFTU8/NkQHOTvAkLP
nrv4YGlwDDZpeKjH2bVNl99S+LthHYr6lQsNt8pynd6emf4Rw4QR9C17unfhrCkI
nFLsEpNnifhrd5gM4ju+QhmjhvStKlP/IfJyeUOOYOter2xw2lI+visBa32bJWYt
4r32yhI3yOlIKPZkmI8qAYq7jjtq7S8XnpzqoBrQnCMMrKZr876bwkJuhLfioKUF
LUYHuzClGtV1bHgicdZ87zFyjJiARAEfO1MZnjT9ntPbKDZPC3GaYYiL/V7OOxiQ
TyK6hiViKfVzyQZf1rlUDX5MU/T6Iaa9aoTiU39jS28bVfZxb/73aP1vtOkqseSC
f6DMeH6w742UJcPAuLqgwQ1ttdwzU57a6Lv7phwiDfmig2zp/5us10q1+xN/nyZU
Cjn2qzcwJItmJwr4nuFkVt0vVzVm9PNik+kvFZWK14A2F5UVNFh8YtrreQF58ycB
Yb3KTP6zFeo1tNETXtlvv4G6gntrqoE/WCSdelUBx4QibNEikKXxCc7QKo4AAndD
3BjRMBPsIfU3XOuOcFTxCGngwoYGoIZrJLnkyhnSZGdojpcjCq1AhPP1jArrWq+w
6Q416fNWgOMVkKhsPLGEJ42Y0+njFE2m1yW93wiDCJbY1Bxw0GMmw1zq2KPzonEA
RxRPkV+VJbodU9FqW7uXN+4p7kIMbJQ6G/jbaOGZcvEnGMHyhs2Ns0z9dR7e4MzW
/DYTrfb2/ezi9TNUvyRGd/RY6Y2G122OiU5vMSFx9JMV8jz4pHweZMyXybIzHK9U
tS4QD78rhw3q11C73Yg5lidJS8kjZ5KfIxqsIrWnUovbZZ0ZM5MzgW/91Q8mwAne
rZIZzFMOoq6JEVpJ16r2lVcm62i1tW5oti65LXTh0sSsZKl+F7Vg6/M9bjlP+qD9
qX6Le5oqmo/ljXdvsT6OxuMx4wL3Bn5U7j7OCUe5Yy8Sk52LbT0hBlV3rE5/jZgD
6mY0d+QbDuBhb2Rg+UdWxTkxhIB38m9R/aMoQQZpCauA8GLQkGPCNK10KL/O9uF6
ozsdWV1jU9iTccmLKN8tHxRMKaHn49YbYM7LL0/r8WXQ2RjF/YVRmcQVmdtt81iO
VX7RY82LGnJWQpKmBzOQe6h38bBgxqWYuNFo/YWZm0OBsRKdXHWczdIJdWKnZ2aZ
fA4l44Y40Qi+xuWcNfkbZQUrHb8HVdUU9RRB8vfmXOI09zCK2fC1L8uWFgpEM3su
jFW2HXADYtNWNvgj+L3D7pvuqgxXGfWwrIg23k4KD+cCApok24aGlaIPFivAem/h
BVwOExqUhJ68hWj5ki2hEe2SbKVlXctmowhC6RFyWJ6BNpY69dEkUXzGr/LYcqkI
jqQ37nPXsUBH1BGHOvMDmhp8f8G1LU5ev4Ju4hm7DWY8K4BDhqretPepe+7UMvjT
hk3UNT/tQi1y5hoRsWv3qo42e7GJikx4Jmi+kAxy6kYd5h5fZ48gQ/8A/ztz4Tvh
7cAi7avKLI/9EiULSUSKQkzjVaSYR1MeTKRxwbc6EvWibKUP8Bcobnwud0dLfJQb
nZvnhUaPG1xYEmoWMLKsxBwMX1ixKwVLlCmil9vm9FKn5vO0FqmXXmZJ3JQFgn/U
JxOmE0zanMXne+eRWxmGfKHTUj6JdJAaaK/KBEen9sqNBKznIFMT4KC/YF+lAo/U
vlWk+cLfF09/DGobOGaGsivbuWP/+Zgl0dNyH0NFQT6UP1enqvbd4MY3UNKMrqIW
5s93lVSxmXYmZJwm8mFc9a7y/Iv5YM1YmbIkC1HTbg66TMQAlMtQ05ckySRkmB3c
nvLMsrAMcvow2Wg2Zto5+v2qB6YiAMfZoKZhSyGedJJ9j+DMKPWHxt0XOC55csoL
2gVOokuORp8WwsPhjpkOTW0YWtkVNUI/hggpLDP5zWYy2GPCYDCwyurzMbGusnFN
auYjcQStGFcM0IfJrMUBDYAeGCp/ynumAzuSFdUO3tTJnMqbT2F1g6ABpcEewVQ6
SmE9qz6VW7lJa9VCEmQCoAvde9hdFVd2ta1w4a9JVeTIwmqzh9hQN0MgxSE8NGBR
B4TDqchuZCsP3rXXLtAb938YUAsOJPfEdBKktpoGR+PT+gUdCZ1qK7vDuP6w9TVd
TvE0FYZixBMeiSoraupwQ4FKmYrw4e+HNZ8zFmoo9ZzCRtG0Fkk11bXengIpzH4T
juoVuzTCnfGLIqBFs1rQyT468sQ2N9CiJmMOdhBRW+3nCNOxMThHyd2VJZV/KlTD
awCsUVpWdoTcuV2tWnSnXGpO311J/tQZwTt5oBKk3kk/CgLEF71VsEXlx8/gTbda
IyrMdKeJJtKHPgIuoXc1zWcDmy/hsy8UKGyjYO2ZFjLAuKvGJPlcjJCIrccUs8En
MWYHVU2VwtTrX9OrXvxXUrV9/jlLb7Gqi0ktaF5MQqTroB20H+ml68/vpBs9s81w
jD9rB99KpAwTkLM0nNGwmG03vfpGpptl0x+9kYpJQIufH/tkEGNKqbNP7u2IGhHb
vp5igJoVSCkkNR7bDb8jLiytmKFlkPcwv7eoZfaj9q3a5nuPry5Td7E8wHDvHakc
gc88pSzcibOqX+6YrW5MNkk5GVZ8HDmDK8LnS8Q7gTahCaDsLh+QlBvEg0MTrvEz
weKN4E2LiQQGNGKYQG2nJPQpJHkZ07qEm10e+YRD7pR4qQhj1g9ZJ0hQloEiA8eo
fjtzWO8UA+Kv/lnfovQQJk2cnI/VRuhZTsbITS/aV4HdT0XOX8qYX+fjbZSUDxGm
jI4s4vjhbNAPLvmqQVCdHQpKqCbTYWTDJGgtLaTI31/EM+LSjaGNiV/GGqNX6eAr
rfvlQyyiTMUiv7KyjNZN4Xq67AQPpmF3BEcnIN/Cwc1oU6BkQihsVPpiWlhqUJ7X
a8PI5+OB5hOyXkRrHW8p53WW20O0BGVqnmGiu0F6a2kd5ygcFaKdR/Yd9Sq+2wms
PjJdaBN/08xc0hy7cdAR77qfTCwUVBkSWGaxPdmu33i41Xw9/4VMB9FC42Yb5c97
o9dcvU4UUwfaocry/sWFUVb+jOKiR8sdSMiwG4sBpsbred0fGMCXASF1aMyh4qdf
ZtQfJMri8LQfnPTrJxvTrdgdzFe1/RZPltavJDVGmw8c4RJij8UE/hoUATV8ZvBt
XK4erZtd+NS+BmqbaArjE2nI59Kc9AIqyJkocgUHAnnDXaTlWuVS20OnQ5MmQW1R
pEF3pQIOtigFoSrwulflhTyANpRj93SRRuUyMC92wJ95BTN9GgdNSetwqyJSNaYD
KBWJa8KRZGc1uyW8c7wXmYVGk9AZcsF/01Xm5nLoCcdFHOdALPhMZVo0R79M6ybn
7ts9G5asi7W/c/vM4QZtHr3VwQdbHL18X1zF2aCm48hRhPlb8gAhxKn+XkGSo93o
hlpUSVPsmu2FV2HqYWYU1kwjEcYdkwgkkSe37W/fNqAEfI3lOCjc2jGnb4P54cBW
TUMlNUrU8oAKkwp510LGdQxNZISpLx7snoWllfHG5GxWfj1hbhf58qNBeQlfXutC
TngBqx0wqgG89waDHnNHZ6xZ3j6YcpAT8CYWY/yIOixDgCfsbBdIA6Rnc9dKOag3
xir03IRt6ShFNko9+LESzyKg2/TStNXHL8mqXh19OQ/diep6T58Mnp7X+8n11kvD
7wtCZiKawXUnCzif4O9gM8pVNcVrUZDnCt211EqoxKXlK/5CQeSErF5OC49yQMIu
dDqNd3zohE/wR7LAFFM7o3VYe/dPMP1fo/aeezgVjkUfj7mTAh1pqJv8cacy62vA
N7ykyLFSU8hGyJxbLEwqV8poB5Ci34UvKwibRSGzKasNoP95ywWtdvcAPCplaMd7
FQXZ+W9v3ScMFWJ9pdQtRQGxG8XDudLZhAFYqz2utBpXH4uypr2FhNMjGQJWhkjZ
z36SSraBi73KOWkvebW3bZtBGzmNKSMnSovXf+13TAvfVDVMFXqYAE7rMc9XqjRe
gtnTq/51N889c5pQOoUYfhBFxOZSv7MRY+NiB4JH8IPMC97HuJByFq7QLa5Z4cUJ
PgVUT7a8ClMld81O6gwQOix1LsXWsjVfL0ulCZv8f1FXHqaEYIKEeGwbG6woK96C
GNO4mtnvGN0xG+cgO8D+rgRhSol6rW1YJY9CVEzl0Y7h6dKqStIHGDmo8cv84429
bSWOkvQ791aTHJEuGmgkknzrZUrGVhsG237A27A6V+sSQOnYZzTjQ0fK9OaOrXwy
cYu02BB782If4UK5J96Ivyt6KDsRs92Rt2AnkfZ3aOvY4YyH2uXe0ZWPaaYCzNIs
TmbuJdtfg5puawPzdwcY9bjdwMrJnNY/gPlmT1NW3mCRjp/vIipMOdan9pM9WFdf
yHV/UovRngnDHCDtAf8qSBV7vmRODxE7VI7VIyS/RZH2Kxp6O2kri0mA/aZJQGdL
r4JqGX1aRh6gXPvYqzWjqbgHPydgYbrprnOSjWoyg213elmNT317BbrJ7Xz3doHX
EH5trpal0KBxixGlBSxDhx7kcSpgb0GDuMSsuV1kPeB7eEuCCKREd/3+RFlb1YsZ
FBykAX1dCTSMFU2d4Wev+KZo8B3BQjGfGdZoK6ac+DeK87kNoNckhh+MFyX72R0Y
yDwtSwm+jm0Yjy55agrGuPaTIM6Pbi4BJDbNJlEEhe/mk7ejmtq4YLR/25wbtOuH
ON1o+ghHaq60TN7LR2xRAh8MHJeq3uaBD0dxOBn3DKMZTOg7d4m8lF1OGSHcnr7T
hkGHnpnfDO5czuvxKkSrmzLKciBEeY1ldfJkKzq/L5+r00q73BIhUvUxiX91H3Pc
/3WhvpocdFu8yZ0INAFFR48sWKvr2EckPHx/Hw/dUuOL9TuKUaaqfd3IhAG8bS3i
/ynPYvGOj7gnbhNQHBkic1LjrjDAKESJGgmSXufd5G+QQAwLfa/L/nphJYoGVpUm
9dW8fiooLEcxQbUF2Bg7rd6ERf4EgkNrly7jD8xMfd0loznG40PPYLWg4FDQcQ82
E/jr5c8MH1jhGVRn9jZYjMpssZcRgZSIwNr30sm966dD99bztwXV7acC6qbEdwjO
SoSiOJ6DQg2E/9KQWwtF/KNxANjmXA7gIyr0IJbn8Z3uZ81hvj55IwcfKUzwTkKs
RMaYpV13X0Eupz4Mc9E0eeIUsCI7ZwAhyVkt3N00MqMdVZsi2oaZ+nfXTYAcJaiN
FxAz3UQL/E7gNdZY89oE0fROLTjHjbtb0csQPFe/lc5sA6Jc4npoJQ21xPYKY7e2
gu9LCbFmrjTuLehXb39VEQVlVeH43FqNuulzIrMr1SDg89SQZX4F22QwAIBMJdVN
c2FqYThi/W2nd3l2ttWWAh7kafIzIZ4eE/aXqZzAyxQHH0cmdD0WGC1wiNNU5IS9
CSbjxWPWfOzrAeaZPJYpsa8B2lzNtkCGvMS7byeI4UX5ZPjOjbe9qnDiTAmFTypK
vn58qpgZZoHHnEi0wEGiDdYU7gAF2WrCvz9Xlzpaw4vAQCXZTLEPnrfcRB4UcUX3
5/iMPExi5Xh12YE6KG8WtsuxK2qfike9iv2bRsmyCVfCoXIabmZq65SZb9dMsQL/
EzSn6AIwnWa0VUlcvy3KNUmmhk598OL8Zq5fUVEgykuIcjl9ch7pxEu7/g12fPhs
jdJAi2joqXJx9FDJ2IV1cYX5JuLeheZkrm/8yHelL2Erw9kEJ4+sWzi3JYfSSzKP
Grcqmch6/yoeVQ6ncCoOpSm5HCynwIsv3jDLrOvaXfzVpG/IPaOPfHk8jmzm6wgN
mn7NJabCnsXm4LnyMGwo5Dem5AP9npNmQsv6e3b/8s71v+Nn8BT0O8Rx4nKK0KWm
GZ83NAv1l8QocZrQLV9FFmV2xEPW3cMZpUjgus9MhwkydLdubs+IJOLZHbds9tvJ
aUSUG2CnI+d7towZ31VxvONmttCufsq6drwp2NyNN3c04iUirulyZDDBC7wTHAUN
xbsYNKc8qTyfoZLSZzAlj9RgFLoqTpGVQNIRuLKRo+aWbUwbnrhiPKH51tftnmQp
HOHZvYMfMj3O7KyCRqUFoaB4NJ+3FFkprUdlPufu9lepp6qnNSBHjjC35NBGYEYo
lgmj1xIJOG4oKJoPxHdmy3ZMDdI1Fqz0JonXUDiFLXqX0JD4eCq/WPk/9gE/PSGh
GebkutxrzWf4Iy4oJV2FQMQTivYKndIwCpzz+mtgRl3OhuEiw/xUEtbIun/2QnAm
KVaMytWJIV7F/WKfx3piWiZkp4CGVf1Wg7MDRMEp3vTWhRfVG+DK9Di08mBErms5
ClIFHqds4daWScV5JqpVESoFvZIyHpID7QLf0tk/W0kXAcre4zMAgHiQlXd1A/Z5
pHqqXzA4G1XUEOxbABQl/wdS5C72Um+zh9jNekuFKCglMGc2sU3ExUTl1/BhVoKs
zREUrYTM72Ea9Py1+Rp+DH96sGmk0d/p0eejTPmUIzyuI8FR5dVjdTSAFzDqLYEZ
lnWw+rOCfH+lQo2EPQ4uVTjNDud6SE8QeTSowvdfs3XGIOXwSqoZeySzKe4UpcJO
gRCKFM7Byr8fMbc+lHFqX7Sfli7+b5bNZWGs1cK3Mfyy4zgFaID3+X4Mly5aMXXq
yvqyPRFxEq+QU7BnpDCMKAuxBLnH5wzoUl6fr1MWNFuC+OkZFAxZL64gr+wrTd6e
xwm6KxCFHgzon948RxW4pSMi29ZX3LB/4B1+JBTC/pYY8SR0fNLSe/7layxuzlWa
3XFB3q8G5p+S730zIN1WYQykrkIy/CWOmLBBZ66JUGfqVUe9Qigpq1ETxKUtcCLm
n1sfdsKXIq4zBpPCRZnPd64GlhryVJOrusCTxKGeqADfkzyuLohkjW6k7WIQxiN6
mamQSFHgJSbbhu0xZdFF4/EEYKxbwI9axErpFvm/FzuCPeAq8NFgL7Zc23y1Na5f
N9DyNHDEUWOhyGqV/oBLmkTrxhKkfcOIEYAGNMZBeQB+7xBJGULb9ZrtCZ6BPKlN
aHQxQRtww+561tLnuq590DyhJ5QC/Y8uYwM2YvXNfMPJSxfAv3LfDHEyNUG/NnQB
7TScvl1XSBPUgekdZXXhXX0aQ3sA4Nljm1WcV8aGKee3OFj7XUZXheKhVBk7YURc
QRPxSnGsK1fNOD2Ui/NWhLqaGJKOpz1N0Vhq1vajedwXCqhlvW3FwEm4UDv2Ni9N
Fp2gZ36KHwmTn8tj8fMWoa0vfscAuXe0wDIwgrijDuS/s0G7IncNeiwtApeLGULp
Nse+Jr164//ILAyEmBRxIUTRSHOv9HpBha+DECsjp61DWuU8qM+qjSOP7QCdlbJx
JEbynAFngs3dkbg3eBlXBnT2Hs03reqkt5S9Ul53nQIjlbc3+9uZcK+45Ne+n60s
nCIcScyZzWoE8gzPcnZqDMTB3XK+TCn9EOqic5vK5TLXWb7T5JPSy/8wNXz01FPB
Dqf+sP00pAU2Q0yl7j3S5pu8pPL+qpSWN9ICVT/vDutS3m+rJNY3ojb8UdDjizdD
w04YENGtaaVokICQ6f9Nvq6n/h7lWJxLiROmvAZcJGHKR860jSf5FiG3SdQouXUG
RGmIm2zTQy9CT+nvv2JmqZweCt68Yz+dtSEblImAcuKZOBBVioIV8WDnVCj2lCaH
0HaZfmiJ3XXebKpNGLIV2IVYWRUaeWJXxSmYthQCc+WQzeS0dWtzwRVhUebkjiKB
fQu+waMh1gtu+/ecBrQU8RaZiBf7TBVi9JBCN7nrCphDYgVaXE0uPExbO/IFzwUw
yUV35qFfGbRNIGx59sLjOxzNaZgDd/FGDe4R1T4yUP0cXOmGykBXxhOo0JiYR53P
Q5CwDljOOdpyrJw+ZDP1i3/I9MNozRLiY0hLgo23ZbqILvHHJykNIlxdyMNwWVAX
cqBDUtVGb4GbT74V/04KaapBn600fOffSor3oCY4ua9DpeaYnBYdY/qHh6l1pcnO
KI4Yaeg1nMgS4qogk0yYshlFZZ4WDmg/XhtNECRrulZvEH40BxyGn8XRaIXKKYKr
iNWk/O+RRay+Kv6stO+1nMSaW5/g4Oit1cosnv8FTWyUMHDqec4HOOGtAOy/H7Cj
tNfN7C7TssC7rqx7+vBZTx1frx0fZ/flsE6tU2ZQjRb2zOWMB1bZmdQthRXtmb9P
ogplh1jbDkuajb4kH2jcNgasD2zlpFlFv4wtS5XeVFMzPh+ZGrkMD9fLL4lQn1re
F+H2GcY180yoNudyUoZZDJXXlgIBM8lQzMxfnDoYhls6OuatMdKZzwlYejMqQdNU
si+bVy9Td30KqoEFvasO+PIwsyCx0sYbRY2TRpAPIm5RtaXp0n7JBLdOycj1spXL
D2fYDTcxxlQQwQs8Do8r+YvGj5e/MhrHuYbpLIuwr7iP5U4NhI+xxLbwUkz0bsy1
R+qdwk+H/0KA/PBH++XuwtlkcWzmm9fLaEWn7Wga2nQ9q+ri5SQQQGLDv7xJJWlk
hoZsI0Vqo8xSeeTH3HKD3WD4ka/QnhIvN7lRPm0HBjtimVZ3LV1ybO1H/D64rH7R
/tLp4OZQsCANPaY3Vt8BrmbjLdkbsmkSL/BYIaLvu7/XhgrT5lAxWczjZN83TojT
uvBKN2SsxhQ7iVv4pCIUmtz2fy1E5hrQSYxIsKYAQb9jFY8yOpWys0AbumV+Zn33
oD+fGrT4glWIZq1RGqLsO5vZGpnm3ru/RZ/ZSrHFc0iIZKfdZt8hgryfSFnJWJT2
1xXhIbOVGZTUJpl8VJCfiG659YqSLGEP6UArJ8NubnL9qUdqx0M4BNBNufVpireb
eNLXtsLzRN+hJ7MnPxYR7Qq8XDZjSHuof4wpoaKP0z4vZkPD+4upehcBGbIuxKV+
J+PniSMCUKGT7a5BGDC+NkHGG6mpagQ3hSXj5mUiJ7KnfKGcZmq8F5pa9Xx0f5fz
aQ/EEVYdmX5dH8843IQK8oSkkXbFAcJkI05klYpH761MA7XtX0sXhZjGdRLucSCS
J1H3Fnr4xytX+KavWdnwf6ybfdiOwQFn7EWouy6EVB7HYbShgzoSDsVwUMEPrrOT
/05bl/812V2ZsMwPCW3YmXgF3WOWCDSh38VUWeEiwDrc25bQKCq2D3Rw5LoelimT
6xYlJHF+1fvUYwlXvnvVzLzeqR9f0bPc7nc0HDUuLPkmadjgkde1DpfqPYAFrjOw
KIa+gTpJuskGPCxhEr6tWHyM7k4bUdB2bU25cmXDr2avBrplrrg6Jb/SPXLLLed+
60J/yvYX4Qg7vy07xPNrZjerfDpAKuzmPVKNnlAjTEauBaNT65sMxewygZ0iHg0Z
JM1lCCptrhpjxKDKEFHcnfZs3chqPYg5bEyXy5ubRHMPR4Qfq03nGoUd1B3cZF7A
bWCuSfMQZ1BzRAK0fNW5jZCYRlGAn+nueAgm5cEFf7833K0mgk9cahApooYw7jN+
ICEIlXYeWCqNHMn+gzFpEZTBGJWk8luYzrVJADrcpH1lGunsg4pmtG0pqE6ZEZBp
ClKQ1dn1mMGhWD3TOe8NWASuCl+TWf7t9saCiNDLj77g/oT3zL7byjp2PwIwnnCM
szVOtfGO+gy/1LXkHl6GpKlHx5uCrio5Z9VSKrGDh6WIcP03nAG7QRn4biexHinj
ifKEYd5rukDnOngTA6qpa+w1jDlogtLRckrNAYJBxhBZ/qIgtM1kTrGuKFq/G4jv
zw5diAIoCI348F0fvNZc1eTiKc+qQGJikig6tLy48IhFYzbJFUuZK271BmsvzF3U
h0EkOb++pyq1B/gv5fpe84d291QcB1qZ0TjcxhLRToZuGyVsKQLTyGSSHEvXyia8
L/K/WoQK7lvRHmX06NlWfBLy+p05Of/IQiFNWvvfh13EHnHtnRQqqpPe8d6hCBwc
cMtwnBuLh3tOWduacTc0QxKZHSyzy14nROFy97UzGlqcS58jkYzgM/5UvfBF/ufw
PFlUK1Z4j1ZIM1nS9OxZWtgrSmYrTDAP4Gxm4Mw7Z+VhIH3MdfKqL7rGNHsIGJHB
SVpTAU2fWx5KqLnQxvSeMysoIi8rmKK2qsfaCFDNkzILcZG66vbKj9vH+MMrNTOn
3AoifxANzPlLp1SNEqVoefqQHfPhUny3jJoZuTSWOG2johW5HQdPz3v3VDHtRUS1
ovzLpfX5wasBCn4t8EE/IZNacAGGX14Cz8spgpd9ZWt9n2xQyv/NQbijWdpFyLUL
9J/kEcfm0QY+V3JOaH2eHgcTs2ZrI3jHf/or1ghQwuhOyiP/K/dJsxwrFOBesZPW
KJijnFZ6vfScdW2lroWQ+X4PFK6JPB19Vqu7r/TEIeYQKO/dtDIAobaYqbmap45y
5p+QiJ6bkAzwlmXXROxIuk5LIBfBdxvKAA7OHcTF9bFsBreO8eDG6pVwsZWwKZKm
6rV6BMeuJHX4Osc1R+xuEkpGelSlzHwKsfOKBkaEBl4r0VMW7xlz2+OsA3MxRZiw
gVZpkXhxBxcThV62bDEg/ac5KKO066ElztOIFQWboW1QrDyrEONZWjWBRlctSLHf
CbzN7eGOO9Z1k2C7cvhipnjovSMfILq3tUJ7fU3S5q4CET3hXFL3CkGzvEWIsgEB
H73hfW4cwEFV4P2a5l42WV+kcMOFXMzK01tcVvOI8eGCWpl1goVk2aPKcH1Dzf1U
stW5arX89UPdcB7f4IEPPSUMqhA8xjYt/3wm5M19EX7iubTPxZYD8fN+EqGzOll0
dcxsX9fLkUo1N1DoBky+GLqZVMyVAsm+yHI/oBDZDjHjntdebhD8XtiBZzdX/FkU
4BV0VMIJM4Ekfp4H2CzstbkuwLWobXHxSAnybxb1nNBriIqcRuvFJMSP9S47P7Kw
y5l8G9aB9d82Ayy/YU4+Wx6r50W8EFtk4cE/GsiNXJK62n4PJa2E4FpcLfQ6dVuo
fVsuSalKvk/h5INmzh4bonE0QTO3BwKYOlDW9smCjRvMNasJOVKbyenhXG44cg5N
cj4NTCp3L8KBvwZOjzmHUtgMVA//dit6O18phNj2Wmjxe0Xp/42pkPOr9gccHNmg
NGESKCFsfVk2rAUYLp9KppwASXaJtEdMW+0qmtLKPZROQZtffGll5tO3VFttu7T2
AFF+bx8Wiji92RTQllI90s3MMVL2Yo4PIf/iheXf1AzaNxWDZ5d7jlW827fZozZP
2a/cImipdzuQUL8ZAIWvUgYfqpK1txiuNzZ6KalmysnLorHpo8p+qmtyPLCITvwv
fW1cOTTG1BUy6bc5V6QvroOi4kvqfxBXIQCfpIzxQXEXwn3rjC+ZDgGu8lo9LXDA
znnp3+fRTXo7y9EM3LwGf+twr4+QG4/H/zUkI8cLfoWlhIWKoBnhhdqw6JV0IidF
RhnWe+y11tQ3G66T+9MbbbXw1c8DbC03ADLJAp2MaYEt4FxWXqaNU5XSjLvWqvxk
hzK1CCnKLSUWSIS6hm0o6FZ+NRl81nlpyoJQiWqjV3LJc+ydvE3m/L5K6WiSMtwo
SWkxc+lZF/6T5lONWVsSshu2FurdB6qwKaV8R2FXUzBlwUxrVQkmXUdHCxwlCXBO
V0JXUFqbscQN8EGlgQUiYLTlJ19yUCkE7H2Hcb4q6Xo4imdltvNL5z+Fx4eQMZTB
V7Id5L+nI2Ic1tMTm6HNjM1oa2vkcNY0n3NOz2FT8gzWpe6IbZOJU+/64DAoA1nU
zT+4JJr4pIJGL81YAPNI7GvOdkPmw1RQ1griO+qd6nPAO8IS7IJDsJT4gjOvhrAj
GX7mqC4Q+ANJBGmcalbWhoEA9kHtrrYtY1CVzbHmeOFc6WFQXzERzNmCb0SV3Nb7
px1NLZI34aGM3HrKEcsQF8x/N+Zfrz0x42ky4ifU1Jd4WD/8taVZTbpY3FTQR2y4
pQ11o4T6hUTZBL62LG7D/dWmoOo3ml4yUuVk9v3uMLTfrgJm8wvJBgMZBLwQr0Wi
ywAlOxPLC/5bo6pom0VHawNCfyIDrxyCJNjX+hcD63nc6rov+n6G8MgRI+3ogD2C
MCYMkQSFysnowRY6CJ4HeRbPZeVE58XPgqlBmMv+FdkQONxCxQvFLIwrIuloBnoU
xlXShDsaIhq7LKN2oeMNAyvjVJal9tbfNC+Du5SzmUOiAlkPInVnmdYipcsPyw/j
tk2SpSYX6BaTZE8pM1BXUXkN9+A/l0l+mtC+eqBL1OLKayA8a/8Z5I/KLlZHntuE
bmsieeZ7pfqdsFxyAH8069n5960r4Vu2mBJuVUu0h9t5eWQDFaJCJoyRLdDfwmAE
1r40EKZx20c/GEPboFlSHFqSy71f+2LTuS3XdOBAdZlKxlfB00O+BY33Njh45jtV
8Udalh4RTI6kJlgLMhxPRZl2U3KgnwvViZYAxoU1UwUmX5GrpEOTu7NWM9j/Beft
6htL1OUobG19P+D3I5R1Qiohzx/AY9gW1K1oXhdVyDtailShiWKG3uK3ObSTV9kT
n918swASGU97/DrgvDIcQwRFmNlx2Oj/lMzUuiNeiDG2lyqYKbMBXyQpc3upotNi
S6i/iZ9PaZ9ShI2baQPn3u24h7DclXw67Ggi9BvUGimbVBxZRhI3lI1K6rpy3/U5
SDuh6BEEWILK02S8gx676OCzocqj24xxlWYwU+8XI5J+GxeMhglJlH7Vp/L19rAh
8p0ZSGQHwNdf+DIKg427UJDcSwhWZgMlcY1LKobi9N8U2ajCkgL/T9bcYCLFYvhy
atkEBo0ZE1Y0nYBPl0mxH346huPWb2W+0g1Zb7qL7pj56vWrqSj9ZPpjPqQ8Dh7b
18uTIREUOQ7o0C8ChkHruM4o0kZLkMVHRGcAXDpGkDaNoC/r9Lb4p6mYdA136DJD
hqtwTxsKCkG9PqccXr6amD7uWecct3AtjT3JUV9LSCJXHYBHgWHzNr0UKagCm7Ru
MP8bc7eLDqy3gDpdWCQSjC5nIDQcc9K/9pq51DNAG+kPqqyk4BZlwp76KOAAJUgU
eUk2OPr+E4yAx4hoqLcOGIWWKBCGgVNQHPih+bans9rjBr3Qk44GfpzIXXYaiONS
aqVGeyFVGyxk2B2nor8lLtTvpcKv4uOhIQufE5NEB3vUucI7tMOLT9kXTrpk3s70
rwvBAgu6PuTjZrah2OXTVd8ROgOosg+Q420k+kgpwqZ2hY3CMQB7u8Qtw9/TRm/H
6x/v+hDY4qPdQAP+gUxoztYDlgiP7YJ3GRbmdJDTIlyBK5pluK8iJQhiJya39pPt
PEM4f0ui2/LM+Dll5pyLuG/Ec7LkC7X656MkbYd2dzDngTtfdvT75a9xqcgUzHea
jR+LrQiNq5m1kqseT3t0hUx6lwCEei5Ha+XFK8FIxy3AEOjH/yYvQXZQPft9DB+1
kkuHUpD4Wlnu8ZBxssqyVuNhU5P3f9qmcfqXrEXXG5ekreaxHjZQG3eu3y0nK1UU
qChRgErorgFjhmSocOz5tkGBldttjQGVtF44RqEZHAP4prSxsgYaDBrLdIBgCgXo
Ige+b6FkdN85mRdb99PDqvs1vF6YGVb5naDABaIPmFPm96xpiEdoaSZLttgL6cGn
9E6JgtiNUT/4+aGck0GGAW0OiWIda1ciUBaeTlb5FlZKy9P5fw6vVupxFsG7d4jh
EMUcgQVb8nRQXQNITrKBjy3Cycym6/gi6gdYssIShJHGwxncM2S7JOKY+R79+Pb5
LrTSE04jw4B3wJ2+NoobKrFQU9NVPaoPnsYnEm+2TYpaIyYlVzC8yqf8QvqdaGYw
3YGuVV7BuHwyRRWjy6gMOgAbpVT3rk/E0MAsOD8Y8l+QcPp/6YjSLTfKOOBZZtxm
rkpZkmxAAG794I4eufDV27TOP1vnSgEA3pielnAGcSEK/Eao8StR81gf0oOTqT6S
CcKGPzC6GGUI7Ajm+BB5C5Hf6uVb3KJ5MH1q0M2BhUMEPGIv9rUMJy7x/YjjIWd+
tuy6JniBkdUgCk9uDUiuruggiI3vnEQ6EytNAiwX0UYiKAq3sriOOug/s7koVba7
S3L8sGh8OZX8i84PGn1VWlHVubPNodJRyAMWOW0F6IqnQt8ydZSpPk6iQyb+9q9n
PB99oYX0X/K3hXrwVFJwX9+Ra6D5P9Dy/pjo32KHyuZLConsTET+sD229cTAMwIQ
brPId0U01i+yQAg7q0KafGevrU9v9n86zuoea5ZldYpOi6XSVxi2h4NRv810UGG2
lI9nH8mPtAC/4OucY6ckG6r/fzLS+7qu5+LvzxhJqy8SKLldUA3kYajCisuSMwQV
ggMtVgDviumB5fBkfRoW1wBJwtmBSQhmrFG30sHwns9FXnxDwbgrwRH5yK7FAnfV
OTJaVE/lO1YlOALktB/Kslr8EaytvQt51DA8K03EAHegDaphpZmdv3D03vHvLBA2
/hbNCZ2IFxtHs3ANzvWnGUFv4ySJOwtpoR35+8tX4NBqhQJYVMcELIv3B/Z1NqI2
2sCvlyTdUTjSDMEibGl/XOI+GxEf8f1Ydf8oWOKt/tYMYI8ZbWdMEolF6z7ySMSG
cU5s1yjWvqWr3c66RSvgQOrrjnGU80XyKVi8IcJB9E7uORJamlCtHcfjkzM48/y/
mBD3esf/BeobmeklnfQufKr8Up0kwSR07tb3eKT2RyLfS9oikd9Vo290phITOWKQ
QGU4bgsP35X8bt7TjzITUqObKYIDRjvfdUnd5UUEm2MQBRS/8Ng+l0B6PjrNhE6Y
z0yo7OVtCL0CYkwtQDqdCV/b10TSixbfe3H6RAGibEFc/qJpazNVIewThvqigT4Q
v0AUKblApxOxBHyvVvpm0oOtUB5Fa5DB+HLP8rpNvUGSEHMCRv8hxK67SaJedT5K
AyUeaSjj/i8mn/MRvNritODoUb7IJx7Y097JyYbpP1gp98Yxc893KIVWGwibETRr
rFY2utMjHdGcJAUnwxexstVGmAIrnp7yL40trxDwnyvke07dEvHVTX0OY0eusa2m
enrNH/LsaiVxJ1EbY3WPG9jRZtiuo8sKTSTIzcuwLByKXezypBVhm2p/pO+jj/Gj
kvimAyvEfv4uUpNc3UQ0W0sPYNv5C2Ee1xA0eCjK3911v8Q6tKNfjesYIYIVPwrW
E92qxSmJqqj/4xBO476kQqs/mX+TLdYXKTJlLwrUx/yTn2gp1AcylwI4qL9Ae8mT
uUIbiJb7vF6mpDI0Y9es3S5W/q7P9aHtRZzDjana26HzQAfpeJBCQEIdDl2Lac1w
909khcAffIdppu10TIZNRWXUSzVpsbrIPwpVoGhOhDbCaQcURnIJjB2id8Zhu4hP
EL2zeo0MWAsKyu0yhnWuwLYsJ1d6fEUvlYf5Ydn19D6pMhg7us2tX1AdLTwjcLv5
u9vWpoEUv+7Z4m3iuNG5QRm5fJvt60FybsirMpf0EDcZo/dDICdbl3fQVk4ST2/R
fFV61kvZ2zOBc6aS65bobiLJUbJAsV4tbJbE3jcMgua9dCnL2A+LQBWaxtoQZ0mM
86fvctfWE72Ufcu1rwSJk6zDnxh8L3h5/oX9l4BKP/am4QAurQ9haGbjdDyPWFMT
TGiAKts/XHmTCFnBXs4sd9E1vlKS79CGqTS/qIHUYRicQ8r5NJCSuGq3VdZwV0we
UFpMSAvXzHiHx77XlSblUNkZxh4K73jeFXdDumIbeWhwfDOPvFDJZD98jJQGgBre
JZ1pHX+NjSkE4asi3kKJpBr/iDR6iJyCdkA0uQy7GY2wnN/272lm6bEOEthvk6fM
DxFjfedWjNNO/8iuq6Q8wVtbcSD3zzAoP9pOpmMNXw26oFC+1dFn5IOdpJJXq6Mh
8g7H81lWJfOEkeIvvSk79iZ9teqlqXdW3b6WvL86E7YqqClbmJG7NLivAwPDGK0N
4ZvqgNrTV3GW/qCLXyyNCQAeiiOup17MuNijamjEnwL/f0mBbfBy5S4X06EhJ18g
HLgL+j1TlJG+4a0GSomwCGtgpS+yXu3tHqhzUvFmaZJb28/1dDA9NEW2v7knU+rn
1XAQXlCfg50pyngJ3c0aElhBaOksys4ppIM+DrW9WzhR2Leubs3gIjubSXPb2MRk
U/P7jOeCGIlKqqcFtRajr5CIWq5a6Uo05CXYR1HHtlak86KhzeLSl3+RDuw6Pemr
TUC7gT29l8pVG+e79vIxlRiZPgizoLwNJs7i7MzuT527SLvE1Nz4ezdXZlsqCj+c
zHR8GbkdbaG762Ws1nGZvezdwnTEgZM9NdY+eA0g81u93xydDnXeJe/fNatDOiH8
lGu2OHfOJsZG1tuJ9vrIK6JUvwSYdO026NwK9fHtbIPw8gu9OvU9PSNyzlo2z6nv
vDKLaZJDuqxpd2HplsHVLIon8gbwVJ4qqBNIF3Hdj58uHN7P5ugPKe8maqTf97Hr
gUBosVuqw62HefWBMxpSFHnXrXH9HAJBunXPCla5gESSL2+FpwRqkj1y7EzmZRBQ
Dd5+G6vw6f3kZ1qsBjyqXDafopdqYUl7bXPFtTkXHWCYnpkFMH6CIKSaHz5PlFmK
VlDxHQSO+CVsqNusu4MXzgENgo7fXNAY6WaSBcjuTMsSWnPaqSTmhRYULt3QAwD0
yvCiqqcZtQ1Bpc5hF9b24+dlp1y0Er4svudRbT+WmYPdRZbbzutXBCpI4D5RssEv
XcTsYbrnTiV8vH2yD0y79dNnMzHa7ppAjks7XV8Z+mBMKm1TKCwXxoscKgDTFki1
fX3c5XMPLJjzubHeLES3bgMs3MN9vA6CIUQXjgx1q4HLt7co0uPoDbq+z87lqDWB
lulYIWG+DJHbmRogyN+sb/bZWcIbZKWOUpRokSBUZakZ1YBojEzObFMjkmveF9BX
UmAkv+qLqlV5Q449eehF0S4EOMzYSA5SZq08iymKIHqdQejwRkfmlGoLQXe58VvJ
SYsuLuTJQuiJmOoSZ9ePcQrHWxqp6eupodIKtQbeOK8AgAxa1u4Wfsb/+PYM3VFw
iuYyXaCjZStA8iUmXiaCT8XHf3Eb7wswrLJKk/wp8Olb0yl+E43jjZyAlNLAZUcL
lnCIjgZQ3mAWDu7W1ubiy4SDdh6mVI9I27eGvEF5EFQLTdrAEf9x3H6L74gIANBW
68dsRFR7OYlu7FD2bfVeN1DExUplSeb4tRHnjkN2cz8RWjhVOY+U16mgzLwMZJ0i
GwKUgxB0i7etg9qvWgqDIznBFCRKNKhFQhmjF5VucyZvfy4RdIxZOIUqdmpxZ8t+
k08Ob422KDSzLL6QJHAtWn1vhk/wLoPm1426bJ1N9ZxkSkb3gi72iMEuTXzp87Am
mpXN3D5PicZ5ry1OVKQ0/Bjnp4AHCPtA/a04cvUUpaMTVPU3y2E2Qwiv6cPXVwXs
A7ZXURu0XerrLpHhp4R4GrVXdasVd5od+35FaYCi2pAkNMRKrQT7EPJfLMuoa2NG
Tshj9DYDok/WhvZdRhL1C5Fa2KASSp3TVi3c/133+j0V8THsvChtpaaW8TYV9OAT
2Gt5IDBDDtmgI3W7PJpoRP2thDToSRMMu1tYHVm1jGddSWEQQ9jgnd/v2oOYnTBd
sPu1LhDeega5WGS3IkT87RDhQ1597C/IWCZj4u7EpBvEP9XrqDXXXZ93iZjATrg/
xgNatE598gF9vu7x1TwcCbG36BqOx4P1et2w5ia1voOLWzkiULEPJJGIXn9qiI56
P4/XmX0EsiMFPCSxkesZ19PzgFe3sf5U/XXDPe9VvqBPtHYMXi3FBCvfwMRbCZKP
tw12t1si5hvUfvbJkwUfzlIandqBZv55Vjhr6fUhKPZfVyG3I73b9PDX/u0G++vg
trbb/0QWwa4gJq19x55iqUEZvvs+WK1yv6AfVeiN6iUIbAWGw5OHUWa96T99HmHs
l2y+sUs3Ow8JcEhrepV48GCf+WmTCwW9LbgwBTtnA2m8ZHseFt4tIsvdTWR216mH
pAbt603/olSQsw5BGaVp+H2et51mQk+qrj0CK6NpLFk1VnGkkD/iThW+76kKRjeL
cGe3QOXH2a4UMuXze6BU4h3VAYcvycO1qil3rEjCWEmKRDyPV0tNONZJa7OtJAWE
GvLFApJZ2KiUxTtmtNNV5SLe2UvVX+SJ1ybra9084sMY6yJUWa/oWRQ29dUGeoVF
lt/tw56uJPh4RE+K8JTzJlU+CIyvWLdoF3tKy4YCvijOmcSNoVxMoJ7Sm5KlbzHa
3g5vdY+3/64LRR5x9JEJH59LqkrxxQSzHDYadw0v4v8gvWx3KPAFo51ULHmK9IlQ
lR/qKNgHCilYT0lJ0n8VumaX9YawLrqhRkJ3T8t2yyk59wZk6APty8NaOec7BfG5
E0itVC2zK4328psW1KRUwSLJ9MLwRnRAbK6qymx19s8LkjhveTYWEc+njaUGPw7D
AgnnIoNU3tJZENOu3OfzfuOSJ/zayLq5BucM82li3NQ5+THVLyi1ZAphYUKrCt/+
5aS56ZBcpuKJ7WbTT+nEp9cfIieo3+4TYwFAofA0JrTvZtlrIcB/o2fgAPW8erDV
C7U9XBWPD0HrzaXa6Rzk0ex3g1GoHktk8NE8wWRbjplvB7nf/IB17BdXYfszUYii
9WIin5enVewT1udOHz4lXFlVw34TeL/EjSkchvoC11dKUwl0GWjySQw8M/z1b8Gw
0LPOFAs/oFA63G78Ok+OANSALwpeeFBgnfotFWpTetbkX3PIjyTWXbt4xPEalQ1h
DxLFTo2ec+K5STYAhTi17HV2LopyrxcqxLtlxx/CGpuylP05glpFxRzZcC+YNpmK
Cx0x7U7xaxh2hheyYIA+iGuRvGOtsEgAT+070D7EvEwnxyNWWvwZznhE/1xs2g9Z
roXOMbgh1xdMIq1w9Uw8jy3EIHTZedXTnqwiPO4zVkxMpnAsfAB+bUZ71FmcycE0
Z2z2bqi8cBW2rqug2qoMzLNHh0zLQWkHXFp22UGBEvizZcIk5p+QroFPyYzcKjno
yqOQSs04is4nBIxPmZSmABMd506XOZGl8mhnEifgJAu1ttRpPjxXyOAyCWRZJR/1
lPdseZiwOHCshDh4R6f4p8+UDK2NMjrZqKTfgz7GRjKLcJ2vCvC9lL/n679rlr4O
wdBzGyRRXIbQY4YxZpCTlo6t/Sx7JEW2REWhxRG5SaNdB7BLpWLJ8gP2XCAqbpLh
ZxsQ+nRZ32XmFNUCh2gKdxNPcDgwwTjmsn6s5+MUpCxpeadu83IMFWOF8iogsLuW
r4vuUdTO7hci86Umo5vSOPq/lTJ7JqrI0v4TlKy/2mhevm4A4METb6Y5yMpTVVIt
KP1w7/XsymBcv6r72dVbZex6URlfXFcgbDg98eP6pC+QTqLV/ebWwsIQNc2c2p/1
Ki+G1741oxw8FlME1fTDYepOgtVxnb58zUi+L4gGQdrCt/C4amlRtC/lY3POpcOC
E0fSPORyw5osPhO8S4T4wc57Jad7Uot24saUZPD6EROct9QGQ6rG/I6hFLEtlr2Q
/jDkKsK6DMJmdbmZ5w+wg30Md1SSJCmvxvtBimHI5v+NLO0FJYpFUYpmDu/wuihX
2KvH2uPHFMyghZaTD1dpEiPnlkH4XUZKB67qJXwv8rnu0zpalmAZmy+Gzojsx7S8
vt8cr/tk2kcRmY9aQpu30OJDcwSSyF+26dVl0QA3Z/fLVdUONDPLovGEAwWypxXY
2uE8jjOuJamqFw8yqALRn8sdk/PM5N6PfX2uzuyCShq1G3Wbah5eAkXDDdtWs9iQ
4nmf0DCuutF2RRvDc0HaMppLqzq+QgKdUAgGdeuFfvyh5UDUkDys1N9gsU3HxSWt
9vFJrTY0NqI8CwO6+bPTJe0FvFMVShpge52SbuBa2HLde3GiQT0ccXvZ61XbbHKI
67egCFoqv0rOW6Bdhlm9GtWFS58m0bZYetyNna1mMkrnWjXHgX7WwltFqETNUu2v
4Le1C0/u7crJTBkhdL9AxFrJwpWHjefzZAufQEDOzKR8k5ABGk2YBHPLsePakrgH
PveotADFMws6tS+IzeB5qJaij7QXmNlzU7qG3W9huS747MVJP3zCgywUiq7jLpno
4/nUftIYxPZfH7C2qFA27Xky6oCNoZTNj0lDgmxOBFoXO0Fm4VZds/MgXsvnRohF
4UUph1h+Jfihnq8Sl+NSmLiQbqPt/SkrfkYKsgF/Q6ljfx9iGljrYruVIG7Sz/0u
D74H98hzChwCAb0RqF3LQ+smspTYqnT7SD3jum384iRrwy41qK+rotkxJfED7vnb
2yeGwB2RX2v/BRECqH73w3Frnh+JLD0hj6Kptv7jLFynhfqif1VxAuE+053hWida
Mc5qOn2Do4UaqT0OOisS/Bo7ED4HRlWvZMUvkDTIiSVBNXq/Aw25GtGMXjLvw4sz
/XPuPWu5YsPjnCieQGZZJsaz1gZ/ohk8Rnsx+dGuqMIPomAK9uzjlYbHLM1RBAZQ
vN9meumMu5mxkz4kMgKOgWCaF8veRjZDPrrLN5dkNb4KZ6hJd3rJx51isN1/aeae
FYHXKFFHSLgYZn794lqThTOYz2QziEaiuCZ7a0tFNyLnWozooS3O8prT73D2vhxZ
noasqvxNtkrzL+42frsHk7c8XFUyQim9+97SdcYGof8eZsL8RyFw1jdOTNkgfuRt
IHsNaUTNweEa9wm8Ls9Y4RrkBiG1R+lVTxu0Z9v3eVdivON16E7kdyicgAAlW4KB
F3lrENMr/6Idtu61MjZZVK86vkSX2qh2It7ynZQrKJQ1UYO2xFMPX+RHM6hcwlfP
Wxf+pe+z+eRbc4AMLUVO4yPJvMFHxjvZQMMbr5YLSsZfyYzBRRNpwYKBIfsu4de4
k5JAuZPd/2ZFthnKHCBszab9+ZtMgB818hjGLoC1F003e0g0/hRsPQcnevYhH2xI
2PJKStMcYwZXgIjsc2qQB0X4tqb6jsg3KmKclqmWAqP1PuQ0t6nsqeWt0OckZG51
9VroMsxq/TYE56c3pdZyQfWh5wvQAfwJkxX5vWdsjJHIDfDbvjHDbHZpXS8nSy8B
OkAPRy/3LVvoCMyj/XJbcvW7OrrkurAyiwFJ8HWxOtb8b9mnzfgGZJ8aiHG9FHjM
Rn8RloCux/n5r/0paXfUpLG/kkgDj5xrOkiS3hv1ZLSva3v9V/6RFvvHrLOKqln3
PWHtBR1H7P2JxVBn2ylyGQ5D9GSWiMv20Bjsv+5DHRCFMefFIHVw5Wo5fC+b7utz
2jEAsl8l1lQ8Tm43A/oo85cctIDFc6CcR7abMIoCYcVbENcqMyVp+p2CAjd3isL4
lm+aJUcSBCZge4qR9ybAkT+BDU6SkM7rQK9TcKcrZUzzi+zHrCp1e06RGvzthNTw
lhirI2FAgPv6xorT91lF4dY8HvX0jzvd1pMQF5ag2wPVZJvjDY+/jjTdC7LriMnB
FTLF1X8Of1Y2wDFYBYPwvcENYjyQJb+hdbmew3/BVvNDFDkXU7rC2HJR2zC2NP7d
wrdnlWpMrHVKgLLr3ZlkSVA99KWHmW/XN6EzLXwtM3T39TRevvG/GYsL0Rpl/1zj
owtW68p07XPkTrPnONPX3HKOPpZxjIIMWeJ2eG6TBnYs4DBbK+kkU9dP8B34hPF/
sGGjqklndQPWCyvwCbDkobNBmRRZepYAK7kPzquT0F6mE60ECzQ6nzRtq6gW21xm
pnEoGfHMDXi7OHQz3otfVBNyUdziycq9HfGeZ4DqM1pN6X5DXna0GrBtAIrNj73f
rMjXZSBCAEX1CFtNbxi1WjtPzu/gwTj3DLJ6sisso9cT99GyBAHXtfpbSf9YpP85
+bbMztJ+up+GnHCQeXJfLF8GORUTNEjn4sCBEZiDV7wNFMj+J2yH3E+waEtDumkA
fD9hcL06faG6RyfEjKxlcxUMhM9lSfED6GeNFF3/0qxS1uKvOrPkk2Ned8wqDGNt
BTQMTTMhwwlnmv+P2IY8Az/UAxTyBuTdntGbAPIR3FR/I+NZdR+8sVWeIK6GH187
9/trQ1RnknRgj4POkzKSc+idOiITSfwMcM+/Pu1pSy3KDOmWDjNZnVeWDddtCXe+
awnmOaEW/vlSIfvjnSLodH/COOUxAWP70Z/sMoecHxsLEx63jeuxYa8YsKYYtDI7
Lo06io61F1bdaSjI3UQLTRpIHS+HkrkaO3h3lpcItAtPmFZiVYmkgsRbfxXOhwJy
lXKnVm8q4Gu9U3Q6PjcbI3ndf6vulR2jYbBUezGxTUJyx+uFLiFRtaARcJ8Bg+MP
Mzo37YDm8qD9sMNzJ9kVhxI+EAOCMmgnQjDzIzJlLYl8hDcz4w0vhX0mJalnDTCR
0WJ5v716jSzydDjICOi6B4U7rYuRP8n5nx697a+TqSucoCEvI22gQo+uAGeiudeE
nFLwlWJhHoT5p6p0q/Ks/gImKZp2TqYPxIGrIUrSxdQh3yoViBv7SXcpmwC1U3pc
OpnL7leJd0tOiLJI2i7hdyqQ6boxxkjOstn9A4jL5EqIhtuOKShV9vjM804tgJYg
U4qL18sElQ/wtb7qAc7xKbfCpv/4+QB/zHBfG0wp4xqV18rzkhKVqJgMQThjMBny
hdakSOokv05bugHUyfFoROwayIO8vln2PAwE0KbyXcatqYi8UbNJ3KRcD0wMTf9p
urbrC5L3YIuc8LoDElJJrU3XpEUFn2L5Wpfbg8uP3V/0crJAmQbjjHxNC+vCZTVR
EFGgmkGXNXneGggeMTMWfhDzR6cNit4q41uG2xK8Qatg1jDWs0QgW8QAzpU/0tN1
pT95Zzw03ufrzytHb0Lzvy8tvAQv7cuQpT/FM7pOV/D0qGDEfFp8pbFf0uwU7yNL
WlX+nZZ8Qf0+7nhlW4cMZ+vViswGzPOb+FT9/7zS6LBT1NHRuDOMaduTaw66UvZx
+xZ2ClfJsQj3gwnVgWEHMJsOM4q6msLIyQMSWhabug0vjlOPq27O4b4catmz76+V
eXUZetK7z7llYM1Bms492tBJ2KxUbcBKC9KBtXyBaAzbxgV4RkJxpPOu8UDZfEPP
k0YfnoAzUoOL1uNHJlz3msVBhzcBJefUkbWsa08WCFVcrg/mxhx8YVIbRcT7JQfo
+83XjMaK3Qng0pKD19FVzeOiBSrVqsJClHL7pQxG0bifO838kAPPC090qx5XEctn
HSrhLzycKE3xSpJuP2xPnoTUEaVWMXN0al8W0gBBFFeQ5wi07nOK9/bHeffCAuuq
E2trZcl4Z4v46jS1QPblHOndcUsQjno4rrDW9xS/6uyLDOBLsST0e6Jxt6iP4DKm
IWf0zPquI8RjBQIr8tuc0R9iaCgpGTTe95DjMX4bhQuBX38EgZClVfhI9dKbSg3d
oYc+A6kQoqQOI/Dll5i6jbpASA7r7H+ODpcrF8B2wF1oBpZnLsM2eyoNLo1Dt0ri
/0C0G4KpAMPegz54LP0QILLQ4mpif8f0nAEyDCB2BdFx0KrntoVb45qIJsRom/JO
+EuoysO946H0De/pVWBMyltNHkXkEE2hsfGHqkCGHd7ved4DRkG8hASQDYWog/G2
xg/r1z8dE5jKclsVRqA7z1/TyYQ5Q30i1yEaMmoULWMhi0yusWZ9Qu6epF5sNo+k
BCecxPH7eqJLYQ19MpWhf8c1ZpTsMQOMFCN0YYYHKO2vhMDhakg9bK3JnkSjgM+u
jF2M8R6ZTnWuM7Ak/8/xqpRLcGUMXww2ozWanTVm3MjZXyLuWuSyjxiSk70IMDpI
c4uNxsIU2TyJhbOsvTyKUnyqqoVn8I0a8qsGOcdf+C5Yk8w2OyJTDUPoyQq2BXFU
oRejUq9/ZLgmo2J7fcZ+1F6RWbrfGfjTw1LgBsVSodkHhiSxVoNwfNQ8sSCCYgEj
ZGpDGHAkxn0l1jxGOorl5Nkfa0AAN34HcxsAvWJlti60EAqm9EDUwqTZGqEftY37
1+fzoSh0FMxsmhHsLMhNcEIww+ZQomWUxQtA/z+8RLkjG2fpnoLtKp6vB58zTpV3
S51EiNCBwA8QKp1Tr6WAqEnKcPK9YIHOGRHNnEFx+kmCnPZj1MoydVTacWSSgr/e
TsfsM7yw51F1Ey91P2IYdOyVyH6+9Yn9FnaQ6ORkKhGnESjrHNViSlFed/NfwIby
5ajrLfFc/tatXUfFX2myxYCBJ03LuY19HIIHHEJUMN51s6FdIJ1wHJT/+Ia+cX+3
DQYLhp6YqrAtJ4Ffll3SsHP2MuJClm/W8iS54UEOa9dXW3O/LO8ZtUX+h3ZGpk/e
VijdKB2CHrpn5OIxYdO+EzDyAHAXK/9eEL+JRB87FlCYT/HBMVYl0Lw2I3jo13KL
x5PNyZ2HVcQ14YQysGCbO3V59GPMkbPepoW7etTRyn6PGGNzi6RyLPMeXN+O0nem
KjHZ0Mwftt+4vr5tF5EO/9EXyV3wFf3qMP7zDeKO6rlvI/4Dhgu7EMMDzLTTe4l0
cjQm9AB9vqG/SeVUV0uFxG40v/w3Bw9UZPaYZxR2f+srWK8W5m7h952jd7XSwBg9
qvv7kWHDdZ07tFrUmziniM/WInY8Eg4JHZ9AKMdI62fr7hemBtMvPbR0uVKvXWEj
TuI0bOTF+RCvrK1ve/EAcGQdqiQORNpKfbzoDay75u5iHUVXqr/Z9I0BeIvi9GNa
rF0JJ16qzfNkbgqzMuAHVsx949XS+M/hc16ABOCSasgE3sqiN5aotuiP9Pw5FxUT
pdvxz5xPk6lZjY/tKtaslyXY5rYCnLpqoe/DGPtlYZehDXgF96IREs3XgNdPv4IN
Gbjx1L+hahicE1pTsllU9gT5QHl46z9/zR7aaitfCKNrNUDL8hDAP1LMMXPOOvVh
WwVmJEkocqmun8Tf0hYi4PcbD/L224ZVSTKzSw4vinf7PnQznCKIhPQq72kZvwzj
lfy9rZzPANuTwQe/dz+LNOEhK7gamGhR/+o/e2gzqQM41vvomVRwk46G4IywjSkD
pozxRs1ENYVJiCA48O33sMT9l+pLSZy8GReB1qM4FXqrx3XDKuWjJU1GfSjP1+kO
6ttll+8b8yqYQL3Zequr9DTHVX5HkXvUDRoqasFkwfEDABa8R4YA3vaKhyicYRMB
LhAYFVmgXZbkYSpmWuRZu4xy//0ur5PNWHJQIe04dQ2H61tJFqyYl5+6C5lerFjZ
343kMxLmRFcHRXqTuBtqSY4erB3+572YPLnFj5Jm5VEY1UzhRkSkm47Fit+Pz92h
NBu42w3f/N0AF2kL0UXhs6vT3N6A1vJtf1OsmZotyAkCDGASnYM1oxWAopEB3G7F
1Aj5W8Pxknp98KHlCF6r2L6aOlKnmnnDGscMM/brh7eQRFeZTpFcVLLltTp3OKOL
AoJ+IdOaK0gNYf2opQ4opdBld/zIbVkZ+8XMRlJXsSX2DquGXW4Lu58Sqj7NW4yr
DiN9Cb6vG+zG5b9wywQCveRoVXUYn+RS+y+iJiUIw3O4mPkJosR7Ym1dsBgRimWf
vK3yX9F9n8s42yzyJvsKGpp64SXfwByrqwVSmky3hnVfEi4jPPOcY96NEukx+JVw
ZfBOysd30Pcfs5sw6nnPhaIRL4aBzPebfg8/YZyLRlaGlyp1ZFxLZ8BS4W29jyZJ
gr7GeXD3p+cUZjPuZHBGLXqsPE+ML1UXYvmDrbfw8hK1d252npBjvJ0fT+hL0UsK
UEZnbvkuXBbGaSEaHhFBT5tbwS9dqepsmPoN8cWqn9KyHVt/3fy6PzRqgwj0zYST
/RlFB58FsyNdUXs0EdBV8cTZ0/RG9rvHkWp0i3N3s11eVNOzpjxuA+9/YIQY5VPH
mskN7OghHx7jlV2XGdRinAwoIY1ohblTlPKMLZKxuUZuEGtMKPK9wUTo3iTNHUQX
aE1QusYbPc32zj5CUqi00LAB8cJcmmZo9sY6OGZTuUMsgIA60yeE77tZ/hfaN7yo
L1sr9twoB8ePqnQv2miuDqynN02hf2wSmRU7BJaxnXYSwl87je6XfUCDrhFWmrnf
AZhvj3WAHLesZh6zQpE1kpRvLf4ytZhD2u0I4gBdE+wnRB6oMqv5ZSvdSCcp89eV
6Ucq8SQ1TqoHPZOU1qHfSnjOOm0WOg3Y0IQpvtILRdCPdhp7fUb9PXxvhcJl2/oI
tJBdGLaasMhfJyFyYmZNvrQbI0huXL1OsCKC7ZBW9WCnCw2BmzIbkb6MKlKECPlN
feTw+ynUzkgpzoo3INrrZGLB1n7oloPvX/02U7iCfbeFyr5rxJNf78Iw3XDzxIrp
Lu8tIqWGE+ZX5MvLtFDXo1TUbOGYJ5IzoCBjEXg8ZkGeHMJdwHmF7JSzyVb0Hj/o
TYT+5LZ19Q4ViNsORkvD2o+HVo3ZdPTz/SDMeSDZ4QThBJ0BOeFnZM0U6+RkNKA4
VyKT/4RdWfGB9LAdCJZ4WpLH+xyjdXGRLR0seC6ylqihCfgPoagqLv3jLg3x/2sM
u1qpemgvLIpHThcyC9bfeQX4+9Iioc+TQwuRl8VaM6bGgdt6IMONtbeGEdLC5o2D
7/1X1RVwvkOhRaf4xv1z53tX2WqxKfTPiYgIxbVjbOrikrOWcJ1XKGwLLiC12EF0
DCmmNiy3P7K4Cf51IcovKjrGkgCM+X4JiUikNSeXJBDOhONA4iARJm6/yqfOVn1I
a6OgUJE8HXYjopJsk9SCxHW+MoijA9FhVdJO8OWcE89AYVd/s0jXqaxdyy552Zjs
58oao5S3X/UbMfxMmM4GKOx8TEwkxtoCYh/kUpRd1yGrBhvTfEus6CRCr2Y3QSgd
Xr65hqOIvTljcgNe5eoTePyeFWk57Y7ekq1RmAYO+siiEK7nEDv7yvD4mMl1FbVy
9KLWGbGsq9Iw7uIEGoNib35zZh+jYbHfSZIPMMFnbKboZx6ZW+zw3SHJ9XFGPi8E
QEHhpCPXxCkIAIHu9hhhf7EkX0wC/Sb7aj/tF5yuSi5zBM/ZdVeTpyn9zGlnrXnR
Tam2Y8FHNn4odJxfODbuZXyCBqVaqiX+BNHd/cYvKK92WhqszMDUJ/GNcPZNMrMN
bwa9DWZvCNmBulRaKjbl+QBMCwWdCDN9SXPC4BN5FPpwGQF9bb/4rGSxnfahMTUG
I9v7tE1wTcsNLVTTloEWVC93dpZDMkC6j3N1JsVV8fDKRhC8Wwk9s7j7r2amGzBn
B16detDj5UYPGJeIvKRF7lDgi6ndVwcU1hj5/VgaZO7S/e6q4EWhT03IydFTTvlv
OWfxSXhzVvave686Zj+mYT5vU2g/D7xcBYJNFSxGTuzvd/KAfvUsqtEc7bvlMKZx
AyoBY8zJP1Tlsm+RqLk/5jFh2u+P6sB0kKqG4rRmP9xoRpogO7A6IXynWYRWW1ag
d4UPb670Xudf90IE/YF/E3wJbfPkCItrm6Up1GHJLJyKu6HHgkVYyHqe4Vm7tHuo
576ofZrJDraSQ1Jv75J4hDTDTl5JbsgYpfAr0NJrdw/dBgvHNkzUf/eoyl7YuyLF
QNNPZLUTmBoQhKPY50y7Xocciq5+Szd4+4Xd5O+4XWk/OFo+LK0yMD9JkdE///99
wnjbKpyeQ8F92GMEHd5dnQaBsiXNfdhpTIkJ1Jbusw0Qk2O6FzI+n8IQBzJQuF7z
sfNE50CWB60OEaTPOci1nj17yzh+en7T/7rJKafPkBneBu4NRj29HNfUUrKO9EeC
nLeiMoiHYWoDlOGgP2IXbJflv6kJWUkBIEaBVKsnW1bM5D2cghzQVK9nPM+U9aFY
KdDukSkj/C0mKec+kwXTUyiIOsc/nCzslTE8dstd8Z7mUR/XBfiX13MDnqnUXOXD
9innfr2lonc2KLdT2KdMc51bUCp5F6pnLK8NBiSEPxdFDu0+Jsxg55N5VnT2ICDr
bVxWuZ8/cHOVetBlSEqAlDJWkhOqbJ+fysOM1ht+B3mtCNGDH4gPHVGhcueWhIuT
Faq9PWUP05Fj5mmi+YPyO00Ccu6RlK+oYbjAcPb59iSQD/oMLW0QcZjXcZQN6qwK
2vGOlL6Yle8Xq2yUIFEOYwQA+epbi7zifZdCHJzl9fP4wYxS8qtbmHu4iQrMajxx
4fGmPirUYvb8Ktuf3htTMgDJoPN3nn4s/QMNuGgKFPI4AKRZBRjdTNRtVuiDYEZX
+BxbqT7VmOUrGkz3XF+hGwEuwyGSkKrB2M4I+XgZ9CR7SqPN9M6LyYx3ZJn4x4BH
fkFgoa0pYWqbRPwkSLw66Ok3FTnXMqMrV+HgUN+u+rduamlu0loA3jDv63BbWcaJ
pLoCMot40clfxji2QcHesgeZO+HLHDeECsf3rvRA0O/KKv9CtWpyUwHGw+gqXoIf
O2TOkdi7VDAuIeokN3k6T3Eiu8ltiDw8JwmDA1fB6avON7jFkVeXCYutotBET8iV
LJoixpi8HURbos09RzOJzjacnN2hBCziEw6MoiEbIPrROHk+CcLTi2By15WkRVBD
rZbGy46BjOGI9DsPGcTiE7WnyolMbTP860GTnTJ7dQ+MmaEkgJUh5sbiOB+hZSAJ
w3B4xdnB/ogrgOlQhoa1jqO+ObB8/Uy0nYgwKSJAeD1pFrC8p3FDgiNE6RFKL50r
67J96ThxcK4LARFYZFAeSSDKYhOuOSKj0MQNQaPbROaRsLKPbCoEyT05aoxgnXCH
QL8zmL5krGLBPfwvLrwP4JuT0RyFf4+YiLL5rVFv0mrPadm4YuG7yrn+SwSJ4PtV
JoAx0qtyisY9HFpUidwk5+14uEKpgig1hjdoojillmUvbwdsoDv7GDYcd+Lo2lsv
/4GAoYc55OapzKxSXfEYJdr0+bcGGJNjvILIpdUdSJr1mZyKZG/vXSTr2r2kAZ0w
j0a6iXanUEunp5sWr/lwJD3QekTmFzOkBUyuD4+ape84+cJivmBjTk7EbvMjlb/p
4AXgU9MgeJqEXDcZmVD7PrE+TRG8B6/MsHTEWg1lW2dQQmLUPgQsqz5q9rlzKPh4
cQWJHEi3uJzebNzXNqWjGu54kA1hhU6NC3LEV2A6+ZWDFyQuzVz461UXJ96UPASa
VEXuM7tdfBYnke/WYlT6rUAlb3V1f64bq595AVHtZsBw9jdoGyN/7fSRzKoZxyho
u9513cLpVoJiBPcWsTEUPbM9Xkb9yfi0SSZAAYBZmtErKOMmdMvksi1p/FeL5AJZ
ytaz4HWK8WfqoIJAGsh2MpmAJY6D5DqldWlVmiXCWv2kYBpR2ae+EAGWen6/NNaw
m4CBplf0ds7dIQgVqARsn6j1LaTJiTR6pmCzOgsyiH76gPSNNKul7up3W95F3Y+8
g52zGHvJnrTyCKn2fYlWRRYYK5ch6o531YKYISSRh7NziDxPm3sos9MdMM7DFYrW
UAyYDYkOczIIYZwk1eQ/xXD0QUrDX32QNHgLptSd/yJtktjomEy6AkwN5pfK7vKg
mGq0lziGbJXRAIqSJ74ucZajw4fjWfIIgjCvBjPYMaP++KF614F4GVlctTvXa8A8
H/0RzqZ8jIGzAcVQGGA/nmhqVlZrHKB0oqXTC4sv1/fw8XToqlw8rKo6JWdJ9yOM
4ktbY2OEpoU70cAoBHKFCA344Qv+P2nLwnFlfR4WGi6Dj2JYjKgdJNsAk9OWum0U
6ejYrdKeURCXYcBr79ZS3UKrIdAKNw84Na1AuBCbN7uEnDGadA3o/ytjGR391oNh
urCHvBYqkbXiTokSuvFG6f4Nyk/x9JaZ+nPY1jYXCEOnCOKwdOcY0/XaZ+1FjoCr
okpgnbdGyRAEU0NKEoj4HWqaAvTzcox8xtPTefLQd+6pbrOx4XoZqoAd0XtriieS
leJcD/WcxyQGWSrBkZnOabyz7JQDMoTs6WGBmEl0pbHuu75ORJqgrRxrUXlJJrtE
Fful21VCXcWyMwD+8pXSdL/EJVANs1rqsy38W751P/noMWq6eTc/q34FypKIt0nf
Q6eqp6xuEEk/7TvCi5H3RWnTPft3uu1a9+pLQpaFhZjLp8rUUBDVEscEJOs7vLdv
POawvHpobSQIwX20Jm3TXWXEuyESQH+u2lS1TAQ0FHIIbmUmOkIkQciaIrYArF6X
Xv+RLWh42WCtfnx8WOoKU2kMo0GLle8mw29KZhUjPB80HdBFnQPUwsfIlkRlXXEr
D7V9eIgGOhyQnRKRtyVIFad92fvQTN5kQCe2D95ExHtfEMNBY9VbCotfLuVrjN2s
vyv5KqXG5tWt554V4uWSmpf1ETsW6kgUipZpvKY9SYiN8QBD7pLyfq7c7EQqFE+Z
L48aC2f/13wgsoL7+EiqRyAcazYdsz0O2oRbZdhYVFzbAtt4caDOzEenZDCkYBZF
UGdu/NHGZJpOvLCwMJGInxHc8tawi2YYimoa1OFgjFnfgtEltzPDkX6JrO+WGeFX
+aiInEVOZ/Q5MjVz/mC49JT/eWngm2Hyx/wgYI8hqq9c6jqO88s2e/htwM+ZqubJ
OcyxDh7bOZR1wnr1x3FHCP5diZStOia0RrOhGYqjXug5xGRntFEnwPj9U4BV2UDb
v2L3keBX4D9Emarx5UkErd7mrtOi5MEulkhOmov8/8vXLNDRhhHEmv7t58VgPpcl
osvbsEJDGORZPX+C6Daz86grNm3cGupjBsNXmeLE11HzmQOB5EZ4nqwGbl4pKVyt
1ys0xWx5K2znsgBZ8WOvUrqja2X4E+jd28q+5EB7E3bi66pHkJ6VKB9cgjIrKS3U
zsXbu7PBiynW5Ww+xOBo/evfYIxMlMbRObgBS7M8FOS4xrozrjN4lq5LoUW3ODCD
3yAynThWNgTWXg+1zFPIN2024YhDP87ZpLPQQrApZk4HEkgCNkRHuKtytSgU0Ne9
8Y6xwlxW32oTrBB6h+k9U+w9kE9MPdBdNpWszwZmdeqSHJ5TaK3H/ohZneilJGdn
SV94sQ+6TfwjcMf+UYEfWNMEYc3m/vS6m8dYTYbfITV/qnInStJN9oHmfWccverC
zZeQFY0X4tFsKf4W+dw+cPCnCcr3geoyPXaXyDAhpolI+jBvsPG2ypj14V//3uze
YOcqYW6pENT70lLbbu1tnfzua23YEkdszyPw1yCQwSLVMFcERv8YFQ72C4LUYwVl
USBGqWDKqCejqnMAQDPAM7CaI++y234+3zRnmOfKAMeaZ40qfViqUUCHIBE02sm9
gIzbd598Kt/m8EFP2KdbHGJgPtJ9I7TBoOeplpST4strFxH4LUymSyBREsPFkSIq
n4yrKcIQFDj5dLRoVRfs1El8qjaGgOuU9pcQ2zr2wwT2IHiDvxueZe6PrUjlvxQE
w3RsM4FvDkZLCKkyhdke4nOR4YSiNGVkhO1qCKTyjB5A9gfKqpcQ43DfSF3GFM25
3MjsnKDXuSxaRG2N0938UUX4ZgeNajyzjGKJnKlicJpisJI8xkTVxU0OxxGIULaU
63xC/YDM2XkIM3KLlrYXSqwarbljAKxzEsdxzU3SINt9uyi/DAEcgBqxVf9m6f4s
Yqz7XlN4Ihd9YXJ/lZ8PCOZlDRSwK8nqwLH1hYaL04b1pqua8cdjIk5obE03cjkc
zigoJx1/Q6HOHpDnm+x1XPi2u8dBNa2fHUPYBQTncnZWmu/ByIf5lBFI+Vu3PoYb
IkymE7YeUF7iOPeOTFNk3xoFJs4il6FFBSY1Vxmr/q4V3rV7r/iqUQnD17y/CUP+
ZnmbZq7qGJbq4cNKJ8w/sEQ8ZDVySDjmRevFGh594wrgI50uZyQtp/enwKvdEmBR
q3XmDIOajaWSTTiKAyDye3RMAGgrEJf7dhy3fGbyv6YpySxw+U83MklUJobDMTwy
3Hgwj6tDYqmNrQdIHiAVcKFJO3GZkgRjKksGmsXEiW2LBuFk/mPFeYb48pfGrzUe
3LR3opRieK1VgmvOWJNbgoWObjcygqj2RTVagnRNuOWTd4ZOEj6CXs19z0kYPQPX
BDwUddqEshy2QGbXXhhQ3rJGJYoqsjXuLvn7YrCPNR09MjAgfSedNaKqMofVl+t9
vh4SKGuXt9HkJmE/Dbx9LQFVv9XKLuLV6zWoaGcQjN/pm4iipemSj0tCX+Lcf7xy
+n2AWT5MsUyZYxP9MqtFcJpHo1JamBxKnk+nEXw6qgL5+MisuRWWfTRYOgtStdPV
qEQIRNTFH2wkLdv6+TDl2uCfFVyZ5go+HN/Z0m9QC4rq9/QX1CVVfRUnAR2ZMpik
SoptoZ0YBPhFHWSOq5cgREw4pe5JNlfwV5Qq0euv9l+o9N1dEBifA+oUAy1enu0+
fj+0NqN/wEpK5LSnxtk9BXEw0m0hUHfYRz725QRoUm2V/xPVZ8nT/Z9G8WmnqyvI
M0xBAR10+p5xXCIPV6vFd195ZZXvjWySmzhW49sgsNxtF5yqefCLe3HH6MCZeCin
MgoA+/PWKaHUbwIZA0z8T4XdSjm4O5R9s0Ig24B6Vq9BxKXMs3FrnaSos1hYHMNc
fuD15NxiNvlD9UB13mUqvcphJ27E+ZZiv6IyKVWHUVW3xNCxGg4I8Tz/9FzPUJnA
8u8ItY4tvfILZIez76y4HP7+zUO+lXNKEK+FdevE267kp0RZfCs6hF9ryiv5aKgc
Enx+e3uH8LbtP9/+7wiWN2Lehm6M60pU1xZ6d+PYmStMDfPtGFXGYaotTqmlYTiz
wox5t9S/PeWmJFskotIqfdrcB9UwqRooepUaxnEqYuAp5N9oWCe+oq3HxARzKZDB
YNWeHUHli7wz0jjqrlq82naTUbWlvHbqyyhh3H9wcDk1DKdSn3iOx4AZnhRwxskt
0no1e2sVtvL5LKjPcaANyiaJnxxgOCY4zWwxqHA9niDXruQK6/b64HC6/11onyAj
Gc63/z5UwPHFx054OCCiUPsbzwm6FPfAzig0Rs8yd4K4MVqeAgA4MfNb180Yq3hJ
VCR36rO79Kb/MoJRabwA+XiyUwwFeXLq6AEJh+8iuqAZa3NuwgwiLKoIkUqcNXAJ
/uYR/yaXTORJg1mhsX5drj2OIBvgxJeuG/6UNqJCsQQNmht34+PMVlqDKK7X1Sgp
pR+/c//QNAKcmew/hqHoQ3RPCbmAGpi7OsHO9Ct3Bn8oFORJn5haiH8++FAEQodL
goPmm/JHRmPhTecmkm1xU1XroROrRwfEjhTPtkP0LaDnCus1tV6F8e3r5lbBfXW4
+JHbF4AMcA2HtWSG8g5HCJQzGuZ3klFtS9WPIOkoiOrDeuOJiEaRG6dun3X+LDrf
PrBEQCE6JfVHl3c67HlQZZ4fn6lJdF6XAst6Op6n+itvIZiqYZpPLJYoD+9Dur+T
1IT3tU3vDPytT8zpZHPCMCdIPBAuhU3qezHgiiS5JYCzH0Z7Yf4vEq0Exo31B3Be
63vDbEeZ4eQjfsbVNoyoBQTM3Ql/lqHnPuHzHSqZqgSeye/SVYymTi+kw7MWn0er
K4HsxDQVjF8YAtv+xbcTul2Mfhe24hNTIzpNQHMHPsdZmsK6fLTpJV2p0t82RO6V
72a3xDqjpf/6gIHFPypYvzcdJuHeHvTOjVK3NcdPDK/RGb3xby1JT8v/IbEnPX/k
MYApiaAHF65Zjw4To93zhQW0ZN4uZPREftXb++wm5O/SCA6JtAWtvMNBevjJbXmI
zZwbBzpBy/FdpZGjaPc6Bgj+in0tru1Dby6+V1KNCY3T7Mhh09c4S3PkwPCkm9lb
aoGhGv0ELKw7+PoqLlaZPbhYQ+cqW5+8nlN6B1/sYfoiA8XdaIzy0OJkCcI53Q0g
n/BqXOL8lUv2ilIPBnnqrT390Mxbl+tT3Srs0O18EGfZW7GMgX4e1qethGRWtruR
V35hHdLoVUi+w+DsP7m/XuZOYy9C/uebyrb66hO4Q8C8h2ylO5Z2rSwYsPM6rvcB
lqBjWEFnvF2bHwgMXDKVJMRctyeuq3GFEIdTSl9QeZ/T59BQsoL6hgB5NoHzMZsG
5dLabuY96XUxKOwL2KQaxRyFRisIyHNbikkP+Bnj+j0Nd5WRj9knxkPKfs28xavD
I3wUcIpUoCz0lu3YVYdmCulQmYJeAipEOqCRJYj6SPyIG0cPJN4I7ZvdDJqogqlc
R06Ih6UYUoZTnVDu9BjJjt0eiH/vloMz1a2EMFw9rRwoyqJUwGAnUZGAhybAeiZq
xWUbmjWYh3+Cj4amefTjHzbY98dSf9XDum8EgParLQ8coeBkKnVOn6UJHZ4Skf4v
+MRzV4/XlKqrgYj4f3t4SFSelWOHpGvI8vV9DJ14mtSMHcJ7R7WBrmeBtZcYwCxe
raVkbcm8GfzEDOdULipkCO9Fn2nVxdIEMXqpQmxBIv3+oOcBxIXsQ1DVe7r8fvOx
yvfRTwY5z2I2Yzevf9PXG3hGIqNY3UFW+cG4+LM3/f3/IIub95+lOz40/y1QHOWo
U58ITdQ7jqj+19gPai3+HXI2quPvJQFqDkJssP+flKMfVgBk2+jnU1Ilp6Cc7Vrc
AqgQsKn7J3xy7Y6jbZs3PTI+WNvRbcZyAtNlvJVRmFWBn6ZEOXuey6dZoJIogT2o
4tuDcnTo3vwZHaI8tEVKwDSnglzmC3AIZmS8/hZoS0xFxkfHGg2y5+L+JPiXigPN
t1r064k8oZqS1n4XM8S/TN5Dk5j4nG3DE9Pc0cjjl7PecNb42KoU5qvXtrBTLJmK
dHQ45AbYUHyxtEgr6BuWmuAhTa67xEH4LZ7iqCtFVBRSWk4GeFeyihvdUV/Diik7
GgzbGcs1ShI0vPo9hGXQL+gltjtGQvs3b0NV7aHla4jmiWyQyhzRkU2QZO2TOhxT
woGmGA2hRtvkwN/6+Mbq4U11MveoxKlXrS32voIfaSSiUjHzERCrNxyUM9br9ogu
397aQV5TfQSHYjO3SCQNbe3j8JZUFVLy1FlQmo15Wu0F95KbKr7ZCCBax81HRjOT
LfNFRadvm4cCqDsspGhkJvPHqoJ/ICcmyvXS48bZbfSwJGo4w7VibOUICMGJkGfj
BPTWDJYZZCkpCIzh5kKnrZc0j/SnOSqwvOlu7IvkV4GLxtXTFrCG4ras8WfC/Kmp
+wVFwUS93fDL97Fpn6XamM7Fcq7V1YsRguoKXxHvwp5ZlbmaUyV1CH7QkMcI50Rf
3IQC2zjtGqXZXkLbC372EGRxqWFg/LU0VaQ+WuukvY0vrPrWrIZFpLYPDf2Bj5vy
nZJ4r7gEp+gtgii4bRkYLMhEuFI4KI/ujv8DBd5RXye5B3gLJfnHU+uXW+b3qLRP
oSjudwX9ohuBiapTpGwyOYJlBCm4PeKApSWNXtFE/PWHl3e0aB7Xdu9qql3Pb2sw
6ZOTT4bbBvfcRcKQMxFK8jFwivdcWciIMsV7HjOApeVx/QE73y8d3f2jA4u4tmwr
20ePPRPFS5v8b7NZxXMXbTUVk8dk3zAn6imK9gSHYLk4hlQnoeP16WWt+hUwdfF0
AxHaHziZl26uteuYAc4sm1THQjYPoxjPH7lpYbY0i4NRe+OFYRC8nXw1rjZ2CnpI
WbfgIbP33oYe3deHxuX/AamH1k2F34nK0q1mgpyk5nfOsdfmTNs/Km+RkbBWCUW6
goxeKbmBd03/eZaOHuZgKjCYV5ixZz3BrXtUXA3JIAdozkBjf0yuTbC2hxXEA52X
IAhEna/3ipI/D0cQPVcjcLSeHM9m9uTG+SeKq/9mQEjdi3tdur5h5s7nYxFhfBx3
EbtALNnwAun0syOlFVs9iekNV94U590KegpJoWbX+6rD6QwM2k7hTEdsyo9qDNZB
5/SqkcApbX6ylbXftgrujDh77FZM1cKhkHofUWEfRzTkIwJYK5gr9hJIDPHL8Eyd
69eghcH1jEEFdaTOhLMgYmo6KckHqcJCLPZ1n4i4Lzqcx6L3LJucekLRh4JOk9n1
29MNrs7c52ENt4k1/jI0IdsVNm9kB8qFGLM/hrT/MDhrqJ3Vut9JjllBVDqDiSSe
HIgJ0eOQe1fETTG+gM8FDmFYpPnM/r8M0te4FCaaBhR2F3pKDWfj5v+S/koWZc4D
oXAQCeuyWFjZHyXmFxm5UmorOG+uLdhd+5/wh8ZBX9datBzZW1riT6q5WtL3kT3A
p5s7yrcCuWTd1KuTPyTSyNHPl7ce8IfbmHsiMRzD9gttParChf6dsXxLIZ6ARj5Z
b3ohueTBJ4qQs5jzvBy00xOcHB4E/ZflECuq36tfaSfHxM7n8IqvAI1MOccWuUky
+7cfviKvM6TD335j9a+jSH7VwbG2EzaVZS4PHIYHivv6M4DXTaLOK/HUccymcuZ2
9DOGw780WMZHTepMqKurYB52T0jJVyX1jYe28KGTwrLB+GLB8h5loAvAUaV/pxdm
pzoAKfNT+BFOSCLZZZOuLmO4+IhROr1pAKdd1b+R/sZ0QMRWJxpUjg1+yx5oMnOR
gWF5c2vsTZ4ediVShn9PPcJJl9qsXvRoTbnXmeWQgaF1/rz9v1nD+w9imnMU5ZdT
xKzNJr8PBwQmDoGuBW2AZgOxG6E0zRD5EM9hbWmqPEql+llQY4aVtXDCIqZ240mm
meykXY6zBWiAqGIudN+A2KSuQS7/dHMHBLukyspbvtF2bIB33ZCvMkAaXItjPRZO
sfO17IyPCWnNWRgpb1CvUwpEFty9buIRIQEu10aYU9jySpfhTu+beVZHZ5f/LoHX
6wEEeG3jSOXvfzVCc0wuH1YT8IA39kSxXMmoyMfLH9Jx7aiIOzHt0lkDDe4tP8Ql
ZAPF5MR3t+jTSWMZ9e7bDy3nC2ZiljS18XxqF6hxm06HaGY1uyGQCcGoSSVCxHdF
oQPOOVXaK2YvK9Mjl8G+vZNfG3WJDB13PT/du3owOrDPr+0rnAX6MTcOGIU0clOH
qMeh7oAsBfr/ioZMZoUqZvRpWR+mbjBj1N/n5RkhjKpm0CWnat2xxcfXIeImOmPa
6xEjivC0OYzgKcG8WhhGjS8bY091wtEmnq7u6TxBq3vT7x/v8EESrPINLy5mSW+C
TyB/hJAOFN8PnH+nsjemcAc3ciQSkbO5EeRQAE4n0lsvj8ruKEErKeL7wypweob2
IwGQTUJkH2vs/GXjyQo9n79k6hN9d1Gn/UnBnz7/C4C8EnNJ6rih/QOSDNR7Z1ga
kNT9mJSMvj91pAi9gxaYHrSPoWxwsTQcycKhqYZoJs8CzLHrCtqzOeQpERhoLL9b
Ik4Ql91QoeYE4HaSn2d0aSoQSk3wuVQ4o5GszS/DnpL/tY1yq2n9vm8dzynRDo8W
peeh6I55IEKEuyR60SVAZTfytNVTnu8q/GwjH0GA9wfR6lpoK9a6ht8x2YB137O0
Z2ZUb0drQNBNUON+3f2rWQedDpsCag5w/3Vnpz0HdyxUiY/emp15rR0/8NE+juIc
Sx8aJVtA6IqK72SpSASejqFgRU/grjMEU1rlBsWpkzmbNzZwpyil+bM3BHXwmAYY
hI+ZDu/LW7zksaGuT8zC6K26C4fP2zxdWL7Jtn3krFANHwbcWLWhwKJ1eZUptjeB
94JXNJfE5zHyIIp3cg/F13978SUnescPdpUnO6trzOp//FUH5YaF+KwJ7SstTsQ9
jZgF5Wui17ew67mhjNv/zKkU6qP+cXnDQxhGE+fCHcO5jq8sy5oOyUyU2qR9Qwbl
YuPOqJOMWt/K5hQHA8kFBCndC/g5DSWxllpl2DdSV5SnOIXChjGLR2Y12BBEj+wB
/dz79Z04y0Vb6+SL7jcYfK468Nh/pr95o4aAIMa1zT+pOiS+DuYnQXN0hLPaTu+a
dZ7P9eTE2+LLchXP3MCKkVmZFwb7o/e5KEha4p3IXphxQrspk/gysy+tdY5cwdhO
fJEMma7Bzy2KAZUxEkmd6sOSR/1V/v4v5Glb1aIqZyuvOHPY++bWjwuREmJ9Ra90
whF8gTI7QQ19SXubEGlYz/gC0EPXc4JW9XgRjSmz4N1W/yaTdcsYiV222Ybj/IgY
bJzsfkT2P1K5IM3PqpFKG3htArkSnYlWDQCvokhvD3EK5dsdUUSY3mahECi2xRsB
Q7dFk5nfRoTxAIFLKNuh3JYCbji0Ddbn5K6nPcs+DS/Kp1f62fs/V78MoqAlWoy/
Zy6wx3zpIghCFwa/Oqo3yKyLTon4ieezQls0S0rZb29zcFvA0yKrlmYJcdJQL71w
z0NbkprQRWGabd1RWA91PC1ghI/2m1VleCWJQ4YjV0dkY15FSyLgYxxyLHYzYbmC
dJYAGZ+5sUPqP+p1pTXi8czdQExwYL9nAL0FI/bzP9mgYlw2h3ArBC+Buyk2J7KZ
KJGvftxkFRvsYAMBdeACHM6uuWi1LVW8FxJYeZMEJTEkjAPi94YnxDRcepIZqHZA
QjsNUdZAvR+st1tM7P39xr1mKFXpL2VrcrASY3z1vxN+elolDuGGD6p0jeukDp6F
wpnR5hxnBZ7xCQwigI/lwm02mEkwYVwKVJtlvROnAaneSciJu0nMGu8SPF0NlHQA
3rSZW2bTecb9KG6AmLyz4GQ8w/hSpJHC6Y3CPWMynRXR/57MWkUjRP1f0wu4kBW6
KDoOEV/UuX8SuBmLirxdLtvn1+7Q3ItFilbhw3U7lgubTuFcPuGXIvYMO95k4HUy
x31GJl1D65pKiqW1QCRyFuBWgk+MU6mJUHKutWl1Sqm+eg/wiGAT70s00YJFtX6u
dst0nSfRXDfuEww3S0gDN5TU91P+wRWxzVQ5rF2o5MaIWYQ8GLV7QMI5EjPUKzdA
SNzG0UiedmPzzQi1qZV8Ak6gLudau5ZciOOY9uqF6cLnc3depeeEgGsCYrr5G1BN
iAm+ilOMU8gqVTHA2C5d7LZPa+Zm7SAFS0fbzgVg2i4B07qFns7tZae1rEcP9ctJ
YTwMp4LZA17+xd34SOhxb8g4KHNOj8ed08FCp/9VGbRIU/hxueaghv8Vn60eTsxL
Xa3B1f4+/YiYL0IyqLdFAogMsJwZMoMP3VQJzAetv+Vu7PTm9LCEB1ZdWA9WMT9T
qHTRJrJPrLqFWgdiEpqiM0t+bdVtu4IQqwVUcrUOsg1zFO1cDlV57eTkGC9Abf65
yMmW0AwTcZlXaD6BqAwHx/AXD9C+RAtNPHKpYN2hPxJW4pq0M13tCOCBruDbDuDN
BSiwXXV3d6BR+1UwBa0JJ02D3HtzSA9pLwxWWTuEKEu/vlbjwjHr4PlaPEf7HkP3
PwCWEohnVRyg2qPwElZ2JryYpNk5HX4y7DOfzW11GYTgvCpz1bwdQysEUOkVASqe
mLrAtw1WMo2n7dWJYHsU89MzSLwKS7QsePZGXEgJfjimFyX7rMmFWZ9M1v1d+KS4
ySb+2bqt2f8R1W+fuKPgXJUgcJpSq7sLGTjte5p/YgrU2kYfSNNBJge3od0EhC6H
AVn/azxM3f4awRkhL0MPON+eiy12U3YrGBzi6DJr02usZ8pFM7oS57jodgaDlVle
gKzw7E6v0hNgk4ep0Oo6nO5GpOaB5YtKAYI13f7n4Ynzuyp09WOvJJSloDvjzeKr
1mFo89hP5+Qfv1lQpxOY+uRLaVHmzIRq/lMhYHYuirsGG2R/zUu6fuj69bPZourF
P0gDUc9P+Vvt33EAAEbDxSQ5Kadb8ZBS2wthELBrpN0Sxszsa1V2LYKQ6ayZMbfz
n5Yn9yT3S6c8AqzNeQngwt02Sb1hIp37xbFmmavWWBM/CsvmVw3Y34KmYet6kAbi
PaPAvns5CSMYAfYU7uK16JEUNvYYs22XYyM4pe2nq9JtTlv/BTdHBnmhEq3pYBSZ
dRBllo2GfoSY2aEtRdDooIjkDcrtf0r171sn4lwFKHWfTF9r81IMoF/sFaXs5GeJ
huBRozTrKt1urX1oTYC3AJIMfIzqI8c4PIcSCk2kqHJMzlk5WXngVdt/kWt6Sa5s
m++cYLewGF/7EfWOcJWCDQxK0RlW97W4bz8OpIDSalXDV/T6JryKQZ+oeLPQVrfJ
jx5Dn96fpuyYdirXXsEcUSTPeaj5uC7wDokuQDCA6uSqIvGgRqSIFy5eE5saM6z6
T36xsPc5hthRhkYxAa1n7u7+pgAKGAFHC7UaexJbZt+NDKvfCq9HA98RYCeDiBBi
i/QILWW6wX3RLLOrI8JuipD4aOKmQZOk7IxkGXIOz4gZ/ZiS0DYFUQDmzZ7o+msb
zI4xQrF+LgABxHiQWOhL5wDXMLhb4F5+6oLJZ2sVuWJOn/g+P+Fxq2k6fohLt+xo
svJ4nXIQZziccs/wQOkjxZJJMU7t5zbnIoUKK2pZ5aQCyMMQf1CRBrisMiuemvqt
haReqmwNcFgfr9BTi7aUU/QYHVzzl1RGzeAc37mow/MLVIprguvO0VZWgWjCWdPD
1YCqCJBsZIi1WlGyhojLNK+hSGVvMWFe7xkhkx/Er+LSjZe+RaSxeBDrk5tCtw4k
RpPIf5jLCPHcczPsgWibqKFkOH+0zkK6sqFTPrkr0c9yTha0hgFb3sPHAGLKM3PJ
+qU8/j4FnrJfV9SLD56icG142PvYKfTTY2XLDm/voCdpjYfG3XVXtl+ndH/QqSm4
WnB3Ohtyf9LC47mWHVWXSJ1uy8YW0vkCcITzRLWKmiXwV+WHebrHxoAQI90cB6bs
lxR3G9kI+I537vY+6Lp9WYjsN4sRUi/GNI4FjvSnwv1rru/MHY0+2OMS1LbfiSTB
yeKTBBCBBWa4wsWcoff9gvl4WfnqFfOds+xKQAc6+Uois85k+NwCSQUqODoXAZBk
gMt5XSFlhtocU/N/J3bYc100gRqwxyDDSJzG4eqjT5g1rpq8YF3uORfdWHt4z/PI
vlX06KRQQ398jue7y1jLKGlUbyfZm0vVNLd7Z5ygyqIQ5esuPKxi1xHzC5srKkNE
FgIz1PHhJ6BL36/kIhadbrpYtX7ZD0H9ng0HSjiMSDoRLejZ8VAOgaRYWlfyx9Nf
2gniIQ8gIPfvoL5mN5xrX6p46ck4cbpPeu3+I4M7BhR+m6pr7jWF5qvxV+YJOMNS
tpHOGm8tg7RftRL/j/r/8GuIhwPUqtk2hqT6ubISnvRcO3OjpjEXNZcDAyyl1IRk
XxBy3y1Z/z3GyPDVFkYs6RkobakjldMwH/zrUsr8JCDGaK0TqEYUStrUoOjbp0un
8WqTbUHm5jFv4ItCEUF4RqLv4HTJgwAfHrmsiq/jw0gJbU8iWDUadyycrUUq9SGi
oL+LVos13faqoe2U8f4HFRN4nkAtDGKv1l360bOEjAEXU39IV64pQq6mK0DezS6s
TQOO05EID/jKycMPo0ERM44ltL9pwUWNMrSXyGf5eKg8obOaNl2zZzKM37KmoUFb
7xwR805+uaYQZXUI0+9fUqBQh4O6SUT2fi0jVccYg4TV9ut/LSujKzU7YCDiYmg8
GmKzSJ+1BYUOV1Qw73mXsgZ/o6b8+GLKqBEUF9ci5lQUzxF1iUeFhgXfDa5ea0D7
9dXNnRJ4omKp0nGfXp2TaoLSITvBVVO23zlLusaNJmLCzLCV6LZYAz582ggE+jjp
MxRTQl5JjOxAT1XaRYew+xyeJyBblnJG3CL3Ig1kwkwzaKwyG+XJTjh6/mdWV8fu
tO+9SAu5snLAqsq/mpzOUfNqG9M+N35dxX9X6q9XcWtinQAimwNEMhXhZahsE6IT
Wl2OzPhz5U6kDb2PG+BYvhBijzjMATvaB8KOYv1atZExnvAkXkZEsdwhztdpQMJl
5VB6WVzS+w9aG83jYpoQeyDKpIE/t089l+oWwn/n7RbVEwDURG1ZhKFKqRSAjsaP
d6cGI5oNMn5dOxXwOKTtAiCuskxACE9VWFfBHYQhD4RrbkQsW4viyVtgO6CnS1gb
kNEcnljus/BWrj3LXQ+UQMOecsUKft6R9UzN3pO4qiK8M1hbl68Mrp8YCWkoELRG
k2Z+1KISoUYJQ0B1oKbv/TW7SrQYlZuzp5zTXykudtruKvFwb+pKxrR+73VHH1uP
YrsL0kIPCk4xE8lqVuFxrvSesGRzwcnwGC7sXke0dVSU/TEri6+GCqthWFufl4OQ
5U9044DFBQ5+Y36FtFvAxU4Q5C0gB3Rhgr5F0DGiNFQey2K1p9nIgW1rK6HSaPp2
kejM1AWq6ogfNY1J3i80oGjZsph9OpC+RPK2CWbnyHW8/I8ZniXqSkE67nDGd2ir
wVqjcTYeJLkiHRtrALtuE7dA0YaPdWLNsDgejrvS9Yfb+XP6R74m43Aqr4KnKD4K
SscY7W9mkiFZtLU5uBfpk2W7RNLH1VmacGenj3OvcjEOUKOnOwdCYYzCTVK0UPVW
xIry7+mRvojW5oG8cvn9xc2AeVOqqGc52sGRZh2/Y1kbOLzIJO/lyK+aF3NcktaN
M2WLQPX7HxjW89C4hTDd/IFRdXdzIgkzxhwwvn/TrLSN8X7bvovVGMOF2U4o8zmE
y/gEs7o4vX5K295dXizx8dE+RXFk9fmZ8Un1c4vzjpbqqS4VazlHia3m2lDbYGf2
8KNlTb2To5PgX1nzcasnws0lexy6ed4bdqzIHEZBlGuKIKzu+BSeb1yIBgI2p23B
kvVsaAmIGmZ9M4koltqSB8D2RLUwd7lHH41KOPUij1ZCJlouSr61CVKc3nSSS8K7
er6Sxgnxcf+ztJ+CSXMwrXdFMgGdQ7Xu3a9HrXV7/TSVCeSpG1JxTo4GG2F2ZjqI
Aj4hnLNQi3EVqIJEBzZdlK8/KK4H4onJ7Vl2Ab7W1slJfuuI2Gw1sSCTDD3SpNth
yzdpqM4WQ9YjaQQSXyPrVpFS++S5WWjNX3ATatvXnyXI932ePrsEB5VebEvjFR+p
WQLvSbhQ2Pl226GmxaFD64BK0GSAhjfpzblOhiU3f02e7s+9aNdjhr3MgPER+d1C
wj+tat14XtLxEmnEjkm93TsIhlsgM4aZI6ZFrw1wX7qEO90gJB0vYbtTbNJfQXR6
o0QdvkpmimZZAyfvuotioFvSSm8UABSr3B94WhpexHLgXfTZGlKtVSejAwBcBGo0
C/8PohkxZgRhE68uJbpBAnzbvQd1tVSZM2FPacEAueHdgdMqCPQ5XopkmGoxWGHO
FRIn+G4zk891aD9grm1RYfvOiwq8FCad0ILctjx6vF/k5h2yoEOUMIqdoqWx47TZ
Vf05koEvatHqTSjE0kizA7SPcIGdJx6Ks2CSW6s7rOTf5CmaaYGmMVgPF9e0OnbX
V3l5nuLygyWsBg8JmVfAExDxWLm0CbPL6Q/MhQh6INsFvnKD6t47RPzmYEzf/256
tImN0V6oZs/r4MUQFGD4pMHH4CmCnE6BYTHQc6pUVvukwEb61DraGYBqkkqFyA7p
DSwPHPe4L1RvnrB5vtZ/0cXpt7jCSFX4Fj/fEi3RvodpkZWlp4yiS7X8+IFBdy3J
foz21kWLKMVRD1kRhTeNBcgJGfAyZMEwfr30zPJ7m1jICAhgF8RCdvFTo/6Sd8xv
GEFt3ny2xsDLY5HGtH1b8HDH63U/oc57xxgBkTaSwF/1Gp/LJgesOVDCpTBFvgxY
CQpVxaGOl+b6wT4ntIJ/C6clORLge0ERN98rqMWN0P/P3vPEkx48eanSu+ppXAYw
42t0Tq/hP+tqQlD5ZJAVRQhdC2aiZRRhEoMBHfMLj91kOESDxLzpc3er4fwVXKD1
yEAKPk5kq9bQFLdqdwC1yp18uJ64KobApmtwaGE6k4sfCdgeSoOzULwbBVtY7Yso
f2706y5l+PAS4Fwg10c+xpuRvEorlx0rQ6uZ9x5pvL+UKlQEKRVFmB0ApKVqPfYj
8m/0Z/u2WChACkiGPqI0sbEzAZZZcN0mfpqmKdFdlyJF7vZCiBw832kMeALLwOX+
DWj9hvgFsonp+z/EW1CefgsbLrKQmFw63vBOokWUpumHW/DzfE3NA0ZdpeY2AHmr
CXN67jfk8b2e6tdhewlcdd9ecIczuKapM5J6Ihb3paaaVopPE7R7IvJ0+GnqVKTj
fsmw0H2Qkf9qxH1eFu3HMPAm+myUPR2HCgv50rLiN2Ibz29ivuktGMShYDZnPWw6
bX0zMM5CEX92Rdq3mIkUG81GereVcNq2fiDmsUAi/NnD8iycmsfQxlKIZ1M9zA4W
HKwPxJCuHtazrbDTHZNBgJAbUs/CxH33dtsI7cTLS4ruDTWurHrRGv1fEmd3wUKD
fhcYdx4howKeTJWpXVLInue5f0OsVrkeWt34Xq09SKSnK2dGC++icw6hUI3R7atE
fynNdOKkEiODp1FdSuzrtkWgZYjG0FD4I6YAN/Y2PqwBj4S+zWKnCDtLrVJUrMUY
5pfkhyNc3PSdjYdXp611crZ3QLF9FzzDfSkcWRH+knYx7uyqfSC9D6mot+NTekTn
a2mfVsdE6oaYk5CMueI8iilwkgerJmqExklO4NI3QvH3dGeB9ONKuEHQwgsr/37F
fDzlrYc6CjX/2Xe3Bd0v1zO+AA+DuwKbR3k5lHD2NxQtaqzew5fTtyVfDtRHPyts
zJ792mikiGSNnB66Fu7g28z6vCBTYZhIxNqz7O8qQ1Qr/Ia1LKx9N1Lbx+KrB/Ru
q/l0zq2qdaSdqtqZWHVXZ8UDRe4hY1GI5IDHL8qvGAW6pIVNO3rO0V/yxA/zma0U
sGsYm8haj693LZGWyacXJH27lUGuglEE0w0v+m8qy9xY5+I34efYbd44tVO/rY5B
VR7B3aYcdrAEt9VxD94iMPIRY8fExm3CngFq+cG81+pZWT2ofTXcnS5Q+IIOIpH7
MYaCMTMl6TUtc19s2fFruFFHGRoR6V3mSzat4fYhqlIPJc1cnNkPvYr083i0ZxFG
7huhcZNhSYT4W0fSeib15N9JMS8F2u4hcMqaTNDNCQb1LR67XlJOZ1i+m3hPLodD
f7R9B+rSSBw5F7hLnsjMExvdrSbBt0zAaPV/SoeDpNGySEUXk49SwOSxm3oCiAfN
xFBHhXHy4e9oRY6CFrr7/4j5xZhhZafbJi7wRklSCNz6XrpbLDAGAYL0tc4dwxPL
Y3bIs/SNGx5awom7PGQ8Yi7EO/aieeVNAiTvYhJ6H8vjKmZfX0McwQ6MyxfkLC2M
d3lFb6RcmZAthH8HS9HN9Ueg0sAkmq41MhRQp1s0OTgV9dDclaKPreUKH/MYRRcc
iIHk7ieqWmEFlz1IqoXg+Vwj2eUHRwHSrx44zfPYAzGk/YfAPOXovme/Cvq8Ir9z
dsA1keqwRYl70OmZ+3gu29bZncsnW2vh5b2gioWuuw6jEA2H5YU1/c+KG2oZc3i+
NpiqV7lXVOv9tfnAT68R8NP47zmtFdnWq2ALUp+lQ1Hztskhj5fQ3QaSPqV0jB0M
mzUukhuoPpGQmbpkmpJSzeF1/w9SNegjoxKkF5LkabePkNmy4zH6uzQMx1aTjVA4
LaMkrNV5A5aekQAhswyunP5X8FtqNcX6s+YdDksUXd1NVFL8W6/kJF2kLp9zB1Mj
XIjCjfyQu8xInAnvMfF1zu/76eLZEAU1sKqF4QFDW2LYbFVqvBLCJWEagRqHLd91
hB/qfntoKm3tHUQOjykZCfjxpn+yYahTcEFV7Xi5l2SUO1JfI3+TnUFyG4wOI8eT
Pxr2YFbuh5lYGp2+wXeNoCVsjM+CdeShsEZRmP6/2pwsafzfLYvglC142NJlom4b
LZcD+Ex4jb49rqhhCurFA0C+LjYVmNyenPuffiPlGcNPVjMGTvyFZtG0J1Qw3j+E
c74Dq3TN204s6BBtvrfaBwGH27iNiNzvnM9jLZbto8DjC19v5dEa8Amqz+1bc05L
G1QsYK9BYS/tqLD8zoFNrfF+oYWsTSfePZdZV9qfm9fVS9/+Xnl4/GKY91rt6ite
w3SV5cWKcJ5EIOugC+6jJT9RoYRsQ1rmCqMMcB2lmrH3MrC1HCNeaNu6OkWvajOl
SdMXaalIuwcp22eJKZzSH9cN18T4y4ZHRVO5BBaLdmUOMx1dnwQ2/LSROnI3gdEp
DVHZxK/Zv41mI8VbXFXVDslC6FZcM92ZJTUvlsqgMgwHsNiV8Tb3jOQcNtlSbHTe
xSTS9H47Xtco8oWQIL5xDPEo4mMPYrM117Tnv+9XZlWpBaivHIJiRUyAoCNQUy12
oMAJCI28gJKDEBYnLdE6JUBf7THHOKLVvZAGIQ8Xmc9FecIIDEhZPOg1e1P9IgNb
sJKpAbsOgGD4A7Wf7L+OIS9pEIxaJiASoVwq3E2NxuFCx45oTNR5pNH0EBmzQLFl
mn+iTjIDg9FpuGMzESxyA3Nt3JnJGmxwrVAfXtpHfvzByxVWLiX9qas/jBrnAT+S
eSsP6ywT+yBcpYYOUYOgMJgFk9o3PTv/zOKN1Pa/BkuFbImHNoieN1UaMRfWbJIc
5YpC0dbesKomL6CpUDYdQJ454Jl9zViI3Ky+EUBh3dziIIB3k0+k8iqk2y0z02kh
4w9+uuPWbQeSheSL0RCHqzzJZZt7HAudrQ0XdVTI+/sGjfgHC8MuzJbfGsR6pUZK
MQZXU7BseZp6E+M0xtSNDD9m7gpFDwIwNHnYsUHyxF6WtUy5NHMMz5BFiFhrO6NW
zg+LFx3V0eWCPHaT5EYev7/a25mBCyI0j1LpaJXD8HPaXpFIXpnKgKmxVdwGruZy
hzCvm2cXjBgEsXX5N0uDU9ayY6kpyxyy+jbkK6n4GwE0WOhABY59O6mir4yZO9H1
m7VVX7sM++21RT2BKjbpbALCuCJSbVBAgQenXSVzdhCnZ00smKMZYLNyMN1rY0UE
PepFQODsncvPUDem42NpE7K3cHwkl2vRpDzpXud8Xv0UGstTMn7rTy2V00ypdpIv
S4PDOEMc4yPHybAcRNVw1nhbOizeDqsaLhejvPA24wfN9loazn1JmOWqXqScRuuE
GkZWQZbF9LKbbg1MJnVxXvH/bMpPYfQqZQqY40b/8wdHc3k0Yi8MLuQBbTX4NxQk
AwIXCCPhQaWpv9kCX1x2AEqQYblRww3WTSsr5idYc8VuiVhU8nKO0sHV2mvWp8Kq
cN5KYg44h5rI2ZnGVvaw4myi178aJ/6w5lrSEAbp9zSXAtDIygV0+azDM5hJIja/
xtk9kYQQmIFX47gQ4XgMRTAvGI9s5foTOCk03IqoR1wYdhmAQRRYksuc0a9LE1Ns
tF6dW+Vvzngb9xbUOjhhUNH5cdN4YmBEilUHxr1TbKsq/0DCePRLAeywllme1UY2
Zv038Y4OZpKkWPwzlmfotyE0yN81vlFkRSGOoZTV6FEJtT6oMF4flCn1o/hPYeiI
tVTYFRcDxtb7wGX1yIbPGr5N1oZngjXb8YQRuqkNgcDZVtds0JOQ39Q7FWUDvujM
7ZlKRnwZutwtDHp7i2snsLxyzsUGQ2t4+Y5Hs66J15zHVj329Hni4HlG72JbxZXd
BsZBPQvVNgFSEvVnN3qAkF0H/cu7J+L293ApJ5C2J8uuic1jfAP3B+PGCbV7G2wm
viqPS1oqCzhucZEpqBCy2kq8RSUjGmweHSH0SHqiEH0/bIAytjYKAXGe40aTQSvi
wzbz3dGT/5aV1LkKL2xpR93qVC4a6cJEpFiAq6A4+Z5Acg3K5603Kxrvj87uC8ky
Qxb191K9EesKZBthXtoYh92Zuu0U9+LujjxxdFR4bFFWuWkvswh6K9haOA2FOVVN
/Hrm/cpVgSzvASPD+SLfZljNSpKGfyhAGa8UWdV51OcEZugFqjtVpM/xGUqV+R6W
l27w/9dhRbfVOHj8gIW/4B/Ci3gnZu9sUNcIpiSoJQymRB3VCEbSpkZ8AKswkQni
gkoCRTZ9JWBQ1AxBD0e6REjxtSwXebmK12grGANSO+Aduhz4AmnxRorVWcYK3Q96
bCv/ErfBnHXUQ4RgeUds4reh5mjSAUc6d2223IYbWUxMn4DBDn/Mo8Uo+TCzZn5Y
IjszrVzpcHiOOU3Te1eJ0xS7Ov+HVubTJQ1Uv2mozBKFaBLXwveR3Y7N+yaH5/L3
vYN3OrVW+Ju4DB665tApZq6JVO1a1XIPq0cOqsEWO7RQXV9MMBG9QjkNFKS6ltEI
8+lQbd+tNWJ8BacgTfmE8xMkKLZxT4zFfRf2PuTIorBC9iLuVBKfGYMK01RUvAvf
kD/Y/RsrTjb5Ul+ze6cGFK2CDXGKX4uYE5VGlrkoJA6FmwCEuDyPZXEdQoRUUN8D
0l/KFZYAgSTGh/0TNcpREaNv2ulo5u0zNXHvyE50av7WXuYMsAbkJivospKAu6/C
P+iHhvtn/BWFaZurEO/Vn4G1jjFYJcw7z9tj9b4uOWDr4+tXz+wQuLINQofi1dPr
2e3ziBFo9uMJTyX2Gx5CPqO9wKBBPtd7mCyL2fdqJecp9fBahQtwQcKbjP1YHd6Q
yLXPedHRnADjNmnq5YpD0KK03l1PGmwXnHlkRjD7BR1jLqfKTT1U7sAPytOUveRC
Nl7Xb2Tt0J/XO6nSqO8+VTJ8z2gsFXaX08yyIBYL0A/BvkAqlo+GP/xiVBR1C5uD
H5bNdb/LiLYK9gkkaTI847wHbWVs14fKbLEKH1hCzBPRKDw4D7SGTpvwkKgdjhE3
thfidy1RFUuBBdL42XQgsCoUpxb0OHlVXM7FMr4P7LUv7+W+AebG1/ylBQ9EOg+J
n0dwewMJrkrWRWaOX5scuhdGAP8JnS7rjZHofodHEySOYUc+UjiQ6+gR3AelIYiX
0SHM2/Ed9kCZEvsuvTzNmCWL/diQflGxFhUmvs9/tUnsE4bDWVM7WqhXVVWN7pRU
NjXJrM0l85GLxL0bYqbqXAjiZWTGZYGFxSv0DeKngG14V3eLYYkcbnFgE61fQdvG
PA9cKG7uLhAuXKulm/fSXtmkgSu1C4J3Sb8I6aljy7VWPtab8fsnayqB16JfRwTD
AAbjAvhqhHsjsyf+hWwMNK/hioYPVCjRDpGXbIDkJ1bM9/LfrGkfIEWsVU2TmdtZ
VZ2ASPG9jtkIp4Aw12vGda8qibAaBy9hKi2MmnYMQlDh9W8nw5TCBKs9UjAsjwVG
sWNZYgTAgr2vVuvSL8lUUZb+ypvQEWkevHul2TkjrHok165oxXzpunrrtxxzCbHP
aMza3GTB6EY2ikVJolhDV1zjKy1tvw8QiuGYS7SPiWm99Wb3VuXb5hJhE8dXq53C
hDWP8NgIWnvrcLcOIZ/A0lJnhZLOulHbLxyog0QDS2hNX7ZDFsszsxSvRDNJaWfb
4zrD3a92xZT27mdl8CbawRvoGYNs/OBvZW2A2FU4F2j19XYuPE9heMyHu9QFd16u
SA8pPFzQOkP/55XY0TjMT/cW3rbtIavlBwLsJW7KXJIdmoJ4UIpuXThrUf4gM048
8d+i/jLBS42gtoP2vT/gON6Fx1vD1lyt6aauAQMcr82ZdOQFtZ/GrgBtktZfNOH4
Sefl9EUf0ZVhqgn0OLQh1/tLMNvqZQZB8zI+/ogv7h6jbdLsdels7mCBAsj4tW+g
KrBTpYgHiyNr35S7JaWVuuRzCH8Y4noofpEk0nr40aK1QoiMG2A3TfIk0kktdSF7
VGJ6+3dkNRyPwTjS7PtnG+fHw1fVCBtB89uYcuPIgLW27AyYbzBRK+3e+mlCTQMT
7pCeBkdkH9C1N6FQMrcytBFfF8MFDbgKuif6N/G2eigpl2gDhF4JO4jUIONfEI89
VR7J6tGynwKR84KxOm7EyNJ/jGLUQ5uu1VjMQXx/kIzmXrosVC6867Z/1bsEaBja
j57qspanNewcl3uJ4voGQgjoiEYRH82pSPaU2I8y4CotwSDumCMU2Bpfysjx7p6d
PkELFMzVBcnqc69IV4FZzd6RTZu93n+CsnFV1XLsnrEdrRwQSQ0bHZ/XvI8eR1rX
wg8f5vtvPso7sbegw9nvqa2Y1D4PwvdAZf/5Lx+43GnEmvaewtNv6bdSkqZff3sk
I+OMdoOLNrccRN/lAZ6Tdl7y7rTysMb5ZddvDT/7r1OMPbk6U8aggLp4Pa+VGjUx
B/e5mCAJ/3fyebqYs2fCtDPIQ+V+ZV4ECd27WrKHaVonqv0ubLc7InZuZWcxs7ri
LxscJ5JhRQX4JZLpUTDXKXPXQSrYds4RlBCf66CYoSAJyUduikt6pVWHHo5RCjor
+YvK1l6BMtbQHm+306PpFK8AvKwXoyzpSEgm7YRpIJvRMGoMAWPKwSe1ixyFQky6
GOtJsooc7kdfx0o5hnJOSRQzET2dsjxOujq1hDU1gWQ9OuhDwvEVOiBt94u3mn1x
oA9rjidQDMXlzPcUzhR8Zpc3VbHDVbgscj3tQxfuj3uEqhqNhgc/FivrlT+/BP3Y
IkaOfTTeSWk79uTSuwMOMfaLbXeQyljWFYoW5dWMD0tnCfdcODrnOOaSi938jeXZ
xi8YxfmnTNQ26Q7ee9TXpCERqcKurPF2csu4OXlPTWlNUpUDItq2M7skC1Hvplfb
uxCvy/lC1ONL6eBbqmvDYTfwknJiYu8qTVndGCmY2IiPUQFfCc4DT7aD6/nPdTZK
Y4i7y1+f5Ot9nxJJZf/+YfcsRkkbJprFa9dOcdbBRQQUlIZ/KpdVx1KSlrcsO15f
S6c5ShcFYjsinQto/599aXkERDB75GaiTrgOYxp33zMmys1I7Pd3+QLL9Vsyv8xQ
Rs9moQFbnuGhsLueCguuRkKPZNhswdqua7Y9D8flp3Xg9Un2ZZWGx+1eFzRB4a2L
f5sNR20SUVXJK+mH35gQT72xTwD+jyB4V3dFBrYMJ24V0rKlWzlt0W8U0J1yBg+V
+oP6GE2cLy2G86Rt9mNhFwXdYUSmYSFu0mlTGcbVtPRf0HeEE3qYk2gxmGeC94AI
QKxn2lGy9OMqcPwH6+hqjHLJ7ooSfFX9z8XO7Ip9jZ8Ka9VE8W6x8+ga4meMq1Is
cGmYJtw+TSBdXouwq8K2p8vInXxy26B1NvZa0c3svZMcp3WQAe4SDRdxpMLSFIT7
vRSQcTgfEt8JL1uszgB+eNr91+LAbrsSKlsuWcjPEzKgeiOTmdzpvt65hgF/rsu9
uIR+cfOhCiXcnVRpZCEWu4PCCmSFcwMk2qv3Imzgz2TReeZB9FGKbn4xnYq5fa43
ubhzh7gM5n72/jS7+nXe3aiDg/rkNrxeF3elhoe5CD7uevxiJr1OMohAZEcSDrKn
Vkyz++vEU6lN6Ja/FvG+KpnhBzdzIT1neL6/rQe94QHZRBjuJFMoUSt+Dg7n+YUH
z/GWs0ZklwxLZc+8lvs2yK18m3tZFSmzrBdT6VpVA8iEozm/QxkEX9MgNgIKyUGi
ln9GS/d1BjRo2qz5iASFutYPmaP9d5pvbC4KjkdW/WFYc3YievB2+VLtFZuecKwc
AysZ/U+xojx7EkCG7YufMlOd3sj1zWZ0bGqvQf+0UN13PjfBRnmXprPyDMhVrU5V
i9IreGZR4zo/JMOILHnh6vRgEun3n8T1BRsRwBOcH5z5fXr5g+cXN09+mQLlbDZj
S6MrZfaSWIJkdBWgcRxEmSfnMa+knuolKqfljFhtW+NluEb4P9oBvgT+HrPgJB6I
AlaQq+dbXpiEm/JFz7PEkKFHlaHAEULjUeqEiglP+UiQog44PpsMBk6A2DMxmKiU
Ra9fiaIYElb6AcbkXaJ4WNByxqU+gLUmrLF6IORdD5vAeNmlQOo2o/hiD1wPerHZ
YDi/Vo65dld0DwTyE0jX564SCA5D+gg9tpM3UuGeU6SY//Y0Um8hHviOstQRK4sy
UQV4ZHWSS7lTwFIYXepziX3jKgvj/P4RL4Zp/4aZIKTvAOPQ7++xzxy+2Eohrg3p
TcVRwj/+XvIRB+atYafhTuIA1wnZKHvtne/kM5kF/7r/97mhxzQUATeLX3FQgQPY
e7yuNlCEsaSmB+u/I/lS6LLergK9KlRVw6CtLpVUVreBSwk4a/rAwEAXOf35D37t
UeG/llxGckmL/9yj9IAoCeCmN54yJ3ER/2ZSeCMgF5OJEl+kgF7CA8I1m/RnOlDh
K/2nYpR0jvRHjExhtzwvK0H0lM0bZuWs5aTUd7071CtCfBVWWvsKueOQSi5oq+0y
JHY9bwavjFLAD2vuiLnoecrmpRIjL2BVx6y07RAdPhphPDcUnAkwroO0IgAywHf/
WWm/L4Gj8cUksxIlNGzKDWI22lxopqMZUCQ5PAO/ZOKL6FxE7yAv3il+Qu9gSE6j
I/Fe0c7i16QSEJfcANjHlDhsW3pG7n7v8464Wo8epHWkTX+sXhZC4NG3uHoSqBh1
ha7YKuLoJtFOQYY6rSqMD5/LRcTkpki0Rca0uRcU1yjlBYeVY0HreWZ9VrEP3+N4
k4+pZWVYgBe3qh8DMhQuVQJo77uW0/W4USuJH5gSiYmzaUeVn7CxjvLajtZKDoa0
FVt9DOB7AXsbpaJDoYRh/AzH3r/3vctRAcWf79h15a9TKl9V/O1HYmKTAtLoCg6E
W8oZmUhcKGyJ1rzjtKaM2Br693E1QIBRWIL19XilEL7MmDHZWF6cfPPAZI50TDU/
zjm9rfJ0ztKIej2dtR8beu60qp/TmPFHHzfrXvSh7A3XyzrhxOfA3aeBHejU1ggR
PoIlBDz5RTak9ZaVUtDRgD/4WMOkoYRBkJoW9U9WDq/f9BTn+v9EmyYkhT8PJQxh
MbfzPo0MVW0nqJqT3s1dwUwUL8V17r95IOVVenStfg+OVL3KAK66oqbHAyPvGmVr
6UIj49+1yuq+LZ0XDiM5kCqFNJc8d8XSA6FaiZ86JI92cwyON1SddmYQPe1CpzQA
6yna2EquU51Z3e15bkW5kQ3RSCzbNvDT8zFhJoGByJ/yYnG9xny08FGoxxnI2dec
9otZa6GPFv8zirtv3LJB/qlhCM8pt14BO/KsbiGhggx7XnJJpifcwVBXjRQqVZwW
1IEQbOw7sF/mZP4qHi6jKxk2AZRJ0N6FhIqKarKg6BneqROoNlWFxb5lqk5ZY05t
VWx7Ed2tGg69zTw7cN76AZHDs28x7R8yBPVfmEupbQRzYll+HO4OV+3Sqm4eajYv
ZDO9BYsbHgs4qQglOdNyX94BfyUGbGdq9psKJRzu+nfaEuy0KXc6C5c2nyUNDUUS
sPkL7hoZtT9dCZElfYPB+5Mp8c5PFivSoNA+nNbnuViu2pO0ZKqxiWY5+oO0Pwm3
ybPUoCeOA3Gu7g8b4N7wg048/3VWgw8wITRfxKHFOjP2kgebaBzHlO9w/mCxnb0H
D4foqAmzCvik3zldMZCyn3xH4IPCbIS6bkxQdfFQhNwKT3gl6t2NWLALXscRh1RB
ePxbIq0LYmlRjkVmysNGg5UBsZS9N+Zfpxa/GIXbd6+eq1pJZeno6Ap/wDFhQXCP
WnbEjnZnJXDmBEcnd222sHOLdjJXjfmdLxdB+uj4vdxnsUaQHcZ4WGz14BxwlMgj
akt8r69py2pVi5RlyYetkmR9M0VoMF1BN8zYtnPLh7521NZ8ORT1cFrB41xc1U6t
+L5tiD6rsoREkY4FKUIlmRcVAQMzwQfeHtoqc5kdVmPTi4Ct9iOW8sYSC+fM6trN
Ffp+aVvdi6gYBWs1AFwJ7Wa+8Zk9OAZmOJHTi+uo/rqJULur3koDfxSlX3VorCfa
wDxtbkYmKV3RTgX0EMPS1+7DJOYNq/i0zVGwPvXZVADMUTJtaxCeSpC0FsORsR+Z
ZlN52NTLrbGO5tfV6dfV1oq2LpPoX4aepwUZPeWpgfqj0TPdxvqtYVoGhNN8Z11l
p8vpvV15EXOwKQqqvdSWAPuJxV9WlKoxQ/PCYcexaqzgGIiEPDi60YDOa1JJfulv
gUJvuSdwbxg8jbK6tg5pYLC3t8nU3Y4+aS82BUCWijCvGZJ5ppn3qSDjYjBEm4uI
y0v8PJsISRBC7AJRjWbbsbIuaT4K027ZPJDnHEVOM17ntiqO11Wa3XLmfZfoF0A3
S2B606gIl609D8OIYFDnyDRiSDFTSoOGR+abboRA65Es/mubr0kyAmBBPcHDXVi/
sA9E6ZUPip71mTmng6EkYSvSoYrDqcEL/SjoOOin4kQ7BCJp2DeFDLXnTAw5ZDpt
O/EArceYyJiPUBeuJQ9/MqOweyLcctm5gUlBfVB2KarYdry/RdNAcgnBrPyT2G21
cXo3R1+S4czOD9m8M4JJ4mKsyTHYPC/z6UiV2D+u1dsDFanr9biXh3q9Y8esUo6A
RuJJYKd3cfWvaJ6ow4ByGVEb3lG+NMBxzuPGmJW4sMmpBAp6Reua0rtEcP9S+CaD
g3kJNHmLp6bKZRgS2W1NtTSaDfFgtRxs9tWFY483p7dCMbI4dtwb8c9MpFWTG47x
Z5CuL4GxPGh5MePuAHDz17OoSjn3bFuSiKKyK/t5bgIaEmwHp7pV8M8rzBfFl/GT
rspU0as7p4ptn/5Mq6HhBxL17+5oUiEM0VX5alT0TFlNXcDzKroljwBpDSewISWy
MOdFto8wKRXanBAnd5WR5ge7JVDCarRe+FH2Qkmitq6gJxfdrFW9Lh3mOXHjLVy6
VSm9V5Q2RwUgOXn/sEDbNGcB6OVGNpsVIM0w5Jv/ucdcVNqRrMeo6XLoo+3fpXkm
IuoTj2G+cQuU/01qOYGt4Gjj9fbvHHEt9naHIdO+42pqORtNXl+4lQfondL/4IzG
QeIvGoCRYGzO4BgPaoSozBl6DR6NVyrRzv7sEfZmbvxgEUz/GpDvDHlM3K0INcpg
/NpbKhCem80Wf1l6HjvBDzp3w+HhL52D6z9naBdfAx+ruVUjfmFxe0GFZ6vdzfvM
wTBLcuQ3ZW7ksq5g4uj9lHN0B2SPzrRGbudaLo1bhas1bGSTjSKKV+3K+hAkrT2u
guIHmEiWq9qDLPVmH0gZAIJVjRXASq8vThgvSjXm4p8IEIjQrnHZEn8Fv3OJ4E6D
c4ApPum73u4SW056A5iUZFb7XvxufMy8Udo5FzPGrPkSahq2dtHJyvAMfzBCsEJ+
rUQiXb7RhkigeRVkXh74fIAGhyq2D6WF+qMTgvz6YPwI9K1zUAtS73a3EWIihMAM
zQ9JimBLdpoCgP03sk4m8rxfpNX/z0pIn0vDfQwsrFHIK+gL/rx18gvSAG8Yv7YR
REdyKQ+vsZFLnCvtm0hrwtivkEVafm+eZ7YHwHFdn+AWgQ2WpQ3WsUq7YDHrrm6u
ymd6szbQx5l3YOfRt6V6mPwVP0t25DgsUz5bFsZM1WLu2J5DTX1Zom5DCbVwxosv
G+mspEFTsNHDWg3YakASHaCjFSlkEzHIzOqI8OEaORn2Upm2dFchsmTcYQhLlcDr
TEbIOgJgTemFN2/O7TwcfHGGwQ5w4ftKWU2qt6Pl7tok3w/PE3/57qV1AbXcDBPR
zwwd9b2zcrXBexJyzz0Nf3nW/czFD/tcwBRqJ1u55ypvsjyTC99vMSbCiMf54s1X
wKrfNZgZAq9Uq+IGoR+s3HxAO6/bLNxMHFRhOj3maPe7ZX5AortpBizY3+pW5au6
zgULR2Q72zRWJAt3X67k/9r2bxxf4gViTuKGbllPNiu75Hh8/ivirIvxFY2/lGOp
eeHDESBdGGXNU78bWXdMWXd+vzUdaDVU1WOyv1uJuIyybT0QvGCxlZGs7/15Ti4L
O+0gpiqj9FbJi8oCTMEq+sneSqdbhWdc6bvGZcF5Sceh+lU50gBkETl4CR0HAhQF
zhy32bo677EKDU9taKXRUUPBx/jkQI0WXkTikCoXfFpx0Vk8dZhpcagV8mb8bW09
3qLXPWQwKCNlvlqFoUuzY3T5FWRWx1+SkKGHb6vJSjv7TvkCDu1idV3MSVpxV7hc
hTj3q0xewOza6ncFmUEeigOLOf6gk/V5ZF8AGSGbpgV3JBGN4PVoNG8qop3zJLhk
YKN3Wqd0wMqMo0TqDkvOoGwHQuMydu3vZjnnUhZVn3nIIe43Yn8S0gGqo34m2Ps8
jox9G6wyW4w3Pz34p0Sx2FMyO8q7g7agIHxn3tr5179Zdo0X+TnNhywUt1TDaOzx
OPv9xoY+dN90hWOVeab1HItocF7OyB4CjAlhg9kIHgQsnCU44DzGTBXinTi+e5w4
HuPN5gMx48aKJBj16ylnwLkKmGXxEPvCco8oD+YXHxQ+s3Y2qcZCJS0VeQ/WiLyK
GvgA2ZEF8UJJp3TZychDBq/9XpDAdK7M0pVZlmcCTHeg+2yx77G9Ay29YtEQSZ/u
W2EigSzanSQdKUx4/kCYw+k8q/+a1kwQfWX2qKdns09PKGF4N4venF/Dwgeuy0KN
GJTrmXbXFK+w53wKSRjW8mdSaeXjUONTguXSj6G+RWxJ3hG5OyNzBPco+M8G4giC
+pmZTa0o9nw0LbaL9RmaCZPeSh8crbcJxXha95dILOWOybxvgXi1cndTcW52U0KA
fDYiIybe/xN2I645jhRGHiXSm1Qzb3hdUsFzFPfJnGdTO0xMy55YTkFMo3a1/q5s
JLgxj74JhAxti0tfcPHOP6LJQPUurc7Zbp9WdAQIfrVEcEzxSD1tZsSMc5beYw9G
8FxRgQkaf5unaE/7ZizLuvP1YDX2uBKpZvfr04t7EAQz9WC74c/h1RKmWBv3e2Ht
qvgUUP3ilLlj5cEW2emY+KWbir9Di0WgLdrz6CzcQirO0/3jUVq+D+BakLr8isbr
Jca3NYksTG0EFZ8eJe61km+5hZ6g2MhPSCHIzA5BvAziX59SMcFHh2yS6NAkvtky
4yRoHxSTNsQLuH4S8M8aLoO5MTbhUZvIajZ8bb3F/R2zuJ4heENn6X9IAZy/mpBk
WVeNkW5vZ5o8f1zgdUUaWdnaCnTYGHsBCT/vFeYyTamxIxyOitDF4mXEa7ChjwyH
MgG4c69h1dkr/BMCEO2mWE3eSSXYyJdwyZZHNyNv6qNTKyBPDgDuLKOo5iSqIO1J
gFvxx+6I6B4WJ27QDrQF2qwlq6BUCV9Rnu/0MGgBVGQu+TXgb5zQsHtP1oOzHiCd
u961dOq0+h7n8deQerO9R9IubYb0A7AaJCGS7gtiG0gtyZbYiUYmFeTq1ai4R5ep
/p9hV4kzwuvlPQtph4DWT5yBxiDjCUEeY4D5+aQwAbrpOpDVs/ePh/lBu846th7/
PxcBdQYKy3lt5rt1pYeM0M1sE22f15GLuxTywOfN/61Lp2WyQEqHt7XHAI8M+x7H
8ZjlZ2dpZU4XrHgPIQCNzKfHddNaRwU4BeWZ6B5MdoZ3WW1ydOLp60cixnEUlN2s
jTErs4uJJxTHezRnO6USZlQhUd8l/b5zjGYf144Zy8yMSlDGk/RF7ye/31HhOPqL
H8jggMvOT15rWSMQTxH6LO2SVogwS+0Trx1i62T5QsUKWlGi8Y9j80r4r1eyH4rw
x89fpcEbfDMTUX/+atTx3Z4zBD5XLWbZlccTn8m7tabMwfRij77yPY28l53RqQ+s
7Io4psezh68cym7p6tSmvc+SEG48aOb8nWZ+6G/mMGMrxyMGFvY27rK8Et9A4xFd
BY5byL8a7acQGnix4UEZplPHoJHmTiw86xy8LJRPoXV+r3qdBsR8H1i/L23In8ic
nYuRHRKKZ9Zp36qzTRhuDx5KcrgyUSo7wnkgXfY2q6A1qk89ozG0Cp5roC9SLNp5
t8MtdgkU4TMgC445QlLzthsT9rzQAy3l6mFo5mX4YBKs7u8aGFJST3uJi485Ott3
q9DMzI9SPHbmcgfP/a6zieJMrkgBwx8q/M4BZ3oKlSwtAkcrMivozxpSNiP/JG3w
fFY02nKMhASil964dcx6JtlCzUggpiaGmYz4/Oduf0W3GbJPsd8y2Oic8Hx+n+TW
5amqmx5Rwq8FESuFNrsitDRUMbMpGRHxWx5QDpGhKFUaRS07do8xBDqcv2oGZEsb
6ghuFoY9JarTt60U3ewRKPNXPGmO1uqlMk2eguS+bHaVeBjb5jbS90wRzzecZueI
6LzRom0qdg3kipkKvQo4bfO38cs0E39hk2d+pMvyvrGJpHAl5Oy28Bf1Aggpw4rR
Mwq+fIV0NuYm9h94XRn+0S6wtt8MQ6ySo6nkCF+qI3yoaKo/Zplov0PDf533rdDt
mIimKU5BjMiP8eZza1yZ3joVQuQMryJi7OiiAqmXzMob1RhWOVX+7k/CTheWUPAz
R9gKrzVZB0mpMgddG8FGa49KoU31pQhZ4Y9FeiIim/9tm0KgRIHdnbpG4ihitlXG
MsGvLx1v3ZAY093aSG4fAdlz0ffT9SzZrEdYgDMmiCS5C0sgHBsQKQnvkRHzbR9T
TqrsSRWDm0lH/Al6UwUHA9bHFASgAALfoJd3w6g7NyQB4Z4S3lV9LvSCNg3Cqhm9
jNAVK6zUO8dS/1b0Z5P2D7kVk7Ek2YNNSBmvbEQzATboyWQRLBr4D2KuGWn27pXg
8RnNH88A4tXfw/imZfdHSKYpFuMRhppM2DIuVFKRg1dnLDegWhfcJxExnGxAnUlo
BVuRqKasrz1HsF1sFVh7GLYmgHk5JF1bB/wXhLH+/I9AYYMronUcD76pEvbAfd12
By1aFdapX8Xbo5KyWosxOOflnvrtHnUHcs1jMTrOY1Bn1E5S6N3wNs0Yy/yPGr/9
rGRzAaNkHghoVAb0hfknxxe06SXukscrtRwF960VPtTQ0fZMXvyClJzJJk/Kk/yr
4CMVFumFZPcK5Ejjz2sUUTUEFgUfDpTcFn9swtdY8HLkzufDTVhkFVlhfeQDWZtM
ts72j4hW7p5oJK97SvbXKWyJkFVIpzgXwNHv27wfiJmTWEkSjA/omtVB/lulaA7n
oiiXm2iqR0/lQF6DcJtzvw4qd3Otz8U0qA71pW0IVVafeAVr0UOsQwrs7xPJ/iY0
g6sdGk9EaJGAPRtTpw9l4gnfj6r7nUgtz5qIgjS57twFyKHQ2KTmI3fNQF96M8J/
hpcmUoop04Bxe0igfOhZkyyzweAuO2y4lF4/uM9FV8vbkJuaWPiEb5fj8mFh06pa
4xLcGfKzJCLuRJm+4LWqYISQdwxE5S0tLnd6LCVFaoqKbXteQ4UWe5TJRR2Q0DrQ
WaFpzHw6RjdN/ydgs8zkLJ13WWAem4eLbZIL2siwo0Ntxt8RrifU0FmJm6lY/325
AmQXVNE8yBH/jZPMAefIHuZ2FGB+YFyrXPzlWPI5hACX7LyfGh7Y+LOveaURqCZ/
nqaTOr8TDT+iF0hwWp+GoVotf1JGbnk33H9xCJqGmXNK7FalNRYxUtXuiZkFXXmS
2bdprsATBnyd3+Hkb+8Q0VH6Ybk31MAZKkR/hGTCw3J0jvPEJVQPgMK6frnzjKgP
SMLyJJXa06Q8wYD/sLbH/B3Idgyd8XkcdVoEudFmGReD/LdipXZF/XJZE3zKeKPC
fvYQ2QIU0tJOlAf6/2wD4SoZRgxb94ASmf16hQdRkwwb/eJwqlQEFJ1byLh3YfF0
JYtIlSPcZpWXdDbuUTVvJq9J/jbVVrVImKJSkH6ptFGojyUlL7VoSErAEzKPkPU1
EjYDOVIUxDTvYT0AN/X0Q3LVetUPYZTSXNOJZUgRj9ExpvpuBSkCkEplfJpU9ldZ
CbDijlM+MZYtdvpBmUxdchljRuzQGe0GSX6g6g4CO4rtdiZJW0N1OBPKr3b4tKfw
zufFmZxCz6ueBLCibFSqQJ8Cf3j1W311IrtW65FE+bxuNUXjBI6u0b2IAe9UjfcM
sdt64u60kxLCPHaE9BqrIwLf19eE2kWd1m9RhPFRxXUgudRFYQ62ukQO2pvwyQao
PalZ3X325bh4/p/Llbyp26enmRf7g3EgywMeAIXllC31EBr/QrhODZ6oKLimoM4m
XbyG0orzqIJ8LrRaPVsVz1Zdz5zKMnONqW+KWU3GbisKdCdwJJfZ0tuGZywk5oW2
0TeV/gT2UZLJ3qmuBWUiN4aeHcdhMOZE3Ov//roVEHaECu1uN6cNTpZSIjnMMx8m
OF/96EgkCK/9EmRg4YcLjbrZYQ+1fqyVXYnpwETTtsEepFXR7psFRjpyHpI3S+oQ
0MGulmEnhibbrQQSOlVFRydVWu8p8uTnjmy7R9d7iy+7OjFAujBidYkOdP2zRwsV
dVebmi5/GnB8vSycE2svBIFLZhI8bvYbQdRXFBYXm8SIGVRL5lI1yX79/TU+zGK9
Nx3a6L4zy9PuuX9+ZhijhAvGb61Fg8WK1iiF4pY0AsFKLvXVvOctY1CK60i8IFOx
7a72oJ2v7jzm24jqJAcBkfaHw6dc1aXa4rH1RjWsXF8cU5Ngkoqez1p3zP0IkL3P
CRiE1v/5OTQXgIViH64Ht2rDg8n8qUjrWlPZsrbCWqz0yWRrst10xn8qp3MnRNRa
5T9wUKBUS2YGsBasAcsA+UaZCclmLscYkYYuUyT4uYWgOqXr2t39zn/eSE0XlgCN
CdIqvXzd3fXPRAIkWj/52cgIEzkzfrhwqS6Obt+ol9sxVKnV+mdbE8TrELNVUBnp
R0LYt1v0ivfiJCQZFaqzV5lkJurJZY1uUrwH9GsQqNBfIEMMOLvceSxWI8d/wbJ4
NLtDMlHEQiOqMdoGzrseQw+zgMPAQdh7c3Beilr1kgIGoU15azF5yaW4JjhByA4g
80azsoXjxPhS5+tdTFoIwMMQtjSvc75SgObCCoswc9/ykK/3Kmv+EMsYRSNoRwkx
Jl+P905Tn6CiisQqvXWmlouOfYhqoQpc7G4HhDrxXgSNqzDGvtqxCT3+WlRhBFn1
T93tFwUDYkaEaCl2swf/2x1s5Objt3miNFxuWJYdWJUDfi/EJhx92vkhJWgVRb8o
59fsryBtEgDJi+CMXNZ7c0OouFR09H2j6IVfckWQilAsmbo+YBA8khdspb4VdEzh
1UEI16RUK2B1y10qXmGa5TEu1DdjTfb9r2sSY4lHGUgQCLrqr5p2cKhbazqLcy36
BmJRZEHaH+x1ejA9I8GkyESSsN9Z0fwGNddjKKTY7L++f45/W0RSILI9RSs+Jf5O
Kn+hTME7CvTK89M8GfYN6Zv7zPhr+JLJfG05lyh2cfi639EXTnlQNfW2170kZSoT
1q/hq+ehqKdnFkmXMrN4Oi80UlKqcFOV/I19nqc9M16OP/vQTwVktsQCrfM6MNj5
ne7sPjCVlhlD0ktaJ7SLxRdOhlHeFSIfIjJDNuj9pO9idfGyiMwkRnfSn9fn9Tjo
GtrxnAemu8fbHWuSLXeWpL4AMACrqlAcz0oJmmgEgFdsG8+MVx0J2yXpqEVk7u8s
KIdZ/gH2izsjEIsz3bZq0a5dOo17V/AzX2U0psYcxoN4UVffRog7Nphva9VaqnPj
ouTiyMTo32tTWfPeV9MMvya38aD6SCNu3ZqfFUDGxULuwz/EnF5BkVQxbUj3GSoz
TSZ+TeGbsZ184oGax7Y0zFXbyvJR+E6Mo9Tda3kmytzzPoXAjeIcgfyc6lvZYeiS
6GCMXEmTjjrkXDooSlHMOAjoa+A0BkwyoT5a/Y1/cy6dMKOP1GRGnp7sFfp6RdoK
+1b46K8hT10i8RR63YQcO19Y5ZkDUyIw8z0u8/FgZA1N/iJ/+2i+2vw8+chODsT2
6N1Nh743oUeZbDhXBfH3estpPRnT6/zlJHzenyTCZGZXD4OobdUmldZm2M+CPmBE
YQc6x7FswTgwn0MyfUjsw9+6ronvTFcMq6dt79KJD5sdrMrUDSCO8uCjeL3Beb8Q
Zb55ldfj6V5vC8KR3wZEsPO9OvwdvwGWH2YLSjohFJYjeKNF/DIHDb3VUthv9YQz
snbwsTFBHHB06IzVOagS1GlN6mt1ztcyC+3Xl3S3MyubCY5s/XrmG6FWFwIp8SW0
HJB4S1lJYFZVapDFcttMvC3PxwTtV+eirlSMMT5HXRiv1F8CjqiGdFJXRZiGJ/Bd
STaW9gTDZLwPrl4s26posYOKFCIlnGFgwLYPY67LvSIylKkaRq6BhHAlwfc7GyC8
kBzG12lDLXy2Agkh8HG9xotAnyslFU8uAtfoL1at3nIQckGohaIuQfWgj61m6ptP
82s9d0i1i26SWlCmSmEyg4Qjw/6vuSNRMfEV4QSPzOO8Z0PDP3h6rk9b7JYvgXSs
sgozLJ0yueZxjPwVSqZG3afOYctxXkI5DiqJsXg70UxonxuyO6Ug4jtzfijZYeQj
PSOr8U9hJ9pPye4V7DylmkOKXZbF7R0iqLKxFb1422CEw/XgoeW5goXJfnMpNfQr
NflwubLfSE3V/yVnyllOr3nd/JczRiEsRLeFQVwDzo7qtTWuX5UQxjoiVbY1Rj8n
H3UdBC4WtT/u0ifcuF1Dh16oxK9u0dqlEnB3J7FWYSS2rqe1SHmuAvjtFYq3c79E
aHV6+myzl6WGPANLzqNQxNXRXGZolQ8aV6ksVdqfE7PgbLhA0VMJOsPBrbSI1ESa
amzsNXRivvEx7jr4egZ3EYaV8tm+kwDDDQk70fGwWwMq/u2uac6WELcHVJtadYRc
JLYXM7+g/drYwbvsVSKS2KYvwrKEkPJ8QoBO0SueM+MRr7Cl/42LToClYfZC8g7y
0BCwM1ua8/DTo83QQEGFw6CHlu/h/H24fZ7hwQaDEK88W+Cjw3KuRPU4hNHHkXED
niek96TUX15DqWOVdd0N59EM+ajf/rqcTKHO7/+auPbWHlL5RDZcQwv//os5yaLF
UcQblll6xranD13yYY+peRJB9RSpUokuhZkLV4E5jP8lzAqG2vMcxwyLMtyllXYa
YHSdd6GC8GjwOgYHjJF5Z9Vd4o7DUdjiaGXf6tEwdsTt4fNqeWs5TyUehMHKEn17
YPO7w11WrJ9jUYyCItMthP17YucB0wvpYd+dHexgPFXiA3xbb582yRWvlrfu/d1G
93ZwjiyTrMSSyl2r6J6mqJo1Iyo/Mei3Pb7o/TxO89QH65xPgcy49RzZKUmeojt8
eYpxGqsrhOaeuA8jqBJBBXP6afvl3LL1f2bQxzWYzhjnRZcGQmplbZmkCfBC4RP4
Y9CYhqEtAAxhqw9tpePNU4zS72sYkUk8kua2Uf9R3CvLQ0s3NZFJfJNWEVKX9Az3
KXhaTa+T+N24ds2Ee6lq+xkuK3RgXxEHN8CQniqo6m3yep0lCPHawAfjxp+n2INP
Lo7ZZE7dIbn1O21SZmIWuK0sBG03EX+6Oy7fklalm1ILAkzB+IB6H6+T9JtqsZ7Y
oVAirwJtgiNcQcQxDCiotC/wH6MSrKmC1saniukWn3Yee5Zvn5sMi2Q3J8VfQ8e/
WAqD/lEAGK3tfcFKDhkUXxmZ2qSQxaICjvqK2XaOFRhbje6uXa9Cdlgl/DSkAH0q
qB7kIxYjUBsfLRbnTNodfoJfAIbKUe3WFD8X3kSCv6kQht935mgbTPmKNwS4VSsN
1GDaoottCNl/I1uMiKle4zCwjFdF0mv6LtYGkOv+FyV++c/7HhIbZym3ZngP9vs0
PH7cHFWRRuO66So6dRzUOH5o8HpPjFkjZvzheLkUi1a0boyKXPc0IAtuCJsqoOHv
icrcooentEp/jc29V0r8OIgOUAOP9Qo5YfZN86yXzmf1j6ABilFXlolK0acYv/38
Dm2j4Swh4jLH3OVZP8olqOTapROb8PsedVumWxKBTlhhZhBn4cMjom0XZH6vhHlZ
/e1FBXMGTSZpUI8rsIkoqudhmnxXt6LKEtAvADMYcWuQlvGGnNkWSA65rPbSUlkX
TOPKgyza2mLuQ1IBcNA+ORx7i05iOHUn+/xxnOPHSVK2hQ0rzseoz1TbIepAJvgO
52VrrVU63gDm7GHyOq84qo1X7oa94wpGbu1m+bWDzKzatemzOGK9PKTFTUzZmTbf
9YBZoOkVyTfQpS9bTzZLAUiAUuc0VVGL6DE9bly5oyuEQWPkCNej4uAJO6mic8F5
DyqWs4/Y55zXpgJIFvUqj2pXyRBpR/5w8WX+kTQq+lSUkbdI5WS3Dsui2gYW8VlZ
/mkrFrJwVH32wvnxbZtUSRRqXa0r08dLCQFAIQN6WLHitkTGxxriEmJM4oIcnpuc
8LcPvQNMGy+bs2U10lzCkBGJQocKPqXtduJ2iBgBuoj9kTLf1iO9ho/bK8kObtfA
D50Rgekk9/LCLs0kXF/VN/NZrmdJ5MGMNOB2uyvjgVomtaOMbdvp253491qAMydu
+R0n0GaFoEx/XPQXPk+n+++fbOdRAeqZ8hkke6yRsvkhoIoMb8TLPmTeraThbTvu
zMWkAHpnH+WuY8n3BZsp9Wps8Z527ZrfogwmRIeUgkummU5L7OkmnzpyA0/80f+y
KU4vaRuoJ/8myWGQ3VsZMo3cp6j6DYf4NsSRbjjx0dtw7QatvRhPDWlHpkBRUDUo
m3itepyjtG2nG57Lk69fyCYELuZDVjy9Qoim8SHAQ8GPPITiILHivFEMGEbqQzxl
GhUqo7R4PmN070VtTthjWWW5AyI7JNzIgXF+ll9AhKzYbdXj/x4uur/jAKXLoc3O
2bOK/mqttAM3//ku4VhiV+4xecs6z4jDan81SBnoWDJDL3vjmamHESV4vzSVfsDB
KXVU9YOQy2J3UVKhP+uJHb3bfsrbPvwfoLwKF4zGIU2yS2tkl2z3Clb5prU7HZ11
Xom4CV50VOc4pMalLJOsci3/fJAWpKnm/FUToo3rnYJP1QRm+S+xZMQvb/ptVVll
y+iKk8g5QNxh6+vxSz9e7hEsUUvoN9GQyt7OsISwx20dOhwfUmhJiXkH/dt2fKCn
5mw16/QBsPuf7JVjVafMT7Lgc+zQj/hZhD/FXP9SOReiFS+FHy79jP4rUjkvTOen
HYuuMpkb/ODtcz82AXfzSYkTeKITFvVP6UCGT2/y0uMkYrtn7T4vIdtR9sT9BGgw
jT+BZqWqCVPtOC1kx1YBHvBWs8XrSawqV1CaJIbbcXUXiT9k4ENInuawrjd1jk8x
7l0XdrpIjymmRrKry56xpXMXC4hcRGuxCC3bGkLxLTWtLcI4DYvXnenWRBRDcw4V
QFFCHLl3dk4+0vemp9JaVndHcDsxDj7XC74xYkFCi4PLb2jtDekMvVGhhYn5bCoO
+FtKE1jxlqLDsGqHcRXAWEqZ2yBwA94QDnypvoSzEsyQg14X1S7vb3qNXIdurG1O
38H7uq9wW9uPQF75htkAMdNK1r137wlj2TQzWtTbr1ISUDaoAYTM60Al98anXvn2
6Q2oWYX5tZkEXqIpsVtxbeHY0InNkJ4oDtPfI/9PQ/UNs+WDEePQBs4RTRHHdqF4
qNUh8GdwdhVIO41BzkP1rBhzLfZYJkQkSjzHHSc16QazymuNRivzyPXkQHr7HfoL
cKFP8vnw8LsQSbp1d7fUdegT9fv4ITxuOE9SzVKtHIfhDbT+HhwDvuEnY1D2NMT3
aXLm4O0lPSkrzuIskxco+PwYdi9uFBnyrXgIyerf0pTykddV+15ldZN6L5fwPT4T
e/xYC80CHlvWKJrSvaN0eHTVcIOh4mMISQI50PJR2aPEch3XnfD72yRsJ1ZDsVkn
xE/FR5McAY8kgkqqu/nBp7RcLZ/3XcU1EPsJkKP38+ynZ6HcoTEUhT/U0MOQAAQp
VTyujYriUjX2o6r+kptnXt0bLiZ3kZcfOg0ZQHcKNqtifFgyJsahquL0v0YhS3uW
ndtqCANS5uRsd8dLytlbHb/CPbzhpuxGyvV1PLwUo4JZgXD8QEPlMboVkttvZQUd
pi8NS8fTrMP/F90xpY8FPJ9XBtZyWqubu07lueDhPMJZWGhbpGhbLDfMuslNe930
IhEfhS2xlPvY4XLeorDuWMW4azNE2sMb7oVIK7ZgEg2CCac+m+VUWEicSKhUcPJs
MBHGVVTO9myqSGzVsLNAyWEAuEEiq0AIUk81cijaDyyAvd18gAnkyzpUjESN+PYs
AEQQBdyjRN11+RSAnYCpr4U+ZQjX+cqAC4BdHQQlMX6CQE7XjyUO2sQwZOs8WNPU
YyIl0pkcw7gJ95dRVE0qy9CnoA2n8OnYxMAr/uWwAnt5iuUKwKZqRoQ88FTcX73t
81ebzCAq6A+Q1NdnDULr1yai2UDNb0N0XLiu6Y3RXjT7fw3bku26cZPSjVDJf/ZC
Qxbwxw/mc9Z/8/N24xz8oiRKKWq7SrMhKAJtEashmJsv1GKdiZ6zbb7ER2hX3R77
i9JjOAqchTc+k2PGjnvtEI+NzdnRzQqUad8/gmwlWsRoBHPlg5weNyszVlZDqoZC
J1wDQ6MHKKwWDnfdqooAj1Ko2b0RVH18d7LEvO0E/OWSLDqR5IgmBFsHHXo+v9/w
SrXIYPXNyw+1JoogskZzJFWS2VDLvs/pBsR4+Oq2d1go7608f5l6DmqRvTMVusjk
LlkKxN2xZytNFLPnheK+NbmkvENKYG1gHDEuAQudT8gCsAJg0PPH+tA6GfcBJbV/
MYxn1JU+BNfSi2bAZ9N4JBwqm4oHuMMIrY507qSTiPgWYj+UVIbc/gjU59sTLHl/
hAO7AsR8JFT4jRiOKTib9smVJLPYB0/G6usLpGmApZjieTjzfAmwsbraHYbpoz1K
shW9sNvNaXfD7BRrSFyr90BnMoCoQ6vmf5EHC6NntxsBbQEwvTnUnK5/ELGJRpIv
cBc5VuOjyuk8DuwZHmy35I3FwVulXQ3ghRI12LmM/NIVLdMSJ8ohkeeNW0qF60as
NU2PAg6I2+faIjziaWasUnLeDJJAcpbGrJGatNOS+ANXRWuICy/vkFn2hTA3t9GU
73gM4ZC9ftGf79UygjIz8IwYcDGYB55SHOxPOtA8Zwlp7zajUTse/yV+faUevRWK
j/pM8FvXJhLKbmTXLXSA5DdCeUQYZfx+LuGkv4b3M/bQ/o3AYDwhZYMaG3uIPZuP
f0v3xp5ZISS1FXmOF0JEd8AkcbaT8F3e5ueVmatd8SdGB+Qji3my2u5PSwWM510c
cgCN8WH3/fM+PKilnE32O1PfpXNDxOnlxgWXCgBGPKtx/88492SVWnsVr8qoh8hK
dd9OioAYDzg9PLd4p/o/mqYYG2RcwSXf6aQemjFvxYbxlNKttdq/xglT6hut534z
MESq/fQ5mMETmF2vWUV18gBLTjhYc2OC1k37zN8dBy/2NmbmjXGQh7scNuHrik1f
rOsUYm2bSb10hIu5uUE/fHl+VNevN/8sNHm+vma7bBbZo/PSQhPxgiylKosyaZC6
yJhSfNaB85uGfo6F0r6NwaVceK5CTZq5bWkuWLRyjcWTnoo0S+J51DAhZvXxQVw/
HvMdtV5CsCXLucxEjbTROwddP5AvKGlOM4jSEEITM0CSKwviRFvHwBFwQRUpOeN8
U09b2VphKd0bxN68ipXM0DDYo7Nz7CHvZ6ozwRn7sHwoR0GaVNjcnooRsQvHAyuX
7dRwn2fclAolwpu0jcyJyntkyNlmb6eXt+HaxYHWCG6keXyj7uBPpqHvrNDK+2ws
x4fjU+mIBYq75r9e3GOfKQRUrxunzfOtfwhy5YOxIRaD3PEVwGeB986fHIIWS/TN
jiYjI34RytIBZihFTvzstItVSLZsxiR3rr5F/64QRBt+D/+UX44ZuReSTBUPv58b
sQj/pnypGgv7LEjyMuDRnHAFjSp60DhqKnxQjrryiDspmdb20eWLy/29JLFNhV1f
Hpp2POjdcgcCRSawGiDJLqtSOkc2yzIfwKrIIkMb1AA5N+y1i5fDBwqSRMsx8WaR
YGUIQlIlEe7bxlnepGfREks+ptB6OV5pmZggMhubiaq8uob/BxVz9RUAqhxB4+jN
9S5EY+yrpYd9761QcOn37KYt73syOa1/ugo69mf7h/4vviskUYw6PxX79QQwGyiU
0xJCAtjgNY8pDRj3Yg4IP4qHx3EENjsyHeuH+A8eRP+QpwyF/gVI6//NAxck/viR
8odH+BSjC356YEXBm9jx8rUR8wbSU9LjatmS4YuhSS5Jymscfj105/WPtfmkK8T6
Jrjc8zifZpdWPl+lTEdjDcspqmVez4Eo/NdQWxVg6nMZ6rKHrqFPJ0C+UxOpjLkW
Z3iT4pJFd1AM7MdV8Xw4uDKTOFxUKAVaEB0Dy4MLqWtTjmYf8KGIbgY0YTGa9DXI
CmlM8C0ecUy6twCrGnO0y+0EN3R32t5DZa/WpaJOeEVoAxOtP9w3vu5yl+RmzWOC
HezQ0F6X55/zgh9Mw+i/0dqTy7IhvmWNUMYa6MS47ZPZw+eOX036fSkMDMLJAFIq
Xy5ntQyl1FpZ+EDQbVOTfI7iQoAHIOMJlQBKqbZ0bUx4CRvPIlwz2ZtImAMn8gfy
L9Gek65jsa45zoVFtaKIxLtQhW7SsjAhF8cY+ef55G4HWByUNnKXIpfOSNSaxaDy
kN1gdAFWsveDGjWrv1JRhULafdCogJMMPiH6/wycbIJMNtZEyOPSZDKqEMu2C+SU
FkFq1PJEyGEzh1S9v/FRw61SpXByvNj6LTDKgBZOA9k9k8d7WLClPaE3idvuf/6O
FhQyHDygcMByWYtDm2fV240W29C/4omFWUE6kRLjFixZDN+WFmQZ5Uo18WeB9pMi
7axW4Ei5NCrcMNXy9SqGMZpzIqhjPQctdUfcHXuZPmql8/mZivjY6M1yMAga3zr6
7O0c8Jig7HMwxGe1NJyLDdKmlLga0jxT12Xuu7rrCoeyNAkd9+cK9lRgVJttHM3B
E6zdgXhmaW7EQXiykEf84VGgayJ+X5I9Pc45pptevjJ6Zmrzk4eaD9liyg8aAc/r
2aAGfQ5PbWXa0TpiDNnUxzzoAA00Mt0gb2pwn+ZMbNI4lcjVjuoDiPceVa83cTiO
nMrhOsRpZW9kkkkhj8j+zCgKsWN3QpT9WufbI/+dZHW1spWCP44X3w8dyrXtscyt
78ehDx4ynyen5cAmEOFSIIegfRmfrxEmy48WfY4wdRvOkHBr/o9NKXHNzfaFqI/3
hAYri3ZWrVzNsGEpUjn6jHeuu5DK84dPUjD9tn93audMCXZgEyDg/Vt6SMIBRBy6
Z3fRuRn26hZSHlO/FfCFCyFPs9P6h9qJBm7kT2wN9phrYT/0iim+CbbYmWhHKAbp
vdMKoPvnjZzvVHyNDgjs5EhC+zVQWw1+W3LaapXfw1m+WZ2i4gu/7ayGk79agk8P
vOKexc3WESrpQr964hQTaahILToW2T9soazkDhRf/ySoB9dO082tSmHAIp+TZWOW
NawXGQg0LoZqWJKDVoR83MsFeCXXQAt2Nil+mJpdAjfMQ9PYYUJw0DRlnYxEd2Aq
90USU5qM67bco+9xPsiYOPIxb5Wte6iqe3WUhNpmJI/lz3gUa6hyJnITFquI+QIX
qKzJw7rGfKUBcSKr2XDYmkG400W6t9zHWGoUX19y27ny6beOHPiQPuSaS6R4XXWw
Gv8R8SuV4TW0jKPfYN1R/ibXrFwx2KvtNv2xMqksswPf/9bgEZLJ8WJUDmGOTezD
EykqAqoDaj669mILquUJ5V9NcVydAw9l7x5bb/PPYAZVLqXK0JxSCS6tL9MCKG/L
2qP5F1mwwuens4sv6n/Q2AxRolF/yt083KxFE09BpuwFF9OoySkMugxyHzKiS48U
SjVRQerDf5PrbHcYWszWNsj4tTUfoAI+mi03IceN6U7CxM0JWvaiVx8KCWDZP2dG
Q0Sas7Ow6FpSz7nPnsjwiFgqC8KxZ1KukARu8HLGvUadV/NjdvrVAQ+OTlNnzIFi
wM1dN5sVjoexC8mm4p33gyTptd6TYa3GITfJ48hW0DKAiUDmqHgerDfljXpqmCg7
iyPnia+lVvcCm6JKrT83XNScY8jDC2C8cucEwWANkXBi32PDTT2DzsEzMpJMQv4s
j7yaQdQ1sfVsrT+ne1UAfi4uh+JebWOWGoqGLbTUw54XP3Z+gFidB6U6sk41IwLv
mceNyFFf0M4iwqm4sHdTFe2ll2yiLqFVWio5w1tcQiK++19Mo+RV+SAnzMJo2NaL
+3rpwO4KHoIT4TftKp4pHngjBYw7f1AcfXI7Pe8nFOAxDJYzD+Kf8h3xdHrGBB2N
zWy3jHv/HpRCPqsgsufrE7zK/jBykn9s0azPoJe2769riisDjh8bjgTDstctGeVF
NaPfhvEMcmTcFaJbchdr6e2LWVsl9j7Lrc+lPr1mjQi5etc36VB4ulcMVS3OH25t
pV1IOwUzy69/k2WMh5f/N8akeXN0H99cmmXnPsiGvLlhGOEUBsCUE0Kzwqn52fT6
pLgcqYx9eHMV8PobcvYPElOqUpk8d6nm9khzLfAjiQ+av6b26o+yGZ81kUpCmF8V
mLsclXo612iLyuHC4HpgOmNnSzOA82vjKVouVEqX3ihWOodjppWFiZJMtuZyWDG8
ZQO9EbS2q0jYtpZ5l/71kAa5vnasXLUo/wsLF/L/b+TR9nvx9vgBZyvFifVT3g7D
BCpdk7g+cFzEYs6dnK1Oz6bo5ePd00A8CyQDRexA16GDCgGXD2bzP9Bt6ZX7my56
pcDbA4jzNbSzNFrMN2iP+k/vPwWWncf3MRwfx3gUIMWpduH0zFFxyEFbEdkrjAMi
PGAJKj7tJ7/3pBQUvvlJygb58tWOCTsLPrYxjeu3lCAU7cDWyzSgqRQhCUgwMDmg
mz2VOhNkLbbnlnCyBKz1g5dLekOvNeyNmpku8evsEk+DqvDRp1zgI/Yh/xjFJQCM
xBTB8UzEmmniBOGgDAd5OwRIW94qv+rTQGgWGPqHa/AR2zZeBGlqKSbhj68LLpSx
HFYP6pjgn8r0Ibmt0NUFuIIAqvxmjldTsg+vlUEKbRPcr05WDrYxUPlunXt60hLC
pJgmI3z5JwCzp47ktZptz9xbQziT2Hc9qd+WZUl0ORCbEHEoAXDXU8zdWXFwr+h5
oAHyrX/kgi7qQBUtqkw54CyuxRrsRO3fflYt53ywXQ/rnYf5/j+o6RmtIYBnq8c7
6OaireZJT4LE81d/VScC5cTSq9/+P0RQ+Era+VJr+gVOvKLUNtonafQY6onxkFbs
Rgz7UsJS5dszCPuhMGtp+lyUAVjVmz5tEuIZtgZ0H53qRW3CiBe2WG61yqnZqEN2
FW6Y3YrnatEiQ65Tx4f6DgTGKsNu7htRZMxhyW6k1zkROnvXKNAag09+xBQyJPTU
SQpGmKgi60REBIPx//9AJQeb7LyFl9pltfDXMbGo5qxm6aulNn+nTSFcp/8gik+3
oZtVD/RJm0WBVosxjbSw7lN7XVuIiUxM6c7/xvO/Jr33ZyxWBlT5JQqNX+bx3l9e
TOyBTgi+4jEhRE0dDyrWiPsE4FNPLyEA9VoYNECV/eQnnTitTORuwEG8jYku6UWS
UFn4BtAltGuZqXpAoF+1M2OdpIdic9q4nWYQSF9g/EwYNQPXktlkk5/8krIzYy2H
xy3wWt6RpbLbkOzKza0IezSfFwISHJhLVF90x5RfNU6tTnHU0APYNGGj7QqSA0nh
vZvaionDaa+Iga2LyoRQPDxT5RJeOhmf1JLJGTnJ4lDQWLqB371eFdkHmihRAPKQ
xDbN3GmTavwKh8Qty+oSW344+EewtXJeeH4W3yendWYNJJyLEwn1wesYI67bpmZy
lGeUQAe13bTFU5F4ZiYb0mZuAQQbmcWQvWgeBIAsmTCR4O1nT8bRmNCD7hAGr6u/
1WjR9fGyaiPH8p0t1U8veAHuEHcjvJKj8Ghzy+yN+frk5k7HFnky5zGS8ioBXAnk
OVKqILmUfP1syid22d+rpj+RwDR2mx8zkjal4gw9pnid8mDM0zxoWPvHVCcE+6Z8
5Cdyd9m46WxnVYC85Oq7FUNRPHMzerhSBArwr0nQm5JLRZhBZZb3Ts+ambMXyOY9
b/gdDVAuOoH0yWRXzWNojqKxS9dFtlbrxWR3uUJsK7G8ScjKzT0BHoBeC6keodGb
L1aGGh1QjZf6jdH2R2/16zl3otbtMm8SzjK6mA/29zuJ67LjvTpj54eK/YeD7YsX
NEr+AzM7rZMuwMxuVZToIQgQeAmX7u2dsg3HAkgf/hrpO7TZ3EoAfn7BZx3MMYtm
NM3zcFNLsKw+var8gHEnPTzX1E735PgMDcSTMYmJSFd5YcXSBkw7RHgTndtao7Wh
IR2ykDUMjKWyzahT82pZr8iNUhJIDtKH84OHaespDPFnZyLDUrYxLaPa/HMFIjCm
LfSVu4sQzM7svIvhbJMRRyxGX18fQXuOlhpMcEKG7APPjTTi4FDff7Mk8t2b0vft
lH6LtpGd3vmBa+R2ut0EQ0y9pzDohW7B0X7gGXDYh+HuH5nUZD1Iltdt9+uNURcN
q3IXC9yoVsnoxUh7rpif7M1YKNGxQRGQHnZiepg11w5UngFBnHSf+RrVzre/l11R
YgoCTdDzz+CdqWfjIgpivKqP2Aw8STfOZ1rF16rN5ekQqnzg2IHmAVR8m+ifOIRf
RnLM2g46Fa3LSg36Tnlqk3a0BPAZLG9E8yf+IFslc646z2gnK04MeuerhwnIfaMj
xLnq06bbC8io+Bw1JExBuPFo0EySdgEXU/O3SdjqYbWrn4Fj4RVlxRGGnerPcSP5
3mIpQpL2TUViz4AY4Y2/3/9QTdPcMNJ0/bUadfAwztOHu22h4+XKACarOtnyGObQ
tHPF7UNlG0GepyhrmF40Fv5VtYQooJUTBofIdtKHRBEn66Y+XDlui0nH571ZPTJ2
SBCPWpB76Q1hEU4CRqry3djMds4wfCRR8AnlxmSgzWEdzol2MlG+lTbqyxisAzUR
XV3VWhTa0JrBV9+6STQTO1ncvQFiRi4WtMZqZcpIbwz4JDHmE8AH8g5IT7prtOSp
KzPmMvxSo/oQjevpWq54ivINQHP7MhqcTMqWwUUyeAM8HRq0bh/XgmjFxh902sXC
cIdILLwYoJ0GiXiIjXciWD2cZvAXgQE2575oKvu643ym+4pNRFebyMq31BysN2NE
A/D8WthD99kTGbcwA9QYO4mrH131QFWZRt3TvHmifaYt5L0CdIBErVewKBdYVY5e
i/9VgpBXdlWJTtKXegxSLpg7kQSLerWgvNM9mOHXPYP9ORr/qM9bn8PKNRLjxuro
Md+sZxpGL5iufB16nPIRutWHHmDQjbUtZcBLov6GlYIJ1JEOVCA7vKydsGREAlCY
fGzDvbb5QecqvcBEb5ubJgLKLG1NOkTCk55qyEN+rFroh88ikgk6MU95qvAc5TNY
t8kOLgkJGMZzpb02jV00v/Nat+QFHRMdbE2FbDylhlRYI9OtQBq3AvYZShwvxiKb
A+6hFsCKk30At+QHZbj/X8AsiOFMPZ6RWIAxzf91QeEFWA/ovsZsEfX3dyQbIKpy
kEHegqw4bsueGcB7Mu4ZlLGEnKBiXOU9jOVstGdfnoZFpifelrDG5VDCTf4aW1Uu
u4ZaUpkU4NXS3T1P25RkGzCPSDm3jsh1JI8gUEASaTZKUcjfO+4fZPg9aIoqjPjF
xTYxBDDu7DBAgNJv7e2uLagupP0FhYUH4RuCrrA8Hm6Rft3pNyuPWYGWcDYzZcBP
/fuiUI/Yy/1oTQGgjHm2x+97I7LhqsD1pjMWM48w2+oac8ksynow/leilt/8lCcA
I/p/StKnQKcZG4fKkGOY3O6dAUS5XN+zVE+LmqKV7zey7uMMzLBGhbIZUF82bFWa
M17Do694I16/7ct8HvonrG+y90czyQKudr+7e+qN5/YiT6K1k5Ggaz1a57avanN2
KAQl+iYfpnkdE7QAzIen0fI4OHwWa2c6u3fvJxXROgqV+iGDpbpaUaqBgTh7hGxG
qCAqx8b1L015NfGL21lQCc0PTzKC5k7aYJIB/XkAS+rOojb+lBYTqvG8BXx5+NZA
bE1TXpsh7Dytle4YhxKR1kYvpAS7rkYhZnMLbrkK3GSTLRw8VHaLX8SDvDLQpIyY
JDH9cWIHyUWyLmf68qwRYy/3H8Opo+ylzLR/Q2goTODMQSgtf9MsVbkt0iSyVTce
48BHWEDI35wKOnYIkzk2oRaMEYcNALzfkoVrtr/emxyuzOSr89qejDPJ5pFFVYr3
KLUyIpxeRXKnyqMTbZxwGkKQ3SA/PwrFb7bOTy5NRZgDO3aIE6bzYpmEM4z++4B/
/XLcEjK3eFREbsVl9bgH4FrycqTSyTevzBoOTYC59ObMvCwVZm5nESzyqb0iq0gV
uGIrPptxt78SY+RYk7DPOpcpv4JeHjNQFFB9MNDftby6ao8BmIogk4RgcU1k/bKj
qZNVRGweCOe6kO9qg4wG7jqmMicpKH1db1DzCyHBGDUn+mIV93l+KSXcrPhQ4cYX
k8/vRWn29dxgzF7bDZk1hWUP/RowFvbq+zs5oHc85AkyH7eiSBnKlfIsdmPOcGKj
emKog0I0x1aANBDR2JZDqVCzkfZDO/a+Ub8LlK8X/VeOda55ZSv3pHWHW42myYQM
2svMtbozcZ2dHpQ+8C8vhbdxWWU8PI856SgNcGWObSyKxZcCSUaW0UQvwhjDHJff
vzXvp4xh9zRi4NG0/1JpNwxgyKliDUuZmK7AyxSiVlngmGZkW9s2BkuXyoqI85z4
+o+FcIX20bZJ5KHuXm2CCl8P2yhOhZpEUOnKARmtFOPALFFHvyoUqHtYbXvordZF
sXAblHUrO/qfQsXEgt9LO3skT6qPi/kibAAqCrpEwPF4PAh//4uVGYu8Ecy6PCV1
aWOGuRA1FsVyOTTVcQhZx2vao/9iUWRJnNuf3EiZ/LMNbb4DC0sIAeMPXTbLxGU9
qeLaAiHH7uGkxJVxXSTBMalC9M+2TlqoXccu6/uOpq04B1s6i1zWxST0HxOBL1Eh
rIfoLghV2BA4DPR8DG193q+tTEx78SqkQ6d7iPm6VfZTk8uqH/FqMpDqugtQVqfV
vDmsiH4a7FWrg8ZzSEIW8Z2nmtQhIdQbR3vo9OXtFGEuUjLPE6j9zCSg5YiSj7Ig
XOZvsUs4SB6LRwlo9p7p3O43nmMpxRvoKJ11g8BTJGiKjxfFA9O5nQ+uXNXqt/Gd
5HMa15RghypDIgrHQIDC6ZZHNO29kFY/aXyH/iOkZiNACwg/j+LFayp/WseNfimy
khm5lwhQ7HOIU4Hhm9MhChR/0sd8x3mGsJyzafYobsbEdydBMeP64c+UswwswEPm
/U9YmHVFDhBdwYl1MTSviDE+h5YgUE9Q0Atq5UOfFRlQX3M1CFMtZvIvJFO0tQBi
0M6niS/7Jbxv0Vf9dMyF3Ewqly1VRtg/XjNaLarVJvVAqz8YYkcsyxjFeTd9/byI
AxRV56W/fZzsAgIfQhh/n9QwXMAouEjAn3iD3zNc0pg/UnnT2fYHgz38xrxKobMS
wA45ZPlK0wrpLCVI5H8Swty5EyFlgTcr16pLpLjRRDcX/yaTag8in9acGalTQFor
aAirr5rSfgBryl+bIT3/XmRg2ImGDGOFFczbQcfFLykSntEyP1a1bIaREZreJdNX
5uOSO926cqfU1eD5S5uHhSGILy7rz1db9kC9qO1305PNE8YvXy/YWF6bPjnsdpnM
bR3f7Y/TcwdLoJBY+LzKWXrxlhLHUAgU/hU3b9oX4q5whluvPQw+evfKUbnZcwgd
0qY47IakI9tlambw8zJjS/8omse3i3DLglKhx0N1Qrqb4ZvPLVu3k+9KhDjEi0Zs
NnxlvRgPh/dQuo8LURhZOGjq3vuh16oROa9VKL/ZDsJsPxR9TARbeM2PLP0wNFaY
+s7HV8RI8+T9oyZI/k4uwuqTh51x55t5bQf1afSbO3synGoRu8cJCmZr3pbFeduo
KdISV3yGqB9v92f6zRkYOQujBm6KiDbIByjCMB+ghvbvlXl19iWFOmyhfqG7CWr7
vGMCsF2V0pF09x0xsJuLLeiW4p9CaOL4jtmw7E47eMzdYajGGk+x7CoAFKyf0KpZ
0yztYAyxoE0JUhmaEicXFh81AFWZDAZ7OJsqYqdBuRyqyIeiv5bBXJgVxtLTilR8
AIt/7NSkYxh8PPPq0F5mHjieXrzeoGJBUSxNbmoGW9IYfKB+ejh8OHtYkiTsf+/l
ds+UkDOkakh8uoEwcsO2H0gnpifbifTVGjju1WkG8ExXoJflGK2FrTOPtTsVg5Oz
LR9GdUe+f793Zf7KXZJBbLt+8x0+4P5T1sNWqB0594zFrObmxT0MeIkYajoXXQ0w
BB9Tv0XSJFzwOzgoWFcoDcN8fnsH67ssgRkmCLUq3FEnwWUs0LwvUf2t69fm04lD
1XIxbfHz/+LTbNn3nax4/d3JKtC8aMo0AtAGZ3Lm+rvKRDKM/fgoQ62d6JwYD3oM
NFPm2sKjdnaNASkpsyUTAbK/AJG/u8m1PSuX3LqTrwY4aBbvfNZaPCwpFuVc6tjj
BEu99Ouva9d7dfaSLMJg01VSXmShe7clV/WI/UkFpFU7Dt9sLa3HS7w2ekAM1Z85
Mog+EX4XmUM6NUWMAeKLWIHH8ocIKmWzUig6WtmX924cluanEKHdgGRTjqp0UaDI
dcoHxI/Cz90oFpzqTnORoWtJxNJc3bLOP0imd3ZpwHgqYeK/eoelGMYnVukGSY5O
rPwMRlyjzmE3BgHs5ozBoEJKwMs6z4L9b5aP4PYNlLGweenD1oqI0teEzQalJzDO
Dlc1z8E+VKPx2VI6MBjnrDP6Yy4GHz+uPwYd1YVJbgYNkONEfdvK0YJw+odbUCvL
PIWwhmP1Ulz8b8VdDQiYcVNdzG19jdsjAd8FH5diZ8Gwhw5KLOUziB6f26NQvkAW
v2ekBUV6FsI05BHO/WLNZ/xi5mVi1ytCQzpdO/Xr668Zw/JwsQ/NZxezQ7jsP7Qh
fjGJ5vzk7a+1jN+f2lADrieFJsuTAFc7WUdbxx3z/Uh1v7dXs3+0Ij5O0HeoA7P8
4aGjKDqpkgEec/8IBttRXiHhy2+2yr25LnjKQC06yX0TEuSmN+KforkNifV1Axkl
saPFHvQW9h8O+5SAUMpwYXHny+2z8qx5cmXhAnB9UFoXpI8X0VbUYPEaEzPiArxh
lKboD1rkVrib4xgz4ZHcKSZg3YllB834Qg19cEVwTl2US1mmcg2wFiesqVnAxP7W
kTXdUBKmQS3byiBZPM9DlDd2N296nyueSKPTxEaMZtONmUDZmc96yqT4uN+3keOS
m64mqEQZyQYFeoo4XNn+U8KgfIADxh3IxhQ1r8/6uHEbCCYPNrDnyKHf3YxwlIyG
Ii6y+LrejnTY0fYaa53V02rHImJVgIhhbSTqWNY1HII89HIZXK4umrNdYCf0SlJf
02V3aaaJDiBXA7VOoShOHoJtLAmaqLknka0pcu7smpzzNJ1sytmmsBJ5xGhiP513
yGfjc6aaTxK7DpesjTs6RKZWQHW5b/KaxA+8abCzcylE0Ha0gWoxVcqILVku9/yi
J0qQKVCd4abtLGVXuz0nq6DQg0ntzH+VsGn8Cl4h3B70U/7iGIRStewP0IUVFrMq
txqCiweBix5n2vWvZPAIaZOGYU4tYYJSbGD5YYx/P7nikbRYshmgb4nnBH6Qia3O
qvfQt9Onit7UDWRimzb17ijuFr5/eSeDhgNRu4VYIAH71kCZcldrXfzOrS4ptSIv
LVjL8OcA6ZJWuA7BjSp3gbgCjsPuX2zYD+0XUpLdrpthfnNbKSXIhwd4bDZ8ESoI
S21iOVs+q8N6gfEhOBuLsPJKB/ZayvnRzGUzX+YCppgQnSaisIUIsR9flWdzlwku
nlxV6eBjyopXSAlFBvFEGqu4bViugzr9SkgrQBBU3/eA6SI2/B142IuyF2Vf7udy
KpbU5HFhlWEP+Ny7Tok0nCv9atEunfzUV/Z1usRv1Fl0hbE1K/2q3aky/YMad88I
AUmy9xvN8VIQsir2PgiNUZON5+D2csr1jeTLPZCYWlShY1OZn6TOYl3f5hKse0Aq
smOPQKPKgkdxnboOhxXQYOcxJVPooRTfMSQneduAl6kOVL7OOGfGvJbz4eLZ7RqA
ZoqPpabWZY0sfSpHLy0EmUSBxIOs2vKvGtQFWJFRFJfgqP65E2nD4dDCiQjUgLSV
vHSlXnfumOJQsP0wGlrcPla3bSSiO7sG7tqqL674RkJlrnrr7DfFZ2Y2wtRLmzcO
K9GIpdGf0BXy55ioAF6zii4q/Sk41tgPU+itLsYJsrMsOpKkfCrIKT058xfXyFmF
lzb9MPjJqsF7fCIWtazrEPHl9cr6V8+3bOtsi1vCRYGivmFm6WQOCOdtbrErfNba
SCTiGVDSZ4DoPjKQBYsIuY0G0R+QB3JdtGfND2I2UJ53qJCHT7dxhtfoRsOOdcl5
NVzWd/jBojvitAZYnuyTclpGPxvN8jMs2c+RdEUEmrbxH4i7J7bNXsSVv+olfWUR
2Wgu3ESnokXT9+SBooZLK/An8zCiqAh/iFP5IO+dRVcJ3gyiB7zpLesSKf+WcZTx
+GfPvROB2iRXVG+c7TSITmQr0Z9bhLz+v4qoRrQJR+uB7PWAa/b+Ixb7sQjaStwU
ctfkqu9CKAyR3eJz3QoQPNi2ivI8lq0GbeQsQFp6qPxZ+lakpjl2KlqjqdRBXDl8
JRjaWlHnqVGdwQDyRAXII6Wir9jgP+3loFy6/Bt4WZjgMUnMPul5CFKoGUSBN4/a
t/XT30dUTemTJkDlygODF70V0Yu+VTxdBmpn2ijn73IC1DT6DNH+Kcf3SG3HGR2+
Lnui692lj/pjlag9Wnm7Eitnmcl/YE/nRcj78kBxTm/rfqG2qKpyKm5uvJRO01mk
kg1F/a0jP5ei7RfnDHEd7/0GJ5YvD+8lzG/5gF+BXBBaPG4a289TQM1AzTbw5jFk
4QycEWc0ht6F1j0dyXXlPgg0FrBKXiufLRxSTLZsW5fna8r/akLc5FPhb1P8+3/q
FPtthi6t/p6ex6Dd3JYbE832a4/PnToBsut7Z12Rj7kJWri4Msj+IdEGewE8Kj8a
o+eMnuNzumI4gfnjbykPVOsmJNUFo9NFgUv0v+ONxpmioVbuiTlTTvYzBZ+d6VWi
Opgs3PMjV0+ZaRmkG22KOYKNJAy0MXyzdqrGkyrKhOpu5zCjBN1ZjzQavUiX+fHr
PEmMH3qNmTvrOrlhVANa414ZFvp/rMLASamOy6flQnww5ncDOjWyTxUfAFVA7nhP
rb/utj/DfSFX7qt8soFY85HUi2G/YxBfcjk8ecYDsGETNaTPP7Meavw+YJD8KHxl
1zx3SiQZ44M9yAKiwtkzxtwN1BnR3pKRZ6JCsm7YqEqSfVltuk9yOD3A03E+T7/J
f/lXAYn3KDQSkQk6TRq0bOmVuBXljCZXvavDDOalf9asOuoKDWZ2uNJqnp+61I90
ILMflVP48piLDoFL30K0WiE7kRVCIXs5Z1qw4WOykGkG0wOJWMOeIJs4i2AiK9Cs
Cdms8ilwfoxLc7VLdH6ZtPvb/l71kJ4CIEOhoANE5Ny0/9RCANbF78IH6z8HhzDS
YbYZdACUsicv0NXag3uQE5ZogqDDHt47EsYFdMvXWgW0pBtCF8ODGPoMy9ypvv97
YOhdfKBQf/MeZZ08WYXGeSzQ9ZQXji9fZrpCj4Jy4anfC7l6J3JS+hTYDnMXbLBi
qIScuqYXs8xRrqeJuIy/R63XcEHcyAeWTEXXZEgVbnIDGLoWLAQjZp6Kvd49Uswb
pfMq4ODtNtWAjUw7fUBvoPU3CHZeJIw7GPF8LoL55/ljxS588f/fFkTr/HyEvJg4
4gVEZGJzNKlm9eteP2a5RTSzN5lrW0e+LxtQG2gLf7jAnU1+du4Gmz5wCT63NxoL
VmH9rpI0/pd0wkFOY1RnLrCZPCv1MHwLMWMUBHh13WgZP5LVyJJ6zUZdCL5hZQKz
KzmJFhM44Cm7ASbLftT2rNq3LWeeEJ/SKrDpJM8NYQj2qJ67zFqzkyuDHZugzpvj
VyH4KxPVLfbd/thficz6+pxUCMjpo3CgsTOCbSQVyjN0KQRU28rdQst/E5hB72kb
fp8oKfefclzD17f8rEFqrQNqWln0OsoddLUkbSxR/OG1N+hTx39US2NXfOV0iBBJ
SsDuXPzDLVskE5i6UMBAqdDdBTh/3TL3o0kDC8Dnj4Tv8KEX63AOpkjku2dOhkzr
ZZ9pZlUQ7HLTLtbHmgHm89+UrFdoCsgt0CrSXl9AkNSMv173vIJKdNmxnmD5mhdt
SGnwSunHwhh6R6IlwlYqwid0G94TFPwOb7QuAXCsgioXxJVJnVe79uDcMmT3qwPK
HvyOijhYHeuntLKOTAwmAD5OkU0oBCjiX6VLCMxiZ5v9vDZn4/qfCD2pKtz9IrhJ
5PM73EZwvKaqXOp9YqHWc2yGrIJvPyR8KgupxMipF/vSP+8/s0IBIs6WHuMGd3Av
Hf5lKfH+gl7zT6Sf08QcEIaNMJVlFzartjZSeuqV5GZrse/mVq8up2sGUqyrNpgW
ZipynH53XUucWrr1LouCQQTW4kZHVw5J9s+GKS0GrA0Rmk0zhVG2pe/Hho5bkaEz
siE9bHHwEeWmUW4HjiElr+hTPhGWKxKu0OtzWw0F5HC41Uu/11Cu4JuAwmmMmbiF
2mssic8A2HIIh9PgzVn/PCDaPeaC67JXsPhdSl6+W62B/rTSFo5QRS4G8QTvtUwX
mWezFO30iihCSR4sYT7+wKyD+yp3qeAFVarnfRndcN2U++du6qLMeTO9eKmkpHvs
SHmJx4vi3zVbAd9p0/GELpnGmpVuJbaGq3b1p8eoq4b2wPEp2qNDPS2eMbasNcYF
eM+pAoSmIRytqitv1JD2RATsXsG6YzAiVD+C1jbNn7+4693CEd4CZHwDLetlFpmj
xTZTAUtdeG9yegF4rZ5Lzp5uhgXOrBTrEc3hJlX6O7ipec49NzsJ2sQUyiIsn7uN
9OI0riD0WHHbFy48hiTSlHgF+hczxYz2P+iOLlFK1twIsEnj6sEOlvY0VoTfvPFb
VtCsiOQ4xy5wOb/TUja4u76H536b9WcsSkGAa3qJ6hswPFUKVnoBUDlNuoskRa2T
Y4S9pH1eFevUhQLtErItPRaKXyZqQoQaqFW3t5j3QrWdBVCAIGYJCJmK+GPR2/B6
gjcfDgpF6BLA56UPyGz6iCjpYwg54o9RK4ZFHTWbarJL/z7Scy8M8BXslQpZOVz3
SRk4zUn1jnqQpeSNZx5pTJlAf16TidTrw5e1Ass4JJcKySXU3ZZimwdtS0uSVd+E
oF3dLxkR5zJSGFTaD+FiosWpSQuGJHt0678/RonLRNMVFTyLLVxZO2jICW+SHz3C
KHba7XwJl7YeqNbMep/qYc0zgMpxosrXvixjgWU5TkwLuNQPouiZEsQsk8uVBvYx
BbCqhRzTe5BxDnrkFAhnuHsHXY4EVsVV8yz9Gn3XFPEEamXoPiVQtjs/gKxwp8AY
P8SlRGI/rmZioRcX9yCnBatmWcJHzqVXWos6WMA7goua/IK6j7bwuuFd4eIt0Pjr
ghLoOTgZBCrHG+bqr75zFGipuONuUlsjSb0f33apdmd9DKq1d6aBuyb936c4Lf0S
nWbzXhnszdbGZE2UHV/6IZU+MvuIkTtObak3xUbMlcUXSK6Qw+TT9LZ/yiJfLEYc
xSMdJke10FU8jozQWlViQIf0GVFKkBhDdY9wRXx35MokbV7pNoossWJr/55oe1IM
CV9BVnSuVQvYBPqFDFM5znxWy0t+HQw4AqO4r0Jwx1/T+ve3HQt9A1x3cvDsasJn
qF2iHXEN44aAHUZoSOmELrGPEFsHuw5d7KzcvNiLBQI//Pm6ek62QXe9miT8PKt6
5k6MfIlGNMDsNBzGKXenBl3jjCIiFR1SrpMaaVEAXKulZpCQlYjBjFnE9/yeKf61
HH7YGx4pT/I7ODD8imUL5Gc5y2uoWNVM9OUWdCvcT8VwFYULc7wnUDOaj5Jop/Yd
Q93JhMpzqyyJR7baRz6qbAN8nOZdvhRtsrPCCucgeoYsau/752QK0wnftqwwiGaF
ucNll2FVNe8f0srzFgmkz+UiwD5rnu1v0aqPdL6zhA7KaMd/l2geMA/gdwUAotgm
aZbR4jcJxf4Ey6XdAWIQLgW0V/C6uYLHoAyktDtAZ+3AnktzRCERWsZ7tgZ/C78y
2Rszsn5I/BKuBjQTudBYLFpUXtCWvXA9MKjiadpLmdD2Nw/I9CGL5+qx+NXxNKtQ
VwkbrSsELqwXOIPFF2xZ4rq+MjhaaSZfrg02PBT7QWWg13heYWlKLqrtJXuMpRQ/
5Nyxbh/liGbKKiNqqJ8J5gQ8CppuM+N73FcoavEmq4/gLB3IMCQ573pxSArfW9cm
riLLgeZYUKwVHnYYKPpsFvLRwAC4SRsmgm63Y8QS0jtcKbnvMjYBBT/PVOUIrfvo
qQaeTI+CG+NDRLrFj/s7+h85HqOsoZdHpEhXHe1ib5vT7ucgHlgokKBd5MocgITl
ZtHE2SJC23BlBQra9tjSuCSFsbPSM7hUFQaAeW9wercJ740KDvcloog2MsdSfGn6
+dmikTVQmlhnKsQKegLboKlx304phnL9lRjYO92QSl91uze1Gqj7bF1B2hxG27KY
DsAaxRLrLQqUKk1prD8WLg0WyaMW1ULjEB3qD1PCLtNpgji1PNapAIo08f/scpU3
GQzLD9q2Kdb32ngl/MHQYdUeqYuZTO1MBqgFqmj3rpx2902dI6v/S3OjuUWvOw1R
uIGCeZt0aiPVZeDMsbugfkJlFYfmgs6lweaE0uU0vUbSRP+iumTKzMVex0otFLQR
ba2sTmhXmfqcbpZLz0NPooL1SGavLW85JU/28MVaYTDuYsr2rbejU6vugPX7NVUd
ezrxyfG8GojDLm+7NdPYXr6S6nU5Nhdrai4YiCWaPH9CKb84zXaLZRjhvzDA1uFs
2cAk2yRwoF6TRB+yi5Kk46Qzu+M3u8oyR7l2z8Jxm8Fk3ALpKPLzXlOToX3XT0Ox
bnlvXh0DdjIqk8Dyu2dy2epCeyPEND5F5PD1IdhYl4iXsLZSKL1g134/Jng2jbSY
NE8+lZ9Iz30IesbBBZ+Tr7G4/5bGv0c0ws/3P3OwTRhBlaSqCaamuUvI3OdC5X/8
WVegVAS8MJTpWItSC3NaQqBovtD5kKz8KfeNEEBF754p/2U9ffS15k+HagS+Ygxp
oXS1hMlSasq8hZ/LdTOdxUzNU/ofcMMMS7V1C8zt3/JjrbZSs9aKqN0TMoB1LKA+
FdiU8mGo3lXSAVXo/HCPQiamz46x6Z2mXrgdZsLTpLBJ08tCrxhfHFoqznBUHcf2
vC86cClYjrbVoUcqBJSdPYR6zzXsSF2qe7jAsSItcbGSp4hLVI6k2UZTEvw0w3hq
cQ8S/MxlJdU2ug9C8T+CneUh8P+FPnkygyAnEgUzUyvutHwrtFpNzJp38x1oHFxH
oUPlfHETNb9aBoyWb42wq84Y9Ju/vdbtXCUPekVSMTzp/P2YXpgiti53Gor/G1sD
jeUPg8xwEZn3DHEugPN3HWQbn2mnVkl7CMPmoS2sYk4Ue9LSOR0xJV58Av7U494g
sPmxrAVgy3qQdfd+6wedK9U7IiFSEaSg3CRBjwOF59iMDdoTnxVq/6q3p32wCwCm
EJijp31PhM5nJT9BEO+7IFD0Lz0TORY78iunfZOA21Odv5WrStf4ITa6MQjDgDul
gOOhQRdpR5MA8aMN4rAKFWWPQJLETdeWBGIH4+swijNDhW47RA6FhClJNVzAk8QA
vkhhLFqd3vcEBZ8kP2bpBy4iAVO7+RLju9LVIEbKnnf3Hy78HiCQ6qjz/qFdOIxC
Zk23rWo0T1SszPDu0I8VEWpRX64mjnpCf3q371Ppf5QssEgB2G/hI8hYEZ/NYZM6
aZhA98blubORvsL8ZidvdFJQDvxeny0PPl9ybw61g+lFwD2o3jVxfMzfi72E9gsb
fmbaYfgmATIU+hAt+FJj1kxL+mb5pMotLXwko8p+6yyJNGoWEso3HNKA6jY1j+8s
Gq+2eT7MKHiNvskua4JXxM8BR5wIL3mZVxlDAnw9pIXyaIZQ9028fNO7RbFgjLrt
ScKzm4I66wXTNIbzUsRnVjljDM1tnb57OpaGds0yB8WLoEnIb5LrAvioaBLT+cyV
pXYRUw0V1n6wY/b/yymFlHJDTgZ8Z6QnWYpcBSDLqms1UrVMJsLKVwLeLL8esV9i
enpvoj3G8xGZ6bMC4DU7nzEUFpKAlKyaQWIonE3BE2Q2v7koxYe1D7xyeCcCzTab
eKsgfusee6AqKqdHIcn6x46KIGPmKwkYTUINnd7Xb4Et9f28eiDCnOWZhRAmGeS/
TP3Ek2bNtheXzoNFM4wTnloITmOk3twj25MXYwXUhSez2eBFaB2HE9FRQVsvfZoR
0fI+64/oiLG0IJfq7z71o+hz0NPN8irt9sFRSVcJNimEyERkx91fXT+ZQ+YLytsW
SsRPbG3XEJDtjVIhjCylB9nKposvUz2u+glRWofaA9BpHWyP+l7Xu9v7vWAP3elV
aS3HFefvpQkrFvqZrtNx97gi3nfZGvdeqGIyg3lccrSGwWY+krq9E9TU+XSsH3UR
GPzX9dsNFrqojsvy9PpxamS9YFS4g0yFC864UIOxyq7gZLAPDBg/Mj4K17sE1l/i
zplhy9BMNRnqoVf7BDBGs6fcI5cOGOILifIwVGihf5eIv+J+5w9OJ0IQ+cqmxcjH
2gMhpzq3J0g/LEEZsnQjK0X4ebiOOCcrT9gSLijR3xobuMVYZ2lhwp5LRgO9zgaq
VkCV51WHTY6G9OAB2ur6FgVw1apIzPA9wTX9oNjawpzPsKsgM5KjJrD8J08+q1p/
OrERzP+ZP/Z17+u9r/NU9jyezxDPyHt+VJ1AF6CjVPkf3ZI47JDjDAb5kiCPyMMn
DG5GWNcbivHc4/o0Uxt420MNk+SY0JMtIZCa/ycdtZ6WA7jxgovbYWMmJfXwgu69
umbaSOM74Aw+Kgxqycbtue4LNyULrHY/n5l0Lz0K9LbVSYu5axjfEyiHj1eQ/CAv
aPqwgGUderCVuFm80Of41tLddJ5odTCUk0RMwV+6+q10v2niNlbNbS00BWGENKJW
Rgc8NJ2+SZLn4cmgK14OOACR9AbNHPVwFlHpQ8hSsb+s7vSpc1KP/1naIsSjuz2c
NrbLJ0I2OyUTTfZYazaGLorjAc2jQ5A138pWgb9Z1fFl6OtJvtfFvXvwL0OgYzk0
qQBSKiVICKfOZnlHMLFIjG7A1o2heYAa6g/W6hnM7jpgafzdn2FW2aa1JR/wLDTt
yPk186pPhF1vhwY9XAqKf5g7MGU+Eu2aa8uITXeQHtOUqBbpNUAC/NPFPYkFxb1i
Uk4hjcAwy0a37rAAwsRCHuDbye2GvT/uLrQnecq0n2HGscjUX5wfhV2rCEDyo0CN
g8jmAX6mzTczGYVGkxbwIQpKrdNoO252Mm03Argf59HhXaGatqAAM9bMMaRX+S7s
kqbNj/6wEPkIuy31aUmPWgdeZ8Elwr8R9XwXpqmS0ZJgxizSLuc2GnbBK2WfJAHq
4PJDghELQ9BAnrRskuI307YMu7JMYn+kTU3o6AAeI8X/75jmOZ7xIRlNxNPgagLL
9GMeQ5885o3D8SDK2YJSCH1D8f9HF0CcrWQyT1B73UXe9cxiF3NqNTurHkMoWIbB
eOZz3/ZEmXN737JhsVzh2coVkg5HituXKcQN/pEpMfeR78KTdqiGBReOw0Crt5B0
lC5e+P3U99bzPfXbz8R83jCZxC3m/dMCKeQyOL3TAiq2cXWfYC8+ADHuISxe8wl3
J6jQsLk1z+VPWyEwwGk03PUvfVEIC9MoHpfOglfx7bJnEEyn8B6tL5tT4mB1uAYj
InIMOwPpbZ1OQjO/yohrdr9NVgEtebkF5LBt+D2cQBQSfuAhdbtCoCMKyTnsaZlC
iXaGF0R+N4ILVQZp0QgWy9W/EaBSHTHMQK1AMYH90OELRjm8qOA53bV/kVOmamt9
TLBrMDj0zelTR3zRCv/LISGbAxOJxWvE3KJ1PQPBAVcw5OqcyhyQCxiRvqg9EOVs
wFIyyG5344ZPV4w+pxTwM6jWcgQIPODms8qMZj35C39umt5WSWbGCBEpbhKnu48j
0sXo87D3YBFgPqUd33cUffFeA8BgKOyuF+Sr+auQpePVpjYxVWAQ8pA18M8pNW66
uB2xxQ32PlQjKO2DWwCx578mvArEtUeKzTWiDRSyjftYM4OvViJ23wFK8S+ScxmS
U96mV6u8DGiCiNNURSNwrs1mX+LReuQoWWIAGIWgC/wP4qa+xQs2fzwjFhUZ0W8e
gkXSZrb0L9jlB2DSpCPcQogtFY+c6UTc6TwlVYDAYN/UMYMKaFTXryl53i2QsdYt
5tv3wOLN9Wca4S5n+xNXlo4ZIKy01CuMqaSIJutuTAdfQJxHBliBPLRGIzW9qnOo
YTm8GluC13yARiWhUeXFXVViM8KlV8O+B0fm8uaLUTch5XUupmdhkcuUjTCdPaIk
YEIDtR3OeJqjPyu9A1NrI/u/Vq3iVbEoisSXYbvO8L2qM8mg5VZZF2xekmrgqZXC
vIMVMUP5Ma4BRNXjIobRMaSAJoVr2w8cptQtjMgNhO15/wqijG3jYY2wq5rkE5/+
cBFbFB+dk0h1eb5BJcdvLQuE+bFVDwE4ujHXOpEwjlZtIUb2UE/aQ8qmJgHjPHV4
lS3cMF7h4XFRqgijhRpmzzgPQrdfxWfgfMc8nD9Koc8zB01SimDjh6QvZ41YG7gP
h/W644UQQV8FHaIHOH26+z26YbtNNWoqYw9nlK9g5rrxMvzLsUeU9g5RyUlDXTaT
r4vVOKo6YOOOv48eLEvj+iB1lSEF2X4DxfUMVJ9DXJSjXqcMgo8VfrEAo9HiuA/h
o4fK9c6zmjfEc0Zm1ztXcSKv2k5iQbSnz2nI9bHNmno98bixnjT8ED/tPwBOU2O3
ncFOF4J7t6hg49NZwz0HATt6tRlm3voRdJALIc4Qn/KE8G8aJS/Sp/yxtnIZQMb6
gGinWu1dZTIe0e+C92M2JdpWCP6VmztwfI02iMTukySs4KUND8ZWrMKSKNdL7/DN
ulQ2WBWzJSujBsafxXfQ7beJm+MykBVQhlDCs21MkZ/l7usbpmdIci0RomsubjSY
EB9mIPzXB4GhyXmObXbsN9HC2TwpXFKO+K0HGSw6VDeUOHxc/TEmmfnhq/Lwf/Vf
QaJXTeNmnKOaeC7C3dL7aBRXBSlWvT73AFcYcRleVFJn/z2HsVG1lBNS1V4lubnu
guUpfbPq9VYz3j3WJdkhCffBW69fj9MBLcLL4alv2XMP01YpM1tkoYdLBMHfkwRb
pQRx/sc86D2RP4iRMyOgjJdwBJwGeULRHdobdQm78OnDOiioq/fZ9NGygjLzMjD0
fvcAR/m3CUsdG0XPjbI8QiZ3nF/OSUuFV/GJqQsbrjhJB6KlkBn3+NpHWay1Kz7m
a4NbUdAYbvuOOKsG322uZ1+AYPkoV4+bEsE2p5QMoDGMlUdRbxYvkfBzw2AbVOlz
O8H9DJeWgJ3vCmyjlrUXELGmW/Nz5A1OcTN48yCllFnxYzXOq11lQp9SbpMfJm0e
gQw5QvW0+eGoQZoZXBj8eZxkOANDUZWRJGRpxqiYbg6siTSoWrQbBgn9MwwBflNU
r1ko2w0xQ0AzQwYc5uzwPIPA3Wpvpfj5TTtrgd7S2AK9zvghEV0nhMOnl6LQmJWd
/AvV4nNwNHSPIahW7iWuR2RiG3MSLELRFdof2kP8flrjLnnOKPXWeI+L6Ula2WF7
EF4zQIQSsSeFhLGgfdOpdpVOcVXpbNCnl1CYt8nwf2EOD4VuFebFoOdcCAD1kXq9
gcvE/c21PQRaaymuMXQW3bUPUCEE2VhPCKJb8x0r7sKqDlots9QVnrf1LNRvc3O3
ngvg6EmSRozLl66tDWTwCzBcDnQonJxQXKYJ9v/VIK5iQBKO82BKlL5h1hNkxkb+
f5nmBsH2LsQxWszUguVoEHdH60VoQrVyje4g7BYrDVzY/6HuNoaiczoG8wvdolcv
iEOoCmBqzCGXIIX143RH0MH1pSmuaTsLLJ00IUu5pZa1zRAYp7uu7t8EvxGZeTPp
FIf1qNqW/lozbSNa/2iusNK4vt/9qUHqGroFvBZTCIMN/obYYVZ0k9nuPgjBD96h
4Hd49WdDfCc5ledz9il3tnvwKvqdg6QalZcZnDr2Q0BdCwBEaPZQh2kLTLK6vYAI
pFUbKRf+OP2CamhTCGB3RNI0e2IM2c44yY45JRXhwY0pSEit0qDkC6H+AaEYIwD9
oBkkiw2AubgjGovr/XWdJSNEGAfcWkOxy+Qf4/g1+Kr0KUEJfxx98EJFWExeIswS
9JRqW/ItLQYIvJWOiEhaUOpab9Mx6e2gwwDEeQ0bne7aiM1gioqf4BNhGtTVRTPa
1m/Ls5J8wZu1ocp5wYwKbQ3vfXCdsMf4I1v4qtk1YcMGvKli4BFhCXABzK8djtou
SH0gO2jIU+zaetNr6KKSKsv/hunoC6fvoA+PKw9p6HoXBVmOdVzNUf1n21FIfDKc
TnoYo6AH2LlOyhYwKloo5KA3RXYHaUqpc7R0kbq9mc4gFYmXDyRXYaDE3RPnOp6K
ULUFSgiV5PcftCjH2yBgOKDeXrZlQ4/le5zX4E2frWI5gJVu/mdxWxLCCZAXy2zH
isB19L/4t4FV+dLCY9/uhzRrKx2Ua1GBi+anDPrqLbndcJyQXw9rJkqiwq6egHrC
zAd+/cHGxgTBtSJU2pmaWI542okbefyEe5JNThT0b850Bs2gCh3nhazW5Qtgr0rT
w+rVxOUaDP8kxwJhIWHHylB7O1Df5qkmjIXrZatORqu3RyCEZnMcP0rr3eFH/a3D
bEI7j7hPLQQgZxKYQteE4y4sEwzEaWGkQ3ewVFC8D5ijq25OaY2v14KTfjzPTgZL
i60hcxCh+k9qyO8G5gso5QjwsyfV8kvYAx6UWheQ3LoYbddDEDuR2ofzjBUgQ+Yh
fV60Hdug9TQc98BMFXOF8V9M8Yz4D9vcy+tlrcw2LthILGFiXg6u1lnSen8mPw+Q
nhMKWI2BBGWnDG7GEbtRMnwmodzlrpL5enT8TV3Av0eZaXpNWZePLn5aMYCasL7G
SeqaW4d2NumSeiSwz+LLReWYUj3qd5Uio9Ydf2XIUv2/cn6HDE0iByxHG3q3XRXX
4yEowqqHgPdzWsXQqNX6HadIvIcFO8uPG6glPYwu+7oPd5eQBv6NWRjkJ+9jZr4P
xM5j29gZKjIsSD2F56DnRgPjuiY0oLhZ720wg5o7UkyZzuUogWex1atFh1CT9zjT
cwKjbrIGybJv9m4aQjY5hqiBrUgcpQsMXDhy0Md8mBGmRBSVKHOYZ+eoi3mUPtkZ
jI2co5dzUxDazi8Lu3fTpoRJ7/xnXG9WRlnIx3khQFQ8GC+5o++jeADxLv76xPz4
o2Ggm8Uo0fNUG6/V38xz6LE5ZDYjiVWXG34Jlc3GBrj5n8Igc2TO4uAHKImYlXU6
n1NpOzvWbXzTgrslGe3YNYtANRaTn+rtHLogUGiApUr3Xi/cnvGO5Wf5jcX7RjmF
HXrmj5+eyicK1znui3HmA8p/XepCfpCXxKfz+AnVL9r2OtD1xNTS5IEEQFLNwU2a
iLd9m+qXFSGhJY0Et4bXEfUG+Ca/CFAJN22j/U/MnOfIHxKHk7c6p6ONDf3N2OMW
Jkd8U7s/SuGrDGrtbcDyInTtA/kv+Tp8Xh7c2m8tvHMrYmGKKZgbHZ8vdhsSv7e8
EbsvgZjh+fmrK60e8QaSiJN2b/87pYL0EKDy5RdHq1VScWlvCwnZH3WKBCg0ee4O
5biV5VGMUkJp3PP09l81MI/gW1loTvi8Do24wxDx6ymo4rwzjT2IgTO6/pXE6D3L
c2iYSJ9+8yKLW3HmrJV2qvnnY0fN8ZfMznMm1E3Ba/wnx0SkYlI53nZxdRN4+sbC
LuY3wEKzXE9vfgXRP9W9ryM7AJVWQZrLfQYjp9Pz1KCaUpeuKdllQu9YqEKp7i7a
hKOgRa3S9LX0CzVPxuzAbUd/AEQzElQVUYXTzirCEpND9jsl7byNf1kc/zAXm8WM
ugEaqPGbOyAMjgn/Y+4RS18ls0P0Wq7mnpbJJXgHZkWdFg5uy0MIkftcrxZD4PqY
RD9CF+nFeacIk6hV3qzowuO+Js5nWGPXvZ6vEDjsl7qxrt7nFdvRDoFILOmdjDUV
+NCMRO9NqZaRACLm0jY440YJqcyOOVLMWRWM8yWBDCAIMA3GhqiHVYlgup2puwxG
Vy1GxXqEBpUvv3hU6BXeAQBmH0FO/497ij5MOhEJLx4poSMC6fsOpKWYZqh8maJY
jUtEu01BCtm8Ny34BO7CHlgYPtP5/xTy1mGW+sw2bPlKKazqFjn7lbc34T6XxC/B
+nfwwpuqLEX6oIW10CvNQtyeFD+oyjNSyK261w7irMbclV8IfFfWw0Xt3vTR4Ghl
8n4lgXOkjRSVp0s220Idg2ONYH0FVpWGmyDINuONyafugXW8fLlFXnJdlZfxnlbJ
M/AU2IddT01yjZLbI7WyhnivXDlEhiRCibZZQwVsoS5OibxObIERFPeRwUrkiFzb
JITz7yjqbYRsRF1kTHrUwkDPn83NjKDtb+SPO2zD2yoqEiHYFf7XHIH2mt+oGtFc
E5x2TvkYMOaLXCR9AYBe/ObJIRvWx+ycggqgtRhlnXdejmhaiAqsmT/wM3ElNYOI
Q/X0RNt5HrUAfTmR4TctYR12ACEU4swjAHFD9A/Rwk5FF9qLd8kAQ1oPsJM3EC09
RWvxmyggGDcx6UPeu65+DilGcFy2PXgvjMt75v9H9xH6t3P2sN3tdwf/MrAdHdGF
y14Ct9VJ3lPHvAiuGwISUXCe/DWVacPuFUY81h0rwALH7HgIywlIQ+H0QF6VaP0X
u7i2YgaYWDWhfbwJT094bxwcxmzQSf7sWvHq882W4MM9Se+jQb68DBMCqqIHH+J5
T2L/8/JY/8X0xPHuS63TsN0mUqSvkpeMe6hMsnEyfeI02WtiDaisUjIH2SNhA4XI
iYKwG0QE5fpe+EESEgxFo51FcLr+AUeFspkpkkqnRSWzaZBPOln5MV84eFwtljHw
VlqDEO6oLYGr57KyzqaZP+W8q6KZQr6inc1Gv+strPWt/pxq9sYInnDXyNh4NMgs
1zJPlDre8DRPREhZRtLKbVWPzV8SZb+jr20jMeDACnbHZyUgF4uAiGKXs1ilo/Pb
j96KYowTcr0Czn4t9DItu0j3vlmxWvRPXyfCkXRvJo+IWZ74qtAdl37jkkDiPgoS
Q8TaWgbw3+nlwW/PtVrNbMfV6SsTA404ulJWSkYs1t5s031OFonpNIgTi522o49w
L5ymFoveGSN2g6msmg7wyCwx8mZqquNLZJPaE3hqfU6ux8lVleZxlLUCZZs6oKFR
YzPRbOXw/XKgEJxorQIyOaPeFBBPlKYcaXwpr+pxYXY2dzenGwB9VRBxEVtLO/Zy
sfJDvciVmmmAxA4VLAXQbbKN87OHC4Hte3XHWTHh5wrBu+tiVUrrroGWgwNTGwgz
57AesPrc+unmLH5XLPloMzu6lrWC0UjzdNrSMt7S7zubSmrdc23e4/XKs6LOz3Vk
KKmGG5eBM/RIrWN/jlPSb1G8B37ovp0uxdCWPOkfeDJT6xcdFDHDn5z/5Y+7z+vZ
FuO9TYo2RHavTgvvUC7t2hg8Iu61XzJh46kTiyGcawpl7H0V6VS69n43vjDkf4Yf
LlD6PiLvVV2GfRx1mFKUfkwpp7Z1gyXRYaf+0nDqsYcdTmbofDitoOAy2zOMUpOh
Qn+Vs7FSYKTik0yEW5fqpKRpoLMeqIDukZ6+U8o+HYqJAdZvnRwWGOVmGTO9VkSE
k9fjZ/Gymm7jDJCRdqV3Lv1ghqgr1DSZqHjeXMeq9PndM3oNINzgvQpegEIgyvpm
dotTntwu+pprcdSqNmmUh5SM7IWtyNvaM2YIEFUsj9LgXjMYmG4EPvIW8CpYQ/pW
ADHtbkYX7T9bqMpnlQkrPIFuIwqi6h0DgkAgTfYDY0TwqBL0AoealGgIKUNhmpVi
tLesvzJZgPQQ5qJvs9U0dl767W2JbdM6x0uTSGnNtMVxbIfrpySXLX2XuPJXn1b/
2UI1VowpUaaX8htfRIRxxFK7JvUty+0s85I2wcRdxSixm3MosOCkj24r8F/6uhTQ
vdMccuYPmNb6FNtK6byIdzA7yf67DAPXD2kqgdkjArTzj9gQxwO75ocZUVSy1ydC
6UkEsIiVqSLl78P4JcYu8EUMdLGTx9otAXoqTzCkz14sCiC8mYiLVm+oaDzgrCNQ
unN8CmEzfymRPzMDaMWonfANSnaGWHACsl8EaITuVCJwRUSyt9/cmKxQYdCr4811
kDAszFPmKff5LUyMUBo4BnSlbxpMnLTyN7y45/9QwfLmFtAUqGnMfNaM2MbcC+/R
ZwNbckhMxEhziURNrKCstlmwY689the001JcL4VK4KHD5VuPmrKsizY4SfKiWEXf
82stcZ+a59/5qcnBtHNgg5pSF8qn3adMIRhXAIhWIW9jqUfbEMuTu7JMds/Vd3Pu
XimtrWoRDoqPqbP/LPab6AoLc3yRdYJuMdmMs+sPqIqLuWVH2Kad7CRjm9agiJjg
bwtzsHCliwZtxp4+lG74/W9tdRE0CH/UXn9GqIfACr9zOtYle7Iv7aRdyQg6I5sG
Z2b+Vtwyk2MY19PI4P5wmZW5oJBbUKN8sRtr+O4N1W7s1QRlXY7eDiqgmZ92mBWv
chLoRik3SGwEUyYI518n5H2vAnH9Z3aW44hPRj5EvzHDa2ENivBUFphES4dAPExV
dNQyc3afefn+Pi4nVcadHBhKQHZkSOidtpKujxUDwuj+R4q2sr/5cVSYtt6eyouV
fFQ8KZvJI4EA/PCD2+Qj8+2bvivlTun0azTcKrRQMMNMYUHXH04ycUISW2ziMkbS
8CYWPJKRZMLj0uEyzobp8lP3IZMaNyE0Fi6+kRxEqUuXD1589aeMFVAUN8ktzmMJ
+q/GFUcpN7GXncjQLdCNRc0YpnrbyRwFqzYcaFJgOvgLe3fAcoxNJHDyVYrqgERU
VUOdVoU7bCJhYEfFniGn3dqxbUg9GhHcqHzk8isD6af+ROA6QB3GgArAMWsA3xN+
wtZBlKLt+nQLVskmsRrhIuVn7oN6m86NSGw1vMnHVOiPWoVd079wPD0OOOHe6DvR
2DC4xJ/LOYpz6ii129LfmD1E8L2xjHIP7zhOR/u5s4mifDWup+5awdDVyVTdcgWs
vtqfmbOXSI9CvjF9z17vjbeCvy9DJDYz8Zkqf0ThY7yuv3lzULZjCqVad3KhwVIN
PXN3cmCkXbIRBZICGnQEXPds+B2PzA1v6LnQoN+EV3wYEEcduIid/+8hyM5H1Ba1
uFAU+IHwEVmd4G3HdH4TWHMke6P3gPwJUui3nH8o+60woT4pd6zYrLo4/5+NDl/p
ivgOCdGOjitWgFRObLYFRVg6YCCypGqOpbXW1T3SAflTbNLqBh+H7cYIkYnVBZWp
ysYZAM+zVqDemHvQHXpxZBgq8taehF1GR/OV/tCa1WdqVCRBkja4O2BK+nTG8Q1Y
wwigONopj9SsEGvD+XfcCh9mskMZJTGfLJPIxkoyyjwnKaJufP+qZFhFh3iaeEt8
zKwEkvKIJJnqtps+z6cu1UrVhqIPlmtyKbgCgKzvM0gqYu80IFg9KJVu3Lr+8ni8
jJZDVaiT/EAK1O1w2G2Z066BROGTWvWMQx5ZxNRFU5bTLkih+4w1yjfRyQ3sd8GG
WDcsAE7/UYBnu+Ouc0RxADp0E93tM1ihw47j1OlKcgzJMdbRYOMZSlNub++g+UDz
tz24vsJ1czL+CxkhKeK/NKVWQ+VeC1zPMO4q+IGzbWmikgRSWssnITUu5TnnEWZR
vC4OSFzW29upCcC07FCzaFuzSwmFURCDxBQaIEzYV3giENizb52+pFXZm8Bf8SOb
6atNLzfY9ql0ZzpBO8RmTh9f8Yh7pJq8Br1aZcNY5mTVaNXD5feeZqwgw7ja0A0R
gwuIPpdq5y6bonf80ExmMTxaOLaxv99DSj26ShTecCdsRJOP4xIexkX5Vh1vnXek
N3ccEWZyqENq3pnL4StW1lBqwW4jweexJ4gP099i5H/ghiC36j9YrBPtI85GiAYO
d8fUpg00f64SNZV2zmLWaB38BQaaPm9lXnUoBa+VZviu5XlD15w+E3wmPC7vvru7
WBiHHW7yC3WkMLzF0Pj1HelGTSxtUCAkotzJPeJ+pAlHQp9hEjJsJyaNma0vuUxL
Rbd2vjG85/Qti3nM4NJ1e4SgPsRPeLx0z0vZlmNInbiRB3C/DBhRIFDGcmCZwd2H
CC7GKTVEALMGvVBjOcQ1PTm41k2VZkGYtyUSsfcbVif3B3SS7Ci0mbqeRBJA/qZM
ogMrMivNx9UAj0LjcOKEIY+SeNFxBCHuXlJbl6Bt51JzKNFLzZihNnKeK3U9jQoH
DdRTx6dLWSfhrD+bMjURKjyEY3DXTFhbJP8tNG4hWYKhotCMx7zzJ6sbaowTgXP+
Svj24Q4DP0BRNNxQd+DFxJKe9n46umrBJ7BYNuh5uJIf721LZF+vbqwFby3tD+/9
krIngSYMioKMmVFHghnXS6vKwD5aXAcln6e5xgsGX57U7O99P2124N5kVhiNzG4M
iq7XAT+SPYFabvJaWkxEeJH9ZbpnY1yeYCwfl87NodvbEwpNdFAtRgo04tmqd6BA
f3JqCGKenF6nviRZpPjdQiNggDfC0DQVDvsoGoaiANivDePAVV8YrQRrA30MaIx+
J5AsVFk7i3x3qaovSzK+bEIbuDiyl9Lq7D8YmJi4IdFH4SfOiHVZVN6IZQWhPQ/f
8f9J3kcNEROTXB3v7GbOCEUEpGqci6yiDqv6DK8nfWuHxCA4onSyptP5MOrbQEa5
y6YWkAYMso/sG/rNLsU33/4ZEj79LpV4qR6+uP9k0SsL8/eg4jfgjkYv1Of8JU6w
I4IcKcpRCkCXZduHJTaeR0aGWIPd9GlPVGgSsNxhfXRnaiqopsGeuO/qXP3lrQev
W/kTGOQxmT/WPLFjCqYxKw5pflPUkM07BhTrfbMz83go3F0LDO9S2Uo6HAlLugOy
EPgWBNKvcRtDhb1hMz0i3q01r1SCLQ748CiSKVz+z+5/jMoE6WDuAnpd9pLrMwj8
2kdWd//oLrANppKaJnm+qB2S7aSL5MES1Q17L0ty9yiaDeirxPk38oDetrAiglJk
JjKXPBujApDhd8gLJkf3ciKaFwoFO4/6Ujd1nRg3yvFpN4R6aI3tWd+7NAhtta3p
tWEd9T8VXyxHWt9A+jDTknyJMwnT6rK7VV+6daI4oPMdgeRqq42CN5gqNewI0tqz
lXMDhp4abo9kso0PiLKr6s3AHc5U1gpmFQnjUL4nybmhjhag+EQLt+K4A2cfJKvM
Kcl0QcqOpFqoZxJJLIOSA8p5OhU1HqXa5vGxBXRtPxrKqHahHqCHY60lpuLaISqP
u7gMe9IzvL6a58Bbh6cyKqrJPDV77Ilc6NgbllJQUIJCfW4+vXR6VJAgeL3aAtqc
vl9to2s++rQ0b5wZt53NVG6dBze+N4uUXtI85BR2cyqZATrxVxUMvbHfNxXgWNA2
vm8lnDKD0SE9aG7XrWpzxgdGLnnrhnlzcBP3ayJbBhGp5+KwIV48rV+4HqLd/VhO
/URDqjtcDIrSSNErrhymwgXuq7bUEkDhk0zYWlhnZGB5s9MTobFIp9jGFYf5kc7w
S7MpmZjnLIstQbQg1PKBNETcjDnzMhFmTl65kckBWLtHcO0+hINWSkH7rWtLS4AW
JmW5dHgtwNoNnS3n3ECh0KDL+BSbx8SrU938CDw2tL/BLjO04dZlRoyfQwSMn7A9
AqJtAr5s5uESQ96gOFt1gLH9esJaOp5dUlikAIJB5Z1AHdCW0Fqyg5gvSNR1NmKK
BNByVnT7ijTJa7iM6pY8sTbAY5pTniCr4OIPDanVX5JKVQBUWeAI/363HMrqJKLh
USwjH/UI/2mI5xhs1BJFR7ZD+CjDCMlnfqytIG1dAAf3LJU3n+X6X6TM2VYZBc/R
MvIamJd479yERzmlvrEZPChrHblvQdJ4MAv+gXThpz08fud1+qh5YaX0DkPNnZM/
KGkT1gnIzpSngCGbsR7S5f9yme7NeSzZzm8FUGHwXTn6ERrfx2zpsYcUxUCgkWwI
6Hnzy1cGH4HCxHKsQhhRhV34uwXn2ea15sID4XfsLnd0c1keC8ARAR8/BmmMpC58
Jskp+Z20O8Apr4tMGPXZpASWJM3WDVApgq0hGvMlmHCs3HvKTJKP9Cc6DKz5yrvV
qzJjtg6fRHJ0n+6Qm+o34WQS8jq5H/NipNH9MNXnH/tvEaQKseffqwPFO9TNg9AB
hgszBR8Pnf3EOx/TVgLT3AH2HUn2ignixnaX49Gg3fjIlJG/QXDwJFnVW7q6Rar+
SUgvLWBSJX0WwcwWORiOxlat1t5GHzLEc7gYSq5JuON/sOg9mM6XBxvj+WMRyK6g
0VrZA7e6x6Z9ZjXRzk7JYGS0F03yDR2qHg7A6hNYUQoXwh1eDUIpQa0B/GSWfGqi
W+Aj8fTqhI1xx4YJqSMsh4Nr9OwlyBksPewoueG/BRa2IKCLFsgj21FSkXKu8xUP
7/I86euDvpjsCWPPk9P26xCmx2/yhRF6B7Zd+midWyOEwzbgtsnJXPDWEVaUMBlx
3/zOsJC81u3KDNCCfBEjXo6DKGPbQYQMv1vR/hTKHeS/jKggryTkX0//SMQ8ywpZ
gSXiMzcZcV/5tqT1zBYBDhNDuElbpvOjaIA9s29qlxhovnWeNCWQGqzs1BEUfk54
jicOFK9DCSgrI5nAlAoJneTdTzl8HdnMGgElM7atwr7ZlMPJtCkZRWOkM0A3GG3m
88Cg5blqOZ/BG59yUvzKzX5YcPLtfqRo16jZJb/OO084RvQw1/cPWA+J8jbEdllB
I/ApznWQMQGL0WYX38PpjuqV/ztzg/9ajdYOvyNa58wimh9ZofVD7xVIm7a4dUiH
7ryZL4bIW5NOSoz79VtQR6N+KDzzolTujiH/qslMWxf/3PbFNSsORpYWIom3GN0q
QtZItQ8Ezs2mt8rcZbxcYf8udEMXjVL9Efso2TBgCvNiehyLuYQqJeBv6W0BEhND
kRRn+yVAwElVx7od0GiF9rZ4UR0iFeiVVM8KoreZYTPx8o5pVtoFB5xNg/92a4wO
+08M9+qIhT5Wch/4cpFGRu9oy0IiQkbJsOcZr/FiRYc9vn3FjkvQdxOphL8wbsWj
xwqIUUh2kgTz6QBvftD1kWFeDcH97o6rtIgg/AHJqsZKV/UNu1rs4n3bvelBz31b
rZOTrMDz2kNOLlc7eY3EyL+27FCpgJMVuXxKCjj0Hg94DRDED8rYGBQHfdxJPmuF
DlTjDdmGRBC2F2J7EB5S8QH0g0dgAOaGOuJIuIBWPHR9g3RVw1tqzG6TzOTAXwOw
BRguHi932UHthTzHPkmi1PmXmoSZRJnrd3ELaoSi3+XK3DMKJG6ibxqBpvmr4IUa
DeHYJ45VhRsuCFi0hBDPEvExWrluKXAoC+OweALBlHPnzaLqbcnHNbKXsjHjnHrO
H/+QjWjlCp4pXyczVgmDRCC8soofDGaF4NKEOnZD8wZ4fToNN6dEDiV9Z4Dk3h44
VfK94Gk6R/lm2djocEsz13vEDYdhQMCwSQcic/qDnlGa3Q71sh80yrci6kWiEdbj
ARTkxkmOdpcpIOZQ1gqzGVX2ZQhmthw5XcTL6LSE1RGthr0fdpE7kNGVw0prLSnF
8w92HnpstHIzkQGt+5oAxeoOcTSSvv9q1oeqd15bUQV+rzkURt1MMDnCNursX77Q
QGgsfz2iGT4NNIWNqqdgVtsu+aoKoU60/hf+YiI1pVZn8C31mfB/GPFHWaTzSzlW
8tws9Q0HQ+MwPoYx0qKILBJ6cNa/ZpPXsRwLv0jKpego89hzenfDcLTiN+x+FN9D
dhmQCFi4ayZvn9OlWmOv8qgOiHJ9JHx4eMhhTcbulEKID7NcBTaqQNntF6WsxNvG
jROPLIY6tC0c/FD0Bi/HrM7Hlw8wZAhsOaYk1F5xlmGvnb8q8jxO7ND5+rEFVRhJ
TZxtKE+V/IcpbqRIMd+Bsw++28Wo0L1GcXmTZysOHLI8Yj124bh+QyhiKe6lG3Ut
8CJAPPmbh738q2qV2zsG/bEh8oITZ3M4W81W78L4DX7zTfxpGSy21rjZVpBxKHuB
j6gyjbejGR2wfbEzdgmkh8BdalAdqzXRaCNedjJoDyuA/0Gwi75R7zc191VUivhS
T3q5I8e5zR9EBX45fShl7mf+7onnnDSunf6nvJL5EeLfercMIcx2mZZ7cbrZeN1J
pkBSleXxTUTfcjh6WK0vvhqcRfr4chKwRXfpGNuNguGvMs4CtAvgx/DVBWeezILl
afi/zhwFHUkdPWZo+2yhVkOnqzjzXF+ApMFQaJfnYwxzuOoJSS3jL+i/+gCeAcca
cFLndXrC5wU8kLpGwLZlgdBEaCnyN2VMoqrhytgucuER6LchVh6Sq2XPTqWYO41O
3As95RXGudzlwsUd7LG6iPegoxSuhe4bpzuUvvPbgteZ0svdDGTUoPfFu+erFr2E
jA6g5gS0aiR9EWY913yM9Ox3Crg/HPWkkIYJCA3LQyqxwI9ITZopPznwiNpO89Va
iJz0/9s4Q6xAp8mKZTYeWLGpXLZYLnbHI3gQCJI6HX2X3uMcqjxBHIgXJqSu+Tko
aqNNgUAzXhOEmnZPFFThc7YuhdFpjXVO+AHucagJGY/O2kxJjEraQqVSGKz+tRAr
a2McpE629zQ0b9imNxYi/er/bpaZXGTA1dj3lNO+dcrra4fyKgOh35KaexfHlUWW
2XSRYcRMBxu0He2y0EjRstPg3Q30T9PigfOK8BqEYlKOxLO4lAF6Vxfd6V3EMWQy
Mot+mrgE5KWgZKeEM17fCIxbWcOaBjTGph6tDRZsUC0Ilnn2uCifUQEeq7kI7Czx
yZJgf9DjFB6eiz5dE936P/bpIqneXpqdNDVIjzrEyvt6fRCVstzRahi5lzKaY9zS
pT3xqZH3S28PXbeop4qPhevVWhr6u7OP5o8IchktNkn9KxUlXFzRukl2xiyv0/CQ
o0xlY+n3fsCJe1znX63TPRfPCXlf7H1b/Tj5THWTArOtb+3XtvNPapQeLXAs/r5G
yyVKpY/YfwPiH+aCGcww9P6vjgWPBFUdpTrzRC1s30HKSMlvjvVanpKRaITe/9Qz
qBNgMaHcsJM1OoMBoKUsqwPzd5bPd13m2TWCTwB30b7vIukTh2L8FdNDVo6toVNV
ALUve9esi5FuKAnCt+PW+4Ao/JQZVi85fgP94bC8qPdm8vbJarL3rjW3NlSghImu
z3hxywLlkvamT/mNxWaJz+dXbZYOZRWiaTbPCuwA3RzM41KzGOpSJ1E83LWXo7Fu
hL5TTO//ecAG2Nxm+UrjSoME92RmVr7IjJvN0t4ZSmLqXCKvv5JoXW5LKu4/Kyhf
BEXZIPUVE8tv+Z9ePnh1soPHBuTJzb2DmdQvxa83grwc7VwYBF/kE+3HKi+nQaK+
BmhEzzRDjkRULDBns1ENacFImd2g3Q5VF9C8Bfiyvg0VxRfHxVLTm3Z60+3aHilA
02eJPZkMXB1heUFmf7vdhVwJjGFGB+vDgl1Bl6S3ifj1gQsbljWz7RY4KbNYSMrz
nsX83iXzeXSXfEr2Th1AZc9mcOi78py6cHNL7e58XYIe1NPYqrkn92UYU+XCLRm7
KyzX0QnSQ8DynrIC9nCHH6pO2pbIzGezUs5KSMos8M+A7YtA4OlStXQRb9omWex2
+2byLVZ2lBT56SWxH0bgrz9NYvaE6YL4bAV9zv/QtqZQxhsO/KisW2+mgC78VpfP
wP1WqxvEWXGCrDHTUWDp1E7knG8oCX6Xqy3/hCNqvO+m26L7H9zGN8ReAjM7AcKU
RYG7ynTYHmlX4xDKkVtKFm5y/Z3rfPJRMcOYQAqfRQ7MbKBiq4GOiBu5I7x7DN8v
Wn4GWzsSjW+NRl50N9WZ8AIelGhk9kV3MqDLFQiYDi/iW3gnQZufAuvhXWjZSQJd
YCgWoSi6iHngy14Ugvzo5zJfxicwGqFshU4BJ3eXrdeb3VSDcapMtrBAojJANGRr
sOwJz9EN3WgdCY6Dl2nJ2lkteG1vDDCfIyDuoUYsRl0EgNmp0fMFUu43DuUysNUH
3v/ijzuKoF3wV6Yr34qph3wA15sEaajyl/Rt76FDsdC43kT1FXY9jQL2PIWaBUHP
e7potzLdIFi6Dep3pCybapRG3UCLKtK46v5z2W3AB3UxSAgmk58NX1vSq9pn/mNq
V181EqBXm63dsCPOKhcf2Yn3mBWvwLqKHdoIsdbL2f9W+0pULSt2nWhc0Qi+RaxO
JGhMHRrwDQmq27D926JsLCA82np4ktr98usSrm62mY0IiIYrAkAy5LTNZWLLgqPE
P78Kg7NP9rgY9WhsJBsxE0JvkqOvP+TUVDjfUyKdt6jTTnGxQyzafG73fSSk9yyh
AqTQQ7TyBKteIlK/fXhdHK3EtUDUFw9azSOweQPH0asDPU5ytNetIlxHgoJVwdzn
fIqNy1JgZ3l3YKwZIBkZ3sB1g1Rw79AdfU0VjwfNCHfDkLhM6zuUSAKsR2QYKi2J
UuYgw2joGe5ge2XuXaxcw+qfxIi+Zau7V6s4PfMHE8G0g2xg6fFIPbffdgAHJgAk
PdKLjiDqAW3A3qhPydKKFKuqmTskvlVsu7mY4C1/pda9WovRKPM0PxZB8rtEQ8OB
wDTdgQX0wHpMPUwcr4fmuZHqW55EAeIyydYe9KBXVJ4ZLYkUSU1TWNqUmzsTmFAV
9N3/RDNUEvkHChpeRUU8xzjwXDGMYWxswtRG9xvSmsfA+ieXMz8VOIk8d6a3Bu2+
kQK/EKaFHh3k/iXqEqBxcV108d4VtG3SiRrQBkapnIZD1OkmEfCRjDkDKiOlMB2P
znbyT962JBOmSVlTLb5LEjvI4bZgQHVrzDF+AVBBHEmOTV0bBE28iivsoCp9GIYO
RxLrH1tbWpHYQewEU2eI9vTe+GU3A85IJn3m5SpRA+Y3rVr2P073Csq/rN4/4vhm
to5GoH5jG+9vCDk0zj5PrpvSCNd+FIP8pAb38Spij60dg5JsL1g2S8Aa8ndUbyPh
eusi+OKzI0M99vGr8pM+ME9fqbZHkGltZooN5mEfQubmfS6EGke5RGOeK69L1IRR
WV7ZJ5545jS9mnbkcPd77+22VN/4EzMWt2jMAPLMvtYTuKAmnBpOhRnknmiOxhva
LYa/x8pPsRMWZKh7ryOe01TSH2aZluidcp5WZxgV1pA+DEa0Qj2mUhT6O8DsVj7c
9Jv2DBD2l7Dtb0clyTfrtIvAW0ti4rYBpZ6tbofwEj8HPosyLwUf3nqO1558DHQ4
5Ii8ejRJbStxyHxwKwf8/eH1R5Mf0WFghFKeblQodupdBAMxjuZzi1M7frTGkxSA
KOjJRwc7ERIULmW/bZptLB3WS21t2RfwPaDwDSlM2+vGNfYreyFNxTz/m6IZxPC5
7UrYCFLV+F2ZKEyhwPydVETK9KIrciPSkn8+fp06JtkDYPHbPVtKXoV7TsCxdsfT
GuYXssCgVev8XyX81jEE3H+H4lRqfeLJDxtst4q4S3CTwvEb9Bm8QgPV+iGw5vdm
Ldz1ioAubctpLbMsXnZtaBAM715abdVfV82AXdOAddPjiTtV2KgMium+jWOynFcG
5aBMERLKfYeOjNUBT32pSOMeznAWk8Yp5pBsUalDLxQ45LlD4b/612J9B5lM535E
OrikmxcVsK27fMSK7H4l/9wFpCr/VoXUag4B5fOBm+VhtPQjCV8W3fcVb6/yBLOb
X0w+34IPMQ95sKLeIZtMbR1ldPh7WQJ8VMibcdmRhSal803Si85A4d4QeNmgu/Gs
wv40xzzKkVuXXH7ghrxykWzSSnUedlTqDT9k6Qn/zU5X9pGd53y1alsGaBmWXtCf
XyLCw8XV+Op9NUOUt5GTrEinLIskZaKmTs6Ey/jeqQ45R4bSlNK2J5i+JQifK8n1
DeNtqePnSQExcS5+cvcs41kD+PcKksIHN2DSYLkc9helPWN9Bis8F0hO4qcutbY0
zneMQYMhKm6EYoxMzYqT5ZOJf/z4YzomLgJFxT34YSo1QtpU9gqUPIIc0WcbzrIj
Ehq5thI0fHUQFE4bsCnB5eUZILiQvm03uCMzQYlIJbVgy/rm75s0B8DF8ytItMdu
TJCwgYQXbdkWH2CPzXHXn7xcd0aRZx6SemAEy+U8DdXo/GDVretweHULWcWlWO2D
FbTkTUL3bCkbFH6QQvSKdJTHF4GnrtvYusydeoNuNMO6dW5C0HrUazKvdG8rdy2B
eq8u964PiLwcvbvJpSO0ThWhUGN6XHwRfw1o7z1W77aYjvSw0wHx1Tq3ewHu08l8
5SusOSJKjVzPsaEsJECT8YsvUQf+oh3W5N1MmOVLp9TWcb+VPV5Kb1uuFA4MIlzy
rhELJf2KR24/gFxYj/gp53CTh8RcpF9082QlqsFR8LexTR5D0Vq+IttUknAQ41Qo
2MoKxH6I/3071jxhf45ywg7bRMyYLHmVopibzAX6UYvkE4KiSaZ6iSFaxfspslxP
dFQ0oSPQS2PlvB75EreIKR6hqqzTEZZqrZnCsDVxP67NnsS0ETFTjaehn76AuKgj
dizr4H0evZ1eWPyqvjRvbHvc6bg5iOEvFe/5kTO65PDf0hzaegsHXmj0Ncta4uLo
EX46WjKNRd4XZtUG9mRWDrfxdTfI6c4ClsBgQcuWoAOeWDWflqFUcucKy2lIL9Cr
QMl7OWIjVqfbuRqCgycI/SoWnqX1uAOAJPBmUEK/AAolDGthB4Io1lrxiP5wmAqY
dzOQ74dKpUPk7esR7Lsr3sOl0X/7jLTN30vTsaMWGT95BFu1Ac9DwrWZ2tmoxKma
d6rZwjqUJK5mAHtmgmvqe5KTltk6L62q7sEihejmBdwm5cy3CbbEB/sTBy89ivyU
fNpNu8RMkaPWSVAs+vU+UtluuFteKfKoqnRwLybY0n7OZf7iBIM1fT3dTZQhG4dk
Zw8DxUMNsOx7y+SOorVBMjVRIuZvOx1fgqTusDnbmyt1rlrE8HutA05l7tii+QQ1
Pgc9pVVj7aEbLm6Qgq6I3spIV6LgU/5k277nmjTjWmy7UesITXu8mysIGuVVR/pc
nImlr1QmQPGcXoz1VYMT9bSQXLUKU6lRERQq1AgVTxCaD16tzNWtErvZ7QX/enjP
O2bldzMLtAtAo2KVExup7XO2Zxc/Rf2sAuI3L+Hd9JrBrfd0UAzgG1M8aKKlX7jp
MbFZCwrRTqzPa7R/fZ9GgAKFW+1ujX6aNnXjAfw0rtANAkSB0ONfLn0Sm5uhzPSO
qtBMyvaSF9xhyDcBnoQooyDCwqn/xQ8C2as70l8If7YVsJJAhnhHw7S3k4w8mis1
mTc064Cak+vrMh5+51jrDy/hyEmf4jHWmXC4oPySRsNjfUJXFOzgc5imrBO6RSUr
+wObMhx7DobXKaweA3sMLdAa49ZdESfEbeYk/fUxAbDRlLEg2eCUvKCoAJ+GXwZK
ZuqSTwL6YqEitsKW2h5eYm0RGijgGcFwTVie1yLAm2zcGDSutqvMN01CCnf6LXtA
7vHf7HxASnrbo+iNNBh4Cqgg8Dsl5RvQmU8juzhHIg0Bw5ZZmWPopF1Ihgt7aZOU
sGprCilGoPFIQd12eW3dicOzwPho5/jUsR4aAXWnT0aJBAuNqUM2rDiVZvs5xAw9
4QZfV8rQo5SPeSZLs6c4qEijyNQKEJokcWBIJsrGHnD+4Ro1GQPni1655IU8039G
PMWQYk2C+CTC5wZd76ZqtDJAzd+1ROwZQr1grOeVrQvC/3UKdtj4smZuxC/bYvJR
63WF+ubk26nESX1/fcBflrmCvxHg18Znqg+91x7oH9WrfCN51hlGWJnE2Kl9Epvo
Vxp91Cq5UV4U+IUEmiL/8dWfwfHQpaQMdtwGkUdFpTeDEyr+hVQZst4HKpBy9Pgc
w5AA5hwUrTZxHmrjllIngWFARTvggLHkKSFdM1wA0fPzeDVPtgnCshGRXKgXxYiD
pCv+kM/2oX8AHHDGLaKBmKAlec2jHx5UetsXS1MBTB9ituei9BtYFKJByDy2e2af
lwizP947wJ/FAsUCCITOVNr+w4qiCamuL6xX/nxIfHdPsoaPRMNugUPUzJkusGbZ
yMYMPhruzWNTDdolo/ENAj6F0pC5NC4LUsl2WtmKKGN3JSx4nhgpKmqym+L1KTLP
fWrfbDgFjm0PjNhTXNW+8m+9XtK318pKyNxd/Id8ZmbBGUGoeg9u42ZGvIpdOJSg
6uYDcvkhtkjFk6opLE7yK4S2VDRsNioPnBJ1oXoMnW4+lMR6V6sfOQxb2H3gGPbI
qKgMlsezctFoSKAmohi6B6a0zXKjJX6aGbSsKhFnhpkhAYH1s+yscwKnS4ft6pkU
uc64QbLd8DHW5SVkR6fzIHtDJyhqra8i0T/dXkqlW5b0PiI3KsfdYtK6xY9jGINt
MKre/o5AGGIJdKJsv/ebTEfF0lxueafP3Y3nmbmo+yiLWg951d92g6+BiYlgM757
3/Ma/tu4+TWuv8+ahoHmuzEWuydGo56KXuc9P4jNCdOuVIPtZa48GPKAGBSTVO1f
02HRoSuJagfln54/l4QIC4kowkIvz6G0ARaMi0rhH2UPzuDunGpc6BaZIMcx02vt
cTT8paQhZN7lHYgvasiFThBkp72r5A/58lUq/oOf5bcKsRkGkQMag/G7gHZXqT7/
WDpTnCoe5bPx6wRJym5D+sZuzbqHLfVGW9qEFnqVcmvl2nxlmWakjx9b15QIcnIK
lHee1DEaNejHTPvI13/eJM48UVl+Q2MB2cmLhdm5J9siSKWXNer//JCag9R+eoaT
tZtqVsZCwniv3+9cjWg79LD5V6cnqWiU4FoSYnFpr8ONsTtrm4WyMEXHDEtmfjoF
tC5cE49mcjuHUYZvzJ91/qpHnVtXRthVdhfkX6nvZy9vuq74tOjc7yKXPZ5F/lWE
M6n1i1/4HYwpjGtTrj/OV9rHTm6J9GvWfI0bTz6KI/IYQJTSNXmDhsUJCeoX6XxW
W/03MUfskB8NTpmG3weNKgtG0kDJLq6fcNKlFh1X2u62N96Gzj4hseTnn3U5sq73
0VLPBTJae0Y2H0RB72VcuYw6dIzT2t9YemIDp+DVTfBNi+C+LMbssS5arWlyDZGl
4FaPyF7pjI0p2+Wm9rDF3WhLXjvi2BStHi8giIL+9ogKv1pxCbE0iPxWyXsLnfcR
T2Wr77NJqClGw00/Itr8NLtnEjZkTYU29lptgrQR7rOfjhuMTKNwJvxGr32WsBR9
tiYA5Z2IY/c+Lp5uRiq6EF+J6xpzdMAYKozZlsLKwGeqqWE1CnOxIBfgnybM9XHP
mV6CzKOhBQ8Pz7j8E8OENfMbXvQ2KsI4eiW3gR++zpZxjJoLXDU5fbr6tuoyKHBE
XXPDKm+lWaLcqwI2zkrPlymcnELLISAaw/Xq+nibmsIlgAHRlIuTGZqUTdrbSmAG
ATkfAIIfvthC5cfRMXQVEHpqXoOJpzx1HpUPmjn2eNhy1rvH2FOSy+gJCu9LxsES
qCxoC9XbgpeK8e4OPmbfp6xMVwuU/TF91FQ+Xc0/HXPdh2XwiqcKYZyKIcxzIEt5
xi5wL+ARSYuGNRSOUIW92uXmG39l+hujdZ/loS1bViZ9s7aCaWlVYO9MXj/c+LqN
Xmin3mQV39y9VuJuJFj1KCSYytLOkB17drHXpSHwN0kbIIIq+m5nKgSsqRNTkvPI
Qo/DRMpdK0z9comlw8fnvnC5bM3A9hpGnricXMvZLNZxMtBbD9QWSva6nlRqnw3S
TVM1lT1GLxgbowHO3WiqkD9zRLbCjp10MnupH9Jjo6hu6JHeknYe9axnqAwl2QaQ
9UEvPwQeQ0+1jVOZ+kKqWSMsSa2WiFsGDvr38ud/Y+YtncFt8P79txPESSUSUtGB
uUbeN5k2S4K64ZJsWu0lSh4rBoh1XCpffFOqzZlcdcwVeydidWPGB1SeKuniW6kf
XR3Bv99T4UuwKCdjkRdO5ocRri+tAlzDSaHV6p72kirser+LzABciX1v8+Aod13h
p/XxdKOswCBYO6zKhoKSZCnxWMqRaV0GI1+/XSrP3gGA6Zrd09DtOadwBqSsJvGe
XcufTY0CgqF7gpq3SoOHez6EKRF43cHecHURx8wuhBd10k9K7S6qLBA7Zt78iLPz
Vvd/Le/WN57PdLu79pun05yZjqisGpu5uq8VTSz1XIneKOMXGAWVmfdaPcGBCRwp
lxZ3dAVckUEPhYc5zRwUDMdInn2REXm66UIkXshgjPa2pQIwXvMSEOLhRWvKVYaa
FOrvV0jfDMOGkMXEXY2/WXNpU/RJMmQ1Z/XVKokgU6WXL69N5gVtua6hcdpMARbd
kjAK4s+5qdZIfk+0/QSlgkXnvBslNKgCppcthNAugETCzrw8zZKL2UtT4ODZEkWE
C9Zg+ktocRWYxdvJ7tPphOBFIIKQzSP+uejXt+u8tlOaWP5/RqE3oGf6LwXAXlPd
5OIiTn89b9xd6aCP/5EMjlyH2lia1L8zynK9b/z1XO6I7VI4Bf02EjSddrHQ0vm2
nFLhpdQzhMXVEX/NjffD50rVl5Ut/EbZb0Lh502+zO1+g3akLlCoCdY+PBUWTu3K
xrDpEOrFl5NJNnJvQZ4Rxjf4g0ZTZx/wPHB5GryPK+LbjZ4aLWC8N9syybi/GgWT
axOdxXjakB/Ta3HzgCuOgndz/FzPU6uW02mUd9vOckA0F6Dzu7i1mPCmmkYR7yeY
dndxKtWk+H8zOVSUiTluhVl33dyj9i6p3no8N1Y9I5hqEeZixhKRmcWlaPsd+X8B
mE4CChhuReMrI/V7+tCFvTBvqLDF8ceUGfaGjpnnlhA6DkVDzFZ7SzsufU57n7Zc
ZkOuafeNsqdrC+TKUwF6RBvBMJwG/aBQ8MSVlR6IfbBMh9IffrJCf1wrKFAhPhyL
v/6bbFMA1vtV+jOI4ueC207ZHHAger2qxOh7kgJx3frIrIVaB2rxbugNy3z1kAo8
PKMzhuZDrTIJzHWehzGz09TJ8BVGZuUyGKdP2wVMC2l8HQO8rys9/e/7eFNrqnmO
dV1upTODx2o+OEh0lhSEKJxB893unzC//NT3Q2cfg8bxVWIsUs97lywfYOfgDNI/
dJ0oJm7IY+1PUZexO1niE+n5wKEjq9PSjSokoBS2Uy5ENd1F7P6MPMEwZuH30Fi9
/sQ11yBHV+Mi2+T40Gp6RNPPWJRCcmeWole13xOZMGJqiWLxxCLMtUyE2kKvH7rX
Und8iwFa8j9fcMeEXeGxSRtk4OIYQdGzD3HsPJP61FL2lMoNaBYCmoGdMnAmzfBt
YUWuJJK1cAMVVpD/gR+2yS37pBh/UimSA3ymUk4t/hZaoBxOwKKkRtfEn2Vi30qd
1G9l+iHZB528RmrYc/bgEFz6FJYdzdGtH4bJJcxHjmkA9Le7JlwRBHi9Dt/I3bAe
ACSLA9QmlwNbid1PFA05lKaLauXpfGo/uYXx7yNGhQ1BJhjx+PXP6oEH9uEBoTr+
KZOKySoVgZeWyYdU40xQbMediExBrGkyPbjumuIBeGyX/e8ImLXD/qoNXY6BGXCi
p7XKNwnizWF4i9FYKWEX3QuBDpy5tCSKXqOzK+VcRPwy89zI3aw1AOT7oXyf/0gr
GSzZM4JzAq/B7k5ppx5W+uapRlbml+rlx5WTqUcT3bpVi2xv1Hy2EVIMRtYHr+Kq
+pMj+TuJxT6FOseLo2vXM4BW2xL4VdIpWSr/YaHc1lCDRZ6iy/7ltgXLR5s9OtLF
Ckj8E3E76eryxh/R/icwhIwt9mjK5OrbS7ENHsypoIhoM3Z2Yrw8NVmhAocN36Uu
LDDXlChFOC+irLrk61SGQAh6z2L7vMqnDX0zQkRfX15YH4OgrxdlpQsLK8hLtrIx
HjjgNjE1QLu+5RWV7IYOInEZPILabWyEVIxE+4Ni03O6FGW0NnT6p0rIAr1UZJx2
aRq0bwV3YD7P3GeRzTxzg0TUy0witUQfVxY07ihpX/zLLHJAE6koYkzkmKswJkWe
zMq1lWL+9IZvuRvcwzCyW53OUc/KqrWcNw+lTbm2JXjVVwacouC82GB0HxFbdaFd
rMV9iI6MzWpjh0qGxpxQj3QElT6eIUhvczjZmhuyiA7oC9uLepup39Uh5hed8aLe
6j4XEmSllID2UQwMIjwqO0ovgx/Fwpz4MbAwqCt9VpLeJrOMttfO7/tf8be6v1AB
YLCwRic/+xvh1PhgLWccm0XghGiEbzL3ef4rEoZAzdscjqOU2Svy1E27o/Uv15vl
qKL/sTJediLTwTps/AMNL+rgTl+Qp1dckhR+/+ildnpwnola4xmwiyzXEL/dVEpH
hcMRatX07ICjGn6139P1BJHbqvZtYgQFErJDPR2r6N/I5mIJYOHxZfpwOhNK78Ds
pQjsTXkHLJCMG2oXkTfpF97y9WwbS5wRzuEy6EwpIlV+yPBOCxonpYm91/C9MpFE
/JM+ZcsVw7PYzC089aq00zFyXpGk12PMcniiAF31f8wcRNO2bB939XORg2XMwdyK
iuQaaHvuIUCXqgIRNAzBMTsmgm8xNOUh+ic2Cyxs2RgvaL7QlrHRYUdQBWu2y56K
5oI0OMGU/aptuVVSzItfl71uByDBbNxg7w7Y4ues3XTBAIKwSyEFC6PYIkD8hwoH
FI6GpuYm4g1cXPgsvUK015gDL/NMw6iU718kgMnP+h3/hvSjYXqUrECHZNmklRwJ
k6E0w43vQWyqzcC/1cu+VW4It7X1YJrTadC+CLzNM44T9fMbJH4crnClG59Gtgri
N05UtgKZe5aigODokApQ16gSmsjuJgYP9p+UI/JxmH0g0wF+ZdeiYu2RMDJAL4Vv
d/czjvqaiG09WCnMca/q33SDQxiGFu9AINuK0iaT2L1gne2WStcVrhg08oK0AET6
fa1LGGXdnw7K3W9oI1IGun1KME9nfOEqTeMZjp5a2bnJpOWr3nCo1TnfzSGyvNB4
DhN/F4kI1FOFkNIGxOwLM/uuSenTOOA5n+tp+BL5rSbUOM5k47lgg9Nr5/JSJvPp
crZPQpDFF+8lZMAtwZRHFRYyINJduYTNq/2+VzaFvJ/mOat1HJLun7OcjZQVn9yc
nKm54HSSz7MqDCYWfwQOU/5kcrpk8nx7wXuOHIeZaN7ZMLp+RH0JiSEVUTmr+h+1
5o9Kv9iPgkt4yMezxqyFgef7ddq9DShRgvXX/ilGPEkm/ibsD03D8T7CBfAQxATi
M3lIeGwLprOfTPRU4vous8ESs1kHpG/zJXpBZlsFaJmc6F6a3tcOU+pH8pFLfzJv
loAYcHXzzi263XesI1GoDhGbvMaom2i1eMG9oRdGJvnbmqbpZi8XdbvG6wUKEcIg
rVzD/uyOH//p+Z94zLo4Ee3EQ/yH04pVuPFVFOQuZA3pO1fdfvAi5MABD3DOeijM
WQ4SSKUi6zvLSb8+wifrinfTcj6Qi/69A+KEHPE1Sf8EHaeCe+8f5DvlZON3GQKo
TOALtcX+dsnT8ltXnOSEFKgtnsLKH7kE/MMf9GGC10vEGBhk4JSTSuhL5R4YwJpQ
LhHeubTSdvWxBbkgXqZzzh4/gMgcs7WjpRmVfwDnC8a7fzdJ0FtHbxFwzATpMhXO
gpP5VGVO7RAxi9ezzkVW/aVaWNsh/2JvYCMxKH2x6ooLtGzwf2fZ9u4e1c69vutD
KbxwV6m7JV9V+a0lVB/e5vjMtsqNVURYy3v/p3bp6XZ596ikdoPnTMwVywpmhErc
MjWjdHQ78J30FAgaQJLObQaWNN3AGUpgin4d1jbs15uMYFbYDc+rxkstHsEitKg3
YNQNpgXhLFJGr+Xv1qM13+wm+10/lyUT2X52wj1aWZlzXILwKZFWgMBuaFXHBYPa
ZmLgR1qcXNuUKE8eh2DB94KAb5AyUqEn1IiplaTDoiXEJ4ApIaZkRAPWdnjQxNPb
bDWgXxJvuZnkC6AXdx829qnALk2W5a2jmc/Lm/+A3fxZIU/E4V1SB2hlrttv3m+C
nCbWwESlPKHVEZ9s8SXJO2X9AqVPrjxjT2nOE0Qxea9M/Z+1TUPOtsLQ0U2ZYwnV
q5jUQTpOOf6rKrbD7mDeKNPf3DyW1psmrGRyNdd5LJ90QDU1CeeE2VTfG9qFCKgy
j1iLZxfRDZmZbr3v/eT9Q8Rjjmsy7aV1pzVEHiK+Y8x4325Vpuiq/JaY/ZUjG9P0
YPYLz4PKQPL/FLO/5U8rC6/z74+OpujMC9s9RL9H3oCG0Iw3oMxLY3ucZFaylB7U
2aqicGdb69pTutXOHZ2HFVuuEHNgIE9s4j/HlQT7C7NbxU8bVqWwVFi58oN+jKiS
6pCYriPLHOVAbMpqGIAefVbutlRDauocu+KEpgLbSkkbOmO9qxbrzZgEQ77L3Nbi
mPwVjdqs/o4jQO9e57+bvq1dMy5/qzup5kcN6DyfQ/ssRUtLpv1dGx0zh/nBcxN7
DKWCJJT22K/keCAwsTXNxYMgY32DiZyTSj4OJUIr+8LWcQXPSMfoW8Ltu2NQLJT1
8W3Ck8nnVpOVIn0acu8n6MAhiA97GO2mWo2hQl04SqM3z4DbIKOzPF/AUXCiBlfw
8fzbk0Vi1A2e/Ja3wRBsEiCzLGKKzQBXNTSUnpsssrSTlwoblIoJ/fDmuTdfpJWB
4354IyTqZjqZqjxalWkO5Bzxj7pjgHwmnxHwJXb374/tEl0qjOsWupz/JnaLUPDo
LLOY+43OeaVdgQdRLImswPS4YW7qeOMW+6m8IyS1UbHn5e4ibMsBknuNPrzrGDH8
3atkpL3ZNpYXxhQs6GwX3MrAwVz1PgjM7rOFBBJ4LP0JnGr34pfI23wug/xd/wXM
Xynrb9GC9BvHI+eP1sm2KwX61wUHyReb1hp+Bl2jkjB7JbxRJYslqWCny0GeYPpY
/Pg0Bo3AY3iQv5tQ4MsCoBFISlJp1PoKZiOEcbcMFiiuq5nXBWVlANF3D16tZVAh
n13I4SgkuhxIGCvS9ByIoa4W8BrxtkYBURrnKOVyixLnOBKBFQDOJiZVOGjwvx81
OYvMrW07adr+132ioDL3kGjMPajnV2TgnA7jIbFlrE8ACoOUHTyp5WGdm4RWOFQa
VGLzTpaRsIwe3+nARRFET1vnNbcA73HXUcMSYnPSWlpiOt+G/c5YDYtB0S97pp/y
/HmrQyYA1/qteb5nF23/tEr9y1pCDDlU1EGlYf1B4fKLNTlCE/nrg7WNC7Qdf9hK
VQxivThUaEIIZmPFMO3PsVF1tgbE30q9joO38K6dkEipzD5LRZGOcHT6f+Y7pcFd
cb+6Ds7X+jaymeYF+ocR6I6gEUOHIFraWdhx5YPnpJNFriZ2DyKj8oxh4W641lsK
IHvoeRsFdVENKK7G5479fHrpK7q/sdqrLkhyb5MvRGNqPdzygcaUxSUaIHzlvnD0
0yFSWUKBnD8r5CbSYCAajIZxmj8NJwMinMh0Ss6w/jZTovnwbMm9RX20cV4lWGwo
c37OTBJbvqXizta7jLhT0YlydxaQe1Ou3TZCaJY71d7REjKfNJY8DCQuQJUeS0bG
wn5LHWoMM/UgzQFIdBpid23+fcSDKUBaUaxFkDXOFITUMxJo+EcXN5tCfdPZ3zd+
2DO3ktL4QQ1pTvQ87c2fm1s7sv44UcPoS4MZ1YzCrX5vRG1DjemGGO31+lfOKYzx
a9iia4vfzWsxxKmO8DwA7oeW0YxsJBNDQ2Y7wi8FjZs3igsNeFNT8ETwbqf00IB7
++zuaX8Q9knktQ7revGjtRKKFWhJhqi5jxCAP4Ta/jSPQpvRR9icyf5ken2kNHuy
8lymEel3I1c0LC5vmbrRFvVjh213bJAY8ghWIdvKi2r1aq5n7/qaFUbq9ZI5BzkZ
rVRbU8NQ+O90/71RyhKpdUIgy+QX1fLiGvEMnlfBls1QABF7kauo66iFIBk+tlBo
OuQxFvqfxdydfoInlr6WEGTMCWIt57MPWqt5+1Oz1AeYfI7d31RielpJHgxehEhp
02+XPRSqJ1iFHDz7+Bk1g5XqjrgLVBjqfJKSkQjpNWiCEz2xU1BthFF2S1C8SWxm
xSObKmnuvima6D1p4KSiBwkvwQOOhRt3SE3aiw9580Um3WS1nrMOV4H/y9qVEBcR
hVp0tJPXIr+YA8DBecaym7AXcqW+XWGNt/z9nTW2UCZR9CAotdeddUQNGHh3WOAx
uSCaZTFfqRZXfnyDou9+/FGy3693eC9yREUGpgP2d3hA1c2V2kuy4NtFIGTzhZq6
tL7K00ke3tgy+TsCsOUMwSLbuYhsXmfkntc2Rc0vM7425ebhK4T6IRH8/d2XvpYh
qMWolGZ7fduZgLC3ift4uUx0E+JmTmyZODfrsYCWtgh7DDKZ636WPfJLN76P90vw
bQRR78vMyv6jauJAhCiYL59sobJtTiukSZygDElpuq+1UETLv6IZcA9r+QXCLojN
+bKHPVCz0TfTxUBa8i2XcrtoZKV4keWB95UKPFI37QgqQnIFAO5N129CUQ3KUzkI
jz/VCWnHpmiJnfeVeX+yObvZcIoaano5kBy/QY9qZrHqlI7PWOyVrZMH880tGJIr
qfWsNr6kaJiGeWuL8hXKnbzoWnZ3ZHzyJz4WAcma0t/CFsO9qkLcX3SAMIzXHmOn
4fVYo3OXZTfNAjhm0Au2GO5vn9cM5cUQDhgnMW1UtUQLBsGv9zc5lFMOzzwq8bUh
pmSBWqNbND1tOxialGWPqPYQphWqJl3SSGAub+1x1vCx/UssjA8B3SkpDYeKyt8g
Z3V3EfP75bDtsVAmsOPH1Lti/V9VDKpVDbt37U5nHOxwzmAhtJbA4v5Zf2dZqbVQ
ZxvlwvveJv40tvrcNJLaEzSvPLDfD1oa6RC+eqAgf79Rn5wos7ZohrQfmWI32i4s
+Fetpr8HfPZlbgD/TxUHcOYT6M4gqgJXRGsS7NV1FMZnt6QQgdQeVZ8DH6tu1dTJ
xvsYiGwWis8HLVhXsHGf5AHnWBXZxwQ9Qz+J+6v/cT2YzgIHjqiXoV4QGLwmKJIw
2JvwJucq4l/usze7nG08vrWui70SyDjwyMOhBjC/YKD13W/DDCkqZzNV5v/wuE6e
+oqlzEVtMqkDpb+g02lKJZRVc4fiGDy0d1t/MFkqFoKZWCdHLKVHuORMn4AcoAoL
R01UUq0LQruIJ4wVrUYK/Vp9OAsxYQ9dr0fiBpZ9vvcB4Wvh/aGDd+QjB13M2Vtm
DVp79u5FHPB5ygFvXkK7RRZyGuvhyUEpFeKmSe6AVSiUERjLFWT/Yu/YRzorCtiK
s0Cc2xihKSKeU4FXQlzODPIes+vNCy7FSYYHPGmi9pl54axrF5KEu7HYNX/lOG8C
AITCuBMA6//0BVZiPvS6+3xrNXzIrqQkg6pp1cefDpet31hbvStJIi2olDhmdsJj
zN6ZKwcql0hXkEmrr4umvUY9NjKZDTB1+AFOTo56SVB1HdViYVGffTwABIRTgV48
9H4BNKcSltUe0McuxTfeyXm/dEDc0Rr1sdtQd18Gf6M+pZYtYjgBYVs300gUdEoe
/my56GESaxpluxzEyfc2QSyJMuWIGM6ty97g4vsxsbwzaCZS95udoS2DwQHY0fHH
FGve62IA2i6fPU1Zrg912+g8FnylJF645ucscKANMV7vSGXzZ22nUpHP5dD0hS5s
RSFgpvDpt0X8lSt6ljHiu5LUyhlC9bTHy2N/CZz0TdBGKAYARNBrn5901kq01PCU
W8CNRa3xUm6n84jPl23pKYwy6vSfokIO5S32idyakClMASKDwwpqmgsHyLC0pD9f
avb0kDN6USLg4Kx9SVW22uY8hKQB0KiQ39kEnr7FoU6XymaAtgkty/Wyl7MuLGVs
pnwEf1+Ug25JgzkY8B5764J7WE+CXiEhN03sDKAIQAxCj0tg8q6JuB2BIrS2l0RG
dggmVgK074soGYUA0Tbh1rU1PqBE43XCb5u06Tqpx8TcseMInSNvUGXcuoT+1F9p
Arcx2XbdAAR768uZre9Kd4YMSUDhJ9xElr+gwk15lVReAEXe9UD5be58ikZQqzw5
tpF6iNDBu5Vcl9ocjFG/lFjkFW321+VKYnjZU8DDs6XXTKRg0med/oFFJGxUxA/V
TvTGGSYBlVWAmG+QK6vdnGL2EnNoDVu141HzR5k+tpx4gEOlVGSVoqV4xOUgxPjH
zATmt/IfKnctvMSmORkSUcIYYjbislQSxE5GcRvgepoxuB1/d/WBHihW0kzaHDNU
je17xpDcjla4EdhfqTGwSQl4NI1lw0SNqsXKyBT6pO6qnflrh+Mf0E+nvUynziJG
i1ehzIgxV0Kbg20E5Gm7OPiM7Pg9T2+dN3Q21qo07HPizDfM9anLEZjAn79z7/Kr
3wljWwHhOgHqCWlfei6OYUS+F1TISyj3puQT+obYUJ5pj0gNB815oAHj24w9MY5v
RRKmrUGvPhs5KJ/GZjlRM8pHuO9a0uIOj0qgQmYXORgjU88c3w6YSrOoXesyLIWk
6AeG2XCpv+vv7vX8bvAK4D8u8RN3jjsRLzRo/o0jK1wF9t/0n9Co/J3Vm6+eIHUV
NC9xgdySp/a6Ij5PBOeTf+HoLQAbXa61ie7Vipm2udpv+PRwfQEOpqKv1NcNmdA0
O6+OsK9k8XIuTg54WDvNNBvf+ZuU96XtNDKqyhZ7hLCrjGXwmoPJLM9MoD4WkFwy
rMeNYVBKQP0S5A+AuZdGMhriUVZb1XkDUVDA4vvBRk2pcuiPFIQbXXXqHreHxIy1
TMGyeqFEGQ/IOqGc3tIxtEdsW9xJD53aCK1jRXtoKffcNQzgu0GgFNLO2/2DVnNA
n7E+jCRWr+xUYNvqh9oyQGsV/73MwFM66SbzprkH8yKhDKbSnf7CU5TKqpJFBmao
V0fw0F9uJxXMWIQsLB5s3M+57j6QaB267lWaDn0ZGfVJMNVRbATcV9ccRWFr0gPk
MXbIRactLyTsB88qWY8i+pdgaBsoE+B68F+OXOpBgYV9U1t2+ldF4ArUinAbqoVz
3V9NKg6fHKWa/aaRXiICApzm3A5AywFke+p6ZR5bNM+AXtnTobvGoCBatWfWC7cz
Iqh8GqvjsSNimDx8MTPwaVh7BULSqDGgm/9A+/fjsDVY6kIE3Q4jjs9kgSYiXRhb
28PTCPLCgRhXVhP6V17j69X+GxI8YPLE1z5ywNQ+5r5n/GrkrcgZT5FgB86B19ou
rGlmoRtTBepn28RjXmG/YO1ARzc7zBwcaZXMv3XMd9Xg0hz1Y/bM1kAUDedrRdpP
Ci7YYKIafpfZWD/m9zm+V6CE7ARP2IB9JWTq0kzibRn5X3zLcUWXjrHlSF5fNaV3
+dAF3jBVWsjPU/r1dZE68f4grCuHQtGOtfzVOmEVOW72tpEw0zKLCw7MiZ3TWEBb
OnlvAhaQSzpECgiYkhAgA4SvzehN5c+gvK+wP5lqccmLQoYfwGDxB/5U59vpgpOo
zVy2EsXGCNlRwlTMgzY30Ot7weXTMkWdC0wU4ZntfBLa4AVWF93oguUbo5iC97ij
EZ3AyabelVo1WP3D3Y77/kY2iHL2GntCAK6Ta0sP6EToNh7XSqzDTadoAWWfJLEY
x1PnXMBotB+lGeCP48AtMqePZ7kHvYQCMaW2ofyq14u81RihHfdJ5dstg47ji9rs
sF4bNDiVPMR9IwIg4TdjqrWJYBPz0U8pULmHh2MVUDqIMPrE9w1AE1eNPZab4aFc
mfJs21JOBPiZV/Yl5+S2xzvBErGpCYRkZDlJskHAE8EW2iokuaqAiNWnPCC70FH4
Clff98UJjsaoT06eg2VyHW/otpasjPxkMtC9gcS7IWhlPbqQDo0xNuSIUOyaLf6C
cp1SPBRF0uGgqod4zG38drdo176XMJit1AsznkeFCIViDAsY/ReHB15+NCtBsq8C
kVSItHS02tUP8sQmGyT/ZaOfmhdpHGqKr3LTm16KoTfJHg2og51D2MH/AzGu39cn
qkZwuVu0XlOfQdARyD6zhZQsrIljYzHbKhAFmiDhinmeQ5xd8aD+w/EPYnXDli96
vRdUS2HvAo8n7H5W8gsoSY8nspj0r/YBq8VQqQ1N4eF3+aNe879WT8AbKK4kZOTP
xQ3eAqqvDWn/8rHt+lcfBiIhSV6XjLOg923ui3XF5R0w0YjSsIkJ8dBoaU176Vfk
9HQTDLp1mk9WEjpVm0r9Ky9BSiE8aZRVEQ77O2jvxds5JikHpjzECC/kpxUrTjv2
SQylKDlT0HzmfcfRqOHp9UJbudxQOPaatJGaUf/Q3EeM2mK7kFUzOY1yk9fqoAIq
/OV7GexcCbSJw/qqjNqa6Kmqtnr6Ors2YGtpvrU4tLS4DDA9fVQh+09AnwLadCeX
bsCMPnBaqkWXOGvu1Lb9Qd0zYdYzucYfNvHUnySG/WFZKRUmrLS+Otg0b+7EvDxe
Gk5SqRY6A23430hPZ/oaIzZ/cYj8vrH/U+WOeTSLV1RbglDoSWdGyxADSVuqc56O
wQ1QSuSib/tCguF/06SpmFi8J/YdIpjxwYg6/hlwaUnDlIdgcav7xYdPZtBonEOd
m3CUdRNywqSgVhdOUCCrgV0Y3jIKGxL3T2E7aAzC5adBX79k7W1UvwB9o/SH8W7S
lo6pG1IoVMiy4FZh/gZIBoUBpvU3YNqKcYHSe0lKMOJVqQMW9vj72wOkIF1ZOieN
K62zJDxLmGBD56yjhoWG81WaNsYKtr0jeYFyZD4oZ0jrBYramtZyPiDk99h4wsy6
INmvrOqZQcMMRbDtawrhTkyTxmGzZtsMTTX2JXFCl2v6FQ1J+rB5D/oEAgsdbG6f
i8OiPIUBGBSD5jCNOA04fE2T8hIwbcok95Qd4liEX2N1RbwDEOx9aGNOH58oxMDj
nOX5kVXCDr7Shr5gqYHy+pZlah6hqRgbEleHykcj+vVFh0r9/qAUH2tbPOxduA0x
Cy/UlFHr2+B0yhWeh64oGpL4Oei1yCLbnuk5U2kcVaotP/h8x79fcl10ThKRnuNn
gazShb5B/A6BEC6wcLS67EhHvdhDNhhkjZ4APFPRCSC5+51/H23mGnSkSC1AbA+X
gVUVN+5DlEqXKTudiaN3bBkq7aO9+lBzFwAeo/tQp8nytKAewojYX0JuHiKFGB3N
Fa6s9NrReN69gnmv2TKT0MYyMImgUBdGvbncoOTqJDtN9GVpV/oSGuJF5Y0DuGWK
ENLsAvea1TyeZOvbHXhH/VhFmtGjlcS7Bly1Q25ZK17Nu2pbWmERUTmQfwcJQeii
eyK5xm/7q9TGXAnARcTuvN68yn0Tdljoi3C4I1CeCTDsmnSThMQ7igQGrd031G1N
qGEqCaOuyeKv1MPIAhREZqxBZHO5suOez35w8m9mIUS2amXH4ejT3EftYlYs/LKI
czSw6scQHSma4WO/TI+tkqvfRGZhKoI71InJd9+AFpVaTmI4c8afkW/nNIa9okh9
q8tEHysCJUzKTk+ljajD46G858gymdp8Rh0UIuYORV1xuVt6FQBKacdM8tia/Jct
SgNp2bmCeIN04uqXAiQMoIShMzPnjVVDo2FudmAM8ux9WCAMPJc/484LK3boYYZd
g+QkalsoAVRnhbeaRH9duN1rYhrBGNXS2Qq6ifdGoDPqCr68A19oGQ61M1FuIdTs
Fh14sSREufvyZpowXbO7N/Hj4lXWholZYYZteJkognSjMWptEMCESCHkIc3yKlxs
6iDMXJThTxRWQm8N0+lprYagkAIfca7nBNQrJP6Lz+zzmqQGRlIUkyNr2VBOX1L0
0G7ZUumIc7dzEGONK8Epl2kpj4lDvrx/khlTXdC9xlhi5AM9pzZD/6+qROxdBnvf
TTzcB2xijySx+ANNnPADJuUCicInKzqtNsvGTp4Y3cb+5VAdGQ8gxxEED5qwHHdY
aJR3yM7OwyKa7hwn8d8P/Ob3apepkEB4PAnzIoQoyM1U1xEgYD+DeJZ4wPHMq34h
t7EpeQd8OzqEKcppTkWmIG4Q4VexTDHfTEWrKaPhPeEJyfEcbBxSFGq4XlVXnKj7
k2Ih2BLBfw3fIpMFCT4LhHGGcDaNOb1MIIIqvhZ0Di/7f6UYraqWEGcMTfqID3WW
osnOHF9ftG5vaaF3TdZgrkLRqrYxECfAD0LxjEA4vBYfHiuVXz82EoD9JWl1bbAf
ePSSNvi+Vk6bMM0sY8ZhELSMArxnnH68EemQdhhsgt4CT91lv+f6vfPhSH2sO9nP
7J/tHgCe30cu/nGyqsP98oxtjTsBspljzRzZbGhnwaWVLY4SlcRyilRRaaXhsHJS
x5TQ2/SBSDI6K4nzRJUfCEbhF85mRtB50RU3xgqHum3VAvhjBtt72zN7EesszuFi
NJM2mJYkIqSagIzlUkyLZV2ftw31XL/Zem3Bf09oKJyTv9+zlnMVAPYzRVemSNNn
oBnhDiDSehh582D5GvIq5Vte01VH98ikTTSKhMhQy0/V+1WtRYznU17xLNL791d/
P1fS5diOW6EVTS98A6aK6d4ToKel+CIP4Sw+75RXEgqNUBpGVkPQONsBcYVvBiMm
egYurmktgExak20o+UvtHYfH7ozjU5yftqPr1cxxcKpS1kRc/lABxh3K8m33+uhT
ntH4DgSVJiY2FrmTZ1Ix96m+nAFgXWt2+rQ6Oa47f7/euwfh+wW53rkMwfwPfAZx
QAb/CQxTEuuL0ZM+mFi/Hrm/TOZBTeSxY5vjzJb6OYzPvqF0nNsalLs63w3+h0G5
A8e28iuryUjQY44YillCfRoNzDkTgNby4lbtgJKd2Hlli/pp8dh6nnaps5b6by0d
ZDD8Do+85jBXqWUEplxU4l7MKDR6b2eFhyiExwnkQtqKJ+/utLsW1q49QBuStQG9
9jjqD55owgdtJSwh7FC0+Qm63uAadr2TSkx4SKK38zDqBjeAzspwVVNkaIRcgut0
MnQg6siBY0ugU4bZZiFXCi2xtJEV6raiOQdkFEeiEh08SB6QGlC9FeZrS4aZK8aU
hHIVONdBi1qxMcsSCIHkMaw3seAU02AX8hfDub7zcqSyjytPuu2F/FG+gkfze40Z
P1kyXeZOLopuQ6W6cr2iEZK5sWn2vGlUeTKlX35/clVOt8HGWAyDXFNuIQ49RMsx
3T2gUZXi1GvfNxhVRZxXYCEYmSrXz68HAf1umSPe0SwikyF2SUJVuMRdnPn/nuqf
g57JywrEubHKDoU6DW24Q62U9kxu0u+47KrvnUmQYe4LwY4yEiGteUD0K9xOwa4+
OhZwIiHIVSe0WiZK0vhJZi8xrg8noj9KGKq+zAXyNljxNMYcwZ6qFXeWrZT9ToYC
XXSKvqux8Oz6SKrHDtQ3h+1cborpbR1qxieBh242brYJzZRHv+Zg2/IqYu8dlGRS
kZUDHoEDZF9DsoJvQHFPDySrxFYrQw61hlp/JZHSL+4HuXofJt5bzsreXpkCc65Y
oycYkvMMSu9h1G/twtO1JLd0SeB/KJGJetf6nbsi/aApZ8LIw9D08Yda+TZ+FtOg
De8sRjOOoM0ag+AVAs2e3A687azRfLm5cWsfpwUewhoSr37ZscDOWmWg+LCISYuZ
tUvvgU8UkKIvUW1uMfcxi64qkRPMtZ/82w5WrBzlBbNM+XieSs75NR5VpILHIvGY
vvYgaD/6tMDWMXnXkaE/1T2W4iW4FGpygDt0fHJE5+gaZb06u5yRZC5uzMAyH6TF
PeazWrlWv9tLpEFFBn8ZgqViT8aJl57ZT2St/C02Ol8woaCivPQk0UM+DYVwkw7v
YniJEERYkNM+x8gjWCv63utZzIlKz7g8b0kTbvcU+SdrcbLQ/6pprKcd72MXXDKS
0cothXEzDoBOygqxOC+8ptOKzBKTgAOUOV9Xf80xVZ8D3sRjFon5xShxtiWtMzSz
0wFx+IQuvOISCOp9EjQzR6UbDpygfE7BGKxfBBNevfLW0KLV8QbJWhn2xaJWf+JE
x89A7qIpqZBllMR0Xt55IPRzcZL5gG4ESfqlRkDXuN1TSgnCeQAR48RyeXF8F2Le
4kdM/Aaj5GYoFqFXs2vOaCfkOeNDYFDQE0NDOJPhCVIMbzjT/dHXZCam73fqhsSY
J+AiXy/9bU2uBAaD/2sI/KyIAe+3PD173tva8oHNrREmy4GpUWXP7TStiKu56suO
a81EaZdd7JNZhlODIUjC2Sep9VbtwNYXHS097DWIDk602YRTjVuIaJDKlIeC53vb
K0xVX3MsNX+i/jQZA+Ie3zmOp2RvfFUUNEZ7303okMwhdHc3Cx1DTnauBLg+9gcX
dxOcoKRkPxvcuDHTAr90iBo9uPwKcnXIkdOAzWkSVvb2VTG+4i4NcfNJEatRMm/7
rZmRy8b098QQPoJBb7SubuAP1LJ5p2yio1FmAJvmGqqBJVfUI1uP6V2Ozds+IOeX
eNdnvnZ7pZg1VsNRqBl8Xa3w3LNOdrXTvuvy1nB1UiJ9jR/MQl1eYXo+crRsLj21
heSjJONV1DjIwZnHTDVvX32khYVL2QysvPdQvqoshx8hqzz9Sst0BJxJfmxeRgV6
810XFhgRrAjgyxXvXUpqMXIU5WBaDYFRMYypEU7qEeB4B900lUjZc/Y0QfDEIu/p
8O7XCR1i2DdcIPUoKyaUHjGl23fcQ2cr/gYWIybXXMuah9BDuXL+Cx0oresXTmZv
Ak6q+iyH3WOJ8P18BWXQGIPCrzoDyR7t/GEcaafHqngWHA+gBxHHDDbBGOmRsfG/
WLoYROvE5tcj2GiIEnNmSwb990u5jShfLawUXywtjLiD723XH/OY1xLjkvcNF4FP
VX/kIIXb7QJ4CMNpxl3Jp0eRpnXiMv4UwCtIDFP7fR8wTUzs0xK9r/Z91YCGVye/
1ZuOXU/48rubVKKn1DJJq0Usu/0vspbCkZhC0fR93W4h5arCwySEpIsxO4PfSK7b
kStfkH+3Fbt+mJ3Q5gTe9/cH8FNEXaQ4AAc/TRtxEnMXBGQO0cxVbX+cuvmxLN7i
DEVAcBru4FN/GWbgNGkqndaQYK9IMNpEMvNwCgIzaO7LWSt8z4YBE/bhKCqSzyc6
uk2+KQzK5W57/eI49Z0xLF1OSBNv0/b9Od50HUjHngDKJ29ikR/H6jC5IQEs822T
HdyN8ONdqdxStUiu5dJ89nAXNkyixEpXqSDQRAUi8VgfI6d60YllVQANyigdv6q/
uC/5B2CNIhQRjC97r8hdK3e1KB9A7Hp52Im7PbgxTJO/sdXddfc/c4kEcDJqg03i
dopYPRH85s5wWW386mUwsJJcqSF1hF15QmRUUnED2uQ0ufSTepfvDJMTD0vBZgJB
JN/IbzQNdQgQurd4kwQW6rTc0eTFdzdiM9cotiLUyeBTYmh0w9QhZV7KYbV+UlC5
hrSz3/FWhS3QUJmmVtfbgvopf6wUZZHSQbmOm+WPez5rYEg9hpcXF2aGSpf4OMQR
+/xYZbdw+sPXGIu0vwIp+XDo8KjPZc4LhlryiqaUpyqoNrVbB6TNV5PhLgr/Y2nR
ZprV02ZDs4YN2WG8cUxCDCyh2I66G1QC3gYe0+nl2XH+HEiGvxVMhA9T4djSWUoC
6dBw+/zf97fzXumi431nnHIY4YNXilTJrAYfYhg+h92k4GYlJqvGaNTrBZrTjFV/
Rz3Qklh1JhCZfx1U99nn6/BvePaAIO3bWA4bEHhadhpctbUHeM2i45redeFE9Z5p
dUozuEYS6qjid8aqQ4dymnrqt+Ur6ZCR+0TyNsZot+CLt7GoF23+TWmjP6eA6Jqe
jXMe7pn4YJetFbyVWvNyklOwOGGWd8izcrVtoI/8WXX+i0vAMG5Yp3EkTu4PCr30
oDiUi8ypLZZfZclMs+LuZL73OIpLnjEXn+kjtK/HtUSrX8EKWMoRfdeeqbVqMij4
fw37kj7pE1iitp6SYYVgI88pc/oIlfaJN83RcgbPLRQ9gUoV6/kNI3QckwK2V4l1
lDfBa01lDv5cPZj3rzfp7M1WxaZ6W990aCUWgiFcnE+396i3MGrBEwK74K+M9IX+
XNeu9fjbhI9Z8CiL+gfUr8TfxxG4f0MpIZLhJoAorDAV+6pB6ghFa5D77xHvAw/t
CRJPnokpsMMru/B/ME+7Hbmq7UT5OFuxBz6RNrTIqhJ0C8X2c9IEtTZVdNZX2o0e
r4cfgeV2KdgvUN6tWHZu7xN4+oa0+kpbT4VV57T3nu7MD28cj5VZWIrAgbfQGgKF
lf/FsTzc67KPBaCJ9ayzmrmVJDLRX7eAgewL4XRw4V9NaAVbUbiIDWLRKx12jPj2
4H8pJ3IUcW/GQb1i4A344G5+vYMZc1zegnZAtjJKKi9S54jMaqf0Ym9VviQxf+iv
Iu15sj8S0mgFklC7upHDMnJAOmY+UjU7D/1NK4NFRb1hUbzTfrJBI8phF6cATXjv
VDlhr3N///IlWHQFi1q5WCsZVnNU3/WHB3Nj+Jqo0MJoH2+T22SMlHRbKo3uN6aF
kQJ1UVS6Cv8sLkWaYrzRfyQ3LjK97X35nxNpkOxNKLJ9e2erWezrmhcel8y4C353
DrDlGpMFOQRMGSjbpcbGBdIScWzCMK/Vtz6bb9QLQ1DHcU9918Zi5gCIogooVVQu
sPuVz0C/XnvEe4+Mh9/EhHfk55+k8ND1aJ29nAgzRaDfn5WTJwhMjj6yDYfRFm7Z
tglGmwlPYnJoCbS26k5xNsb+FEPDlJ8f6RT3zKJzXYLns2tm8MEwy2bWIR3nyi/u
h/1hwdnfavdacgFT1+Rc+F/vl6/bS9/IZpdTUNO20hgKcUW2QzIq05mbAEeQKaM+
WZ46Ukoxpqd55cimFtMQtPCi3zpn9FyURN9NYnBiyuhhmkdOyEhzrHS5q/Yl51BF
YujxHxZOnAemEPsrpkdDjI/Lj3P6GqYW97w9Dl754VfQbFPVLtsLvd8udoARZARX
QTV212nV51u3PTN3stQ+Sru7xiPylJthjuysks4H3vkXCDmilAo+bJqalW/ssyoF
Mroa1nqeykgw2L7V491Wm8omP1JTe7e689+sApg+BskTi1Gu8YXn3RiXKVvFLUTH
rQ+ezJR3sHnj1PnXGwmSWbfx7EuCQBMVynY/1j4naDpEyzCdpEjjbzCvdUnKxG8C
1o8AL1yUjSq0edPK1yqdGsWJ9WgvIxdhWfc8Cs6ru78YZi+xY78E5GE0BVuOoHNR
Ic6EQ1E8EQDRUknq3fqDYFSDIwNhEld6UWDolVppFMYiWd03Xh3rvU7JR+yfkNjB
45o8yzZ5JmN5uuGx2luCsi1/4cgs/r691RqmLGeE/vTyg+5Kbl63e9u58xTgb3AU
KzsjmpXYcdokybzL1EEhEqZ/eOTYBLhoy+AFps3e0bqucbYi25FVvrlNX+VLfz1N
CVNPIOuJXXAMHTXEctjqdHYpLTpt1nwIn3LYopIPvwFNfxp6b05Kc49rE4pm5raK
77T7pF34pgiDvOU1d96vaqM5GBev2MOe2YVucU7jyCJzEttXYxnWXgiuBVBe4Qp/
DeZ4Q/FUcKOF11wyZWhJjX730/y50/XggiOIRslt4qGWkq41i7ru2GAb11zShAAk
wYJEefG+kqTlDjcIkhmn2SBZvKArqjMHdYMHyFscYcuNnkDetu7G/HBs89Okdt9p
PKBdmsgfS961Y6VENPjZgaoVn4f+oxbqVGSnO4gaFU2I/SXkcm4X79Ue0tzGB4hI
s5EdW7scA+I+x5l9d/yuBNnPumbwC27e2Z0cwQGT+JruGje8SrgC0UCjzfQMew3S
CRV7fl5h+3raLVQkqDe1+m6dwj1869cv12PdCba6jiRO8UmlAyVBdyDXQiU7CjG0
vpm9CavkDrnVBgdPzG4ADhVz52PoosZTzUUPimbU8qEnxTx0FaRZZZlqMXgM6Cju
e8+6bRL3VHdki1q0rgmpSAeBcvEbuS0yA4Q8pJVtmnE84HvrprwIp5aBxI8NJX/w
CescMrNCreV+5zbl17i0/DTw+BS1soG12FQMGuvoyd/GZiUzlnT9eVrNKnFDTJGc
aqrY3/X0jquf+zJNZLgcLhAf5xHLQdgZTAKW+4UNCOCxQIGPGVCjSdt4S/oHO2+g
8DtsK3Gw8OwJyE6Xxeh6439hwLpT7qniEFXYTmvHe4TdLS91T8YQ5z6nlr9quyD/
Nk4pbxfe9yqkGbut3iB2YeEA9dOwolPgiIcqw7M9/aiD3YHL5/bXKknbggSJivGm
o1lOkITw6sqqyEdXoJTMoaURVDobyHai+KFzagxI6XZgnnCtOvjAhVgOZfQk9e4P
Mk44usVpsKmpLtYa4GO4s8T/Ain/D/yT0Mxxfyf5NN1Vyur1eo7yvdK8MUeIuNPx
AMQ2Gq59m+R3ALn+y9jkjOJRPgRJhKy1UldQL3LLbztiJxr+tRXQ6/78JIcAzuPZ
Dva0+KNcD8FuZkmrbNqjTByCnbi4g8A1ulCaDdBemK78QGaHJtIJnMQHRor0cXLL
Ph1Xfwm1oTYHHVJHdeZ48lz7FClfjZTxSbfaSpSpUqxs29fnSVjmshvdOM0KTpK3
hq6dsezi2fYEm1rcAEAp1gz45o/h9IcKuDpnZw/CFng+54UT5iaeEvHIPxLc6aKx
EgrA9Guaau+jDySmvkOnz7Iv+R4M8+u8URHfyGHZZ7mnMrOJdv4qfW/Wqy1ThOIA
agObWeZepXhtvklg4D0nVaMmyNErkBTdYxc309hTB8lZeEGHYBHrK9uRMNPOOxGa
af7SbNOD1SmUfGkNxa5bPYWo9+y/wKXgfEV9F3MqlU6VisApXLLByrkWTCuSllO3
1uN2JJlsphmweR9Ee9C7uvhDMZ8AHnKBzafAVmYMSLjR8xsRP9bbxHreZGyxm173
/rdorFi9+0o/yX7j9liuDOA2VTollXtLann9l4uaJkA1G5SUgyljTaYjgGbWZG8t
ckbT+BF4Zr04GrDCPHLW7RgeYkVamsf9/y5PGbQEtBUJYXNnBuSw5iMGf4Ly/faC
7/CFgwUj6FfEBjHXPsvIQvaYQ5QAEnATS7rq0Vc4NSyA74wUWZ4EgOM+w4MtIc65
8FXuv4Cd5qY+3VUQRJOcm6ve7E/0GfI1iHhD8UjrdgJ892kFbWVmibwGX5QXNSu1
g6vzdLrUVgqWcUaTzDOFd9MIcdv2oaxLB7XXjxwK1x7X3srD987R6wKHVkjyoMgl
DQBXjSxGDMB4HaaYQVmSQbxyBaqCyn1/bOIyBd1uZ4040uyVed7LcW9gghUKU+MI
wouqNwznAyXR/5ZeNknKiOvUWvWvvr616GjmoyZpwZwNI9YSKlG91JMsAiDfCav3
HTRCyULZKogJbUVWQYWuAeJ4D/gob7tNbu9pU/tHiYpCOmjd5Ke5GROKBnI/pg/S
EQgpZTtFdJamnnCgh6HiopdNCyzBgbBryGE/+wIK2QqvVbVAN5IOvuKEKuzmFGLW
6nuqvK+ljfjZk7wBwRllJfn7NYzwir9CPlRVnu2nG89hCKj0wTYIa84mtJu8diaO
vXHl8D3P4rtu1aG0boyJbvflePgcxE67tZmZ4i1Lf8YHhy4978wbLi5t9St9nsSz
q0B1IEEAM+d0jCNuGzNmhjQEQnp52EHYJXQsZVhbpLb/eO4T0YCHDB79TaUIIKYu
f0F0s4aFTD3c4/2FnP8nzbPGsuODPMra+EfUqMKNxbYJhykgFiIVkr3WcvaFlcsU
ilCwOe6IlqTBW3F61kmDsz74ub8GUMB5weXD6DuToODawKxGSD1Jnnw8qmTDwQAS
iQUR8qN1CDY1htzTYssfE+bH/t53PokbxNcwOH8ADJ2WPPdilz22HRJPfQ/6V4RO
g4rC9tIXA39FURm19u7peQvrxKUZhOH8dyEjeN6V5jmoYowDZTVn/tKGGzVxm5wh
P/q/LyFD+OSWTYlJm1TzB4JBZneXP1J//dWUdzRu22Hf4FlbRui9W/Q1MK6old7t
T2I/lO4dJRPg2I3jQNjVPxE603mOliVEgr2fpoOgEV3hEeHKCtlQbCcNNuLP3Wiw
SfrroVRYIbZ7Xkx3IrKkqkIgpMLS0H8RJHXqqD6gn/pi8GfyICCpEOBoUc7ds/b6
O/LNecb05jNhF8WFiqBwRjVACmu4yOayGyXzFBCFsR10ZC9YBvCK7iuGgvTB0g2T
HFyIT0zgWcJk7o3XGD63ZAO0C6tkZARDc0r4F6WyrJR7RnYwLfQIAoECZlzPMj8d
PjYc7LsXQZKEbcclBHVxhDKrLXL3l6yETkgqSyJ7Y0RQ58PK3+Mje2UF4nJM3U5Z
+9aNy2iKxu5SSc1fDyIuwigbJwSZd9B2MhQzRsClLC8TEimLsU/Zmi+cAxdHYxlI
CbF7D95v6ZtXJw497OsteUSDBfclg4hs4N6yKRhJaUgRN3GEv3Y7zgJQpZ8hzojE
DjV/xe9HvQjvOTLZJkt6djleo7GseGn5rB+YFhg4e1u8QjWz6ZfSAw0tzx3v6kfm
tM77fLOkS5FZJ6hMOl2W36rtrYUJjd+lUOOMWd3OVI2l0wVd1aQlq2RUGC+pFQiu
FkwXDQ4Q9mS373bAKHOzfwD1dL7muntftCAff/g7KQzCNaFB+dgj6p2uYRzAN2Ju
BBk+sf+oV9Y8CxejhGcepnT8f5PQpswBHG1LZ7gIDFImDTdoRyjI2JmwWg5itxhn
qmGdtEK66DyoBzuoDM3C/8OIOnCn4wpiAcFzYp6DJuECnotFkhg9SZ9WTFwblcdY
VWJ0XebUghT3RWCSmc+kpbAzdWSUANMAPv0DqfDkOMc9JPprf1wIxgCIomUgrzum
YMizplnUrW3LiYzJlwmx5PXur9FmbMOOg4DAvLNT8srFDl187UBMuO9UJA5oxJf2
wOZsvG2zK8DJcA1/A5PAFJ3z/QgV3MUfYqZiPTBvD71oqxs4smKa7RbrUKSifOgk
VH1nWWCX3FONPRurt0Q6NowjLpsTE8SPbP4/Xi73wDn8xCDUUXp8UosA0lqdTIK1
1xDEZu+VE4Ld/DDgPrmVDfeWrKZicv/3uoKoujjShEgh5rsb6Mn+Pi6RzvaI1AeH
TxyJ2wmt5L2oJ7VGLYCZLFYxYvmZTahkcuqz1qVgD4qNjhp31UDcw6AincRSmHr9
/I3APTH2RikqykHO522fIk15MhuGFDgiKE+fnRouhLlQ5c5XWckgbbb1Bc/ZcrtJ
Kmsp1T/kHiJ9zhhfSGpRWr3FmnLeep/bPAzO8BjiWQonej8xTU7WTSFNaP0dE/U6
wfUWps7rjwJZm7cGhO/wqoSeXjiv5e8PSC93VDRK7jhouALVYwHpos2Nj80wLgv4
Ajt7HIMJYZhx00LYiclGVtPl3Ovg1UYMG8JZZXZlq+f/4wa0phg+CLvk5iBEBCC3
OLl2UwJoUSmMgurpAV5D7Wy0xBwefyfZyUJOID1LUSQIqGaep/jGzKT0G50G1c5Q
hFBpwvjcKPRPv+NpnK2dyc33YQuiPLNTRh7T+ptNiVU9E8uGTuNw7llDPVvvozyI
lc+ReuFaxSUok6Hu1w0qWMmllaMpi6PZnLof5ML0N0GFUtpkZYh8vkPnqpWeRz9n
R4H1YTrc9GWxUbYdRS6OEdiEMdHLZeJ9sGHTDPWV8bKVy2VMB59dUCXFgSlFbyEu
z8JM06rGBcZBiSepKGkzRrr5sQtRMwqWCcFv60F8ZusTlmtc7i0UMP3PQ7ghAxUo
ltSDGxs1Z9F96rZ1WOntqMAEqHAaWJaUjNQm+QGFFSFhR4vmJHqGoe6U4BiZh0rt
q6y66XbYYH2TH0LQcrV1DFFBU1kxFo6eX3WSnjR+gGCyWFkL05w0ecM6dO7iAFql
DgR4KoFvA+qxHd64bySeKXAASQJyTO14ej0FaS4bpvcBaE9r7LhqET2iqE3OPkFo
104r4w00+cv+ypfg2TLoypowDdJjw/XTVmD0wDYH4yFysuY1OgLpsDp2L19DTCwf
XucT22MDPyC4gxD8v114laAL8KMdf52GwZ169xfbvbA8iZACniqZBPCP/yaoI9+U
n+pM3d7emyxCR5EWzBYicbqEp101eEHfwR3CfJeKOBZGMoQyXntCZVYq4zfJBr/D
ylm3x+9xz6Zs3vAeMX5ux5H1VWA92e/KRkh9KO4ehK9pIVpLkgOPDcfeXR2Z3WKF
ejzN1CazqRTbawisGLvtC85APsN8bIQ2NB7DlNgnfcX6yPiittK4nzfPb0c3tBGz
MiexQV/OHAcx2bGzZnDybCYQlI4rNqmIpEpOmuLW5sT2ImTmdPOVFr/IhUcn2SV5
ynGRnkomw6JN2DZZgBoe462T/SBhEGWkWtf2+7NaiMMurWGlMHekZvtczucXIvfu
PiivBg48KB02BhqqJ3nUyhkJfYWOge61x29FAPA6+FiKYcKLG42ufdl0SgfQfVHf
jpRnLMFSaZMMYsfQQoiiSiDjA4oYPfHtVBwlhTRIm6cjb9ludeqNR0vPkdOnAcnX
TS32LYemNNb2YJW9gwaVFShSRaH6bWRCXpKeZo8PTlNwcaTqWRqvKBHIQeCLv3XF
tn6yTzkpJWIi/O6vGumoeFbqLrat/00HlEjGMMwxvVdzYYImDbjeCaDpa9MwS21V
uz5X2/4fxwZbw0dXvyh4PfK/VPsNttPhgDlLiWyCxCBCy2Uhx3EdZgWd68s+UP/Q
Jsq24sUL2hZgiwqvdqAlUMjfsCR8S/1c1G7tUrtfwN4WOgXann0vH41SeM16v0H3
PFFYMa4sfbIxVaRTLQnDZKkEwPMud/d0CF04MmJPiTNjkPyvUMSRHf5VxeYGm/ZB
K1JQwKKPtL8xQnsVGzj9LLlKswkGrko6XDiAcTMWmLJjw/WTfme+/5kTOR0xZxDX
mAm89nScpBUHeU3pQBkR6XhHmQ/hJe5Eh7swDVx8kRKRQ69EGutKZeL4TR38z84/
c5kzq0NyL3gReIcILeiB+Mc5VHieSEOzhagDG00VmK+MwOj1gliG1qwrxZO23DSy
N94xO9psr86fjGCtLPaTkIIIjvWHbmsPOuT6fKKSzjvRzDjuDnTOTcjD50sSwgFf
yePLF4NF2UgEiAlAoer1LRoaIF5cUyC7e0M4+qNSYZ6ANutWDT3AJqfjlAujiVvO
+LK9jPBaaxJTwmo8+qxhy7A22Wga19yaBtToFtdCVcpyPofZJYim11UmxgIhXfVn
/gzhU6qH0i6ep2q3J5D6MIEJTEou7zBaqngtyJ8bYojUK7MTlpV4l6PPCv+ByToL
UYQIJFNWrys+oVAQvlHteuF88b2eX/5ybGZQC1Xbf9ryGy9alU/rB8RnLGIZCmAr
cUPjHhamRArreud9WWF34yNsWoMfT9r9kg8LeSZPfv2iOgNcznDNqJ8g3O0us/0G
8TlBoCpGm6WLp6nxA+jNeTvdXZFP4PmcRoUJEtz0hY6Vn/P+Fh/jynAn+67mXlBz
JW7U4SqFP4CIRrIlysjODgLHpWrPHOSPfEXJ1iZ/rWT4b8amBnBSyUabSQthOjco
JB7+0awQoGEWrYNoBwzWwoXdyufT8aTU6k6LZPLkthVk5DFZxUjmVZd2Ss7TPDzc
owVryu4i1AnIwxiP9Fmbl6Zf6JtVe+2Onv88wDDX5ApNH9buESTKjqn4wJiz8jf1
htzEIIGJ5n6pCpdzLL8+nE/6+eyb/HULos6At7N9iZPv9Zmk6h5ZycsTVOMSQBdO
8Z2wzI3XkTLG6zcr+DOsEXwRVYqCaJw4S47ldIqdVYIDuU31bo52scaWraeBroiV
Kpi65cqz2AsF/SSzY45WQELdBbz7EYM1plZAv42PHq8k1TI+D25c/I1XBQJqGnkO
WfTz68YJPFi79FJNtqpthfIm11zWYOZG/E6+LVGe4gLqRF/tQhfjdHv4ygNmxwBf
5FeakLIqt2SBIS95duxoXd7zk3NOa0Ju1UVuCeFv9N0NONwISjti++5yDY1e4JIn
C4GMxraINPwOoVUT2wcYHjREXlD8x+IoGF99RG4vkxEO28AuRxf4KFjMFK3N8iep
8do+2M04MB1hvMuz6tmgmWIYGbFKDYDaP7yqjCPROuDWtXJ6vrdI8t/YGFhDyONU
BtdMghbOP1XW5Ofle24t7cXr0GKzLvHdHOFMqFae/kMNXN6SprNT7SysHW868FBt
t+ObYjRQSXndpJkIjBViYs4LsWlEBhqMy6RrfEsCyPxdOBkMtcvOXHVcIV8JWU9h
fSRyBaOrYnLXjRv14TzKkcYK0HeC4fzt3ERIe+PTd7a5JwwIGWrH9X7Bme3toicK
AaPvVypJd5ZNV1/pCacItqlitpBmk1GNw+zeWZtt+nbgbqBsueeLmo1JLYXaUQTV
twaY4ykjIDcwD2e2NFfPfumAzDBuu3rU1WIjdXgPLT+qhGhh88vcyA2oofID0Ol9
31t4ZSQE5z5+9jagGxhafgmO0Ik7pw+5FOToAMQZGNH/Om7p8RjAIb3MNkiV+s6T
vnE7mGUeqEu1XyNmNLFx+bEVEy0GIfJH2bLyaLjDU9a/2EhHxPs9+W1LCKgZ0nUk
XoNAyIZadiMc5CrqkGQaM3Ea43RkOs/xmmgjcHSPoqlhQ1Q8UO2q50fHCZt43xBn
9PKIts6ndN+mNr69hyrg4IcVM8P0D3fCsCcgHtto6WfQq3/k3K0D6Xtyy4HcIk02
6urA1f7+f4dhhgROXekbsnhz0PvhHtYDoniSHfxDeygrMkUFCL9Z+uJJ4kRC5Me5
8PTf4HdA3PKImcLTwn4pNQRb1SobQMeDy3Xo1vV8gVC2pbYyZCZOaq/75p0vNsDW
AKZ20FxF4TQdHklLUvdQHcHJn9uR83nOrab4Oa4kpfwC949lLGOO3OgWsRas+RFw
Sz12bcA6Q4gTQsLiTwTSt42ZXuDzNVG8C86p008LJgZCU3fq/vjPCMiFPRXh74gZ
foqv8o8Bq5iRI3hfqt1/aiPAbdSKgCBh2lseBTuMw1Pr7JFekfFGkMKJRUjaUktZ
SZMIL3st/ajAT2zSbs35E+N9VdFTcSXHCt9gWQSGFPttPT+x/7m9/GEOPofGsblp
fsvdJ9DTDeiuXt1oTT2/nXEnHjSGI20DQ+esqUi89sYjO08qhwT/LLgZt1HitjOw
0bMnKvZR8PT6z0pHueemyd1TBFQYAn+zhdbiKfQ1cvht4BqIQH/UsN9VH0PhRtZS
PmGkhObPBF4mE/1doHOXnvGAWo/1xfrKiAhB02aE9fGPB+AQ6aG9amgmKHkjKqQj
9zlx3b/3AAXimf8KXuRbGhpdYy9ZlAbOjAujz/Z817jlqSAXqfMuxMLagcMmRWAm
i1W6dhO4dLBkVmryw16Jhk/xFbtCayGCKrOorc+Ovy93WsImXQsBQ1/BjOucmYWt
0tzL03V50quwpnRvduDyxVExm0Hta4rzJV/H84Bm0jmVgvWyEs6Yit/yr8Ph9CSR
65Rtbcj34NIBicoNTfamyUsrVtKOCl7NLh+B5rtvj3w+uVCjyVwpFveUmggJBqWP
j6opclHeCWK1D+3JZO1iWaHfUGeFPYAqyzeUzfAdS0Zwy3UgYnyIF9PFP5eOanMh
L7KRR6nhE7F+W3OUtZ8y2HSnxjof2PPnlfkiADtA02OVLkfECeTAaLo3BjhuzNPK
E6BcuekKUorR5iQ13ESEExSL70TNRSKLHsQnmpZQl+vJFM8NmbbDknStPO3SMaUe
Xupop8LmC48tiudDvYUz13bSMOcf4fPZYS7V1gw4ROmskJFI3EUQdUn+IB7s9inL
4A6kSr5qGUN8TybhbnKpIjiVnsvWgFBd1QpPiskM9Y5/+eYBT/ibZvEHnaS1X7IP
CbZAP+tsL1PEEOoaxXq49O7vISfDcKUeJAITFtJVjx/0Y+4/ZJ6GqQ/VzZRneDn4
PvV62t61m346qniv6LteTR3PgO9Syi8Re5mxIB+jqFOsL3gpTDNN4WJcJ3WAcx26
epItqvqZ7Yt45PRnOIISPlOh9MC7nnVNyEhQV94FQOVaEIZrczmpmI3jdQnRqyim
dTIyANKj/t2OFM3P1bPK8ZON5BEm+th1M3WZEFFw+oYwwvFjvo1NuhoxKbKB24s9
OuFmnq7qwW6dJu/6BBTrTJFrIB6IMsepQFpeFzlm7GJSLnKP2AHb6Q92Tr7pQ9q1
/IfMgLHmUoRA0QNdqimofETSO7M3tdtmALoAvlLGlmQNazSb+RRXc7F0uDOHK3QC
kRtFM3vnndW/q/CQmHfgC1NF8bo7qyjI7G7aLnW4n6GvkXZByO2ndVqbj4rvWLyc
qsFkcGlnnP1cLqjpvbRQ7zOSj+NNh9HWhGJ3rFKy2rkKCp2rZY9gPOvhz2uhvj5S
MBkQ5EaoUvoi47NeSKvKGF37O79IVMpXZrlsfgnJ9ShqCm5RO3BOFmjf9IEcrx9h
bpK4tLJp9AEG185iO9vu96GDqxY0VzBknaERK1GEl/ta9FuHYot86hHO5JCTuk21
oU6DDrw+m1mg/DViUtcKiIvz4BAM4ucj/CBg472BgOi54G+le1xW00yQ2n5v8kpI
UTRqD727nWAofHy0oTKmShC2jDOuMp6e41Y+4WKOscEboRyVG9fA7jOnOINQn2eD
wdnt0u01bf+QbsR+KWZshVDI9qLUopadOPUTfWXsOw01bOj15WyWxD/D4mKh5XRr
VU/6wYVAubXoRzhM1xU68hTU/OBXtgvwh80rZ0E6P59e3V6SBS/AoshxVCPqIF0o
YyTqHy5RlmKS5PWwd8lIvpHmqOLkZ1Fi7P9QhsrS1sF9TnRWVZjxmUKvTLUhnX83
wC96RTtCio2iHwwW9GWWdBcE2C2Iek09GDYsLms/tw7C0Tb4wo/gAXjJjrtGRZrN
2Hhfr23PPednwTPIF1uzRMkVCgmmcfr6FY38KJG4tCY6bjs9k5OQiHsCD7aNN2TI
BVTmL2DGiOwMg/a8Kdo4YcKGQDYyPWgvz931GHVWqTUfuIlHVv7YC2RegXkwtgep
iMc0WZ8/jRcK5rNjFu0QGE1btCCyo6m9BQXSsZAGbD+wwrEf8b4CyYABco5qZfN/
C6lHUnyrgEdVZThdCQOlU0lh9rrMJ/ca709LIZu1JgQlKlrBwlmK3NzJ0Et3pACF
fIAMKlMZCftJSNwqCQlhJoOezWUDYXMf3joEJstysxQIr6kv5tPx1ZQ3VQriUvPQ
jYaIfjjgSBufzfQ+5k3GC8W2YNg1RFwzeDas0AN9nSV+W+hgM/YBqI/F7YJz36kr
uxZQZfd0oRDbEP2rnpsRLWG5Ox8lO5OCdweftzhJT3tLebo6ABL9LixPIMesr37+
Dy7noxLOBDYYU8wdB8Hjxj/a4MdaVqatGCQrBV47WfiN+w7jnNhcMjSwddH4JxYH
qEyrFAeAgNFH5xORP5ZV0Q7JpcsNypCdJZPXO0qRxCej1IGhewQBe25hNoZLQ2Jq
AmeX+z19T/BsHEN/gGCTHcBWCsfXl21jEhnymg/BBpdKPH2KIudLVUG2LDPd0rlU
iGk6J9J4X/kDZ+iK7QZJW8rBYtVKkTuPh4srKgh0o7M7QstB3ERmjw2BlJlGcBJM
4mtkvr8D3zY4KM8DjxzFwxJ3O7l74N3XKCC1p5e94GIoq8xrZhMuIVg8xNPCDUaN
asQOWIavL75to1H6tEmX0DzMfYUkSRYOxkvx+6iG4s16YzEkm3/IelMvfgcB4U0u
+nMS/I7mtexGqA1XGKc9+kQZbdvocQZ/YzHKXFWjjfjMtQhCyfnUkrBET2hM9R/h
7QW74qfmgsTET6rqdTLCyexKUUx7BbYRftLx5pDVFZ076hFli5Pb7nyMyIRrF7j2
vSVSve5o4EzprjRpOADXQ8FtFsZJ0EsrKaUUsoGoiIuKNuK/6Ti9WMqmutQHO/6s
1nQxsiTtlQmY90Xjk1/dfMMCEVNpNAUG6VZPcTJamYlCCs8aZrjC4a5wXVUPzXaU
MEVGKbgb6M2kQ6iOlMkZMh6Oai0n2nBjf+s+pbP9QC7K/PoWWNxmQzqsDGOj07Dq
muQmS6G94PmSQTVM5F5WcKd75ye/QbxCjOP0Q9hE+eVJZr9Hq0b1YBS5A0PWkhZG
R3WhSdsX/4QxnQVysOfeddIy2LukuQLADN0LfKCJr1MOU9WAWc6zMcDDMe80bwrX
JvzcUEXWRF4pO18sXLaOGObjsXkku3N7iXF4w9qSNw+u928ghQ3jc/rmxS7pPk8c
3aoyqzLVxqvwTggnRh9dVBFxN/cBXuTu38wqL5qJBMZtMkXUb7vhFI4eUj3OfrxY
AEGvs4lQ3XH1XRvq7mgERuX2NPgTsFYRl4JwrY4Z9wt2ssQ/pHasXEQsrVIVxFiL
zH/FAtPXVr7oLdXcoxw2rXQu3EIcMMTnWQvm0N8jQUCZIdVRHDuY98vnZq+/lJfM
S3Q3YiTfVkTW147E9cD0pvbkKBsk4aG6s6icd+EPrpWeo54kvj1UYUL4A+JOzW4S
cdKLjVVuhABnwgeOFga2AtHmoTN9LwD5MzPD6aB8iV8sThKboSYAlCFOv3S8qlE3
SeszqqET8n6Cm2ejG8UAoODI4n+/oUizy+CDnQHbtVOsph4nIRSoeqfEy5xctaTE
1CO+fz4M/UlQWbUs26BP0NshtLyHQat3CXQuEqPaXu6k/OCYmC0KQlI/YsyBwHo4
I8pm9xA9N74f0E+RIyh20NFrYdeEEYD+gDHGIUbScqclg+ntyobNOCTU2J/MWYTG
NeAds8XQe3r7A9VRk69Egh52Q6X1J107/+pvI8KqDyXhaHYGj07NdGTG0vpVwM/G
mbjBQZVsPXskcEcu/KVLIMXwegsLVsTfwEwfX0GBrL+NGMrBY0M0cO5CqgPlDK96
uIb75jVmdhbR67gnRLicM3uNPYCAtu05ERACY1GCrAxhybLauEdw1lC0a82as82b
uGClPgTvFhI9JYE7vQb13I6IfVArWlfsJIKTaMqy0jnm5sp3BoVA0tMlOFAvUuzl
sD/pMttSuFqkxuAK+YobY4Cc0d8H64LqriEaobZ8ZkwFfs7dFiSVEDcUdKuMwVFX
tsfrwkzE6tzeC1JVmUQ8dM8PvrrwpNfAtibK98YyiBY2gDIjTQGb+pnxBEwp2jgz
uIFTvWnfJV8G5v6RWBpg99jO6vHbzNnfElg6543iaAc6MoRRdG/owM9y+BI8GcpN
SKEN1y5kalwiSwAFKFI1BlkPWMDz5owDT1TPIiTXL51gpROoIPm/bu31EyQu0V90
Rz3Y/rBvCsNwJTZxb30gWhe37UgM4wk35V+NDdK6tZZUHiBQjN+j5cVVNmQsAOQc
OKAaJ+PMcsnLwGETiSZyjn/PWWcCokfm/PQxKr1kZgK9VFlRNUtS6SgRXYpI8Tdj
lk5Jv7XWc3eKI1EbmG7qr/aS9xxObeUzam6SDReJrqo7kL4xx4aCdsk+p8DROf8w
B4LXL2gn8vY5oAUBDmGO96WJEEjlnY6RzUd2dVHJZVoQm5qz1dEyafiq1HRA0fTX
jAQ98Anw9B8qfxH8VqFHi0AZAkf7e8A14giMC/4B2Hdv6kIBYdAe05YPgsgAALfR
5BBlAYeKAGRRd2WLCQ2Skyb42MMqncjyzrA/puuaiQEiTVrY/bRBRd7jiI9FHPgg
jtW0kOO6NLjXVe0Vch7aIss0SvQLvXUw6xch+IaB5tbfSL2Cyfb2uQBtYd1nmW6r
Eqi65Hybu/V2CFiZw46T+d8czTxG9eSGdqxvviQsC0aKnHBkXsTzPCujDqzLxBNj
oCBMcCTfcc5Ri/tfelufbmc+Hvtu8pLqyJryC8KpKsu9AwDdhvs5WDDRxmcqtvY5
Ad3/JoRSPJgz8taohjZzGbz78CxLU8qVMPJqzBa67L+S2fHIm/MnzzUV+qkUy/wZ
JmeUUzpi75sCIXkgPxKfao8nRunQpA9lvhKnLsljbPpfrJaOYdlcvIOj5o7Z6OCd
lfrVYsCV3zzVbQf5G1aESU3ZjjvPQe0IVkd01yBLhlk8X9gnBhgi0KHY3pHfDS6Q
u45DnYXXUDxdC/YqSqFDJUhmZ+VFFeFCiIV+fiVCwBNPwKfI54gFYS/8IQZ3n2XE
BEUv+dSphkcLh1ZcLuOBQ8537VUnM0pLF5nxNC177hBpVvpURjz8ciwM6l9v5XNb
7umfI3WmxTg4rmm4FW8gr5CGFbr84MlwXFkK+tdUKo2O3fNMqXWWWw7cg40IKd+P
zYj8a5XlIuguRAwqktCzZNF1aNCOLTTv/dRYTRdKO8rDF3vIRrViUDxmldFiMnud
gK9BxbL09DArUSqpJoCP0bY1BMPSybRdodta8yUpOdAebx80TjEA+K4mKE/30Juy
xchX7NgVQp2afLTccRzBWbxZ3/7DmhTMbVVtuuAQOvH0BRdC7ZvqD2XzxCQU/oUA
ju19q+SCvjQrna3tSVM1iwk+IhGcAzcpW37EyTjaJNAJvIakVn1fvC3I0dY7Y45T
bMzTtsg+rmD7sIKz/7XurdKj14bvfxpCwR3vmkmPO6xSdsxl08xgbqmRqvR1uveJ
MHHf3m39wITw55YofE3S3GBHiN8Tdp1Jlsn4kylJF/PeDMWY7uD/KD6sQqYzpfGy
A9YQfc6IVafNnfW9PUzOCmcdN+Oo+4LvKWZ3E7JGoE24Z6Jvd+NQyZsXuX2F/eki
5QNlmcbLubh20dJ9O5lwjAdI/2RP6oJ+PZlEfiJWPu10q6h5RUJ/I5nqDtwXfqxY
1qmjW8M6M9iKoTsXPL56ojgA6c3MyWd3KdA7+8SoGnzQUe/4O9pQBf6C5gOldZ/8
vhCmkblD9wW3GzYZDzHKWX7sxdLlA/sIDaNidsDY4/EWWH5V79eZnQ7QseeC4H/H
bVNw7zO9hJPD6s9Ip2X+P1vb8mqCUrCnGXxFGWaZNI0grVOUhpvOOyfaUN6os9CX
belnqakZVn/LguZFqKgAO4VL6Nh4W/ae+C5VoRRrb8goZk2u8ZlYxe8HZ/TwkRkv
ETkJhAyiAmgXCLteGb5SylbSJvCU34vQzGuMaTKqn1t/DF2ytOM6WU5oI5oUkeQ5
8xWWHRxktWgfyTtBFfAUbMwS6Qy031BF2MM13yLAYuCxcuPfKr/arAymh1kO9w/4
MsFJkcMT87P19NVxsuhgH0HJnr0sguAWZN0akUQG10x79DS+R33vhODBvc9zaifq
vwp0dLja3kS8hf9dftOMO9uIYx9PoB7yI+WO8DasUtH1e4WXmDvm814aXpQ52/62
uLPlUb+bLAWm1CJa3nxwO6e+Qpn1YkAh0JRyVx8/bhWTJOXDQZli8Z1w1YkwTdP8
l3DOseyyIK4tJR1bioDMIVECt+kF3I299IVEoiP7r9eYvKSThSHhwCPWgaBOwK+l
cC4lP/DD0zKjUBrd3kAlMU7ntV4qoHqWwsdcdpxOxIGZvHLSJpBiPP2K8Va5l3wR
cEhf9ivt/GYpDyA5UWlZiqNgEkHTzouAud+tM320SO4E3x6TwQBwV2dRfhYGvVtW
UFu/1+TW6B4NXgwg/DTEjBLYE+B3uvCZ8BKA8QCSMme4HdejhwQGZ+Nrxt6uUo3R
mE+cOzJiDWIitOqMgdPijb1l7UdX5Zj3q+iK09/5CMvbKj2d+qup03BqfRA/yMgB
ov6x8cMt3HesGimehp/Gle5vZCki7SUuF19KXoIvDovzdT+a7LFN7BWIF6aj59WC
xOReSIScYNU7PwirS9OPAvd2K0j2MnAjlKc12wJ2CYsee3/i6TJ35x3rW+F490dz
ZV5e8d8tJQget6z7nlBlO5H5YTs0em8BRCtwBqxQGCSN0Icaw0nSX5efELd/et4k
I5otENs/TAmGdC4qfQ3YLUMFsI0LpneK0v1K1BwZPQsVamJHHLB5EjYR8fJHdeAB
nM8Eh0qNFdBnLE2PnXvMajijY/KJH/uteKc8SRl0SYoZZUNWUbU9Lk01EWqbNJeo
HZabUzhAWEsNVjfzVzFm+1zoKGLjBRCGDBlrthNbuifIULoeo1FNmwUxM9r5Y9rI
nWAYjLcpaKJyqVq+KtKqwdu3k1k4lokMd+dCj/WfQx16k4BBRMTBYlhVd9ftWYMX
DAsaARkY9nf2aYDnuzjBZ8sEqnLBriINI5Qxh4/JFb7gqaY5UWpMSxL8WufthQPs
ydF18alPuiiSHLEFjqzRf7qe8E4i95hJYAQJSS36nl9HBL1GW3U/D9076CYpM4FU
HryqOy1UeK3nDPzxhrdK3J+5fGAnDcrn0ehXOeBzd9w6+jS/uOOC7GVAvMhxZrrl
P3ejSXjtRR1aZsIYE3mHKsKQBU//PX0pMWUw0+JgYbXfoCmr+hpPvpmb6C21Ofgd
L2a8cqiDNqnmIxxI7XflEX+Jmwr5Hilg94EdDR8XfENga2zlF2w6+8GUggkFPzum
oXASfku6XHi1FMzgNoXSUNrv3fwSf06GHcjklZ1x6aDKcw4oj9Zr98zvvmXIk9wA
7CpLaf2sx2h/09lmDE76ITzt3rDMIVnEewOH1VcUNt2qEZ/nq0DFvO6PWxt2a3OA
TfWhEu415YkU5iHNydzYJig1FcMwt2bJaWAFZrKFiTc9vZ2hRskw0546UwVryNtR
cQUKPdV9alQIJukP1TgxcHG8I09d9LetEp0N+0ndg7UQ4l1ixPjKWuZcPQnTKNNu
aruCmd2UzwaGRTUbzm9OXb64LMDbW+Lag0L8yV8t//uX9FzsRZxkNeNRSTwP7EiQ
xw9IDkhBRKeXtL6uAdf0d3jsCvKd6e4sr7CdH4AOWXF0hzr6BT98qVMbteZoqtgH
7M/AER6CIyT/mFWeyiAcQ/UPRF7Jg+exwEantGnxMDHbOGDV5Fc6YVLNhSBUy38+
rt/W53ZAb39I9bNEzCwNmNCxufXFf4V2UEbqdb5ClZR4obYHDrOiHMP2H6SOvLXm
qruto2dCGzymOrDzIY0uxxD1Pe92d2Ts0hyocktckFMDKRqEXaWe0gQG3Lrk80v1
rP1Nhmv47FzEWgIFQtdzWjBYayrX+RGkR2ZgNPWDRfJiT8Ln6jpaCTDH8RoePino
2K2JVJ5Bx7t9aimZnnT8TBObB1Ix0qa/sMO/1SajhbVgfqZ1UoGaHKjbsng/pd/g
PV+t0Q4cp1bVaXIYAzWOxNMysk5tOV/jA0QF5PmDCUH4Vjrm+xjcAiggh/gZvsMY
CiKfeQD2n19/rkpL2hiNmmKiWNXTjxepKcqrqUD7ebKEIgY4zrz3bSi37b31VZu9
dLb1Hikb8TE5Cg+RtmezEv0/3S9/PFIJDxqIdRUlj02QmdOL+rabUEz0debZ6mKV
WWuKwzfTZ+k1NpDcRg/mzMmhucK1A4iv1xuYxWubH782+0ES6+us9ADmchVt7QpL
qPNNxcdcPtBrwYp1D/AmQJFovMBQjOIIIJ9S8thQ26IDSnIYMem1SObn9mRDPgme
Pj3lZIJvGP9t9o+ed7j0esJv4W09I6A34pR2+6dP5vXLhdmS2ywOmJazLabWExEA
nTE8f5EDpeyrgfkecan5pAEwroEF+k4qVgDvNUEV0PBLpqSzJCyQeT7DQEf47hCj
yeiR+WolFmzDrfAMo1rK9vAsRBP8kjDR6DTcycFvXEF7u9KpKYOxnt0zpBf/FCfo
W4r8Zfzo+gzjx2MN7YXYln0zTnmDKU1Lhrg5ZizDWXxxw0q/YcQzM/737czEis6h
HnhcH+TQdCsWFM7+t1s4b591oZSN8907TEJmqf/A6CzHtuu3kTsV/5vOvJRahyIk
ppYWGjitT9gMrHiWZmiJZQbHBCcg0ruzJSWBYYV8bTXmTh0zsAouN27OUm7P8Np3
AzYEFZD6tGz3nvN1qBOZY0pm4BDiaMgI5QaDZtI+WI7bxBZ8RXOySA9PFxbMlidZ
wx73G43T7S+L5Bt8Hq74adRIJmaQzJyL/Hu2IcYN6YYkGFmI0J2P+wBsERt/mLW2
NJivZk6CBHH9Y7NU6cPFG8GVhsYpLsjYa9TU2y8Vidn4dnLztv6DYntG2Bi6TYC3
EJE1KCi5l9Az7k08kq5e4p1iK6/ePAXVi5qOBWXPvpSGj58zSayZDtKqqw1nTZGD
GsfSxYHoZhsbu/nMVPh84NcUg8QKPtwz+JBtRGsfUkx1ACmomqOK8FoQnLyKk/4M
QZOzAj+sj/SuRM0MiJSxs2tDiCtZUY8VzbE8t+U7/IK8XqsiRvZjn9Rp+wNOJ7It
zCVnLzOcDUTAJCw+iHRuAEgY1x5lt8XwYEVoJHOqyuPGSZKiuXNyROPkSHUA9PIz
WxCE9aMJSfxNvjt2eMTHIaqHMbN+ki0B++F0SCtT3wlCsXuy65Ckecjofz02aNVy
hL1KMqvRwPQqjphmyA/ZS+rYdWYiSufBwWGxII2GJQ8ofmDT0paieo/sjbzhOCgS
G1MjOc+fjVuimdgdvqZdGQgdoD/KI1JQ2FsxJ5hQ2o611WNIOK/Rb3dyoW+Ks6vp
JAnSKmtmDXtLa0xPbjBUSpCdq+/Q+Uh3Gnq3Qq+gmS58mMQ0H8gwJWoQjub0dJ9F
/P/sQCt0j2mkoHRpW6XIK4bOhjA4RoV3whg7VmQDT/4EaGuw3uGoX/F4ayk/69ct
coF36/SY0FmR6fh0JDQuIP/kroUuRf04O69NWga5kkvQFe7fbUKsca/BPXSuRce2
PfYiFSiW/xXbtCNFmSFnNo/sJXcSDIsQeNHlgsbc6TwjmEPWwgLpScLLCZBGm64Z
mTfFFz3NoiCPTDuTHwEIhmcQxPr8DHdT8sbDgU6/FOrpnEGWR8J7Hf/uvgf7Zsuc
mUmrFWjGQvcVIFbfx+xG1f8orNGj/VrZi9o7a2mWGFc2qCcI484r/FVRkUQnz52X
jtxn62hBPK/mLSnmXaKks3qy7jfBb795I3pCKItOeu0SudvaVDczV4jk2BfdpL3j
YSUwNi3Ua2JPsiY5OlsowHcg7o2RzTAnCfeOPju/O+UavrmBdE9e4+/CG72bSnlV
uyi0N8y/041yi0ZNG3ktugzYAEtThemW1dPuZ7OpGO53lvD72xqEJhxqyt2A4hgl
ZZC9XvflpSMb16LGv2c8Zti+C6ybar3zFo7PNH8mnq3Wy0WCqwJ1KOCoM9rS7hXz
DwHDOSfbIfsEUXD1gWXHZTMhqJX/kh3hwryGRuTiiqhq33ZbE3A+7hGQwfsd0rnH
TBFHFuhrkuSgUAh+9cmoEAVtDxcrfoVpH3YPXaKSBDGKCnW4WqulsEHKccVDhSD+
tTvZszka/ynbCpViKR2DtirV3JGgqV+ahTgpkcRmREc/vZcxUu+qgChJUUygkAdZ
rwJNuEiFs2arwJyxsNaQtXwdsKzJkpTlBJ/67mB+rt9MlZ42Tu8riFTQGOZ8MD/9
tYtU+rEbFqQXyvcK2B3q+wueEjjGobFL+gB7J1TcckREWF78RnElmmQQX3A3CTHN
7S7FJFt7JurPdfn3w87gCoDYBrQljPVybUIZfm8Ki8JApsPybNsv2ey/+BlWO4XC
Rs8l9UHG6N+afKVSwze4Zi8leqdRD71BkHa9S33sax7Y6xPGliEtcB3bFBpwCnwy
DU/8vgCaY4cMh7/bRhmyPbHq42rWMvbSif+6HczCtz/igUs0eKSaJvpba1ufzZU9
VpIs3xydWaHKvkYvk5qRd76akMEjxgKFGeRiotu3DII42imnamjbYNJzOZw0uxrj
SLhsLzX0E70PUvWETwMCYEwjWMTewgdQJvGMRKIBY3sBHqEwRazEnUiBVdpbY5/I
ffGBLabGHDLR158N6V6esLz8yCOKb8UnmEyeh5bmmaPPy4Q0Kot3HsZSLWf8omdE
p5J0Fcmfr27V1/Wr3Kw1lcYDL0fXySzVJ6Mt9fsZtpIqpTquhS8xd3HgTPTX+s4w
Qz7ymdz0735aVt7gZypYvL7K8EO6RhWB/p6/5Q5AygKqLpCPp53BZwyEymfEAO+l
XNGlXpQvsCwhiJJxHqr639RGBYN73XlwvG8YUEtb8Hh6as0Bwp5RLw81qSgvsqNZ
57wmimHvJIKSzVtgXKfq0LSU7hVfLVmijwf3pFukMjkpadq2Z4T8tccgAn+bc7Kd
kDgo+OPbmT7l0OqHdCz4mQy2dbAZDVegYnuFRv+y6nkLKM2NA1jWpJd+Qg5GyKEl
gflFDS1ZSQvLiQ0dcPXFnx3cCJbdk2xlJRtunmswdS0vTNOnLDitQQRXEWX4YNnG
11fmZpk00SsXUpde7hY0cahm383xVGMeTf1uJiHKyFO1DU1eKR9ol56dS0E9SlU6
hPm9K1IUhc67VauCfme1/sa9VpxPNU5cL/+1wk6S1K9StVzCI+0SPi6CvLNl2iUM
LiNV1RPJcg2QUUEdtW0EEqhhO8x7uifyx6zbaaWp9tpRdhGbHxKH2dDEULi7d3+L
vCA/3hr2Udi33kuaXW/TK5mxj3F/KK3ERMEh87zDCfaPkfFnuhuV7ToHFFTddXKd
92UxwPpwq9FRNifROiU/2VvvQZQIqDUBAm2mscLJP66MEg4NHLrDMp+4lfUYOkbT
bmAvsSDrF9ePzkOOdU5RcVio0ejJwZjdOHVEC/8VlEM6op3v38d+p1RCVKUg6MV2
Iik/REWnmv+EnGThWe2bDNCqNOkpVfbWbNvVFqV4lqxb2qLvl6mculBXbj+C7fK2
8l8HmPEqYulRaWymDRTRqPBemi6oq8lKJixi33r4mTNHt8d0kV0mojVC5g1v5MME
p/Dc/htU1RNnBzCodjc01JVzc4M/QuNJrt6XMdbPLQwRFGOWS48zLA9kHMyHUwYi
IqZSs9cMlvU5lFvDE9mL/0CO+GtT9i9JQxNqBrbmKLQPBGHkLu2j0+q3itI1HLiO
6yvpHEPSbVWSNQ0m4oa/+anxHd5wTgo7JHq3oWE/ofMEkHDfGgrfmqR3lHMVbpuc
xzfRE/ZLQuzUv1ZYvVVdXX8wtylcwo3Bm5+G6Dd2Orqii6XjEaW9LCWSe3a4+TTE
7fog9bDCIf9rVG7pewkb+1A2b5TDzsjZbAVHf8TPbxgbTXckW6P0BtU2xJxEUMKO
9Vjo2oDVOBdulJU6JWx/Z2fzSCYumfMaop4pu1pvM7CR3u8f4z4pR4zcqfpRf+vK
Dz6lNU2HEK0qvmnnyxqm4P4xbgpf+hdcaBSIZHSM2MVxwnw+Zqw2Iq7/MBRunEa6
tLZeghUodD1Ljykth4yfYTqhJGQeo+oN9JnGo0YgepAdqVj4gFIpnjn4BCjM2Tvp
6YpqHrBkIdfBVqyc18tVCeDsnZTZzKb0FFQ/QuG+/Nxa+Oe4sbqUDTVGnv0Jg1FR
nTbgWhOEMMrhcnNXG22RJ6k7hs/9MxxgmxPOm8JdR9LdKYIHww241FkIxAUQQJkW
5E7u22EWhaStb2L6xsZc0yz0Xeik+efk4hWGwJK5OPpAPiihz9izebc3pcePsjF0
b9l4w9ZMuBXCGtPcxqPMTwrMJpaNBBPEM3EnVmK3dGYVGmYZBvVz/8HvD91LIWMK
pURhTyIZHIkIqKV+4oeUZpIrpP1x84Bdz4jyqQk2KkWRMmaYmDXNVtWeHlQxaIOW
kAdTjPbbqgiz8S1wUsDBnQlQVv3rzcAWTtt1KM1TTfeF6uf3bkHYVIfRczbehVX2
EqSAjbUYmDZ6Fh8rNAgb3RCNIlC9gp9VzXZD0fo+qWMeGZ6Ce+Fo8vsQa6QPgCIK
j5VmvuPl5IDALgP2fzcaX9GFCe4mDwprgFKDHrzS5rQ4Zg8qvPmzWxrkhnFvry/l
MGn34U62bc8DM37EkrPuPNmnJWJGqmsgvz1k9WZWJLAM9C//dPx9wrpIuDMvwbOB
9lqgK7P9l8x+yZ+TxpWYqh+T3M53lEP1e2+7QBSz1ddTZat/KEColtraSuw/Ju8s
GgEJBJSGZN8/2YZv/PZr9yVTdUZtAqONePxz+KRmCgPTFPIg5k9ESVGBrjBZNg3s
j3QB8v7Brw0Oj2rpNFsyqs5nLAZH4czwylQhMoXX+WBkK7RviTyidyFH/capxk03
B2/03wcviYyKlXjOK1YsN2whcs//or9Ie3V7otzB4vwyxDWsnyvadslReoOk67Fa
voLvljgOf7mqGQ+RBThSvvwMg1Y++54ACSGT/kPej5GyuJTbxyKyctJcvfGaoe30
LH9Td+00P6hl7Y7egBIywGVSlV1lxkIMCZy/qgmSllb6W/5+HhrIm1vkBvw22Qis
65zL0uAgqVf+HD520SrONzq38gfccd+1Rvi4iGxmagme8l/d9GLlPN6CYK+npRm+
8fbP3RE8pX3zqie2u2zG/CRjQX9YDyys4JPu7BKI8j32P1vuKL5tcAUZgMvalvdO
iN3XWVZCCk7kQVbZxmTN8xKVR5QAtuHZTxWg+l/WyxHDQy7hylmXuXqEPqfk9Hy9
G6Bpb75aK6RiGj0ZcpwTbDfsIlF5DNvxlHvBs0cLRiaxs8y0tBtl2KVMgRmpiNT2
i7u/RviE06GBnmv7t5akYDoQ0FVt7H30XmIltIygUyFaGaoYCqzs8sJ2cPo1F1ZM
CqShPnmJjmpmPRtUU/DW95RR/Nxj3ZmXh9+wydguNdQK5VIOLIJdyfQOgRPD/NZi
OdkDtxzrFCVVpkN4duqybC3ZOt2dSOKyxf4eQ/Lr4EezqO6r7ZBgKaFQE5AeQeay
Tv2nTdu6t4ypC/rA9qFRlv+OFBlxSSJ8kAIVXhzLYag+fFBF9k2L4qTK+J/qPMry
zIuWMd32yjsczKYPWcpuw7mM3OJ6Zv6BoGa8EATbrzjsDlDZnsHZUQPDs+EcW5K8
HAD0cqqoZGtSzaZ1BEZGAOANfg95795HkSjPHkv73LM1IokmXQPF/TBwiUtV0PJa
CBeXTXCdA+5tfS/G9tP9fSjErqmgwTtCpZlh0zIh3y9WHCAGAHU7199gAYcUY7sz
54eE/hpO4urum0+iLt4z2UosH6shygmqao9+zS5fOsSDANC8bIjKehrT1XHGZidJ
vgp95PAETdIom4qukSXfvJ2hCI7/Uz036Jv9MYM/ch0ZW2vslixNYk/xadt6PUPT
M9dPAXn+5bp6Fzo3SyYGenH45gMIrGFR0weWR7zyfYJ6hxOaQ6r+yN6begMgoxx9
2OSQ8A6q59B+EUg77LXUSODgKYT5fpcyJ6a+tMP6ojy4FD3j9ET701ll2KxCULrC
U/tfvtYdDzlQYTnTNkvKzOIqrRzRhGAZqDcIZ4epCZBNKwMRCSJJnvF4OuXEC/io
FVVoqs2V2gsd1NUf77Z2GyEIQH/Z2N2S9Es1dT40WepiM//A1XZOdNesgxk3yNLu
xNouqfjtlI01RJD6e8xEcyqKcyJPIwPfZe/oQvkaD4xuY8BmbM862Jsp2gECjrbG
DtqZgseXr4nWOUxAFZyCGzWP04w5jh9YED+x2YYLYWgnUuFoZ+bW0pKtuYHy9dmu
EC1PYtkTQuSDkI329W4wxNmUpKVGXmhtMp/ngr346Pk1nYNJgiXAQNrsO0Xgb8UO
vz5epsdb4l770Q7Tkv719yTsi/ZMjm6agZ0KftmF8+mA0qov5f5ob16lV1NVyOUB
nYVZSC++brJhk6kPDlgvKWZ0q+5iykrssDXA8JJAB3H9yFexRhWzM4kVdJw1GevE
E9JrSzs6RlSayGgNRvmew4+eKoxhRCm+azYLbtrKVSuakzbVBfqHLpsNdEEPmFHz
7g8WT/3JruVzRJYZ1f/gX3pMBUwvGySYszuB8NQbf3r18IW0HmD4VNiAr/rQB1x7
Da1GNgj3bQJIJW+vpPHOIBUc21cvEF3cgQkTAZyDBoAG/2NFmvdrU/Q9ycUySlQX
TAGclgHq7mzwTQJyRmNt0ijINQmHsNA7ARymioBM1ROCiEQ4oBqKLpzfdYTgk2hE
IZuoj6oSaKsCZNIKYPhTtdnGy0XfvrgHd0n6h6Ou/BgOdvOJPMSdU/IcYm5IvBC7
U+b8ut6pOg7hm+xdmsO4ddSRjwVW8GgkP+Q6MH+kHdhDNS4Gs4c4Huv4X2tTW/Cg
IfwS6ck9MR3xHmJeKVSABrTRU5eoLRHXQy11p1tQ7ITfSD9MetJtHvHo4xwqCwMg
tE+pzRibeOgdVkmYR/PALxbMBCGGt9TO5ZwZq2QZkPmLBxryZ8zwj+RNWP81+ZQT
HHMKaSBCO8sob9AUI7iiArOgSOE31dm18p8QNjgOXni0DA02BSYARjZogpexUtCN
hUNWvNFOjWekkpNvgEj2AxqTRiRUST4bodLySVTtEU92Bf7bPJiyw7DjHXVtD9Hj
KpnMbnOY0Qr1l6fbrKPMU5P4Vj+e/BRfqmAyo2CpU7VrI9ZMhOuahT96Ojz3VyFK
zmin9z1mr+qcrWywq/js3arPmfGxePQ+K/1u22spi6iDT+ccmYQXOALhhPrxpeS/
XZFNOF4tkvEh0o0Dys9iWE5CIutf5PIZ6+Xr9wKdVZI3hiiRhRqT/NHbQ/e0AXvE
9yNmLwjKYICqeOWSk1vYaLb2WQJXf6XVtdn3/Qhtj2XqHnPcx8pcd+EDC4JxgiRv
C4zti0qcT2sjCIy5Jr76R5yoFmf7XOhz/4zhfvIRBw2JXgjNbeoQeXgvPKIByg+u
3BnqZcMbIX40Hqf4NG98JcdUVhD7D77V2mzGqKWriLVHCE24NLdexI+eAQ3KQb7Z
sOwD5Yg8w0jzIVCtYdwSM/DE39ZpnrFvjkMce48OI4w+YxGJfxrQU8/ZWU2I6v16
bKjiigGasmzKXC0IoJfcEq2Ek5OX5b1ycY5aKENYqOPc2Rvck25fPycasnsIoowa
sgJZyQwlqt/uSWv7B8olOSuZJQyiQ7jXchZQo5hNGqD0Pn+jK7RGenPsTuHe/JHL
OtLqSd2I+xZDCzIOmJHLGjLSazGq4qGvsGCOSQFLmMonW4T33csbWw9196gwrIrh
7YyHAOGRf6A60l2wmAByaL39dZgVLEzv1oTDCmBHjjv4e8h7JkUS4Ms+cz1Mca8R
pzgpjwdbFPFnXk58IO0vk/A1E63N63Q+au0pNgMOpvF03bUyJCjM+lnBrS8f7gmm
U9pRLrEH1k9lebCyYUEev7rPF58UcZ2OQcKHY7vVJoiCod3GyFLpKUB94ebIxQcH
cKhtS6tQ2ny8ADaUsyXh2Zxq+U8OtEMwp5Ip1PAJsL3N9yOdvZOL23YijVKN8kjZ
HtNgTzMh4EBuOtcW530iV5GPlLNU5OXanCtOZeZvGJpMzDSKO8UxmRuLZIocWXHG
uj4nSFmiMGjg+/3BGfJHr6JT4W63HrDpsIiggYd/7BW2NARNJIJcyLms8aIRqxJ0
uTxBUZyoGpazS9ZFhlZr8rUBrT0f3x2rMuIqGtcwnR8a2Xz2cRW2ezoKJjcP70n7
sweU6kTIeFfpsXqwtz5vecqJsoF+kumHIg4IptG4j7Ve7+okkIzzXUOfYY6Nmszg
opI5A2YbnD7NjAVLKjr9HN4/bUPYyhhPXMd7FzY+IoBJ18sHXQz5sdfY1Xrm54Nv
4KiNeoXeRJVi9TSOY4J/8Yljrq4GYapf13jC9STgl4zNgfw02T/Tm2CDc7klSSbw
e8zb2sDhF7knuAnztZnqgStLgOJxi4ts8PCSV3HFkP5/1xkIcJ4qqEGhT4fJeCuc
bcKqsCHx3WfGt3vWCatxdEs1UC0uD1Q2Kq6VKcoRuOVFELqb3F3Bo6T9txlzQgSS
1v7cqxf63R+a2vgYYP3x9dZ2x/2ZkMFxQr7ZoQGFw+NdGBpqC0HhUUxt1HUbN2iu
IL4N5emSRD2vHu+a8zCRgKvN29tTYknw39Nq+UJH9xZbYQ+RqD46otTuvOO+stZ3
DRTSnoLz15yH8qJL6Mza3scH5KAR3LAz0kCqWOkzHdENoBPMMUvOBS/Ku0voDg8B
QsXrfPefaYiSCvc8oYWpx+iiU4xd6+907bkvBcN2eyy0lARaf7KY0iCW/tVYXqN5
QVoE78nRzQdIL5UTcso5l4DrPCxPV9Vtg0x3ATIrEluLFr21W0dvSvIxkOe4kDmQ
fzMSRVSv2P7y0rC12zY6+eqOe2SfFSM5+UlhzcmfpnKiky23XPPPN9NPw3+nqOMz
AhcdbJoG8l62OemMQlhmnbeJJS1bbD6GsQUKnQ137/AxktNB8igjMqxLof49Ei8G
+XJEAyHYKn9HrMT5kAhJDP5/V676NWEOMLJcIkMElNXEaDGBZwwlzSpdXk97tu9l
oepNCmjvAMIWA5zAIq3RjbW+3jCo5sSDwicgiFaEd43j0IujqvKxfLuXwZn1KrIH
m9Z9GQJS4ICQTnHB8+zKOfp2/b9YBjd7gqVPANKh9x/OjXFA9iv/DIc+xSP6r8KI
5XAyjjfrJ/KuicGkw4YinSRu2XNqYK/ueSPhP1I6JBT/yJwny6JcHakyPPeneqOT
NkwR7duhPXc6I98aaQY3ohYyhjwQ0BRfUgJIt07uF+FJxasJAZnyhMhnCStYDIoe
XE0A9aQPcFpk09XlfggB874ennp0Bh2I/Ko61aEImEWmTKraz1Nv6QLQC6eVDByt
yblAzynJ4CNcrhdMooE2q+YC61TsrZubEe8CTsElXCTux9XZraUW+cUg+5mD5Trw
u2OZmClFor4HzOkmOOtuBY1XYbmgSBFq3GgyHAeDeDrij+hf2qGTMK/XF/1XBC/r
WStUi4Wy1x/S1lnLcM8bi7dRSW/ioqaH38kbo4NILGmJ+2elNAZUiowT6oeC7jq/
6ASgz9+2B2BCfRCQvqZtY94YjsiYTycOARv5WqTnn4IG4uKPPttNEtakZL2TW8sM
Y1/0TgVWicCA+uzMHlXehXqCdBcN7BClSnQI5EGkTslgwEDKv1pB9LihX5Tf6HkC
aWI62QDswZUcVGPhluaWk65RH34M0qBHAWijig6EHjCdMvTvr02RaITfpjhhDoB7
kL29WkKj/855og5eCOqixMQxzc2+mvX66dSXSjF9vBYxH7qsUUCCr9SYCi23yisr
iRWzSqWZcrSGq/n1KcPqSCVTxWeNJFevavS4W/fz5ysvvG8zr2pDhtIW/93PSlfr
p99rDeYYDCAwFYL36i3lkgOVbluRpatHfowy1gY1guZCI3WAQfRaf7xpk6POgkoh
AAEKS/QaO4zbBj15Le+z3nZi8IEzFqTpNKc2lYYwyU8bKo3x2zGAwNzARV7xV84Q
FpDmhtghc4oEfjW1v25+HOrAy709LXscvH69j/eCnjYBoBYb1GnVEQhtWmSWxm+Q
9ndWjImuHcHxSoPAZIJTFo1yo/T/WEe4iVmCE7o2ogdobfBOMFpE5dW0GCV3R0jG
WtdLTqyoXrjVCcmkWj+I3LJTALDyxRzOZKQbNZqb0+7zsFqYhSuiTAeFY7j0I0Kt
9yMRwY+N0uMHm11+FlmYXoVaMbBl+gyqXxkE16X9gsuZceY1J7IQ+U+4su1KsCrS
/nKj0PNq3+8u5NMdC/WH5B7SaZ/moDfXmreF0cTbJD7J9mWjSAT3b0ui18PBAHjW
ROBVnDTpksqy63ObWxiqq3AanDGTJR3CbcLMn6OwMOA476FEqRtcJDRn3qQgYWOa
dP4ne0FLTJQppDoJhVzOG0U1CofAFcLTAosJZHGbHMjOREVxpUfSD9HsiL89mV8o
50mFVauWPfn438ZjU2wS7Xjmc1NvSTuRalsyYN6TwstGwBH9R4/rRCzL6TueVEwx
NNTFWHnAARAXDQdvNFnN25HS/6utrF43ys4OVYnzqFPepFkKmryh//0Z21X4ne1Z
U9W2JABSSzXxYrV3z2KA2HrWAQDVppQqYc8fqIckQ3s7rQsKa9CkIMXXloChS+Nz
fkwFzzcnQj9P7Kzud5MuCpS3ACsCrJQRCa0eE+Lxf3z+9rqCpflaXWNvq+puB5G2
IyboprA+nTJ/K2j96vwqwFlVCoHoRfRI6dvnHl2/3S3kHUL66am7ryEfPzxwUYkl
SgGX5JbXL63NJMuY5GZ+Mjn6ubdAyDDemNBntgvGX+Gmf8QRjSkrSaXVJ14FaQn+
R6Tj8+wBXJo0QdiJ3jQyO0eQ3047BuogoV2sxuh3pqQfhrQAYGiO93DztCfejzOZ
DBhaqN2fj0zqJsbvjg6aRn/GrHgsBlL/0Qatwd5Ct4F+h0rhknPz6bI3xkRqZeRC
meVxU1W104sL4Y3WUr3yhK3H1fOjMzHxbqbLPaudKN5YaLsFlJ4xspbq17wGMB+d
nYdPRhWB4+WdrQLlF6dmDvsVNjNyDpF/d7CuYtcbgB3L7/ZJevKwwG/gLlEiZI5O
xZoqDFiM01ftP9wfq+iJ78vlTinXBE1n2uu6EPSRZZkgAV0jrMTf7oWDdC3jtewR
ARb1Ftkml+xQAYjh1ZqXy8WpEVnbFMN0e/DUCGvmqo0/DYwOOqD3Vuxe74HggZ7u
sc1pwgFhNIqKsuiH9E+mr+7Trh5OQYhBO85oCTvHYwIvLUmnGGJo9sDPqp774v7D
tkNg8Gcm+BIzrokahxV3FPAj2ICgwcnuV9XFPF/3bs997UJd+qpv4algle+D1Lmd
a1kxTJPA7yQm7GYvz9ge4HhiSY7tqbCydpzT1cAP+xTGvks0cENxoP5GSf1rYLE2
X5/3T8eHpkJB7PvEY3WJ6iYx5FhFUr7+ub87vruZNI5g4ILNre+pO5L5zuo6jdFI
5dtr+C2lAs/ryTntdhsSGVCZpq8OI3WVBqI4vn/2j6ohml5Wu1VJKR+KretHKM4X
tcUuW8rrI3jIgraZfxVrK/m2tP+u+5IoxKixN1pA57vYDjeD1Aaj9a2jWXwnWG8W
i3HppZTg8wsbKswxTFxXr/XlzjrXdEoVDciMlTAeR2w1C+glOJppObSDyrCLFNjf
KOywL2K8/hol+SZTCw0OAeuAnq04QKEYYsoLSmo6LwINZTq8IrZXYKO59QF8QQXH
PuIxmzwtw3yS0BaKyBxNeA92dDvAmxV3GeA92jll1F+xu69naSIei93ZnjofJGQJ
AC6eJZ5FCeL8i/y2XPZJz7zHYHEVMub/JJQKgMREjgnphSPgAC7PWZPofnhOzpzq
2m2v93w18fKyqTcqcQtDVKJyaKglRelXishIOokDAlnQ9vCG2mqmfP4vuFkjyvFE
+EOuH88CLBk95KB87erLggWY9BgmRTgnRu2N1hxqivBW8As1w98M3AW0AxB5kaHi
dwOQOQK3WrQQELja1hqd+xTnq9eHV2ZgBdBROjNYVcbtUKcfcv18INTjeRLoTKNS
FstPhiSOhphS7L7LMXyB4BU7NPPtGB/AnYNoFIclybKpUm+D+EcDHrX7zfCCnLfu
qgI8opZtelsKTED/2pP1bZ47ux18r7EBEYzZ6+ixaKK8U97xv0huDRtkwdjA/B5H
CxC+egTPN+ltSzowE7hu3qMk2TIru2fe6uetPgO6XHbN3zb2TVg3XPfNOnjibJfe
wQXKwnkSAzDerwooYpRtrM7kxlXGPc5wXSExgbhqZAjfwg4K3zRbxNKd2RjPKdBJ
76bfIdq3ZGKTk2R9+3F2Zv+/v35tNqIvTT6XXy0txITo7PsN/to3gIoiCXhzJQyM
6LtTAY4pQiRL6uVmJmSWLI7X4gQvvMmQ6dSlS8khcIZB7t9wvh8Yg+yciWHnPxAE
0KQAUTPaZfS6YywL1vrHsCCoCn5BWvWW3T50uQg9v2jilmMyJ4nWRbcjus0H4Alz
1cka9inmzOb2QCEAhfaYR0w0SLmksUw/L8Y+oYtIDEfi7VcLdfM8W4RZquj3CuNx
B7w1RcE8eYro/DzVkUOei3p+osVZnh9DTtOKtanBpm5zhwMLBYybnUJNlktTRMxK
Eu+L5f7PXmrYPnWbVew9uD3gkU2neulOrs1wS1x4FZne8Iz7cgPsYWpPM5mfX+bP
dQ0a9JA3kh0HKHshLz/YktiJbPkoGJbWOqUI2h484TzOvopv2akIPpGZj1ec1Nv/
ue/mVQzSISlXTH/KwKseZQ4a7VL+9Jf3NNXCMjTNzeZ1RkSbNYlAIBoaGdD9pZJh
82+7t0cBvBgZsRMnG9uIp2hHn5bYkjtreR1Cne4cqd3cWsD4k8w/e+wPTDwK7Rtp
apHMWu/kMVcGds0y7/MGPLQCYPRWR7D2QDpYVilNgY/N/zhlfXq6zyGeMfmYejHd
aPH5bSrv5fBLiFzT6QaKAndoUY9tMFQL+mYAMB/i5WlsSTTFz1qVXXRIf9dHDRnA
9CqZhrjNTOmvxWn37qhegmJX1y+pDP3eSfZd9pLwAarMX29qOVxakYse7ZkGlvfQ
qHk4hFdeNg+S0T8LeGqp2foZ8Twa+8WcHNM+T5nve7E2AXYjnYU9PwoJf0RH9B0/
XwkPZhZb0AY3JtGgikKVDUIHR6SSlRqpeZcPf9G7iPWx5itndQ/I0P7a2y+3mzOr
h7KyqUNkKE17kzIbixJXs5sxpqXGHF+3hD+9J5To1aDhHsI8Is+qxaXvlwufcNUH
hL4OwZtL7FSQhKDOGCgXZPBo9VvVNQjJ7sSxUz+6H+RdBvdyQ9BbEd+YX/zhTaoO
0nd9F+6IA7dA8Hs0tt3YZvMF379HibvPnakHKHj+AK7O5N3M/zPlD5JBMyEaifpg
j+gk6aPttqmnehei+Y3IB3EhOeegsJ7az6N7xcpf/pc1+I/6qOLnQwnwXDqvXC5R
zYkjXj7HrKL9K95zUuIbANu96F3duIP3tTxXykWwpwaZtChvOI5C5RSIXCkvGNI/
HUzwlKz+c9L0Ozw0kUIV4rB+FDODlaMRT3ZpcDx0zaeClYvyXcs5aK24wntOJ6xO
tZ218BEitF6FtISGNal7Ro9+LVodSBNo4+DqMr2fkFu1dJ2xzt/FeWHIS6w9goCT
+N0gh2spe3gwOdX/vMOYgaEO+FWvaSTbWlbiIsn5JwiyS4aUFX8yqgy85lgGRMXJ
MyV5WAXp0H5AsEByJzUMe14vKhk7FCZTVgoxjTyZtJhNbZi5dS56eS4o+giIGT8p
zr1o6ATv8QdyWuJQ9uaEywfsK5FIcQRESyqDvcMqDmcNosZLKjdoIWq8XpxcxoHR
ZdHwy+sZ6FIjc3qso3z8oLMvbbvj8ev+r3HjDJwReRs2DGpdYaG7OLmPYYt5vzNM
5HGRtS6R3qd0fasZr0F7VyoeZidY3YPRi3YLm6b/1OhoPky/KJPbl9R1InxmAUu4
wvXvF0TDY86H9iVJ9gGEKrEkmUtyrnVzfUGUv3R1ToPg/Yij+FTnyv0aqKESNdv0
9Qe61UHn+AGawzHobXmbiyz7l/7ouNVIUUrXiWAWrJbr6q4YEzuaFP/qyGZctPs1
ldrNTs4nJ/Cf9A2eGfOIIaUBxP6DVud+EpOe8WTPqhWUu82z9A3G8ODr5F1Bz18H
fOTXNbH+6lvuMD3vVyTqGvLf7FEdrRg7BsYIdBwguCT3sPwHaK6GvrslMbjdbNOg
dzUgpj5pkicocphWNhfmy/AReXZ/JqHqgO4LAJCOQ4nPi7RIGwq8PLjUdfuqAW7m
cC4GMvyvf8jBCa7iMP3OGYUaDEjLkLJhP9ZCnmXhM8l3KoOTlvkrmylCEJbohXPM
6WqrUYgvueOT2Kp4XFRApKRXhjXQzGqhcZcSMkjges5wPNzsnNkjvK/CrlGPP/Rm
PelxHd+fVGjjfPDCvjm5sx1DUq0v/TcFtfU7/oR19epAKiC9mRUO2XHotK+UHxZW
dsu/H4+8QFDh4zxKvxpshZ0m0by2wDhmssF31V3UBFnBoqt+7hpcpzcv7vtJKFjb
psD1w/Drh5NZO/0t6wPcN60w4zIjnXki8ZiLznnIjkuZMAjvxet/0fPfdamZ52pb
EL8OaLJeFLaOQGx3OHChTBd3FNlQg+6Zi2wTZQ3kSjaGOq48KmzX0ADPOyMqMc5X
yhvv6isJ9Qn242uoedBXz1dhjnlUqFFkl+eFisqGyP9BFezjqCNsgRoOBM384Zwv
WBSjWTR+QJXmp5GHGeROAAGdhfpqiXjZvkDCMxmrQ29HWM2i6IPx9iPOloyl/PxH
hmS6/xHnd0vYYxpp/e7oLFlohZA9+12qRicZl+7UYO2DInpyTeFBVgfLIQstU7wo
kxUymHWb3/rJ85vxd2z4QOzLOVjNmklxGPonNhS2a+/o7pmjmi0/LoMATnYSxgrC
MiL8lcDvkgHjI7gK0QzxmGB4LZV9eaKCWqI5UCIsqVkXbuEOxHF+lxYYZdRr9LoC
J6/OseTIuk8AeBjHkpfhVfD0Ek2CS0Rwi5PXS1VNOMe8J/0ZS1JxQ2XjIHDhw8G/
tJubWjRbHDwT5Gc4p/OOKl2j8v7tKJO7cdb+kdz8Jic5f1DwVaZlZ1LtC8PWnixS
BC2Hef2bRWq+P4prurmX1xnW3CpD+InjK8O2HdE3pKg0grq9pnarTZPeTDUuMZnm
Fky/X5lc1nClyxB6WVCkzMxZKypjLkcU4hBOLI6Pzqdeo+d69tnVGGNl/um/eIbJ
BeQfnfDj3OQreeoBWmktNgd+2tWxOseShg38bcZJMWG2aOHlX5mkPZHw6Nzk2mRp
Y8FeflOpB51G+8Jixy7F6rUz6HHJgl6qXNR3rcpMDvuBCMuNMd+VK6cUEj0sAmPg
687vsy4L94AsAXYJ38ppNsCGzXLafvgD0Yx8OBknbLIP2j/xyttWaFDip/VOiubK
OxTd5cK5X13r3rjI7jIBN1QrAX/R6gxfBWrVZAoIO3MRs8BmCOq6evnQEEOW7c62
F1MfJwPksvOGXxP8VeXgQTAnY+n7oHjTr9HLchoHOWaouMBCA7B5kUIY7qK/3fZy
ewthQe9vCtcH1FW4CwlE8xvv2+VPmSago/59xnqbhy2V9onJnqdWYoICLivVYwPD
gprMOlQsvJTBIy29+NQ7ETHl3cVUH/b2ny40rvgINaOB5R1jSjNbd/S28nh+nfGO
J0CKok1quPC8FW+zUN6DTv1xzstMU7p3M8S75s6nWnvMKFRNNZhjUJN5MIxEE+Rj
Q8PRUZtMJ2B+97Zko4so4PqGvGu5a2g/6TPX8UtMn74id8cIooeijAE34Kw3yXQj
MFs12VS4waGm/Awvr4LM4mfT8xwQlZ71uPdrzpJQaW2EAnsqddJw79YC9HmhH9lt
Xzl+4z2taSrYLwMaZV3kdW0P8/PSt31iOq6UPBnCT2J3y9/KrmlFintt18byX59v
zK+tve7cekG4KV4KEtMDeLPeDR74iLQlz4y4nmCdxAq3EO+ZqXR01azNsv7z6kkx
lBdoCUtyR74qf/OSFvIM29lqEKgWbDiYC4uCJ8sSiItiAWQMXeCCXaGzt6+pU2aX
fc1RLNAXi2GJmyCg/Rqqr5MkXj6AHXEzoUFfplLrglLcdNqfRX1N2+UCPQrEl5x/
GfKUJlFIvMlLDKHZAGsXshczo2qhZxNW94IOY3KFtWpdvfZUWsSufWiLE1+rRZ9/
UuFIYIp9kgQ1iQbqK+EF25Nspe89pvFU1QxZc0F562sNWCHgvpRgw25CjjCdsor2
vicC0pSrTv7kWKEV2ferj9hxnktpQV30ntiZ+Zd8NmzhIWaZ/6W4oteGE5YDXQ1o
FWk9CZOt9Y3KgR8wUY1Q/BnuOQn/BMgVkwkszxexCNxlpmbR1lelZOF7uKc8PRsZ
yzQVImDMT+Sue65vFMumI1/dmbsS8P+C1aGM3QFCr/Kj2sET74r4IgSk8vJdKCv1
P8iXidupqZWNvnQ1uMtF7T76qnqLP0ksmSrSJktP49SwR1zoYeFavnW6je8MogBB
M7rOapCKA2VEGfU1h04toEoQNVLcH1c2P49HMvQDhxPd1P2vrUre2u5cIPAxLI04
Hd2uMw0q4G5d8onp1qjLFBvKvA6jHN3/18SbaPeaN3u36UXJVaL0xXu8QuMp/6qD
SiSNerSr3d4BGC3bHpBpJgLS2PR3pztoZ6/UsAxLmx+wqYwwSIfrbRxVI5vu5bq8
tbPqzZUVH2IXwPWvPoHzH1vvsOntkwZutS25Lml0KOoWxyxWDpk9FM533G8GihTn
1gMWFZXOCOSzPdW3YiT/Wz8OIny4V4RsoV7xUHRNkcMKzn3N7rCw0DRAcNofe4ZA
NvRfzsm3qCasZ5AqXHCA5MFR1JQ40+ZBnfBpskcN0NQbYLDBlyUYiLUgLAsWku9P
UG5V4Ur9kKpPZj3QzpoD+3JzpJX5/GRlpiIgclOQC/C16DIhOIHjipg4Y608Ha01
o0IirkDC4tlhy1I+vM8br7+reLh67qSJ9UN/Sz+Qpd/ZGNrnS3KqeE0DK58bhN28
H9Kr3nt/+9dqrF2LBmaz2Pv6VcLn8DULazJyGqtqLVEqLSXBFHEtWXWtrZAUI6WA
G2DvzHPvxq7eELh8sDkaCYTVLxno2Owzx46ZVnkg+bA8MRod8o+1YR1/ZYngjqsh
JkVy02o2gr9O8/Nwclk9FuBOhE8qjj74VlKbmBasIkbbCh04RceC/ce9b5S/w6IR
UB3LFCGPFyuAWwBTZyAr8OBvFUxu2I+3ukjdr9GKdGoGmccjENbpe552M3o8Z9i3
vWhnkx/LYFiRPabOchXzpUn9ZZxLG6+wjCSY4yg4AzImI7hvb9bkAVpHbDIgeWx3
z+9NdvNrN0a8JCz2mTmTH8LjOSU6aQ+0StLa0TrP5nzXk1m4NE+F2wCMHXBHD2uC
9EyDvvRr3O43nyc9QWtA+yOVyJH4hcjuGF0WLZJqeuQP8M39IHW22CROHKi54HgH
g2m9UtWEyN1n0FfY4uyAjFSOiDaplOBZw0ObX3d2MlRRlhKa8CKx5l0EVjg7GpwS
1Wo1hZeoFHDT02Nd48MNIOxr/Rpa0iYRHfl4AXz+6X/c9KYW3LFtq+TmE2/FOsRM
kTc/Q6RNmkTFiZOHkT2w8kbOrckuJD/w5U/2DYkm/kwWwCD6S2j0Vur/w7rtbxKM
rzbaaDeFVkNgBw5STUcEE0okzz0oF02TDiJGv7VkO1IHuk8Np0/YV1z1AGCX3EFx
TWcYgm5fVeoq8CbptjuKcyn8G3oFWoLbH+WrPSpI2TqVAy4IsrhuPOJoU3I3FDkJ
RVjSbIDL9wOfO0sT5xh9TBH9qzWtPUliv8Ma9PnMPoyFWeTZpyvrmYKMXetpcPem
+OHxDvT1j0icLJw8nyiNDLiewvPaZeiTR2FmN76qJxiFoU35Y68N45YbM5DhzR+W
56HkXkHHgBNKHNYwA8kAP8zf7eKLtl+iVb4VglFOyKoiKRqagcGoVb3PNzpjpVUk
KlhmGx9o72iDq8/fl0rRIf69ps4/AyxojHC/betlhucgRXrcqTG+iUBShvd98BSa
6viCEoL6NAcMELsJ3PKUwFU830JoFOU6riLlYu7wA1rO3VIAubBg0tsI5nQK2Z/n
zgR59CWqJvRbFtkuo/3rnktjlJqZU7zE7FjuCKdRwhQQ25Zp66f2yxsc/XF/dVye
SlWg25yxSVTuYFU8IrInG+w5mBwTWXdBt4Bwzx+yZ6UC3UqgmtEA0zv4FFD3MPDp
Ldj5Eu0T50OY8ARVyScKyxOOs1J2O51Ex5Bdj/FNDtjZ6l6KGL4/fR8rtd8lDIrf
bRqsx8FpRbTooFmZM7LOioYXznlczMTwl+Wws8FVwcky2Bl22RISd1IiE0yP4sqW
coZBMj5epW/ZVfUefjZxJiS0Q4fKUx3ecAIbYEchYrpUqxdhxF0ST4GvEusrSxfl
ZVKsBipy1DmN09USF8kKKvenMPwhXhNIDeIHN6Xhb9kiB8l4+x9ejDMdlu2UK+dA
ykV/vQV7nNeGnV7aEehXBt+glTezBKqL57RbxVD7t47uUz6Z3tyJacTN9KFs0gyC
y0NGKyYkTjXqXFMG7ttNoJyV9PhXrMzHFYfHHi2M6SOxudON6CTDi6VtGWUZ9WlT
1tX+6CMkYG2iIXrH5ykx4KBXH90avCTCpV2WY3ZM1VtWR1zj4M09Wpco4K+saorT
jBlck5fColHkd+V2yy099/qfA7KU7PY5jp1Efqv59c3nYrO/Sf/OHcKW0fPdI69s
WJlxIFkT/fh166PEdj8KJpJsrH4MTakbvFl3FJ3Ex4qeLmfW77+CDgcz93ww0Pay
SxHRZxr6/W7s16ls2vj9p1kRe3txzXwkfj2YwQ1qHcxgJMdzMVuqxlcTE+t9X4I7
u3hxj7bMeY1EJ2HZn3RNqD242HUXn/TBfEdzMg4rc1KfpZjMoroNzHya7frbzwFT
TqKGw1a8n9ydpGzT/sFOX9brdreMeZseWoOj6YVIBDJ6T6/2RMtgWevUsiaG9Xrr
LujV4xm32tM+A7Q3jInydZDgPw6Qz2HRfld2w/wk/1Yu/GkR3Egbw/8hsQVJRAhZ
luH5Rzx9aE4bsSbLMu3yqpMQxKfdLqhXPjTBfU/Z9zEBnny8LkrW27olyzwsM2O+
LH24VYrgWZ/hCMqbfrHaZaA3cgcmlmHK/H0IYKYCLdCI08pg1Tfijm7c1wOcLR0T
8/e4S3NYPfLX8Y8ffPrW/DtsggJ6sNF72oxgN5+/OxmzAtjoTSBkr7moQbNRwPVI
2Kr976JAPBRuJ4sLTQXvUwMIKzq5BjRVQUB3xS3Aog6ZcIbJbx6ryhjLQkuhTJug
bbmvvJ5VtW/mfzlEseT79D505vnrMUUBlo0SpaW9mcmETKMag9u9PsYu3Fo6P+Pc
ZAYH7jOplMpqc/z8OTJfRWdcUEoVM0lOynDF7DJ5CvSTAht0En9IX3fBAP/K2zG9
LPYFSVt625Ge3qhMOYN+fkAMLDBANasiJG0/1ezeHI+rT+Ymg+2S3ukmxzJoNJEj
P8QfopC6zTu27/jJcWTJFxlcOB582y0fy8RGtWl6Wk/IXg2pr6PAuO3/H1LpC6Mh
TPcYh2OdnwkhmMy093WEwa8mzrGsHKZszAJRDHa17rAP2lPSNw5dD0AqTcfqgD7m
2gibaBZjuGUsSuWzFqYNqJx3ZdGSp+6McPTz/AO5akv+wy9cWt+smbBJbtv4TEz3
YL++HC8A6MJP2dFeDVGZgo8KIm5Kq+MIwNruoBEWdzXXAY1ThmF6OM6nJXDo5Nyw
qSKebHwuMQ/Vq7oWH2U4lJ/oR3Ic8nmXASytA1TAg7PQgIHEBAJNNFtFYRNwQkHX
mFZC6QDgZ1Dom2z7zlyAXqM9b2HhUvBgs9joVhETWsjgaS5iKoWEnbKF7NwFmsYk
uQVU42wIZLb3io8/PCGotHsfgcuPFyqjGgp7z4xcl613EkCT/uENNJVnu0MW6hkN
pIX7+TcKiK15akvJP2Yhr3V1Fwp9nndTJuQfq/D5ggSfJFGiHgVOwgGc8qXjxTlH
vb+eCUM6qdmo0JgPKpIs/TNrrw/wt40ENIaQzxuhj8RQInczhtFfN0tQHtwdIDkz
nn1m0Mv7lRKEuucYN2ubTeig3xIsZ6G5g9OZ9o1PIFonEp/5fiA8k/6ecBjXXmeX
wmUFmIRnDexeS+o8zEVicv4302uG8T4MGLvEzzczXYG1jxKR8nGFlznvqpTavBwO
TRQdk9H2//zKWv617jZTdxuquKGEYbmKeVoEYEdxp6OIhMYoBbtrhsOhKxr6nehd
0Pqrpj0G5WPAkVQjphgaLz1wP1wpWKu/XB7IuL+9X7WnGHaaiUEsQBGGnvsq9ycC
lB8jL0btahMIN/RH4nZ066Ev1pycJEN/QhvZ344wRkcKOviq0oIpy6ppKE8bKygS
DC2TtJcttt3BaBb6BDUzZaSRWijfocuK3cbY3aqrDuN7sQA5bAqep8BNjiUdgLN7
E/Sq861jMCF6crfZKGiSneWCdL1oZgAm/zn6Tp7HVj+KxnFisF8f1EWqDwZmihft
U80p1lGgWELEB2NcF/XSNypivVGVSmooVIna5/geO//H0xfCHPulL4oLdAL1ZsWA
jhXQNU23znz4nRRASkts5vuYFLHYcWHCGHXqbeGntgSGx7asOU0NRrfTif/M75fj
X3IfVww6sYZFHkOLucwTb3NNkBHMnKeBFd8Nn0/1vGZaQwRNU5DPharHLkxj6M+U
FUX4us2VsCeToQ5pD2XaYCSkUYL6zJokLgsGCVB/ZdxdPrB3t//b6ADKRJPl8aOm
Pctg4jKMOY9LHvEUlEIoJQy2FomwbD/OKXgNJb+yMNRyj/kzLGk7r9AuVQ0W/vHI
txsecqDUXuUDXH0oj3GU0uki2bC5VUbfY4wBu1DVXOCvQxN3mJbLoiS4EzWl3Xuq
8YelRa0wzXHiEWZx3PmXtzMxUzXR6bLFATnUwYVAl8T90++8fR61dkXAvNns2Cd9
xHmAlPLpItaVFOfJ/6q68nIvf9kBz6/KuuoU0sPkmsSPxY+3Bs4PSc1asyaDZ6lY
2G4z6MZNvEa+8cs9+pGIVYr4fEfgv9coKclH1lSZTF6MohwXyGFqkjQMbOksPqwZ
widQTmUFsor2pX8I5r0gu61m39yXxsqA4sOswZcdm7+gszKEVE0affotHJ8g7R5Y
Y9BfvRgD6ZRH1jL3Yw1H1SVR26Sf9jA4mckFwCPkpvXb1fyVSj+Tj0Ec4vA52Axj
FASPSkF9p3lsH9gFEXtKhnKlpXoC/6rOIT+omSXD9NVlAH6Nr8epKk+ejCV3kRp1
XQeXcXIYzYZCUkYaEK8nh05CSZEI6ZZQ/JInA2/uj0ZAWDlVKr43Vw4U8C+EQnzF
d4CQHDTEaoMoRYcKAARqwFWPm7lErMdo/Cefx2eIPGD4KwiucJw/M2iD/5ECnXgW
S6BJPt0tnux0ERYwrxwaIKU2fUsIyq4NeV9/PSKjCPa/Ou5Pa9MB6NLSV36aWI29
VmnHfz2FVevfljPG9MNyxoSn8JuEo1IJePquAUwxEkjvR91+wHy4CgnFT2Gozlcn
gzTkOCntwvX8N0HxQzZyN+DgKQa5WQNanxwM81CnXGJ5xDscu2d9+fg60eaYEuKi
UMGEQsQ0eLWNh0+8JhIOtsFKu2ujQdDWTWYC2Dt4C6R5EwfsLs2xLpXLjyjgfrsb
2t3GRopZaQebMwqsnC0X9Ck0IK+hHPXQrRgO2B5AHHzGVnafHO+Ttnm5k9ATnO9+
V5uGRX8fvwLagmPJp/3O7R5sS2d/qzTRgf1SwhlCizm4bvkI0RcUtOrvFqbfD4qJ
kgvzwMNM4LNENgO+D/yLh6upBpU1A9AdWbVeR2G4aFv4Ar+oBt1wsmUgHcsE/U8c
v3fWsJtkNW6Rc++MxmKnDyzHWB4rfyzM4pPcMBfHQz6vtj0l+ayGzZ1CZ6CfeGR+
yxT3ulNr62ALOSyKRxkJafx18Sb4jrfYt0GDI4cV3Q7uYbxmSL5dsWmEOTmHGXo0
DNhVvuiHqZ+swV8la9DMcriMFQYcLWIbeKzqqMIpSiJF9FCnKvuRE1tFm66eN0MU
I+D5CKbKKQgxcWMYjwejpnjjuAuMwZJ13rmcyAPWKekB33eni7hcnBCARKfEbB+i
+PsCWYuU/i033bMJuscsJ2fTAcL8VCiO2WZ4kA5f4kxvMI0FAIKbQ+KkIpsEQWLY
quIjJzxvmGZljV7c+9Dj2I0rIZHIQGP1e2MbzkMynPHrE/Zn+hVZO4c4NdsSbd8X
4UGInP/yIqfprhhIvqj2tLHxKPmJeEXAuYGKzyDDm+gbcBuxqRxO27k02xSYBHNT
4GXtm9Z6Pc/PleStQpBmcdOdiGY4WnYHgcpDRyWxI5moaIBTORIr2M6jiE9lSQrO
YzjChD7H41blbrdqDhTSQcXXM0dcz9LeS2e6u0phJRcpwlzuXu2q0Q3/WtwdOp/T
BuZ6MPZbi/SPQ28z6wCPKPcrx343xfI+zM/fGzVchO5tA6DW1o6XZELy5ekoVyTG
Eu+347DrfbVEgHqA2athfyoyc3SRY2L4RFMaIvelosnBqowj2TmEp9TD3/hRjqhy
eD24TXgOGs2wuNlF75idpW8s4fNuxFaZw3Ob2FSjwWmnQjhr6n3WrwqKnxXSBNHB
QKBkVq4wRdzC46w2gMDI5nqskt1NQg1uHi/QmxwelZpOfqGKSdJmY63MTEA8/yaq
stdSSfLkM9LrOvJCPvWd+jAm8DLHBPdNn6V+SN2naiLI65wpuLcs1ukeq4xwPV3E
Kux/zcY7Cc30gNqmFd3GP+3ldJys8rmp6TXfSUy9wmvRl+03VahlglFzuyzZep6C
3+qf9cbzPduDpQXHyrovgb3/uCVSfB9gNICl7NlWRPk3GDDk9dSYuMXczjQ5nH+t
dcLSNJkkyF0VOdlPw9x+Cn2zaFBdXTeW1rG3fI/9o9NyUyjE3IHMANQa4p2F3Ul1
vG9SqJwIi5UmzyCMeCfyIfA0sWqQ4/+D+oXikqlD3aRWGJLJ+wGXGGdKzGa7lT5h
1gmGFz8vFb0Q0mgZA2J0mSUqWR+PzPc+JzfOoqCXpXEACy3Ph92ua8ehAgZrxKEz
lTFZlEjuoJvnoUNXAfnMfpqxfXHW39vS0NngQfsdbaEcjo7bmo2Vkjwa64gnN2wo
0yl66viUWpOi3zdo3h1GRaecCiuFpyBI8rE6FqZPAWyitn3i5thV0B1vW2S0K64a
SQYQICTzwdW+S5uSeE3nlzFCo7U0JFIqNgrRDZI2Y3F74IQFaYrVLES5J7e+EqeF
X1QXRlM1WwGjbt4lKXWerGUWlTvHwla2HdfNU6Mn6zJ9hZvDMwv16sF5dUnB3R4e
wei1VzAVxbLgzJPdu9qp1S54THW6PkJnmkaTtisEV0hWVVyjXPB+oEPhS+n3bw5n
zQ23K1j12OJ2o39Q5lPXPLgEC/XhpdM9ww2KVvxzJQ+BiqWTYyJk7efWoyom0D9s
xSPLNwGzqgvXD7QsJkL8GpOpgZq/MFrV20xQVzMJOkBlEZkxzSlSVwnzMeinSLwk
I9zbH+LymNTB9Lv8aUCdFJmNJDWdX0xcB3EVQ35GoIhND2mbLzgBPZNZYTy2q7f+
4SSY5aR3x7pkr25BdL9N0h+aB1uM8HeQN/V+0COJr1uA2sscV/F2zKDo5MJ0blUX
0GjykqEBqbJi8ov2qUax0WB3JvKJswzGup6LHHxObdCGsk9D9GFnStjq4YLLxzwt
kZB4hjqEGt4cLGIf7uTqhaYNN2bWnAgpwNyhpbom7hlPHSzLspm5MC6T8UJl1Htq
VcuQ7VCRAc1+eYe0qILQsZ3XXeqEyA1lYabZja1Z1uBiKiW6QYRPKCxZhH2IdNat
yjwUjPcrdheUrsz0nL8/Zpyl59P+/BmKcEJBW88SpvK6sfsfKmLs9lGNzO3AHIJT
ePeBrrIynKuN1981NTc0nq3Qd3M++N6UV4qmfwhSMlQsE/VuQYdV0ZDVHwU79+EF
OZH8xCRpTqB+uoAqYmhtJUHSmOaTk0NBB0QNcbWnzFOl6yz/BxFWQvmRwJFOZP41
IYuR5FAl8MablB3vHnjqey/d4Ebiu9WcLSiFq2IbNJZfQb4TQsCFVMeV7rJMFMag
8IoVpMmJFXR/K3PB/okwOWDeaCjLgHlPFRytrBNCQIAIf3lpXoWhm9w2tjn5Zp8N
TPKhd9ygE58OwotKF2GDmJFPkBnIhPOpM0C0m3A9ndTilrdEkudcE0+S8PR8V22n
HbpRhvNp1Ejb0RW9FT+i0K7JrND8rKFY06toaFbzrpi2r4wuDTs6zS/cHJa35CAp
4l/TqLQxbFMjvSYS/gyqPHHgrX6aRFBpIng4YNT+bouMT23lLLONmkFx6nMj3cFO
OhYPJNFQsXMtjW3QTq735yH4SzSmDfX31ogK4XMtSjAdfU0yFqI5zahycE0pZgSF
Dg4shzcUvH43kE4p1lAatIFMNA3WZRsPh0NMk6GxGLth9L3KF57Rb5FkFdDQMRnp
MJIDkTf6e7EbmZ+XeFqlRM68NhVG1KCyAZvYEcfZ6qOMp17mb6UxmYH591Fe0cBr
E7STd36QggQb0BuwTY61tFWdxEyxJQwRx/Q27iC5jXO42sUbnKYko8mYEwX/xQCG
VfuBvAxTDGtBr/vAQGMK8ePJgxdf+44hfTQB5QqG2Cbz9qKZwtVcpVt83m1kUz5O
JAa5jdRNF3uzhm7ODUL8VHSOdViAKbkQ/HuCqARqS45A4gCsKInIMOKIciDn9rpb
hrIXJOBzF7o8UWDuWTYqArtFey8eNAZcDry4ROUWm3qev+HAHXwU04hhmFJ1pc90
QYwiq+bdDJ//Nz54fZt4tBrHMc1kVxPfxBg9UdkKJciHxxkAzT5gV/KmXj9h7240
zxGqc0uP2jIGx5OSDvxuzdHhrNWTxESIlJKE+i2jK9ZGaktRurw6DIZ3Nf/0jcMF
+rVpv35+L6LsyqXOzKpGlKl41opS5KYyBpM37xkJ8unXMcI4kzkSds+TQdo5ZGCX
Nk9y4OMAvMfagaxdpojMcft5KL633/2x28UX+ebzuYugpuaKjd5fJycxMnYi/KoU
DMLwBWsRRCy2qgsthObvOVzhyTxBd1gkus5A2SPLSMI6+AueBDhlinsZfqY7nZ39
v68sZfIUPCuairXeCuT9KGcFfOytOTvEK5cyFAdKo/dDvT/TclfEewJvhcjj3C36
Ecbmnaifl6aP6fcnsbHw7+41Q4tpyQ1Un/a/7nkz7N5trQtx+5q5/jpu/KVAUSEW
RRn/LqZ1tf3CBxH32Q73oT4fYOe3/HNj9dJ8HwbUrIUWKYUsyO4X8V7fYVgXpnsz
C2yRocsd1az3dMbH4f66pTDzb6cIwZgtal32IT8XhZ6hSPeNMS1brgUICMdy3mqy
u8v/9NIWJjUoXv8HIGZ4P2EiJtnE++7bFJf//jZobIzdMfULgAa3IpDoVcEVeBZF
WgnQFleKuZE+jLfUJ8I098nD8UgPII0ltQGIxCKRAeVs465uBH1axwZ3pNPYmw+P
q5X8yWoJKffyx+GmU9ww0Z4LbD9FoLZQuXFI+rdATDXLDnZ2uMJwRfhLD2yv2Giw
Ip1SbYfR96Pjk0op7kxLOYc7cRRapcJMsjKL5xUsS/w3K2UKRg1kWGtLjGOAc1r2
WW/mk4p3Gs7hZbgV6U29M/knP+ctVg/FWsido5LiTRjs/0YNt6QIFgenc+eP1jgJ
AA1b/T6yQTBeM7nda6fBkxw6szp+kDWC0gT6qfLosL3vJs6KeUvF+Nq0C47KDcaH
4xzfbHURLbnlsDhzLrIlqL27G4/UNIfBJmYSLmQ7tCZ5oneRK+oD0Cdb/7o4W0c/
Hzjv8NHF27wqsDqiTBEaDepSqHYtPEIMxvveqffQssGYrVCO/+mICi9MiTwMSgqB
ykI00KF8rNxXM7GlhTwuoJxq/JOqHtiUVhBMqi3fKaliB5/zjVnf12omN6bPf8VZ
bVPHUm5VY3XeOBNVvpSwJfL8/o0FThfgRFWwzJaR80ajo6S5ZdOhVx15ugboV9+K
ZAPTM2+a1OfSOcC7B+ethqSUn4tDv7gaOSCIIWV70y2GcjvRV+fxKOvNu46yoWBg
Be1K2RaTfiFqPHZygNfAh+E1z+enyXkKXGAmueXIEOqjd/CqsKSHlWGYGJG8TXBu
hX7uLwgJrNnYPGJCLXkcE9CkNzpG40qZIGBa/N16qRSfCsEkUi1lK0XYs3+PtbFv
+RIGtoegfPdDe6hZWS0ZKec7ro5WF0/Y2Z9R4IjGaRgXizL5/YF64sP30kKtVCRp
5XVS8cC+PHaryT7NpsAWAx3g5XHkES+J3Uy0mF9lj/XPwkA/fEVFCWTPOl+D6/N1
5tO3aX2excN5+IrD64XiouRPVBJVABixL3JducFTps3Yya641GUa9HDkyBALM6Sc
4z81rgsXjN93b6tM6cmroBf6bgrEi/FtLGmeW2RPUB413u7Tl/okVu1bRsZaJptf
AsmdyUY/s8w7/sI5NBynoq7drSUFN3IEhXiDrudA6dQUauthek23KseL2cHSzIP8
Q91OIY4W9ZrA9JPUeGZvvr6EWbgSsfhIBMXoIgY+GVcFigpMFC+MvMb0gAbSl4E2
0pp2OMyJXO/T167mieayN2bBrCoO+E1JwC7vcsqrbG9bsVZvYgqRoqZm5L4E78Ce
O7PvbNeM8KRU/Bs9kGHjDjjs6SY7ydgZATK7md+edtd88o6U06KdsR7oYZsTi6pP
g5R8qrvMpa/iofK/Et9FNFd0hJs2ge8+h79FVti6iiNGjeUYAjeqHR8lbIN9Nvui
8mAg1/F+4rKB5IVE0qRspbG32zFQCZwsAED3mXkJQgt6ch5OLbNvnK1bTuwFkZdz
/+U8cJ3kdErTcLyozi97lmlOST7ixBw0qwfNdbA9tC/9dmSL7izIod7sMmJ/NrBJ
g8PEPeJEcIdrfIxF3M4n3LynHUlNRbsynK9GoveUeFheN2PQV76vp0TaKRwJNFxl
AGl58IzD3fh+EZkYhlMKI/jUUVwuS2z/cuSAtmRDIhZSuYnEzpx4dyQPB1yQT+DS
DlAcYiA5eL3wFTv63elApPSJy+Zqx0HmHMoa68N+WyoyKSGlnNTnWwdll6Gb1jpl
r5gdTLiXvZCyLFWZrWa725xPyk/KnJDP427wwYvHGf7xtrM8/Dzhds6L1fnMdz3X
coYTwEO/I6AISto9nbjC2b74svjXMtGFpKFfOvNeAzWakZ0d/VxxfKVXyLdfmmZx
8U5WnwzfLyWVIj132CoCIotRz8vhQ76yEAwYEiI+cE78c0WryoOj+H3pIPXswfS3
aZvhKR1W/pJy7C+XTIY+mJm/tbiAnTNclV/m29BSa/HlOFRPDZJNSjP2PZrSqANn
S+zYF7mM9pLO6bfhi/H70LZ7goApZ8JC/S8z2DiU+R4KUDPfWUZOlKmng9UM9s8F
kgcmyB5ZpXO+1kmNFXroBp9jvs8jEgLrzRBJS3HbEJtKP3WMdjskCCnBhXRnq5Oh
d/w/Z2BfrYAAtfiE+F79vABwxEEbwlVP1hrd2DvDaN23sQpJ843dvgIGz0B9I9Dy
B7Ei2nlwMZ/GMkbDtLTyA2OFwuH0YZosN3bsieU0XWdsQbBAmn+caB1U9YxEu9JL
45Lx3beTHVJd1mOr4gl7f/c35Hj0dONb+Uv0AY2TiSzlm35qPVs0OV24zAtF+E8A
PFKgaKCF97/f9GyUnOQ35ksxmxOAC91XHudu9wtK2dkeDCXZYLFPm5HPWI52Z3OQ
Smq5yk3Pdztte8eoRtC/WxUlw3NvbHm4r+A5CtzatTBNUWL/endRCELWre/Bd039
lq+YtiHSeNr51u9Kv26Zpj3OyHa8s5sFqc39+x8P3rErt8TLkQnYswZgmHy+H/0o
IHK5jL7elY5anEUSaimxIm7NDGp51ALwbmC1mF6eZnJ2nImYlBh6CUCFLdYu2QLQ
TqQv3Cbn9pn1/jzbwGcz2+dWIJTRlcDyqQERA1szPm4IL7wVARJzISFKevajo+yK
WHoud8l2SXzt8SqGu1u8jw2L/ZQlGu3gpkU2hSHT2teMG1GAgfrjDIh27+/Kjt3d
X+knnc5YPTFyJIiUVr//5qWo5HylvDcvXBnQjezlqMoaYFkeGmVcGDs6HbwxWjcZ
eASC9OiuUvO4KiX7azqoIPCdA78iLE9FfmYFVhFN4vJJpP8E3hQYIPhCdOlpmSiT
czYmYGzQGx8bJk9lBLIgDyKzzVC5Fh7x/Qyn1yHh0Vc6uIPTX+jGM8bCj3NFof+Z
jFnKWW4xo1FStQbU5QZwZJPdSUOgjCmnlcj1Pofs6uc82Hiw1Vbssh2r2uZ4MLry
e3FC/IYLXvOZF+/zFwQ9z3FrOUK30c5FDKTgTcpFzX8v+rO8tCRhvXhHAMUqYWKi
D34l7LpRHd3gjH6br1go97/LF0KKe2DRhkDGi/ziI4tJuvlRMu+AvIHchlQbcAXy
Ih/OzcJGomVDUV8nOB8vwiSvy6tClVKb5In0457Ar58imhPAj0q2JM0a0Sm/nsXD
Bg9k6TzBiR+6Q0roV4ueElE+UJ9QTofRMqd7I9n/PBqFrBbaOTrwUwSmLddTtPk+
ftHPhc6D20dT8KBBhwWbG5qanSXcviezlvBfyopEZ4nw3zStJnogchkd7wK6jYG1
HNyD1Tgm8Jk1r2FSZesjY96kwfCXT9dgOckOJJEyQt0Fpy5Hb2fNudBhdRts0SGR
hs2v6lHk9z4WY8j6GZdFJM6KLu97nRkv4pSD2d2sPQMj8q6U89rEPH4ozVl2MOLA
Ug8o4M4btxeieD6g+ONR2565aBGqHEEbC3GOy3/GTlKUwYodnXv5aPbKwT3US1k8
3yBBugy6ekLI5WbjrwESElSVVh4uoEnFp3mWktxf3EmzTwYR8c+9ZfL8+XZWj7iA
x6UluAOyJro3JQaWILl9JAy/BhNrytUVNsQvcRM4bkAk5ZiA4WkkKbAznW9vXNyb
3o4FnJB8FZrAg9/QGzVs/8s1LmlAJEpKXp0HrfdcR4yELOcZmkz3b4ydi5Ngj1QC
W+Lv9+Q8/kXwHt4eFsDjZZnZqZAOynJnI8sDqLQlS8x6rrhDOgUXj42w2+5414xH
/KX+Z6ajOUaCV+CpLqAH3ht6qyZtBfURHfl6WV6G5Ep76VA/Y2neUoxzFlK5POfM
vyghPRiGnCwGk/TRzfjpa5NhJg8zdbAnsAboJ2AkCEo4sPWXEZqjJ0vFcdw6+/bj
F+oyUhZW22Xf+ZtDktONFk3kYZ5Fp9Ztq1RzlRuPsGzVaI95f0qhi+9JYOyMZnbO
sg1yhQi6X//Aj6EEZS64zeRkjJ3q7IadT+g+gL+vrK4haZ99FDCgnHK3/BzOKeDV
njtl+NK5TfQkgaLmVDesKPzBvU/6qN3tysxM8+ItG4EXS1g6mp6yfl3v3Xy4BmrA
b0E7g9GR2dJLzK3t5hZ+Qs8qX2rJ1vZULvSt3+Flw4GAL0+2xVzLYTyAbY+tN+pv
3HU7iGrBJSdxgWyzstIH9dW62B+tTjUwUFGUHhgPLG/YbEyw8i06kRDV2X4ohf9/
KgzW8OGJcTYKBrMR+ez/LfT0XyDh+S5o+o/iWbkvqyS66Jm/tW60Razy91Kmwduw
RIJD9U5eyrmaZDSESQH6sVNe+IDFRIP0tdHA6vpJOdktHrCJjBSk+1+rkDxmHYEl
SURFLwBsr4tHlvLmQA+xiWeRxFMSkm341xLiYLcww+AmyLy6/g1pl0SxSnWxKYL/
PQqzR07K/OYPsxP3/yEhbRBQ9gt1+2DTWlObp14KrpJJiMe0mR1oF115FI/jId4o
S7SmJ4XFkLNjz5QAE0WnLJhFgonHX4q6pVygpt8DKth/mKn4z+r+mUFvWN3dS9PV
lY7j3EpC6J4efvKPz+J8VHg08EuNxO0aQ352Ex7qO1ZNVfuNIokXTRLEWeaBVwjT
MJd7/bGxmzWCtFiGGdwH1FQL0qHJAbEs/qo3nFHcfBPJekBXP0zqAEdtvRRMPNNq
nI5iqRsuUl760LqrvM21U6fPVeDjsbUko9r8XyB/Zoac5AJpkOY1AINF6FawfGiS
QlEJcBIARyabZpnmtllOk+Eblke7iaRNtb6UOXoLnOat/dv9jQt7hGWDfT4ctBsY
/p97dOnCtexpsE1XXGLJxKbQY6X0uq/4vnbGC/GJNN3QjGzQihum6007SWMKoea8
zbGdZc42zh13FBHzl0OlaqaaB2Po1Zy4vYii46YWoG7Sdz1vAVrJ59v8zxedqrVm
aM2pJ4DcMUiHx4hSBRdjteVfyQgHq6pIYDJBsWlckk3H9wywKm/ENm0rXUW7rJsR
1ze4cQJHs/YGP4lD69J6JL3qtWf/Vw/ClEdh59cUdmDQBNjKGrD5kfTSogOnsLjb
cViMYY2jP3ENVpYXv9Pj04TaCdRk+0d2NbJCQ2g3wijNWzEtnoZ4jg61cQzVJo2O
meHYnaA7s09I5V35+sUU/yiMAV0bPpAFvOQnvUfGNRngvbUkzI+ftry6XS11GKmg
F2yoQen1AMxbRadc+VGUd/rxwaYFUbz+4q5hihGWP61Jxii3GeBr7sYDPTbL21wF
EpkzOL31f5DgwR9Z+It/Gx48+M8aJIba23nrgmbpBVSuldp9CqJmndEtdcpHtiI+
Oq3oE8bm+8BpzTj+RLS29vkGaxLwnP3Rfn03zDlolDoaulWgrJGDnAExM/bGxPdw
DUVp2FJhWRlSe3yfBgeVmoRtcTbahxY3LdTiUvD2rFL+/nd/qGa8IHGeUwBChl0x
pbdzxNVMkzPbbFFVFuxYUm8+NJQX7DEBsuU5E+IdTK4yufNR3utwpGRBZA0i2nc8
eS30o5TMEy1ZXilLAKgp1ajqHkSfOZwN7aNNOokxPQlByC6wcxi39vThFKwWMJam
HesJ18XwphltPzTjKct5e+3dfqZhhSYaBvgtz3sU/2FXXrV/u+liu3+dyo2P9yhc
0S7SvEEquMB+E8v2hBGAyHgFSAyxCxw4dV7FjfTQGkvKwIYDm01d9s6AByd973DP
cQ7WPS5eVzuhqFX49CFd8oyGPw24219aLRnyWhr2ijuT7PgFFAJaKsCbFXiMBr9s
AP0NR5q/BMXgGmbV4iSLsFwHENNMruC0n3YqiTKxCmDXIaKYMUxEFA+EtRrGlJNY
smewBxhJM6df9jLbTWl3kVrmH4cZnAbWaSP9pjeW790tu0aYzEO3WSUCu/hj2jW2
2zFyUDXd1NKSUYlLs9h39AHG86Ct9pbH4g/gcwmqOapWmwZAHhDnZMBi5Fq3BanE
29ljbw/Webfoj/+iwIVw3hd+66I9yQzzvnyS5JOe+C1QRB194loFI/m0A2OsZ4Ts
W+PRi6YzrEWQviMmmb9A9u/MPxE+dyAYyzTVAZureFia+Ph0kJ5ied6syYm2RRIn
HwIWJbNPSW1QAD5nPBia8vxx1T4wgRZDLRrSCtTZpvrrRHCytUhMt+VkMe+XL7oW
ow31BJJkHpqCenv1oEaFeagto0KVzdgOJU7lF92qBjF3QvsoHTQ7lo5Lz3bxHK8f
xGc6vAt8etWFwdfeKQmpt8UUjOAnGDZhIR5k8z4BfW3uKSVOhedht+CF03HAdjcA
nI9Yp/ce1lXXvsRwnmZ7+YQV52jncs0T64XTlHS0EyKh9if9MUNWuWnFFJmUqxSl
SZYJ0RfcA2tvrQswoO/YtH8Q4cBRnw+XlCvlPZ4fA8wRRWJZlEJiMvlL0EP/iiQO
gMXGdqyvPzOpyCwXg0tBfpeYC9B6MRGaMW8s9rTozNaP7kHpiLiGjvcCR3eWj99z
hPVHMwwOnvZ7Tk461OBLAFQqriOf1Ld3VuYkh+K8ZSrnpXGUCAW/qF7Mxmg1+8hc
SMvBXFF2bo9XDZGnHJ143s9/rj8b3dA+GCLqjhHwaJwAFbFXcd4eei7dNuBp8jIB
koeiYazvc/BqFI0Pz4N0eE5ashC7EkSLU640xxCtbHuDvBfTTTN1SoW4xi5xDBJ3
sgwbBTKLYVnRyT1h5uyO4Rl+n1qG2h87Qkg13sObzk5D+XCx3AU/WRKK79NAsvAo
634sfbbGbBqhdGCT1B2FTrO/RfIGKMpkAODe5AKrj+sZVoqsLYHysDumRHILP+gi
FpL3QjQQg3zVaSwkHFUrcwAJwk/PvreufHKnImQphs2TqQ8vgzvqhfcYJB0IzBVH
schSdm0+N3FVnsiVle24zjnqDrNblB8iBGR2XtMp9j0ekvRWSNhi6JBysW81/lXl
pGNlv4H01FnvN3J7x1n8cmvnMAOUMUzR2/D1sv314gKnZLe1ytlUzj7zf9DgfzzE
rMiNyGd48CZRmkjaUFoeYpdIQMReEV7hviEC+4maStVBHFE+rGL0uJmZdzj/nqlC
4HvLK/lfBGG1qE8MqEbmrxk7e1lb9aoR9/bplTEclTigg79ShXa7HmqvSqeti7lr
e1n0ixrGGE5N1rVionsbmQHdaZHFNNI4jBv/NtNOcae0FmBz23T3gtoGA1CiRsm8
ysub7xejreAwSYcKjQRFC/j//jj3ElfS68U3TpPAlGiVOOLiYiYMEbkzKqFSVv7n
1ZaH9SuI2F4SStcak5rHwJeCJ0/bECNjk4OnUV4Ubxsq8F7CNyu2HTbrF+MyIh1L
QLiRrYTPLytxKp4kvIWPrm4fVdGKKfc9eeABi2bhAz8wUO2pK/ddg57ZPT4R+KyZ
zExa/rDNOEEubY3ON+7ICfboO38rABzZl3eoK0XaqAMF57Gvz1OWPVzrhosQ79uh
tmR3ScTyqt3sZLFH5RVRhAB/OyJOup6b6EvFvX9xGaTR2wNH2/9DmCUe5yvVq9G0
QbWrEzVn0CKjMtXVkeMri2OH3+tJhHDrlcigLWslyidvkdCBXvKqDZWGMhepLG8q
4lodUlgRHup/h+MgLNr4GTo+evits1S11zARdjrUUxmvLu6udhKthBbvcfsRA2TN
o/OxpgdbQOkrQ0mX5Rgl+5VzOf53RTR3W3byAtcaBXrlZhcIBXcSVvY++eGXeEKW
4rmr8bKijTMo6r20rtCOpPKvO4Lyb/EvZ/y4wB5daSemsOQOas+77eZC5u0Gru6B
OLEPxYWYVJ2Qw5wkAJagpOxaUl2evZ1NpBcWXr6FyEK08HX8f94MKiKu4DnQco9j
exW9wj97KDFZNEi7kPaCJ8AIJaLjnhJQVPw/dk6/YGVq+3CIAXn2HVixQ2CSsvtN
ZMvPTaZ37pwliGsduDkbQgLYGbEwpUMDDY6lv/0T3Vl8GddIvfysCDa37Eu8HAmB
3AFTJGCAZ0VnLChlUDyzfAoIPtPs5gZjJJfMugUXgrj/0FTqbwn6NXZowiA09Gz7
NtkuuHprWldhCf0lTXaI2QDc9cZ2nEBWKVtWwygf7OPX+T08/5jilUAsoL0kG2+P
FxVyEOgFMPA9DUVrY3UoAG4OokwBDQMx/sLLaloplpaBXnu1zYr1zG6AoPuJshrH
w4konqucuRtRZv8eWBpHMvX/PHFfnrSDfsnuAVWp978r71PvkLgodnD8yLlEbVb9
RhBWVqv8lQBTrz1/lnukHaAz7U7JMxmS/wq5lkvxiUQ279tjuVE2xnB+o1Kmr7qN
Z7WeV9wrDBVovmAEAP+nZPhvOy9YXygFo/VEjA463iqX0dmKXm3O5stTJM5JLapl
UpLhko4e0foBhC8mGFf1tzPvgjleZSn9uR7EeFYW33uH457fKquSJ6lE6szPn90I
/bzwxvMEaGahMrPG6wUzeWv0Qbh8ue57u5FcrHiGRgi6n621uuNBEG6rWE8Y2q7O
aVcE0wWbeSQT7t36r4IQ3EOzONKfZqiS14BwA3YCxGQ5/w7WbxWEgH87BdBqgWHT
6blsrpx76+uxheLjcLwuI09JzqrRB1enk3lyKlwhxsMC4Zr41c4WO5iD9FcDofdQ
+leM9lhToKav9hHjk/QiifeqXcp2Hg5K7tF/1AIs4yuhH2R0i+aeXWDmEMMnkbRF
1VXw0UzA2PPUeHYwAWHLONfnNhcs1CvtMxw5bbc5nT8MV1Ictz14/AtVUicuCS65
wuWP/7DNL0d6Tgq8nYZaI0maSb85oD9ZnSaNmURRjselrzZk4IcmpULjc+o37kpm
SJVNnINeG5TvYD/BqAQ5IdejlTY8AcxJODYCXbzCueLrlrmNOqCHKqXT0onOwZiF
gtUucG5elUx6pvPrvK4SUYQ8ySmXjLIMWxBW7qgy/wS1vFG5W7F4BfUorjZ2pu0Y
M8MTd3a2ilYON8XLpOSGZd+X4X9YzMs02yylM1cRZb89+TF2Ri3Jn3IqEnPrWF9l
NHYkeTSeC0eL9ZOX3wpHsZLxzjOU70yNMKJmEVSu99y8HdrUDhF2hB07+rhN0qho
XvlEjs206FfNMQnkfBpgZZaBnmEXCwsBzgdu6ZXT+UxDPBuOwf9qMApDeqWhZSWH
Gsc9HuT8tHoJ7SVf9x6Xq6GLy0L0k8J4XtdSrrUbZHRX2shkdnbHWYZTt1QndxeF
y22sBiU9qbADkTDUdQe1uM6w81RA2kq1lrA/Y1sJLNTXoe+TRG9pKvBwHb7knFn4
7v0fKf7F+MOvyc3h2FSJm+A4IibF7ypxfB+uUjscslNcBi1PHAqaXZIjLXAajERf
SmGC4Zr5k/Hs9vQ0CoETrdnanwbsLjssPi62eWP2ghuj5epiqCbXoqQpPEgsNW2b
6caba60RrgycZMfE7+buluhnTrzNS5f87BuaP6naVgr9Axh2uRRenMYSYFqBQ3pD
1V0KO322by2Gg4CE1N5ZABYs6I0HsWVH7yCJCdd6vCx7tK1ITK4LpXO8JU1LQZaN
wzs7kecrSldHhcN3aOdS1pr2sa5aicvxS73bgVPOoUG7D5AAmOQOClXdloLkOdj6
0CRDUZVj30Hc9rX6Zz933+bnGyow0AKbmzNoO3M6RADimcN/hBN5lm3YMXbmaIrE
bM+iiqY+s9AWFTlOIkoLXOFRXwhay8RkL5LTt+tEgw9s+4J/63skcP6TBmHeuWYW
Z7GpGvlmuyHUZAv7rCzQaNGpb8c7ApOd6SHm8b5UPAGUEJnzP1HYMCA8016WXvMj
uA1zOUAZA7WF0aRrHrw6Qn2zVQzkdN6ZmIDYJ/F2icjgWkyzUu1YFsXcko70V0kF
lAcAYldYcAOIMLQMtNhMti0xMT9yUNRix068G6+dRvXVf0frZUi/qd17N2rm2foI
LR4pViD3OfXOY7ka5Kapf/AeWeAW9UvVF0Yp/6OKSlpQNI+bd9v7/bXEko606xK9
yxA7pFuWH1DWet+vd+RcUddDl2xV8uuO8uijpTsHyUzIPjZhHBiNSorFHjlLA5hr
KrZ1MnYPbVj2q459YvCvq/ttN3uZh/OHUiCRpuIe1iCMTeLIrc84AG16dY0XasgO
L+33C15Vfq/5oPijUFBvFBZTFkXgxCr5USKHBnJFxDiiFBW63AQFi85GFCQeRcMn
mx2wq0kWsKCJ9kxqHPfdf+RrtA/+BGgqF4AZLqCmuCAFVHvr/y12xWLRGyo092Na
LLCuyZATxA0ZmDxhfv04hqTlcwepttYQRl8FVfN+3PCaZ+G2PpDZPIdHnRwlb4vC
nTS03MD1vRlsE7BK0kpWg8BC+qaWulLFbE9/WF6lwWdDmCMy3F9cpbmaYXRtTZNh
8jdY0O5e8Ifnq01jQYoJcnMR3dJPNr2cHdfQPVumPg3vg2UZCe1xmlgzxbUMQA9A
yxuxlZHePK3yGVX5C+nahzVuNSK14J3p7ASI6NtODoFgLyTshZ+cHzFxqo67j1M7
S93GXLgRV8FL6TU58UAAZnVrHOM+ltl89bd3Ef6cylpNrMu1SbclR+2wd9ItT66J
BTIhZ/jiEXtG1/evheIsg0IhdgqA1gB5mFONUpEhTTsEQSiBZUPe9Ivi8420NfCm
I1h+RuKWZuEa6scPXBn23rWvkWCKVgWcg/P+WluBj7VgQOGAKW92t4vyhWQiA4Sk
tq1isVYgwwl2nCgnmuM/j3Uvat/fSwfB6F1HPbcrNNMFf5KaHrgoXK3xQRUZj7F1
mO8ZInjvn70PIWRc089cpCFD5KJr4C7qtWlncAnh8C1B0HQgOhdagYWTCt0cCvkQ
sPEYDaLKeizzZmqVqdNPgYSk8IMazC4rQGm/Ci6A88ePZiSX5DdQNQE7tWKxI9Jo
FqfBvrZQQkP+GME8ibJuIydjYwynw7pkJcqMkgeXtXRoPlB9FPU4UNPgFPESH3tz
SSLbByXqTsx+Rcja/7gYFyUNPwDAHbBymbNOc+oGLwZmUTZFero800ypsKr6TTKi
Deh4aoueRpcQYzk+IYSA7YlE6SAtQhgKeIoTCvofq4Zb8TzxR2+jkjkRcPd5PQdj
WTvCgDDP2DK1rDXhGjiKqbIdrZAg8H0DY05iWpuvcHuYnbPT6PDk53nJv5LvlSsR
95lOS7l30fotWYRmNRaVULhlw0814XBy9XSO4bXgSb9Pt2/tLc+RZyfDU+LAx+FG
j3cK/4Dp2LrKNo2QUKFF7SLaQ+KRv/X7miDdgXTQ56siG9tYxGcVSAqDyVf/JtFK
yRK2ULxIe9UBJKo1O/E8unJD+VqopSReidcEh2LHTSW5muI4sED0stxQkf5GZf7Y
P8VXSsSb47kIxDLiPhq7tU0jJwaeCfomUJbDke6jly2WmIJU3VEvtoy5vtY8/HLj
p7alt9rpUwJNA6PUGmM8UWa8w9yE5AnifOHhhIuGNu/w0geSP2C9/Mq0qHk1eDlF
69vhEkEH3XJDr5YQCy2EhglutBgi6pnE54ZUKM5JRHKjV+GU50o0zCb0JTU4eTdC
v7i5hfHRgKnA1FL2fdbDv/mq/pZIBVZZ4J4mlNSYVEeLjP8SRcqHQ28xBuxujaGT
vkVvCSB2a2TLYpMYx10qr6X4aw0fREjWd8KCTAIP8v/ajhczBcfWdIimSozWi1Mb
G0ZJmiJJELHBQBj9/zgUN30c+MUzcIF8VMvfzBcEPL48lzusEWfSbgCnSIKNkhkS
TMxpR0q/Ul+AyFXqFNcQi+rGU/otcrvvFy2wOa7sE+8nCJ4OMHkUqBh5q4Mvknt9
HkjkzYcvFrchw+vs1qDf/sED22f1e7lnNIsjuF62hOcxLcGwBV4MPodfhno0WBaP
T3Efxy8Wj1RFp7O/v/Ao5Lnb96L2khNfnuXItUPBhemxV9VcGYTrPgBuqU3tZnW2
F9YlSwa2lTpiog/UhtE3nhRdk9LPLIG7xuesNTurb1ivC5XX+IvXL1IwIaPli4TO
hgee/AlSmTConbDJANPURpH+FYG5vlojKOPcZ8+0Iubo3CK3UbsdRnbDBwiTsXJL
ddJ1cl4npkgwxi8YaemyplbyPDf87LdeNkSSdPGyhHF9ZxlM4tHuh5ZDmijgUBFX
fwuSX/F8Gl1d17LpQXm8It+iCsnVGOMZsfwUE5zEcG1DQqwFyEbmuDFKeGXw+Gt4
SPyKe2kkr8310+/e/sHvlq5HCJ4CudhthW969BgLJnO1xKb4lhbfiq/Rur/Ai5Ch
ZpygUqhi7A29JHixNLQZRtgC9uOid6nTv+jK1i/l267BXmjVa4/qiR5dppa0Ar8g
eHWjVdg2HpKpVPD5ijCTtDjOWbxK3eNThmjwo62b929l20iMQAB36xr0r/pugXz5
cE0tNqc9fkT+Yx5wvqvRb2eOwv2Kv4cvV7Rg9BGXeecHzPxOaXKVBTIqb7MZMeDl
g5UWTnaMmGaQrN1jgBgFq4k3OUCacoMHzooCFzxFa6iUia8sFN4P5xNd89BaT+Oz
FMN8VleGHRwjqlgoxlmi5gQ7p0ASDdAmCX/amIztYpR2/+BrrvHIFTgMMDfVbaDt
tdHaHbR4+n2TlXiNOrphhUBGUL7tPfzpDlYcC4YMgg9FrcZj92HFuQ6NJR2FZGMY
iA5inuChQduYtKFpWslWRLDksZPmpUh5VGc7tl7AmoMHVFB1JAmze33jTfSO/pHN
Nkz5mIS4xv0hdDlcb/v20Xnr5xLXTG/1d8fqo1QA9YLxObnK6FgEa2CZ2in+wuO2
rxQ3xZbn6Cttg9+e04RF/fjGWRg8OYjpgRpo4ErXqXbtWR+5jzLfluk/Nq/A6g2q
akRQI6MJwjKaQa5AWAvHs3BLlF8hu4ok6j7VHnj/jKPdZBi9/Ea8lA6wK+zv7YDd
uWU2TIGK6mPP9KURJT1IiiYwrm/3dGBp//XCTDwX3bPpZplt0Ur9eH+GMu+dixf2
iJBwBjjcvDqRd1CELIy9AZycreflGtBt4b5xzyLxvZpe5v4YfgsKqeid4FG9G3OI
m17dkMy8nYhVAICIexIgRCktysBlBQyFZhyD0p0D9wFE32bjQ9+yW2IfI7CwOITL
Yq7knjH6FTrgpe0BTQMruMC65DjLmJFEmCUYUnpuUssyF7W/Xl4UMx0mPJ8kNk23
NlpC7SSM4Ci4CUqE4hcCgxKyAEMzJIamMgiSSGz2kbJLcJ92HlhC1RHcd6Lb+f7e
Qw507DJqiXZMUSf0qE3Vs6vEsbaZJ0ei8brw+ngjqGfiM9kcndoBeu8vL2r8pMnr
LiiHTG1qWU+l4COuIz3kAdtJHEOmd2Io0C8R8gAt9S2vk6FNHFWUTdq1/ItTwO4+
Me0Wufj9ZSlsx52U1Q94bG344mMHLNxsqhoaS46HDMjmhrNIO3WK4/1zMay//2Ah
wcd2EFKPiG/QQCfoHVgbhJpz1tZHv9X99kLsOSxt4o+5mld0NDlexD0fjFtB1IvI
L/IDyJeZe/HQ+zd3uahTGsF5iJmfEb4zckpEaLtuq/PxaDxHegd0cGebiIVUuvDf
iIKxWz55WNtaR5RICGZKHHBxgOeikga3FjBa6nKol+dQAp+nKtZmUjVo/HxyAqkx
JaDJBV49t9Wlnj7arqs449KCwQsnKJPVGe3iUGT8E1VLblMpobANPt1CS0GgkhSC
TWg7M8KjdAn87AfzE1iRM3lUYaFu/WbESLO1T0yH+4a0a9MrQEBlOPwETKPIjOWN
FTRN58DkuXZoIU3HsWEgi1J9gjA4CGjvr1/VfjkNE58KdUKK1NwYdEE6BlgT69Nc
Ej0SLoemCWquIkp7vqMzzfy6XoOP9ZfasgBuR1N0nrO8dcvQYtLS1kCB/Q3TRp0s
uHMeaw87laqErho0rLDFVtxcQYFtzsFtcUgrhNdYcia0LJflDnSB3aD4DHWCHx5O
GqgiNbSLmw5DKCdvIkCHts45fAmukl/2dM2aOThU5d5+8Iy3R5la5uZKJ8ooUk9k
k1zvZqY8mxqaQpXNGYVfERNVvFEdO0o7F4lBIItfPOcGZyq/R6Xm82QP8g+/qoFH
VVhYD8UNy7Spd/77wm0NXJcmrj72xd2A/kuaYUtvIsSOJN97KFjWSJrMBMJhz8Lr
jr5DHtHgj48VzJ7uGiQdvQCpzjqMbk3SL1RpS6WEE1NGvXXsfwcciqXTpZGyKgWS
fy2jGcsSWnZ+76LYo57emB6bnqKMvq5KwOc6PGJW02BvlKEx+a36pWTdjHIQm0I8
+3qpm5pCqdJpteFVLHqNXb9mqe0Ev3BXcM/QCbDuUHxjvvkOU/lm2erRljEHABwt
b3LaopRDNHRphKA40E4L0mK/ErrOyZyvyuFMfSxleJFi+saA+Tw1CqoUg3DxlAxK
TBrHlinv0bEhz+PegHRGtoCY5T1mhtH/GLKIp/GfU1GMMso5PjEfbqeyMiZitg2d
s0/Z7cPRM4SnchdFlPr19GiWrGVf1R+C7ygs55wEerPrRUVJN19pn3ct676WuhwL
Szu3+XN4jmSfW8qDJ+Ska4Ra9olLDPfeWvI67nPtD8H+ZTNV4yTXGIGLIagOE/Z9
tIciKb5446mNbLGPnNXFHKVoRs16MPCHm4wCsXOD5Sw73VJzx02/FYLwiROFZZB3
Un/k0DpMYdyjsQ3xmfnLWhN7ed8A9YRZeZfCpgsYvCuOQUrpoBzFo4Z1BP6IRom7
MDErSu3Ua94j/aU05Frhpd4+qFTKTEU8GeTKOJLLe1E/QAsWaB5WGesRGNZ31jb6
SBp+4pfC4Js41KZRyziS14s4I3ACc+EjFbTFkPBvAG1c4SlQGnufX6vyoHQDw6Vg
oHiQAP9PL/j/toozCJBJ3uvJbn04NPH/0y/k5yHcv3ziTY8o5QgxPkEd7rv9BuPG
DDdoNL/BaL6s+1yoQ84CX2GLZb0zKrod2konHZuReiwtJ43iRStVLus8VzagI4s4
njsPz+SJsFWSJNM5fTEr6GYF4leUQnQbrkZzEpmSsVfC/CFKog+NT28Dy6hyLsxK
2Q6rULjGOMMEoNQrCLOftzIYINE6BFKrhy+uNchI1ldr0KTwr5mYUuex5IHxsqY7
Ayy6OWVcWiJ+7Tig8wuSxSqFCs+Kmj5vQCzIJVCnbSdH6BcZo1PxE5gwdHxRxD+s
pLrvMlpTWZJpAClKCMAAa2qMb0kHZemANZiqP1y8s/iazodPmNKxSalYhlUDeJc8
NcV5FdipRfC1zWnXPZKcaW2zb1w3Gkq/zlPRCQMMv4nAr7lcfhbwa5eaR6NysIFV
L/SloHdt4EZauz3S/pvKsO9y5iNWSR5b7jlaSFPD/MCrqoSBiH1tj5+QUF9bZSVJ
+5lcMntwTrtdctD36ExnxvxtauKnHiCBLB/UQ62Jaom2mtridG++t3F8mU9BzVQC
vcocrmggtAb4dYnCm24yvi0939QQ4e02UMrKVetNOod5tFeYtvOgo8vUyK5lbjnA
OGEhSy1z1OzsxXmYExHu3J9ljwfHyuN7D0wtJgDMvBPYeADgpx/rh/R2ltRMVB8X
UAUnU8PuLVWGk8IlPQQHErJK2o5ghNpTszOLWK+NyTcMZT7LpvQXYNWnceV/NZTR
pFBP76cHICntt+nO+GWaAT5gqTuwdR3U2DbdfnWnoz2IyggxEE4EeTLxKXN6oolm
NDs/4Ix4lO3acAphFZpeXIscLUfhaBsGSAZcDIZyhlJGcN2V8/9/hbal4fK65MvL
jv+4C7yu/m9wvNbhMISWiXG8ohwNFbAIbFAsQBiCUPQdV8aocuw8HO9zskEqAY6I
leIeScej9rWU+uhawYXKoR4YnI6yktUYu8qxkWjb1mJREbcWHPHics2osaTrljz9
Gw75k0SJyoFOUi+dfGIiCZWk8Uvey7sLWm/USg/lLAi9JsHZyGEwStOMlwqzTLlR
Js2AVZ7lc7Q/1FrRdf+0mR95N+1iORrFwdKFxkacCpVgq/dVgTEhWf3tIKL3geTW
E6qoeFgeB30lKGnqSJZ5yz4Rp+WtDSJszsSxSur08LlyzAQKSFPH6kJnDxLA90lk
+ZbEkkZYcaYiHwM68UV/QC+0GrnkuY29rPyP20wbgkWqq1e0VvSuQZ8n3SlS41+t
4aIELODsoP8dzDZAdvdx+3S8yUzzzHMxZdBqw+5Fnv6ZdPKx9GPiABlvoytW6466
DQ168mRLE4t+zCbcDrAdu07HqrpEbwU2ZYuJsbi44Oy8PQK3BL1hGAk+rF21cH1K
R7/gSewyd8s1zlXC83g6aZeR6W97Bt0ThOgUIXJFGMbxiVAOr9YIrhneComTXYVK
R47KujIulHgLq7stjB91Uu64quUtCa9OSQ731TuAqEpfjPoGpOBH2dPmVNDgg8Cd
qJTMOQRCgc6qiN0Q3ZVqF9uGWyF4QMAvCU9p94+uc44xiawIeQqzFT33ssYHbJ35
r00XVYF774t+A8Gsd9Ivp7+I2mLAxsoyfiSNxm/wzwPXGvdDpioKQ7z4Dz7RCj/j
faKUVlomMd/lXRj2kU98gSZGTHjBEGdxglJJySf3UuAWyBPoLd0/JDonRgdwKQX0
l4CHn94rmGB33jp7+pOnLTdUNnbR+nfqjBFduQxN/jJcRkUnwsjuyatr+cpqqBjC
tkDoNuCVGKSggg6t++M+Fbs7/AZg6+OoohqmNIKSGtPRpfVQ6pSmnVyiCek9Hob6
l/1Fl+vsCAJribWG1BlWf6RMxxogZLaG4PlWp2yk4XC3WJs4s0mlo3iQosn3jT+2
Gc5AOiTnG08WtAKpowfDqsjwpw74jX424sRe5QraXF3kqK8HTRFIEP6JPSHOEl6/
MXgnUswLLnJWlDKf8FliKRAk5R8pKszZmAA+4QVWOJ9gBwrdappq4bcQH4b+Ctlc
TO0xc1VpFwrpsF6V1pwKq40kTD6n/7wOS/VOo+rxkaU3HJ0bwijy2HUN+fZb552+
hTdAFKKWD04O1qczEV7VWRM3Q2E+V3qbKdWpVTVsvFiUE8UhXjm6+Iahy65YLkbL
ZAWruBpkYbqjCo6ZnhyRoQMF6fJIVbgkG8CjzpkUvkB5e8/wEWJo9vbPIo1+4Zn0
h9mQ9NBtmWuj7LfOUEzDBrWq3ZRTDUMr+4o9Y2irqNIFdq1HcMKjqur0CrYOxSXe
plXvIIa+VkbeMBlFJZ0umbBVJ811ekqZ7F+tCwhw3jKgCaw64QEf+i9pyPK6B6uL
UInXnsVeSa6M3BHksqPUlm4fpsmL8fBhDQGygs0xwxEzT4LMYnDvE6LOKv0tpfPl
voKpGAwXBa5AvHmqWJMl5Ob6Xi1ksy+twAF/9wBvQWqt3ef9NjhbSI/8Smh1tk4o
QTVs3Dnm22vX2h0LUhTbQRQJbjqHjYw05Qwm+wBPvnyvlpVPwDewzC+Tn+PVO0la
tqfYgUVyFla3VF7gy7yv85AZpCBc/LWK2E7xsNavMp2ghjVhBlAGO98laf/9pILW
W2kvUUSxFkuKRDIsI9+wrmUIsaGWxoCMy30AcPsZGl47wbmVVDSmHe+ct9SMuhQj
e0+ypkIXfTMyWpIymqU9JC7n1X4Z5zuO01FP2SAzk89orZArj/yoFSmWCFueJuGB
mB0gDx0JCruNQ0/zdzF/iLmrW5d+5z4hE/O3fUHNg0drqIlUpBpQu7kGx4HmJsad
HWZBT8d9Jii1CUhpMB/QES34PrDpzHsIZw69sATAMf4uI5J/Zu7egumHNjieGRA0
vFhQH+W+yN/dVZE4MkQgoTlbKRvgLlNJd+nsBJ85J2cu4Eg8HN754QQh8bjpCEWj
OX773BpGkyzJ0PrHt04vHtaCJZnzq756bedx+1Se7Q2l6mvgnu2DYLm0+SYtK0iB
wH60e2OulYoShIiZ92k7OccoeJZZAYFbvmrHrbG/C8pjNOlyJbLWhePqba6sAScs
KR9vc5Xgclr5ZqdoIe84+3FAjTkn+S6isEaDtDgs7xOxpvpAoZWwcLTQ7cGebna0
dBYfj5xENIAxArshgOgUh91s0amfnnfEGgc5Fpbbfm5inyiFDNup/ZmeA3xMYjZq
ZFUGZprzea7743zaOdiR85pcp6ikOSBnp4WG0PEdmRaVy/qlFXprlCCF60/nbqzn
GImNpkVSM1k06kaWFSaqOnUUYaOjlDRrijIHIDb8hfoi/RDyWr8d6FXwb+1SWHyx
h6lmkKDXepi2dY6PWytzVZ2kVnpbHgNttVXtfWbmBh8NTP3FBXulKZgkeDZ8ycKV
N1ODez8UExTiDMBwddnszhQwX5UzRbN8DLjQmuPl8yi+3a/kjt5rK2zVqb0/tVO0
5JWgC2oUQ8d2PlnE3j5Ke16WHAQ19TrjI/TfKzXxOAugrDzR+H6XFQtkJy9Bmpil
3kWcUY+CEuFj3DRUa8baEmCiv+dE2EB0yAgDoecbLLftyXUvqbQwzgp7QOT5DldR
EGSP2DNT81RJGXjbApeRKZNDqwjoYzTVBuHrrt7yFBuCiJvc6Sq3A77/z68sNQxc
se+ZrGWC0sAoOqursDcEwygEIBgINzSG/Hlc6AbElzkcyw56gx0xuIzOdzW5WKbm
4anVK4xehtDyCh/lXm5XCbDbz3k0XXABhZHwHE790jBdd0C2XaRX3jrc8w0MHjV1
K+Oefc+WOVM3Hi7ekCxWHiQWvATafyT2lFWv4Y0xUy4x+S8jmNRQIMjRD16gw3lu
YRBHg35uSxSzKvKtDsgzvgL5cMge99PPVwBbGLhJj7eaNgt1QdkD2jujmNc2Gy7p
7+Ge/NKYDEvZSMUn0bBqd93/pxTxCow7SAF+gbFX1LerAg2AYYBi2lBFmF6IABLv
dgrm4zTfDg9v5b1x5yezimL11pcYqwL6pbtYJNYxDYMbBunU1zUxXJ7Bk217qZF6
q+J5q4//Ez20z48oKMOASiwr/OCLPFWk/PAlJ7aE+UBXJdOYPApWcDUD03h7+OoX
fw5ZT35DuAtzdLtbmQto82ngnDVy92xUvGiEFO+mF8PM7fhLBFq00SFVsWfKxxLJ
xkeKQy62X6/wDYNlvv7yMloNqFHYgsbKdDDv9Pht/v09yRu5uLQR19niagFpMfyX
/o2qin59mjEC3FI+p6mj/YUsvgqD4RgAbpoW+hpEWKq2fXfjVGFRdAexZckkMEhK
johrUTssG9L7WArbcC7UQz8STCOfh+icwRXewGzI6j3j/cv8hf6ON5rcyHtnGZxR
bD2YQ7hT8RD8xrV3H1rI0rcwutZGdMI5CKlb2Zk1WQ/wg2zgqC+n3rvnbrvfLXF1
dpJXyHvzQv1FNhqkEQM/P1RbsG+ckAY93kieAIMMl1p6QT/nfOXlfClnAd7tmcf2
N9BDIFuamFNew68FbbZNhq43QuGX5gXom5UmSlDMgt+Hf/364MkvZQGDegls3tD8
WwJaFDh+fIi8bBeaIf7VeFdoa9xiRi3Ichlxioch4rW/5CXgUb5BCGBmtDo2eunY
23gROvv3UQk/pnnKNLMR9orMEhjlVxJDdCdOFwS47sWwiUD8bucby14LNCAx3Vog
4T4+yXlIo8Fh4UJHdI4+/NLgg3oNvDGDkH2H4Cfy1MN5/Itv2O2V8hHJVqFncq4e
BXRFifLCVArQB6xTs8UMbLGuym9Qr60s+Efl+UHhAQNbIjJGvkXWDwtVOXClz5lN
ETElEw7PFslVz00n8p6sN4LHTuoXZgPZU8DHZJEBzmFex2W3wReu1xjHEcOKlYNy
7eJTP694O8pyma0HiVfEJGQAK3UnYLKNcwp4qZ+2CtnNoWJtWsNd61kmgd43+sHP
96NDKVIYMw62Km8WWzQfNWj6v9UTZxNLgqy0HHkG7uni3c3oIe9Or3SYs02y9Xvl
wmX+X8Xr0E9Z8VrgCO14HMi3R0Dn99Yqauqs/to5f3ayPuJzXZcNC+Fo1lWAUKvy
K9ySvDt7CfQJqfnzRvRbmOFaAeehphgwXSbeTejhAYhSMAETV9PErymSrUrHRU8o
z3esYO5UngH6dYV8R3shQ4qHLBik2MmusweIN6u58DGRQUiIi7v2teCJVyUnv8kc
p70wgl1D7uzt4kIbSdhFbzhLoLt3FfI9FFEC6YzIs+aeW55piL+kWg9dxe/Lbgvm
xxCmrgG9WAK3noBjSXQsAuOaxlel58dmuwZBviffLv9MYUsR8SqM68J88tVadYe9
QRfUpVZnvh58JQ11PCUaBOT6C+ON6I/6ctR4Y7mdXZ0tpJ1flEeQ0ZN6vIfmNqFU
bRMcTnZpLBnvpM38IVy++iZz31XdhljHGBC1CuwxrhJnCj3tBSiN56dU7WfMTXeN
Ok8IL1IJy1uk53R9YE/zvYwZlfg4kn9TRH0oMGWUKlRvMPf3BZsboX7rZW2Nh1me
BOyyIo8nrUd84ScQlWBQxI4C8N92aYA0fNrn+TNA6NKnycZl94l/S3pkJoM6vAlL
dgSaz9hTA76L7d12k0PlJSV8CWobnJQb25XbN2uLI9TTFCvgcm7elhohgD/bG7Pe
nLnK91G39HdlIj+CWVDhl8Y5VUsp6BSRO5Oh8tDBoO1r9skNU2PRX4e5EcphqLq7
q3yn7ZscTJRHYgHLCgSuo76GxhO+RQSayrNvnUFMGsbusqwscEUyvqt9QZ13K3wE
9T/SqMbh7miXNPUDpdM4pIPUv51jBHG/OoNLX3CEri7Jh7pl42R+MB/I7rTzFUui
q+3lstOF3+5D7NP6zP9xpdJtvNAKTraj0TraoM7iTuHkYLRoErxw7IZ1QpGq+Wo4
HmPaBcHKUNi9C9jEjrywKyfwCkrczojvCc/L8+A/tyjTFMfZc96kEbLBXsy8meBQ
bxNY4QXcJYoRETubWei6VPSXYu5oIfaV6dJnBQ6QwxRIbh+6WO732WeDnjAQjzvO
ZVMBxqW2ZlHmJADsCSf12NqEtLWkhT5OYZ8+pvvcRKKtxoyHK1FuN3wjchpqaOsG
/1x8NzhrqL0ylfkx0S2FOymI94YGsiBM5WMqS+en3eGbxYfb0eZapn/BBeV5/5uA
UcO4xcRSDLqvUgQ9jXt+yL5tHvNe7wzlrFT4unEgSJJQ1V1TfNqYvrbKvRAR2jMF
dmrcfgUmw+NePy92kpDDtFveBn0/gY+OidFR7QWoAx3k4Pr7u9DYL0vQCB5ruFx9
5Z1+cIqxVrGYf8zqsji9oIGq+E4/PB5la6ffklSQfT6J1rZ3G8Ow594Y/6YYayo0
Vyrb3NEueWkdmSPYbgeU/m4FgU5I4EnmXSx0LeUqBI/ImShwmnWcbStXW799bsLB
R0rWChgmw8JFBwc+4CBRw4uVRDXyHN1cLnYNoAqlDp9MlkbBYJLFp7FmBDkMhg9v
b+/qZTWmUuocSbeopawJoBGHcXDNAu7F9l73OdfK/MSPjQwNQMpO0KBeTo3+D7VY
XfV0oYA+9zdxr7NOC7UB0rN9PvwDg34YDx/YwZmaU05MSPBDH087xPRvWIwB0TMJ
Xr7mIH+/kYjOuQZpE++5qDfUiFVPempdtjDrTdf+gCeARcRtubAXS3cjHjafd0Xd
5TMQpWb5B1t9mEIcJ6ebDwSnK2fK3o9QsoDYKsqqD80/zckkpI5GUAJY/O55U5mJ
uu2TWl2yc4o6mYJrIQYMghMRNZOvqXdXMuXSDZGNLh3KtyVz4mwhiECdtxxzvTB1
RugvfarVhdnpUrNowNqbSdEMiXMv287f4Lh69P7rtmNw3cjHGzTmnrhBtuVI1Dyl
i0MNi/KPwgCRzbu2terh6r1FMntL/wmyXCviJPcai0xS4e5zaq5jrxhKvDgDM9li
mw65WWTKAPeFmcD8up7cVKJlcmnJD6hZfeovRGfIKKXS3/aIbGyB3AKshTXrwPmx
pr0IESDMOOTuVWherZheMVRknNSl8ZSH9212R/AfdJArS+2QYkYpLU+XpQdAcvGb
bvz72MULy/9oJq1s1Ppa7ZUrUBIh2KjBDZp7Zh9ixyTJTjDhjAWIUHNwR7rB7BX8
91ulqcFImwCW98t8Yy/IEOHj+V2UsLNtUACLQ6tMnKpv5G28ND4MIYMDutGZK4fh
zYtzjiQnH40+IqnQBD/EwA78WVV8EtaQz+hPyTq2aqELLUzG0G2g1ROlQDugD46h
DHH9w04CPOOTFxjhhZZBdu/6fH1glAGr1qiALIIN+puOtD/TetIZvGvH6rjzS85d
QtYqoyl8NUuwt7wQvR5cs7kTvmORuvknyhtNOyyDxGlQpIoi3JUuG5rSe+QLpZPW
TQfi2GWGd4/xfj2u7yaU0f7FWW5Gw7+x6qQXkmYt6YdZ9t+UnwTV1ADO9EBDyyul
tIM3JY5iQZ4YVV9/TS154W+/psJ2iAwOnlh/UVQjNDOK/nEglkIBBKWkXJIen9OO
MZ7iS4UKE7RREd1MYpEJWYr/zp8VSBcU5rOqDfaRTRgGWIweaBbSDav2vjZx7vs7
h3Jc0K60t/D3TwKIxrKYC8FbPkscqhnmJWc9Sbz0V1zo4/okid8OG5o/OQqHV7xo
AsI9sNhhawqIkDoOpa5Wm5GClCMVFIM01YxsxGu5SpvwBVdEoSlk3AzSU34D4kgx
pfOSOfpxyVpNTFIHK/R+9jS+XnVPH3nazt60QAs7AXcXvBIyb5wIK7LqpaUeET+L
rwwKbhtOlyFn5nrnN0lWnJGuZ/RAP3LOTLkuB6zLUaEv7Tmvj0CAQNqWONV8wYM/
q1mhqWgH1QACqSaBTSVirTFiw6rhDfs4LRZxTHIvIegxSV4+p6d5tFG5TkYI3bPb
1YyU0LnUiI6Kwmu8a0HCjrHGgKFVln1EPmYYHrI7R8UnTHiJZZCHJ48CCtw6b4aF
SHtzDGNLEnW5Y/X/K/v0xPa60LL/iKCbg8dJTLrbhiFTHPEvLzawf+BQLU2zKoA0
evBvVjZxWiDVoWDUP1AVvnW3A7d2sjBc01eTwQe9wXAaHhJmuBJoi9A1Vr4q5GyN
zdy983eDIzjzxgFOjSHfjjKY9JbdW8sDEwFnYkNVww3yHb3s4RU3QdHPYgeQF3Rw
cSsCgD+apv1OcOIffWRMmaAsWCR497kLUUVhwbga5/sJq1Y0aMllqaeu7EJz4TTf
7ZOPzKErFhO7L9HQ00JHELkbzv/ym8azLO7qZRLACRxsmFgllsd+6VbtjE1lZjYx
qqVzRbcX9eOj3gWNBY2r3ufKOAxuLZpSN/3pnB4Q4gxPTIcS8xigfrrYode8SBxQ
Qf4QRvYHJIMsyjpfTNYYJFSKBKUwy7l/6QSzXbGHl6on3nXBSjMAt0oFuYCfkIHB
7JkPycGV4zC5thWPD97YSW5wj0E8pGzlMiyl2M3azKz4B8GuWWqsmrhzgLeh928C
uPn4N3u7RARWD4kkrjQ5tipwgkMn+qxYsG/tePhLp58MI8FrqWFbbMPlDFnHatxA
JaLQAZfaWqPx+7I6fTKNGj5E1+Ify/OuAo8i9a4S7kwtPpgcbs+GsLSstBUWuReK
OoZlwAcZZ4zxGHJg1cEIEjVcBU8Qvs3Kio8y6Em2v5mJywbLqhJIgrRZPcoIHadj
aA9ugDkjLVU7CaV0EsALrQpOBuYTZVyS2rCCsA+j8MrzVyTT8pPDtsKqzWAZDQVP
lMJcPEa/UfikGDwy8sHaAb1EfBPejRKHYIymjMMF4Jwxw1K9kCxnnJvYxDBsirW1
o6zaN4Txdw+Wm5SLhgxpsF02/gfH30P5/yQ1wOy+Jb0s665rd1nN/HqlHtLacLbb
zmkKx4ndWH3sDMnLv/pUZ7ZRHVbyIzmAKgEKsizuV7u/Ti+olvtffrtgsgnqq52x
5WipD8bvqriaL1oYeq4StOytVKJicR9Z0HI0XMDP5GspqEML/fYJr8UMM2q3EAwO
tx16usem5U9S/blJ6Blbyrsn6IG9VaCx/YOvpz/SzO03rtaGbBI/q7zhcWP3ukMl
nHB/bZ3Y/IoRrmUqNQ5u4iHGk3a87sDhXmPLBmGB4F0GfLudKk5gmyNYCe4v1WEz
aF72g4rDWM3FdG2N437JN0xo5yZVB4T/vfhCIoDVYbbvad8y7M6s0hPD0IoYzZ7Z
MkpgdPD4oBTPO/Q5I23KJ8wWgC1yFrmqg85YsDwE5kJe90g4AHNfv/gq5uEL8yZL
l+iyAAyfqXj73/7GIyN5usOuB1kXoFPRpUYcGYhdfYytmX+tlUVbnm83UIlVYLgI
rjAho+kGeK80Rk4D5aTwBt29jti7wgrMmo0CRAYKh6jBGRVbWt+ppLMsNf3rLG6F
FNxUoXoYrlDlmaWpJNaijOmwJVhUbwL3WmhlCr8uqF+xdRfC/G84oVMvxuJABYtW
NkUAMnFk8Wg/ye8Zb8z97Bys8CZwwGeREn3CoymvZdafetO8FQ3VTbHZGK7PKNQh
VGRgjh//gczPhaYuG+u+GHbZTuDZ3K/wFbZdsppnJqfKDXDZWF2ECHOiNLadrg6+
AUX92QYqNc4IdGWBKHj1/S1HKUWDkGdQgrQ5PHRFEir9af/E8QXHrmzs194uoKO/
y4s/r2ssYqKtZ+XckHwsL9PcBsItCWPUkbuSNdgDeOJbgSzV0uL67ezc3D3bFNaA
2MoZ/A+UJ0Y/re/VW0eQc3WksyY84uNEtVvGHJ6S/D10R5TckjEUNbQI0jiY+mRn
wHmduQ3EC1VN9ukG7pjcVqlW5hjh0FYVwPgbpjDeTvRSZhpf3zIXdNcxbR5BoLOy
5njs+0DOtDKSamAQQ4D/41r/vSQiR2Y4/vCePEo67vt1JQEVPOg0V9QNnaIu21Ch
HxrfbCUPdBpqZ3KaCvHKNNtKc9gsgSIZYkQlksAb8E+DS99h157da3ukN7Cdg4GV
ohrN3dOkJQSnIDoNxaD26PNFWzoLPFQXiFwDafDRtGkluZBai6j6fGyLGWw52Hgo
i7XrProybpELeG4T74oxZnfX/aFXsVmK2zcn3y6AftLp21DvZG0Bb4ChMHWxnSR0
c3sSLIavDpyMZXgajywSxJ8vuf/wVzwk/bpzwq6lnuK49pkfAVMX3KNSygZPn+7L
xAEzrsYlkBJ2kWfAn5ktmkstfg2MyaLyISeYJR6puL8wshUT0TfH9HBOyPHRqW4Z
qKnVubMgPLnXVu+h4QEzaFMpRireOkAXCutdB35u8MdOaM3Y8mH37Rr7frnzk8Wv
f+4xUyjYrjLuR/d8lY06x+skHRuV/5nWLiHUZx6owPVzWkFX4h7MWL6vMZg2eu9G
aR9wM+hyPOjUCZOgvNm0SSJvX85Pe1tOtvZVaxHG3imNpvSZEOrGYVeM56TqTbri
/g//7+cUl8s7xISFQZwS7pn+SP1ffI1QEaFBhOm71dGDAd5PWiPBBX8YUV0h9Cbf
Villz0WW5ilre3DVsmgs2v2YmH9Ki3tnf6zoauhrqE8625ls2JaIEjfX3/UeDiEK
KvvDVq0OmxmZw6oUQ9mej2NNBaVHu8amvDPYuQ6kZrbrV1SlYTOHThu2IMkILJPJ
1Fy9FWlW7NvCJZSegie8u4LFfF6rGrdEPde7FK7g4WZE7P2F5K2UfM27p6wIgEkn
Z93611f2p/tcdkhe5CkTVfBuElgWvkhdImEMzkr7O4g2V9CVc4SbA+MOeW7r3fpw
vjaq/u3TQZGlhNw+1BvOUTlkGYjx1WftrGBARxnqz2EP+p/mDW+wSoN2xs5fF9cl
ziH4UuD8rBqda2Z2iMD04ZZIG1omBejEGtw2+ZnV5AKuKQjpvxc0LP+8u8YePGmO
zdWhVtScNHThO+l2nC97/So0p4O1gpbt4CE+xCXrIp/uSEgB2vU4w9dws97kL0lr
33GG2JBh7o/PUupj02aCuOZhBglN4p0L9W4vgI/wlFZLexksopsrexAUh2atzSXf
dN2ypsH9LUgClf9tUxVGry8AhkuUp8oTH3jHT95IHwGP5H2KvCa8cKy/Gujtp/EC
lQD3/bB8N5yG9GZU7FrMlbv5ExLcLP2MGNBzit6mzbzGgCbUZ/h0TJPOtLuWkvOS
AQ9CJS0A447vsgx5lZHIQB89QxGnrk3LLHiwgurEivAjkoZlV2wAsv2yYpwfuwyY
xR9oApUBFYnQ+LsW8xc0c3zEAjrmGDiJhMySKDKIN0KVRrUzqIiwIsXZWjl4IZUX
rmB2CVtkeT5ENIG74aJOyBkfuRo5wBjkxRmIsdT0wEZbK97AWgU3UJgoPEfoqmfb
yp+0mGXTX1AxpUsHh1fyNVABKKXI+nNV3+SrXAjl772xF1rcgYcKXHOD8gjRg3KZ
QmKQojw28mv3W8S9bXpZAploYp50+EfxBoYlBUWqzzg6ehia4a62MvIjTaG/OdHX
Ac9Jag8K0OuDXkx7WAnHsCm4Z3o+Qoh4fVtXzJSRSgsUR0qXg/mARCnb73mNw4xK
GJTpq3E5zoTvTyeCU6nE5CExgJq4F2of43MXQcBYKVTAQQZbcGTcY5ZsXAHCKuwE
Rcz3i2OMKkZ7fA/LSZ59pXvzNvHIVKgYYeQa1tMpsuo3iWQ2oVbLWfwdCi+/O9Yr
pA1f2aXhgvtI9QD9q0ieTxilG0IIGZEMxE2y89bDdIKS4VajfVPVY0+G0uxF/s82
UrPa+FOl5oTtsCz+ldCXcSCudg2QWHUmzTBoQC1FQRlPARM/bEfBocyrFDuwkhrU
SMxbtYDuTxq+GM6KEwi29E8FoIS70Yv8JPwZb40AMSNoFT2zpQZM+1075XJjbwkw
KR9l6aZefl9TB7dD8SuvqW2tUdhM+AXrMYTQJvq+SoXNQD1ciQBgkU9WW2aKVnkw
E7fFdS7U+E34P7rKD9/fqBnqrh5asboXLcTIybbvAii16GHHwX7qvbZ5QcTTux3X
xphjUiKsb7vUYtKBUhbq6dqmKrbqafWaaMbwUVi1THs5autEcgJGpupi8OdKSF+a
l28MxHhyveDnZ5iGyW4A9TIEu/nl+DWmMqjrJSbEmUgHStJ9YL7GPiuF7NK6MCGD
5RjMh0zTEp+20QNG4/8Rn8CyKgoNs5Svz5DgHYXzH31uuSCmax1Zj53x+X0JmuI9
dvgXhAES963PgnQO/xtdtyOT7uN3QAZK0zw2RpzjN74DxRkmP4AwDrQ/so244gt+
nnAAwBCOTalV5znPJclDhxWCTwuApofrdkdD6+/S/oSQwGozJrsjMR+nzemWaCb8
72LmR5kO1SH09wyrFyZrx9Avnq33tcpXd2JxvXHu3dfQSVcQ1p7rjtu9DOywu9Ve
KEycyYtS8Grs1dpD7sorxz5LrTpLSg1gD0duQcq9VgqarhhfW8npGE6mre7oN+rV
ENSii7hFOo1hZx3YJW0OIPKyWPmXM6UWMJxqvuhmR6d3ozx1JzB8cTnb7J63Iaye
Qn5g8VfcbaLhHAXs/yYObZqlvh9YXnhTtnPs0unOSHWsHMS3A+lB+ibZxBTl/9FC
MfeG4JqJtvERRY4foINTtJMCUJG9L805w9JdZVHMGNEN+oHRomSZTOsJEHCjA9C7
iIw1Muk9kcSNyILByklpW3AhlWq9CmpQrRPE1pcOIvBvLbGEZJQym1lN6GQRXRi2
56vAxMDAGog9Pa6HZOyXOr2UN8olzo6bGc2kdEYs8/Ti8vBrlLlg5a71x70LBVsH
dm9k/xSAqBpmqV0wtpFI6JGdOaI7VxdFyAnojFE8WcHAqbIoASFvPgAWL6XAEnEJ
a7MJlP+u7uGNd7P6rEK2V72G7qQkjALmUV4bBJxhc3trao+Icq/I6m8QNTyGfs6P
UGnYKsFHW/wyYML+zCziOpdUc/xHRnX8JTF7/3RXFYQjdgEnTRQfniesiRkeaDfT
g3WFZHBZgqAOJ7SCir3uj7GQuGuwyrkkOmk+Br5ZwPR1PCVPM+DyRFPckzy8OlRX
Ew+4wWcJXRRn+mrV5YHriluUi0aqWJCvJN5CgtgJAcKPKcUMVLF7MeFKLNsT5RDs
z+MFnCD3u6O5r8LBjM5sNUwtUbNuUhoZrO4dSdIsrnbMNFYkZ45PJmtZvyE6Cyps
RNMutjvUH2l4tF82VN2NotVAiNH4fNsj2483p5RlVq4RXzXlWzpm0tbYa+2ut+A9
FpNc62cVOEgkHrPto0Ub9r17wU5PX4rchB0NOzzmczSWSqCTGdITaeVXpRGIWnz1
r+Mc18Z4ZGM+qOOPbLO+IKe3gSB7Rlr3IhYLISrIryPEVjbNOJ/GDylrK9g1WxxQ
rHSKwXCelr+8Rng142+prLztYqsV0yfsF/IpbBjGDkU8HtsA2jmkuOVdl7Y/oti+
omHPPdZ26OtknlDGzvFj+VXPlD7lHqKyAUrMiziiDZgyP11gMxDRi0E9K7AGJzOc
lDSZOzCWbARYCJkI5OKtwmW2vIK6zag6JeLXWSAKR0p+pPWem1kEENwDg9bZ9qav
wSCxhrC5S8DmWsNO8w50WmK/0GorJeR0c/3rPXWnG8Q6FZeaesAsSSib5WwsYlDz
x6YDIufLs1iJKmh7SSAReUgyyJKmXxhpV8TnIvYWlrahAP+/kY7Vr5GN3XYWtC3Y
a0oIYJnQKv0gzFmC3ujgkvvcHDO4Htti4XRtz3IxKD9KHQ3DpHqUu1/bg+8MZu/B
zrE8KoVTTUn18iCulETlNHZxYurxETJdpUil2p0Z/TmkTTM1Ad2GhDILo5Plms9B
iwzATKcARn28KnGCAjOM/DkeyzoxFAESlGQjnH9J9iPTuP6BFP/k0vAzx3fU0QUs
Nf65FRwAMklda/esc9VvxRvce7MpGuxDBo2QGdlC8oApgApNkSN46wAO3BdyMDq1
tU4NtPQFeiKd5ZOfaPHgddj7x4AbIeViH9l0b2Dt68uSnrfvC7uLKylnDOVa5mN+
lcIUmj3OFiz3FLUCWDlcrj7W1RoDLcVQX5J6srokRXdI9QW4z+wkezUpcpXEa+pG
03Ioh3rmuPAKVmT2IZjT/ukr3yhI9EaT0SsgkqyeOjJQ5ajDyOi6EA6riFZK/E9n
ZkKF+SIrgZqe7m6FgbZrAmGpfNDqprN1zB20yjI/oh0OPZGzu6iRS7MbegDf5kJy
dxAbMRl95Ys0qJUJrIYuzUDY6n6s9OWtbX4MGrbwHCb2V8nhhkXNU6CGnUtRtLff
cK9e6NIUTqSg7vMqc+6TmJdnk/SJNW0y0LcD9pjZSXRGKa03D/R8MP/3eL4lH09u
QLH5yZ6lE3OsVxz0xh1vznbC/kdfVK6fwfQvZSOsq08oaSXpgzaghHQNu8DcHWfV
tpNCqDBYJn0DTCIZK1KOgrirwVyCa9vNwWyQlvEfSBWIW33e0/5jnTZFgZOCW8kK
2wBsTUOTbxFRXF61VjnqqGWAuxJNS62Yr/jkFtYbhTXT9ifiCpI06sjGdvt7RRyW
NDl6lOt9W44LNCE4ZAEc5V1YFihRmK45fkhe17zDvViNoC5RQCdTY/Bljskqe9WH
kOFErJjJNY+tVBxoM1WaH3YZ6A3BvZ0YnmWRgullgQBR5DgYnV+C6+D4w78Ovoz8
krOfuYsn3scb2vEwiz9WIMcRE1V319scquemIx9xT5uFjJqDgDxK/aCpQKkFKNJM
/X8aiaRI1NN+bsyXg95bIBrhTe6kRCXNptIVr9NEsgoEniMUmcIN+0f8m7NfByCq
1UKMjbeR8yIgviUyh2+FloUwENyQJgXMsuS34DrEqNz2iidznoEUxs6aBRM5LJJk
coa0/df+uYRaY6nXSlHy0llItGP7L/EeaZ6ya9c+9O40DWWa5obOLjVn2/CyK4NK
iyUpEVlqJvs/2/BUQ65PM5WqGcU8mnylFhlRBI9PkEIrQhyXk+vGhycCB7JQzBbO
SeRutJDxODR/FMoDGCPFvIbcTLF4CDqoVMewIX/oR70KKgjgpNZ+K4BnSLmqtuYQ
8llfbsGJz28ptGAYRQTktT0JjZUO25bEgqnEpMsxFH8OKNP/a9eannyXO6oYrcsp
XyFVtFj1d1bCdKXTGYyqiWFlprZ1TVBKBi8DhL2ZSro7g+OKXHmXssnyZRj1cJ4Y
OGJzoL9ExvbVqBqMXmSjid07pigWOi9tt6UbQLxxNJqUa1CxNoU04yIHibIm8Q2K
My0+9d9x2LGR63qPGiiucPwEktzy5FAI03j1xJ5YDPFs/y2lfaxe/zRc3MHvclzb
Y9GSvUJXww0M8oOrpJWhI11WNwRNvZwmv+g/pAHyFkOjp8Y0CQdZ3DZm9Jt6nix6
hvW1oe0DtGZYRpBPpSoONgy3wDewNmc6P8WPKRytHsWeQFa+n95uhny3jOEv5Tsl
pJaeeXjryK7zW5DI2iadkcxk/ObTrRjP64fbv5hSwq+S+AgdiKVxp9l4NihUkpxy
geM/IABjIki8HPa2wGVL7oAOF3rhSNXITdN0knvRZxkIVMSTtkyB/B6IUJ7WG45g
MnKKtMJVRi3nI6JhnbrKVeUl49t1onn/MCoi125A07bM3lqRAeyQWwsKjvzqu+WI
ftE087p2bUG4rtuNJE7RbYx+xYC4F2dX/oyAMAXciO9OUEaDen/cO0iq27VgMKLt
uJsXcC70MU6fVegFu5AEPTiT+bXdPzMJDwAJ+TbBRGJU3GBbRG/oA0rkzds8Ciem
un30HZuOd67tkVZJRbgzGoj15xvry+J1R2kWMxA159fGzMfr4VkJZ6okIC/1m0HA
i6Evdk3Z9Y/Rlxmuh/907ETKKflDQsoG0rl2SUaCVA7lJ2pecJPaVlUbhwbu2aQ4
wXBWBel1kbS6VE6BiptNIqqwhLcnU/JiDFA+fdnj+QIY7/AoFHrFltWDbqffLMiW
8nBshI7gKVOcAOJmR9kJ+UClk11jdsJQz3Oj80U1ffXc9jwT3QOYSlOk7lMqLa4k
HSU8R5RKYNdOS0G+uX9Fso8Mk8KiK1RoP4kfLwegi+q7FDSCj3y0OGC7bezBoGJz
L/n/WnK7GhoxrDrEIobm9NdBZYspjawjSA0yV92i4ATmySNq0muarNaM3Hdzeoci
092x+PQelnF5PjM7MN6oIRLJuIFGme/bP8UQS0WS6KtQGTYGoaaF/xwfWQCf7Hl1
SVjDgMW9Kzr4vzsUOYOmR/QW5mWWrEYaiSrFyZe230JkWIHz4PuMzPETFb/kDaAf
zkqIjlesHwSyUl+y6999b825JdOYQ72BPDxHocbe//fN3Ii63eFlYTX8mDCLBJkA
tNxrD5/n88BckbAZO+LV5vireY8reDt9q9H1oQ9YVTigTTV1lh1JD64e2Dlkbfr9
hhw8VhaLOBtBv0CW6pTPjoAbJmb8DEFSMRyVDvf31n9iEapKbnYIQJEP5l5CBi5D
D18IFFP6MlQsG+ewPMmiexyGnldyqQt3BwNZAbafqdwUUMeFIywTKopmA3hE6en/
Q2byzgo//Bim20RO5/3dJihCPJHHJHF7vqiGjl6wbjq+zLVEijRgokC4GG6dvvkJ
dSvdLkrlJOtXIB/Fz0SQ/k0m7+wU+Z6PBfOTsgbciTmXQy8PrCHmCLRJjnysYITU
vXjEuyNoJKzJxXUw9+IYA5Ei+MSF6mHwDjkg9zuFOBIkEJTgFAxOVI/AB+2Al0/U
DhRfdMf2N+e/0GQx/bU+KwPiV3dMM9E2iHTGQwT+SueOBRvsdwTmTpukrJ8T5WJB
3ntuffNFr1/ntBKaOQqeJacFyyLZipsaN5fp3qyUjq+P/1VHjDOy/p/vs3zmAR69
yHIL/HmQwixoPHxYpcgSGCuZbrHdLXGLwSJNtkZo2Ev71uDXk95AYbUE8ejlUOi0
b30DmDE+kXtEERNVNkvsKYqWJ/uQMZIcE2Nx+87j74RHRXD+70XNF/G4+ewR1Vsk
owUolA63Gun1ILV3NMKOzjewiHx2DCXE7pRSfg/mpVMfk6Abih6ENQxznKMl/psg
ehgBuKPb6fFvNGagQpJH+ApdNKfyq0c/96Zpg8eR92DIIjYT5CWU2OqBDzNQpTGL
ZbmGDUrArdkSDbppvCDzpAXgMg0oiUCwGoKVfBOEctCeW74P4rOtPprjmSxniPCb
53CVNyBoxVRb8dBWs6+gFCmP5AwzsgDoffhdpCgurKm7UrrBJNFvmzNRu+5PN/o/
/UMZN/DI2dyBbwL3ZU/vGBdkJklh5PGolZQGLIB6D8hSMH6idPoZSiD6/JVlsnxv
QQlndATdykvNIIYyi7s7zZae4BTcQxOMwSpMXYQbYe6O06Ny7B/sxo3HW2UzNmFA
OUk4AP1E4NQkbgs7+z7feyaUfksgzVlWzI1J/zRZVZ5RxvVEzcTh2aWQylABn2cD
kl0vc5gNMVkoy7rKlwoWFisEpPDWL29GfoOgv+19k2xAgC7eNNNz1RrDA1De7Crg
twQTa13Y1Mmjlq2P1v1ucoUP7KhosbGjFEnj/stQGTTZCV2iHCgB51S7Fbt8J7vJ
HgvbPxjljxg9II/ZgErwZBfWhEANe2Nq6c3X+v0BAYVtt8YT14/dqDkRFzVEQ2c+
CqC+iCkZsTnij3s/1R94YxQZKv+Odbk/4WDkNmAQHnEeRF13wwZYC52VQOcd4ZoO
wiOuoG46PYH2SDdcJzw/6DgwDycm0ilwRCRdwQgJxECcgn/Piq5NiwguikRspILe
Ty/sreAJbUF/xZ9T8lnl/yNieRSMZAVcdyR8zBJC3WLaLwxcq/bi8cOMaGCkgzo1
qlrJW8F5e85ID3c13At3FHaarmb2ppKq8TO5fVUziOtFrilZAileDKpo/9/reunK
Varn5KysYUSg3DbMTTMSH22GIxJ0qx4nRvADrLrMD51oe1AyZJ+PAGUrEkuBfVFD
wLzZ/iSexfkP0W3yTJ9czhLJm+DRU/ee3b0qDkOt8/DMKjasGX03239XaGc/z1ts
6hr7SyeacwkTU1KePEY/svvzVtxt1Z+thY0g8nA34wYol+AE86/QdMBFpZSEZgQu
r5eXf/r2OzSs/E7WV5SUoHCukFhlQbBQInuvnwuKqGq6wHY283ykZph95JQL69z4
PZ7k0LR15dc7vedIDKZej16WnpbiE4CeJTVzbmXRLt5dIKmRgidSmFkEJ8bv92n0
0XEeyr3sP2zYllhjARxYRCvgyZIQ5kldE5Df3+XXv4walwi2W6qQFtkXBtrKNQ4j
FN2fY80ZPkVMLxyWobpLgU4J+8u2v2HX24skLmSA3xiCSjrVy8ExEd5lGLxY3Mjg
CiVHKQ25CmBeNvMnsRMOXjjtzQRusTPM9KmZkwevqHOLsoTlKUfs8hGRZLxS9PT6
y89p9dZuLNiTWLwyRIb4D3sCkjCKA/oKP+b7PFGvmhtBONQ0kpO7LTZBp0/TF/ME
HoobXepb4jFv54Ab8XzbFPnxRBRdg5gVtC7zq+jRgP+D8FCoCsrt2UUKNfTMEzOm
AxEM6vw5uirZGt7DBt7KnMKFZb+91Y1cGu/ab3hrIjOjWS99U36vpmcDb0MawLO5
HUZlLWlzFk5IcJo5rvaWMLz1UZjblLRz/tKqgc30aqVs/19/O7ZUmA8sbGijrlfe
OWDxW2YpTaq8yWtL2/YXp82tOLYL5wj4tE833NCawyxJLqetyQQuB9wXodW44+OL
tybt3OuBR6d9Gvf9W3F9hr9NP0j+3puzSNYvXdaWJu68CcJvlWCOmYJ52qt21pnb
84rz1oRQIAH+qQvB3ytWvWmRuGRf0K2vMPT6bkLJ+huIXSgbVo7bc6daVqCSet9d
6uHtaWmOmlco91SzJsF7eCiSsEQC7cWyV8KzMvDKiFiD52hyex3HXGarLg8n1t2R
PSs4gqKReq/n13rvOQKK2+bXnhNyX/kiSnlCYVgd/djuFLGKgfzp1f2in7Ve7Y7V
B8Riu55I4cCTXGZOfImSoSwA4zn/1b2SrJy6GJ01tRjhRS0EmIe/4fnUJRLqpXTI
DQbHTHvOUclFDcEEwUQOmOFlPzsPlqhQYBnmX5QzNNAy/hAH8PO06hqUMxVB4iSp
RAc1+FepcWVomhyznTvS9qPkF9awmdHKos1O1nKUQ78OAeDEUOFnUJIoGLrn2//d
a4GWrULM8l4TrqI/uQcaOprTJMrwTUVTF92+HF62IpmJEeGHR2j5pLHd4/HUNt/x
KTyXWrzcsWIwJm2jZF8rz1gbKZaBytOM/2S1z7F1UsvPXCPzyIEhNwojp5a/O+Cz
PfnFD+Vx4nHqfp6hq2Fw1NyD8vCsf4FP3vwHIwEONaebH5kPOvsUDXDkK7ZaBQdX
RTKgLWR0vSE0T52Lg5bMeDQ9xQQDlSTJGSCxKXR6K/42g1Vl42aPXMSukWGQpK6r
C5mhrs2S4FjKzXjzgA3afdz8R1bZ7OzqH+QwmPX/acUsk3sn4xP9Jhy9uzW6/Jkx
kQ1Z3oy1rqWpasbp/efqYt86pb4Y72xqWlJ6dU0ynYg2XXbb2KuZNet7528UlK4c
4lmz+Pkgx4tgdW6hpx6XMbRX0uFCdKDbbpUNexfrbM28qDfUVEzGlJmDkUfME4mX
YpxjHSuw10zp5qW5o6nOb3O7g6/n2v6ORKOr2eKrKoV5OfYrec0w1106jPpXHClV
izj4gA6MCEFC8+BY3UFt7GzooirqkR1weSdNb6tit1wwvfnzlLIbiQ5/sZQ/BDE1
Ar3Jff56Xyp2geimXKMIJFyybaGR+ws0gj0dfYtMWrmb46hV6vCnlg1DP0xWDv/3
do08jUeB/STflayDHfurHrc7v3WNPkLM3m8U0X+1n4j1+smF2yvTg9UhRq3Wch/z
XroTO9VQEmXl9JfLLw1GQdUMdiUSfgV1b7ZYEdseg/IAy9a3jG50ZG9RIRVCAFBx
1kG8jnRVrmaQ/GikGcaVTVvhhuRqo8jku+zJtCvA97mY6J03i2jSk0g/U8/4jAYL
QKmI0HRkhzbl7/Zr0k48Gbl89YKz02WyciMZzuPZwE5eu/Ujff+KIpz2NBmTluYg
NTqToCQUyhgiRfpENb/io2xr2vNBoaa6uzbYW/iYk2SmXVQkFKu9w5750bvcYMwo
Jo1WO0/ujCKsnvfonT26CaxRyUZko0fQwgXw21wBodP9HNDvRFQxhXGwPo7JbS2f
nXr5/Zy7ODGVnFIyrAhE7Y/4JoXiLn9lLMZuuPpjjQi/freQlRdmQJapvNpVBRIS
L6HONeI40DV8zru0AOGQmRHcNeftf9NA2q+BnpRy6luB7FWiQrYk1RHrJjNmG6OA
rGjDJvpv1A9YkcEKBNzI+fS7n/PHh/yEEFIDiJmXtT8uiQHwMBI5T3uhURW0tZTR
WVETmc4gmAjz+kOSHY0LlXJoEdpoeotEf+Nf/EkePvawA09FdENmXImF4fGg1iAx
YBJmdLiUhpUs+Ds2HnMuim8EILayZ/Ak6ZOowySUIDxdYcW0KNiu6TSX+FxGXUWG
SyobQTNQu55HkIEcYZUiWqoSsOx1XVBCQLOMbwisA5D2cY2imRf/lrMzxmqRi1zg
1NwPDOiNLi7n+U/50Md+LLcksm4UkqftPipNb/RYEBzFxgAO+U/my73bNPhaaSR8
A13JEByVQ1LRLFaBaFlLJtS9VI1o/vNG+/59LUnYPQSzQaWUrF6C6MR4oi1T5xxc
KlxrDcqcUGZlrMxv+yZnOAzTvrHyyO9dLfTLTxvt6l6ay6ViFbv4KVYtBLIMgPNc
jjNCEQ0Xal6q7/ic0spAq/db+CuBJidNLvBQWtHQi8qmRHRqIvOXrjDKkAhevVpo
62I0t8f7w/y+RJ+rcQPUhaxy4UU7RAblwU6YlP9pBqRj7/ohMK+x69z2vH9/zZJl
rg0FwGVjOumTMJxL1H83yhWX9qu/Aotf7RFzImG2vSfE4eCM2xT42pFVHWyY6/rO
YAjFw5HPplV/qidq53Cgk6pA9AkLwTBnVXyYN8qj48hvnpA0bKY4uhLfGNOfMZzE
tEIPUN6TDClpyh5QqM4QJVBdc1nqVbYrTXFMlh05XqPsRNSnMmXYtYLoE9V1XrNH
fh3ovdDuZfVS7GngjdvGkz4lfUXK2aoAj8XJoIlt/vBCdMuF5/bzC+lWVDIjHMkI
mhfYkz+mgMtiqETegGLG6KPJqvnKjFITxRdp4Fnyowy2NH/4+niiuAOKgIAKtwfp
MB6EYKUyPlf0PtX2hGRFvkW7jrc85Won7H6tTf2kbOsdL3XQ7mIYucblUdcpRB6j
uYVunwEG+v54jFau6V/SNmsX7Wqy4ZO35W+n7V7/2GjIGKMvFx3tNIanCihFaajA
248nwg90BuXSSwxsd1FjW7edsB9AF8XIud8pCM6UjGtIkcszUk6BNZhPLFn47Tc+
5E6gZJWMwZ9GsRVHoaPWXw/RwXdc/Eqxrqm7KtxILVvWuyUetgPyDJ9GK6iDoDu2
scj4FVrJz5xm/Ilaj3nZ2pn/dTFmsP8WuULYOFLOqM6WiyqLZ25uoaHtufwZX5ui
pCgJaylSybteF57IDvR9hGMvY6YfwEB9oFQ2xum/WAAkkKwWmJrmUsFQMq29hxaU
SZiCbOIoyxTgB8o85F7x4x+1QFcY47CmVALAfeGVraRixwdyXvEyE/YMXElX6883
4tcObKkohQvt5VF4FcjNnP7UprgBRVHlFFwX78Mwg/bFaW6UrznN2JMXcDR1TB0V
P5R9mFRq+4UFJhQAGW17vj2k4FXlDKrLIpMO1tLuq3xjScvihyNb7wm4zsRO0Zfj
vPwn0RNK8Xg5DcUp5cmLbOqZLzXnhIVQ3XMd2fvPfUFBRNrMS9s90HIxIuHB6eA7
DFl/QmQM2KTUv2XQ8L0wJ11467/vlN18JL0SxrDyfwZeyxLOcMwy6SNRqk3of+yB
GKNHZ4UzHWMT3UunSahvSblDJUxIFxk3yuIlcwj9SnaUArk67GIsa6Ef3W57h67h
0VVtma8r7Mv717JE+QW8BlihOqE7lOxNrxpLFMYMHLRWZOJZUUMXn4LhxJtKayRK
LMapF7WQINPEtDNZi0zuZbt0fjp4Sm3bNLHsBEqt7L8OdU43Qakhlx7grdGsCrOo
5EkiTQjAm9d6lLjv2G8OBlaVXi9Mo4hYW7ZVBzA4DJptyDgiiMJOIIOunRYu7kBq
ajEg6iMuJ0WtOgqCOCEg2lKXY77tIYINbhzHu+rdiGFJeTeYdcSOWxV7KJ0PSA/j
7DOzA1kkd85nKLHq4uPBOGRjJfKDlboBtrALtIqFNY7tOzLyINinghnRW53HAo3d
JSeE1C1cHTqOup5VkSEY440vV6Y9mbRvJimV8G5n8axNqaNyoBVGl8x+olXCaTwD
SdWW9hf5A99wZkM7ppfb7/n7D0cDNYDYjDfqlSZsG3OhbnOUhXt5kc2Ucj23ljOB
GzyuZFP60d9BSwS2SocKF9pN9eChsE2LKPEp33Hpq2oPeoVoR1/sIKNgqlJCjtOE
FxQa0KIc7u058KHd0Gm8gC5sWeUm44lr41+svDE0h+L+8aQbrud+9Of/HxJywNCE
Rn8QpF8eJ2z/y11/uAL7Bx698lJLiVEHY+0KL5m9jRBTyCCJyiwdrOiE78X+w2XO
wFxK+PGL3YsZktYxAM3ugeinFR8zfwOcITRrzDzTNymd/aym+iB2nqUBfPbJh/Ok
tgnehDhffvKd/fN3uiPbsf4SRbRNNqmUe20RGNBbsObymGoGMzgooaN/6bYXiOD9
9xiTyU8AZZplThVFD5bR5mu01TC+Z+fXotoM8q6V4SbIdWhc02ImvZtfiUFxSFzO
2A+Upj3UdlSp3dJGKe5c0thhVt9wgWeLjP0Zubv2+exhM7zL/54GR7vT96Hja6EY
pFdkK0ZJjucdjbeNHkMAOR/LNny5vinc8xrWe9o3hRk+4HbAVPyiTfVtoY1rmBdj
BJxe8nirSjzsG8NXvLjhijX25R68efL1yUQjmIvUIcJ3FjXRGlj+DJvJnebDj+jJ
SKYNaa3LoMjMvAii8ZEJtrxjCWM7px/kGJqFm/oK0n/zf/uYcPddEiKWMvLkstUR
2E191wti8ba3KTvJPE4g6Rcn6vOqLMijFsJMIY5aP7eVdbuxFVz1jkFTDJnT25BS
2y35vr4veyeBb3jcM42pL6leSkWcBXnYgQkpbGn2k1SNlUyDvNRggAkKU6pL8K9v
hxKoF/sIe1ng6dSpqe181lxonzmgr7aQNGMFtjMfOd1OTT/lHvcI/nKh1nmjcmx8
4cwbveIK0uWminh+v6NJYneR4/curotBJpJ2rNrBFWl0Ni16FHdn+vUVj4LBqddl
m8prSJeIYKg2PcBum8Ubxx1CKUSy7IltBDhBbn/OYjbTiEBtYC/mDwJHPSHbo12Y
O3K7Cc+fdJiXpBurorsv2ArxiOhevnfM4CsHIuFPHaxOu0u1Lnh1loBxXnwYqRwY
Lv8c+AoceYDqz4OVur58vrGICsZHSex/U5r8t6WclsGgPz037FAaBVqaTDxNKiJm
B898mT0VVTDRvy1XrAr8LPhiBil8K8L2hpoYXIYEJPsojuQCfOJP7hcTT9Dq6n21
4pJzVdKMMZyis9M0Frrys3aPUlKDhVgmsmlz8posfrgJRV5MrZcOf1FtlMrbIb74
HEoSylM5lLCvraJg6NE4Dwp503vkLYbGYTLDGkEx/SVV/YIrL8KKNleK+7NL8H44
Cg9yRyZEOR00YiD0nijglllhluEPZUoTz8wtduXtWfwlzelY7KEHekFQGE6rq/Nz
rup9A6sdTA9kv0bS9UzN0O0wgEIF2ElKJAdQdG56jBcAfBTt4KrOrmg0LXxQSx9D
n+W0WL5VGJ9cIVoyqGpb3ybr9/zaWOiZtl81YwiYMav5iup34Vche46m603QUf3d
aE70Fy5LrN7KoMFIIxTQO28esAseEAqIg1yGztAQDi0GL8mU1nhMVTnQAl8ONMKz
jmJ48ohV/tXyc8r17H7PgWBYX4xWk4WJQ3+rUmJ/UiD35HWGsXc6s+elX9mKkwXR
6qDnT2gmwyYlSzRc4//NxEfJcZ6kkdzONVFMLmzs79v1eiqvjSIWFoiTt4GpMKLn
xuJD7otho0AiVMCg7uQHiZ0iyCOsaPOvB0dAlnknXrNFXgAUCnO7cG8Xq64giayZ
45iP54ufc801qYqGGIVfrqoUEiYw6+ElpWvFAOzZaugil5paKpUFtc6AsJs0pAoj
puNqBd/S3Q2Zwb61kkWHCMWTrUsfy57Xsiu3hj83qFZAyKfNsqxda17YN5TDSB5E
CMwAsquUOHLX3ftMgRRZ7a8/Rpy/ytjZSkHO4PdfcjDu9LM9spGP+2KFAlx6rbej
BgYsXVmGbyl79X6/UyIkhkBb7QDm8UzrsOOOVV2bCiCYS9kyuOwVi4Nu83gcJWBx
cJru9vY97f2ldHE3C2xZvj+EQPgfHxEF4tGAh7p0lqdWP7oksZJuFUGrP93lzmmK
b4wPNh/0LfW2Yd41mDM/3c2+tMfCRDdCOoi0HXCl2AAa0M6jqPR8Bqyu3qf7DTvf
GwuKPIvpfANmcc6Yk4TfZsckENwGyEUOshxKKcbAmrBef4xJWyjJDU7SkzAqiIfE
q02PPxqznh9OltwKLg4bpZ+Xb/KXxScOpOZb5/TKuG7qiiw31RbcdT8fbIqftK2g
IFR8ULv0yJOCWqPocfz+XpOGhxnhgvQeVQF/F/UT0D/7lbrnybyswtLm0A2bOnue
Xk0YAsG0UH7clxduEa9J84FTQp9b8AncJf1WitfQNOMnS72u5LQqdGudwKANikfj
PTwBEFtQ8a9e+UXtd+W0Cw0g38sqNYWylHTwllr+mk2As/NYi9io5SgL4gvVxlwN
hLiBTN90WEepCEUL/DAiXeF9BBF/5EoIxaKuoDzUeKsMUu/Qd4HWtwmlv4JfOsN9
s1Pul5HDJpk8uLjJfqgoCuEDXttaPuQ1QbAZNWOp0smqk+fQib1jKtB+afC9+MwP
OwJapzxSRoeJRAA0ouytgDLPvJy/Tg+jzGRhnH8ZrTkpOugpfNo/4Xbg1W9KNQZa
F/kqrcGWVVMOAQdlQUBPhQzVGyF7RBYIVG0BQsuzevwtIm9ZRJQ5GYKoAZLP8Ycd
FM+wnIDaH8+opvRsuEZHqwpDgluO+uDHOaEHz9WE0XHygYB5NWKZxB7FburqOfbh
mqhYXw5aE2WK+M6l7vK/iWdSx9i7omR3QSRxF0lIkX0mVO+1b/JIzOhrmzXIEpTg
MEYpOcVV5tMiqiIAXUmc+dYuAZgJUK/GlazI9C0HXv/sOKcnC2wTMdHczS89eKVX
UN+xPF6p1VUr5n9/5sxmFdWTPDgy0+TLFJ+/cIbMyNjQspHa9gH/6sHrLrhLWey0
gjrbWZmp6edqD1ADIa7w9xhcCzTQswdaptHpZf6BuCoKqU6ro259ZmjUG4CV9h/R
s0qeHKA7dP0RimJIumlRAI5PhdoJ4BrcOb7JIhA0h9+Zy5m3MS1Jf09a+ih2N5vV
NM8gMnyDziGI4Fr745XAT74A5PxFh6H60ixfOrrK1n549t/EOcciLHuuqZNhCEd3
7HaWmLD7a8WOPoUi97+c7HyitblZQhCLBwSr5my8EmYxFsiQmlrlTybaEhCoiI8V
AdwIfceeEuJwPELdC/ANN4lU2j3or8leXDoGyPETVRopdi6NitQ2nvloNzss3173
JVajj7l0NG/Q+naLufxCr7u6HqyDMVGfd8eI7w9JsEv+9EhutmthiMn0h7V6EYBB
Jau8CGf5aQ6StTRsLck8WuBGo+EcukACjkgKFT1j+O6iRS5gQKo+zv0Fkh94noFA
35Byl3ImgC9g7gF10wZmDD10WH+Kq45A6aLrFkQiDN/2GoviPcw781pF7zan36tR
SuRlnsHiWWDXzhcrPZFaj0BrY81bW5YYa8RRzeNEKbiD9OVSZjwNBxgw3wQYzQi/
6zgdpolxNtCPkzhzpBjFdbceZhKCSs1UsoMAZVL2nN+sEAlpu+Z4xgo/PbVJF2AP
WYQC2vXrO/qlzme4ndnlBBxoaUy19AoqOl68LrmL+Ka0rRhHeo3FyLm2DA7przch
cXKGgH3DO+jIm4m0l31vriTymd0shx7QH3M9RA1aUSmYXQ459Jsl0l/bGvChijN8
GI/DyWItqGKMYfmi2qO/mqLmFBMVnGHMHYBqA7DLfftSLMqJLLAmxeBxo610WiYs
9H5haiPFv2YHpDOP2cei/56VksTdgWd+nJFm1th5SugD2mDKm8PuhKGym1vckDIN
J1ZOQQSaB3nDGUq2myyA5DGSg9rt/B9VWUiY5KiIoLb0R4rPlXtu0P1Hisd675qH
770UX7WESBS7Kk+4LYZaOT5lx7Otb1gM6FRe5aM+ua/1ia+8dyYpbRT8BYd1Bd7e
QgXJMzWj9u3naDDZTJmzoWxC/jHOB7cbeqLFaFks1FG8tiqOSb547vNQ7EK201Oz
usfD1anH3fDAhpAvv0j4eB0Vg9aG7n+38bzDlFXtpY7nx7DRI/LVr6j00JmoF/E+
nsipUBzT5irIW2UR9DyR2ui544UTv6Lhhye05OSMx8BEQa9l3MqhXPPvXL7eNLTX
ghIW4UMsUAJmZy9lFE4qg+4xcZag+/mjIH5Ux8XCFAjMmKDfGXn6ZtPxE3NnCDvZ
oXamuO3KQRk+3+tX0IZ0ubm7+3T+DgLK8nQVZdTM0LywhLB3civ4NOIYbOCqbzZW
eWZldSRVyAPP/tAYv1TakomVSzSL/CI+oBi/BerFxVukXfdh27VLShmw+j6bDoDR
LH+TuN3YWUZ1EB01bUsohs82Dh0o0wVrx6yOiErOJnsb4oox9UZRbgLO0RxGm0xZ
gGg+ZNmmZc3lXlUwQBwS/WalvaYZ/qB7nLGleDS6yscqe/6co8MYT2XXwnYYHAWu
z+gxtWNbbweSPZ9XEAO4tlw4YZ/SqxnMHxAAlKS2opsI51xHkPHCFKGBanFqqWl1
lX3oMTj0PuGK/Trd3TRkmtk2MlUdmODKX4JmhFLQ85xH8XyRklmMCa5obLO8l79E
H6Ypb+AvQa584H4Bs5I3syZiS3K/Iim+xqAH+0/WORtfsAKvZDWeUHwb8v6AaStR
ujViFXUCylsTrIXDnd2CthLfTCa3zJ0nbrX1qAx0+no5ng6gzkH9uYHAl3e0GCE2
iNaMJvH9qoSDhxB5wPgkGo5PpKvkBwIIzBMfYjKs4b0q30pydppANFckXHBKMIyS
IvoSd4w5amBNxDHRoFEghKCwa3rGxGQkGweEg49pGE/JRvbeBT6XNu3Ow4UjOOeJ
P46WsQskDOWEpU/CMrvS22bjb/Y31U31MxG7hknQKAX4Nm3AZ6vT76HZKW3bDG45
jRkuk2vuH+W2619LZavsEVo89v37CzKbBsVAxzszoLeUHJiwp3r0Hl5IOvVSmS0K
Ep4i4eP0D7DE18jxJmXxsBd2QIP1MPvMX4R212H5qD/2CZ5hbce1Pwj3t0L8QAeb
n6tpFgZjYCZWgRyd4Tv6cwMTTdtGszMRXD6/zFuJFtDaQXE55Qz5S8XzxVUuoMGu
AVZkAeMRKt3fvSY7qUR0CMg0CUBVBYTXI0FfaNrhzbGQCP0beQvugeRCqmLw67+f
4eAQoFrpPQN3rCEUZgcx/M/AWf450PfItmBpWhqDLDOzd0Eesv1THuYwB81LRH4k
+Tk/7Yydc/6HxeNgPu44aBqt3u3a6fbFjIDFitJgplcGH7k8Kixv52Hu2ijUDpTU
DHqgv0AC7f8mio8KfUEmnLDwLju9vNpKa3UIAf5pfoHHe5vO78hkar0desT65NG4
evLx7ATx4+MZ53g+ktNsEYZFK2+UbNJHltrgrIhXe7vsqwoDFYa5Losbn9PeeI1p
7cFhjUzL+1vv9c/iF3vWIo1JB57Ipct9v9DEOTBZgGu1PgytrAZVkeKDCWdskLC4
ZYTOXUIasBQOKjYkly3PHDZN3COQcUrZ2N7t88yRKBz2V1jb+8VU7HlLBgDoxaAk
sN9m2KqvYRTNEx8CEGQSyJb70W2o0tYguImyiceBQu8MpiL+Q79S0XNh8mRaUPuv
q6XLx1m66QDMcO0fEFljDqNAvB94veTZqQnsJ76YtwbIi5sTEz7zqOQYHy8npBio
+qEWlYbWJWmXMylqxVMolaBOaNFwVkJ/h2y1JfJyp5hGlq717ADKmCTKAZksUc8o
WvbWhmkEeHeMaIfM6YQJMXBniEMVuUmSoE0yhAIPmTY+bi64iKgkj2RJkJRp8mPB
ep7WqqogDpKQ6hWAyAyv/7n2uZI2OKsqyo0Ef+DUvd7j8pfFgnw9lCu7TYh41GVJ
Ru0IBY2qzkcNFlQDOFJLfnYvJ8rORj6hpeSaG9u1qwXXy44D3l3yttGkbn4DGulC
7kWRrRWJsB8YNXJW7Z4o9JfAdGVB/xSBZw/HfVWa4tS5q8PcajjmXydzBe6lH8SK
5piIsgD+OduMy/z21BfrWy+Hh19SKWfIxHulGxLgaV5Zv+6U11NEnJsD9BiQLhMs
s4VJPr05Suji/P2t/PFQYdKP53WJrGRkueF920Q5Mg3EnCVd0HVG2kpBOEnfWTHP
XnfbJSk5TlaqekNPKN3vZZ2hw7w8cj673LmpGiQfzMBGUttn0Fkw1PjEzOqS7iji
rYGXwfIOKOAXSmJhuqjX2HUOvrWS/SBfh7GbeCW1cxt+Zn1xoMYeYAiC4Ms5/yOp
wac4BecxuphJPoeF2/fyFTTQC8l91WyRDYGlPMAGMxrxpfda+NOg4udPBbvsnNaX
fAQ5Owu0ITk85PYZE7jn/rXOFPOtU68hJ6d3FqDPmU84VISKsBNbslXraxJjP4DT
OxcoOw2Fu5j+Ptk9wPvHcS9aYMaXeSipqCbU7JWqcpHDcqDP22I0VBJ87CpxRxJb
Hj8Z6DRk+51VAQbbUPo1jaDW6C1kWk879UhePudXQDBumdWh8ZLfRl5UqhiMF8Tf
az6jeFKWA6tHFCU+bQl524XG9dNtrvuUExnFBz3wJq4bRN4X9UHRoenr9BiYm4gX
S0mIHYQxLbYddttVUrKW/btw5T1df+cKTPFvS6YovTItMvOZ4fbv4/tf39ToQ/Wt
GmLqlkB0cIk+YpqE2QjVd34IaNElFqi23niGFIaoA0qR+J4zEPQDbUR2baU9l2vA
uBFdBzWb4VrjELm1EAxIEX3CviArJXISuJqsPpLbj5zmw8td7Eq45Kx92k0Zn65i
ODzJJdtCfc02ld9JKnRwgMNuu+R+/tmzeO716kKbxqwEYqsWL7H3u719vnvSOjnm
22BMFbyTrefw1irIQnq9na2XYmhTr+XHqVlIB5b1JB+nIbxl+mZ1Iio7sKATkRGm
fPV85YtbD9VkPIoB00MtOjpVJhuqi/IZx8UbyWLOpEbu8tTu7L1IjreDpwbH+Rb/
W4Uig2uAjC4oSeeg++q1TvqVOTSupfPnPaIpsjowxHSQef5QD4lkqrf2888p8TH3
1mjHcHOVRgcHNI7tRDFooMopFCRJ+PhGK58zXNUrz4f7ue1gPK+v+cft0CVgzPoC
5yIfL3ExGX5Lo/VJu04Xxi1ncIxJWV3tpW4MHcC16x0PJcm4VA3SlNuccOejpnuY
Sa9oUQBdcxE1zbY+D6qqSGNbTau6ws1VBY28B/xvC/kP2oxXXfl8s9kvcbgh9lS+
UNu58AxUXWBWIRmzUTRL41B48gvvBqJisjAIfsl9D6/ANzSB5eYsRPrezn1rAFVI
LuhL8emB7GduCoFKmqF5F+nwV3qIGN6hoIaNQFvYbNbpkdpjZOSXPtPnyp+kTML1
S0nPcKFJFMNkLrq50WYON94LQGuK6lNCItyyJnXIfTikMT9LqOedDDX/P5DcWRDi
RV7O7kcQaqtN+thHIA1ezbLPW3i4xf9ZK3EKIkhiPHZEe1FuxyTZwlmGYgiZ9++R
MMjfhvGuGffp71Rw9Zxx8ImlR+NBm9YenuWUGNcASvVN+lpkDGZNUs3lbiQwe5ZS
WIdCsFQ/qZTTShxqS/X8BMWq9DsRY5L9tFvQvcjkq/mptUAPImHG7Ohl0raFeFug
bBihWsIASQkKgqEzCN9tfGJ49RVrdm3DeSBWH3ECz8/WHG41JcZbIIE2CztCsCOK
1MAcxDGPd9mIc7gG2UVneuimihhY4wGaMVJeRQn5a2az788n4sro1k9VN8NqkQJd
vmQFK5Zsf+QkUcRzI9H/wiFdh5cj4WnuR1vuGLtrchLCkUUiqw8lWsvsecPGD6Fx
MGbsWVYq/6lOHb3aHhMatiNDLXbpAYs1UoiOLxEtBX9JuQcSkhqP6YBsD0bQMMit
WQjVMr3M/CB9KbgHU7w/0smqleEPH0R14K9K9fq26u6SgL1qHaB8pZ6YltCKuwSp
JarXOGg8vIR1/PsNsrzYRDfc4dUf2qQ3l4/Q8hTtTuk392WrimYX8VwdxwECuuZL
UK1EaGignNposbBmZhYFivxb+XR+OuSa+Xxs85qiRG1LXfGASMX5tQQo3bpSQlj1
cno+e5JWU3KVpF5o7obDZdfPOGdmB5NxwHFVdIMZR4tJxDGxgfKmzhgQRxUiaJj1
JSI6rmToZctyhwKPAqXO6sLJ4ZboGxieUTCTOdbNUb2uAGZvtKLsyDg4uBy7LRyE
sO6WZGk5JeRpMPhdE/UsNnJdxz7qZuVRy27/zTTWr92v4m7IPEukON0u2NvtvTHl
A/EE6Cmf8EVjLsBTMOOd3OSE4DuE4pYNakEhJTmrurShH7ZV6F5Bp2YzE5r82Fmv
NFeBWQc/6ksyCDDrKpBu9/JtV0baVvgLtZyGVXqXTxVlnmwdGaU2EK8kPvqQEO8o
PVAFS38HV6KvRhOlfI/pZBsqY3C1piKo6/7G+9Nt69d1qJ/kcwR7YhvFQKw79Bnk
e4387qgyc4oIE04TYVpeHr/H+3P4pFA+f3qOgBw+oMvCWiOvtICMrdmeQjgSHRQa
K7tUsWoF5IMhZjJvI32NfLfwza+uNyEDOc/agPEVF47CqBkvQn5krTv0tWlLlJ2w
+kypDXF4zTbAdBhDrJnlblJxmig+zOHaYTL63N06Rp0EOYCY7WGyZ5BP8sfHJoz+
eQj5FJsmVhXMT8ScQr+gNrhb/p3hFnUU2P83e2HAcXwW0oAe/piWnkG7qb+r8UfW
x+zBwDRVAIcek+xu05ZhBNbO4bXdg0nvt5zFXCmRpS9CFGTN+hbLr5+qYR3Tja2c
045GZVYuaF5inYh6vEG6xGdJ3aiVbYPnbUI23+n7Hu8ns0XixJZj0hte2pdUeQYL
nAU3yXaLuS2Yj1c/Jyw5Zc2zSvWoFo4OQF7np7qmOFjSpW++wu0a5vqjJQPVyb4D
e/p4uwlH19Y1sn5HGYY5JHdZSCYQhgztHk5uWmcR77AkK/L2+JPgq6dugriVbB+p
VhCwBnKZvTjMDdYei0hhznRVSrSBbitXeJJ0Hzh2bzEQo/9cxZfsW5/eINi9aAXv
7E/JS4H5mo2mpVxWvsiPhghlGl5KTb9E2CVO69dJ//IOtfVzp+XeFEIXtDWrVAs9
PO2LqsBpmN3gleMtLTfwD1BFQ/wwYfsEd411SyBXke+jBlpFww6GomvsKcbS7Kp0
fAAW/k485hza6d+oFWxOhUapX7iIThoIaUjzEYKj10wbRON7GPYf+F11s1UeX/LJ
4hSoPLcXQBtXuVJFqPj77GcR+SunOqz+FhNvFF0on7NSCHPmfvaarBbrwOHUfphs
QKaBfa3naKZFm9gvG4gFZw8h7KzdcxBNkRyQSeUBtQ9O2ZgkuzrCiE4ezVdi1M9C
kPRTlQE5CYwmT4h8bivHoYtX1TNHJ5cCZgOO0jyFgNoR4apfxwpf9vZlFfLGfWlE
ub2/DVdLYjBiB6Q/mwkTORn/bnOgDH8bUUknxA9Pj0pGXaghQ9d+214l4z0lPpjC
vIHFHgFPFSJ6Y0Jm7xCarmIyKIu0hDlQZfezJ4FR7qeQEBDxY2vRDp/vlqVlEtjB
cCNGnXUR0+RE2HbVUiropfHekzM+N1sD0z8vfTLDkmUWYKY+2hskZnPKALsPHysV
NyXmafb+XQn3V9M8U1Z9nekkjeVx0XIWwYeeqp7QHxpNdqY8TPkw4wvsXO3zz5Hr
WZ2iiL/9LZI2mUDVz4HWNDGMLvnqgfxXV4aX1NE5X8Nj5dj1w+qG6xLdhjKAFdlq
t59LSWHozXyQt+71kZWiqc+gGlDGjERC28YmLk4umHvNgL8qaBGkvW3SWpb8OtD3
k11a5qpwi10A2tyDr5mUV6DmrtxruPMgEcNJF55pvwpGd+ZeZVXg9s2tw/nmbcVG
Vk+2e0IY741JHvv2JrmsQU1s3vEYWBEqDcY5mGukJjbTZQ1zSFfkHBEhPpT1DEQU
8kcZ0RNe1NFCyVACBRJ57SEQPPA/NYNBqQ7nQ7rGwsFHa/d7tBkp2iqYj9i553uZ
1mUDbWfRnQROOyno2ebN0e53K661qTyuizAPakn473DjqR3H/rmLp6hC/OB0rBro
9cNI9FJaMNMc+IG1mdr7UEr8sU5LCBD4U3PLkOqLNFP/AND1a81pjbJI3/MIBBpi
j2pJspB67lhUFWVQM4gLAxmlTdTCZt3y+0cMg3xTWGCF9iupmLek0R294+zH5Ppm
anjpfYkyBTyniLlw0lvEZ5L2IC5SO6wsleC2I+2dd4oILILIKBbwiSdeGCWJQWev
jiF720jmSJTLpLCmBcvQXC97/Ag5voUjNHllMTAk7iya4GWuEssVYxeMtfEacF1Z
ejHD9fPuBnq905gHHalieI1PCkpPFyWVJTzVbFDO3chHtbMcvnpVrgNcDC3B6oNJ
blgNs09tAd0ieyGWuCBUp3cgUXnp9FSsnLd5HQ5esPYHeh6cwY2Vdw9CFeOfI4NU
ZCL3L7BZmBKQOPS45ra0MK5Cv9h51/Khpq0r0ZdmRMQOK6x5398NIYt2rNKjqAP5
2ED5cCHQ0QmnOINJILgOU5Ypg4deGQcbQ9jwifR8p1hI4WaV2jHzPtrD/hrXUwLy
fvm8ClDhW4bZk/JKX5g12mQgzNWb9Rf37IGmnsHtiCaEoV7QtnhbndBVmcEeElbW
ZL4Ef5a5FHLjXpnNHQC/26q68/ECc/ORutzJngmEuvQgiwfnxTzxULUVC9K4Bcu/
pkbQ0YRRa6f2p7UKvPDGZjNCNLYlO9PGlZUdA5zh2/8NQN8by2KtgYDsKLcC9Czs
+CSHLrdwvN7aUCEZygJX5tJGCCsY+v1QtxZ7TtpFMzGErXM0Fa9qcMN/RB67KF1B
SyvWT3HLWDmjqZeWvfEHkdzqzPIXCRHPYVnxUSXxzUi+9y+AmisB7e+hIMGBYNME
hZuI3e1jSNksb4M/vDdvrJz3/S4Ggz4UZkpNoys6u46Gjuyg7/6o4BZ+GNRVW4ZD
Jmbz17Ui52SYzLVEw2FsKul/9Uft1ebKI4OnYr6Jl9ZmXMJdZkoMFOKzgHm+tPva
u4j3h9iMwv/RBscIM9kHoWBBUi11BuWUXaXYA4+YJue/XHBg6NSKADQBP5pKZZ9Q
WGffoBRh+I1GPcrU/T+sG8/BY87LmZXjjksoiL8tzl5j/g54Nbtg37jwQvDHn3fp
kJfMczilAyeKDpzFrf9BXiFOpXGIhGF5PxOuUwp9geJlE1+6v/e5iyHms4p/PrmI
zl3sq7nnOGKYmsiepo8QJiZ8jsExg1z13Q0K84+Q95EwFSRFbN3zJizmZ4GIqgMs
r0TBMGrOB15G+WO97VdWwQrg5hZxkJfwNWkxFhsqsepp5DiYZ+fJXekXKL/6eer6
Q7E6e/7AWwRtBazlEHsoQt7/ANdVhtA4hFCIb22HuHaVWJFRybuT5xemTyqcHwFU
7MxThs+UN03flFYXXn4Q35nO5LlRFA6WEqH5qgtiFHAsJ/DyMtNe4lq7Vz+5gG3D
XunJfqUtk3y8JwpCyfOyUi0Og6VZCRIsurtK0N5uw/+BqkoAmnjveUTYQDcJ2kPg
ekTgQeDVXEuiQXIqNMQjWkrDsW1ZaARAZexVcOb/V0VoJlP+nnZ2V3OQCp12BmUZ
mTnKv0zYtNskngURSLVG7agGGTvnuJU6QAenKU3F5+/k9yoz2J5VutPXb2BDwsYi
kTmD87XqiIjTQekEnbRKFtfpSptwzD7h/0937OpiNCmTmw1O56sM/Mw1aOd7OM5O
cDt/BxCuLjW9p1Vd4Kd1WYpstMmc5UF64rZWyBPpNNjx/XAlvmF9z2AZHf/bhKi8
FhZpvfIDYw0gC5Z/l6V5GxKU3uzjOx1OTY9CGnoZJ0vI6uxYX7Md8neYv5P9ZQBZ
ravFqEHUFW91tnPkPKcf9vO9pJizpMbvwtxcdb2UkHmu/LF/sPXB7Z0DAEiKIDSD
pVQB5jqDbsKSxWNaplx3EIOrYPVVt7K4ejtyndCZwRaObJ8w3yIjeiOxHjE7EsFh
P4b9Ft/f+R55TFNW4SGLelP1mm17thym1pZo4Vg62vbsPWkRUdVZbfPgtD4GzuPN
qIIlzUpZo5YyKuBDvc29blBreqP1V+ScVlTACcrCWom9UEUms2flLfOGIQst/C4U
BunWVjanoULX7f4lmC+C/uAFufJtD/wvU3UJhmniln9usjEvpCcactH0Lw3i5l/y
r/y/977+Kygix6+oay4UWNGe7NZE73dca5+BuK4I/2OvWwOd2S+pfrfF0dO3j6Pg
30uLxA9lFgDhPgrLIXZrT2SL1CbcBAWn9q2/OUpFf2oCzlXO1ojluO7bxqk8MnwI
zlBHbTyEA4mjZvOWM7c1XxZXT4kkM0ENTFKwnfpXdFfU25/D977FoPHU1w1Q2A+f
FZFnTXM4L+Wa55HhHPhsQi0XW8ECcBAQb1LiUUesIdruSOGzovYU0pxYGdhLeRR/
eieOp1jF9QN9mf4oLHsu8ab6ya9wYPOzAgjVcbSdQ9+PpWjYdXUnMMP31DfAZ2dg
wXGZwWSv2YsBWJ9II5tuywWCvGvcYhzcdVeVg3486A2DTL16IlyWvCws5EhJzw5m
nmWpDRYc90GZscG2JbyKvkYGZGTYVzT9tDt5YYrm3badhcUvlyjkqbj70nryBEbG
X6PtA54WYuhOIJU+8aO0tyzJh2sm8QqrXvZe07nyLGKazWgzwaiC1tzXaXq4HV+u
lA0SCPY9kdQncOZ+g1S9CJG5RtLLjvM5PxSrRLtm/L7xwAcq7EnL/7G1KOWoQrdc
jK6e5s7gYA09Ey5CBdwiyhth61tfH2XXkPvGJEkXKjr3M7VHspCmWW4KoqyVPe8y
lxlxu40RCWZ+yZi6xtMeXIqaKwYAA15sy7LRItRFrQZUZzg8OSP9JNv725Hm8q1l
WjB7+uCNfj0WHZ17xrD8pFORE7PTGOsj5Wyipq8YLau+6V8M27iNil4U9/uWVKxd
ujJeywyGpqW9cgGpvM+sWsJVOIOsUC0SiBRbnKD7QvgXQGd4H7E2HaGMzBZUVy63
QGnb/KZtqtGQdhuNUWpMx5NJYJiWh4aQeMaikNySLr0OBJAiMJf1jinC4ZpO8RI7
OdZM+O0OH8PVB54zGjr42ckUcVm5+odV+JdlrDfQntza7Lqvm6p/Zw6VDOKrxknw
toP+X0DsBsDBn4FtKpharnrh5TlwgL+jVriRPUNE37PlJcvo9eHGxWAc9JGbK00i
MWY58SExvPEIcIb38DcmMxvvUfr2wqIOd5uxhF7l6JIu0y145WUIx3OToThIWfFz
CrhXI8t2sjlnD9/T9X47YRCoJ6Nq1RuDhvB3VFV4IVNeVO8zwZa2lDJWfYrlarI2
FMDPPZsHmzMtHci7qrxIlNYcdSbKHce7FrvH1AN1lCmaMSsq0zk7oyU7R05McP5y
uN6TQBTbviEsZOmr+duBUHMvmxGZSkMvfzqZ9zGq4zVdvL0VuQsGGlQP3pcmsWNX
hqdHufF9qIaFWWT2ZI8Ofne0bHl8thYPPd6CO+vuFZbfLTavp1af+fLkpEDVNaM+
BZ3fc6a6FuANId/ZqpBFEKCcJNljr99g4NFAbVhCDFuMMBSnnqdiRJHGvBXyxTP5
R+EkM+KUZJsyjSu+KrNDt7p7Xnj+zRissR2DvBYxGltJMKyrlkaE4MRsK3Yq6T9U
eeAWSZGj67NLesnp5dYgAvVt1GLYj5NyKWkzdunhdv9DDSBmUDC3QUYVfk6Ts5c4
yRf91YJWSK7yBbD0M3LOPcLLpfrX6f9QgKTFxmgqDW/US8nk53jBrHYl8kdhov+T
aO9J+6+BbMJki/egcMoZERlcpzryNTSsOnTVJN55J1yxhWBVJf8NgXLPnPHQk6Ab
rk+XvLXSpO68llzvMQz0mptnkLAofB9ZpPHCjspmUX/kQl4PYCSPLFbYy88uGf+k
6rl7xA3Ra33Oih6RVTui3R3ID/qJepHBTrzO//BPX2GhqOa1gUJ3N5CxIPke2uIO
FBUD9ENZjNH4AIyEdnA2AjhYzLlzfxMrk+QfyY7r8LtaWVwwdS235rkNnMb6jTIx
OF8DdCOWEYsNiP7BmQymzqCToYD1yN40QeVpQm0WXoANblWhp5ovqrg6njE+d0xV
Y/xXN61EPJ8a4ki3OFgfe2WPt2ZqNQDqHjmWPdWQu5DQjSo7VIjEdVHKix2RxgIy
FwflQLnMEtXbQI/Y30fitZY9i3kI3E3jojdmV9VKtvr/yW93w1wR8Du9Rr9uqJcc
zvznGHRtVKFDiL4w4nYeEhmPjtoBLF7p+mrv1Eb2/p7rGTTMfDvriIAy4cj390HW
ry8P7wabnHGrnQB547vsZOVNtevZFmK0jm3xTMKVmIWgbdVoEOmUjcEe6UnLQgsy
u6EUjOW90JMBf82ZL1dAhf6AwEWSrVDCC6mi4M9lXRqgScxm267OkL2CuzjyXicq
zs/MBqrW93UgLiPbLSr4HqHvkJMbVRNmPqs/VetKza0MACz++w3lniZtjfF/Ymfk
NJTWZJOMNlq4Y8k8bCM8rG0HkMGM1BYDjvCZ4e80HAyHzvfg0kL+PcTRHF0dkaTG
kI4qAwnrL3x3EWOq5kS6cyu6GpTIodYuRQabNhqZPdVDzz1IasBN5lQ+sDRCnZKV
AgB8zWz5bi9gjRR480o9hlj9RiGZWW+sbHQJTwPf1sNhCADsbcnBe4PiFk9RI3p6
Sn++8noudpVudTXMb6w8XEh1fW3/8NLldJT6uorfhC2YeLRGiE8FMGn+Gdb5bJrE
cmHKdKxia8+yQO3Awjzy48rnWvdU7s1lnN9ZY+Fr9CwrtfzQa2mekf6E+gqIHBkb
YlCWys1CYBjgyqvmEANrGq7YZRHzIaMZZ1C2YheH6ilw5/f3OD1hHRGPga4LBAc8
QuNbnj47df8QI28BFRzF4dNgrcOawAFGpP2LHAxD9FEoXnWaP/2fZDPxmj2kRMZu
ekg37O6txDmzms8ew5aDdupdlqNtDtMFrMnr+RHw7nsdQvykHMUNfbu4npvqEOmf
R70zaJ/l+CBOkYIDg2j87xwCkghXsMK/lju9Xsy9mQulJOoKDW485AN20HvKmXWl
PjJNrkRC8GohaK7pEsn/I2vx60FdAtvs/4Su+uIgLH6tcHf46R4oFBdcsjzqKem6
wOYp7NblYLuTU/OriUCHfpjYzBEWPTd5xt/fx6GXz5yBvYuhbRj9cp8PG48+7REg
E1G8dKnFK0fPZsuTINSW4RXucYc4y7q/7t0xEDQtQe0Ym+d8qjIsA2CRP0CmDTkp
EEcflGusYKnw1lgp4UqSSBbgtoVa7AP3KZo11GxcTgpFkUjBKZ8bRRLXlUeahGJz
7WmgZlaKR8SUObyQlWqZF26dOOibL+Q/SsM5sYX4TKIysEff0jEEeyadV9PZuqxF
IZBgFntoogqcd4+rULPhRoE72IrX0dTUMexvvR+E+esZpAekQcHT42PfQtCawS9+
sq1xfuwaJxOdPpKwwiviZ8fl6oE2f/W9npTdCoBtKLIMJVmbD/fn6MawE9likrEf
kV08QvRaKocpLB2aP3AI8v+npQvvpbBZkcc26X+j9xo6ourwjBx49fRN95GRQ0I9
kt+ksoTn0YLqC8qJEIr989qpkdGdNSUJ0LkPZhbFAoP8Fsrew2srdSnqcusJiHqm
2cWYI0Drkj8noE0PfgnqWyvN4JlOtZnOgsSeWuk0pTLKk+ZH/1j5ewN6XkrCJ2G7
lkmYvL6Kf3px5MQjAipeToQHioXenV2n3Ttb91GES79RWTj4VYW3zD2oNNvU2DQ3
65ZjVbQYSFUJiwNiwG6XvkuUnBNkEwZz/A6XaC4AjznE+J7aHfHpeiqp375YuZ+H
azz04WyrqsgQ+LAlAGc5JuY24LMwdhYnctnPuPXreUvmc9u3cB1EvRPHdEn4e3Pw
WocG5/FJTdzMwPqbf4/3KSfDi4udPKsVTVzMiFEzrQmH6qvjt2BVvzC1VCKnp8S5
c6Zb92ClTYxa2W12QEDT7nXPWY18GvMCzfvPd/xGCqrVs2wyWOFeQ4irS5R+EVw7
JurvgX10Nuv7Vdy9lj8+eqo+hxfnH1XlPRSOIpGCyiYtqhWtVYwKwvZgIxy7fZyq
TGziG6bJwZV+Ox78sTb/atuaRCp66T+8qoS912XHHXpEn6SZiduXGduiFn6VR3YX
HhrLUKS5VzT+TXuZY7T9puJJ6PnzEaG6ZpteKWhN7eYdMHg74lJKwlF8Q196x8Ed
sWzJRFFhzWAtOrzvagdLkZkJJ10vQlnUobq59YvQsyyY1xlSJe6Y4rUq4AFghWSa
N46VbNJ2XD0KBz+gOjNeoVoV5nEYhe2mngQEbn7b6CtQSM5v3OcuxoQfQ2YKdS1a
DlYv6qyVW/QlrYP48h+M4farA//eIeW3m/qE7FuVPeZyZo9iOUZRTKBcCyMLiME0
eLHSMAAgzjUSvOnIKXyy1MRM1+MY4j5jRVaMhP0nWtaI/035oUbHGjHEEwl5IAiv
BnVEEgmy+SLyqD7g6KxFVR4y1y4TIXzhFpS2fO3/mx7/2EbhSFLz2UI4GJCw1skh
ga9Iu7bAs2w4BPW4qtbm8E8ZFUDnGVkFNOHsLwXmeAXE9XPPScqBivsPk6xnel1Q
b9C5To0S/NXrSNYJ0JreCGrDwlFCuZ6/WTUP4mrIbvj3/us12FJbUi2u0eACtUSA
ONARUweTebbmHSZ3pexEdj9tbDJTuT7DyOCS3+uzUmino7QpmLJGx0kPeaPCL3i1
1L10r3+ZNeKqLdodsiMM5kBB0FDjW7EDYynskrPdJr9Uyk6nn9oiNU/5B3bRQyNN
9Jef0O0AZIgy5yUscLpDLlSrilVvZ+pF+0cPjc2gricj2jpWORn3/qGagoKNA/73
as7JozQv3PjrT5V4/d2N/GauPP06aakQNj+bo3/mQFijJa1Xp5VWaPlN2evjF2sX
ddDDShCKkMmpRkVyYQX0yb1rbmITd3FluBArXfjQFCjNdP0qBRTYut1gYbvMbId1
SkzG25x936lFZZ/ysnPvbB3QqJOLxj+eUeRgbnp5XZHrMgZ1c3J6vGtln3Geqdye
pGLALa8evjkxfASZh+YCWRAlZZCts+S6fC6JiAf/I//+PnT98tqRPsRbydB2l+1R
q2zB/0fO/ssG69Ei+m87xM3u2hdka8GNQ/7/fMOGVOhFywfAKbsW/G0QV/sBizse
mgDzlkB8Segv3hNI3butof444Nai95on42XpQEAzzwuF/hhBazttJeqqwq0fCtDM
8RIeMytqwaodjD4ynXDMv+09kn8uefF0bWVj6hhWHkp7NOeCXeZ89RnLyPlP44el
CD2hiXJ0UM5vBBf5pDuZ1r+3MLVdYGSV1vIyeWCDTxanYOmzIXRJ/nUmeiEOxykh
rmvMaMjxGymzVK15s0cJxAqBCH5PeYzizJvNmbLgs0OwQ56ZtyBA6zULLm9MTd+D
0XCKHCsFOdRwv4nXe7BftbK11eSWYnrwt/O8XplG8k1GOlQBdKMOXAqPXIaZMJck
Solo/pxRYAa0jEV1URM7Nx9cmdmJUhGavKIkg1KvFXAgcK/WOcnavn4m0BB1vi6g
GPF/tyhNNQZyfFCymgbBwdrneOVkgbLN0BRxHFlPU86Y7KwljTC/llOJwOYLMAO1
MZ9vzFu7jP+dMSS1hU/PGpN9/VPteEsOB5nsS5GgwNPAt2G1wuWdC9Vv2d95wuRI
P49nNxUG6rUes/WWH3DKr6giojcJocEj5sVWPsYuQ7WGHzzlWWpb+orMUp6kuwxT
62GaBm7HqB8SeiMA6JCmlgG0lojd9thl0+kobSJILSkiY6v2iSLcY+R88AWKNHFt
s4Knrfwzi1LFxetBOiXA7LB/cpC8sUfWtqWlDELRzCgBw9rrS3j3gw1QOkdWI3Od
ECA8Ac4PQ3OKBFoeL/WkGaJQg0wFrw6sYjllxHGDy9Hd/mEp6xu6i9lkPgAITP5T
JpByNbfGDX2Bph1nBKQF9RdUXeIM1kbj9T7crjgZBq7ZqwzH0t7MC3lRp/WAxPz+
ZNCshLDJZ5kaKTQcQ36Eprm+DcRYeOdcr4IkE3rhmbjPe6KuSCoohmmlR3wgBzks
Tjal91hAIHnPEOj2wZsIQiSZZG28mM3fLvpxqsL3X0Aq95DdcEBkCaA9vaUZuGLU
FxDkKqY3G4YBJItM60lVTm9RZVP8n2eN8giaOEhKXNYEXCjyKeXgTBYB7bmrNcCs
8V3dp9ghmXDR7IT/QS8UfYtZ7nnNYLEanprvwPvTkoXpuolDU7Ap6nm6MSMxrORi
nABdYhl6DXRCBwEm9hb/itg7guQLF0/lNc+VfTKK++4pYerXlEyNmoS9kshw7/9c
KIATc7iS1YTXLI0zX+e7k+kjcyq28AP3kToG/Xb1cumDya37n8j8VSTm+Sg1zvF3
nsTRe5gZ9V6Ap0I4aVRoyt4NZgDrYZyJpeEIi7CbPFw+b4TinIzks31WqA5f0Uja
ATAXxt0NqLeUDvqUROlCqPEob95dq0OmuKdAJW8zNs0SaD4tBW8q+6/3Qur8RxxD
Oc7wXd/DiM6d0plDdMDxwNRsg8HpZW54Xc0HLLgaMijTXTFxdD0suY5laEz5jcdB
7aocRZCMOPya95VhKWGFBk5zW7L1yYIXeGEFNUBd8ARWaa2/tuCbIdmsZkQJk9hm
fd+vnn0I9dcMZmqN2NuI4PwBWZbd9QU7PUidu/pJg638Hpaiu7loMicVqUKG56CY
e+bwj+68jJ9c/B/o7mkbmdlFz1H8YHJ1HMjilgot4ghrCtdbTUdTTbobvAPhKTYz
anUQs9EqQJtNP8mciTbNn93cp5XO6fdMj4Rq9j9eEe87dzPyuTNN/1PR2hSTsqRC
m0R0SW5435a9RtaZ3e1AKYlQYlSJvtAMC27Y+54xcOTYtC8r/7vIDPOlwIw/Sl/A
yJVJ+lWmN6ZZmcy6AJhgM7gSwTmL7jTriCvBz/hjT9xHya+mPIGB1XwJKfeyIEKO
5Ug3zwVZGWj3bg2Dahd7UmwqT+UvLuj0TAWO2PHAH+ByLkkA5qoxNZ0MzB0P8/Mm
JDXfgjZx0MxpvSNtHNMQpo9QAtHqQAn2dIYLLYtpDtOTzMA9ya5q6O1YjvqQl/Gl
yi7CKeBLeWalwEqn5KV2yr1fKy8iGOdOHx+E06BIRhOuCXaM5slVYKhT789R3miq
Y0BnrtDgabw9JcWJO62YJzZ3eYQQKjEVBlwcem64pbMyFJQ/1c40o0mdxP5vK41s
KrDJ70HeMG2YXnMjfkFAIo8mKcE8Mtew8LACBSmzwOiagj5d2fXRZctAg4U4oKRj
I/svGHu3G8fSJ554On6y0hS98I3wjJsHiZdLgu0e5k4pLzB2XJjD2jz7vlRzRdLf
iAi/36j8+ncKprxqYRDnsoRlgi97JsZ4UMT3yvhgOH8OmwVOgxF4PQGAmFUopVMI
mEw1gsRqsF/Cs9mC1OUgvjQ0ZsgXAshCxXYOu635A8yqmOujsSv474V3fmqDE0du
/HSXsHmKY/TxIyJyJYQmm13ru+4VIIPmR33zUMzWCmSeLXlV5YnU+hWVIZdXChGe
t1ofxS+vuFpsFmwhOgnLBR9EQpGXg+J/rkBfN0lDy+XUVLzT5NJ7cU7h2lS3JKey
nw+VWdrFJ9/tJJ36/hT6E3k8CM6T2K6929b7gx6Ngto0+KzZH3N0sn6nO349Cl4n
eNJw6YlQck+OkXc4kYpivq6tinuEbcnmIcv+xXdvWtbByFb5RnbKgfr9ZT7rDoR9
vt0EelLk77w3S4UKU46OtWCHHp98nP/bCZY3KasMN1WRBsamx8B5RTJGQNA4M+Rl
Ais4q6OXjnXTclfTv9SJZB2dPfS+/E5w7hptsYl3lYDnXclzOe9SKw7HOau32VAL
JfSTuQ9HSKUgM9zM1B3mAXiJn/LdAKkyJssZ4m/xUGJVyT/eWiDctYCi9DL6HZSN
QqVcY6ecQt/9hHirmQNR8TYSGDpANs7eZLIRmw6iCE/uVnCeRUqrSIUKzwi6nMKy
d52wlSZ1xRYNp9pUEC/hMslIIRJLzA7IGwYea/z07XBe5fnGAKwBLF08huojMkKg
l0hbUDNS74i/7C1QHVtXTwkWwTfQQ45kldV/JNSnd87yBlafsi9kKt51tM8fe/vc
MemdUiBR7ontRF+l8SU6Z0iFyeyudu6fQeVCNmUAFuocIpMTTXJiJbtenZhekhsd
TlV7ZZ6Kyig4G7EOfc8xsn/EQ/5iBMCu2WWKc5CL3JzM6Fn5RHqZF4yIVb1Xcwa6
soFn2LS3OY2ZSgWaHEsgesjVQSFrC9wOjsCHXf+xx4OJR8l7JSoXJdoNZkqs7FD/
hkRHCzoIuY4rD7yDvpao8LKfT6n1n3i/MqMAExcqgLgJx99QQRdvsObJzYPE6qOt
xWHaXtfEH/P2aTiiy2zzOE2yWB0EiZnRNR0rArcR3czmGKSl+V9HBP1J80JI+EYl
df5BEPfrPfZDkHN8OQurEDr5nNS6+iSVu3/9LZlx1h+sHTl0qzEl4Hy10SDK3fh6
JP+oI2vWKxj052dZJZTV7KbiTskhEjgc6/T+X6Swgz++Yms8TgCeEdlDklUR5geQ
R4PwAOacXJwT3ELZg//fU/kMcQ20cOxRblwU9iB4kOZktAVtGha5GnXG3ptlWLec
J5++sMWi9slb79A+cbzAokUWwe/MXBHQHYttDSoooDjgoQjy+l6FlzYQ5fmUIRoI
HT0qDISCG3KjIxOe/z+IHaFT9f0OVhm/YFBgDJvgx6nM4oTLNPhtXLr06kSELuTr
1v5zfWGOjV5jJjPbCZmlbb7JxVp+HvYXqI9hlKbgm9Icau/vNeYOuH/XPuAeEOAU
gNus+pw4BUjKwS+dnLYe5ImEeNTWPKA2L9+ZKWQA7X2t54PHqKJ+AeHEB5DZr9jt
K9Q5UPPd/bXcHmtF2vUe7O3EwKkQMG8OERrBI/3BU8ws2jWVmHdYv/gy6d5Q8ocU
MBnZLMGmFTRg+SZRTaM14MHrCAIwWg5hMr9FfJX0i35+Hgna0+14WFmoePT8i84W
cHA6r/4Gw1E6rbrHAQ7yD3zSfpMs6eeKFtPrfj4hSdiU5Dp1ob5IzCc1xBt4BvEq
yQcSVvDJP84aatLqXbMg/g8K1cCJ2Q/aqZI8UbdrcGSLcBoUgXLBO3ow6alFB1wQ
0KKzmd/vTPUDqPE6CCp5x2mir2rqt+pIJhhR3PIwxVxMsZYhs05ksbH8Jqq3rK6K
JNaMRo9J0QeXtprQzqe3k82O52XTkxaMuq8oioC8TJXFHDYdpDqg7xEVFraXMWwO
b/lECfPdhNK53FL7qGlYuQBC7xK0Fsh+owy/b1EerckD3r87nPCQ75hnP4fUmHvR
QcPN7DDTC2/h0l7SC/iviv350vqeDdCiesZcG1PJ7CkPjqG3gBicujZ9FlcKsvFu
j8pn3QeznGmzj44J9ldf+yWO5oPc9Bzr4ZE7O6DiOT0aYdWrNtWz7z/pXTw7nsrg
6rB4RGzWa4yNYT/fdXzb0W+ch3QKYhlNayU//RUkVbKBEeRcXAFHRt3tnDCjueXA
vD2oK0vT/NkBc+qoIeDbtLJvq6iJ4WovX0euv7JL/b3FDVk9Of4OnqM/hvFiGLjT
dJqwCLdbPMKi/d5hvaBPgnd5+h9SfJvohfkLwc1cFykwFy1eGTrLBbJ15FqdRDkj
5UCmGV9isMTD+9w5NrW6+CNKdXjAGY0a6m7E/ca2+CLe5gEVdiwSywP20dP/0UG3
9eNv9dPvOa2jGdG0M5VY/WfiD0GTYBbsKmRHJtmRraKeQn/wr2jF4oDU47LP7HMp
PvFsh9BY3T44G/+LQkyB4ugDmY5snAQeblJlbji53g7ytudEARxxrd14/xjtkyRu
tnJ79wuAdypoAuMIBTkNdnyQAC+A257Uo9lu2L8PVGYbZKjNFGR4o3DdQHqaA+iy
N5Kc6WZTGM0iuMddEdGyMQ6ixuOkT7TYd0HZ1PNXUOL2mmeZOPbwcBRH59e81ZP4
8fgjZPLU2aYtyXJRsXrKk9exuy+GJNhbb9ABBYKUfXD9t1XH3Yghz5Zv49VhrelH
1PnY/ssFmLdETGxEgrRRwrMYadPHswRYicGwOpY1OPy9Oiy8S7opWGrhABCCpIqO
cNF0iBFI/Gk6qmCQHEBtEbrfrPdL8+g1hOmi5iZT/OI7McYH3cAY7PcZLxDhXuVF
GEnXoB8Gq1GY/C92OMwAGpLeMhGdlnZ7KN3Ih3GlQwaF9SSMb+CUj12KaRNBggU9
HkMX1qU164Auah/ycXVhiidgD/x4DLVvBER6l58nMY1v5jW1xiEEEDEuNYIAWnNp
QGLPRxRlsNC/cfUAQ0c6Jq6s3aJf/RUThMIOy+OyssXLCsq8WuCWF+XPerOsVFd2
DWhuOeulzKZY17KKZa+1D3y7wVv/I8CCkNaROfns2NvQAYxGRdkwDsO5aEUm0l6g
HPUtVYRv1M9tbPb5jUZRtEzwJAm/raTCQZTGo4hlYwHO4CDJL7/If0hrYygIBtu4
qLHr1DenPQkr9+yXB64x9Cd8ePnWAWtqGP30NR6mRAqlRPoPZfZqftyGDJiEE8dT
WX8f2clKmRw+ctHOUcAoc3Z1yIUn9q9IvaeDFyBiTSSQmVoMw0fSkEtNveua5yoE
iEfoVObsailDYDsUBMwR0pNjJnlORhj0rSPVhz3/WkEC4rm4pDmrSMy9JA4hctfv
jiwn251eDuy69mZN9jbZyyTLBzRzM7KAYmsYdN5g+jc1iKrvLqd6VdUAkTrMLAZ2
pgKzQ17XJUdt2/mMDG4oKADrkDFRGe9RIf1fw/RF1yIxav8bgvL18QMx7Gmz/7eU
C+BQZiRA5bSkCWJwNHWh/kjDcWrm+yFUwVugSkOr4xsB981miA0VjwpGUCoA5QQB
4NyncvbDcAYlL3S/VHtkuXpzvwtJtaXSeLUQj4C0UQC71MKdrmnDgnCFhM2iH1HC
W70iD2f3UAkrqIGirzdaTg0p+WYY5Lcg9YVoAhyKRGhyY3qmXTcNgl0ilsxO3Xtq
pz++I/vcFNNw7cFc52dXHnOExkRw3QB1LKV4f1TL1jSTeqvANYRJiQfvfV3qUWOb
H0R8vdT5GheJckgCTnk2wHCI2vMoCJDaSOY5TVhRcg2OuDv8RPO2o9YFa71K9RYl
aYvo3jjMPrmzeHspWjC6mC/AwTVBqXSE9nFnYLlwwYq8YdJsywEF5IyIOOFgMLW1
Masr8RVDA6dllZ7OC0jqwrNhrukOc6C05ZMeF2PXbqo22032usWCo6mSRv6xcRTN
9xho5Xz4EwM5vC27djO9xbaofneFeX30afHGIjryTjcXqs+33EIpD01nmYchUQ44
IMz4y0FqoXwNw3P4/pAh/q+LGLI23ELfXBzs/frGz2V/Jw9d1OzG/kpEpIBxUBdu
VQ3mF44uayTe6vRliWQWgiVYYr0NfIc+I6EDdXOlFMjBbMR1KYYAY6OGvQa1uetZ
fk7XbTQ0OaJqNQy1Igr2Z/dA+EeM5FshHoB4QElRN7B/InDB/1L4qEVzkL0M8zh0
TTK/qTZwrVCne9i+hXUmODpDx9BMNKG081q+jgitvzzfobjPokHp/srabTi/7qvY
0XjBBqRo6bf2HPeO7msb+PqM7EOw6EWkhvF19ijTzZ9clCU8QEmYvZFXVKH98abx
wEmAz7L1e+xKhc8OHdkxc9MsmZmOtW3DOYZRSsQrdsXNuDKtB7eM2stiCiMivYr0
3Tp6Tno3AZ+ra6Y/5UiiNkamaMOMRuuqBpVHxdq4ri8QtJXRNOH/Mc08tBq/5c8c
fq2InfIbdmkiIgdjf5N0c9qSHfLnD7j2TD9uI5eFEPlcqEgQ6U57RXNkyNkQfXPj
bqwDv6YumBaq51d5N7S5hE9gYwmadYMajd5Sm1IELbC6yKKToB/3XmPBz+NkbYJD
bu3VlrC1JZM7/OMUM9KYI4zGNp7tfWlW8UWOIeE9R5xSMbYg3qb8wyfnb6wMfI+6
B1scv/MEYeSBjmCpiTsydzYYfZPnV4S3Vh1aqTt3UWBedXfw/XBmQompWWmqGpHB
3mHmC2sFhX8RqHdPIs0hDQGHNyxiE5ZWbmkroaiWMQk/7F8x/FhDbL9WZv+yvTxc
v86Iu/calX1ayp7VMvjSq0vQcSQsmY7XqLqp/eWODOEO8g2LKGifaWEN6PkODgAH
86EUDOJf5k1167cHjVjvblUzxXr1Cd0ai3JcIfOqVj9F124aAboxBP1GjaD1wxWq
vfto4otpiXf4WAVZPlphSgUEMZt7y6SxSpNb9k04Eb+g+nxEN+5/9gegB2Sg6EA6
aEA+ehzcVDdWm6fxSXPfHRc17FIjLOjElpPzAFGGEXEA+Y8VnWGvR/eLdWDS7X8u
2IpJSUeo6k9UH70AG8cp124afsrxSyW3yUv15kNoVsrgAcCmItKhflVUlGf1sQpL
QdOM7UVDQFWzZqlbBlx8U9nndg3AQOPFnsezsgp+IoBh2fdSoaCfThaMr8pTb0gB
XDL+1VfQ91wS7HeBNWq293W8gX0dSQEx4Icw1Nz3OIBzBjKGoqD4UDDe9TtPi1F9
3g16Lde7xz400D9tztKSnGV7effAOkODZpjgg0z1TI6vJMQVIO+K5ot7EIewHthq
L+wvkETegs3M7kv1qgORuQEdRo1/Vds2aqFwrrU2iwrS4FcqhvAzcgfCgSQU9Hn1
kDL0EXyb+KNGFAT5RTcxXakIjrtKFdRCm5abHIYQrMaQB3e04RFucXu4o0Q+zdXg
k6xql8yBz3CDgashwKqFDiwEcjPzeqNLLiQggsn0OxYPf9G66u6LmbmWV91f8/Qm
qTIFNPeHNtaq25disCQS3KVeN6RioUCxfjNz74scrMn2jRW620crd6yjLeR1GCLw
oOwOvg3O7W8DIIdBNeneYac8Nr4XgcQ6xvCi5TXoYVV83EFNXDkdWPaWF9TYygBJ
wETXIBNlLZVXznalTTYAkNxHBywaHAucpSYk/qU8VQ85+ahGk6KCUB9eedKkdLjP
veSR47KU2hWnfqvS90At5mPlI/xGRwOirtLAK9SdU6dDSwGmtJbOBdYkrLTRugkB
Yimv+Pizhcz43wq76grhzwB2eLPGKCNF11qvKG1z1ia4PDDSa80d7RDKkzt1Hh7d
kWmEzO0t1ZklYGFiaPmhg+fWGkWS3mHL851RAF7GMy6qzWrMnZXX1TZl+98Kg7cq
SCkul7DojsTFqtA/Yl7VIqODkcKCpBFQlSsvpx5YCyNBr0h1XEjGOScw8XkJLDIh
nM1jCD8JEdDYReem0ej8ZH85cLC942ZaThQepw1DrTSQWorOx9ut+gMGd7bZ74+r
U11KDZxxmpLhirQZxcdN5fGbZ+/woPuub+At4Ny6DcBGzm/QLnNRXUuQhy9FHPjJ
QhxR61xMpEAKhtH7YRSMSqnYGvlbpcPFmgK32llGSuqMn5h5IV0ueo8uVvt69yHm
zVGFYr63V3dK7auvlcJfzfb2kPUw60+l9+qIu6z2sDj/1KAHB6TdpgcVSGDuYtc4
bxOITqDWkfb+URMEbFRaEk1y8h7LUvK6xDYPs0uWkaK0UWmWMwlF4tIrao6LcdHD
TAJnVUNhguPLQBhMecf8cg/UEfCyKTQknl7U6F3iWWm0TjOFA7eutZsCV04der9H
1rkZRgXT/icIQkreHVtQ0g99YLyiqL966f9tHMQ1BTOkGEiOtZvwtSf6tkzHiDBe
3Lkdsvg4YPzaExzMKg9dCq8Rfuf8YEgzfulTa1YJtlzCTylfpg7Xh1+mYpWeIymO
UG2MmoVCuKWdtelZmkV1P8CZgb/O8Puow0zNsXSApitXJm+UhCanPw3SDMuiDpE3
r+yV4w8i0iZPccdiGw7RX8BKBsqJ8bK/47K3h7ehfta4qjXlP+J0ZmnGkAHy7spN
0I1h5YATrGEvAp4CBC6pRbyhZo2f+IGCQxjw5HIwn22qPeO8I9fd4KGDZcAGl0bA
FmxBIyyAwGtiTLnx24Eov1a90aIrC7ZGMIiqpY0xbLWPzy0WlLqGaluaXHGZTFKq
b1aHzjY0qHJqNVY4yp3X/c3SEOU4tPvwMAdY4pP7cyycqmwCLryiuibu+N3P98O/
9p8BxiFvwPfCqrtmzW5eVP4VlpcApFLD/UvZQ4qYIcA4t3DzvhUdkSxYddClrIiQ
L+QkmR6QdXU8SNCejgdBPN5bhtrvtm8vbFTIBXRnxhBvNlcEAMPN2KwzChk+rVYB
dIpPXc9Gm+W2MRTTed8lQdL08rkJ5sn+tafTSbshxn4LoxH9mKA6VABEOqzXTj0i
J2AHVRIC629mNODamMTSQ6Dm0+zlxV3TKOn8zGTpC3buTcfZ6jZncupljJgsEdLf
TSee33fgc6cOTNQxjSVLNQkB+kNr4FtQcPCOMqaIDq1UDzJ7yxZThcjsuwKpNCm4
tGkHvLzGjAP5RhoGURWmZtUNb/1FUSVhLt8nzBw78hGHHAghKl4WDI8gjzZD954w
2Rk/svHLS6QfviMEIAkpYgO/n1QG6VDA9dkqZu8eisWM5lOR/Kt7ijv4dqjktU6c
K38O62+21Hjj/3HyzCSlXTDeulKXO1t2GfCwzFe4Rrt2KFcXRhh8pZT1cecGJWom
HOLQZwXEZBvL83c1BwTNEgzkVzwh/tuFRSx5/vAilRO6btc/L+Wxs+WeQYc72qaw
5GT4OocsuVIcGa4G+thWelFsufBiqLocOAfcq8ZU9IXJQ4gCV2UPivBEottjh4OF
Ji5JBKL5n6P+h+gzKaPDBgBlaum/X/+r3FjfVF7NtXnCQHjdKp8/TuKzQ4Ty6pVS
8MYxYas+NGWkDUYp4GBMhQm6QEjoP5V3n29XFjUIkpk7Dno+KrtZjcRV8AYFLHyK
tlgoJ03M7pwhkbHCbhjHfLfbLILQlADIauHwPpU1X0B5glOZxpnSeEt55BgHipTN
S275t8Q2TMEpwQCQ2r3VuFMLjH/h2hIGXZeSggfeMSHBGxhgueAT+1jlLmSOe4IO
Vtex7dd8HnTls1WXqVzJqwZgYTzqHmsU6V4pBfK+BGUTrILA1P5f6ukG12OcGYNg
eRvEnbKRnw9DGdU9t/VFCa+YP2EnGeewCGlUvuSijJe9MyevqsNpi2hBll8ZLzqT
WvI2XbF5rF86saA2XMnaCcgseFhhyr/uwZx/fdCny6jAzPQcB2Dk3i/4jM34pi33
V49YzRCW0jh0uY8Vs28fjWz/894vFzTGDaa5Z5XZtestlqCvUqOKtWGJHcIgo5BV
A6ag7kQj6Gs6b72VaquuBiCzzUt3wyw6k+EXQLwtG87JlCTysDEZHOEFRL/bj3nq
BFf4dWWCxJKmjQX3KZYKiiU2+CjoXCtWPkpziX7wP6LyEoupF/mhNqlcatfLyM6C
H7qWIl9NuiETuOVDqj6Txupr7wk5UioCRqEdMzOUbBkSoIdSSRhmlX1hURwRDY6o
8DC6jDsU3m3ShjzpMA+ILDKSchmGTugCT3sgmlSzQQiT768m5NK0rXGvoj/oNibA
Dh0Kq9S+lSbNI8YaWLVSFvMHDObSs2CCnbQ/O//bmPNLM3W/oGAyfws6Ox3+SH1t
d5PnyFLo/5DRUryLKAjyFFbk60vE2O1XBrb4D6GUcE7Af8VLnF3naycl7kLnw1Lo
XBuqPoQsOJGnk6KE8K/RXG8S2/EatBr2tRxNrwZMoWlh4kdzOAazoEtSOCuikHG0
Lh9uVsOcMtsbHzw2p3k24VOIE6Qfl0no4aa9Is3URemCRP08wO+6952WjO3BV3YD
mnA6SWyXIGIyhf/Psnch/vRTsvc5uQ2OxQmkCxNxvO5fnVbQlJojby5TQq1bs7YT
rOUwYFi1ptP7gKgZhB73myetlmoS/OUcOD4VZ8Qhgp5dqU1fWlnxl6e4eMwJrdAF
ke3t7hK+f/i+Auq/mJ+a+A8GhDwN0uXXkb8OyX50sJ+00Q5pVYghuHDd/nnP6f6C
jy2eQDexTj/u6T++xmBKE7v6RJ5bLGC+GpILPvDccj2Ej2RwhAe8gtfarBWltMXn
jc7L242C/e96EHAljYsLns+s4gUI2c2Qzr75XWats72DTDETqJEronW06PSwt22o
HM5YnysCsSHBZ0FZXtfiRnCB2xmH1gNHrfOwfiJs/bsUEiSNQ17vqvGmZ3QlMSqe
elC3T1a9LSOD1PQXjU2Vw86WBR97KSA4nlZzi+FiUCbg0r6vJSHB7I4+HGdPFbbg
fv4Ka/oEgxGgj832BWZoh3Nc8PY7LlwY7xe7TxZa9TzfKC8FqoRFYnLmnhFR1Eas
FLxCZ9Jqfwtkr2DIID2T71VZp0ojVCXRA3ChgodXPJwkiz4FMrGs1cs0Z7j8wbII
nhnqn5Ojstmt74zf9hEVB0xTU2a91a1qG7T4HxeIHfiCt36vqAIUD+3Kebf/UHAn
qoW8uLqOwS6lccNcjopwvainEPp8u5t3i4p28pspSIxGZn99UJl7aH8M5h5KiIed
qlYVKDZt0TloSpYpWc/FslGkSwAKCEXj2PoLAejp0Gy9fDjdJADxXK7b+AC0s8uD
mXJW0zlXrSbnjqrUWaBVGPfqo18AzRlXAoZUD4jPmVznxnpqPRjhG7ODc4hH8m3p
ItIlKqkJp7rR7RwxvKgmhdXWKDwBp7S6xChEbtAjNBx9O7kSljLV9VYHI1ZO6acs
XVgFAMNWYbEjWYniRHhDWoNwqUOu17UYnz77WSLfGIH4FuBv37b+znA0NqOPbYBp
iRdyyTonIWta6W4/kzEa62kgXWl1H0uX+nYwD2B393CVWjAvDeC5RmA9w/ZWd1jR
HWkVRrH+RDFnjmNNTspDwcECUVtyMkv+qX6bOrcCVTUq/mwEV8DHJSDp8idm8oBU
T0TyX7VBV/heXVOYy67g60tDKoWQTG7u9YkCxPgINJl9DGKVEeI8o7fRZ7D/qbY4
ulT+3yRjaTxZ1W7nuLq7RdxIhnawBW/eXeYqyPhUliN6HCy2vDFP2Qj8uP2MN6GV
Ct1lYpP4vOh14d2/F8+hQ3vIq9oOT+FAAnmJhC5f0NE9DVeH02id8hkuZTYQIZLB
tzqWOt7CbARFeqSKcoKkpLj2Vk/aPPgrpt/P8hWWkoafn+sqxP3Dxu08ArmE3ZCw
EQ0AsGL5K5gU3bYOAkI1rbaiGNCAUWi5SMHzEQCkdX7TNV2ZEdEU4fP61Eqj3pLc
z8Dfia7q3M12ecxMcEzZPS0bJiLGRFWq9jqZDNdOhY735PliEZ4zSp2eEABEWp0i
aq9tmxFi6BV8U35Biu+YLcl3DA3x0D9Pg4l7C1KGkxTFnA5ChF2rOsU1lTEAgZbi
d5QXE7CkW1TC7SgaNiG/gKsCcnLWAGMtEpyh5tZp/bkosnhGDM4tam2oshkUPwfm
VgMq8DOQbSnobGYUtqZn8oEmjCGypv59w/vBSK2O0muTKEMa8Chy8FdtXNXcQjK8
wxBRZz0Cec6aVrhcN5CNbvxlMpm1IKJVYIKE6c3tTR4MaJn3b3GvsxVJHPLIvWib
2YHdxClYunclFV/92io9tleoiOWqt3zS+0XUuacsg0023XzRo8w9kcNZ+b+jxnXK
UpAZr4ZocZn/OEVeDGorNOlskQu+ILtO+zJ8FNeb+nY7nIBk7t6lxljHgc+KrfF3
ZuEEnHPDa1Ei+/8kLVQraBGIcOQljppYhLdFba87hPoa6e52VltLwFpa06TAaeVb
pT8lFAQsuHkLyGWXukPHJkODCycmqcKud88liutYV5Jiht3nkZtcLUg5yQ/Dt/n6
wxt4k3rcBg2MuDv1PDJnSt09m2NIT0OJUYbJuTuwMgVs1UHzWqqfusObfwLI4qSp
svMYoVwHBH9Mm5fkILiwyKCG6ES9BEjdc9CwGR/UQov2UotHZp/4Vq049gYD5sde
wXVFUEfzX8rqLwzs6+eln4wta1VpA4btB5F7WGe2LT7Q4SLxI8tboUYkh5pp25Ek
fMsNGDQQF6NKuaUUJq6U4fxBh83DjTTpy8M1TGNvrrJTrRRVmNOxTC8evlThl/8/
B/DUhx1vVF28goi6YWe6dE+d3a2N4fgIDRk46YRKI30qA4ipPlq5Gf/6nVP6FD4e
AP/kihuM77L/pwxBmBrYsI5Lh1rZJCO4whRBsM57DdPZ5DQ98cywW/YUGHEPb8iy
9At7ttj6bS0qAY7IY+ReM5k1zkK4htQ+zi+VrRqtjI+5okAC54jLaHQYTOHbBfXd
6MsbNp722JXJ5Ke8MzKUvA4Kg1Yujv2ZabKMmJSno5bSHXD/lAe31MYBf0avEq/Z
zu16ugRW3MCjyVVSgJClN1uQxWf0yOKfQf8EMjH37DzQSMfzsYNMgdRA8FyXRVEN
7z0LCyJ8Zz0VZYWNBrm2bKt8rGEt9oZ5ZQvoPTO3dzQmFm2R1HJKkeYWlYbyk5/o
jaZxVNYLDg+z2GmUU6WwqNTlHKCEuEYlbK7Obyo3pVkitugNBbPGuF7Mmity/vox
LiXyfBhiQwwt2ZT9kfjhv/uMwexJzjI2GU5fM8ZlhzyfQRBx884b06A5Rtifz5Tu
4LPCFVPaWTUSfXGruA9xEwo7ClpIHu8ceH9Sv2l75xJs/jpg2e+ZUMAEw2mqfcrR
0A5wB77QURCGYopl6RP/zWx0NY8V+qdE3dCAEJPEZ36x/vYC45Mu2RucHK0tLaFn
pG4CHMiSeJB9BS/ieo5fI+N2Iw1KGfmISc0I+6kXAUcdzVhMkaM8TGQptyVlAWbr
rqD3xBBevH0c3ILM6yK9MIJj/DSRyi5cgYBhJZyawXyncm3uJY9MZS54+LWq6Ldu
uYk1XYBagGgxKMHpYdJRsUtxsmHJIjHiCODQA4NDkTzsybVT7vbI5lEWuKB/DEZA
I551D6bED0kIAcfxxvfTeLzlKPbRjRVDi9DIv5PmJjx3PV3b2yY/8m/LZpUa3QwO
9JRuxXH5LDsoMd+5hMtWR2Ma0mPJbJNsmTGD6swWCIcYVO/Dq3UnIA5ARxvpQit6
OB+b0OC9FvF/6/8uzLLcFMxfqLnh1CjDAkzxTPi6YVDpofC29u6k1kL55634P+Y1
ZSXutIZ9sKs37zxlcIQo9LG3wVSAiLWVstjZviYU2Z5neyY6kY28eNkV2k0HqqCC
LNeSnJm/Gjo24BwTkziPMnt+LyhAgBKMgJws3BKLC8ufPD6gePFbbAIV0bn3uvIB
jCkpaC3J5Q4K8YjoVTdrHKM3pxEN9B8sN1DPReNwGJ6mDM2oARKPkgyeem9TAISJ
RiX2uasZuS4jkmN/LGrnZDJOjJs2gZ/GnzhzE0c4qcIGcvuzoxYnJHSWYzwvrxlD
NOA+UJLyFVw7jFPAt8AJwMbRsi2Z6jPDnLJ8kOZ2vXm6mrrSb7r8/PoPemiapuC+
lt53Hfzbsqszmf9GIXQEbLYBXbbVmldPqeSiNgq+fkr+zD8BR95i+l2TNumAX0XH
W2+X7mfS+F8zeMS92Th8U8tihj0T19xsoAZrU9Io4hTNt5l1QiSyXrS/OP72eY2I
qRzw+MamPh7STpxzx/cxUA81uw2j446Ijg4O+oC7NVovVvPGqD5WcnXBx/yhfRfs
qyZMduBkf/dvecDZ6Ne34WKrGM8yv6eZE/MK4cuShAkGt/ryvtrcwkZJl/+Mfibc
+JWttrBZ/hmMbHImOE72IrYfWLgoI7LZUJ+E/65cvm58I8kJjHIucV/QD2aIcZ/h
IpLiLnn2ZLnVB/Uei0RumD+SERgH1a45dq1usSL5OHPtnuAjT+3DDFXrNHAoHn+u
Uk+mf4EEDDWOXP1Tf1mpmT1WvfPCW4FakZZRD4H6BEuMymbrObKXtZ4apImPyhUF
oPoE2CFwbLd7MB2uy0TiRTABrW1yZOt+oe1Zc7fqBRFAzrI4jgI7bBd26hv0sSrB
2hY2NAou1p+PHNhAxr1oQIFzFjAKmyzbrf/uOhh1Pok5nNmxEWdcianoO3mSQcLD
pItWf6jIlp/g1gF4qOb8/Gapx6MzQ7jJ2c1yt0Bbu8oamh1bq3octNXU9c92yuZ2
A18EUOxVlGKhEg7311Nc+8YD4mj21w7q+c1tOb4N9xmWaZcHugkdZ4GAIImpzwUc
Gys+DnuE7zHcC6/+S8SkI5E/6Rhr2Lymk0t5J8GYEM2i8ruZa9nWW3B2o8JsLIdb
A2MqM+OlsUKjxZrTKrqDp/m4tmVh3O2qoRF6x80P8e2vgAcM7u5fA9qen8sAwubf
PwTzLAh1fW8pJumgI3FK7G03Ow3T3EbsdhV7jBbxRy7Kol3j2Xhx1PW9Agb5BSxd
yo9DxIdTQjPjhCOGv+JDWeVJpt1CGsRuVGVwuFd6HEbxyqjYTOUjbYlmIUSBIVEf
NcCP4T7EUhBzRgKxZHziVXAiwduM6Ur4Px7ow6cHcrDsz1G0/gcphz9scg4i12Y+
k1Dtq2AlDehlmK67acTAs+ow4Owbmkq2ZFT9OyWyqHMWacfzo8I7uWTFovhGvbYD
nxKLYxeP7TIA4/hzcGTvavRQxKBTDWRoOVaZ+/KHK5O+P5bZfKUpPxVAK/foljxq
5zHU7WM3cxrIR8X3jOgupGD4+C5NZG01FCw8RC+x6g/X1Eqh38X4Xls41Aixur+t
zuoSzWtXOAIZGOsdC+bTLTE8mi6HxK1MzSN6Q7VPn6TjuCqqU1GUn6SRZNEKECjX
PD3dL+10JbEOGl9mL3SrX2ku2xwl4dix8mm30yE1t7Og9G4U24z83U1qmhyt3WE5
21WZfVnNyriAyz93m9Jpn8mCs7Oy+dLPkp7QAatjpBwPHBsl9zX9hrF9HsfZemyY
5+Y77D0e9vTHGU5XYzN4nW0twE3xIDWYcYV/nfPynq7vhn7Cb7lpKrSruvLPsVYF
s0A/zw+4lwQfCCvGYVyenZV5fXLPM70o7yzEvjlPFoekyKLCdQjcdmzLyIpoXszY
m2PCn4Kg6km82U7P2LXBdjwLP2jJJupBd9tp8baKvKvtF5zLDdFRSRDmryg7ijNu
vjeJS5f7y6/+29q1X+45RbQxoyXjHnVZsm8Y4F/B37kfz2VfQrBbebWj8DGzpIuj
a7xmEt13I7JKN66yResOtMGfyjWPYltmUD0YhG5dMtuNo2nS3dK/odoAL+bOvmOm
0sy9DIkFCbjke8R98Ucy0haj4Rrp+Ibk8Nt9WoRmRK7mwI1ixE/Yor5vw6BnLgpx
TH4ewaKJfLwESox5bbg8/XTuBz8Q6XI2xbxGwL0RACAB9z1ujCKqfdOat96fNFvu
1klsgF6uMCstXg6otgTgeUsiw1YEw4NQqA7qJR9r6ozG5YLuy66htBLRk0VHBlgf
rfPCKaUX3MNXzJHf4jVrqpSJb+VSt1Kqj8PYZ00K99AIor7pjTY6lgz32Vn1bhPd
hx5mEHs2GMfSg3d2PZ9WWR0JruwLw8Ye9oE6p7nqxqxLevqMt1IVzxvExPUYG0Wm
FiFr08ZlmLxeFxR2chDBMZ+UmemKvgq3ZsXEzBSY8VpaVwnpddQVukFJ04ddE5AX
wZykjbYtDvTbSEXaETaSCi4MvMuYk4fK3HGwjv0nP1AIoSXR+TwIozARgBXWpU/o
tktYmCA5nSbHpSdw4a/S8RTeirtg58FcvGUpgckq+d8O0NOTjgq77YBx/p6JKUK+
3Mrz4NGtS6Z93S2n8gD/sJApQUrXjxI9r/tgInh3ZBQ437ri1iuN5dO+SeLc0/Ba
/nEPdz0b8Z4V8R7LIZertjmIfInJec4KbcnkQ3VGzqP0+OsaUk0qN9nkjFLmOjSb
ag4Jm+v+H6wCaa2rXOZafMf33e+QriU2qPjqH60CY6tKlpfEeM3HSE1g0vFONZpI
9dMUewOcxBW8IUoNW2bCQumIjrJFiq7lPRpqhVe89WfCo1ixBKy+zlqsD+21NYrO
LCARaTFqM2FwaUmmZmMlxRxEGFHDEh2bd+9gFEKbqps/XMGGSeOIr6jm1skQAzQU
lcDJp5Rob7+WzyPL1SfHx0lFqMUFW6qKYqs82X+iQ+gYfrVmBAbotFeI/HjmNl7N
VNHqbSq/8E2C8cAhLXN3pdgCpfcH/c/T8j2OJ0vakrNdHDe5PoOvimJWnc4gJKVL
EjMkJ/r1moQZDA5D12XuidYLTrzbiWJkMFv9iIpT0RlhL7oL1+Fo0fq8RHVPhhzT
CQT8ZUZnAQbcZ5TsaUb/sEURfBjqP0Zqe/OUKi4Z3n9muVcsbBnsXJYCZryywbyf
jI1P1GDcXPQB7aMBeWGwO+sDY0LlsedEBMG/CFLpvC0gTa28kYMITeMQySRGhCqf
aqo1pzztNgND3utY/ByoLI5lWjien1DFttA0pytbssGf7AOKN5ZXq4VktErTlQQn
1VgOFLqObj/LbAk8MDyE1Prtrj3HWkMHIsOCRstC0Et1GfcOftmGgVaLf4ojuuyw
Ut8CYQBaIyPlYdJr+RO7J/3XsLXDDMDy8YhpIWogHn501MMAWG7D/BwKqy34T6WQ
XHeSyv1/nC7QHMF6egFtTq/qgtBYGiho9ZrRR2BNe1Ff4HefZjXmqcOh5ac/z2B3
DdQ9VelB7YdadJ/aclGsfDZk0uI6vj/AZBOtoD5q0l0MSodC4iOJhLew/j21Bg0K
EJ3ZsnA+m6ma3b5CH/4OjddbU6RALEtZnTauXKYrmPrrvDW3pMuOvrj25LSnOEEQ
JUst0NLj8xuBeX6ig/IbI59gQpY0FLptQNAof+v5FiTbGtLI+o5Qo6XHgfCLZlaU
K+UTQ3SeFdBBGbytIwSAew7iSAMt264MzHjKEvFiaTjDwctO5dyEMZzkkXbGzqnu
47qPxRDJr3I2xbFWTGBFwxtiEm4knkFzzRN4DOvVpDyHabLtsPjC0aWzqlScBvY+
g5Fn8aPtwmgux6eQDwxx9aVROP99l5eqmJpA5n9TdYQN/wmO3NnAkLN3HgdONqdi
fmLuXh30QILge43i+fl+4nDPZhiwjoLuoNa0joGYeKCGxW0B4Z3MZ6bfeJJeJ27c
ukPOPjECkOJfrLwjpexbH8hRqswnbetvMJ/GOUVqPFByS6XKsIJ7nOceQVlDMo1A
Q8ZZpjRd9oz2FPxXyygl2YCFgHkhQNo6KVNeyTpxS9eNGCd5FSF7Sq+R7Fnk6ww0
v/ZtoRPqVc1QyWX64K3dZiaDmTe8ulVvt7rzqeXAYtK2o3u+BDXIrFLW+2eobRmD
Uzl+3I9FiLEqT803/XKCoMi+8HV6wmjG9W5f8QaSSeIJQ2sN5Szy8Lc65+SonbPO
R+7uPNAfqOnkDTr1xVaN/RC97c9BuHEv1KbhfMmMaAF9vr7FRdnzm/3uVZmOVCOB
jpHKMBC6f31tZvs0nK99al/biyQxGt8yGeL+WqqAS0/G01oYPfOG1VqddpFFP+LQ
yMu1SZ+oJM6tJT/+esQFhm2XpmUTLsvSNgMPALmq/fabaeU6oa7uATwXr7zBSYuS
c2OY1auk+OqIUAK470HUegYFkZ10usPnGfd42IcQzGTW32BDPU1iXzX+lZhBPrua
kOyKSq8hm0B1r3ZQNl1cFJxZNE+UAbTwQoFSAw58DWJDvRRt0pa4sm5ANamspOvv
/KvttwwKuRLXSXTsGLppCRyFCO9+UoWeBE1+bBWLQcuNGllviGOgECZWOf5TgSrF
cb11S6z46oR5kR8EDCIU8zKGI5HQ8CULM+176UOSa8yCJqadDFgk2/cCIBBMPRZy
XvbI/Rb4yPLyuk9t/DBCwN+hwlydGW9FhlMXtU7DoYYqGm8sjHnk0U9+VPlwRHri
dfnYdV0tEzcYaF5bMY0CkfDxKYF1KUrdxbz7HmWv+s/jTyJfSsd2diFyZ9e2Io+X
WOO/K/q7Z5kb/Q4a3hLei6Y8KXkRfINj78KALvyOk1du7bjdqVgIXHbAhzteqQWX
Fsolnr6BPdbCLHUfHWKVfatMkoNfY8dGgZ191mJxRZefKvB/G92FPNu26UQyoyys
RJA2hlYgoId4YMkyXcPyftssH8TVHPvcYUnTOg5+DAAhtzpp2C1LGG0cD3PyP5Ny
4qguB7ROeZD1PuGu9daeHCWzWeY/o5OLxQ13d/SnvjEH/e9T6SA7tzWLd92fjixd
9bAVgxzo8uCsc3UOgcbeWjXTnfX9eBtNiP13u1bL95XoXb4TOojy3kYJlHlCsZXz
RmvQbJ7c71p5arFGfrE7wFOAOOSpi4xMj5IDE+MrMlTpCqcvzTs2+jn38BZIpMDN
vYeO/R25rNbbE2erMb0Th0g7gBWoodH6k8wRt4XVhhDBb8SmNDGg2Kdnqpj7OHQl
Y3KCAm3vapczxTgd2NlCEmywdC0vqZmTTqQH0pXhb5L2yUe8fRR5yZWiwGEkUhDk
Djcxs99VdbyAbbv/ulTPeWRAVCVpYAxSiJYWFnleg8B/FTVRizMQFl6ML89heTe/
vFSjyBBpoF+tX4XbDFfVoqLPmC9sbsZc0eWL+Hzas5fh037Cdmy/4ivOTkT0Vppf
fJPS2m/BraIDL1l6ETJgRBH0O3VSixWP7FMc06YpRnBEdxVi7M5oeYgnkH/Gi8K4
aXwFmjsRKkxvHNPlCAz8w0HC85EK3Oc8nCCVFnxcV+TKnBmJBPt247mr5ioCs2QB
jKf9Mt9JtH4LZkf9Xa3LT7ZFWuNks3Fj1YwV5CjHeJJePs/hZPQNucKBziBmpNl/
Sk+beDInwZEBQrUiRVn/dDRU7Qs4KC11+NESWyN/RHsIhMWhOMPaj2juu5f9rqsO
sdX0JCc/QOnNpKE/WG6vwtWQPtZgPRuGehhL7Sdn2MMCdZdDCiGqzzXpvysYOSE+
kSoxJjTPDw/ppNq1kSPefow93K8B7eotmmqnS8G0L5mQZf06Oj/ZyqnxrVYt8App
Vbpu0rzpSAFILOKA340U8N/JaYYwYpo/Q3v5P7Oighb6T0ueRKm77aTrJEX7oK3O
rQaaCrmgjSSdI4Fj2k/dfvTxS0gAy1aOChIAYf6mWoivomBxK+zh/CK0J2fID4ax
hQWDxuhmBfYxrkVkMXftq/v9QkcQyp4tu3OOSfYtCK9QBauc8LvpLVsuKsdp52O/
s7Ramk3g4fHG3B5jLDJcVa2gCUVBmi791WCuacZPV2wUB47if0Slvr+wYUdAcGlk
Bg/k9t9fzT29YNdblc1PA4yUbqitIjbbzdjYmgVgdW1wsv1mwbSe4QATpz60Dya0
NOpGOYGD5Pm/jauq566dGzuqSy/wRbz1ZScjzKKiRqHvHDNXZhxY7hGRIZ8qCFd5
4MpmFDDTVKmdAsYy9meyNFInF0rC9KQIneTHuHTmuzZGHN1jBSeS6DAp9f5EzFKU
jk/iTLHblSWggwIZw1gQi20Ef0zZzG5NXvfwoE4Jaz+ksZj3/ZQGh3vgIEQvKB/q
ZzmyNy8oTOIgGf2/AGhKQsjRo8zVrKmsdMDfyZ/oM0LVpdvnPT+9mzHjdXQ7/zXV
IOUb2TgOyeCd00ORMG5q+AA9emOP8jlOfFIYjlaEjbi9j5veP3MI9vTuHaJDjFFO
dbtgViZaT/3vwqK//1W1afU6s0hPj//gYy/2zzhx9lrADkGpxlnAaaVTsIkJj5Uf
4rIzHVFIkrYYc1FCFKOztj9KdKnNj9P5cOc4AYnYdrDHdBmIYCkDqYYrfP3v/inV
795t1NXzZBBUoEknA93GSw6kdBTSlHX5faT/AbcL+ZZBov/a+ZS3DA/i5i11jcM4
uK5/RO6w0k0pTCGWWHAeIQn22krP3z/YZBXuXePvST5MApB1Iat2uEhSbQtyJFhn
4NGjzBEYRbVNLCbW2pY6nsrpA1VpkodUtQElIUWrCGDGZxXRERgVJyw9AeUhvCZZ
m3UxwUq1aO46xygRHku2v6ATzhYG27udhky9gqd64HXcPC+FFQRD/Jd/sqqyF9Zo
4793OSbiUBcNfXhDYP45THDJ5yKvlCVWgaQYqK4J4d87NL7EGVmhoF24wOT7YBa8
NbLl+e+63/zP306OjHZlT8KN9owIG+hFm+Yt3NNEUHW8lrAOK6ZCqtGnUoHuFV/g
qRQn+2Z7WR1TVO/2hZN0XU2JKlhxXxX5bzNj0vvIgZMv+2bTS1jUck/TvZB93TUb
MJepfsiU4FajjFqjuT70QUnlbt/MEOSOq4CJhBGBCUCWtvkm1mq2z4iyatM5WRr/
0YVn/0EpnHNUzlXPvOQsVaWxO4cbSo8lmguDKjcNUgXqb4p1v1YrVyACBlrDgBp2
3jOKrDW2eCJi8qlg9tKAmO9AO+b2jc2zfcgtKAzpTjZdo3hcPEZK6oaBhfTTudnE
iIGgK9mtwKAdv07DbflzL36IbKwk68+eIHKuZAGo08RJixjAAvG+bu6wn2zdhtBJ
wfTrG0JQtpmNfVZpNY+pRovLtUPELT8x5LiCVii/kxwy27vTAjbyNU0zQBhXCmOQ
zoz5d8r/zUmVXreoVQ7HhXgaN2VU7v3aXDM95UPTj8gHIzoowSBxyEJ27wGzuSjr
cUAzxE3+2d1CXmcnbS7LL/HKOnm7BR23MpdsaTRq8oE+jegMRVds/YiCgqnVmwEQ
VJTdbAHA7Sy9QihxEmI82r2zJlBdnbrbSroprkzIes/crduqBStGxtgSOzKwDozD
lr/RStkbzNRS/I4S7oTujT5Lyrf0UOPcf4ulEG2lz5KQBqyrmNHku5j54nBuQ1El
9WBPp67onDkDyNH0TQyYYy5a/hs4401yve/aer2G1IK2xdlHsFQnITZpHBMd+p25
IPhSNObu++pC3de30PJAuDzB6EGziawZ5X3HRo1M6YtayoFc66ZAuHcpdwn2dUcC
zP4EGivllsuxDNqwhPBMAoxAA4EopN+y9OKXB8s6Sdkt7xuFb8iPWIDXgELrvE/q
HIkzJuCky2TJpgkVPzpUQKQw2ebgT1q8YWh/PkK/4LicaEZZSYv40jJb/rG9uIM0
6i79sG6LLdkbqWvPnuo8oHBpNPCdPW7DBPGG9zNeJ2kkFHOMgYtZID9rdg4F5Zht
s2tH+ES2216JOpFoCtyzwvHMVdBcUx1Br2wl0LMV0bPfYmsRpTVPQxDE1lX+ObKO
KiEgKE3u93xVS2NKVaDGkJIyBaO7ZFjHWaocYM5JV5YXpcUksXrn+ul8A37blPrP
aBhlqkOPI9RijapQjJcN0RVJbMoLYYoG/Cx6dv9yCW3N95/cbMZZm7lAUnlEk5ni
l971tp+LC09Jsr52Da+zl2/xNVHVuFhg0z/286ZFbYCvERj0LU8VctJADMeFFI8+
Bi2J7FZt+yRKVGz7EQV8geST5vP6XdARP063rjI1lzYFphcWWp+DCczWD9kyxauC
aKnvlHVSwd3DLf9raQgUILrl7CnGviRiXxn4FmDf5+kIrsUAnDKH5hHL8zqpM5Uy
xqZ6p7z6Dg3LRcg/VibK/rgf8dIFzTyaQdX4pyG1z6kL7o3eqPzMTjVC/3vI07R3
yC7WrgHMK0diMsBMa7KSTozZTPmGEOkP6aq2+8AD+nXl8sWPr1vo5iL5+Pdua33p
uoVGUeSSTtJDtAA6R/Gzq7hPnKKNV7JJSqkK5b0+nuRUr+wbBxN6u9evE5Vu2rwK
Sq1nk6MLXnuqQXakqCg/jWpaEcvarqBzh7Gxq1UTq1aeR/vtSE1kGxofIdEYcB9H
5GYIFFz2jR97DrOD/Xx0VI5nJRQiTsbw8vSV3ZYbaWyRRdmuDqh3LnbDZfHKeO56
KfS8m7pw/pzxlqzyAblDHzMDAyBadws5nCmtRYWbj8TX9uNIZCQXNmjLso/tZN7g
wl6UfEqv/RTbI7MjmfaRVd2OzNGABOw5S5kjS/+2hcVgHfyKAheMqGGVVGkUJpxW
VachNmQzKE1yGrKuj8LcjKM0RDsZzNmvahNcuBfhHEyGezskwrmqTDEaEFXjr64W
T6MriJh5f8zdJDtmYhM6RJsRffIqcb7tz7QlC6z7xHLyqDhR6KqpRLy/h9kH3+RM
WFV3MuzjbdODVzTVeDSs8gy96aj8JorrVqStZxN5ZiCZH4/3HgNAu7QKUzuCvrbX
i2BVutmbUwjMr7g72a8XkjkQzEH3fMzqsWasr9to9dceEfMpqFXXGbi7EIxx0MMr
aFmeX1t62Y6O4QnMj1xRT9XNlAy59HHKZGAFAW+UwCDXzcgH3d0FqL93VCaLv11U
q95XAvAyr+U59K2DGlhUES4AkQQFcffgrtZbaO0QhHwE9Co2O9KS9+0a5FTO8EUB
5SWap9BwtisD8RWfytgJ/u8cLLHbIE7s348CXyrBFELe/MjJPnC30ey+VN4PeXQP
MH/zR2fNhXiRBLWJrkSV7IfE3CRVX6ecyAJWarmPQdNAem/kSMNIfB/gqg8YZlUB
7iYah+7tPsQDx0E0hMnYyaxGqHbzguW+8eF/47udI8z/+qEJKUYnRedPdxuHPoD2
WFiJzcFmEILoOTAW3c8XxMUF+fSLaXtkhNy4VAphFUxu3PnixYP4R5ZIY7fiy8fh
U8KZBOvg6ywn3p7vO3fbY0rIU9VwnibXafils+UCdXNQhjiNp39LMMtcU/oAKyuP
LWLG7CRfGIuBYTJNBfmzDBb5Sp2AdwgHAjFLuQQzQXzLbXiBN2+yXHYltxFCX27x
86X81gS2VhEp4rahXAlnfYgyYNFWJv2hxRwj4pif+D9/wMaN7YwvGGrKi0yZ9UMB
O79NCJfn7S/YruovBPSK5gYrEO83Hjx5TYVSx9zWk/dJK7XwujMyEBaE67i2qjS0
CPHlr3jr5KPVoq+ZMEHMNpei03eiRonCtES3sKYRYRQXWqf4B0lxodOW2vi6hP5b
Q/Lqv+Nz2Rc8IoN7TFa4r1JfcSP1jswkccycpTEO5F9fK91PPB3TeTte08Rh5vcC
cRxDni2FRkJVBcCmkKs1V+EfL0jW2CLlmQh7M8odPL8Lx2QuLC3JO/MOX9wP4Vuo
pKL3gEh6yf9lA1wzRVbw6Gi3ZXatJuTfT829JXMqws2EfAoXMdXj2ARUiNQNNCL4
W+ZMUncTLfDRbex5qINt5VaADVc5hsv5kBt0Bq3NJJpc/uIJM/S0HcOIyAi3H+6h
T8dRMt2ip1NK/G2wCddRRedpDI0x0QE43EApmYuJmiGnp0sPRPPVMEwAMKCXIF5L
Qd+hrFqcEIrINqd+gTcjBn3gwQjgfr72TAR9DHa4LUzbxK9TK7Z/OxJndGEMYGjR
a4SX49MADDAg2X9JykaMCRwkFcNWQzkFkSJy9JcFOMTRHHmnHZzGrhe3Psob6oVX
9KGZHpxSrIEotCKxHXmXXW1OlYrMmcI3mawxiFaZdTtQJrBN7kxqiw/PZ7WHNMba
z5q9TbULqQhGZy+DRPx1Ne80xOrGfYY/nPnnkQBndnSceJPPBQjIGRbE7z4tNn1b
69+nKgsJvOQtZv1mWm7UBdTDaiL8A1ORKB5h1HyUVA+mH+V0FrDpwW4eFP0jeZV4
tLk/gvkxJ2DiXmNaEXZXRxaYwEf1ZePU6F/0yWfIomD6YAi/VtaaM0sfSe2+PVwn
HLEZivUils0yS8ON7XjrJH/n6J1ayTRMFcDZEHMk6by8RY4VJXsECzCryPbVDdna
KzdBVTKwXv5rduzySqIM650Bt+xoQ12JVKihdQbWhOjq22WufYZPeS5InmTnU2xa
Oqmjb/y6MCinAC1fB0O48m1+ToeUX7n0aw2ct0HiqMLfqd3uGcADuaTk/4CW4eXi
mFqj6GARU21V0Tgzt9/be5MbifDaGv64j7DUyggozVJVapMyAwePYCx3ChX/RqZX
Kon1uQ8kTJSIJKPovFHdXKh4RcY0c3qwo1FnaPoM9YH3E8P0geHQOD8jTtF92ymA
lRWyAs/bqDhcUqJ4CKEXGfzh7v/f3w0vJAMDT7t1tVd2mk0ZKkyZls4n05g+4PHg
i6+0rQ1AlnJONVKJMeoZOUg2xqzCQKgLsBRAax/w8mWrv8+YeLWe1mewYnHlf/6Q
rsBfwN6ME5Re9d/Js8eEyYho1EZHQluyCQxf5XvFuouWB+WUhCzyF/eKPVVbdWT3
sPbHqMkb7AgDoUAuYP/ap3KvDJ+lPBR+S7yBwHRsgdwJ4d+2txunpqhK0aApGFZS
FZv/2k82DjuJ3s5NuHGHXGrryjXT4woXD4gXTLWffOQDkj/F6KMSXrTJ0Vw8irqx
4YkhPRxBW/B4lj9QC/WHDjWAAI60b6V9wgMFI7DfwoWlFkHKEiYF9mPnY/mBpf+K
OrKj81OZDrlyh8KD0VA37BHlzWMWWZ71uj2amrYTrGhCwyciyXTXUnSbi0NgTPLk
QGPdJrZhRdE0i4FgSTq1wJWAxK9CFzogbj6nPfSpBlq3nynG39zRIGFrdqSFHjce
R3Ct3rSa/KCi+p4l9ru+QLg+YX/JSuOVkD0mJHxEBcJZTYmUddLb2doEn7VxFr3A
Kmxn0yBT/lOe+Jcs4RZrbPxj2npaBgDC8bdAXV5Yr9Lyra+TwskE7yvoChrxWL+M
w7uwflNT8/VyR4RvPEgF945r4sZ83IpADKvfgPvnowWcZ7qTro6BT87GTs9yz3ys
1gfnVtnY3G0LTZFSCzm39OtecN/FW9s4PV0B9rZGQEYi/Vi9T1SAinpLaV4hlZcX
QuAzlARcPxos8v0dWc84z6gUZ8pEk7kksyE9aFGawE0bzrHk2H0h6Vu2KRyxIkr1
Ab9JoMSPfR8+tRXOoNokqT/C0tpkKgo6PWb6WFUWKzmol3O0iJXLcKnNmUeqFy3A
5rywbyp4+/MUmy2ZWLqOFqswX32btdD0mgpH7G/pcGzJL40klHUMQGpph73xmz5N
Yr8+pO9ASBVogj25ST6u6m517oGdx0fbyp4sCQLp+uK/B4pyOIlp7ec58fBkstst
40TE2unTXN0HVPScLt4Bp//mLoGIRwyu9ZIzTCEmvv5d38jiK5LCJJ2N85vOO+nJ
AfA1XkkhzqWVzwlBmDg20Azwfxxc4Ivz6Edp5GHzqtKs1mAYeBQ0il0aMzCXF/0Q
pxepJsUe14qzLkDsitXLQT7FFqX++WETxNs0yOj4uMqejiPQtCYFpqrJB6HnfAOJ
kbFnEuG8nTR9dCKQODzkh0cgZG0H5JgbbJFNjdty3gq5yeB3AFueJ9xwHYC641c7
dEvQCUwNRGDlg9weVnznjCL+D34l+r+PpXTHv2xSY5tnMLdVECWiZZqG4EKpSEgk
A6N9J80bFL0ayCZsXQxcqtG/SyVLjLJtI00VmKTMwYpc1GYugG1BAlITyLdbk2kh
3XpkgK8nl50v0UStZ7hmiXiuf5lh6iN4TpS+zQ3JAV5m0Qoa6siy+wDXO4FPCH66
f+PlYfZ1bwoCS2b0QKCT32NBKFZn7SFB6aAlKxDbmGeYlC36mo0oG+ufw/cSafbF
TuxF+gSX2ziD+fGIEul4fUsH8JEJX2MTFLZkvqdlRSHsDY/OB0cOZT6qeg7QdN/+
bVBrX2l34/8mIJRXFrWh2mfJxHLbAXCZDWczMrhbSKkabWinlXZpVW6PVkuiCnmi
FTBvIYeXemvyc4cOLLmCUzrtFmAsqfXYmW1swIYBj7aji+TrJOGqGrAEupPO6vOn
VHDhftPIwuER7AeDpY0hwNYADZmutiUGdHcve+gmrZC/AXq4CWgxjOYvTAc84pHW
wLb/6kG60oSYYfQqcJ1MF5o56uMyoZ7gM/oPm/ViWdmxTfSCu1OcIc0HsurCdpKv
3OuxkOR1QqEF/HtMEgLO6dDrslY60kqlUMSY10yUdrwpGKoZqMkqhnK7jWHG3xqb
F+Q3RpLh7zN34X3zJzt2veegAiWWEsyEFmfV2Wn95kKAeeow1SvT+pTzPdypdL7t
757SQhdXLHnacIqx+BIJpiv3ZtVR8NLOaWaem0edq6MP482a4iBmgOzrJDkjSSuL
eWwjm48A2KSPzoXViE41g+JJERqJMCv1BaHcazS7PBxI6vaC5PI40E7avTxsAtQj
sdMyn9Le4x+N4QjSlxFsX/F0eHBihISFe0O9I3xkABDXPwo8e+VF7FjHFILgUmhP
ez2dr4kzx0PkFSG63Zo3RvVu9+omI8f7gng/DP53n1ukAwEofVmZKYwI+FFpXQ4s
mDzit+AlOlZCk7h3VenKwuHy+HCdAokG1dP9/2Cv/9iuDkNtgA2hvC6ZSeQ0EbNR
Hqa9OdQPyaDoQVstDAAOrBMteiB9eD7LoKknupmzFiedTBMRGs+1vEnVPvGCh8dv
a16EGveVIaa2js5hFP7FnP+eRDLdV0ZLpZIc1lLFeLixtxgyXqrT0i9hTizMO1Kq
AmLmFLUoJbzEeo8p3WxbWWy8YkBbFMCYNPYF5qnbgRIFKNXJ3TDIrrMa3nU3zOdY
iwegs3bu2YbfI7NhmNYAtpVSYTGVTcQGdMt8pVSOO5s/QIMPq9NuCdYEeROKGO4n
ameEcI978n7ro5A/gRcfNkrWj3D3/FqJcLoXisHxV3rArJfrS/i2Nvr+2XFZuezP
EuhVOabxpAk3mHBGOHhXqCL60lbaejDT5eJPjq7ZI7eE2aoqA/LeIB0leeoAJmb3
t0l0mfYWYkEMJu1Ezx+VF62Um7ibRs+JyyUcNwQTOzSSBdr7oV+XABpvdnkkQgzY
E+RP/0bKomU+CqjpyCP24Qa6Aha7z21E1JIJz5OU3+pgh/8dTt4nDsxI92OVZUVk
9tIZjkfCYFIkAir/dXG7eAsA8rPIV6HnO5lfGDBtvdVSnGKnKdcO6kqi4CRIMHuh
eWAKw5gqhkzvoLRt8LBC6x3Rghrg+kS3HdJN20N4SkN9Ki8hylTyvJLbHzBno+8B
gFh6WRIXLGMS/3TpmfEQRjBB6tn/yAXyK1T1IddjxeyTm4rnEGAYwBfEt5rjnV/R
jM2T+7chM3WTg70UXmELcLZw5D5yfS+7uGD0Y11MO+S5+d5S3TWSakWPJ7P/PBRx
R6RoNJiGnvPX/LVlZQaONN2jogUs3ujr5E3h/LKdRAkGwQ2moFYdlCyqyjHnrmlx
jxDyQF73BzWozyl7mU7+r4G1NGJgRgGJKld++mlEwVdSBmGfTkFuwlmog5qG69BU
p4qHbHvf70pt5KZE7u2Gt/L0de7sMUUz3UQV3USzYAqjfvpVXJumlhM4gYsVuqO9
VVa4WwxRb32pVfJDxuTL0S5HhnLk9x+lgMfnPrTIoQuHu0MOU/dCbBLMdIzDXldv
9Lk/ftTPiJY9cGbmjcQFtaFQlCe6T2+fNaGJqysMT9hXowwfKVviO6/+mjgbwkIQ
cp7U8bEbKil8MnaeVNYKqecUSw90deM32GnN4WEXyGgQCcfeRlf/2xm5yH8e9YNT
efgwhWxMM/Tg9trl1SjmJkat2BOztbCac0lQEzV8oJlCCIfNYreKa6DMsQGbRWMf
mDzhvBTRiGF/d/cFduXsQfiK2bfXpPg0erqzQDU/xgY0L7CkcrOnX0jwaaaHpkKb
TcU/BZRfGZnJ7FmJyN09tgnOX92DL6A9pD/wZA42e8JkIu5R+cLRcX4CdJw0EZK0
vTJIClOck5zUtN0CYw9UuHaGXegwfPO9Kx4yGxmADCXrLlocZuHkKifwsQdXJWxq
pk6beFLEFC/QuRU2/tFQHeZF9XPBiGEUcDi0jzWppxMXAndFAfiOb0A+UUSBVhhE
G3MsEYQSst43MsE901TpMWDFopmwlB4INesJzYXuJZmqbi4G6cgVTSWy7TuxQL0J
UjtY41jgFFDHwEcNTD2RSisbpvYUMY+5sRIvfnw1IgK7u2/BcHgSQqWi7nWZFzbP
G75A8/Wm1rhApVZ6TcudLvavAWjaqC6BtEC9IeqtCuJZoDGtDuKp+SZFOOck0VwF
KnR42aJ1eEadpe3Jo5ANVDmIO59R2HcUPM2s+LGSOWtq7D8P1qACAF5RErj0NFuh
JEQFoqBxJRMYFdJ9YXE4WY3G4NcKKsZFg0ssIvmmiTvVj02U35L7R3y8W2B9XwMF
8g9+PzdDpuRcMb8VGrvBn2jiz/cnJXg3q/EmWMfiBw5uXU2Jrz1vIEWgn/WcNUPV
zoyUCpfhMxCrgwroTXUWlgMEfzkHNA6v0QJh5eY0j+qCabxVxwvonAK/f+gvyY3E
S19NsdktJD2az1v8nDEIKrr0KsofbmI7kFyhTXSAZMiL+2ZNVSkPN5Zfooopu18P
tinqS/3oiF7C16z6Vf31Y9PSBwp/mVdcb+ZqZIGLuMoaI7dcb4KRCptxcGyiGitn
/I8h8WQetblWtNNbxH98+M0k0/3o1sqdtTiiyhIuhDXzwsfuxcayMEAxQxhYJpbi
3WBWPkLmIMpABBMUQ5gEaQOKsXDwqstVUddTWVBx/iq/g+LMZtYYYPbCGRJMpeIn
FJUhRyIKVZuUa7Cz0RkIfFLcfx5XXY9DiyZJQJ1JpvuYME2QnWbT+b3EDZQ2JCu7
RVS78alkhoGgZx0W+45Et3K/waLNT7MydmM4B9hJJzsjUzt7tlCe0+2tPZT0e639
kVc31/9M5eC2KxyVy4HuriCuIEoYpbRLMNpbBRBeJzxBLwcLlbj/QktQl7s1KhP0
l/9bHF1pLVp+HcU1lWCdcSo6H18NmHa9v/SU49OzMnXFeiKeDz/xTNO/6e9bT+k0
VkNrlL4KACjVWyvylJSn+mo3yXLPydepaQssYrOkPFm7HdUOt2ZdgvwxESUeB7lD
+vMnM1DJzP5PDKbImYlMhCKM9AJectz3VagxuOY0EXHB0Q4C+b2IYnicaBwTpiWW
hKHrZXEHiAT8T0pqw/nySN/Y5uPgSPXueRDpotHrsz8Mf5e8d3UcB/3NVoT5TkMI
BaDiWDogNxNO85VGAIst0d/EV3PhAQl5l+70CIXErix56izUic9fnnUWUpnKNEGu
HfQn3iM/xUrAyEBYwx1zQVTn3WKGg4kYoDsCxyE8+S+sM6n0Jnaivydt06bhoPlf
Fl2ASf8RzvZ1Ynh/S9CVCdu4pw63Z+7Le9LxzmkTwPR+y/2dcfLilIuWO2JtOQ12
vl79pYGMKpvfqA/zI/L3IadsLtYD4JUjIMn/CzxfRd8qnYR910+Tcq+pwzT52Rwt
T6487OckqQexuV+P3TLMu0hnDN/5371TT7cT2wQIS5aPRyzRDX7hr94nXjf1tuwL
eQ1FJSSsx65EdfGDu5gj3OMf8A+3GNmF+8sJR/35Ntc0nR7Phwy/av2iWMK8XFA1
Edjzc0vGgeW9fowYzxzFOWSMnUX0qQX2TiH3ny1RKhjarE+ZLoN3JFAZwS01+9p4
B7DseGj1d2gzQkaycy50CxKWDIUyIAv5c2NbeEEwtYtppIriosGqtbwv7HcVqaUC
RbZUF/oHd8Mc1VOVBUdGquEBFrBAdxZACkbRYO3PYwgn3vPNELnqxsnwGplyjsSz
E1dDVJODTl0MHVs/XWXSB1iftPjHIE3BgZsUxo44rVYVn2sBy78Pn5dvMCbNQrJ5
h7klgy2dmghWpQi282JcpLpphJvj1gYJWrp01VwRpxQ/90BSNV9UfdwYHfEqJjFw
6xtFg7wE9wqwVTxlkRqOd85CV9816HXUiWIK4kpBua+s9S7xuSG/r7ZtsRmv6Qvb
VlfBa/PE/ok2EYFsCowutKbpWA0mfZXcJ/TdGak1XwrFo4NL3il/tl7WybczfDR6
/RTcEvmanWrKRxHRwvAOhrTM87W7Mo0g2Aa+NJXN3ySAL5WMYW5dxsvWkLFsYnkE
NQ2GjQSMt/ELdcG+Bq9Lqqtj71UoepWcXC4kg9SkhBT3XdNZlv4hn82pv0aiOl5c
sBkruAuKa69aidEmKdKJ1k6uxqTpzmfYiBi3yR8AdKXrH5jUQ5c3S8053iZ22cqp
KzSpREtNjTRaV9UAtTEnCYYcWx2eqbuZCQjFepXwENgzMaFO1AjraG5I3v5WNit0
Zc14NY1L/yon5DVXBx0RiTe5GBz80wXtjCHpyDsNJ/5wamzVTSH2xMOZsuiPv2ag
ciojZOpOLggiwwiNDj3599q5hK4k+K38whf7KRwG0amFsaF2NmbGSHOgR99OESzq
tV5mPKd1A/8o+UtmU14sXwWlLoHi9kRvslxgL+uPh+zr3sphGSOLdE/zJJXv0evI
VjWzAx/i55FGiyyBTqZ+9F9/UaU+WDfyrK/ZDNlAJz0qogF6BJd7zdETaB30YtBV
EgGByc8DJNW8+pNcaPEBKGdd26ETI2pgm+F8cyNOoBV/KsuzwNtXR0jXUmhccVKC
n03EiAEaCuOU4ciJdC6XxKyyaJnAtVS5YGBvpKmDWB4SsiBgWsGQ2tN77ncaAv+6
RdfAV7+EqK+BLCMh4EGZzVGWw2FxDXSh9x0NQFYUCoObToxEFfrxc4V6WOEYKNVm
E5xwhQizL8OBS8iqkHUbAO/1ymRb7N38yhWEqf/8VC0Yrxph7CUqpXNZQ6Yd6y+s
ZGMp+q2QpsOKeuiuIqFLsWig8HUhx8cJh0vNwqhnYN6ygBzMiNOqGbwP+nDUy6ws
KIGDXawhReuIkPPIRlz6cRCvzhkIYYneB+z3HT0AVAHeeb4SxLIo+3K/xfe3ej4S
0aspmi6P2lhjk7bpTrn/WahXJIjOL9LBuboTQp7oZbGtLrwAbV8rxm/vD33XYoPY
zGYfHJxijm1d+X2ynUlZ3g8Z8b2FUInMjIpHDvENe8XvJajliao9ZeK9XhYA3QTN
sSANe2fQhlB1ch3cgdLdfJ3v3Ox8og4jVlaH5Kcu8GzdPgzqmX4/0mpTqE/Fuy2W
Qy6D9F1CuT8ZVbIErwh4Bu6gGFzMz/gYLqmOwVXdmvxJbRmtoGVV+HHGJNStTN0Y
2UN+ISK6tT4ZGqQTYvFTcjU9qpaDaaf7ujUGIj54nLYdc2cQKV8qPHB9WNbJmo0f
B5g/ZY482ceuUAKLMxXQxDT0Z4SfO9Po824AHNMOoSrlU1g2hNIvXpuBry7PgBKL
pwKryuUHOBlW47Pvta60x+KTx10LarHL6tLTIb2Uk82k6qTgmu7Wxc9kevDrWyF0
aa4X7kupr+Xm3FDs3Vm5p1okptT0uvyV5DJl0bao71JBefGAwQHM17oLY2SoruBa
2yuQFQvon/Uw9176OvBEyVLkpWzQpjVD6AcJUxf637mnFxhAiP3Fe3nra7QYM8eD
DPU15OTtctnfZUJo7wcuxinAOWMcj5aPLTHclwmLpF7FAhLVf9jZo9t822mLaaU4
bp2YXe06/66+l+WvZQ8Nsq+AYkqIM2hmPVj+l85puiNxf8kaC8GIK0k9O4wsMJ7T
d+F6IEgL6Ge/C7O2QdyOQscN/zfs4lz58vlYMAVTREj7FWXbODW4qz6kPzsfuWIZ
gk02U6HSiRTD46/UEkBl7Kll8tUgNyi/zH2llPvJGTISu9hON5GHGkT0l1VvcPgS
pm9neEThvrZarNzg1gdU5BB2gt6Ks/bMh809FICvkGjoikVOwhot7q/gWlopjydu
mWTgfnyr2Si14+l682eSa6ROZbmkUEcwO3hSyMXhU6z8gHZjFwUebSTi9Nwt70zG
36d+bYxLHS05JD2YnrZARKeHp6zKkQSMjQ6Fsn2QNgA1n3o6Kn+6KFGCrpk+XVTU
SRc9I5+NzaoE2miHYM/lIZORq7KUlKnX9FFu74UVpxaxDqY9SU++JRq3m6oGNHmz
FJntLq2d4ExhFdVUIyYppaR1EQfRdg2xEKswRdz1ZpcwDzBkecle41npOmtNIzl7
d7AXbCI2Ke3ngHlYPTBWDsRZeuGdbQHaYVwc/vmdD9EOq63lmYXPMef+YkGO3wjC
8nNdoNjYu76qS+QlOZXBiQLNVQSLQO5buVtKDcorU8fc7I9YTBZJ1hLcf1EmKdDX
1DANFQdJQbd+M0t4iipxnhecA7xUiAI5MrCGVTjXlj6SOt6jW2h1nOEnbzLvrGmU
rs3KBxp/EgmwOZc8mpNH3g7THxgrvEpQIcva8aEiiLj630ShLkStYm0io5cl46RI
7nu4IN8STTLVAML0BFDqUYwfIRPBCKnFqL8WQcxcoQgDig6qMW45CxvS1V0OrlC0
aNYeVlvHBu8l3Omvsz054qp/UqafvxDE3ZBnZ0cvJUyXKUQBydX+z/AQICh++ST7
DajFNS95JftalUFqEuVXPirz4fDwB1Sz+JFXs2MiAIKGj4bH81YsNt3dHsxD9R5K
Y546V7TsILaVVRvrFlzTsUQEaia/HlwXJboev5BdBJB5uqaC8rGYhSlNbF7SZhmI
Wos7qdb4VQ6x8N+M2qjIWRMVnLPaIkvwagKPyiw9NiMvLWXptbv3UlcekyhzOu+f
6Eg7/KozntrZD+rIVJivJAacJNqVupCo4Fu9ttdgSs484Rf37E93+heaijwuWubS
e08ZstpYH0MLtatHguhhnSWJ0NwiEaiRQM+MfH9kAla0El3c2g9zYeKhF5evNGyd
TEXfm3W+DDEpXd5NbZ7H+at87dQd+TxSXX5GZDA5pqhq+edYcYPL9dEKoZsYW/RY
DMb05gewxRtB0kYA0cbZbg1FQmYZEDuVsIMaQqJB/M42revaRVjCx9ahksBFkmwI
IKDh9900vAmbQgmLB+NkI3Ud3V5/mQba5yH/43nBZNTPNJe9SXKHk1Woh5/9kChE
lUlOhJy0y9Yup1EtN8RPerL5DoHAV9fCyIwi+ElOXeQ+Ob5O84t3yn31IsY1LJYr
oJjB8fzbawA1hUJ+1GZTUo5px2kzxpnq9CPgl682gPuVBGrOf+r/8diZByzDnw1X
QAm/vscSMy1vABMLsUVR4vtf2ICasA9zMDcqThU3lB3KddO+ByRYLJcmgBH0KaIU
hO6/aV+LUm7uREhZwnup2L7A3VwmBMeuha5gwu89P2V2f54Ir/byw2jbS9kbkjpF
EURXpw/iKD8ynk2xl6WWwg/2LvJzJsBCVT0QUL6O0Vvk0DyiX+sw4q0ws3Krow6g
hz8tD2U2Jzqs62PCmRkR6yNAqKWn7APMNYnKenNUPMpH+OAdoFH2TPnr0514dCQy
xpxbFVLMjIKbHoiCeA67b1hzy/E+fvbxxK1tk/qBl862FMEk+X2MC9sqWxAv/Rew
tnNMT6Ao1vAVUhxNTWvXuyUAO4PID2c2JzWhkws010l2QwfNGRC2DdYpmAzcs8NI
xL6MN2DIdlMEQwmlCNtuJDej1qjSbK6KwvHO+NPq0QQWDQv5Ex5cz77ImfhhckeY
yNxukwbKvHmAuCAzooDqRbNU7r3pw5axqbCc5qbc+z61Z3jGUybrRelLnSgkKd1K
O1G0LTKBgpKAfAJgvUK38im2qWXQCdhPNeB4J0BUn0KCU2vGaBdJYsdl/PYo8bLn
CsqicOFGch/0Q4Xn2xxS5STQBiEANl4DJftT9M8oijjLOu6q1wX0Jpq5kX9mxczH
5HsJb7ivPc9u+tXrItaW+DO6A893i+dn9dNw4+0fHyHuzMV5HRGpJapxNLrXWZwt
eWUhVsZBO4f/6QxYRpM6EWxgNBliiXdp0n8D3T8CePpMwPIJU4pf7uI8v1wkTXbm
ORWW22AZEiR3yb9PxtSES5TaYP5j/PP4TGZh55vl4Fd4eQTli2RK1jfYz02I+8NN
qBse/oc8usrSE3VSkDgxN1B0JnVq1chZy8W/DO2Y0FWDJNi9UBepP5wXPcmiJjmI
RrFXiYL+7ZRXBwFmY9CP46WSO7TL0TwjGRpb2zJW2z1UefZZ/UkPRdA+M7sgqFhj
IY9/FGYbUxVIhZe1yDv3nPH4FvjEppxYDNYBMCmUzVdwk+GeKvVwZ6cVlRNC5DNx
t1a8m/vFiSM08ELOdQ/h/a5nVTJ6+sz5q2cvnN4I0g/EX7fNN5yFAXsSI7WvjuFM
jwltJGCXHjY2LPRBazggOvtW0akXXXSnfHmyTC19Ee1xZAxtk4571nRYC3n23GU4
McXREvCvL55RUs10UP3c7WIV19aNLFjBBVlXCoO3rXEE+J4/D/Ptzwfz8TePSdCB
zJ2SHtM8au9H5nVhVdjG1l3bqotyIbIiCWNiYf5hWHIEoogi51OlWT1U01yc/n29
bcuL92+5KwstdfkX7ngTPvwFfck2JtBZt31gevpan6wMXYYyTPaXcKovg6HnYX94
ihAt9rFJmUsVOefntv3m96CbwNH2M1lQbh/KRtdGo6JWd+Mgq4YHRyot1GwWphhp
nFaXqzb1NERd777JlPRf7F2Ij5Prn+7Z1NTXYKlAo+/qrIRXBV3FHbonn1uC33tz
qvlv+6QiuqG+nXS3gpIc+WTd5dz3Vbjpy1ZYnz97ZzNzgJYW0bP/RxjEuaiGHK82
BOc5dpiCN8DtcEW3OZgPKVvZcoolz4fqBnZ8w09fqjkWkigsAWsnzfdQ1Z5Gx3of
et759VQCKTTU64AB11x+scpWl7SDGWF7LcH+QfbspjUPEwRLT0/g+Q68FXuQIGhq
RmLowkaZnVV1wHSwkIrAdx9O0ObcFss/lvvV/C/z6Y9Z87yBQGq75frWwMPfp5F3
R1Tc9GPsFbROPMtVD97kj0lOvacs1TWCsRqiE89J5hQOmQgJmLDmM3acN8P3wNUK
a2QchestVKDJNZuy/mkPwcbOpEp7FwlbjaBPPlfhjrTr9MqK9WarP/K2mJiwQW7Y
sYxU8Q1q+p5TRHpnCem1g6fS+vJQbtWI388MJOoXIRXscPvlwEbvylRsG26+Mhzd
4nsijflsxaqnwDTvnbIgpPuLAEkCC1V+B3err1yRkvajAtnk5+Y4+66rM8JDROGQ
trOR+ZfALKPbWoHjm5/ZMQ0m2NBygVMmjHVv6VKykOz9DYWf1el9mFvh8MCPH9TU
LWKFMWfjbVe8/puw0k2i7OEd0Agxkk1RWKB5of3Cc1H4IZBgKaeHL/jtXOPcriHR
InR2hBdj1H2CuCmqn+dgBhyL9PDD9rZmPH/7H2XjGawA8PyM+E8X2zCTZLEjH1+D
hw1vpZqE/7msfN4HAw39YhOff619RwSeOT7vSFu3Y7pjyDYXng2BlYM67UNj9mhx
6IpYVmNj+axuQ31ldHcYHoSDLe/QS82djk0xhtPl7OVD2ZYiy4VARFX9hoOeqYug
PHl7RArLKYI3S61afryXJXc1pkMFkgWUw1ue5ibCzJwtQ9y9LjnbZUiPU5Y+thsZ
10eQlZ9GoFXfQpjlpisYNAuNQ5UpcXtp5ubmeCorvgMpgBV/6J66HAIPbL/Nrra1
JSRZlZBCbkz+tMIaKBV9mSBuSyq/nSlNTmUy8b1P2s8zFIcj7GYkeh5mMfaE5iJN
pHh05GBQjkbtF6CR9yBsUgs09R+AtX91gOHGBfI0HfDMkU12XLeax/BA5plsdp97
PnSSZVr5jH4y1o5gYaPWbPuIaKOPyFSnDC0cQ9c9QYaOFOpgm/dlJB98Us6E7BIU
yEVeIoLAxGMYxRj2th5aHQ8RQRlE+KAEPGuip+zglV966g5Nv8x0jytY+OUmC9XK
hguIKU96b0kBl672QncltdEvvs+PXEW+liZTPY+Kinlpzx3+ivjJsVzXzGSVeamz
JTqcs0qPWRPJCD0slZe83vmnMApXQaPPw60PrY4019rri/TGnYRKURUF14LhqQiT
LghYPzE7ZAe0OkOhSWsFnQVCanUjL8dFXjyWTpckGAmpCJkWS6HdfOLoSYBYGoyF
kTOR8s/i9bvbGJmlNDVrem/QG0DmGELxWhVdtdAAsypFh6K43M+IK8ZPo5WKYEp+
7O7nvmc+nBCnWRuZnQoqyCPM2VVVLpqex4t9uGZPsVyfEx0HloNSPtbOAEjMUJIP
CzpkErE7SV3x0g5NmW0Fm1eeROfoAsL33c2ov0vkmdO7YrAfrZjpBifC7Gtir246
Rej33Ttx23ZKlQAGfbZ9i0tsn+selGYJSuAcH538kxBYhedIfsOpGUoDbrFbNehu
kKIyprFQKcSQjSiFMPSGJJSabhxFpLJ9nRYgq8nIlRR7ufgOv3hC/wV4lmGM7fSO
psZb99iM/wz92Rzj1jjvv3pgEp/2V2aZc/ZoYlcIOT5rQ6+NNvtCAY5U5n/FaqpK
kn7P36YhlUpcdlrbCDHjhS7/YZ0H5vdhHxb6svOvJK1n1+eTOuStQuoS2Z1St7E3
iAUoJfROAVyC9h46OK8+rH9z189Zu7az4uX4BrS0c6wc/xJPLasOG00vBGFfMapl
vQ739DK6ayzHnJMQBdsbp9ewA+RSsk6Ve+GVqgKD3E/CWg7tC1WvhMopAZmrC1i4
CD0iOcgjoRX2DyQYrdvyJduAIFttN6YV/5QqxSYAB0HGyOGGTBo4XtWRUqOJ19Kn
OuSyYPLT5DROGzl8wnoUBry8shO5RFdYxLLDKREbRbDE6j79NvC8UxFHFb+1KuST
yOsbOly5s/yEVlazm3GHFD6Xpp37JSXw0b08ntc14jNNzqo1KhTVRlprYlnEGNjJ
8dm/dEEut9hBgPxVDCYSZ1Pq97iQWbBVSnVN+Z55U7n58eKVTchIlSG/UAbJMN6J
utMrWGBj8DABCVq4evqrKrw4/Vex1sVmKJDqhcYwMowU0mzP8jm+BT27KyLTn84I
Y4dlNvw60ruYGlAgc8JVveYdTOSxFWo0QVo3wqLXrRNRMezqJHPIB6EldR0hzBNA
7La9JMosgAjJEAngJX6DCpBFWhqJ5EfQGURFd4lW3VXi209r15LnRTYjChQbvLk7
FFcRCvUSAYcMoI821Uc7TIIotOTITV0+odvOuItiy1axv5qr7abKx0k6Th7b3DFc
lU74dzXmjhthNdBIIQ6f61RfxePZQK8gk6QKtI+MNtmigGR7fDqIdogr2umOj1jm
RX9tU+TUazpKj95319oWtMjcjriy1icLLi/vz5ZA8tb+DDiV1frW4+xCtpn76VDF
EJUGSqtf04/turtv0Lom/li8D9HOHnarTovdzmbhib712rkOX7fHWfTMd7qQJelv
zY+l83CeaGNvbv/Az1GIqeZ7VDTv43hwZWussHvPWUHvplhxrCPS9/Ykc86XYVOk
XCTJM33LvmAbIerYY78/30wL3bHboTbSKBGLdItZvW1mQJUNvTQU+kXT75sonRty
cQv0ExRq+cAAZ4ufROh/jNHdF7x2S/5njQZQoTyUcZ0WWNM3SeLgzMTf7Kut9eKS
StMNMy0uNQ7yAebMZCxUvd7ywuCB88e20M1OcR9pqR0j/fa+FCh2ZEu67diYIz6Z
Ob7J3C0RJ7D6k+RxYJVaXK6yiOJIlMLfoAOW47oJPFsrK2uHA38TeSCIO83PHj6X
HJN73SrXnVi1VVtOOKt6XViySqZjlUhbOopNcFFCyONePCydEBK27WpP08ij+pY6
wRLo5doXASqMRDb0NjXLfXLaJLrYy2vyea8Gt5G5IpoM3s/szpyOLC70AcY46iP1
k1UI4sBS8UNOd4NBZR6LOBAnQT4EKqZaY/aoYFMtui0iTT4HRTKoqr61TF1dsWwb
2t1y6otunVnkE0QYcsHNISEvUMJznvavg8vCde6KIE7pMWAGFmSDsL6zl07Xx1iU
990xINKTbUKkWJYHNAmkMa/JiSi1dH++TTtcQN5XLbbT2xNlNiV2mGKr1MIXS1RR
SspS+GGLtX4d+nPnhfpbHSE5jfw67AfxNansSmYi6eqNNc/XosMuzN5jBDceNPNg
7JbXQECRlqhguL3dblb4/aaRYRdnTBEVIXKNq+7dOiAwFWx7z5/sBPRQWr4vtRDz
aQlriShUFd3vRr7cLVOhUnIHOxuvPz+Kbb1r+qAWMAjZ4mL5xKvrreGlfBPfRxS1
Ga0ITo2l0JT/EX8WFc48MiGwj3cl0XvVN1xclloKiaYNM1j6/gp04mWTIgRwgnIb
1Ji//l+oQsHdU+NUTdhNLtXauIJJqsIPMXXA660JXDNeoP0qad352y9vm7aoliwF
j32U6eZLYJuKIpReHmWHOzGsbe3Y6Qu5lEp9RTX7/EOjANI8QlN1DVNO8vkSmeWX
n9jYKdLQRWT9zHbrYfFDCgUewpsbSsiV5ExAfbZy0Gro2LTkqxbEEK6oYckp8h4S
mJxLDDghX0WZnlM/pbSuZB+aV6N+UXDg/2AEIt8rA2FY+6fjYuMKz5z8CrxTaFbt
ja34P34AAwAW6MKh5MMJOUJM/KKkBE+ByM90a3lfXMmyDcbNnZAYXKi9EdKXfdTx
kwQGowwvxUjc5Hf/O9knh6s4iMZoW0zYWASD8q99EsGlENy/KsNhY4Z8ud+IENHe
YWGOg5II2koG9n4XJmHKFn62QYv6hqJ+wgTJr3gpIQIEpG92sVhrKpjA5vQw8Vue
zGXHk+qH6Rp4auaIWC1wxUY5UDecPXhvvotvz2Zm2trT61fUQZthCdqcPnNhRJdV
I3DK2imMHPMUORa6ed1roHPe7h/M+1daXn2Ds6RDjb8H/s+LnlfODiwrOZ8dvblS
rVFG8QO0d8byou2KZOLPTdcLroZUGfsrHcBNB5pbqgJpfMKXv8XpFG62XJMfa7XS
rsIKwRQeXGcy8lsJxsNSouryFUl71VABAx9nV6+Vr4VcZnnIsO7374iMQa8pJtHQ
FnfE3VR712NpXlsif91jf8lJnAYL8b9079DDRqigstalGowyKlgUCGdGM8hhlBFb
DW02s6IHYMgPeAZ5bRzBZGwrnh2GsXEmWwGwvzsVgF4FTLPevL6aKlmYgT95Bq/X
7vDl4YLL82hZTPt50FfhxzYdcxozybD2SSAFUR+VNAK1dtnK39WicaMhSSFHvc7p
yZKCnmOd1S2ujUzg9xTAeDr1gyBon+zndc6xTycPIBY562pVQ9sZcFWWiDZEWMQX
NiwClDabL0Xzs45AYxLQM2spHQWQhdzjizNiGTgm8aJrArltmYjL22i0NJhKdRoN
zEnbv3iDuhH4S2PRotkzbGa6py/K6QEVILcUHMSZwohHQ41cHvKjBJjO321rX1qe
8l+P4Fevp7WVv8VEU9VmF7SH9Wp+IKUmKPr6rcBocIX0aeKIrxBsor54R2kpisWs
JqRnAPHGQKud9fJOKpxvG7EP9aUnTxPJqESiY21sdD2v0yWJAn95QL8GGUdlKcUU
j9OSMpI/QltT3HRU7WzbHpEobJZEYOaBuaZbbGBelWfyCOMAwVnRTjDTDSjh/RR2
vfYBO14/G37+QG0/eHRrA1GFrIcc/N6BXiyfPNekLq8QL9VdcXjkDYnF+0m/20oa
AyEbl9XzS1qDlaXVV2Je9snSSX3TyyLxmq+VRrenDoDwH275u9iKfUUzKUNzZaOA
Kac1httwe0t9t/Pl1B4V7IpeeqiS6RxnHA6R9MyUL/ujrAKElm4PU1F3BbbZZEa2
p8mhMdY7L1jd8v/DJfp9lgzaK0UktipZJVZNtne5iveWRMDF4XTa1zNiM9GbHIdc
fzchG0N8/ZJCiKoWQGm1gt9CPtNEfk69YEa7XvpcqmCWHcVgOsB//C+PXlOtXShT
MZDGu3fjtwV8y4mTvG0zEOvhD0e+SPfezI80fd5OF1I9FHQlSVB3sGaidpkC6zxw
/NwhqpPDPuwD9NQ7+W4ZqJWXlxFa4VwcHcTd+1ooHkGXlxLeaw+lNWKQhO6Gy4tJ
rwJqngGAUBBWG4nALS/Wbk++Ry9L/zllSHArEn1B8M2i7/3blBUEhrLHhBO1m9Q1
7lf7XDUuztbrcOc/jcPRVTJdSVaDFLuCw+waVBBdbendYPUVm/dzpnHiIsk9x9KH
FZHU7zZW0DErcegdp8d0Ig+eVme6rDR1v5YHROvEZ/RnuggMHeQh83ppb9FRAcIO
3m99O1qzTVyGb3/hsQ7BnYOSM4Jn9uVe4MZESoaghq/O4Ep41CneVbJfQ0iyH6AT
ZXbU5XbXYV5eBYWVYfA+fGnSP1f9W4/yF3qE16fB/S/XgiVNEk6fMY2z+RagUlFr
aBqe6H7synwTnUl2hTxSgs5eArQl4lJjt4/R6DxdyrdfT7nw7CUOHd8gMFqPamEY
JSVmVzRVaHhyJkywCGGGydtAcR89/L7a+4dpS8riEu228PDCOioCvej/suOfkT/G
kIMHm31F6DLmh7NRyXBfEaurA2VgZNKyx0Bz33IGUtoulDb0s6u9xqWzzsA2pZ7Z
UOuTzcHYujbpDOPKUGXzK6X91f3/ZAOIqlw84+zBcYPgwyjn+LbdajOimvogZ2xK
V/VQk8Xew+Qgt8KeFNQAFsIri5R/656vReBpe77/qUFgeXS3pgUsRpDcDHrCpEpB
cFkV+D6L8FaHJ30A2UtTSLwolDbGyyQI6ioENKdTcS9s9A3msUkPJbCUECVL1PES
IBuGhgQ++D2xk62+tOV1osasZJ8csXFy2KHfIl0K6UXSOpw/pC6ygZEfMTsW+0QB
PORBD0Xy7ftjausDHCcmyDLxEUpjxUryMwVojADdyc4QAe6MRVlzuSvdnwCot7j6
N0hPGskoJzsmqY4qBrso9/2i11g7cSuMoyOy/4U62qjjEZ/jTnlLgiPjHJvolNdz
XdeEG5KB4Zy/EbDMVlszGpNL07PxXmbNgDbf1ttwaa9kYJ48FFEwP7lbTsEIntcz
Kn4BanzyFdXVgLJvyzBn89PRUGWDgrEXOXetYfN4+Uj43w0eYpcwA38QVY0Gxv6J
pz39bm1LHe1G64pXq4ajgjO1ngZuboieVc4w+bKRuS/FihbhNQ2+ARuo3F0QaLDK
I1iX6N4TuCiGXZFnpDpQDM3ZNCAKp3rY8NSr6173iMrLBSwmQ9V85gicLwwv5kHt
zWbXGfbkJpwRzka7+MHElq78OicXXhtcCM4ojl5n5UidukCXwntb5UxjIEd1Q/6Q
NUu1TDZIqQFct/yEVOpi8I6zbEt+2IepxDj7MVf/RE0xT1frAJ1KuolJEpxuqRKB
AIPeXjx9YoWxQi8pgz8BJZY47c0ZyyHSAE6T7NUvtjQc3GwePnxJ15XE8PlqBly7
cB0LSdb/dbgdlwcz9ajUy6bE0W0nVWEnOjY/HM5OmunHc/XsTpRSbGayPAvRIAPQ
iI4KA4XJFCcPkBKT8/F6EN4DGAq1HJu/1hpEG4346Q5S3ruBsshlhAs0OTcm7ZN4
BKFrv360dY3n4kOEKqe0L+SGOnMh6OX57RqIfzODljOdZkI0kAflLyKw/dVdjajM
GjomDNN/X8mlp1sz6wEz1tWvFZiSMKnTNc5oxYNzyqas69B2XeELwa5AvT8tgH2v
ZxOIBHFXEocRTHbNNvdDMtwTEwIe5dKdabSTjwoF1JI0Q0UbCauk3lGcSh3hDhYp
+PLFYaYnOazb7vNXFp8EMv0PU54liqUNR+XJOAgCYkCNtT1Vqof+EnQXcKWJZGGi
7jHAYsBWqvM/MW4dUMS2didErRxQSZTDPsDNf5oKCcZy1Wtp1SQ1EWy04SbiB3ya
KXxpZIyEnVwpd5E+NAS5AOnifBk/ErzZxdhtPJav3QjBslS53iskUFDtMKFuMP/n
+ZH/ypA4ZHcGnuB0B3B3fe2JgBELNuWUuZ9rcloZ0jBXSCZNemUpJE2nwPWSe1N/
jOSoKH+IH7m/FqGWQjlnPQ4gawv3LcAOxBfALKnzbj8lyOZfpaIf5Gjr+gzzBFoG
0/MiPwRUdX1DmLzwAC54rWa0a0o6spp/wVAKBA4p6t7R9eqZ5w5GbtyxzdUmNIVB
9sty5wGZMXL8rx7ekyhvhUeCTL0S1VmtCfxdwVdwj9H1hoa7Bi+51ZoR6j2dXhxF
CFq+/4mUbyKiPFNUX6xmXH8ZDZTymCQyWO9tI9l1FhAG7Z9DipkpMtbxGSB1QXCQ
CRp/olvgC4Fe+azXxCUwdaaOGDNYkWy3WVwHgxlgHHc98J7lTBBUucVuUCkHGL4j
aGzzg18SA+a5WsmsUIEJL8+wDxp/AOsJacPyeDyluhk8danjhxukwZZzeEOf77g8
2Amkj9wFEpFXoP2kc7zj+NUK4odP0raZucLR6TZMib92Cq1xs9NPi//pwtIKibSf
O9POUBZlZ27+OTP9Ag+3iQn6Xk3O73BATJSzUktV66oDw9v+vhHegmAc9qA+Rbvx
tHpmgH93W2+/L08iumriKd1UohWbahMJD3wQ6WTlO3B5NDlQDrlnulDryo2+SuRI
ZCgeTvns26Mxyi3dYe1MPLlmCWtuP2lBtJsnHoSOvJHpZqDCzLu7cklCJ8Ebe56f
gewjyIrlfiExvvE1MMq8ewJrwGnUSQ2sdceICVXe+Z5qmtd04KyquuVGwmHpbMEU
54Zw79+wUDGpwYH98BgCuP4uqF599QT5OH8+Vjez7OuMdz5I77442dnsTGgE6TG9
DIcyAM1eNBQbJJD3Ifw2Yu9QWVb9Nu+PwBvk+wcC7DGamX3+QXHhA8xk9js87JDY
urbKTUcLeZQPh+twSky2iURPT1Rgntrn8oQG9ec2AaI9tK6LkTg5gNa2LXH8ER7E
yt/JHKyPwp9fZ8oigIBnF4sLSLFtDux+ayHlor3PVJz4t8DfSTDzxN1zOsuUbN8d
DMNyx52kEU7lhVKZZWLIPqYXGbCldduuM3bQ6mLZcb0VLIk5omLX94UffvGrV5XS
ryFfkRd4H7/L7Lho394y1/0nR8u75qq65nM29SiGwDb3xDfGW4DKJnLxn0OZPKDx
pW7q9HbQpSTZ9AY40X8eUYYJrACAA69eqW96tNi/+2K9qSVQlYlyrVotCVDBSvmK
C6TltAvTc6c9wKqvjqCXZfiURVfqf6qNIXnG3knQIuq0X3tcwQGkHxyc9VYLJalg
LwJcc6dF+Jfvu8qz9P1D6qaklHpHKGS4wJrGyy3Zvnvzn4/d9+3Y4UwQrCdJH0FC
LulZv3IWRY0hX9jHL3509E4gWU4RI8tgShc1y26p20Zx+9Pxx0x85ALjP5GHcU9y
CsZoRPV9MU3/QCDYcXZaVOve5bG2PsqWTDP9DezP3oOR32nNQQADt2rR6oD2g7Jp
RIJjcrX6CMRq6/s5yUvPlCIAiMNlZancq6qOIRUJrUOD0IP5O62vNWduxjlt0GtZ
BzVLeA9WQA0VZjVr68jtWTPsok7bluzbD/psGq80n/ImzvJvFN52xigIjYRFhDDS
vIZcp0Qakh/rc8mPNVGK/N5CHmrbACjvaIB8yHY3zzYA4zi14qPLY4y8vjpz+UF9
DuTT5+cRpT8wfjOuwBpUQ9dsaukYFyrvnDCYOh8xGZZhrHRDV1BVXlbxE1mJMr3d
Mr7SGH2WLjIk/2/SjnIH28Knu8023GGopSnMMzcdyBCUyXoVpqzLs3lOpqBMhF5t
+XuWtNGav2k3xS+md3OEGCR1XCnsYUxI8mBwUCp25vwxTqyyJK+oec6AlfNdY/gH
oRZeeCMYppEj5n39AhLrnL9FiBU73+aLk6i1Cw8eY7hzRqnJv9U8oyGVAkogLxKT
vkL1Fwi74iQqZr5fl+VBGpcp7KlyCuesm241rRqDUuVghvbxr72zasUGlTcWHA2q
vNRw8PiEb8rbaFAD37IxwNbq0CpihkPWdShDORQmtyixDYOoAsRBaarkuiBw91ct
nMFxVgLWO4gZ65kX+03vXEckX+EtPivViNW/+Uu1uCBOwhBESxTj+8TZ398Zr3he
O1YRsCV/jP0/kjpdWZag5LBI1lnPDGIUto/j3QRZ6xvsrLZatapYSN+CSHePdZbB
e2rkm/UHqvNGrBUW3t/BDQ683JL4ESJ9p9dAE5hcpK/W3Z3P4fAKUjhJhCSfwBrF
mpn6qfVZwJTlgN2aWrVzAooyKkI36ejRapcwz4U2cERzYYhWLqk24wum7dux87m9
+LpSahgpck2Wy66JFYDs2CyJ6V9XVFxIFKVrbvWp0pkW2j/Hy6pp6kjaUP/dbpd6
ssCuFKXe9Q2n4JDjbUn0fM8uhBx7xu+z+b4oZ6OA/ti0L7xt6kkEW64a9ROOE//e
vpfKbt/Jn8MpmDO7+Gv2puqKjjRSSEkLu43o14eEk83xLXZeqvsHwlTn0h3yYe70
X9sqP+jAwxG3//ieDz/GszIScX4Q9S/0f7lOGQKcuZhqI4p/yEetRI5dM8kzEEkJ
txdTdIQt3XuybUhWW7Slrvo+5xnAET2em6RZCxTvJLz6b7EzGms8l1MlSOgnS3vB
mdx3xF5K2cNwYHukZ5HFJz2ZaXqu17ofwy2HL21frjR61r9GTEyR9AcJ6G6Ld0Af
MKDagKvPQqsU74ZbDIcM0MsYUlZM0XscKiT8cWSUnxNwz5BHBpKYkJQb2/V+fuHA
NmsKcXi0/0YPf3FfCY92U3fwLQlfy5BAalVTWTMXhoGUc9CPd2L7bxDsq1srTT/e
QuJNA7uVcALZuGppvIcq2nh7a60dvXIk9zGjz+Ib4o/rGjsjAtUpo1RpFBEjcnO9
xzvFxsdx4JZ1GJuNTZ3TqlyP+Ar579mycryhdYATqNDoaRPlKioTrHFlycWj7Rjt
FKsvHp34Pj43x9p1UteKu+rdINkMbchly5w5qia+xxrGjUjBtpsYPVmdrMJY9VX/
wWSpbxP61yXIHyjgq51NZm5W+Ylgu5Kc1Gm9VhZtQoGBdR9hFhqvXlQb6DYKXLRO
4AX8mXsVOwokvDuArs5+U3+c9gvpfkixQR6WaaoQGbAwNkqSGRmrmYBWG7SUTvde
tGseJovmt3OJVfCQ00qIIYYiyhVesmC8GNm4XMcSTH9PPsn7a/HhSh9eAyzwoGHH
2iWWHRNCRGWkcW068DAyBnPhdnNhSX1JvfDGGfzV7OBuwdO67qUeFta0W778NTAA
KfYHPKGg7UuAnpQq5Pj9qkw++fepNbzgcm8rB3GOLyywOjVifFrdkYNQF/dENX6M
ci9uKGXDWZsNw9+fD0mewUI0qR7Uz1IzJYHqiulZC2mmCO/08TqcT14l8BnwRGiD
f5tsppse0Kna+pVzBR4ncIqNw9JEW/mbzrqrViCfJE+Ijf3R7UsjfhC9AoSEePqW
2A/0e7G94ZyXV0gmq+6HyKUoq4XtEP5azqIyg1WeguPEAcWvNUGnoW1y7qeKerNI
ofkNpKAJJlmpNVl9hiXrWMJONM3WxMqY2GCAwYKb1QXM2opBrDlk9LOdwux7dqDX
9L03MLUtg5V+rrsmqd3Szf1TxsbU1QbMNJYv+7c/fZI/AMsX2uzD46dZy5GmcHOm
uHMWNQ4Su0+yDevOtzk22bZM/+rZQaNpxW6pVW+tevby6znp5MfQXF4t4IeqkJqs
TE67KCCiZWzACA8vCPLO8YNPeG10TF2TBjiQUYwL5Ye/GPMNtn1BuD70PIBFAubQ
58UJG1HW6a+IIxDzYCrH2DKRl5mch/35RFmC3httbT2NSyHnrSqzfkg0eJMk+Iy2
Z0jAGmaaVrFRpodhrmMwHG8xZG9eWuNM0J2X/rxD8WjCJ7Pl7X8NwjJ3UYUjcJrp
IDqZjvnTQtbyB1/2+cAd3ib7A026UBD0QA+MDoG9IT0VZmVOdoTXNTT5BTSh0gYG
Inea/zHfWqkIwDtfDk3Uin3XbmblWRbVcKBe/mRVj9yinGQnkkU99cXN/9flT3aQ
6oknjGx5Wuv/zNrbgily6+l32PZEDKTIHUCOWdjQkFjszPFLxnu7TxOxYZrLKD9S
e63et6PUVsfLsQFvn4bbtcFnBQV950NAMIXaoZJNKPxXULmr/2rKP+p6H8kd0V5r
F5bijS+rnPZP0EXnK/561ndpEYvQggdMaK5rLTi84Yb0GAffGyZYz4bACYyWu3/t
XeSpkDZrDT66OL7HFqgx1fIJALxDd0NU+HwkDor5CzLg29b3txZd2ZcAOSDqJ5Bl
BKPOTd66mmWKWiZkcSbPa0LHOTR4kGZ5Wew+SFcjsIr1th+yU+bgOA0G1cly4fhh
kZlZYMclxLwzjyJPruQKj7HYAPI1/xu+J+HB0wJ8kquGrxpj3iVPikT62BeZBuI8
I+AHk9P1HEV7fb6j0w5r8lKKaq3n96fMPavA/4/XqbvLfsFn010C/oDYxKtFRR8p
DAmZsovshG9Iy3C0XLKUWUg9XKP3vt9PEyYNaJFy+T+MFlUJYx7V1VshUxzutZY0
VCJae2X8ZEc+0lPSxN05UXbf1fUdm9a8jPcodYWLGM95mjPs5ZlHezwXj04CViF3
ppb2vswGJlsp7saR45gWmpf9TgY0hKXb2pWG6v0ZbSvFdj48iBEW+blXZknaUZj3
lcXlOYOYSiRe4qvocS1EAWfIInLzO3+k//9euMIkA6CIlmtZ4Eh006vNeyZzatTq
l3Q6fUfncxLI9A/1lptDnT7rsZd7HvAYjzgJ559nmpPFcORjveZ3uiICBxFfE9iO
GGrpWR2cmngfaWH7bJZImErM8aiILLt6kDn2NT9XpFRddMVKQ1Aakb4MOCvxZvph
rbC+FlvILiA9+y2llrB5SbQO0H5YOF6TwqBJVXJuXkG65oZ9+gparqz1oSkcaeI1
oT3Ze8bu4rG2jAoh1b+Ye0AuFGOG6XUIY6G65iwl6OwM5tr8cy+HvKMx3oKMTiF+
7u371DMTZnAnbcRXIaXJIulRmL9o7CtSLq6jNvPQr2mVXA17WPppcIhbPiNjr279
jaLzlLR5ZNq0DYmxo+nNqhlFWmCXSy9Cn7+BOm9rDl8+DJeD4ktApWQHuyAMwKzW
MFd8xjcgx3Zl3/x9DYPObh8L9tlSI5U46/YyQ4qWxzwoyfdT5yWHUYOkEoQM55jE
oI4DVwmD/rrqzj2GzSJxc5NLzBH8+Off9LN/hUPxjWsFe9139SfwmJnKbT1uLJ51
gQ24EU1JiJWLBqHiLPx/0ajpYIom7l4Ar4dbO90R6ZeYTlKpz9/CB/yyaZ667izm
0T8iIN0In3OiO14F3oAcb0qIRz5mbioZtdLlMww24RTMHU0ucPLWcyhq8pm2A3Ui
7aO87EY0Uao5JJjtFgziilSWpwEwPpocPwCbEzhAdo2SxlEYDh844TPd6qnBHkWo
ESuGL+rV4E+NADj1408TTePcHIQ6ryUeloIQqU60b8c87GagTCFocItFei9ZM538
QqCZHOBgxErZOzBnsl+s08/T6uXjIpmRpVGdP0BlIltLf5UqVf80HZMHTJxa+w5q
w1w4beW03TduEL6NRxXrW6xZE5uuTSE4p+w83+hucAi5thGb/Pd0FtYPEGfBKWu+
ZhHOyvZQErA6dhQeCiuxx5+XQXRcguNXgmOJJH0MJj+QLpT5XOMFJLeg9E9e8fCb
iQepAS5Kl6VyjppoFfN8xVX2R79urs28ij+bNZQVbJhikPm22NzzF4l41cdQ1SDx
BXw42w+orgGTQ2QY2a5kSZwBPF/k2yMAoDlMNrXMHebHAkVViRkgJk/Jh5SB5drc
9rs+gmZPOD42ppA295hInqrDChFOEcEw1fgmOsl3jnxRKyb+Fma7CiJphw5ftgn/
CwLONq97Qz+YqgLM9SRLwM86RNViFN9rqorq6qcNtZ0o8MgZ//sfDAmoZ5a20UMK
80LwDZ/rg6Vli6IF/7P476qtPWEsRYyhowkVkLy+j40+H9ZpUvCyKcPRYGxRENyG
wWNbizNwn0s028YF1GZINRE3BkryTNo3DYcFnJE6KXVxd0L/k52wby3VoOF58045
52AiweKnNNP7Hy1tJ48sAxbUR9Rfa9haQCEitqFYcUZgTf/GgpzC+5gqufD1Gp+S
HtIQaVVeSD1HyNzjRjTy7lCbOgUg0ks5nkeZugoWr4QaVeTWmr3rKYCVxbgPaoco
kZ3GmOXQy/jHV4llO7YFr0olG6iCuW74Vi2/xmPWAd9TYIF+NX8/poezq0Y8sWRU
H4Ghd9oQqc6q6FbM6dvN3aIbShoy4Fcq+9y6136wHFfi61J/q5b6QHSpkx7qwDa6
LxdD49snAxXDumifrGzXKT2WNqfymp36RuvBxAQN6E04IbiXwTaHnx6/bD5ha3+N
urFyKBlp6Pk75QXA7RSpPhcKpyRvpVjWOKyyi/qVbSqyC23FrVZkRIoSvps1+yLp
FHxUov4WkoSVivBpQZqLJLuNsFAZB+X+DBhzKEtcMCgGsSKFT+1S0ThkuETQ1YcE
Eqf8+FImRr1PHMVg/UTHDMKiIAKkYpK4lsYbBiQI8ocPiJLs60MHxABVzHXXW2zC
PxM2W/5jb98rCmpQ3eCmlBFNbZ2ehKyZ8XcHC+K+++OT5vg5KXZx63o+wv9IyEfa
l64GKaB4uzQ2uH/J88aBHeZUjH1wIVoky6/emS4lt4hnPs7Bp8pfn3sCljHCiIuz
ShPFKE4MqCd8+2DQk+sVLZxH56AdygxN+kSjfqmFBo/19is9+IyyrkBbihrHYZU7
ltDTDAYODSrlCOZm+2YPyvLeNjgYmULdUgGXGQpJn741oyrgyXb2PkE4O+3nbd72
z2WdqyyLM+nxFMS4dG8q8h2eu56qrsGH0vBlUC8/7bY0CGpWe44NOmQY3sp0l2ea
mOop/XyoebeGING6mZ+rmO+KY5/nmDuCzDI5OSazor4bGUXY0RAwmtgDtjTJcPcV
UXxuQMkdQhd+LqW+FhcHg9NMMEXFNA5oqTFFhMCI3bDYB9es6L6uynvQJMoqPD6I
NoovR7l/c7geWmxdOnDmdgmw7FHAM8+uoy2RYMnbtCU/RplTbyYbMzvNdGKX2N7T
oJ0BGlk1tonk8ZV03FOe+KrJJDtHd/7m+jFBViyYXIWjcroBNpFQ/2MX8gfmHxwo
1cpVLiFykckA2uiD9a2DxS4ACbptB6FhTNikpx+S3hyXJgVGvTLWKKJPceA7P62w
4Zy3ITsq+O4CB+9KkQca2OtYMw1hh++WrrklHuIdhDdKYHKbmJqB7wBkPvEPsJKf
R3saZa6Gnr8bWYCy4cE2kMCz//bnsLYn2VrxB/uqLsHBmmbXZfw374tv3O7woUEh
+88c/WgBQnmH1ekDLzuqO05slzl6CKnywGj6WcWaqZnXiyWqwOiMF7NAGLRvT6A0
pYociLb1bxcu5FEivSjllCdx30zcuAUTlQo8/yg1tbXZEVy2ZxpFP/yExlWIOdJZ
orkMPXfc0phSBdm1ajqlNTMC5r8jScVVYlofE1XG4QrPWfkJPM3ECg5qBrdm+sJd
CdvnbWBeOap6qvRVmJqatP2Fj2IOvbyyu4go/LFyoUVSISXKP8imv/DUsa3nl22y
tTcVztlicLUbCAPcmKrS4kpSo+GgvE3gE+8s9W11rBjcKXPnu4AmlzzWjH98bWss
QemDH5KveqC8PjLFxuS0zDry2DCAoaixeg/5cEmaXBMGQnwW65KTjzfFM6/wyLYS
aKQL99n2UQ+xCHUU2yUnQXAQd9Y4sx+WIUNPjYl3J8mbJX2WNvlucURLGn4aQNMj
dTYhIjK+uuzWqcxUSNkTEFu7KFSNrefPfaow4yszTIFV/fDKvoyP5qo55Rnbooe6
/Qo3y+mgIcVOrNnqSFBg8DsJrfLWndD8mULhkPkws2kyi0GLi+e/Nqk46XJqPPpB
Qh7DaKjwIxWU4b54cB2lOwqIucLXlOwnks1wB0LNf4kF3q8bHf2/0DiF1lqmcV9k
Eqwd2D56tG3ZwjY9/zcs8+z/nndOIfj/uvcJqRYCuLfIY0FBmc5yL6HTRBRsV4AF
etif38RHDeblpqDEOKFk4vo4ycoMTdzE6J4dnJgpQoI/RLr9nwrlQ01PI5iyKxw7
67bT8HWS9peel4QEwRpOTADynuInnmpfewVaeLagnfnpHHv+LgV355zQ/w9eGGJK
4G+ezmEdg7PxzRiizFjPh0MC5lCO4l5MwFcpFTcJSnK6RC2YK6hXSPXBlsWK5Osj
eOTNOEJPqTFy86azwKnv/RWUH6MddiSmJqJfiHRsFcFnxJ9nmcLg6lC7lGvuLWsL
nv1dBNs/jWrSXLYST/ZTYNy2CGD5eJ7DjwAFSu3eRS+6dfrNSqr87mgQw8Oi9E/9
vkg6By7UBY1lpXnpNCrrlQKT6Z2Qt37quAHPrFUgBElcOge2nVYYkEUHSATcaXzG
lKsNUlvyYI48UrZUKndCU0t+1Q7gCFThRC9Y8P6Qpg8WDdMOCGJMz4XEShTcPW4q
slNZAAGRFxpoHjSBmkYYnyHklybgu3BiQZnSZ/IuXUdUkvDmP5MZZqUhAdJdvBdu
vd+YqSRioEpFc0t9GjFkxzDAqp3ye5GpY8P3RLarz4USw6FUjvpopCo5PYdXX3Mt
wQEEZ40EeCBAMsPrBOqt5FTqvsloR2pqGLiseYweplA6F+CZvYTwozsaaJm1Qfii
et/Pb6nly0OsGMMy7sWCRzhqTXZh08hBrpLmk/6ygHioj4rTVn1+a1EJMeXOEGtb
BS3cSuHrqG6Thbalyk1qc1eEcHyc6t+IMbMDopMT0sVz+PsSZnuZT5v70eWwNQ1r
M+S4FY89V+YhLjUXLyYcvFuyhF/2SFqhl1f3GCchn+hYpYFW/Es8i/3obAr3ESxz
rm+vbc/9daVmSVWFXyVjM93QPEGG4DwPkzf+ksj/stsNKQ++3otvh3S0xCP9fox8
qu6B40pnuUab/Z8fRp7fN51i5BR7yN265IAp8AOi65DmyY9vGUKloFsMKcLKc24b
D/tbFDly64T292QygxrYnFLfW7EgAEf+slAWbtcdNdSiCfvz8rn5L0z1VwGwGFwT
nFRe6zMooisGODg1N94nFsSyLx2mNNattRe8AUlPOzEp5G2bNcml7hsmtP692CjV
2nGbpHqpgr0oQAPz/RPzyPyCjhlLl3zvENy1JtJwTWT4anb8fVMiAvMsMqLSxbyG
KGE+x7blgJ6Pc6UFyd0upSe0eCXgLqNrVR5g7by6giQ4MquWrlFZLJdhTCqfoDjd
zhMXX4b+0IeP6Oraj4H6cxcsfJad3jbzcZvinKyQ95uKFO3CHLvkQtOs3qJara3D
ipRm0kaOkVy7cLvpxRf6qQETqI79NqLJsbWEyRC5GX4FSIvomqsVNGqBOqWMruT6
g4RbzNd+rcvnUNq42Tlk6aQdvzcfkOt1rP9rqwqpYft62IE3gg1m+/SHfddf++oy
b19/lOWtKB17wngWfq4j5yWscwjb6hXD+VODKBHQxZgtm6sjYUwpP+FzWbzN3QCI
oYCJCI1k/hI9qJ2zmKW6WMi3Iy6tTMJkn/5na0BNAnwhnXHa6Gp+ObU8+iPK4iM1
RkTidxf6X2s5wTnRhny0C+TdduKeiaNmZs5c8EgI4G2W4BJORh7qI/ZnzyoMCR8T
ggpM6GpU3Px2GAMW4usIrzMzTGrsgGKCQU+EECbQspTtxVI8Yz2YeaS88zzB7uUU
ra9NF2XivQZqEBB4gbjXpGgs9Zl2SiVvceVcH+FbKyTa16zT3++baTDS/PGf97pi
6aPmUoxko4zkPEXr9bxdOGiFvKovqxdyJvlPY2a46k2gqolYXn/o6BzVX8kDrpQW
cb1af/em5PwOsKQ8DL6w3khdEifcjNC2XEuxNjCpqiiulgbq+1elmIRsYyx7PWEt
ut9hJbiLrNiE6cJF2Hq4vFvR2yq8QK40TY4NxwQ36wWfQtgqE3Sw5TSGeWMz1ChN
fiJ2JV0ILBvHShEj3fR8uKgsCLL+pYIS+PyNW1jFmVLid1jTn+F25Jumvp1z83C1
c/YB16H4hNxXp21vOTJ8jgBKtwhFZA7NCKDV1aX4C/qVxnxNxokGVgE+x6gMTalj
euAwl1i4i+Z0U8u3cjiNinBfpqeIeBJALBSV+YqQpgTu1Big8KD2RPd6s+L7KOrY
DAsWpSx+Esb76WndSUfHKlYMGTNm4FYMlGzWcgb46e11NJA37rtqjXqvuGVekIMv
FwCGjMaYLBACyxheLxsuqibMFcerQc1uo0BTkH+uhOKyJ7uOU/gtdj9CRNznVYTI
nJmj/UPfS9YoaxAOU1D4SxCF6ZSvdferuWVJJDxuh5OLL7AHM4TPHMHOTfcW7xxT
d5B5JSoOYwcySEBnWQaJseoiqBLCGAWSoTWlqg7pTRmXuzolN8cGaVcixyK0iRYY
W2DbWMievMm9Zov15GU9zohnPxd5p60+Msya1ivX0fEmaQdhEk4l7K0ehO5UZ8N6
swWhBqwnS9ThflXdeeBPaIbkUlEAVp06VLbHMerzgbefkyzkJJ0q6Ragu9NzQwi6
AbbOHLaMEFMjnFNy0k5iB931h6s7Uh3O3eujj2VZHjbO7TVEo3vunxiZbySi4/Jx
r0fdO7wmAGeJnqMQmCvQM5oz021JNqXqWqZcyh77r8nNtmc6xaefIvcm1IILF009
AN2BC+x/9nrIJu+Q8pkHk7JZjU8WZvJs3S/O3PdihKdBfOs6G0nAUz4sGt7qyXnv
iZWN2JLdk/eemgIphhEhQvHqdKrev/K9mhW/8a16BkbijNR9Yw9SVMg1IWVGeza2
+089pwBNzFNFSvIcjXeoiV4jIzA/EZNUtz+k3JIvEQhFGLneNfhjCYog1+dOhK3k
Nm4zJ6cJVV0YoPHRVy1vtKV72WuE+uu43ZddTf/SBghusP67tMDglxbExV4dCvb0
Wgc/uFMFsBDCymevShdAQVjcdxApCvgutbk16nN8XsX5nULbsvUdDXmz6EHm7GiP
jiONAcE6RgePrYGnITBn9Kl5v7eWaqBLCIRnWkRiuPSahpe2DJJAqtoDNfsODYj7
/shUYQ1dto6hSlBwYg2g1nHnou//srgOfTVNL/wRdz6ye7X6gQdRagJ0ajSf3Adq
B9iGpOV11LiNjye6P9UXaRzZM+Z0Tf1lpg4x3rboe0JsDasH8/8LHqUkvYDcN43D
S6OcrQKZOj9lCgmPzXRxhsX7Q9LM5mZmNbaCoK0BnSeHqVMpLdAxaycULp8ijgO+
hgGL/FktyjScE0D6p1PXtXhKfE7ND2cTw8eUnF8OHs2fx+2ixMnvsI+b+MuOeMeh
lGgRJreM2ANkUNwr9tiRuiN/YeP8/fXYmBy6qVmlNiPthgtVuUPAAFtv+SdpsuiD
rnWc/kIOR68LuCpOeZXCJK6gVKv/LKK6bdtTlkaVc/n69tp7l+VcZC8uyBGGyMfm
QC3SuiBM/63mdb1DW0Icor+lUemAxCYntKlUVRwBXH5ykrvjitf/6MqS+OvuPeSV
Yhv9pSyKgMOJ7a+AnEHGbwOafctjjgmuRuyzA1yn+7SaTw5RexEUuZv2WnFIC2DV
Ob+kVEaIVDqYuAGXNE8xf553C4eOY+zvva8e9wSiWekHp7/vE2YK0cZsKaa+R7xl
AxZFkGXyFpCXCGEBTrAqqMaA6LVScId22jvt99wiDxfbORecpTm813X5V5dWMk1A
7MKJOPRVjaLDOL9t/P3k4EMwGemn1AcAxHRTjamybp6NVzh4e00BPm0O/h73xwsM
W4U9XnedKqTS099xIDTSCFRQIFDfXJL+Vi5h+ZfvYBO4D4bH/mPBtDoKofFcSGpT
YPosjazp/+c2t5tt4Si60bVy6YUUX6b+oNo4W3/BKX4cfuv+Z9fJGedWxn1uQ/5h
8MbFqnVYStzlfcxF0SmI240ZHxML6334rxylYZYVuBc5oJRj3cCNo0kjku7Jh+Zo
PLNs3GZkjMeWgVk8tQmKIGl7nmUSVt9Zh5P1YlDwnHeelTbDIlpIob3/V+xHt6Lg
Dy/9IXMUa9Ja9yEF71upJpXd3IrbUsFkf52hz2UCHLNUEXL6qv36kCkm9LWO+sua
LseBXDbPTlO+F4CtP1gZpCNQPH18hLLKrxq7BicGsaf6dqB4GGLYuFacjlKnU2No
muj+voM/sZyyrMfWCtC3Qeug8zmf0FcraEIbQ7py8FqFGZpd4RcgmzDIfSma8me0
awWovN7uWN2ok4hOjeie5qKpEkavBaCMNe0kg6oZBeAzH+rdLN4YIfSNkV21VtZB
hngOLO+vqyqEsxynhElS1MAHkUuLXuE61WbyuzRpCZoTTRl5fgZcOuuFvfY7XuS1
JrQ5ahu+CFfJMqw7zPitpUpo6L0/GYMK58xzRgVkwIEDL6b3zyJ/BU3v9XPptmZf
gCZF/MyiIhnyTmYGi0pMJmXFphDk5c9CXUHxIzxp8+KIUyMzhVw9FiSpgunIBNuA
wcugqghoXL6YoazZYWyNRpVuuEfiHhvCRD7Lsqsz4bndWlTaljYKX8Fxvv+bkgJN
9kUIyd3NBkxsCWPP9Lm0oVVWNfeIDFSojvLb5iKE3dFXKp+UEELL1LsJi0NqxSBM
2yXqEfJdXLENCCm5546adLRhoA+r5naC7dilktIGYCJni8oV9FFI8ABfgxxXg+4w
CrMH/FpWt5G811SoGIgiITi0XtzsK6x61RmUle/wENKTfHibUSjVBI/cvLXyRPsI
Lqdp5srLfK6GIpmLPLJzMfr9D0kJW9RH6SZ0T2FKR1JvIa44mGON3g4ELhUBLaKh
oNUah3fJf4eg83AI2tSNGJGuidPuoluf8VfUcglx1vgPzLMA8/9vAPAFQ70PZ/Tm
C6pgpL4NvWPjF2ijIhrlVLKpHj11rMGztBocnsgAWWuZ62SbE9US6HQignFF6mBK
/CTSQ+kZFifPICBH0+zLKjRiv8tIYL9bFRya7/LbHnH84Cn9OvrZnCwwaZC3ryjj
lSXYMBt+F9T+dHxOHEUl/uCB/vjy3pu3WOrIYNv897Y6af5UOhxne4rf0V6L8QVH
vK2Mnt+MV2GAEwuwLHs5/EsNvF3cwdLtKah0QFKYoiG52tq8ul9LA2abLP0wqLwg
CVcDBPxu6kLNXWrPBAih70zmy13Q/u9Jqo/Z5VQyLFrFQLrb3ajuomMoNx+zB1xs
6EsXLEd2WrZd2CaJaTXMQ0tZP/TJkktgoij5A7fwTt9WMahBdXAJ8ZbPxc7fDtQV
wgOxFojhC56nFHd6qBerXcgGbFqgbTrDh/q0MM/SPZ+RgD+RYf8YROds53km99U+
50w5zHyE92yUlUjKQR99HZ/FZ2Smh3Y21DI1O+px8Z2vjJcQCjeR8rVz2Q/36Xmy
W7g8GXtcide5Dps5AZ06txLXcOtny5MEt6UXwiXMTJRb8nvweRRTtBpW9NBcgz+9
Z89zg4ehQFVy9+QuWob6b8BAae2CJgDFH9VSxiJ0V0UOFbPinOu3l6ykbCIbU+h5
tpgAfwIjQKrTaSZSQFwKNDa+riRzw4OHoe/vYYfP24CZDwDh/8FcBK5a6K5JMYZv
DApSZO2hLuE23K50LbAlfIHIzzuyIw+W5qYidSF7fcB58hAz+eCijV6758P0m4ov
Ufu5SpPqM5rfFRCBPnARypfE6i4EnJR/JBp8DUTm/Ha2/GYC5bSc/KjFXCVUmySi
WaSxZzEc8rZq0Qp/SETm/jm4MMqqO13fPm2P6MZHC+TfEKYewmCBD1qAufIBvO//
5rKoXQX0A2sxIzV+dpqyIpKicoXh2mGYW5+66irqCldZA5CCBacpKpTP2GovyEDw
J82reHBEGDoDmuh6oPv1zUiP2yUMWKJFS/feZdA0dYHmJOplUwf8QSAb7sK6G3wX
/tqNvEP0jakTrzR8vnHMXcHs2bavMn/E8QD/Zbb+koTa5lfnzqWEaTbJd09UguiS
sccCh4W8fGkQcEBy0yCH8PyTwh+6T562ZguN0P9SlogTWzbfwib41/7NTNsdHLDG
5g9rd8Z46y7tIyFXhrAxb3sFYmnGtBLJ82g6EMmaAyfNzwLDbC23IaISM16+UzgE
HVVKXm8hKYXfkJTJZZiErREFPvPxbJhtZ92jTo38dlQOPHKK1ZEhUmmoN4w99F+Y
RSN9NbCK40UnrhVHzTKvcioURMC6YMZ65AhoYOddBrURsJgS5HV04REWEHwEQx8s
AjJMMhQhTA5NMvS36w6gWPvzyVTJ79LVF4B8OxMbnbt5VzAtTbxhHnXZ+suXrHHx
E+JyaQPOkHmeqYUgY1N1JN04Orf0RhZgEe51E7VpSJLbXEGhVwZeJfV+yOiHs4Q0
oSwb7sBPYu4l/AmuAbSfp5C1qUtTOYNRJjb1kUU6nDo1YUJInPEVsq9a3ep7qDxi
Iuuf7ac3aWHKzQP0xxryGeqsGVJqdRL3weBV5WjXTJA3vJZoJf6pPPDBFIEmG38P
bFaC2TQef/kiHZH8AQ0mnX1etbjrDA5KfExyMMTHreLQq4sQHD1wY3xBBTOwbkl2
WDeMLGx5oCoH5XwTrg/p560r3BqxlZx0P4LpC6towoM0mdJFvFlqN3scO0S/gj0x
XQo6EDiY0STzeRwlfQpQPFwZEgTNCmRV4urTOhuZa4u7RR17KNzcCyjgVdkrBuzm
pb/nSMo+yyCLMjpKNscWxfqk+m/q1BJtVNXDJ0mkHMWq/x9SUaoS3h53mwDNvjHX
S/o2bktkThEHR9CgXRN2+kImvor9rARaPXuCcQMmSeGaTWZL2imhKSaEkhyhS4dc
hVh0rdOtWgxbDB8FCwi08BXjxxvyqTASHT8ecR/FIAd/w+/2v68z4G35Ur0D764a
s8zMtCdRICRN/KmtUKA2arF6sdCcgaE4YC9ChlD/VSR2HM9wUonDlC78/8h1/H5p
u5mk76XT07Wr3+BhJff30nLt/i1lIL+2jZCIQQ3D5FbygjfhLH6taAKy/G4vQ4/V
sFANEYP4uYiJ5UFc4QI+usEYy/V8HP4+D70FBc+frbbOQadeyMYt5eVBQK9UAtms
dB2SnP5bspHOF06mf6py85Ewxv3l/4UBy4vkSU5U2O1VCcA6Zy6jIpzhHLEEXTQO
o648I9z0yTpqVSr9TWQnxgfX8tN8H5u9dYP+0Djmgl86lw7ZZBMJn0lh7h47cSv1
RYLtUt9I6yfCpIn6CTg9JJghL8oy0GDO4mG8qHrb6q20f6YqTzyq3Ogxvtfw79dY
Ru3K80QmVmopqFKTYvimXN7WFlFAUjJwZLV8g+pUhE0PA2xmVjGg7AFC7Xwlbdn2
1QNIqi8jtNwdhJ2dUDFR4dJJtfeyhiDK0bLLokdmiHWt6AcJcl5xbBn/nGioHAB0
vmeoFVqImW/+wV1lsaQOWc/3xjhICBD0/xy8rt1obR43rChqXNndpong/30E3K9x
apPLlCSZ/3JbuVyUuyuCQcmzDgUtDdCThYAWymPk4fK3CjhP2v3JNL6rgrmxxceL
r/p7jQYwMHI6JEd98KhmofNx3p0r8vUtt6vjq1qgzC8rN+812c5BRh8OoIg6vonO
VBCikdcfvncFLDR2FlPH7Di9sywPvTLg00V/5xCwPc3Gc5dCxasV5QlQPpsMOZgh
xIc2LXHcnhCppSsaWuFFirKeZHRlkJAS2eD50bCKXXm9x5Kv0eGFkIHsIqgzRbVs
92sJhWpt5I1inIx1m7tcORpXWbN+805AkDl/EfJ7x5UoOeMCVlMl935SI4J/58q1
iNkG5pdEwsNIFrXx9y1VglAzfhmHGqUtrKE6+wEmmmxHYdjQxgZjMqE8DF1D0jgH
ORuKQp0jQPap1d0RaF+mLjudXHwHjeAGRG+xIPR1tyYH+bNQew+z6EWf0wbnZai3
F3X8tCRdUiCg9Ybk8GEjLHS74TattrQ1j30KBJ6yaxlZV/ECRm9LVScBkN3ciy5m
ka2iP6nk/yTeOX+pHgPqTGH60SgDa7i6Ronaq9gLWxf9VknbkrhhzfScaSB8+xUF
YZUz9DB5BKH4mHPt6Ik05N0eSQE7tjZOyp3LSZYDCwZBJCRCBz8QLMG66xHsA8bb
7CqmWvhO6pAsfuvKkhPyVy9WdFCYnimdItA1eBzcxyL/cInlPVmH9iSvG1FKkfUl
3XdEH+Xci8eAgWkG0MQlWXA2ARRsTAXAuBw06Ou/TBkdG+eNPKyfWl17gyb4iSDt
AX1WYWFaupCUXHGwkoYXpkCVg1vPB2LhvpfInc2oLJPuLLbsdUsbuRP28CVkbNnd
OeM0LaIjv21w1ZcRyePqn/6pk1jnsUTgRoNwh1qcf1QyLMxn0Qyw45HuYgIzd6Qi
12pMaXV6gnBrhP1ikwkIampQAkTUXvJiI8K8iDpl0rKoRgwLVB9EAxp39GLXBDqo
9rzClv6xHeUYInYqZUvADmRfIaUAJJXeuXw8J2u/uWPmw13r7zffFCUYt/vmMpQC
/9kvVwhl0D7t5KgSpyTz5qlEXZTaONbIv/XuzpyELSEA8eCsabHqpfRIR0l1Gi4g
MPHQo+S52VEzQXta+BzVugEp2G9AHcp/mR1uI8viguREna/68dG7UMWlcxai7wFn
L0275pVitLjWrLJRFiYoIZS9Sv6q6AS/VDPryR9Ur5Hqax2tjSKSxmB170JmCrot
ddKgvDLIefVr1+KJtk24g0OuzvFqiQP3o5COnJeKrt6Tc0+KERoG6XVoUPhSjbO8
/J5X4sD+KO59zLJ7vNSGRV8AmQQmyRZjv5v66WhNHiIcCmVLIEfHxxMAmXH3mwf8
DXI21RQEKfmffWhQr7uHsZT24jrnQpLSAC6jX1D7Y4sfoRdNXzeBJxNVbgG94j03
vCTF9sQ93/CSgFmWwGKdSzMm8lN8fl6ohSPZB1EUFoW7jv7KWQwiL9EZa1i0Yy3s
eZxkkCOXPtKuLHgIwLLF6xzvZJyT2qGXPfwDBmhSyBuX6wLZgQxSk+VDBQNe3cSg
ewMuyUO6om5XlxP6J6QSX2C1QowiHf/ErcS05uUPjHfaOpkGaswIsbV1yDSHeRqt
iioKOnnkeNyWd/MKDImhN+8xK3CqtQzV6p5NRCS1jnHdY2HxL+FEyuL4OY9HHmh0
rs27EIAUqDUYyKEvyzXfCXy1YfRTdl0BgYrJvNfJbmt/igYf4hsKWZOTWL6C1BsD
hN7UydIv73gVKKuhyHv0WeVgQthkUIXxTMvxLW5UW6Pd872JZsp7f4Si5+BUBGkD
9gxDjyIK1sd7HarahZLCiPI/HSVCn14CMvcFvn6TALB1KjezxD/MwaoIoyMvXyPJ
0Vb79ZBba3TJa6RT38QDgvrksulOlGiAszZHCUfe0kGkSkPY6li/Uaak7umFZk1o
YE/NY58TnRAyNxOjfDF9AAmHTLcWb2kNnAG9ZU/PgToXY5cMDbfeOcNQq1yyemg0
lxIsQWde9c1e/oWqDU2TodTYfTAugYgMKGglPs5sYXbQVNTPbSxSTRw5qk8wCotn
D5Xuj7l3OJZ091uc9YLplSLIfEbqZKc1cK9ghDDVAuK/j8htEQoq03hg0CoFHo39
3jK/k//0/oFB27PLZSiEtFbBkHKfOOa8ScW/TfOtSlO2JwTDXrgcE73Rk78sOk5z
PLWvd6UvJHxVYEm+q5XVOPHLn5u3ymKQ6OR3h3nUFdqWU5K6qMdI2tLfcAYlu2KL
uitOiBwcEGFQqzX1x+7VrP3ZN7mP95W9S0rszu/a/Zx2gvrscvsmvTibwBSFxWMe
uruKH8qjYrVw2pSgBJ2s9xbTElFDBt8R94Qjp42a//BWUQVN54bSOFo7bZqgTnlk
lq0Ktzibo2As3AJ1SROn+xYi2dxegZQCJByIcBvHsj8qCTpm0YbjxXNPXxe3cP3f
Zr2S2fVK2kmIY2rRBsghKuZ5iu+QF7kuV9hjFmwsRDU8E1wjxygz3U+o+er2PWMQ
jM5MHAw5A7q7Pspv8/wYLjCrgKAmTx540MlA85BPs4egvNjXTJ8SUQ1mw5eBLXsb
lryTjvHxQXfXBJdi1VAx+4DJR5KYOopPN5QiaXRZUY/P4ho1msZkvW2DyNy681ZQ
yaZ+AoTHfM6ideV3naJR9DH3zFj0lmfXH2kRu/9wjll+WeHtu+2peEKWJ94t9yeO
/yrh+YMtLJjZAQFzQGtgxt96WvlRRejERjcnzPhlMZajS52irCkuZRuPcsracI5e
hFL7Md1nVhxjZrGqQmjly8rCNghD+MWKnzC8gu2gGLMOW0dBLtkIQFbqZtk+xYt1
KL+V9DRR1nbmsc5+lR0Fcjvt9lSqNEYCqVvaousWdwvHCucAsHPYhcHtxMvSlfPM
JXhnv72LtzjtmxjttvB+5qMyZ2Ll9VrESA5BpbWuQZybHFSYIMauwMSlnHqQMMK4
6Klixk7QFzyNbWTLDjQMZORNQXmJ0CLRvvCrl79W6k3HMt0vRS51513sYSiOk39R
glhA4YMwaR2H7t6uw0Fjw2JHSAzZi4ld3ertyJuR5uwSiQ6rS+os6x80Jps2EsnL
IhV7i9rdIdmxA34f1FPijgoTbA95bKN841SiQ8M24L2NulWS8jhHnHb4t1HgX1fU
DL/dyOSDzoWHaLJMPGk2d46iZK6LX1jAIxSDoQiOcI8/vi7iWb9KnwysvV1D21dK
y5QbMCNBK93BCrMjZMPNodnJDxJZ3cDssY5qG64HI6wdKBYQ2h1dWEaiyHS13m84
2bPrSPH16+Q13ZI5b4hyjF+GOXoveI0mY8bexEH8Xn8rZdwDsXj76wOuEA+Ihyz6
CRVtw0oBskuU0Na5/ID4mSWpWG87QQ0BIAxewyQ0wZRwpGDiFq0v+ElW0mh6A3Zv
zpH1p2qFbdcQWOBAEqH7kFVHRg+LxbejHCmrwUASsBHcoa60UckunCh9zrX0uyaA
pPUyA7WSoaW7D4gDwtDaU3xAzbuxBE8qZnRBiGfAc9Qpn2QMBaSFuDhRkhdfrGJ4
8rBtcho87XQyCf1czzKijUuIv6lrCRFXuoLsQymddc1z+PEFO5fh2W+qItWmIIWZ
VMRWwsbpXx+PFsGjrF90nv2dUxKVRIbxppafVAkOfJHliH2D5Py9okYr9tCqbGFn
nxjasNGkjOTO1bqq1ZPgIMyCrY70M5WZbb03j0k9do1M13TGkja7TwqHAZS8NZYX
+HWSRts73ej1p2vwq0A+6IgAhEx0KsyJJtMK4f6+O+0vHpAlbFSxLehc0b6ND/KP
dzTxlzyqnZ+b90rowL+qRnkF5ko4m3WXN9ZQl/hVUU/eEc8FyrCUFtbxNIm2joVk
Mm5uHAx8ueVYQ8Cquv+UjmzGa66hCU9am+dy2f4uYzJ5HBDE5F/jDspX9iZ1jntk
K83ZVHwMq41fklHUCDGp+lV+Q1x7Kt2qlH3cq/6Wu/IS7wvKjQNSg60vXRI3ZA9K
/YnblxXnJZ1aXWsp7ZIpIJeUcZm+cbnib6EDzT2Qpy3s0UMZS+3B71m/rlAdbkGw
mJVofFIfqD039ZTSRUBRJw5AFJj4LIgriPhJ6bfk6fe5phUuiEMQ9iW82FnM/c/E
6gSmlrPbSQd82DmuWwsHodQ++wtKNFXCekx6kFf77wTVgxlDcNUWcYk2N50lUKqn
6/g6vrukN2Vk+9gNwEmDpDC5BAuvnQU9GJIVS1Tn1KMSbFJ/BlFeMVhbcoa5HfDh
dD9hmI0DEPdxnoqk2PWi+yJck84tDFgyC4oNCu8chHquEwVAOUtyeVUCxdObsWtI
/kjcf2Z5Kz7/OK0mJopos3/59gqBd7E44p9bPwEHkgVFpSdIRgS9k2kOBlMA8Ock
Ga0Ddz0Tw346UN4rvfpriY9uEtPOw+eFztLgm0ItqsNTtBv1o1ymWslGXOtipati
Ma3bJpMe9vS8vBJSxXUv2PruoKZbBKp91hkr+0Ws5PtjnpHKq86XnH55EAs984yp
s0lBwql9o+/6zC2vTtmgkSvwxqUQQqXyNCSPreR4O8kbroJueT16OsAMAkwuEMn8
3xNjkJ7saJyUDtNHKFsIbfP585oOQvIQAs0BVwFaMBThgKEBDKDCgAWYdWygsFt4
Ihfbbto9eksvx/GwMMRmCs5V4ZmSg5HKOxOUMasTUtov6bkFREK3k24vHoDrc/Yx
l1gUGIQAKVZEtrriFUdjib+U/BeC+R+sTGzSO/NzoTJr/th8PeX4CDcUTYvtN9Mk
7MWklHL5TjLmRhMs8v3aB/nq3PDcB1RnmYlXiTTEfI+8RsnngCDBq3tvXaHqzEeo
o8gK0YH4gVzuxO7Sw5ATlp9HNFY1Z5h7OPRt+GcYVWX75SUpgP/DI0TyKtIxR/ML
j/r2lzDwtTIsb8r+2riOYRpdvlkanwKmEeMiFVh72shP4gmpAtI0xDkAT/K+v193
KdTEqWqOYRg2WF3nvyyTJGOWIGDe4CXt0h8NHaROSpFTRK9L+xBm3JOYwhy18x7Z
+CJ1xnWUulK8KnlS1NyvXswJMtUmm/Sh2GR98Ucvtx3LTSGR55vJntSX7H0MGL9r
Q4nvHBUSeeU+wDdonmVMQuz2I2xgau93WOiE3bikpM0i1BCwAxXiF/UMoC/1iakb
cGZainKHkIuQxcB9T5Ao/sWrrT1v+u2bRLKe5kl9eHXdUkOSa0xbDvBDpMLI1fvQ
MlbkuR4fHnSzXCFfKSsfusdmF361IazCzaeQar+lYXmC9zhMaWEsCbf/Uw9bMMYS
8V9cJY2w6Hj5ux8B7XyNoe4Nygyv8/TS9/uG5AGroLSRBO0/7dmMX5qe7yV8L1Tc
r0K/zXEZS8KibVm5qsjW56uK8oKeYNUyIukrAoR9T/NbgHdBDg+u6nGArROFY1sZ
bIohd6BiWCoz/r+Qiz0LvvnFroAmjHmwXN+KSse0QopgE09gMXy9woTFpATkK9I5
Jep4/qZ6i7ZVjoEJnTudMiPKbuT8H7r5oVTlwDCoDEP1c1qGY5JpWXT1Uu3d1NG1
p8tAROjU8IPTj/lfrY910Tt1agroWIoJ++ahmC70biCnFbtImOG9yEqMBcVnF7D9
xwPB/g23jOxhFpdx89cml8Nq/WgasecXW8G0eV9Ss14G/00OkpViYR5gdsErODq7
6tIwTMRxRV01/qZMVQo8bvtMk2ige2NyZ0OvvJzwSFgJZ0fIljdxP57iFSnErcgf
1dmu1JPW5lhdlDK9KuuZkmyUilQCLkJLrol5aQ2+l79o01EJYbt2CkhJZnPHnFJG
wV3fYahirPYGTuVdUFScyl2j8q7+5LuIAP9mE7qwpVjEQaIsqvyhgxn6LHJRk3RL
+dt+ACKEn2QlVApdT7ujqOZEnFMYEFbO3up0r3Me0M68ekWjPobbJ1DTxhXkMwqU
a2rogeqk+KiWFXEGDEKoCzRc2QRW91zcrYBBe0hGVNiv72DN/HDvLLerBWNQ52ks
5bICcJ3Gv/b2mqkwfovK/z2Q4xcce6gmiWw31vF2sWlKu2Qct2LQwdPsuVMpt6mm
zycmi0PPsVuD43fQZBXN97gcYTl6U8jow6eNcCsZntX7MK6DYmPKchPONE48TDLs
NXLp2I1NkH4SEtwHK/eJCotWJmg9Aabwo6SKoic8o3P7x9+MvzTEFt7WPrXAao3w
5aTYgXdPPptw67amdNkaWRi/0O/cABZ/t3ROHPPN0gKB1OAZQDzwU1U1Zftq7tUS
iUpWz8OWA7S3d4pJz6vi4KrWD0EXsEpnSmt+FYQJNuIgKvW9K7U/urgDP2tRgXFU
7UJTrewTxdGrJRlfh10ALPPPllp+hIFCbS4mSlk4lCNd726mbhA4xc476CMguQU/
zdD2FzAPgKWUjElILoKTAgaqYFEe2zQ/u+OjLwzo9Eaf38QgcU/JnGwp49G4AWrf
hLuRCO/kgtgZZV4BVFYvP/CLs7R4J9lrskV95m/PTfcsr3WiZfmROFWMqYUKrxHQ
5GJ7ijtKOQLhA4FxXigWtywfc7La8lRQXNjFuW/D2YXdi3CpjBunxST+vtZ/9aax
DN9WVB3Fjkv83DDAlPN4CTmffzNRrh3vLN5lH7KNsViRY8i0nIvnZ4YvzS4HuSpI
RPZ7Lp+FNFbrVvPb0K+wel6aGn6rAYgO1MUhyGc590hopMjCxJ0/T7adISjoBqzo
g7LTzz+nJJdsL7yH8dWZV1oNZmgiurmYSlFYaZlW+83Gr9MxEVbKlHLFv37fR8gH
OsWpEh2PyGwfqvokcAmqFqntzbs3FKjIiV2P8MZvzsB56FzPzpEUo4MicxIIOEZD
S8xY+Wc2rNcnLANMjEvQ/GNqOnWdyz3hQFD4TLsFmg4TmPkfge+l4Qz3sil5CCwM
X6SUF3ETBDF/DdlPlfl5GP/ggbjgrONtFqt4pbdNTjOOUhEboUP0osHVP2T/kAuN
rk2m6k+THrY1hOxzZt6V1uQ8+hgsx3t2TGLTqVWDVgfNIk9Tuuc3SYRsy8X5GTaM
3fQY7Asb7bfXf/APJNQ1bAUrOjoiNsC9eIGHYAYb8SljqXPZYa2d1Kv2UqWDUkPy
zqrpcPsMkpfKQEViII7skMlIfEgzTtCLq3VoUpdPSxE1o92VNMPumQZeNuc6oqC6
PPCt4dSGJI0W36T6o2cHfMYHf2fHQ7yEUPYVCwYUJQosSaVkCFzry2GQK0w1VaA7
BjfeJfQkbViHznjCiSroTIc0DSnq9/o46XWfo7h6OzgjXu+EW7NkYKE9XS6UPc+Q
l4WKpafbLQy/FiPEmD7MNlqHRicNdaUHTfKROqkXte+vTXBE0j0++qzQHIv2rrGx
KdF3RrM8jFzjtEnlFCqeDQ6GcAE70lTP7mDdUbJr27DeM10DwiVQmV/14gSqQqZv
eA2W7Xwc8h1thacvNX+MzPq5PD0+EMtfyJ9G+IALR3KdgNToOKjmPQ8M3fFMryxh
/uZzk1X53NI1dDEBHy4h5Z2ls4QWPSaFIUtusoJqJHI9LR0SvR6VIs2wloUD54XN
Ne1kwqkMYF4Chz38wOiy9oxTF3VDqkFWvmnEu/4QVats6fVoUSmMn4Nlj8hW5NTE
blMIn4BryNey4fdetU1GJgGWu52gyZ11299ZUPDVDJmg6Y3wpvIrD+xWkEiwqhPk
2xKg8YpSAK3P52d9A4Vzh1JGIwa+h4D7t/HKKEfRf3EG/XEPrGq9GuXNZ+ETAMD4
lTCp2kS05mRKQUPpWgoO5aBJQrJccNBf7WqkVEj8K+e7DTV4bq8zujIPIAqrZsIY
bQKrs4FlISr00yClNsWiR37n0YlUmMygsj7a+Btd/OfNa7eELc6PnRdJDDuRcbu6
7Cm2PNuXm+PZZn4ybcdDH3KSg6vofAGCjew9h6DgGC8VX2tUjz/F9e4zbKBdxwD/
lcp0bRq5R4n93wUY7jnmfjEU1m1FtdIymhQo6rblczSFxqmusCmDAzsxvshX2C0l
jqqJ7XfyDwl82e0FmW5ff1lpWKhpqQen3ZoM1/Nht8PV+wgI5h/uxC4ayuIhZ5cT
ojE8IeTOSlu3j2iyQDnWeOxl2WMkpKdMln4g/9y5CUHQu8/WSOci8ukojxf2UQvZ
1xzOuFtbP1h3VSPa4GW7l4n4JiUYbf7aiB+YSQ83E+NGvtynj2xs3+mqMM2dVix3
ip67P6bZ5x1IjmsG+788Y/LkO8+4qzBcKf/g+GO30YB7fKq1YrH50AQH6urAy5t7
H2f8nm27TSXaD0TW39gHpN9yXLzAxJmz+d+g3StrV4Nh3zhstguDxogajkVT7U3Z
czeIr95G0fgrw2pnrztj2Piajh6lsCKPAZn4HYAUzmNeswW9EzxNtu7aSHbYTHlb
GrLRCwNmpxNktiQlmctuinvtzIruB5SRfxG9Rdg9wWDMh3M6ngv4YBO9L8Ud/yN/
pwp/U1ox5vlIknPXfThTjNk6Zq9MymCP23dha8nNiMn01ZRgura4fmuOMdxCYkG1
Gn6kp/+IsRHBHD9ef64ctmy9QXrElB+msENb9Aic8ktJa21lmmpotPG2boG35jvp
mtVMUc/mNgYQo9sslLvuJb0/Ugp46dkeEUF4Cixm2WnVigS9lAYU6lxG2WOk8803
VReozA7m18BIO4ZfVxxj30bFgI6Faf0fD4YVI3CB+c/o6vnf8L6e/VAc4/0rXkcr
MUp8gEBIQuCGeVwqMB1Ri67LtsIdEVLyPPew7ICx/bRglOxSF7nBlddJE0RqBZ+v
WiUaWmfOVBFvslrewXmPv50ecZT87DtJaM+cr7bKQtXUE2JODOgJxhflzNZXNSc6
z79o5HzqfZ2ph/DZ/t0Ksqd8ewAkIWXXojMMlgtPERe+mLutGwKdXEcQNYu01U18
EtJPAzzVrBl2K+D+ZpQp6nub6owqjbu3Gh+sZMnJhsA7xYwnekoQxI2aj+4AJ8sl
kyPEqMMcvS0jooBBxp/1aJb57WxgDop5c2TP/xQ4tsF3d2lloE/2kPbJEMG8mxSq
RFlhRAjOTENPRd+GkU9F5PDv778vK2Ojis3jCldwXSHAPBMBXI9UiDW9SSNfrkde
ANj7bkNcJ1OhHpdR02x/O+TJBfODpkBwN33nDcHh4HMTI2rjN2s9y1d5eDKOjsUy
FPNDDeg5HWV9tP1RYpkwb4byilVn8kXw2t3gUSTPAsy3mnhirOPf+QGXy0sifzJ9
4Qsva4vR/oDoi4Ruyy5TLJGggMD0/MCfWlAhLP1MJ6ReGQ6zB/ZoxT4aDt8TE6d9
VUd9ySKn/705l4fKHvSkaUE+7ZMciK1TBlne53LXDEiVQpfosv0GblVVwIAVy6o5
XbFUcf072/nWGZrJdgXS+HzDPocdLMF5OVTRKlfWDaJu4vINzK7pPhWfVG9/ciOi
J24/1jCDwgOydkEUKAhOO1p4iV+Wq2igEGDRffIpl86ix2lsf1mhtS0wedMII7KE
PhA/OAOznYvoLZRjScHYAH5Lq+w2WR5A2mlcE6yYUGemiHCya/e8P3VDx9RrQXtK
ZGBgFR3yon6J3vMlLkxyH1ZuWjLAvb6QazHcmc3Up/c1j5pcoFZftbmVxLWDTE8K
/wjFQ2lYjCaU9rSz+TncaMUm++0V8c+fnlyeYNJuMY+3Qy0RvTNOqukwESq6BcVZ
m6MLHhOqgxJVaxmJ6t+VAfitzlayG+6b6B9aD+iT1s8+od2Hk+sCAJIZU25pu6ua
ykg974MiSt35xbwfPD1vDgOFY7Tn2H5m1978d5ras8A8Fi7OA5iR314EXyl4Wpv1
sbz0b/BiKF8vxvdwBa4cavXg8bAZKmybFJiXw7hrspEvAk6Rel06y4xaMmqOzQQu
YiI3tBj2RIJ8+vX1ZjqiWN8MXWlGjOQg5OeIp0HKlRANQofZHRfTxr5Q50FCgOvG
8/mZpvmhLdlp4UIpBSQu35L1C5vVPeGP3+H8XYey9IS4L8L7ESssV+RLrq0bhF5E
3EPWvjhL6xf8eNwFg7u0Os8E7ZN4p8cVVeopmlge/KtxIqFSSbYGphedM0UFSigm
kXCxiw6UA+HWTA6byzMzA7XtFluFOpJO0GfFcqP4nDI9+IuUuZm13UtFRUwFiln6
WM2Ix+Rx+Lc0GH5CHktnm43lFFGZEVvNomXIdJKqX5c8Oq1p94kjyfOTSBmGZPWW
oz9MZmAAfPBar9cuLCM4VlRPtW+tQZeLZgSHjcLP6cxtVJ+AbSkKxr4SShcqb1fm
HpUri7QXOunUmfo7gckLPURI85t4HbxGMKDw0jknxe5C6bncHUENKPVNf+B2UtGb
p8A4FQHu0B1gKkjZfza/ezQw9DnwHG6LU28qZPT5GfPOjUfQ6le/PxNRPyDDZRtJ
vQgWVP2/sZD5mFTlOR3vhbkGU/WysimRqcqd1g6jLUvQIIBD+M2zeCoK8ItBu/kq
FDinXwWFO3lbsVIkECWmSxf076bH01TmvRFbw9gZ/2TJfcgrwxkZg4sV6Nm8+Go0
82qqJI9J7J7NfRgZI6kvdktEkFndpbTfWmTKICOxTJLChZtp6H4UFtnOPUOP65y1
h3BZDD4myud80jzeWByvNXphin98aaYnn+j/Cs5P8ptQvYp1YwkB4BzjS+rsvITg
ahabw0Zh0Sx+WonfGv2fSwU940pdsFhOAkm2xcs4/VBvgiofks0acdoCbAxXOxMM
5QMNfFKUtVnP5lvN4ZeEqGL5WsizyipPJXywHb7galN4gyF+Ff4S8+9+tlk8Iuv6
pWjG6EZoNO6mbLcppJmtRseFJlrtUmH3TZPUDvqFYZlwrbEmwYPtULuLL+3sJvXs
Oz70DkrFfWbYGumFR9QWIbwNIYGmpG9IMIjk8AZ1QAd/LgAXeW89OfCufx4lDHJ1
xYdWchwJYDmUWDDvYnhJk0A9WUKr/8EJyzTWjTcroCOCdfKa2jvsY/kbzuUutycc
bV5x/ThtVe2yaQ1ogKc2CgqNcrfaLOuULJBfTn5stSQ5zA4eMUT2nHmDtLSUXtQy
5xGl96TP683XU3PALL0KlNxRafDCWOnW1tzAAynwMgRbIecjCZjiVceVi5RNjs+z
ulhUQmqciMPYsxbO84akVLQ9xvys0/rSQsaZUHbUVuQYmZQqCrXmgY5A4eMbbSPZ
w0xBxg0pKTJsHrC8qBDdkZyQC6tpesqqn5thY5Yob9xb22xOyuVxzsLuxZQ4oB0D
MSxbs7x2p5ey15NM0ikpV67+FZAXQ+rsbeXSK7MgcSD32HXdufpLvu5PVkMS1TkC
KF7/J2UW4ZjeQejs0JSWz2MYM7tp5R96K7fJ0aJtz3pR1RBT4hsdh2Lqeg/ekBe4
mwGvlkECygK/oA2vFqSCgQPSMlXUI6BmrurewWEsspQoqomnERvG2WHvQ334vblq
Svsy1SesNzHZSCgGGCN88v3FRVQ5x7ke9F2OrMjRypWyQYJT5IN3n7eA/ZWuXo+q
yKVyeHHDhHVQXs7lnRBx5gJSpmWjJv8JpADR+0xBZpCOY2e9ouszCAj9YA2+WuCE
5i2RBH7I9pO8f0OCTIEoUNcvtIxIbmvhHQPazy6jUrSo+gd9oHe6Y7GtCNXo3i3r
9UQoOwPA1UQkxIbg5ok3d3rnUonD7I7Em8/Foz5/x7PYuoktFCODlsI/rnXuIAdO
5E9rydV8J52FzXTQsNVgvbRB+6cam4FlG59NSbLR0SkJOnV88bOGiIvEpusiKIqY
FRHcLu+3jhmYLbTH59txrNEbc7XDdzH6ooyXohMaAnwJ4qKOh5FOKv3Lvxz6YpZy
F+QUacotQ4TwlGpFqd2Oi61ZuMGDM7G9z7Xw+APbkDs5qFDd3CdP5ekwKmNOFago
Fq18+XBzp29+eKqXa6+M8oN5tZrGxoFAqlrXibt/uxdp+e8/qYL4cqZAkc+EG7Hu
ODaEfUrNf4BMkAponw8iXM3Yl6ngM4qA/lnB5TEY+Ml/Md9Xniqgcpa1gTgSl6EB
Ig953ljO3Jnu9ovrbo/hrMz95gYPOMA1LiMx14B+xcFFIDB7i2s/TlzzMAyQ/KGH
U7wiFV4UdPXj24MTYoiSpXxgb0vWvkgRqNeIpCMQORa1bySZak49g4Sm9h//iM0S
MoS2CDz2rLrFB7BWLdn2nNbuB/ZtrRGZmQljRNGXMPaGvM9IqNiewXD2a2qLtuJ9
xWncwUnTFy+anvm0g084Z4byh4ZgZD6P1ugBy3aDB1lh8zTGqLKyz1S06vQ5v/EP
beI010ZWM4fHPSGWoTfdofJf8h61YHJUENoMVmQE4RIR/e4PRYEuiUcN3C2gXmSS
RmzyO7ZyoMYJPMtQTg05ETMcq3Yk/cBVhi5Le/M5HvsgTnzxItTNe07naINl6akA
YkwTF/q+uGz2vs/cSrmr/ZIAdZh9MIMyE4YwoW+wm9U4aQM8t5Sf55jszM5I9iyu
bgTTmMNUcxFx6j16KbgCpyyL4JHEyuuOzmfASNQ3jnJAvhhlyM90gjGXW73K2993
nNqnrSsCqhGjiJkZqjogfzv26TNzqe5cdTAy7OmAvMTc/+hS8GfhZgMIkRM/jVml
0dwS0BGeJSO1sGr0UM8Q7/kwiS9OejSOvzJKCOPOzc/SpOuAGQtSTSbDHHxmHv9b
rIf7Y/m4a4DNPGTr0B9V19TGzL+8s0vXR6t5Fc7P/45bBIqtzsdTuVTgb5A88I7Y
t/TwWzgFV3c0xPGThrVSpFE1ZckxJR+mp2C4RjHBrfDzrwTf1JVl9s5i9bD7JRfN
vAjvV20Rst0uRCb2rNvtH8ucLaHCT2OB9mTB23Jgdy8/hDpzJObcJiVbYPxD3IGS
HoHFnd6lir148/qFET208qFkTWD9355Qullj0WKDyvEdblrr+35F1XbDFKAmVY9n
L68lz4RCU+J+ME/oojUivrkQQ6fSuoMD4/cGZ2rxDsMho2y2r4LjDS2b2z60AuM1
fo4qULW+/QEAE4Lf9TZGsrK5SPBmw5+4nXAubh/LBPDFSxU/0tzAabz64KTLA40i
HjXrvS29VHeQOLfjAD2YjIL0nV8mg3IiBIBtkQI/0JSJSjgQLz1OJ8U00PVexqS1
fs0l3naTZW00OiPiwrXz9zSTOX/4SKPB1ipQbvEdTyx3DCdfHNlDcoOLm4Y5D9Tw
HVtdc+JuZyYBsDNkhGcD3UMhE6+r/3n2270qJnmSQZuoIdOzPq/q2sJpLSAOfhcJ
A1av6+on+vVoP2UIdEJsxJPU8Vg10eHI3HZXOnh/eR/1zPnbeY5pd6VBxVlPOv6A
UbfjnJFQusK+ZwyvnCQsFu8/xhKwohDzxbdC9mTNgeDAPXXJm2Jo7HYumZHI5Fqm
LktBWOvH+AnfLtm3rSB7AwEldFMYJJTNxrVkhwn2RaNEU/0oKQgvXh5Y93djy7Xg
crZOwHSfkbsqWtH5HdDxuCyZjHn1WzaML6MVZXlhI5I2pEyLjJX8mm/qM38srqoj
Z6xWm7EHGC6zo25mo2sqV9e9PuVdkpTaYyeWBpFsrIWCleDqFgTGj4UNR6/ulWv4
QGzUWsZMLr/9FBMBqKG5arSpergfyN8x7YWylnOEvleAVvp7IpURI8jmN+Ix77wX
VftR617D9H0VDm6EAhOZn7xWDpGKuU0UkBeu7EVogW7TajXVXwVJx7yogjZHyI/S
LejR3kGzepXToU6QgQ9x8eX667JmSvkiS15ZTRgY+Uqiufhmko+hU6zBNp345zP3
Q/8ILd4SfRL9sdiLqyrn0z4hnQ3g7GJlpeJOf8Jsw3/xIkZrE4oJoJ2RSRxA7GMM
imbixv1BcH7aVVk8rJ+TqxpnJihyeu9zSkBGW+Ahf8E79+xZFBZKzL4TtQqTRK1o
sXlA9w7/3JaDyhJNweOXZSuaMfA51l6b/wPtnGeIfUVLxku/sbBN/gLiOLolC9qr
SRWY6PCwXpTW6La0qXZCA0kyI8tL5JWpW7zj5eEuLn1+CKAxsfvTXQR0VTW1196W
f52DEiSTyui8R/4rQJX+KDxlPJ401TBCwkOq70wQbK/RohNKsxRn1LYtt1OVA1ho
fcJSqIysfcf4cIs8oHTqQrBQ3LQwBcEiX6R0skSxK/nnHDSclCSSlvqcEQdVlRm2
eWz5aoLrv/BFV7y8/8sZuC8nAen8wr6jQkWcQLBbs4TD5NPKZKFgu0PTIDHNZQOv
kSmU5LE9Kw+tjPPBTNHI92JOrNrsTT2CPyMmupI29X85aqh6V7QnZGi258siMvG3
O+PS6AW6yg1Ree9Dx6qENoBw6lN9LGpSanGxINfrYTvrangRt+nD4jcbgpv9IUJC
2JBW4HPC4Dh3gkb3jM0bmxKcCgsa+plq1aff9hcjQnVALSi7N+J51cSvlNfvUBMu
vjbS+wmO/xIqmoBkk8eyFkPdgiHpHuCAF6RwD6pqDIR87oCtXwoFGHPPQswyW4Uj
JtTcotpOZPrgqfdjiTz6kzuc3dufMvA8zrk6BCooeNHYrNiBuNaRrThQWkrP8uQi
+Ykj9CYtD+CCmco7bCyTA+Cca5ljkr8NeBIEKxNHwx5tfwNgqc6b11g3VV63wcBy
4dm9LCak7I4GBAD1aC0/7AF+xAq3CX5T+KlGx7VefaUCWTakd8/WDF3fJgNsqzai
FtPBHvYDPq3f5vn5DQo58bt8ck4o1PcOLoU648FoyBtjZpuuSlYf4yezGn1bDUUe
AkSEZArDuv+p7iyeJPPwm7Hvf9M682e5enWQ0LtUYEtTszLFfbeR6nLv5gCAdt+n
2h+EtP6sbmMjOayBUAskgGjq9jScnayTK0htHvy6w3Q5v92Dug4k9YblHbTUvQV2
XvdcG34no3RkqNsHJnkffIrG3/K3fbH/N1vn/N2rc+/Nl5eOSIWmMProBcGa1poi
c9AJk9ZJm/k2QdqSheGstS1JmDfUlD2OzUeqFkKyboxIP2KQqBH9nJguMkf1Eh1a
W20OywskJicKJDV+huPZKfn1IvNmMr+FgqQ76MPE0fj7sXbGduuYhhN3izE7LeTR
wj48MuPsdftzK5bNYCOSyJaL6II3i+5m6gFWQDIizxNXzCUUOA1LWXJ/hwKuzEw9
ZHsSfpiYyUBa0uDqsVZ3PhYloVBz8EVksnpmq3uY4SfP+Vf9ySBKly0Y2mBgxIvm
75lXaMF6GXYSDq2cY3p9dYSYaSpOI4FdSv9+wQIGyjtUAuAe/SWaonyfBIvU/pMV
TN92797M1KM2wQ/zF5vj/Xmex+2xbIr0pBPz562M0L54vZOazHUMqnJCYPyPuFEX
+6Clmne7WvriJDouR2KOX5oYlrRiRc1apP5t5PJHLWkmfyGfFr93Idr9GzmZLurk
SYEczq/4XCF00pNwu1M6xL6x7V5murKeRTdzxHi4BXRmfK0QBMqjcZWtl4kTttEV
n7Lvo/u8Dzb8Bn6zAqYRE+6LfbTRGVM2yNM5NdwyMAOpJw6RERmoSuPuNYd6Y9kS
HhYMo6fWRwwG8UaxljXGFoAKg0TNlBziSi8bttI5yCOeGrd3h2aracjfS0N6Z5hn
vxkdB/QAOBw+iweTFNrenCRxu9grX7bsOYRSlTJzvlJFPIVcNrXDbdWfC6vIybOC
uRET8+51LUOQ5v0xokANYO/FOQAxAB09yDXk0JlHZ0hsRs7j68cS63RMvGWSk6Es
k4uzho6udrMrUosOnJF6dJrFJbTZ4KolC6etMTG4DSGM+C2+JAJg1q2Z8A2/Pb2c
ZsFlRTuJr7X0451f22BSC8WJJJP4kQhp53t31q7q0Y904ELOZSDCRW2Hrm0xy4f0
wby/XWJt3oz7M54DsVblqCjjZPc+LwcR5cziuZ65qxkiL4YBMpeXeNT5UaEZIedQ
txlBQDx9tNQVybNqI7S+U6x12hFtsBM/lNexqG9PBGsZwz+6lwAxTjFqnI0MQM3a
zgW8W58nIrZElKRr8HE1WOITXMdhOvX9WdERedTWCUCbFHs4Rm/GxtE3uhBhRY6q
Uj8RIbGn33uPvvYf2ytQqtjlKr2db66wC2GCIg+QPQOArcy4P+uz4a+PBWT+eTs7
yybOg1sWCDKECltBPkSsVODvk35G4Y5I3QyDfJ/LDKPvFEYtGr7jbvpwiMSu+s0z
8ct5Q6HTivLtmAB1L3DcL8Kz/d2fGmSsmsr5JKi0Q5xoBjG3l+ZMFtofe3iXxbkw
LTx0xCnqnCIRj49JC9Rx2Bs9GNlu2FEFiwish2HYU9LtCrjnQ+urygR8YaG/xw82
zl67nasm/6J2R68FFvrJQ3uNkJCHXo2MKA1TEhthI6sgoJQWEu+RMltr7+8P9HwR
e2tu0U1kanvhvlHWOsSA3qVIg5jiUASCR7Tito43UrKWNBzUOkr2EUkhVaLQinFu
4OEv+MMZf+X2MJ+1DedCHifzlzrUf/fNeRJ+NQcRfUG6JcME1J0iqhVn9la46fg9
A/AQs5cQILck3lCL3ILlLEF5AQxdqloo75ZfMk2eQfhnqTddflNDP8NVIUvT9lVN
FQn2lzHStxD34sh1gwpuTf4MDJQ0tKGsWLLIkby2ugMw4EsSY5HihcpNAmXlvRYY
y36mtKCo8B+nMLQoyvGGWA8vDn6BNJ0z7TO7QmSUXsP8oql32jxj74U+B6ycWN+7
WTi0Ac8jt7fUA0ue5fcaK6AEfO37wv10ME77SgsUwu2N/NjsaIG7MkilklfpKHb9
7cq1CTATEAduu3nn+xjf29cuTwUt1pHT3zmE8DoY8CUT9ll4o+uUYJqQeYHmid5g
eJp3eEEcfAuDwuNanXuTNNe0ZdftEVB+q06dIyyOo5u++tQwuhUAmIfPQOojQc0b
Mt2deszyHIQUia5kQILYQunIHrUXDdxoOhaVqAYwKkXXoJ3RNjSxtYWta3D5DoM8
3vi0gQw5OofJ45zubv5Swx7KGM9wOkxyG1vYJ4VbbzWaCflFoJTPxIASOd6A13a6
QS9K7vptTUGy2rqn4orXfQesKvRqDHlCJVFVUkybhvaT1nHCwOp8EDWhoQIngUGe
W5sdxJQYMZWlk66V5YQRU3Bqy5gxSVXsiEoW7p4mxaRcOmo8FXBX1hKlJ6bR48P8
Hp5sNj85VYMxCtJh7Q1esVBDH7G8EsEWDGzl4pkgdKb0aAo7QzoLFxICyJLPTC3q
tGE83HKbXmW93bQTqzLENTInG0aqDfQGa+B0pTFh7+wCCLBIDbFdnntISAQFEefI
4QHrgQFoU/79TJWIKQGFDyiJ1VhB4Jl/Mlk2l5UGD5eGR6TsaeNpj3YYUZnc1q8L
Bu6YCu5eDizqKMle+M6HZY/quZswoYch++sER5B8w+0XPByc5lhtK0dJc33bS4PE
GMvIwDKArwyctlK/DQ1sqjHRkiYQvZecYLuNMEjZiv9rbBKdaNYzZgZ9afMoMHXf
NKSVbk5s2F3hr4hu/IpHoaT5P+TAUhXNBYKKpkrOZbJcUCsk49qniLnfNivzVS4H
ZL6LrWklzxmxFRnQWVDqGZ3eewRStxK4D4uF+42gW+Ue0xUJLCNUmitxX0LzLxZr
zczKrxvfFZxqtsomBWeuxS7mKdw5yldwhhO5Dkyi/Jdy2XzAUR2QYGrZ1YbFrwku
/cjRFg6MMXiTQWXeE8y0K4uRV4LHxIWiKz6HrCGFDG22e3AisYB8jrqkwyeI27AB
IOBd6vp3rmjPSA0P7XY7n717luDubNgjy+91bMyGVTzdJNt+H+kuMQ5jBf27rjK+
yGXuE2Vj2F2tntfaEmbh7L7umWG/6arI3W3n0yZxtAQpd8hJzAWqC1/lPok26Udl
ZGFS3mc3cVwoefYtkwMskj4UZ18rtWMD8ru1ik21OC8X/RhrTLwp0MkAwcaRksMJ
Da2QlO/XXrfBeWOtemtktOz2HXhDwRha9Sr6HpjEUbTOy1hDrU5tEuvFY8gt1HZz
LEq6D+Pgqp7DE66s8bkpEXU0AVCwYuqKCzSWboXW8210EliDaJX59hOtmQfdfvul
toSozzyoSkF0imTfhe0jVnNxXlTOexYLcjHAyLzX+EUFjE2BnWAxpIqWeMTh2rAS
O18xiso+sg9mM/u+R1AFg8lee5nLl77r9JtgwYx5JCmG73Dmm3iJ6LgZsCYuYq+f
T+EGELKR+0mXdjBhSx39YNpbAqsOFeAodjZkrM1QHRks6eAAm+/odYNrFUbdMsZy
almac5vu6RTD+tIpENlQ6ZqKFmEjLqt5q+iLLOvxR4hZveecUxxPtmD9tcPjy5i8
ptQuHUV+sFhKWCATHme7yHryb/eg5xYquiopotTJosJcHz/ogE95DF+RFzikeFpx
GS6neBvQ+pkGzeMi6Dsdy88usqtLC2cM8BfwSbYUDM+6bgFpEWY1+UyFG/cuYZdA
qdhfB5adPqL+50W5ckBaH/YovB/QXutcYvzGbnVRN+GBUbKahcCAaeTJCE1qBYjc
6la5hXnMqbl236cROTwRFSWJELWwieYEeODObzVEC7ng+I8T2+TqMiLw2H6QAzR/
ThD9qvLXCrjoCogVw6gwErivwoHmkcXPSnzFmD8WGRiadobxxi5TntUu+fhHO/UK
+I7QpdzPKwpBMkki3kAXZuhf51mapjvhe+5RvraS/agQD1RDswpkI6C1mmNKMKL8
TJW8VR+kZEkbdWdOiENf5o+IwQOvya1mtEWJ/qSFlRytzVu9sgXav6glK+ZmVEzO
FKgDcak1kF9e/5G9WBqfMhm27o1r1cg5FAyF3aM9cgZ9marouC0bDkEA2B/tTFdl
L4j8sHAK1OC1tcrpJKTyY2jiyAERSAiSsbmNpD5VBurDq9lq5DFt52kvJ+Fm+qtP
ZyW03E8otlTbhyxBBG6VIoVsHqfA+N9+KMFPe4LG5JVS6xuksge4mzbPYRuIj2eK
0Efn0nTNnct4VAcGQYH2RAGzm592ec4hAP7GwW8Ya3tqDFod2cXTXdkxNgihsFYp
WpX8lEdB7cETgbzwHpYUnPOwlzcJRywLcBRbjDqtadxgsrfAHeLj9WaQ7jA4/XsU
VVDn54X0oHE2I6uWu2hQQ39CaHTZZKqun9mdHoIYY0COc48Z/AeBNzs27aUaBDC9
Niha6MPw2AQuRYeURwH05vuPNML+lYi0GoTnKRl6UU+oJagttMcTbVqVSJIrGAyG
KF0k8ZOZzkDqhBak0y6nIOTR4dpbdGpmM8WNfRD7Uyhbu+0WtBFB/ov5hLiteRzj
EgZ5uqGxvzVhVK5MdPgty7ZzjFgSmeYeIfUd6Y8U5NDKZn9TJXb+2d2oPr2Kt6N9
yIqgy+aVraDvDMTJiYNX+L7OmwSutwTGjGcTP0nXu9H6a7b7OTSrNXU8XoDhWge1
FKKoNLyboIU3BcbJjCRFfFvMoW48+vZUV6ns+b31xTyIWvJJoKOIZeH+ClAz7t99
gGVzH1bz8OC6rVvHgeTYHE26aOnA+Fa/wnSG2OHdsS4CE5tHtiJHirRuiSfxicb2
gz69sqsBuPC+iPy+hhOYVAK5+CsEpsJsiPE/Dra4esyrgo0vr7F+SXm3bXKwUcqb
Bgsl7fQOkbWH0Uj8ztr9lSm9WaQ8GJSRUeamkfOLEdeSffnwbQcGL3qQbi4KhSPr
SP/TXU810c2cfa9R5R+11hIfoNA6HokuiJur31BIcp9T7TbBZfwptas/ky4eQcsn
ocyezwSDfwIWWnAUMlnEmcA9G7+A/OvCgj2HUFLR3I2ZCITTAHC96a9YWPZQ8bNJ
yvemtC7fr7Fn/dFwVIGQTZRtqVV2Hni7OFrTNx2KrnIiq83l+DLGbUQDkybEm5MA
wi+dggSHFrgGwuhH4F30W15aYK420+MG79mdm4iNmmwRQBpO3D3Fv3t0mJBKTVbO
my/HBiKa5rm3QPWUKlFaoaioRX1T21zIlNPgmwcHsbMluRglXtu8jFmAmMWowbgz
ANpTbPGtzLCXSJyYkg2UGhbHb/FfWTepUvAQ3QEeLEna4+Nkw3iPs8PkYAV0QZtu
BLFRcnPfc6YmGlhmxVfre8kMeYNQ8dJSdgCNAgP/EdRq6A1Dmjbk1tKT0qMJ6M8w
E/+EnSkYTXBqC8LC9POE1YFJJQrHHXnk0zev/yv+xIU/9Nx3uegKd7J6cG8fLOET
P+CK6yEIQkY3V3oa6kEQCpPDwuj9V3QJpcOvrZucGWLSl2pTpPtIonr9dreTDpSx
W1GkUm4yJ0lYqdcPjAopR4JHRJEGtpNr3GiR7751Vfpj7m5OizYxwEHaCEcGlBvP
i5Rzy+8o12iMBSIrF6cU/hzBqt0zT3MSB9vnyGLDpHB/EfY6hiPwYGJF5BZbKm1n
HDMv8x4Kq/Bk3AlkbPiJsy8ThRCvd1CkHywNo4pw7yASzS/c6OE6BOTIBP6sgSsi
WkL2Y5r+n8ttUOhBbGvhZmbYq2D44lX6EHuI+HisBNFAQZE17HDnaZEnxsPa0YgG
6frnKdn+PX10Dtuk7ly55hZd+0z8wD6TTuGfWhHDwZ76QfiRsm7E8T1xp69GuecN
KjRkINrWQzizFsZz3HQZTxz9COHVTMeKSOm+6ab7oVZ/3IO6EQuH7bAIKzWsDOLG
pxeCsh5d14DcBrbW8/JM7Z5eBs1zazsVpNr3M0/VhJN9cKKgkBH7T2zD453CHcpn
Gr4j7pvUQ4X++osyTLy4jxHtYrB5JsoAsOfpOgEPzPtplwtuuL70/evwRkoHGgPC
eoyCKNyZ9KtpXMYKK/pltDySZmVehP6m84DqGDC1d5PUdkXcKqDa/sk3NFd/cYCT
TK5b1MjOBX6WsZBh0a8TmNBncLOn14BxaVI3UxPr3c20PHTUKyTCBbwiPcV2OhX5
2YPS3jlkuzZhj98hKoXEUez1zbLVWKhg9PAjilsaEUwlvl8T31JXwRTq0tTS4q/p
+LK315UCq0VnGKA/k9myyY9ns3TvVMEU/i/4kqYt3vtsC0LKxuj8NXsGcdUwIwdi
JpH03cB6pzEM4EOGJj+OkJzo+5mh+HDuXBfjHD5QkPPslPfKOOAedgwGmb5RQVLd
8KrSzzW8FS/ljWkfRqx5VcoDiBX08AGhs7BlY8jGdbT+Hj+UD1LudZaSaYfAwu9Y
XOX5W/fP7Y9qiocu7nPvtcnUs6CI4wxDkqv3JH4iZzHnxZx7Kaznld6c6Fh5lP2W
bfmQ5hgejynIEdS0MFf8nYnq4q3Y99GqseVT61aC9tOBRJjye8tff9KJ2+Ho2KJc
BazqwnKyKziiEuVBKWADe40EdxTihvjsJLyszNseZKdL1YGBEc+tBu2mFvWxh+j1
TBILb9JaPbjMS5zzPXC0snW+Bx/SexlkELTfB94mp2x/wVvL3Ak4cZME3zAwSLIM
nzk/Bpwu1a7l0KM044ldpBod8zYSkrhoetC7lSqtUI2csavYh7Tg0KfWcEs9ZdJp
Lt9/Tv2zPWjQZlTekQKOYAucDO4DRAlyo1OkkeMEtzxEcPWxRH+w0XmCuYv33BTw
tuEXO+rfO/DU37CCEyI5CSGfLsHAlGUoASN4Q4QsiFfDi9yXDu7sPvIjQ6o4kQbS
BnbOeDlKVD0YJA8RzRkiZ+N5mAehlcx1R4ZoCQVUnyrv2RtWAMWhcxN6gG/Z2ppF
2rE/m+nLezrTxD6wrQlnlVB4YrZLNR+SWzwLWZlZ8qwCWQAf7Ka3HOIOqifs6RAm
Si0Byh5qRGRpEkgnrUEgUQi4q2DHc8iKTeG0PAzOPm7QUJnTaQ+b/ISQzvCIBJCm
xNEZxwVkGEqPkR03Myf0PcozGpMz+ygDWjbRelhqbPak7N+b45h4qZDOyDjBefoL
ZpSHqSlbAdqyVEUau5qjU5I8Vu4EUL7cs8d9MSLacBCEmk5bMG22kRXDBVEIpbvn
xbPq1pSoc+eboDpuiUqNYftQbBZsCalVj3QDRF88JesgjJgPkvytwGXbE3h4FuDE
QrHZdQXWG5gYXeYNmfyhAsEx1SQo+u0w7JIVKyMxTFxTZPpJkmgsF580IyrjiPKV
aWOb5sd273ChWEyLpxdVLYBVY73b0iicXo2UFyrrMELHjeKV49CNfo1CkezEWyz0
F0GuYqtDQXsB0Z49sLHZuvpPN8w9Ky334ccC5c57WiJhC/JIBcZMN0SRc0xKWyIT
8GowQ7Wi6jkxAZoFjexnQk8Hn2pUKRCptAZ1qGuU0G1v8hwulFzRSQIEe7GufDFM
q31mFZP8IkzsljMO3cTcdeMPyILXXy7Su4KY6ws1Mu09QOSW2/6Y3zS8NlbQ2QbA
obXkp2s7o0LiZLXY/rx6RvM4JBKNnO8ql9XFF9lOahUMCrPQBxomWUhOt9brEHIH
Bh3PFGiJcX6EalTbgtQUE4/tk+Nm83ltoK3qHdV5W/xV6gKp/tqCv+1itpXfSTSN
jyPpJT/cCgxL1EPjxWT6gX0CWn6hRQOxblGyZ2HV3NIQSogycLmyktts5bhPJMei
mcRs0HLXJzebwktK6MSUH/Kqb9FGdGvsFcJyOdCtEJQFHtXipbeB47DSr6lmupOw
JUqTN4/CqPPmiZxC2XEINSCBLJyAYCFIFA73dTmCRNxWjKa+QrqjWMGEXuj4QEjV
3rtnlkt/19qUSEzbub/RlA7jmKdE1WRAevCgKJZdK+5pR1Pe1Lrnobcly1r0ra5P
MYCIOfMWxqGQ3isAzYttrPD85Lh7Gv6mefU4ZqZ8HngOrTBXXMbSkyS+U2KXYCZe
aRATkb9hTL8KWXR/6onUhGZZzXOEaEhpwj02zM9EHaJOtWGP3WdPfntXTf4dWVDg
PQgli3lepunvZyWYPKM5S52f6u7o3+eD+Xk1Fn6lr98tT+i0duOAbGcXIp4WLIMa
17hxFWmp/uvZWAKtpknTbiCp3HGvlp+2E4OKPZQiYXE3IeVS/TyeoVXHCLrmb1Va
u0rlp9QTjI+jQtu5HYPHMxPb/bWG+SD1nKvwxivq1cYq6YRF2oA9nIhL4EEn2+5s
l0++sB2aNqg4n/h27Ti3vhGN6GobGwKyQD+mn7R1oWPSHkG1WnHhOf2jE9dslPzu
gdIqfYuPmIe/UACGs0OzaobX7YZmESDVIhf64Yh7sykvkAngLTEs8VwOgqKID1SE
G9EAy5LFYT9eeM7juS6O29cWqwmgRL7ZUvRmf6RldX2W7N7gc6xlyua0VH/sDf2W
vsngBv6NgGvfo6dUWdh82rBoz7L1INeI9WKesFskIhe1lwxgip/x4nuef4jSMFSc
yWXLkA0XSLvILuJCMNtboJfcwYOfYUWc1B/LiPF0248O5DJ+baAgsHjgvrr6i+vz
NYlQVy/fd6eJK2tQ7bWsKtbtFpIakLa0of6x+fkB/K4HafGNxy51uR8Zk9GoP6Ka
NB5c+NIYMd2nERM/Q7CnWoHANiNVGCryYh0N/qb9C2cSSsJv54L5oavOk8UmOrnU
Y9Ebdykyzdej6mRo6Qm90HfdEnRltHv9NX/nLhSyf4lEI2of4lDq1u9+Fb8Vhist
BaRohB93Xfy4Sx6yXbXM4C9sd8VCEM7FUnFdYUmhQfIrfQHsmbxFeYtmwJ8asSmg
y3Eveqh6DBt6DDnSG+mryW10E+rPkC9VygLbLPQOJaj/7/XJGYa88TV4W6E5kKlE
pGd1kPtZ49KLIBSVcGTqZKxRiSfcSLUdxJgNwwIgdPdj1OJV2PQ26U7UAgK51kVX
+R+b9GY0XhLolWKPOY9Yl+5E/U1YFwuQbjioqZiIUHiHFa4lCRfuZq3GKUNKm6Ul
ETGFb9TSSO9wFp8R2zs4nD2RLR/xE6s4uk4fVg0v4dciOZuWyiZdi2J6JwKEoOzd
Twhx6OXZQ+d74jcugoW0oLYEo+kF4nBxzgSFWl00r+d70HzkCtIqroevt5g1hww+
SHQGzeT6UTkQVxQPlpG0no8wO0rD4nq8jC+MTdows+XoBr/MqQO0fOMJwJyQ2BYb
r089n12RGbZ2HWMQ+IwkUt4Ef5iwk2jzHqVhpUQJ7tyUmwU7FvrEsvoh0EIyZ1c3
Uo6W4endTRVvgFZf4TZ88bE7b/eJE1XTGbxSoLgfsvlhXPN4149w3Rd9W8XmGMZ6
GXIXVGcHvLh85DhTDIGue58ryCJnqQoDBYhufhs7+La65fh3La5GPD5AWRmAYEFJ
0Xpk2owmwsOtagsnBaY+dL55Y3ifaMwHSRqOebaMT+5RKi3P0Z7AfGCmLgCsXlkc
c1D0MHNaVkDgouaUBRNijYH4BG9yi0Dd3UKplsCmiiFCDFo2eezr4YnU047jE7CF
uIcIORZsb6PXCugDiCDwJBCCGrhLuZDQj3qH+DqUnlrrStWS/nSNUWC9whk466Mr
Ul1dag9dj64cJnEInGNYITNi9DSQ8/er594J9b5d1MGywWNvDCdzmrUqOKvzP1tj
sa5Gqg1BlrXNswGspoR9w3sgMCvKjGYXsQJEhH+jO89QE8PYNDwS/udlG0XI1Pq2
lh+l/ki02jEWPQnhX6XKCupLGvd/ibwfwvNlq+NoWH0lX/3zgUhUqdJZyxziLLS1
DwmDkIRikXGKLKaDktl8yIZ4ZhQ18A5JGXIPtQ1tHHqnA+D14TpcIqVEw4DrzmSV
A6PVFawJOijwIy9Mwj3qn+pzzqBy8lxV2stAxRNUImLy+urHKJs8gJ1ZgL88AMIx
pZUvBvTW/DcYJOV66F6cuVKSTjmiatybx9FMvfKISXQ7LriDDaRjvic8GOrfsLv6
a4phBXKsebeVoRJwrCf64n9K7guWJJpqYGIo5gm8wAqK2Xcboa4r7waqPj5pUDcu
kFh7q0noEt4KjbSGoxMfuzQ/kMYyp0xoPtOkRNiuQYtCp/Ya/ZaPsap8+vvz+H/f
QSlkl84XplQBMCDYtYFLK43Q72YIPDAX9zYRYLLWFSg4ulVgRpY5SlhWnqwLLEtL
0XJFFR78H0ipqnl/mgO2GzYcfyD1DJQ0tyBjZO8Wx8K0uuQrWArl3OVfcMel3WFj
89n6zFs6/V0HCCB73Gy6QVd5HNnGjIgTnCoXk8DBc7wNaR7450VI+RXPG6bNMH85
sz2CRXBifzW+L1DVll0yCJKXu68qgqzBiKdtUOG0fATiIw07QZ1L7gH1UnBi30eS
v63X4xHgBaiq3SM0WoG7UPCTYoyTIPXuc899eQuUjFcV2mYIPv5FdNYsMEgSmc6X
hqO8F1+UEL8RfT2cKaO0T4BGuqtiKm5P8rWIlmPXRrbWyIVFNzzYfIh88Nyo6qUN
t2x/oh9jnp+hLokNKYlb2nfOqrEnaFw1tENAcvdF5GVUu0joVgmRAcGvDE2FWx4/
/ZEz/JDYEhMUG0sxLIBOOSwvTqbnpdmofz/v/BIzxfJLuQOm9yRBYmSIDFOX4k0s
IvD6PMwfrGJCO5WAeRYpLwIDS/x+V4+8twzGYJiwHCGXiSq/rc8IR/U++PrWDVzD
ZomZwdwjmnGrsWMshv1pltMqtncd/KPxfN/FYwMAq0Xp8jLqMHJmP1ByyHsfk8UF
HhiQrOlwSCH0caDrBIYP/yJiDyNWCUCLLHuXw38P4eM8NKJOHxuqZ8Uz3VvMzpZ/
fmce8mCjUiM6FNZAk15l0p0so86x3wUaJOMprNbBgsKxeVIEaH1ahxklX1BzED5c
hzKE+oB/1K7mvOHnhWwPqcrHm22rvWl8+UnsC9E8S6IUuLxdbVTVOi0hCd3VpJAd
n9Ztwx7zsdxd8IBgFgGGoZJwyFi7NG9VUEkQR45UzjRa7DymXHP6BqQpxK5lrCyu
fJeOWV9GsCXov8EjjtGg3H2cEvaMbocCF0dBjuZ21ZGHTRyAJC1tuWDhYGcFCK/I
V704C8TuFTgs/b5qd12c3stjwvXL9DK4OIRgyNr8eGrJHdFKiw6JwevGniFzbpFe
5+vfpVckx94HesB8tDmkSr89XW6qJb/4akpAsSw9JOz3HPl3bZU4fBZ1l8WQhCRF
CCJf5BP1ssW0TPcWNyT1jAwIJVmBmonUUIEmIviQ3sQ2pmhHAbrrKWKf6TbQGfDF
gkY9Gv8T1yYsMHxHCdmOk9WIexKzD29MfR1qlAQHLc1F4lDGi/78jR95QYth1PgU
29VF5R3cwcgmPUtNf1E9IY/qNrLi85jBoCgZ0m/NZrikGZrrThFJW5yBjLBdaxGh
7KA7zLW6R//SMvqPaT4fo0LPO/rUS/agL3u6hREEC+P0xepW4CcFvEsifS+cEajT
7wVIJZ6QVJsi+8gB47e9Jzn+jfAL1B8M3h3ARAjkdRLMi7n4w0ud/v/ejMNbLh/z
bXUiCTsXT/us07FkhQEdETe5mBL6+mEWSzYM9Sjd5U6j3EwPiT1MB0IjdFseLQ3C
awNXGCqT6JmyUpDb1RasxfihA2fPaYr3SB0Wi1NbgCfKJFOrOnF8O6DDe828y0gp
NyQbMy2qWdA+Z5/43B2oxT5kgebwc1L0zV1+F8a87/wS5h1xyxdHVLW44X2v97Sa
Li4fbQfB8RqQtyD1MSbNdzS3U4e3UgyMuikq3BUNiE6R3x5euEjkI8Ne8qgZi07k
wYznO99M+xh109Jr3hV3qwSSpS+CJkA1bQbdBcm0djCVOkwV8qsJpGG8WJ0nFM7n
0OswygpVbS022TOvQXW84vCB6IQ5ReAu2z5gSEUrOHNvn127jjIxb3b4GUVoSM9Z
Kr5nziufWR3bukSEMmOpXOBck8pc0etKxUNJSpax9wU/ragZUtPvDG7cKJrtiuHz
cWyJCTyNOtHu19FeyoxBw7S1+M7oG6zi0VFvd96HY5qQx7saIt9RQepSr3iSw5rW
CNNw5xRySMDiKXyBtnGkGUL5Mi3/QBmG2desNHpEEm1MCehTrgcT5ZJNvhqexgd2
x9xbCmpNdZDhr1tdhjRya0yUQewQ3nV5S1KLLPIIMCJoXMnQg1QIOp/TQRuj2x68
a9CdDc2CYteyHLUJ+68fHkGsjlQ0GpUu3SrOFIzXWAfoKdLbatx+mrrEXXwt3qVG
Iir/63ksV40dDRQ3LpVvm55DZYQxCeoAnDTZ1KWjdH3ztK+4PKefp6u58+VPvCbh
Y62ixc5Eb7T24jLdNTwzJOv9292rWm3a7i0yxQeO1XD1mKxWCEWrAFS2sbWQLdMW
evrEodDWdGKLQSq5PYeX5z1XUjX2bjJtdIy04YivekL+yQfELylXYVl9hJRdqR3W
xeThIqiSAtXVN6C62ulPpFgzz3d93CSd5lYTwGeOk/jspKQVHwBrJxwUpDfMoLRR
ICDVdJA1eHOZ6NQY8lCpMGjHcv9Kuup8oy2sV3NJa+GXp0qz24UYVFnld3vlCQ/Y
noIZPQNhgd/4mEuyE4pTUrXZEgU+MU5bwGESxI88OzPR5KkwtZtXNpiEAYFw4r+Q
cE+Om0qNsXHD/BRD23BGGKfTVMhbR6l3wq+pzpL28i5+JAFDNXhjZ085OrDC9db7
TRqp6pCtZ4PltG9uG6uYhxlR0KN2rDFgRL7avaY03eG83AsSDDx10KrR0809tAGN
UxFFWSObyrhxTDHZE7Fvmokek9uty4cOcKe2+KZktUwK/sNZGuxLXhqB2wbNLLgO
nwLOPTFLn/w9wTCybcoHyO5MHOb2AjPSXMY3nOmWR+uffIPqPxHOFe4kX5a7IY2y
JI+aiqLU9FMisjyD3SXsJS8ZiQvPtAsx3BRIWyOrfSj5o5YnANBEBLon9FBCbZtR
Me2Xg4kJGK36VfK6BGaJXKKi6zlbtJLI1xHUN+F4D3XRDI9KLK7p++5NeSlnqo/S
wGPCtZukmZUlI6QI7+ebcNAGcHMRQbTzPn/g/rpzL/NSQ8jZN8fczx7tvSIZ7a/z
ltN5ZV2tj9D0oTDRWMnSrpdEwHQkIaGhqeNoPqfqC/qDszSPl8PZa89F/Ax6Opux
WCDXGLyZjhEGYdYzOKZx0Gf4swYbXUrIFt5xMBLXEnTCV+RTHjXSNvZ66/B9ZxYA
pWp2ktouJVDZ6gh4epjOCGZR2nD74WWR+16nGJQHHLDzPcuT2zpGoRQHDwaOnLdw
Z5wYqrkuse47A2KK4zkzVPm0A/pFaq025vz7CrkRfqmvfDLZtlcN1M1TqUEtA+f0
9ffz+EiMfTb479QfwncBz5/rN9GWtUkRmE3t2WXShGaJhygwKA+DLw4m+gr4KsnJ
vr+IC1W+YOwFnHcQtHMZmwrudyjYB526EFCYWISllQ4BfMxiSdWtWVwY63BVg6qP
aBwYj+NYcQeeAKK76IfG26LcB9nZ9gaZeBJ9CBO7plQExVaPstYYJf9tXwRn/SrM
8f+E95qMg237jlwY6KfqxFGPBUGBo/xklhfv8eMEcyu++I64rreRm8ZOPNU/lczv
GCMd6J/Iz6P2QSXYx3w0pXNLRZbSO4KxJEYpxZrfUyCGRsxyjPkcqJrEHQ2Dhe1r
hHgCNmxKAx3ow3nLrPbT767CNe2UF0uf6hxPnuY4NQUOGiw8ewRj72p5EPkfgo0G
V2lgbK5/Qt0o1o89KJqpy7ueheXtWLpvlkdUP8unYNIkmzIXT1TBaU+5vIwJ2zve
A0NzDQ7j+ALankTJcNKamg00IiPnaCbSsyZB8r9d61JWt5zVNFtFoo6WxNVeqa8K
7TNySYZmpWXwFn5UFfPugUrh9V+6rfKXVZcAb3qh7WSyFc4cCSV9JaiVk/oK2VYD
1bI2oYSdDQ7wonmDM9NA8mKX2bPq4WmaItuKdiOdGlLwqhyolCFPZBbS0auNjEG8
EBBPB5YYvVz7e9+SREf/SGLFy4nQoiS4Ae6Uf2QlpOuobYKh+Obgo61ZXYgeNQVq
xS3odUnkqkRUecnO+PY0uSlldTvRcvFieNXN1VMa2DuqQ+j4hq0Sof7Gl+hPFPFv
ZnUFyJU+uRycMGfkrpePncTOKpGUrJq6Ij8xoTz2dKAjGxM/EXWTAFRQS0ufByr8
VTJOHkuxQv4mtCRqe/AToUEgilFc3POojX+pobrxIQucQDUVOw/tmbAsNLLHbYfl
ERAEr7cldNdYMwlvvgB9ClW5U4DS6+AFW6NEsoWFlDlKUd1rt1myeQKgTZ71GbWO
S/BRc3pt/mtgsF8wpN/8dskw5RszRCNgBi5ikX92m3fNoTWR8jxS9dE8I6qPXnHU
+F6Xv6nzcYYu3rxlZZ0sz7DHBLCIDF35hA+ljNGywnuaR667tit/rSgqmN+OKW7E
oqDUvQ/XRbjcLRzh0L3EnKXPw1kNslmPjXynKy7dNZgCokxsqXCSqKH2QSfefkgn
QQzW7+k6wP0SdwDt27RuRTT9IDy6+2erbr8/yTg2jvN1H6qottoRgu+MSrl3OYln
4ivRGoD7xNvXIwPuf7qw3eJbFhHroUlsmE0Pm5R98uGqUB7W+8ZK5BimNtKJSR6o
4g8vtZ+uc5lvKZFkKt/nC+43XYFflr9teiri9xk9iYcAO/PrEkZ9A7t9cDfsJREU
u2ccU3WnqnuJ5JccZFO/fsndhdmiRJrOaH1/SPkm9EdxalXXsT+bf/HhnXF8tpW8
6ylTQpzduAXg0gGjMNvbJ7KffOj+kBkucCfX84eAElI/axgB12pbeXSf+x8Uf2cm
7RnhZQHW3tkiaWv/nenisr+wNS9O/EMQLDLNDm0p9Akpyu6lcLNv23WJBFhPsvuF
o94Z7pVSy3BtooszvZv+QI9J2csHCsJktwBoPiGHQ+gIovFUmeFsQdf7f81HYmIm
mlU6y9omSXk3/Hc4QX08E1YWfFhTN8MY68bdDDSLT78NzcAbqPqZ7b/JKUkuVCHo
hL+MTUzSGjtqztkRzviukFyvSBs0fqP5xiRuTpdD3hGZEGa+YnSK8M9atWmDCWJX
wOEpH4if9pCsj4HgqU9/jmVFB4dOfYaK55seg47hfEsKeCT3I7Vu2I3W0Ut+EJ1o
EQoJfZXPcPEIeRiKDo8RckPbgbTMfkcDQpXArh8c8bxHJsVq/Ro7UIA/TJ/83Wx6
Yhsopuip64XOP7iYhFu5UmN0UDIB3wqtS7wFw3FZrZkv8v/hLsvcjfwSXHCuIE9B
+VRtDjyEute1LD83zOpPT7xabt6jxtFtWdqn9nJh8MxqK06Q0K9IQQ+04FOqdkAj
E/iSXt/btXtVnbi5CH/S0LQhRPUDhhbjOsvjOSO6asfmqV5n56kVtAsiTPnKE3ib
TJRgNAfkSwVlGJFup9Cdj+IsaGjT+Gabz+BWtutsUiEqdjjUjZb5hekIfwEoZlL5
txOzgw7YpdBrSOUYQ7agPGtxDOnkF3TdqhW7HnzSpCi2t+fqVPNm06Nu8xoz0osu
aUNWD2/v61O7MjpFlsCvdYSw51k92jn6X/aVuA1Nl0ilT0eGjahsKlP483DCNAku
u1ANXhc8PaTAHzdFA52JU6ExAsL9iYQQn/rMM26oxh94Tceyo3w6IuNR1dJz1Hgd
1D17PQonm/Tts7wX6SOH75ddB+QCx5qG7/+kAogXvRMKinQLJA846gaSK+9iBsLE
QZqPaQ772sqWfXRse8SVhD0zqUiQOrUQkD6RbkF7qhfwzJh6Vvtd2c43o8b/LRBr
TCuTll0lIfvuaSDK4ebjyXWbtZkOrVJNDfYuVo9wUr/ZoH8C2YaK1EO/XmvYi5je
8ivAvlQTSHf/tYYDoa9EJXmBMC6i5XvP+pp9tmyd4kN59znorpB3ux/NaWGxAfdH
/rqJRxy5sMNG9XyN/e8mB4Y4gX0L3ZGvxfzGmoaZLLRkXNZxP6o4rQC0EStdyrHz
PgKbe1iRI02ArTZ02NO5KOUuBsJaSpJIHs2aLqazFrm/r5QwNICmL1nuQ9R8GUEq
IZNTWtiNVRrjg9U2iGh8JLUv8oj119LGwDsTJw6p/BmgVmGGlf04+Io/TvmE0N+D
8yxP0C3YnqezV+Qv5+9pT13Y3ryjxsM18WeoQEvaIWe/n0cD81feL77ld0KNdrei
eKZwCKEozg841jzODhl0cN/if7VfGKnnbRbBlOONGNkFLACxZoq7sk1xGvOEHpnh
VrbT9jkdtpNBp1m86rJxjRi9AnodqEkqxOUT7UiqEk0zDKpR4I4rILtmT3kvkZ8i
R7Z2VjzhOwLjZms96QDpST9YSva1not/AtFKRouREtaBD/BciaxnDPRFXVZoWhjg
jRSBkAR1TNhkF9SlAIX5eKKt/YqOOByjMPOmlNOA/Zywqvjjo2+gGho74bLTydAC
4LJnGL/pWWYesFZhm/6+exg0+xsFmva+RmieMLDpMWFzD6uQnINydC8SSwAToJs4
TuStuCi4ZDK+gA0k9srUgbtJxGaTFpePzkFoCfk6ro/tg8mPlC5dP1RaJloC6Sqi
7a4zeGa+qroIddeNcm1gHW0zYfyoWme/1MOO7BN4lelPc52sQC6zo5TLfw4rJQGv
glen0/7N/cWaTDwQdyYwvqiiQxS70Q6vg3HAjj+v8S1fW1HELo6MfjuSMLsp0Ckx
DPj8wqwAxJ/j5EjEH+BF08WIB1lwwfw2hKwlhCutP6Bq1ITRZJZIpFsoH6K8PPTA
YALLwQNapKV9Y7TrfqZjP8wtqaRZIejlq9g2h1R1Ohkn+Q9Q/r4CT4i89MnUXezH
MhI38eOAHFRJbFIgucpR2bunDVntK1NZ9wjnBP9YtyRbBKwl9lUstDxFhGnsnQoV
TqsF9ZRAWXA2YidjCGJAADwrkPcf44SBR0otNpdYNnavOAGEx7g/PXbaICl95qVW
1om4UaL6Q6EL/EGfMs7UjqWYGh+lbhsjBQ6KeQNCJvsolPADCnKZ9Vivi/Fc/4/c
x4hvrudqbwvr2HFZ7s7OsAnccDaXwGt7tAPijc2Znc4CjUJ+WXbDhvYkerKQklk/
VJup/QGQQj+n0xScPEIzQbdVslBVyHG8LYyG3/sBrxygr694Cyp49VCH4S6ORk7q
UuXULxambyzLfFi0SoJ9O1Hcf9Tlg4L5pQHogLvKMX0YOns5kQRZkRW3PuOmUunV
8s9JmTsZyyV2oBYIMQyJhcVn8OjO842zS3dooPe2vETPb0ziB4c3J066HnmdjtH5
lXu6vsLr+lkODy73/j3d8IqVaMBQW46Y6C+1qDYjZj6BoDFSbQS1TQHnfJfgDwnN
+YnR6K1mfWmf4Iu+ecd8Ydeb3Sc2PVrR4MrtEmQp58JM3TOhhRZKCC/A21rTNmm8
FcC9QfoIe3NwjjiEMqieIDE7vxPIOAicGNT8v6xWcgh7iCHjLcojeqDGG4GQbTph
tLARAbJAKdIHN+59J9XXm51yHP8Zb8/OXEty7YBHYv4+GhKKzFIbUL3rSNU3G7QG
V2FJpUSmXcgSeJeLIxZ0LddKntDDAW+gNKikvZshQZd6UOOiJJsl+S5rNAHYWGGD
uLW9Ydw2x+Ab9IrGKgfSR7s+KPqmPWBj+mz1VpE5WAaAaR5KPR5DqWBCkcaR8yV+
pb04QSJ67f9pirzDMXvCnHVF7HsDwS88aFOBewUI9hXM7FYN3q0gdx0nEmFKKV8k
TK6ytbMqP+U4BNhX7Oyh8GM6dy5NNghzFGG/uPlGasvVV6vDiLQ5UM4jzV4mx/tZ
doTKri5lRyVYjY54qcRNwivPCSkU6jtw9HERH6jqCjpWzFk2lp6LWc5W3euNlUSH
YnYLeD+81pdvnJsjfkns8vkAJrM8+gWR7QuwcyHfYAy11DrfJbQFvFLc0YlpB3dc
x6n9wOcEYpknsfpenEm+s61xg116yrY9VjzMdgYTdNkBIHwvSZIHHUTSgl0eBI8d
ij4/RgJmzlWOh02GTDD4uwaN+U2kFKRvFN0+trykhUqbG97Hn5+OoxRYQXvFgaBZ
4AY+xzU82J9paCpQr4KSKio0D3xYzaMnKYGH4XZG3nY6Y2yv8bP9GUCgzHeXoCOM
8D/ldc2qTCJ+ccIrokR+30jWEhiU6RUx4Bvvi6ks/4bhqmFymj8y9cA9uYeP4x1j
PADKkNefFWPqrzWFbnwVvCrLEX2Jz9uTWgT2+/psKLnPrHshNF57yPS3ldLC7vot
WAbB3AuMqZeRQjquzUextcFjXzBOe8H9dXg4kM4eqF0KerX9Z3hPTnk+uPZ5T5JD
p7HWkSbVfSqs17tSR36KXmV1StYEFdW/Vr2B/dloCW+CnimkJJWrzYxFbZ3y8ljS
NxGgVzKiTovp+/A3NWocGGrTLyPeN4A0t66hzyoopkxRMvXqko8N0gHGWZgmyYR5
6GUEs/22t4ZyWV4NjICydJ6ZQCdKPjpQDOdHapukcnUEh01T+s6qGq5xUoRtBSJg
rQFPGSaWUR1q3wZF1QckA1bzAqubHwGG4l2OTlcYcjmyoiUPCmYoTxXmAp6XSotR
hOV7CVqj4mygt80NbYB12UfB5hk+9Sfv/Dn2KEs7XuewzxRwQ5W4g7wRquLhY8E5
P/QHfxALhQW6MHxWm1gjW6AG4mv8yHiUlrErbCDcAAbFbOm361mw8m4ucjVTarqV
amSt02ZHnAwfXiXYW4iNFl+gtALjEG+YjIYAice/89D+UWyw2NAa4VyVT/I8Aqag
5K0n3tAgcpaBnWPNjBiAOap/7RXa7mCg9TimEPOAnvFEzdP5QhIK1Z+X1N1zrcWZ
HJMGGA/G1znpZZyMpF5knPgkBkfcD0anP8NxNDf4gtv2upPrj+775HV4xZP82EcN
y2iIPqnm42ALW0DRR+Nuf3r0ju47Sm2QkiURTOIlFuZi0+gBdmSFg4fWYYPR3bkD
mC3QO7EMR+AsjXBJcRFkYWrBy8cTHwTT6DSmPIXaCG9zsZVMNWD+A18xvUMq7kIu
ClRcnD0aUM1Gr80jTtp/TSNQiRPh0JhIZ1FpRHSF4zRn2TjQ78xNDqWXab2nsKk0
XGVKl2wKEj5W90J4Y5+KR58R4sAQ/Sw4dtP7Q3nLOPMRMS4b1upJT4qfTf3wQ9OZ
o8undOA+T0fWG5mqSoi97SWUvYcxTTnURiKkiNvnIYp/0Kpill125Xqe3DevvI/c
pWWHDFgKnP6RmLCcLsgLnaKH5fiWh47EUqB/OD/u5JAi4M9OMeB5EbpzYlVkUqRg
ylYSoHgeCpg8ejhGRu1SnPbAiCDpVWjEOXqtbuWT5hqNTzNcftVNlyhZtzjt2Gx8
kXo98N4Yi3XIESUHfFUAjce11CcQx+9byW939QYtSx0BglN4dZ1Do74Mt3xwGliN
nns30HwCiu81ZUrkuVj8zqegCqvGfFsAbw6B04G884SoBB+U33DaJdy4uqgTuLPw
gSetvB/4775e8gYotWPFz0yhfWnDJGAnBQJDsIcl4BbXyvLxKhHi7+OqI1HkLRR3
k3cXnYMeNJAC4PR8Nl9yG+WdvUIqTuBNmRrP1Bv7OZsKIK0voffGly7HRQVJM8yE
djXtZ2/ET5/HHG4tu0t1NeT6gEU1W8/wO6OinBF5D/MXgeJ9JKb4U8lC6zIYDXE2
ZI990yIuSZ6kUANbUucByzVo/LFkjk4F7iXZgSoNVlw+gfxtltF4V1efhTNXkGKm
SBR9HDDXoPuniI+g2l5egmRmyW/AJWLiXusoljZ+DsS4OyINV4yxaGwhC2/FRsiH
9T1HlJnhlUt+o8QCL507gMB5Tw+fiouerCTDaH7TM9VP4vgQWTGOz0R0psFdBZbw
Lfgi4hFVFV3m0X6+kgQ/A5XZwY5dyWnSnKC+bG5gkx1fXKvhYCe21lPQjMd3z3hP
tbgLqFGUFCmxvRNS1IqvfOUbsdwvS1fShwQVNBn+LUKtmFaZSfH9k9BzvtPC7hZW
fTXeQcGUm51ipKKFWtr8q/x01HspQ2yz6D48ocD0rAPyrC1PSSb6OMPfzFSui+3r
9qxIjLIFSa+qOz5ROav5bTo0dXpvjEA47RbhjL4qe3Ea54JwxszrIXKNhApZxnNH
lG++Bl3XtF2wDJYS5S34VL8yRed5JlH1vrogSMAY/BCJwOPc9pew3gnG5t49iRcY
Bn9/65U4QymlHUWY/l+UgrGDqcdNb/sBTPQweFPOIvZKYjZgeIACS7wXup7a0K5o
WwuyoVfCTnQDOFZGEszE7+c22+WsAsREjDk9S/meGtcJu1YwwZZcNam9c6Ojh9Do
ZQRvEikrFyQAAaswtCBc1SSwE76YR+ZgmKikkDSR5RwUYfDohiMdL5xAQSbuq3Vk
i6HLvszqW9NjD/rEQkw74DVN9OIME/bkUTc337CckrtzYVJcWFxI76yzYrAPvbsw
ZNFldAvp568iHD786LAqVr4SXoT4MR99lEU9FSVZPIoe7AxOg9nq5UWErpCGGgAi
tyM1rnc7JfSFj2WZK0uaetm/PbCfkPgm/f1zyxxSGxfxaLid8uFd/TPO+OB2yfrT
YEWYO7zf8pfrvJqe3B9bbaE9Zg3PPbCZj6NSaVRgXAQN0cPFSt1ZG1C7CsQveX+P
9gDQFSnkro30T4pbwmo+DZUwvTLEkTsGeJU2s4zLnjStpr77dRqX4ddBEgSWcqS9
99LKdMisQ3ed5GWr0K+QICdGNz6ueUhsk4gX6vkRQY1/1dCw/4OKUqSshpk5GXj4
Oi6G9ELvdzugeb5m/DkMUswW8SkKR4HKU/PYnN04hUFF1g7+NFqjVKHhikwsYAag
LWD/kW+UexzoUW9KrK7MME3Jnlj/fi715HI7G/wPzyA3dcitEeRNcHp//2A8BlCE
Ue72rBqjxfwpivJPDWOsyP5psGFsXVw70ZtCRrzDGgj7M1mWQMrEVAFDj0KI2fWv
MJUtQdg22+cVs58cupzi5oMcL/2SaYA1HfU5DZ4rm20a1DHloXZDMi7PERIWzadU
bKN2jurvW1bwYVA20zYDcvZb691D3THOE+OXLpMpSHJcnoviWARIPSirW+Hz+aBm
i2CE82d6gWkJ2l7ZdL7UQKH+VsKSyaiGWwMxbNFt8SRw/JY3jEnpbB5N/W29EDfQ
kl9RsNkMuHadYK7RCh9eDejmUWvitdE6R3fVYepSAqqBLPIbbH118P3/2L8xg7VX
dowJBKXTCj29SgpuFK3WjIXbe93WD3t8A5jFHkVmCpEEG95261uUT0196JheWaXS
jE3Xpf3nnm8IVu/v2OvbEr/aklQFUkyHGMC+IcOZLi/8/I7XIzBKNYOImyu5UJTV
4DnSqH9JxgIJmXndU+52Ei5Ldon7CycpNkkOfs+PuolxLyA8FA8zlU6VH7MwIe8N
VQvb7qzKdSiBDT4e4PMXbnJ5KEbVD0nmA/14z+G9eihL3fK8JJnFw9wi5PSp1q4V
uyYqUQrYNf5Wa9bLtKEq6KbTaqUv1X0oXu9nzOAWwllfGny1SCinSNvbwr5uGv8/
uaUZLPi8EeHu6nu0sj4WJk9k8GRzRJcnu/ibKJzZJAwzL32oy0CsCCdRfFtd550M
G9de6+ko2jAPVd9znQ0l0i6/TqyJsWYXJjCJHPlPYulhKOKiYI787nJq6ZDUeO7b
VwRZ+txZoulgvJ3neUw+qohHQxEN7+KeN0eMkB+Z77I3XFnIFre1HXwty4M36SaF
qjOiKBal+faSgBFQJ5yzNrGY/cmb4rg7Ys85QPcb/OQiXE73bGgIj9JNutNI+8tg
yFJoWsFIFX4nHb+zkiIDYKQbQ99Sz3eeDvTlN96DL8xPiUqWMMeBJHv9C9d/0grb
D6Z6RxlmtQhw/Kir+56Si+WVytbgmDTPOGRDOPeMVOJmcb6GsMGOgYcPUHIy7Wa4
wczz2zTWgfJcu4IMXb8R3v63Hp01HzejGLChim89LS9GhStxe7kkMLZ/0GdBpaGZ
WmXhEIW7Cd6aqeHN4x83JhjEm85raYsSznbbedGhiRgTooZqmQotyEblyJ63bWAR
xz/1mcv94qN+bknmh7Pbm05IUQzlxQ3FyNec/avlogqLOmxjTDI4bYhO5LTMuDhZ
4vmFyUuuLhsPzUaExu9LiYTFWIIZz+6IzLoGphjXgs6p6Sdqx3XWE+e4fDIik5HV
Al5ZE/DRx4Y+u0GXHrDPfS/uecQafZHFuh60cXXP/hKAkheyNQCe+EHiB7wSVe2d
Yd1OJ73ZEghDNPWsWS7ac3tIvMnh4qaaUTbLTVpLzEiqKVN70lpj/iNAXHbGqQ5P
ZUTOcFQlxRKDBN+KMwVJ+24k5rteO1kn5QjIDQuARG1jtMN/cFVjWNBy5/HwsH23
ZtKV/Hcl7GydDFxcmpdW1SWbR/iKFcFkj/6djGEt7coK9AN0lHMKN2dcGYYYJKvk
y6EtlO2g00c7vh8euBaGyvNDGKyuYS5dFuQ0eqvOBnnsHwP8ZvH13O4K7UPg0+mL
sZqU4DxNsNfML/3Xgyvp9DCHl74wDhzUgxVdL2uevpmUMZ2r8X/6jEPvgxKdIuLG
fDC2qpYbJUH5F8+SvczO4t733NIva1ouEZgJyI4ng74fZFFLnsG4E2SRKIqPHpmZ
NPKCEEHi/OVwo4vZi5+aLrrMC83IfoJzKfySMh14BuGUq/Pmeuz0NnLjfCs2k1eg
Tu84pnZRqxAII1pnx3UFcgEdb42HS666gy2pPXO/Yv0UK8d7KjtuNXuP+NNQBeLv
cNjGuPPrlTDFEifyH4AFn5IkHAY8EguY9iRvRLocXg1rW8p933SYA+lhW4ylsXsy
5/z4nmVGu4ipI/4whyxUuYJnNJObVCOD8LgRSVBVvBwqWox81ShI+dtNS9RnlT8s
gg5FoBVUnK31njs3BoGHY0c6gcDububrATecC05s4c8pECgIwmWKomFqM7K6uUI9
ccBD7U24J4+e7VCN4/T9RShbH2jzDZQPjDdzZ9Bstp4T7Hvfyq4eLWtd/y+9wlpc
oTVzDAMIU7+NwUf1thkQ0vRebiawM8b6bATSfcvNAfgl4fVLu4+KFm/3cNL5RoKL
oj8Y+bGUj1gMZrZXWttz+fpzSZwm1R7J0NCxf4rEEsPHa9NGqmGWU73UmTWe68WI
8sWO7CaKOIBItR0BLDB9ZuqPSo/VKNHs5hn6tqrheipt0/+Qb25jZMkOcsT7dr9K
gj7p8aoLxiK9fYhy2nLbS4I/8qBekpG+AdxBmukJxQswWExEXkymOo5IytMONuvW
Sr0/ZcvcBMhIl+aN7eNISh5G59jyg9p5UOce5Hn3T3yEW60gLmcvHoN4+WgW2GcP
H+L+vE1HVDk/K/IFz2kmMBGs2XETRVsDL4/EqrkQ77/jy53z8wDTVkxH5RiKvR/g
6QJurbp4MCIZ8gUxcv1IJGo2igtif89wpNBXWpsLkOtf+BJOx+d25Cv+/A6IlLYo
1kZR1fJ+tShvsqUT1w1lHuNpSPkCEN32ckrVNIINlOerJqSlKtxrAN2kznQ2bJ+4
bXdcGQFhIkeYlz9hrp3PC8FX6k6dLOpIjL99qCEuq6e5xMx+7hbusils8l5HCunz
Qgy/TtmMuyI/Lo5CtAdUSJU8yar/vSX7MnmATnfSFOOyGgBT93syDkqvAQMM0oy+
y5JrY9sQYz70hSokdmoFWC89UFpU8VAOVfVbQZ/eWZq2qS1iPI28uwlfMPczKqFf
zQrRJrt+u1RapfrIQrwZkNLzq6wGXaqa/f2cJ52WhO5AL+bDt0ecS0/ozpbbgf1Z
DQgbmynkRpDO+KhKLWG2t0PPD7UpeWkrzOEuLL6bMO6lgpPcNIf41bkUTYLTpaWL
qDvpgfRatbCBwA2ii0OWTbspong3pFacCCmjjhBtorTLMmN3K1K7Xc0ah+9+GPl8
2VWvBvR4q064A+F6qzVtDAS7LeNfKwA5aTn7U9vrwikUT7S9ZF9ZIeDcwlenTDIC
VvjWz8IT0gw2y2wsOHQWp8xYiejpf+5MnK+jsHbEe4Sb0TbBJbrSUVyG2N3EaWX+
1fgdReYjD7EwB8Z6n/Cfdqt5O4imJyQ6WBbeqacBoNuPOc4I+BMbU5knmg0EQA9U
638L7npBRD9YFEEhr93Z2f/+971EfBHsbsDPKJhGYyte/AX3yoHJCrQfwggCBV6n
PkmxtT3P/G4ph6LGSAXe8XgQeUm0fzln/qYryD7ZonNK8Hh/wSO9SOGmPI+SJja6
jYN8P7iVaLlEhp1CPe9qENLkFqbQcvSVL1r/8fMwEwxx4uSxO9mxzHq9uO6AaE4y
u/KG+KN+11S5iU1fr5yriarJjTY6obj3rUjqhriuhsiBtoTOpeayVpk0LqPpfYsN
ZNBiVdahxbMQKO94XUG0QKW8KPGu5l74IHt983T4iSuP3CWyQaVLEBIVMMuahr2d
wNYaEWcGcRzB9NV9ugN70H1tKKqYpXZnnrQaKyvboj7nD80rSV55OPuBNzqTrBiy
ajYtKrnuyX4aVIHvCV0Ps0VMNLETzK8l+gz/Ru5XzMuxKCTrwbkpkaFlMm2zc2t7
AL0JkJ4LK88GO0Cixw/tCIvurqjmtYn0lFmn8kuQnKt62K+g0n4qtIUr1H2rBfjZ
evRDdbSjXntS7mn5l6mQ+Wiy8KaAzsinQr47w1QzdjkF6gm5p9ZZDqyBckBeeeCK
dSf0eoWrb8L2fVs+2NVArqxvQQw7Zbld7Hhv589h7ICjGlnGKFFQabbjX0Nue6CX
I+YrnSrL6k/nAx7clzsxoREiMA3ttLs8XNu/r/QZitKl+8q/4Qlq+lLfazaC4tiK
8eFKDDbyTRud9qiq5TDVXrQTlNT+/czWdQ1oMMnE7Iv8Tmw2ei12lQYzRqunO5rB
j0apuGNRDRejDvaTXBeSMaDNH9bl9HqD+HSaltRqZ4TW4h555E8ieUCcHzZFwbdq
t0h0tZyNEF1POG2dpLdRDd0nlksoFJJQwYVCGUrsZzZfMuMhYl46t8voJAAmMn1E
YL4BZR8unQn4Y73VFyGvZ/LlHmPB6/KNCn53nRTxUrv8WqVddvBxYHuMP2ACXR1m
LnXbRtFUm76lN8L0XMEaAIGgbdEgMBW2m0t/8g+rVBVEeTrRdjK5nzjRAY96YA66
IzyIiao/vgMmYwmeUe/Oo+RWnRLOMDhdzBcG7f4Jgww1sVBpVEF0/oZ6pOCsh6st
1n0M7F4kBhj2hn3Z2XtwCKjGygMuom7ztBSM5OAvWU/FhpLo8R1kQ+TcfNg2+hlY
PKeyQx//mP5z2kgQPHhsPYW2dbJtK7KXn5V7O3tcwK+UBI0XyCcf4wh8JAyNHyvb
6O5AphA/Ua3ZlAmYKGDNFISFAWgrVyA0M4pX4wYnjDbRhgx+x3OZ2qqs0Ck6lz5c
XZOOuzGMmhchIrmU19yDuSuARSkbhtHtThlY/wZAmDQRTZGU/Kprx6m+Lcn6HBE+
fMUsFAhvO9o2N0FKPzFIvKsa20sr9SH5gWHcNOZY4xNBp2nIBEiJ3auHdY84lPhn
fP2RbgCQStSiMZQiqmgLMc3+vvAVgmT7XNV3DMFIo/tRK/QoQQPDuzJ5YZLBoQEf
WkTeT4SuNvtH6nuchw/KWZN2KZ8cQGK8JvBhGpQ6Xji6hXNFvFr4RwtD0fUJxSIq
6Ec9iVg0ozM/u440Z7hqsHLtinrMxIF62kHya2YOoOe/Qa6snrjFpzdtXJnl5z3N
Ab53GoSwKGw7afGW6w9JMBPl04763HTa1zZxNdl82/8fvDrxdv4DALX6vB+Z7JFe
9qXPJkDAI/riWtLgZkWzedPHYULroojtbccduD/bVBNlztdrenVNDztKfODmBtJB
6mH0YACdlmkh1gCDJr+cuSYL4G2dMV3q9mdHf0zLv4o77MCfAliRQQHM/siO0NaW
JwmvzJDxUz8CYSF3rKrnstCvYcIWYQP8/riZelcruSEx2Djtyii2590uCw3SXMb5
X+qgmtgMl3w5sOW+JTM+EGuLJUrrkZTZwiP55WZlEoDI2wjVKqvhvXxXnRRq6DcR
2EGSaH3Zjl2irb8sj2I2nIE9PV2FBqdMQkcwzCnCEAQRqPw57+QWuZTB8ewBgI5P
PqrJdPlkcH9NSeMmUswLv5e98OK70oTkBPWrflKdBA6gfl7LhgzI9m/SgMZ5xvRR
RAY6HZKwsc6oF2ZxN0Ri0YxL9iqHWOLROo7JgZfluvU/p7+ohet8YU/RU01ibOZT
v+ZGfKo9CXu9roAT0USBbEjFs0V45hW90o2eOydVN+66k0U9Ft0sr2BPVvBM0UlK
RLS1h2GcPeJi9DQ67x8PdscZYvKe0lcNgt65zB2hfGw3FG3EVbTxwUWW3EpHPEVc
2iEKbcWhZkZge8lpBvTFYJEnXM0IWv4sQrj236QRgTQ+RX0aDfxguo4wpFbNPc0N
d9Am/PkccdpY6hefs4YLewuI2gKM+O3Bm17AcuWw+96skurM+df+aNZKS6FIExGs
CtIUKuiF9lFn5TTTJXUyPF4jR+4O9IG/Imgy7WnGseeoki2MUDUiS2RNplneN1tx
NjiQeVXlWp8+6B92P+D93v/0k82uv7VlHvgcGNYkwHZMcxyx7W0xpD94qL/bYi5z
zUpP4bZ9tyThnD4BA5QNzDmYTHMAKa+3I4IRHScFqQVua7hbNc8NLIToptpufpl+
z1zIenGYURj6em2cqF7NYH84vDq5kBkb11fNTTZ1u/2vDQRr6Zj0VFKjlwwRB7Az
RB4MHpauKwAoYVFSFFXg33nKSgsmdpcu0Tl9kXXvbfPOkUWMrnkFubRureAWpYCm
vOtYdqiid7DaPm9Wzx3AIawboujn/LF1C36cZFoPKKAAYiGXyVfshj+zSd+cAWdQ
yrRQGTFDligOZC7Ek4dAKxf8CPl+c95GMIKy81BO5jOyCJE/uQXTFWgc3hsZVqQM
XrGcsw+4UsYBo39e3Xl82T9nCMfOrNgP7gTOqjsX4Lgks5Qn/uKSsrbuJGwaGZ2m
q537FlI3BdlKjdW9N9fIAbGoH4aczm/fFVcCo6ieiAU+WenWs7kRai+WpnrbFJmh
NvAB1BEYTMvQ5RInIOBRl6HKzdowetGi4vQI0rEf6FnCFNKcgiDQSEOs7/7dMHLX
ZeEh45VZROjbXJkCVicA59WvHH4chXyyDhME5cuyY0mUtZicgWEPbwSyymAn10Op
nK7WRHbMv3icBLdTOm8QwGXIkbWKjEwg/h3GLS9mvzaEcBEMgD194JL9VLd5i3wK
dkb0OZ17y5VIRa/YBfflEMhjcVk88vrG1l9i9wzW/YIkmnLbisWr+dQ8YfRRCnt2
0fcKCyGOnyqUaFaYBFGKMBroZvPqUdfQ223L81yMcHLvg0IOrjlxtYEPvdLg8U4a
ieMQt8CKWdCiY+gOjp8xcw+mZNbvJ3Ijj/AvUXut1mbdkiwCREurKO95buov0CPL
XzphLBkoTq5ww3Vx4nweORdCeM7NVwjDg//BmHQ5WgdLU0kfrZA0LUp+PLcQpAfw
XkvSdOV5XW3wZnsP03ftnaz2jKirCIgkubYxIz/10I5GKOnE4+gHrRaQByt0yc1T
zhU4x/TucWTPRNiyyg4HY11TLy20WR9aE/IHmFm32OupW0FVuqw9TNt5mZLrcp2y
fN3axOgmG4Y5veQ7NnM5mGwLFJUKq+j86398FXyGgiqHv9wkeueFaYcDSwf0KjeX
QP4GtRfl2cZ9wAYEEcMZrg4cod2Gxft47XMxsg51Izvg+9FiQ1VxLq9bAnSGfE4g
liiLEI1a7bODmuU/IzioCVOGKauA8ezCVGBj44yD19AvRAfbUUrnmbM9Q6udPvu5
8pYnYu5f3sjd5ZwrrURXXaf5McYTaqHU19SJI7BFwXmuf5s6QtaY0UjxPt1CeWiq
m8Fy1KY/HqYtqFV4PZeHkV9TM8bT9pLjX46cQi7dhXGQG+QGTPqyaHge44ou3UN2
qDe3o8FVstQWspbhpZiAz6dDaSgnmFY962rjbEPgy9U7M55B1aapKPBzQ7ALK98a
clYFk+ij6jkjIJSmlsefBaEEKJXgWWQudOIq4L8bBMLRZv1722pAP0EnD83/YI6K
OVvDPtbfC2GbGojBmCGmz5HIIDf2BNbPdTkxA3f7DUXLIYWHp3knaNaXN4uF0PB+
PFIBxJSyLLEKSbIapPXIYSO0oJnLxEaEqAfsv+rZS3DY1SspOAVGsPUq8uDvnkYH
hPQ7GvHkRi5l5qVMWL9laQJqvrzxJv1wa89RngOjt9lkfacHLZmmLnAUSSs5se1g
Bmt4CUkmCEXtzA6uyLABuT3+f5t8p/68RUjWAtl+9arhp6a7myO5ABHcEB8jmWO4
OIfgjc8pMcu4+IE90lShu58+QVnjhrktFdYS+YVcDm+FQx0y4KfkyiswZb4/2g6p
KaCmYlrOcwYwqCVblNStfwaRzmJebVqObRG3DFknHY0a3HOgHNZSrZ08WPUUinxs
yd6pHtMSMqV3CRkgXgx679CymUsHNp0CvTiW7KXWTpam0DM+dcrxS9V/jsy2at1C
/0nzxTmJhNTa9axX2U17tHLug9qOhQGsZmqJBDN89S/ulk6vUfX+RtPk0fG3yU8C
geUfgNCCn4x3yCOYRhB+6+i7wI5W9sLXSkL/GVGHWzLkDCo4zzsXoGQX72qLZykU
QzwMVOhLrPxqbRPb2RfUbIKzts+yZ98xv6vorpWEycO+ljVGrcaYRfHZfkjb244T
toNBeHTW8ijNqQPl0yZzpSuTksJ7cl5yfF4F7IpHLNLA3C0bEbheG0/xutO56LK6
EKBR+Whygb8tgoRCBUDMVd26jK8h8dXLiLg6o3WwMIG8mDBN0lfF5vqmbyRoUbwG
+gCN9cL0YHApVO4V/RNJebSKPxX504bGaizexzoVXH92U6vVZ0vZxuSf2495oF4U
wa9Vc7ijIgFvjQva8m8pz+ASJoN2evsXuoN4aiZ7Sl2ae6gNwm+wsUhl8NsWW9BZ
XFPxNjVfMvlPIzyy+0L/eIvZpVigpWDMT1dG0s71zjUtzCuVihZr56zddNzbfOqW
QdWo8ac9/a/ebB8w/PWYPjwDnQiv0ktgnwtcAuCzh7d8EM0kJzHTU3F/Ui/0Y6NE
cIqh17aRjfAAPIijoVlCwuyvQBTAKej1j9zQoKl2E8VheiIlvwGgaZerUOYvR6Gc
+4G1FPQxvmNJf1+bgeTXI223V9PNDWeK3qE9a+TFwFtufduflNzCLwtJ+L6aGKen
cM0QFjuMj/FQKSdPksVKOObITmP436tTQmFVSnGhA1+KlCQ6gVxoZZbnlmpehTFH
tWj6UVJkvVq5/WV5zi6gwQQH/sv32gWx+SMu6mXPMVxF+Pn4GaTAM2W2t5ov4pVT
0GdsjO5rYqoigZzJFH98/b0l7NvDbZaVGkeWxDhnhHNFfMZ/N7T7jR5FMqo0+UfY
5xhUO3u8zwbP3Y+FWw3hqE51HoFJULck05T45uMQzgJu0KP5D3LFjZdN4lWc53W/
GM4NoQU5I+yCRN6dnW1KRJS87gbpyJJY6hiSGrSb4IUdGQYSVdulrVcJb/ZoFIk0
qgv3qPhQmrweeYx3ePXM25QhaSZq8R3doziQLzFmr2JMOuA4Dny/dMyXnv+C5FJ5
xK9rWGc/xNnSWZVf7cZdqmXfUFmMCmN21225KhPTapds8Y8kqCA+DCZNR/jP+5/s
lZYxqQdE2TKd2lapkgTxl3mYyH7pk9IF4n9bOIrmoVW4xWiX8UqZbOkRevFFJAdY
gwAzV3BkGndATnp/LgUqoMUtNcT2HG6TiBPQh0fhZ4ZNvRKn5ugkxkt8v9oM5THt
T9Uq/Q/crUR71V0/Zz92LwdP7k3oYoToDsInY2Wm8hIfdErJc/1r2WSH2AY6omen
rattLvRyKJvTR8Rpxc55klNPf/ApBkoXTJGn+zjAo5qjIL1JtRaeODke/ZX8Mf46
40lZXW6166jM6HeVX4LlT6ZHl9gblYeZ3hfEwEiH78uBsEiG4D6Bxcp8JRqyxeaz
6FAHvZPtwgBJUhxfhEY+AueAYp+cICoK23IK1K+QXv/RfnUdA+upZybpdNrfppO9
HrFzySywCL2SCgNLTdUgXI8i1FHXixihyk8Nb/+8vChw3QgNK34ofkcaGkIvQ3sy
nhQzesSUjsgMYlnO4Fg0aU1EQeYZF7UYOu1+CzqLjQQ92/j43J75CJTrRA+YQ0tA
jyuOFIBniryPnrJGxP92RkIftHYyKYCQKMS9H2XoxixV1QoOLwRaRzKHxSbfNRfD
Biun1RwT9/cyNUNR8+KbiwideXjc9T91bW5s2ZqNMAoSl25ZR/0tuQ4Oh8g25TwY
T9pVnWCxCgqgLB0hU3gmtAwHYtuGcEvhGIJNM8A9LEdsyv0GKyck75b8WVolSxmZ
e/b2SgR88JHwayXY5pGyhA2KNfuPClPNIvBhGYUy9FZGXlJkorLH9JpMsdsAF2l9
igQWFSHwu6c23wWORx0wIXrPxcFR6PAxQBlH+DrtDCGfn0KJIzVO8tOJ5hU9NNId
Au3ZMLVNjEUF0mHVq259ZuNFuyRA/Ox1nVcMvG8CHZGAW6D8I9OdC8jDtIZ5O7Ia
aT8h7K04ieV44vMmnlK4vJxODZkEJ8dPRAqC4OmCKPKCQ2fmS6VhpW18D6+gRb1l
aBEKbVVKDgr5WUXDGiwHcWK1D833eHefPgEhwTTbI13iGLmICsOC+dvnm8UcI7GY
v/NQyqoRD49SSxev7lUie8VpJJNIwQ8rmOvD4sdO5qDypVdTtGVgoFz5Hin3avKa
f0IUvgoxCFzBrosFwX68+YveSuBCn5R5YNbPZQZEGXElcn6S0prM58bgPPO2o01f
eChH3aXma4rOYm2QoEBbaiD85KU5W/q+j1O1zf/zoVKSDAbk4QR8dFlz6nHIFJos
AcU+eUKRLAtD7MExGH47jicg5qCvloNEv+wF0FK0L5rDqCsZfi+OUxnCoEoSBkuT
jNwcKEFAMiBjIjXMDEI7E6RP/kQpqjPTb6Y/RUkvGbYGYwrWqsAxfAxdEdr5Q0pj
ckER34dnxzXq68SEY5MEq5ymEtgRogl1w2eTPxG+IpI/xCmMmAqsGZyesswQhCf1
0VihMe+Hnm7puSQYaZLIALN8F3ROahqJ/6p1v86WA+2Zr/fSa/dADbtFBDkDXEYv
hH7zukqFn/8LIifHpao3/s6VBULYb1nR6c2FbIydpO6anWURow/EpGhy/YMTOuLl
zVQyam8O7R3VGrq2PR7D0D8PYrONV0WColbO1f4R30JXnJETvsb5xiBCI4cRSax8
BboIvMT4xp9Mw6O+0OSGkM8OfyISjipNBpRqu1safwW1NrFkxdCw7l8dW8dLUapJ
OcAuhIHxqJUMK5xXm5Kwn8lpdXX0l6kiyQfCCQTx3r5UZHQRSGs+lBdH4rkidUhi
ZwzO3P9n5DdTr9UVQdpBzXPPxyB+a1lbFcnjonBCpF5MVCuvqNZVc37sDz+qxmVt
KAEJTLI5xHJcCK9lU8XTgk2sT3oR8s8zugfUQiek+uCGjL1TOM+i3tLKSsnFNnR4
5Tkud/4dH+Wx6/4Q+Mi3MwyWFzZtu3brZ6oj2TJrGTjoZAv4sCPXbZ4bPehhP/0t
d1BLd2PXYFkXHiq9/9D17yEzAEmGIYiWYECvEwo+8paqmlGenswuP7IfL7M2CHmb
i3+4tpkxw+JPoUzIMJYse9nH07XhPXW0EqlkQAGcd8PFKG4qnw9sy165j8elxfOQ
NmD7s0La5+9t6YUUgkCRrUCPd8C5rn/hDUsS4hk4fQcT6F7M1GpL0ucQ72IviutT
GZPadKPYtlqyPhEjJ2lGqojlBmzN2aavv0eikjGMUKSkt5piIflD3PwPHE6/S9Zc
yl5M+5gG21QqYU/QycjroB9X7N8lVY8NoQCSUIs3tEqSvJ397kHfBu5f75Fz7+AO
fgK/Lt/UhVFl+GuxN1blr/SjJ0M6S7hogd/RAqnyC8dtXOxsAEi0MLEoIpKfmajb
0Cz9c796KCzTS/7VFDpVrYLN7jKSbRrtiEaYlkLZo2u67B5DJMlq9itHTB9gHcZ4
RoCVo/eu4bTkGsJhjR4O4yqrhNjDCkumLGpjd2xYXt45sJVwsZzGRteLT6IXJaHm
EWPOKrIXI7qgJlk3lSIQPGivF3aThHn9eD7MTmclZp+RS/6TycYk7ElLrXZL6/8S
aE6YEOIxIseVM50MkTwS4GoYBlJ3MWmi/NnBU9DZJXGNZ5kVW6DXda9smfEEmGdd
hTPuZmef+xzUbE6c87FLQYC2xLCCfubZrg7zHcOEBNAlipginCks3yspArP5yLzS
PGBZOociOB9HDKF2yn3loDim3D7Vgk6mGd/yerFy5jFodzJzzKokEf2b4pSk+hY3
ZeKwbCx+IldhYJJINzvXdJN+GO3e0iv5ZFf5cCzk7hw/hm/SocUeu+al1YnfDws5
j7sQAzMHJE3mJQEXlQv/k1YUs31l9yD7uoO9RB0Y2DFZbzxAG8e3NNI5CDCxE2t2
8AMCp/+9na5rXTruvzvCq0PSSIJTKF0s/B+3iDlntvsP79l6UBwxOxT+GtRTe0ww
XzKt6+LaSsl9IQam3pqBEYvS6BlIYRj9gRIfdRVwC0L5d0kOrnFHc7ybTZgMZs0+
c3eCdO+9UzzHW64eU+BpcgfLbIWp99RFwHPMKzGL5uo/MfzjsOUBbvR/Y2vb8uXO
u8jpKQWMid3g4hWezyRh3OooW6mZ/ZGC6pusX6XDgUZpXI8dXplKRivnrPrAw7Ol
nY2wdgmYr4kw/ug9KwveBUcCh6ZFy2gR3hL3WOIait2ACS6FQq+PRZCsjBJa89Th
S9lGs0pRRwoqkvKgAumlVWGxqVyElc9Tji6bDlSBJcU3BSoYPs9VI2NEQx9ufA5d
U1pH/gyob6AUP5vl9A60ymji2pnWztNF04TED9CFFSQTva4Dj9712AgR6lBo3kq0
m6E2Jq0zRYtk4hlGElFi5e5VXDI9Oi2NSA10ky/pyTm3+IpOPyLNugwgINd7agFW
bLxvAajCvzxlylEskYFEgz5oB8rqR/2NCn1Bu/3yIc8hJFAEQgv7yM0ek3ZPOFRZ
vNBIFjAT9lzQE8gVtbS6hs0AP++9Q/Z1sEZmz2eMSDEsoyYT3nn/bDs/lqJNBnEV
k9N+RDvanhnTd3WpsWCQ0/v4AoQXQ2up0iV5I9lPYhyX6XY/YcIzyAP2RErt9Wbm
fP1GlFrbLsvJyYbjoa6f4OJgKIwymr5lu1N91L+12O4pYbPPZ5nx+EHrP5LwaGUD
fRMWGVVeJ34o5v2BtecPa4lcNDuoeoG1M03i1STmxls7xnFy6rIRtV2/RByLtaOG
KjUMnmCMtnWbv1vB2BBT0egvgc+DWbY2/wK30P6wVEGd8eRf/UNTeb780I2XK1Yk
LKeY1uOYmPpZ11RsVTzBkNXNTiC5ILrREw/DtFtAQfoq9KIuQZxSbx67OCUb4GJD
X5IRwbtaXiboXIOcRtNJcOFfM4kOZju4zFVEJpulCiCqMSOuDt/V0IA6NQMtS5as
f4mjj0bXPZ+K+XmUJMHoB4ImCXp/OCPkEpKV1diOPt2ZRcqqxqinDHR4QhcwIq5h
Ugz+4QKz/eNuxgpRS1gvDcbl4rN50PB6kxeC3S/nZxCzjih+PAFzhVsYtizHBXFV
W2oWma+60ejJSvYnIY8Ti80WixtRKw9QHaA5DGPJR5InFksqyun2yVCHEckq1Jvn
KrMXZYZdLvnWv6ZoQp4gE560sjmdbE2pSB3Br4r00YCRB9k95wEBJwSu71R707Gr
43H4yAoSd4tQVcx+TlB1hL+thnngYunHKVgoNVc1R58AV3x5kEpiByswmOCVUEj6
w+FqV9ZEQ49wG6DCFWdynwBVgiVP1qessnI4iGHbkIK6Z4B9SX6OJQNOLxfNQ7BG
J3LuVuHqOVjdrOqYl99I5ZW8QXoHi3FsSDevEZ8e30d3s8Y/Kz9LE5TacyliM2jd
A4hLj4Q5qvSemhnz6kBGNM57fpQkGh1K1A8Hjkheg67ROOEIOqsdFJVbkIXnsm9o
aiYe7m6q1JGpZKvD6pVJWsH9d6QIgYsyutgOxmCdvZchjYfmWPw3PjF7HRmDG3h8
8YiRv7LT806S7odPjQy2a1to7bJ3q1HX4be2z7R4qwNd+ODVs/bR5vVenxV89AZV
Pw6ywpNIpr6I+XzHnbtTq0aSSsJHPA08pFnSpkzaflZAKqRHOt5fvAyff/9tnKMv
z3a39NMmR9rIaG93ZJXhDfm21sou4g+yhF+3BpsXoay0acuiChHxO9QXNLiq1aHG
EADKOL9dEj2k0CN1gUi5FGaR417O62lo+7lgDecaRJEhNZZgA3aYkbikzHf6TzZE
CHEN3DHYXLCcsGf3O6goBmMNiiR57uMX0Zrzn1kmuq1QhJSQPQryqTV7/tR01oUl
73M8wBzmN97XJMfKbHA6gI8lqu3QfEnjGL+1ImjciVHh/lW77FtGyPDOLEvldt8c
Gww/hfwWSSQV3n5LBf8CTI8tLbncxdJttujTmdGusTZsxKaU+MbL8xdDzuL0vlp6
j46vMB79ABJgH0bzZhQA2JX59kXQOS0+xY98v++opyf/f15TAIcgl/5gtqoCgu2y
Dq1j1Uzu5wgfmU9dYAhqED8+ub9vhrpSTLrsAB13ldgdjLSzsTWpBbvKzu1jhp/W
tDJXyIRAu9EQWQjada7ui+6vx7Ke6KTedYYFFqahW1BMQB1VeOcCjNnWrxv4KL4f
KWy7DDh4/E+XvhRxAoTXI+oNhUTxfo9HJ28OKwTNcRiwfR4qfUiU5f4D8ThuLTZs
KUxBQ089Ngqm4D3Ayg3UnHdu9bfHx5dNTSpdMmyrpM7sWSnKfKcMWRcHRToPBhKz
a73oXLHVuLctS2couVzhGAwdf/Qu9Cvzs9T3Rw2KnPckh2HNhmSR0FPb+n4ByCKm
RrSqYPXfYwBB/lhC9PWh0dNQA7U/z9imSOZQZjXfBO7N9MGViOzIa7CBJWykefto
eOLYDNmrnxr4MF7cF5BGynQsPGuN9oaJZQ2ZMUUjJDJmJpUMRcZO6BttSKLUhSeb
cMrPMn3bOCixVLTXZ26Fy7FSmTUiyT3TOXAHIrLeU9S3PzcMJEDqJFpnXizs2n5u
LBIWzyzda195xY3184DCM1RVWQ6blI65Q9WrykC2ouXSqU8yEmHkm+izr4TvpN5s
hvyzniEPhLuT2Yx/AObijqp29w4K030VWXK9OFHFqsRoyeeM+RTXdhY0ErogYW96
VRFYR5UdWH9IQUWJLbo+qgjp6Qs3K5jbKsC/SV0jyUorGo21V4BN5hRPf+T0PkAu
eS9sPD9aEOit9F7U5L/76lbpclfFsL9VktauXuF+qBuTZHvvU8ZYgPAzfavqwrvB
8ktjrIsjY5mc02I03jmUxv0GM/c83Oq4oLrZtzO/xCqDuUaTZuSBBRnleNsemT/Y
UZLcmxMYl9P4YCzhGHKrvIimg/0kJX67SBlADyuw182O0+CpkG3pHC8XYMbqkjRv
63q3l4OHbtRlmyFzzUq8Cqyp1tRtOU7Z+isMQUtkTXwbDH2XCwVf8BzKnv9qwnn5
j62Km6a2fryYR5FviEsxvkWJkfgz98wtDp9f6eWqWYsxJQCHFB/pwqucwnO5knsH
EXdMrGsLxKRfY9n9oVgBY9aXDUETNUuIUQSaaJrtP80C1wWYKa/QMnU8IFsQfS1r
zOwshSKkCfNS4n6RinRUq+z4Dy7qOmhbldasVgZw5KEMfBQIrnsbrrXww6g4H6fv
s8tqSSOKPytXLg4dazG5dDcAYuxe8KXVM8SpgMRaSsoQGaKNu6cO/4FthNzvIHDc
8x6oaNrMMn9J/+cBsDfshwA8a4iNogDUwK+k1nNDDxdH9LWTI/tDLQQG8FyZO6la
44nUT9sxZC1zAu3ltLGPU0l7y8x0xRWYF72q1cTIOAgi54/DHZKpDIbr6thkMt9D
YknxT4iECpGGDYg/5mhURiGo/Uq+3Ami3hBhj2j/5oF0RzbOHHLn/6MVcVg0ZNd/
Z14rCW+vHIu2bO5ptgY4rYcPPqtoXxEvQsxqNlVTR6N1Tabi4vGfAwZU5cGQo1ZW
IKns1jmIwRwQ1EBX8kGGnMFDad42WIXVH3Br+bFIeEbirbaK556rEV11587shQ9h
Yv43Op8+v4ZKMMnPgN2Q5+T1xKLy1X8ZcpvLZivlzlzYUKGmUGn2kgDEWnWoi51E
kJADJ0FAquF1RwPStMV8nsRTrobhHxa/o52D9I4gsK2JfxAdludXYGJ/+s3aXAHa
zFnK18IjaTwQO1k05knM3KZoHFBKcifd2+wdvbFNoBGp8Qi/Gr4V0CucMKEL9JCv
Irwq67VFg9UZtXt8uQPf4P866qenUJ9ITQttr1E5prcwBrQhTI5hQlaikUrmAaUL
PxaNylm5do7NxdjT8NlvR+lWSd912ciBlKz/NilNPftOlstzDJPTbyr1W02UGooU
+rWkXiP5WH6RAp8Rv1aSNOIIEFrOHsvpLCZ90NxMY9WDqfX4CKCoz3jtEUoKhIrw
qQdrAL2iO9zzHbsOHF7CEI+nDulIiDdgcK9UW1ON/IAvkZB6sV6cg7BoGlXm2vn2
Bs2dOOr1jPoHKlurie85rIbqrWsy6NHZaQhJjcoMoBHRnhbLodv5YRzzwIEdo7UQ
USa5MWsda2pJmUHOYeMnwubOo19IMVY0DgbpbhMqFSqipfprwRwk6e12/T6wLpAm
HqE304jX8P2ZSpFUvEjGPYgpfdFFqUVoZmW+k1XxyVMmrNZycxwuUI4f29XfG1Je
oHDwgLQlygONBNr6+Uthsug/i5dXPGTPdwc1R6Wi4jLbqlqqYcaLnNbjsJV4h7Vv
xDpUZ2wadAtDYRQNTxj0u3oZqfQVAwK2MyAhAnX1lQPHtiXg5cjAAZFjx+eiDF2h
ysL9PmdlIrrtS9H8jy4G83Jj3+7oQ4t20G/WxGzU/ajUrZcPyxWzK3fdX9DOS3ZA
fhAVJPar4XG2b3KkKRoVvvVMgw7yGR+XWOdUR2ksTwCaKsEFxeXtaScfZrPij8EL
wzEzoobGoxQY6Nf6E9/kZwxKZYT0WDv/NEhw06O6EEhnEoIYnI5s+xKq+amnRcp7
tFhTeNs7/zdo4ecVw8VpGTe7L7jFcFLB4+eRbwI8wbFiEZSyP+Kj0M+6FEf1PSYu
tXscP2DVYNen9DUyguBp5h3ipE8/HKmQPH7E/sQa9HxuDsJmGIzMEgBiJZ1+t6lF
rsCXHm0Ad5iJYiiTcSy7TnhTe2MlhX3kq1xIiiSwDT+ihHkaMVlQPxBDHd98EZFA
vFTInvp2HuOwDbXM5eDpRSD36WvhYBAJ5GJ/1S17B6x60e7C49SXwumgLmZVUedr
mSoWm8/yr5nIBwMD+Rxh5/ocBJ1DIkkrPIBTWBUG8X0j9GnenXiIwF3S2X3nD4km
YLphndsazolxpG4fOGhpcBMbVEnePPRdA1IFRsKPGxLgW/bLNhT+kWkMkghGmRZ8
8SvocMvpeenOOGCOCmiFrD/aDoQ4jOCYJJjYrFGx9lDRIhXrYKz/41HlRUCFa1Zv
638L1TnwzXsra7HOtCtoFGD3wpaE6v/7NcCcQB+yzkbLvsHRuKjDlzNKrsyW/PUg
yUNSeNHNsqutkfSk9vRXoa2KrwV5oFByhIhFxDiBpeED9zouzVUkFYbMaDhfJIuj
x+bOf3EipG3aaDz8zrnAz6M/2VAGV7WhVYfYKzuIAtmNz/nnUDc82es3og9SH5CK
tjVFqG2/p/bHzMNb6t/3x9818dpdXzxSZQnGWLn40TwiSPdGMEDWmblrBVFkyq9o
gfMyA37hP7rbReX8LPMFPkHBuIaPqUFStdMrKQvD32DdRQntmA6VW6gLKTo2kK1g
ezZQQuU5V2q4+aJTUxFnreg0s7jn8bl88V5EVKwihQgKlqD7MsVNyOAbAq3R8zqZ
v/Vq6kMyPf1ibnLYfBKst6N58sZbW/aTDR8FfD4IWVcOg2kCOODDnaDYrH77Pcn0
IyYbPgsEb7vdNBQosNeyJ9CQ2FBo4t4bld8WG3WmqIgNQ+DHUmorgdo3hVvENN3b
Gc/+p7eiH4kffmKAGpU7wlhf+GvyM1UEkcNL7kiIefJiVgUlxDOtD6wCy0q8FgPm
cIiNDu3hjnpQcsk2tWXLebO4YEWj9y1YDRZsW5dIM8rhya7mLaBUj6wnNrZYlJxI
Vk6G5oXs+gniItuUY8IFKS2NMprcLw6ADBmiW1QpnxmWwkURhqXNW1pB6i1N05vl
0rkqP63+UL+hUAQnyeFtvjDrdWOsG8VIyFLr4wA3sXsvE4NvtFxQhGyJxsKDQgNQ
nu7vPWso1vJ9R2pjSAWdbdGaQUhuWS+dXSi9ADAm9ixu6uPklmulMephn7bEXUED
d1J6SOQrHZtEF25bC4T+pn/esl7B640LxZz7brv9kVNSa6TFFO5JOcX9FlhYyMDs
gpM8pSkVh5z4g7BkR1OVGRo2VIfqrs5xlu7vEEftxdwUrduq6He0KTiC7leAEjB2
JB4BlYRYySRwe3Jk9JlrKvflRs4JV5NimhPDPi3i60aMH84VsFZQeVfDCngJeJLm
GvU+1GwkszIYjWUMZhJzjwRvY4aC2u24212rJdgND3LQ8hN50ZBmDoUeSByQKb6c
eIy5LpIiSab9XHRkS96kmx6sX5KI7OeZ5Zhq7EkqpkRkOLrLHX7bgVBtajFTFIjz
ZS4CYCA5JPVFiSPvWNXYjqDRGeERw8UP5x/duu1YvckQ1bMQESD8obwjcfmAn5LZ
RbtCzHyeCXYWmG9OEjzrXt+A5wopo0H6NygOzTlISBnBbByJrc4trFSHFJiIMgBH
qYc4h30a4dl14vQqR1CWrRWFmlpYFvrzSqI2DIxTdjFwTWdTGF4aRPjJt112sZ2x
NSgYWWa8crsDo4iE7a6+OsRJBEodS2V9vOIx0eCIaXXPNcXLukZ4UGSijlJAy5RR
ifq5N+5Yn68E4deetk115W+EY5GC4pSkfhQMkcjyXTMSPe6ZrPIZVFWdwxHCahGQ
fKkbUyJjBl8IHkbcBXiIj9M3Mcqd/PYMC3AU2Ny1Gvk0XcOLCNJDZ0WoXgy+4tP1
p5b5aOtGpUAjQyr+lUw2OWS/Clq07nBqRbxgqmQlP0Qg4jRWcILMNwxjKJSBc7BA
07UHgaWXVJLjSU5KeXwTQynRbuqWFrDI9C4IN+S8YYsQKxMULLeoAV4RzACErrpW
0oGvtKcdrmjRqMYfQnYwtqRByF9zy4YXZ7tlfDhTCeDKAOVGHJ1JHhB2V9YiE+d8
RW6bsLq4P/0H0wlCw7sv0ZmwmFsOVeKcEhur/YEz7GEXxR58pF6p+oSHbQxd9S4J
yo1WkDfDtj+X2c9lx7jRgXHfZpS8x5uBZXnzjlMhSX4lsOATAU53i61yjyBt4h0X
CYU7/kSl+1Ili5VskQqaf2+guOPLrp2o4CAGVZuK4LohIJ21Wmc1r2j0rkiqlCeA
DDpQIhxvjAcIuV11ZEX2xARJTm/pvXBWMXBNr2Lu1YmYw4xOq8q2asodbmmag122
IE6gxUgkMIorzLgTpdTAB7pm9WOE0NjSDZ4kiE5ZbBsk7z3lIdBdFgofawN9uqpl
P4LubUfupnOO24BR+7/09BA8Uab5NuFBlqnP8g54aKyQsGsPzOB8kHF8pqAOYNo8
4QF9Sstlc8fTawkphgYPlfYdnMuf87OMzvFKFJ5i/LgQIkWqyU2fqvUxL5Ruz00h
QiynTCNepZtOPVVwK1tKepcMKEBU+Fl04LxmhzJz5gyR0D6kOoNcg7Qaly3GgcKN
H8IFKOPPOn/nhB3rYW9i+n/aTraaqPRI41ZR5uOhkr+AoJDto2zO6NE1teGOHDmd
WCKBX56xQDGmIoEZKvLF1FSh7EA9CL+f1HusWfKFlThvjjS0UsCFWvdwjRqAod78
5ez0pjFQPrkWSD29UNco4GdbMVacQDhBLvHvdhVsJ2GqqX+1j+ztsCYhDHvl5W9r
ZP2bJdunSy5obICPhxYnlMNFB/YCLOpPeDodcJqt9EinwfJ48qXGVCzl+WQ3pfdN
KyfPJC55rJ+7eBRcNyS2ewK4cOGoi/UJKNi/N7BrfsYAT0m9UDqABfHogS7LTY/e
i7/yo2qyU3++Y2+hAjgGIVGCbYu3+NPGr/M6IFNvJVUn1txLznGo4ljY3WZaaAhq
0SJsi35KYb09Gu1oqn2fYOOmk8dDZuRc+giZj7CdyzONi60CdINjTiNE87vrPDvP
kH1r8Z6bcPrmCImqNl1sp7SrHx7Hqw+AUctZ3gsb3RP1DvIFvPwqn47bdtQNfAKA
KhES1HoknjtPX8NtiIMJ0XhhCd4mscTnPZW9ukEdRCueV/wxwuoEEclakDMgoX5G
QFoTfUncICIYcychZWj1QW2/F5rpuQNDXAbKB40YTFi3Y3rPsEgyx8lLO1QTR1b3
hdoIeu2FuolKnwpSSdK1RmfgFBwK/mauLOyWJSFS78oIgIixP9wKCo6HnUUdEqsO
M0RcqLWH7AvobTyH24t6mAx2xaHX6FbAX47BIUt6jJ4MW4oJn1kE3EMOvke9TIkV
gqHvyc21yJ8XXamVqhnm6hypQMltzaGlGzYc9dVLLuNsQeDe40bQkjFqTtJQpd8w
SuIUGzluEYGyWmw/DCtF4x5YYdPN5OkM5RvNPoHcInXUCQ1/rHlZco2QhhXxMTjz
x7jzkKeWycR0fCjmHVshEPePeuzqVaoLWa6jfOF8Jv6YPiJfzTx1oQvmAFAmtZ82
cZP2oDUDwTYTHe1SO01tR3OBhLpLKOyyii8ZByZe0yUlU1iXA3ogVgBLFN5ujFXi
oQ47m/vm86x+ok8tsoMBBVlaOQLSUuUHNTbbZcIpn4L/MAKD+RgA6J3ojG8uc+PY
fZMLffDqjbFiSLDDbjE6doR0KUK0f7k4q0qEnvxLx/xqeLbfffvb1QDX2Pr8Bqq9
VXiKa70Cu9rM9yg4KnO/4g4gr8sPyofGBdXg0quDw8049suxF7GdTsrFU5G/1PkB
W+CzhuXnGiHG1bMbyKNEw/GK8cQit4mTVYn4nlOiXs90M4I3hNTOf55XoHZraXKx
E+wku55xagp9cYGKm74tQMnIx7QXklDB3tyOvi08NoyEV985l4HZGb7X8FlHie0k
+rPzW7sm+td/P2zwjaWw+1r88vn7UJZJANTChYfKfSEBI3TbCTcexs1d099xUcG4
MKjQD/aKjbLG2mVaGMOG+HAytpi9sN1GAXMyzi+Q58iipUfH4nL+LslmQS7A8UmH
lJ42qjFuhRC8ZmTfpHxblcIyEeIHD295rdwAk0dZrOcO0SY2/UpQVD+OkyoYmoxV
bg9IGLC/nEGEuxFbqMXdRvPT32ky0y0jj/dZ4b05bwwpiRywVWQqwmEdxKn9e/Bp
VDTeA5XwQj0dlsv8aGzY/SFv/PvuvgfibDbLQRt1psYN1BZS2gNVYhBkWGz5kUm3
nVvhFJpDlGwoP0q7UDAPueHoHpDPcLC1mLYbj1Ga06pSyktSsNSmmE9KaNK1eSKU
piTi8Vr4S3j1OdiKhc2xRB+7QEul9jITipTzazhuYfWdPaDA92XvZz9Iye7DJ0qF
pip4+o/kaavf38K1nuiilL2fdmy7TykpDhKi52Vg6oL+ANlvTs3+9AZ4OO2SzZFB
TTwJXnnhy4sy3EmaMeuCCT2tR7eIxSxrEJ0hBFg8kKE5BT50JjKerhtk1l1klK4u
JVa4ZJ9w5o36XVDzH+PEYxSWMBQ3mM7kp1JdA2numwTN/KoLuCkat9eItGHg7SiA
/z1ENq8sf6wvl70wFlQ6JxN4dWewcx54CAcdRpxFDwx+7LieZ77wiz/gT4i+d5sv
hPSqhebnXA4XetwOc4Z/u+7lqg0sYVbwIT2O4ARnps+eaBxsxUqDXQuZp022SYww
GbQCbMzOzTLWS0HlQhxHZz1AcQ3/sa7clYOYrv/+ib73jPyb4eJ1O7zExiEO5ads
9cZlwz8vtMFLZ2E0z2A0uge17mc8BcRfER22BQNgBlvDuOlXmmI9MIwkHEFsPQXX
Z7CzbW0R2vt+0p2qgxB96ZFomq0N8llNY9Mbu8fd+3KNxL0D0BhTbMdGWgtA33dS
jCuzpRC1RkmZ2WhKwL6k5SvWtH1SJE+DaOjRy8Wl0T9pu6HUq8jWC7MKhCDEQBZF
BkOmxKu2nDUn3xnRG/Xut626faL+dNsEV7Hdu3hYisX0H61XmzX8ew0Jn4yHkfnk
diO/swQgm7AQT9gIGlp7/O+YNkZAxfgZ9RHp9exAC525FZOW4yTXkdGorGqhcjE9
6uE2AxFU36c6d5r/gyvJK3dWjYUAie+q3q97xm0Lm9PoEijshIlRm0/DEa3aOdUk
Rto1WIwwCRsgkwXJKTJQDpAmtwDvPYM0qsM/cA3zg4ltigXauN9eC/Faqq/LgM2X
7259Z/HZsmSlTIAVo4JvBIrmT/EeRqoEwzQEJwPm+2nwiPPf6gQ1h/B58x2G/5Dv
d+Gm8DuP+PE/KvzsvPJYwLQ+C6WvxcOSsoPb6Cu8JM9bqVfEd/JhDS77j7cZ/g2N
fHLt6AMHzvrzwifCy2vEMZupAFKPgA7fJ0lOXJkGRNLSGUZnqHlgMhKtdQhCQHRR
Hz1V1+Z2g5eKWYSmO8shmbhgTP4ulywW3KpE+j4YeBT7z5V6Qxp2hJhOgDIS+bco
bzHfV7EcDtDpI5iGJrCfltXqWUi64lt2sOnZ52Dr5HGPdcK4KNaceh8SsuGQBN5k
1jHm5dl2EZtCUmfyYc4I7Rrv9pbjj6XcyF2YiL7mOKoktTGXST6NGvKBUy76NQ9R
KtOe+azpyR9409nHlAIE/Bc9xuaZw1hLCiE25/8KSvVsDvpFKbDUkRpV0NxKVX9E
Po38BZS1g467kEhemRTB+VLAFDqYLh8Xsw53iIpB6xO9u5GVUKXBnqraWpvn6qrG
rJ5Sf2fbiN1DeGmnA9w1EVQYv5XmoPjHcKWTnRUXWHXlSPsUka9WUKnj1sUOsrlt
dFt0Y0BTGUySVQdhI5hZill6wpZ2+jV0PxqaxarrOoQxPxPEOXFoO4vWwT5xOijY
oc/nbj12A+55BqPSLA4psOcjEpOnH1+hnaOphnlPgKflMpUfgbJxdd7B5nNmUOm3
BLWShWJUIGTpQLMLzVdggBzH7IzSr8M3rXjBJe5JbZr3JiDiwh1C3YbcnBYJQGJQ
Us97SAbFaGXek5cQbn03w/85/+KNZ29pZvGXjvdeCjaDKjicTvNzWj7xCTclZe6k
9ftK5gRymu7nh0zpspLGS4E5oRJrYzRm6QcsimJ8aU7PoctSH0iRVGx5kRsBzbSY
MboVFaY9ZirjxyHc+b1tQrfKPY+GG6xbZTYtxC8f+gZIrxENWf1yT/4I4qk4NbqI
UPqR1e1Jmf4HYgSAripe8/dNpvfE1hIRd2xZZBjp1QTP++vaLzeD2p/U9QCnyUfG
um7MJh2ov6XEbngXNwv2OnFDcUapuod7ELf2UCh0MsOgPUrS7psJQQn8if96Cf91
65CqsACkt5a+fEFQ73PV6ujMqzug4/2IzaTOeiMN+Y01Qi1ZUwGyCYzisoG13jhF
+Q3Cfp0HX1+kK1FQDCaBAoeaA64neCVDi16+BfPW2GJq2P8NCehdZOM6RKRSRPat
Oscc15ZP82K0joEKcFVVpiAQKhWnXnxWaGgave3OJb7X3CZ/NIfq34KO0a+P7zRu
zXpVbXBYR4cb+ebBedR465o4QiRimmkOubs1cHLqjYx+mb8tug0iNGule4QVsd/a
6EJLj4OH2vUmXmFZbW9SrcVY6/nUZwEjwJ/h4bNtyXjcVznb2u3xxkgXBIAGSzvT
LzjWXD/KK2yiZ2mbpz+qCpDba8Tv5jhf4lMnERVi2RndLSCX/koifB9ABU7x3mLm
sLNf0Zdi7NE9AMJNew6uM9mzlV018PzAoawSaXwKXoYOnld9qiCJ68imWTtxQoDi
uayChMpegSGm/3n7wX41nJN2HJ6dMdNvoQOZ/dolA52jqxDo9BTvevKwRDV8cVtf
AcHTMDOpJsMEFuOzJOncPsNRs/f77Dwgf9I4zm9Ac31zJzrV3uCITvGanIHWq200
70xSAZY1b3Sa5DhzngvDlNm9RGn+7q08Ac8F92YO3idoAEiXImy3eA+54EEYVCMG
D/HcupwDUy5UWv6PpG1Ku8q74CwSjnB0eq48Q24aj01surm0/EBfFpz7+d08UmQl
p1P6THR4T9oOoOGRs+alTcCUBuxkH1MxZcG9SeCcw/RhoxDxn+MO4tWbWk4ZvtB1
0Ny3UbVZagsZN8TgCN9zDFf6by1TZqHgg4s+jakG4PbMtvXrAz4u5ToQAMNc3kT/
dPsiCJKj5ZzBzneO3PAQbSt7lWTqWYcyPOQ4Q2L4n/H8QilCKWwfmvftuHjq2inu
RKOTTyPpo6d7qXRPLbigROIO2ZeXOHhex6h/ho6J9UKJgLacGz1GRTZdzvp60ttm
4xX74fFDWQp7ESWBchRsFpvWPWA5AmhJx6x2kit4SCcm+IYFx0XIpl9csQsGkPtp
RiYdCkC2vJGwauNUKmw5hFGufpcwdfa6duFtJu0qmDnqNneET9+nrdn+vXJqBimx
kg8vq+g3Oo652hK85UZWQnzdq384zXYHh/R/zP17e9auLswrT3vMEV0fJNAZz/oI
Rj+Av1DGlUvuZg4yLgpiHumCx7OgBxX0B5BH3EqnfkWTU5H4S+b3sgdsXI9zfVOn
4Phsit8Kg6Gs7/pBLmzeXe6wmL2gRMGFGX3nSSVmmOaopzYtA4IYhOXD16aPsKwh
giLhN0pG+x5Q+X9sKPfkqO7yER8a2+TPZvSBOOj0IljPYTcL54y/YUXeKEcXSo6w
Ufs9odHP53ipNtQuIyLceL0QAkiys/3YpJtolQ+RZxieIr5CDKaxYwaTedmh5uZq
/o+szWbl7bQ2It04yBeuPGZkFRawFEwjIo9rkmyoliSk4hYYtbPXXwTxgC4Aaltb
QSs/jAhU+In6GnLRKJj5UYvSPi3A2sDcj+qENcJMim+LqFkEbE1wRNdiQE+ENPyc
DMXn6uQl2bAvncXAJz3g/6BIDqR53wk8LO4EvxWd9xf6NX/U4tfB67Y8qvICTfWJ
kxfB4o8Xx+xx02AhD7n8dUbTkGC6k9CXIdoeVnAYgHu1OyoIoXiN/MVUbwGk2FTa
H+m1bWHG3HR8c4uzsrXYrAzwfzJzJpXfgBp/08tin05m1CA4XqHWnOuT1hIFsoWP
RwcYBw/NH+Ium4BwLqG7gShBSspSxL5dc5R8C1AC7Hs4+ZXSDMSEGcrgXqOnrepV
IWkl9OkFIAumUi0/vftOPf+dVmaBR/sFBAoXD0WqH4fVPtVhX6ucu8n8qZIrlTH9
PGv/QdL3wHI3UcOHynx4wYnrWgAyxIvN+XD4nCZTC+ZP0ZsMNNyQ9O7o9QABlbpn
LTzzZ+/cvgYSu5ruwERXjrQ8TGN50VhFAPYmNzr7KMDx5gCQzEYm610UX7oAPjAA
NhU23W/+VLookeGIlfkRjKp4AEwQ197RrKTr4rn/JN7/PMYpHlJIhujiAIcxdOY/
QbOedpPKDNKpCvFK0F+H949Le4dAq8F6hwEUFmnWfC/mionWk3g+hSqfALBc1eq2
edrjGwyW3LPQWcNdozk8aM/FkCb+05a2+HpmM8tDFxGwffqVL2jVnGNUe/Fr/D1E
Mv7hlkGkGDucqFs1K6G+a1kE+2k0M6GBp/3KNSBj9xdyPbvbjhpsf5br0ZD+c7Ge
t6kCGgWR3zLc2FMz4alCAHiFEkon26/k1ND+wIYXwz/RpvGZocK/FAMPKJ61G/jh
bRp4iMeC2y0IK/Qyc0Bx5LujDqPKzXWEo5jmmnJa4mf70DfWPcN4WiB3JVm492dm
KXAy6+ML12qu6HEUkq8/X7XypQgEYdWo8/wrypgJNYGXr+/JHZhz+fvo2ep9G6gL
Od1neB4ewecrswyf5CrZFhk9wgLkYRTt08BylvSmZA6k+dDQVMIxdKAfmtCvfMSi
ZhmKuRS5RuSkWxGB9zU3xkPRnIuuZHY9f3FteX89T71F+YMMY0QEOEY0LLmMotH4
5ANIQ/i2vsn3Rf+QoDgY9KqnfQaP3ogiznkpk4ODc1eYhdwG5ZB0UsLU/m4dHm+n
LHzo5xhK6jGbPLD2a8C/V0qZBDdhcYbi2hFbtIpQ3dEpLoQCNepWE2SPxsS4h6O3
zdP/jK4nb3xSGn1kZACDR7mTMHTFDXh74tJ+fFzOil6U1UGBeRANuGoHARDcPrA5
DQ8CnwT8d19kWmB2MuyrJoM0JqntjuquVGIv/kOPigTWRl6dW9UOWTicwgl+00ze
rfaXsXG0jEfDz2wb4WgnW0e15+0Jzgm540oIgIsH7FqPSLmMrvOPCY2JDCdJDMoT
gnFahpjLKayc2VVD1tSlD16hv6n9Oau95Qlnd8T1/l2K10l7G/sxAWotZI4lkXz2
meYOMudCMhvwLmhb/yjs312zk10Ds14GPCZ/8TmhmSLsarw4IzNKOySi6vGb5SVY
IQ7oFoREyJF1uN8Ry55FQAqkK5CwpV9CoOedSuN0WyvHd1pzcL6S6cZGbrm4TSJ9
jDX2ud6hYfiraZoc63naYHVSAhrc7V2WoQJChNxJrc2r1QxNh6UGmz+/rvE5CfRR
hltwiym3pVoVVCLlIGX0WOEwmlrsxIubNIO9f+AogHZPensWZI8K0hG9lC5sn7B0
dMppiu608q6hHDePIzXkZ+IyVHMobi73FYpS1xQQEuVWfumR9gKO38dZWNIalPd0
FSdxe84urHhfgZzdX8b8Zukja7iu6hp1COSKYGbRfWlCnuhYd8yOgnGJedn0QuoZ
+H8sxeMaOaXUikY+r1yYlltP2lbJnFdpXUXJVFRy0+Xy8qv6tIfCXHPi9ZhB81U1
FEr6HtkV37hy1IV2IF7oe8Mnz8jsJgaOBQtzRaBudkjA2+wKMfRziT4Sw/nSjUbS
/DmLxQ12oZJZ/99no+pVl1+LbwAbAyJQR/UFJLx83i8xqbHZ7W3i9WXimWdyJO2t
NyZ9PRTawz3VfMY+boOa6uFZvhdsu3KmpkiF3EALHcfF7m6wI60IwTaqeo37DcLK
Y40N30hrFQsefM2PyJvzuq1bBP2jUlAhcRwpFv80TwvU44/tGjcFEu4NItQZIv3K
LsA6VMj83tVk9DhQ9LDw99SjdoQCxbnirfEhMWQIjyj8sk14Y6vvy4ABRMZvlfKW
Pyi+MvLj+mN8j+heuugFR4GVAeuLJ/cgUXX7sEa/WsYbC/9Ml8i+6RL6xmZVm4ng
IT1B9KKAvHF35xVvERwFijkjJTCTn+K7UxglVq2dJTrpFj0nznlpvt4IPN83xgYj
mHE5rxFrO3oVcXPxPf/x3StejZjEWM022YXSFNC7G4OUQ5A9kn4nsxvHXZZbgAgj
Dhqjq3+H6Vo5oW6VYLBnhouiB4LPn8a7dfhkDifnBv2wss3wT53AnLiEG7K+dTae
nDK7ud+98ceYE5s55YGsWe8xi8LfFtAcWoihGAOs3lWe+ZDLfv551aG8U2AmOcNx
f5djl2rLNqo7VBUoSPOwBY6wLmCh2eTSkv8mJW8tCquxoluQ29bEg7GJR+cvXXzd
/54Wfty0GdnJ3J0P5a+LIZy4HvNToaja6xQjeAapFzMwrIhXNFvoLjdKPL3fa4nl
FIEuEU6pa1pFIu61MrrODTjK7w9U1DmPnu8JuQIgzZnQloBeMQsVOcHnvCxbOgXg
Y1yvk0/vytumrRYBoF7vGBen++OOnxoIa7mv0K+Pu0ZulHEyhkW1sKvaq3g7jmU1
aUnjzaP3QkAcaP+Zrf3pqz4mTpTWvOwDrdj4CbzW1X6pcNUHfnRzDqhFmah2SnwB
Y3O/k1bpsxTQW99DlrXYrGf0kEUbaYnHnGLT8Y9ciaXXQG5gUxx0zDmT1GGoEf71
Ly6P50x03CyLhsl/PddzhAViX+271CG0fMHcB/hOs4mS1Snm8/JNoUmx8iFFyh8L
nnFGvHF75zEDRGumzBpYehCPtZ5N+5JNpgKPL0squVEQ6KP0kzl4O8u3LPl4uq2i
iLRvKyCk1iP+BW+6JeoKOF4M+EuLLhbee4JrWsQJYDh88CsAJ1sleLxUl7eYdCfU
xJr8vMZ5Yq3/nkSmAvg2s66MHpOt7Iuaw5VQBYGl4N4fqw9FkDKBvMuQSVKlm97Y
vxK/04B7LgXefKRttgBctHNRiMLdSZAA1KeCSLoau0SyfSWGePWOETEoAOiS5bA2
Xi8nImdslrbVezGIsNhVtnTBikIP3q2VohFRM6xnC7PpLhtbZHo3tvgyl3wEpn/N
2//oTxarqw1NRjacLi0hzI7Uj0ZgTcFgZ9UtG8gBYlarVzHmS2ezd2aFfJZ6zrPQ
0pFpAguZnWVt6PMH8j752cb9EK/lOJhVxSQY7GIGhWC2egg2f7cYlhuF14WFtjSL
P5j1XWije2aQHYBFWcfI2/8a1EDqHVH0Ib+CoYolD1wmTJaZoG5BB6gz9k5PRddd
bKRu0M6hiluAaDx4AJwbRpPqA918j91f/Qny2uql188x3I6hqPHsE2KrLT5N/K1C
FAouSzhTJBAIVDBqfqSvoCf4Oa+KBfPgKC7q+b0/Cd1999OcGcIV0U9iarJxeB2v
kNNl4a8I94DtXVtcknVxNJC43bni0wA/PuEPlVvRlyDt3kVLa1ICan8LD2Z+nKvJ
XI+VZEO/ubCNrh7I9mu1lbLEwrFHJRNjZxvckquq2Wca3R+o4R0ipGoD59U4ch7k
n2jZlRhOpG2DboE9ELdMjeAP/jrjmmCqov6lBF45MyRxtNbj/HhwXXmkqEIrcNN0
z4kzHJsNuPJduhCGY4XoIlYKLPwt2CufCqHD8YzCg+JgHvcqP1j1lGKmn1/7vIkz
IInwiaMElomgOPrKZuW+BfE/Xfkync/JNpmr8YylcdTgU1UY/ZBJAJ2Y5D/452xu
MrqI5w5FJeXcnAm8Z6lvwtRhe2dt2qmr910s8pXT8e2lcq/Dy/ipNMnLhwN8jgOp
stv5pmVei9sVdZ6mV2xmJ0HRbpYiMtKAfdIR/NM6HJZ/uchESJxVMSgAIzxY3OrI
qNA4gtVKQuMKrtS0JjUHrR8zjOlL34kXD14vMT5TAUNt3IEiS4qKxepxGoyO+HPL
YoH8U0lvNoE6XqUtnrpEbmGabSbmyWDwhMsWvuZ3rOE3kxk9iEFV6nlxyLKm+GIq
art3ejKBkBXn9ZJh5cBxsokTipgynAWsgtL3L/X+KUbNhJwlG1AD4wTw1KE1poVj
JbwYYlxN0aoN+P7vBZmfeHPnqWWA+nwTYyt0QkXlFl6Dy4IvygTg2DZOwSUfW8rq
LrhJG+Att5yY65dWGjZ0UmkuUgQoyOv1RoqftKPYgq53UMl2U7ieV5BVFyhqIyHT
dDU19UJzNQHciwTV7K9oJ5kwkpqfWy53t+9S3OE+zR37TZYa2gjtm4GKk01IqiJ+
4QQOp6yiJCE1DnXGZ3LxmpPzJek9TpwgjegFeYPZGhOVJORVv5+rjiJwVIFZGngq
MBKOxuLfEbkak3Pt0xiCP6d8XUtPlPsln4MvuUQcqbpPox3Gj68UTEDJXKvhFDFE
ok/fGE0OCJIM08qNZAEChhqDhZXSHbotXIfYF9xiKLGPvOGHUdo5hSBP5rDKsH6j
76AbGPir+s/p/nP60L6MvJyxf7rLtv6Lkuria5GqJ4L3/HD4AK8yORg02VzlkJJr
PZgOME4x0EJqFgu2qOaOHsqJoCpsvn5jBF6rXlaRM2feejySNqDog+JGaaodibqm
ZaJb61TGb3qr6XAwQfG6+RPWcDEqjARJpCTnmfwxz5RWL+z9yHnEIMgJ+mos4eQI
ldogpJ/Q2pMM4rwD4LkVnJpo6V35EljCxaCNSe0TCW1y4Q/fKr6WLaGfmSQpCe4s
154xScuYbx8iGaXTCeVcDofWasQnbQ5zntxinx5U0MWAWxVdaChxEqXnNvetneqb
JC6Bdu9apuzIXp0kRfkMIMLkNQeZYyim2HXuxUYu8EIPzXv+P9XvYYTGXpZjaxQd
xIzW30KSMSAkMHqLCVAtlxc6gpWICj83nP9xgA+NMlXehtmYVXwehEgMZ4AgA+tC
k3i9kXOIFXQJM6PIHLGiRsfwUGl6vN50DLd4VBKeSKHoIfB+KM8PvW92UVGUKL8O
9aPC6V01ffwfr63nofIvvArSmb3DvFd+5eCd0DniZfPb80HsHO55aIz/TNCAK4vS
VthaPa/J9lGN82/Xo3dluKhIOiYKYp0pDEsKCMI7C1pSqZL92GjqJlqM64/tuB47
j2kJHNjDRCy5dn2Acn9PbFDErT9E8wOUxciTCXAxzxUZWkYoM9GYef5PFlC+offN
Or4FlNwSeRbiTxKlI8jt2EO0E3PxYpMxMCh5zftPw3LT0yOiSFKEhnHfUc9ruVpW
FYYgQ/H57YPtZOiJtgSmyj9P4Cd3ySOWbv90UFaBy14adhptnD7N1dLZJorAAClC
fSwTJShWalhxz8GR031zoLsVuikjkprUWX/TytGP65A3Idyzm8X3JIpS7togz5Ik
VU3sppCF7n+updjyVLDgcisVWUxRp4KoIpotRg1V2FiBiZFeti1U26mFmIBTKLJX
wyq+VS6peexulWv2+8VruXw4eRchFOfa3W9PPieQL8KYK3uWCdci3DWSp51KHeqI
x64eQHbwDgSW2T2lIv+WAfGEIbccw7ymjsUQyg00d5INbB9WDJgwX033cyF0/KZ9
bxdUQe2i7HE87QvE4qUtEkX1jbsQUvlEbMbguUYRYgJUZgz7VHt+meql33QYinPi
LYo2/4cFb0eMjLMf6Taz9f4mBL1h3bnalpeSZdvAvWmWmxIHm85/O3FrKApIXrBg
cluVDtF4S3B2X3R6n8PdH5AlI8VehzuyCEuF+8P5fWg0+2E+HyQ9/M/kvGjcJcKe
h8iWiKe/a8U6pQhG//CqyHa7DhyEtA0yH7ZjAmsFZBah/jx0aWX+dmilUJOizIkl
D/35kmlSAx8A5JxMiKpTLJbb57hvXiQzP07u5nZhy/OlbheV1lWvetCulUFxBYBz
dndJd2vaWuALphOdtcX7KZnGh1+hBh10YjIwJjiX7g/ORXU0w9Q4s0YnWLcxbyhU
OuLs/S4VVJSXlwkO9cDPShX8uRBHiJipzScnBdZEiSzexhr5qpkYmBIWtUiyC9Mq
xSMCgpHnhH9qw26u9SB9me2xCN6gJZvwWD/vvxSub4mUE4OO0xTJQWF2Sdduuyz6
feVlZE8Hd5wZmzWok7um9QtOGEcQmPWjCDjPy/QK7Zzke9cJGoN0h03Zbl68HHCp
1/wv+xjiF5a0IKdNQEryWutIDz2SGjmjcO0p/AM5HqLr3yUMeZRjfzQ3eL27hrRR
eHXj3Ank0vN7OFDAvGOpXWnbqMW170608ZwIVeAVsEDCRsdsAMs5UK38je6BcI2/
SSgwylH6kdPsHHNzo+sTJegJgPB0QH2ieQakWuebDJyapDT9cqoLqo9pZsQ64RXU
hEoIvCo0mTGzK5XUeCCXa6j9pxuUnX7360BGu0OhHBO7feGFdpucnML8TfRhVC5Q
nc+8pYUZC/Ff/2HlYt56U13dmWdM0R90dqhYMrOrKcNGa+eWLYQn+g3+q/v5eIp/
R/77OzVfZTO2LSTCVIpMeDFVwOGnBl4Tai2R7Wp1JWLI7KM7PjwMWM8oEisrW226
c4VqmaFUpyiopMK+hoq3C3pLfCO6RZzUWMOswq3j8a9RLCZLlInURfrsgUadv7kv
RWNAqb2hgdJuxihVtO8hckt2/jKr0kT/TdDQ1pdau6KkTIeW+QLejyCpEuUYIQ00
m3R0gjzZGfUqGH3VqaU2FXLN1+ze4kneg1CREVodRdP76HYknVvGW1uNLEfTQSJk
qVJ7XMH5kcMRJ6nxwAJ7QGRdysYKIgA2A8GiMwYAJtdgJi+hBGNkAXgw7Y0P+Q1T
S+WcUeRPcVQ83sVTzxwWaFU1RC7YOuyJHMUOW2GJWxPZwz3/vY4Iriv0wSS5j4xy
4mcikX2rJ10QITwVY80ZLGeIl4AUFifa1kpsWlLrRxea0S1wV+oNVAJkH/fTxqN+
btclL3tiwC5bLf8RrCeQNJh+gg+I3yZP0X1DsM58XU0FgqC5lzZKi7L50DrWVVOC
4xM1/9hM/CAJRjYKODuAsmd3U14l98jm+j2GC0jtyOSv726HybjZ3VpGgCYm4wDV
X7AxuQInkueISQY25T46LZPUCbLiRXsWUDmx21h6SHqMYNae4j6fMLLH1JNlBI1v
shtjjf23BbOxqWwdTRBHIJe5p733HDI+qgtQtFVibx93hkUY67CJQLYhNw0QbB6F
xVOLuQp4MrqQAYx+5GryF6Up8mLyV82ih8ESoxb4C6+QOBES37PS7v+XaFN9u3Tr
nbSzMVULjGjy6HAzEFzQWGtJDryQvavmrPGBuYd9uNwU09EjgyoxSeSnhRuhwGDx
XSxqQN4vcDpRePelZ1BG5gW+EVw+Uo3HTZ0vIS1IziMdypEW6YWVXQWdoXM/gY28
xF/kwOS3NDoZGWnhIYLwQGdS7kDe2nTiVRYtTTo3XaD2IRKpaXa3mkHkS0nVaZhr
f+gwEJa9Wp2QKK0NOeQ6IA8oi4pZg8zG+G7B3uHR1+lI/u0uD0OrnhZ0uyV6Egvs
wvKe8SWD4hSLGy8v6sxsEM3ubZItauGepxDBs4oSsDvgMeHOYoO76HIt9GseONnY
aIXEy4rWLMILVV6ex7n+or6xPOqKxZ3YLK1LFvuP7FJEB4E3ZumJZSRSrE+eqnMV
BGbK+0elU3w0Sx0O0IL0Sawzg4PfjxrIs2gvC6Ig+aKQjFzcAO3qBFMIHb1LX9DN
lel94kmtn+AIRHq2CUBIXkxM+a58Ce3G64gNgdIr+gLOxMahOXldHL+Uz9IM3MhU
mHA8X66cEzJqtTVXPD3dQjSFCxgX6HSOTRLCdo3sdl83kxe9orUWetmzHIwZayoG
z08AmDf8SJQXK+w0dxvOe6Qt2Kjyo5lOqEl3ndpDXKnci31l30GFLhLc0kC4Juc9
VC+DfLpfsJAUa5DZRDQNeNK+6cUTPRFaSDxewIG8spGfl+wq7FhndeZPRKQWIbGg
oPJwDez+om6WqnD4OLfE69c6NHZdinjRWHObr4P/4ROwG/TahQ2ENsI2BFmu5cHa
3g0uJTQcMSbjpY5GcHEpRES/VSbXURQCm8pHYRKPIcDXB/wC3wnbCrCYqHKYXCD1
llusAVOuT1lLcV7dT3bKluXC9j7PHKhfBzoTDc4SkvfN3IxUpP7iUktHG4oUqowe
hINpE6AIQ76N/4zVfT/7lrhTFlpAE7yxizRyTQY7YNclQzvvKenJdCYsWwuDOdxa
Kv6ioQz3k+Kuzzj5cAvqP1QxBdSBxm9AjbMyXUULd9SgyxkQUTeop/JZBogW08Zd
C22tfKCZIx7lIQ2owFnxoeybfWU6LZ0ue84nk2hcVtiqp7YthnBmYMfN6JmyR/9e
UpiwLRtBYnaQBPUp4VZxUdAbANSwVj5V5hQ23IB9YAIwqMc6ZgceYeEtLxlHwdv7
XU1Y1uf4CGU7ojoT72hGiDeqg2hugMpUMeuKx5Z9L5fWonX1D40P5UNwwrfRL/NZ
x4F/NAf16XT40ATTdrVHSzMPgyJDIuqi6cb2pCd51OdjOqeMZB2RhlX54MgDs1tJ
J4TiaJnZHGQuDRxPrlV9CDuKUwSC5SKVfIGaqcaZ7WlyHldarrtcJ7b8slLPE4uS
OUetVWrtfSUMTnzzoruBJAiSD36iyvTcEzuFYvqx4gcP7HNjc/DBxWgsp2hfu1bE
gltsxWmW5JFsDEoPi2AoIavofMQUX9nL8GzYhdqXldxflUYxFGNfxlEnG1Q3Jxg3
TFSDJh+5CZDnniC1Y4IsT7mpMQ/vvUkEEuIhiYHFyDk2R0sPt5obUW6IwpUgfXH9
fXFltQYTEsjYpyNFj0RcE6KyKnepXXWpO3FW68LrF4jLpQx/KvyxibNwzl1BOEV+
2m9cnB8LVqrcPDojc5xeL2obDffLo2r8UUIP39vOFZ6j5+ebDUPGogI/92GmHnfm
Lq89/SZiZdqIM+KEBt7OPlCyWQn2weh3ffXPn6BqdybEjiSHVZYD1MArwfDICB1H
UeT85Keb2ud418IXqn3pouRfts9EdpkaRZU2ZIteeeR4tr2aINJO3XWPB/oKNSuK
MI2xktvCiJWkreSC2MWv9DnEUUSn4zFjIrKUPv7G/uL3yQiBesIYHVdi58BoHKmt
ozuX6Jnp9apt03bsCMLxt7zEs3Wskobe1Ljm0RLSbjfr3SkMUD4dwyb/KWUg4CkU
0obcbo1B8x5v8BeJL4PxVo7MeVILfFjF0v36yvhMRMwlxFX7pYsEX+BFXTdATERG
kvUrL1T/cA5OT+57+vIhua+vFgC+6YzOrV0dSJsofv56ni5uab93Ifq14JrhNSDY
b82vFF4jfct8zJng+laB2rERh05yECC51YE8o/HpCKvF6DPn20dTDFUYHKBU0aDu
/eqYuQgIux+PG4o1aKyVKkKXZsvL698o5XQfPtP4Bun3OLMyjC6mbRKA/EwXVbWq
38HiJcE61mj2WEY482E61/pGeFQ6npW6h3XlIrxHOnIAYLO7DmAyJSYCZhjZIlCD
U9m4bU5oaguE8rDphUe39gLKaXKplvxxg82ND0Yy11yzyfsVzEqiwtgL5p+tx64t
luyolOw3ZqeI3KI/5FEg6ig42yufa193YPG0RkpcrzxQps6GaW/mEGGq0R/0QQbp
EFrfgEZS1jR+OVZc6zFYOI0++hFMHV5SZxpNjD1SDpu+iS3SXl6GRa3kVY3+Aafp
8t/58KdkkMlNy2NCziGLjhPKf8+3+q/uGqsfrTc2bbZFwcKbh8oGBSDXRfOTWjf7
TZ4l0022zcqdTvCGdDi376Y/dNtcI9OHFyIBh9KK1y1MJHH+uQahx5/mI6zGVdC4
0VslwcnanHU2Y4o3wO8QEHFid4iMqHWzEEDV5UWB58qa9WP21NYz/A+8ZGHO/6Ku
2yRgZjDTYILfEACbEn5qBEuFBnQYRWWhNsjSEVo6X0iFrudWcdxom5b6iY+8aW9z
Q28OY0yQLQqBeZErkqQzQVurJZpgyoJ6/yg67csaBGd5lYKoQlf0ukIyPmKGhpEM
EzZNvcXXsANwRF2pP5HGmiCjPADW7TKl0Mm9UPq7JZdnKie7NFQnIpiMqVZLdqhK
uYCEKI21lQk/Epzs795ydarZCeaFtZZKA58rN0mcAyZy3prdG9Sc9k2EdMSvMjB1
tKhY/G8aCriDD4+98YmtTl+nq/o702dnkKOaHRBdJQLA5zXxy85oHxRfJRHEr3tb
1lHe8JJ3Z61vRjkWjIniuWqRlPgCdMqwuZLk00lDTByOifqv74+yv93YQuL8xOIB
9AYy4tJknednWlpsREJu2cOlh0ObR2gV+vLFNBQBR8xZ6Z8BUmxf8Q9WqQWcGbOU
dzpxZJNNwNvVPzzf/0qYsL7oZpdglHEQiZxFURaXOzpj8YQScEB5fG6Ui23phfa5
KLsernhyCB++hcuj4HJJLZtzOYcpSkLjtlIPrapFnjd7HJbV6+sCTthWn+fzF5Yq
lHaSktuR66xciy64gi1AMKDJ90yDidoqPARUszfwKgoU1M8E7dqYJoekMxHGKgmq
fUUmz7pgTGIBfk+U/AOV2dFwi9wyJhwwyrlO+mbCEC7sG+BwLv1Zb6wxcDct1TJ5
P0hkggHdG22ikzS4RE/yuF/dRO3xgRSLgaP+sv8HC1WfXkNQaDCyVhaoRgGd8fzA
ltjk5JxI4+J6zvVaWcUmaMxSZS50O+AebN0JgJdw6ppdjOa9pgvn6fHLl0iV+zRQ
1IvnyLULr31DYc7YcdoWS+fPsR7HJXNfkbCo15qxEr0A6f/rnZozfFlZxD4tu/wJ
qkTZzgeGh3aejgk1fmvLRuLRpntbLGmzzUnAgraER8LsS9X+oPPa3cmO7cnDX/uf
SI0xwVuvf0wA/+H70WEZ/giatNaXiWx2dhAxj3SIWQEg5ZdiJK7zUJsySe/sxKod
QNzvfFk0BFHHS/E+RQF8Jvp4Srz1EqpLBuSaSjQWk9chVi7uMO5zAh3Y9a+tHMIe
anMcBt74TSZX8/s6wP+IZBO4hxmf3si7OneZ1bT04cqmvn50mAHRLWBXNyN0zxJC
7OZkfGcxSj5vfi8kFxM3qIpBkoYmWEEF1wITVufzNLljIsTeuFH/ett65HD3+41X
feLOrKDStn1oISP9xA99KT0gdKIFAxNfGS2S6eTnumDSTcXYSFmxUuC1rfFRprEC
ezvVI69yOvlE3uD80dQGRGFo3FYzHfzMNldrzmnrNrD+HhcxqgsJ7gKdzmBXst++
wnH3LvK2mcB2PTq3G3RPZ9BciJFhtMvbOpjgPdRFvoD03VUxLPPxgvdyRoAC8Hcs
PrR+smfqRqgdW0XTGeKO3SLCFmcsJ1U7blpm2NCaO5B57kS8ubmZ9glyhmGPzPwk
J3CQdF6aL4S1Qf+BHXONckeSNEVbFPAJ9zN39EwKuEyM7dcDPW2/vHKGH8KS9ZfO
8g85YLEB/tJPd3OX0CWB8AU8GaSLRXgMN+ZBArK6zFF3cmJDkkNguKqkHTGzO6ay
YMfu11Cs0isu2aLgo38g1f86g1PgcMZ9MLZ+BK34R8qs1slZn5WHXtvFoXkq+B18
c87ke22ifvmLO5qaqwWH8L9FDQomWaNMQ+GNsPaxhJWtRxNRpKj1qUbNijXt8DBl
5BuhzYubu6VXkYf+v8LZRr3LSFLSrKateiydkDw3ZsEfIxzjrVVEiNQy4EtHWg1x
0kdUcu/wbNhqs11UOzWkO+Tlf5v7bqmcJ7wFmuIkcYbxMcW+TK8NfdxLyCvOBXgl
oatSGyT4cz5MBU4Zt+Glq6Qm069wH4pUG7MLUn7N2Iprq+eTBWYr5EzompaJUzV1
SeMtcU4h8LV/SgymagQ5QWdIUuI4WwL1UtGQZO9oC0esPxkEjeCV6gHCUrmnG+ns
kmd8aejX49it9EFZlOsxKvct9ov0Q/hnpU24lEpEciXt4K1ojXR92GBQ6q3+KtgT
c9f591OZFulob+5XbBsOAIncR7pQQCDUT+yh6y8rj8YyCYXIl2PBlymAD2iQo8/p
ACm4smweQliAytPeIE+43am+K2lEIc+bFK7qWyBxJFJL5I0pxtPgmxqcJeHn0P92
+1oksCgcZjAkTNMTCuy2bJqa3q0woBq2ntbRwGI9yQ7Rfcl2N7cCK7mOOC8VNroa
rXYN67DiLCGf2S+TLsmtwSeixrAtn7tyLkK1+0xQn4kYq86GmsIo6S94YLUAX3OV
/gMoVFHQOOaQeGZjYL8EQYcPRQLhF72niaw/6KNjfdqSWoSOWavTnlfMzCmy3Dpw
IAY7qXLxne8zWVSXu3nMAajxNrukl1Z2Q9Nd9NbkzfLSLtvBdtWhK3gIVNOk9flv
mGIP1EMTCp/KYhfzxCXB970gFn01BkXjdy44naeAgd+tsVZlrRCAJAfSp6cvxTzn
sqoxqWegjLhvkDi0m9O7i226Huoh2T/YQ6qD7PFhgWPjJLx8CCKqs9H+dYeZHd+b
Zq4TqXIX2WXcEtklMNG4j8YrcRSyQuyamvZj9BoEVU5h0c6t3en9SxKt+cX5O80v
DZGoe9v+RhGDMu8b5vrljCZuNtX4VJk+VF80Oa9HCrGWhJmaNLj7nMJzKBSJrEZQ
eUPKSi1xaBDNg+lKG/dz/tElpe823jfJf0LpeMwWFY7HK7+d+cR4BNym8vog/+0h
ylySP2bAhuNEUJWbU21dNPvEjkwgNx/kSwzXWUi49voC3201C4Q9Uw6G3xdCWln/
9favG9BcOp9uDcG1TIz6hlaErknbmfroKF6nGkLJmhlkACba6FWV1bCKxtGAHIg6
7pWIZJVavGbBxAQXtp8YlOxy+slwx+DhgzsJLQqBleQ6dx/PEImRO1ZWl98csnP1
0mowZkUxSJK2QP96uTSuAQOArxg2SI0aUtyuwXzH6LR87S6/uGwzNwxIeSz4JpFh
s29d5p1oBNk3vnubrG4cru9iagVGMGgQGDgNDwbqsFQ/daPHeLNmmrsT6ckmSQC2
K2om8fRZYQqDLS1nyjyGI45uo4DWDJYwKdTLh2Nj1RYOvcTxrft2V0MrPhbq3p9j
b3vSakCfvevLnped+aPIbyk0wK3/jAMpCVH61ekQmkKbZ6SkCx9w8e9NKYVJOPZV
QDVu7zntgIL+h/QuwTjJMJ7hKitXw5vFBlDeHTdNuQ3r5JxVfdV/mWjvD3/ZbdFp
eJh3UGrN3Hb103Ix8l7kxqCMaaPAhYjJMlunwJEKadUDh8pS5Sr/gDHpYJufCD42
FVlkvb9nh6cylsfE04nuuRSxz1PwlC+xxcpbbHPkt2tY/lbOaKKH2jxwvKvdVBU8
l4buKIhTcdAF8Xiklcs/NxcPrVVpKikmrbpcOxdLnEOwFJJE/8SrVUAVl1ZJn1tK
kc6vxshMRbQ6OsHWNwdsdOZWcflxwuZctznuee8qN2P8UmdLSgSpq3EG2fRmbc3h
6ya1oQqaE7eoaRtoU0iG0Za3EEHyd9y8+YS+uGrvGXMqbZAudMu4Bp1+CV8CqWZh
Wu7PLxdOsuwSeTI/hviSW66bmHIWQ3yEOWJM9ApdUvi1VCpkzMw8O7Wdw0ztXAm5
axNbJJ8Fx102gMA3iS0j0oOAbFswqOpTlGdVE/gb0CM4nrYTkWKMKV24Mv8IQGJR
RjWa09FqEk6cV/f/nVtRGjun3iZVjXNlyXLotapLnM5OnejkczduQnEDSCAUTJaN
rhiMSqaWJPUfKaAKmHc26iZNMtffyHEK6p56FhOdOY2X2DmVgGUu2p3pYkZOkhBk
q8VeRoiiSDGrHDixiv41PHzSQE7+eoADZEPEA+Y8/BRYKINN02ZAxNjVF1l47MuI
pMUFp+UD863ufNXd4Z0l7lBgibCqZ0sKiqeQwVXPAsqTpVFFHXjey3zEjWRwip5a
9nnmHsJDhSvS6gC/7sjP725d+t9YTn1/0LbxB8LmjKWwt9SsPCLLMLI2VGEnvv7U
ic3VMCqJ062Cfv9bpvp20ICpQVWcKgx3bEp8vegtOykSmGsG75YroMsUZWPsIivt
eiMpYElMebjRgEKq9hNI91ixHzuaQDQEkAK/C0Qp6/4Vdnis2Aofqf8Vn5Ne2x9p
vFBJdT28BWUDmiI0GOG9decEvz6b71aiblGCe1psU1Ah3tapE8zElihCVhAx790p
HRYAy2aVGxiymgeIpAKAbjR76+KUZ8xzidujraLE+s/Rd/YKeBCnZIr1yhgjV7gh
j+8zlfVEgIlaU0pEPxEbIIkxfhCIQmlh9BW3P53r4Dobktn7o6cZ6LALFek42AVk
OSxYE6gmSJYUaorme2gDJ7N7C1KD70zyAhKxeIc8BO2uJB42JjNZ7ha8xklxy2Ax
jqNNlE7InOJns5i06G/gyLzhUXkt2JB8BmggOcdooi8DRQdY7lucIjDuHESh/vm8
MLNSKieqdKZxVj0wunCLrId/PUvS2buOAZutbeIHn0v4h/b+ia2SOT2soqCa/64U
Df1xcLcQO+URNKg39lOwi+8jVv0gLfTTMf1CsJ5GNFE0/Lxd/QYAFp1qyJnxv1Ig
ZHPeJ7T+nfGLvZGv6FdymfbsZkCT16y/C81uAPBkFDjjDT7IxY4BtAO0zep0uTtG
gHvuTKG7bP7JgPgiuhdZ1LoJENbO7xBumhOQkNsbyGWloAGvQCzwAE2lApQ2tyei
ZMo0ib4BoAJE5q46B09bJ26Th3xHU2m4KN0Gw56PDmvir2UXqu9ZodcZXt827rnN
sCH5+/+VMaSdx8twSXpdpB76a32iYXSSNjCXRHtwFYubOkzZAZArFmhy52YGMrxG
jrrEcPzsFkEZkr5VrWjvSuV9vuwM5iWqygHXQaZnv6WLUmipe8VpJccNcAcBc9Af
suEFW23cbBBFCq8XagEArhz/qyHmfdRbQKkQyLeA/kBkhQ4ZqUMa3LXFP2tteoLV
s9RHyY7EISCfZC7qlZEzW5Sabnrkx9SZK0qU3D+eyz3+oYQws8jX66Y0wZtTE1mA
R0b0RY7xRs4buV/UTpOWLL01+FM2GaasLdKMVaPzRYM7DiN1dXdjXJBpL2MhUil9
/pR7116fujzIBxd2zV1++1Meii8UOTERqr29rNiDytSQXDnudC68QjlEFfFpOj26
blis3GFJAn6vIjU5eAhb+gbAVFoyCvkFY7IA2pVDDQE9HOBALmlw+yj8w7eSaSRB
agKH06Vq3pDqia8gqGsazbp9+nNvVhvGpEpqxCrwiLAsBLz2zJufZMvz+r08D3i3
hSMaY8UJ8HkAx5gJq4Sqq8NR6rJcPCxDHdxoN8jYZ702gYndidw9TciH0q80aliC
3gniX/gPC6Nve0hlTWo77gXthnG7uEWb/II4xgdn3t/EvnKrsCsAJIq1E3C9oYun
WZC7R0XUo3q/2wbg53vg1qct/PDG76nHy8SrnBP7owWkXHDr+10JCXC2Grw0L5oj
nLJo2rxMqE38+0IQ0e11AZ+4lNd2EDh0kHnIw1dAWY13V+f2FPxeRyD9mndI3sUk
PcoaBChnwhpNMNE2x+2uryUGX6tqzQ21ehKXfAiFyhzJC8isTb+f1IYaZNKWaQll
MODKlGwLNeIt8z1l06FyNksYPUsWiEfNECflTmSjzLfM8gRAKQd47ZbvYGJHr+Dy
8w9iDU1SF6CURLM1/Fd024uF75CEdsulbv9BapPrGLKhKBAR4/gJh09xUpWtoT8k
ALB8pi5T0BLSTVRwoA1EGLhQm3pifk857UsKaUH8yfABe/lJIqXAsb5S+ewYie1k
ykz3nVBAlwqdrQ0mxGb5e0x+lRn7vtwG19/xkSvjmDx85MF0oDebGjkh9u6G1rLL
MaLKKaU/Hm3Znv8AsMC7mXVXtwWxW+v5tDdPVw9uZN2jextlVL0fqewP8b5FDtOZ
Zi8LsbRYWNw5r4+fPyWHFUmzOJjScb1lb0GcwheQGkM+0Mgk+ELyKpG9bARU+SAe
NIza5DgaUk2b6Mdnlsm6LcKzRI/PvQTEgOq35sf+u/nwasq5VQUc/N6TPswNcfxP
rd9qPdWZP6HYP3udWZxkcq9SKZnoUF3ytgnn1FDpAz/JuhLXKGaMRWNDUe+2RkLL
EIiG1EpRRDmAL6eMNg+tQqwPc9zXFhbUxWthCQtTXUYxNc4SxkJ34rT01PVBqWIU
OP2K3YgvDHlseTFwkSf4vPR5YfhSdnO0Mwb0+GwaApF7fnUHioKdnZwK6/e9BPqJ
xjAyJT0N72ZkKOVT4pX+bfobdKuuwYHsYIHvIHRc4RaPJ7Kc6qeIkvQNHrQcCM6w
c5szJrwFRDUScSzv5ypbBShPZ+ctTDZ6zyRdwxfIpT+ahH8yvCsj2YTPtqeRUPRc
M7L6KO76clnX2iQIEFGw1qfWXwdW9hVyIDSfoAO3iQHPIeaOTso/fFqgYlZsJgm3
99Ka2PoyQEBQ+5qR6A3xt2Oxv0HmGbSO3bZuqIbDD3PH1cmVAp4GmpPQ/ArYY2py
ZDP9qqeKsmEQ+TObhBJrcyz9cuW++zEfgfowfDJIl8ildFw9b+KmTYpTaHrzJJ7s
+ACWEW7e39MlhFo+OzXKMCo6nVipcaVijOUM7OYgcg6G/w0kzO1QZF20lmr9hY68
/zH4bFLgfKtZliRj2Gv4iSbICwDcNzw4ZPvdU9XNjpIXha6yGW0CNxOYrgyeQAQH
RnGRfg9nan8F1lCxpxPTB4tUd86HsG0+DCjOF6mnXQ5aSB6g2nON0PYf9x1358Nb
VKPzwcyhUxJG2BPi3o+zM68XOw2lDYxyeg/2l2gkOb3AG9qgFi3byZbnrLYt1wMU
Qo2bgcijUHsajJiIAVzbWFr2cyOTEtDMgSOOY1S8MLvZ293xa2nvYXk8/FpwLlwx
Kpy5epGBf8QuLQIxmVkYQsKU6EHDNiWIOz4XPcnyTo/MfQ6RrHHOtjHbbza5gNsI
Lv0Hj8humrOTaRzl+uvK5NzTbgB9uCWJYgoaPtKojQ5O0PQJyohILsdW+PUSVCLn
IIkfQzC239uhKHjstThAiDbEUYBm6ZGRJc+fvIj6Dr++F0kzQP9+2mYmj+SycZBn
31Z+qE/joSI5YH5pGFAArl3fQoIIgrsX354TxQvZX9l2vCTCdWyE1iID9i0gn34K
NZhnhiffI9wGC5iQrIBa2Y6FqlMrmnAfrC/2SYJNrRWsNrortDQzHePQ5VagrPpP
AuNohFM0CK2O7kUEGnQZDFSY1IGeX3CVNm5rNCG60nLUTj8L8Sj5JFnPIZUtQDsC
1bNyPZ7vExp+YpbSEFM5b5LgCOdS/uN4DOYFwd+BB9aVKPw6UyE8h+e84WdU/GCm
e1FMdEeZLrHvXHRXhNxCtn0yA0bCT/S8Yh0BiVUYt+/LHtHEjNPiRxzNimH5OPRl
tJ+b54iI2wGE4cdZ6bZwxxqWEMm6pPCBPeUd+E5FMsNDVHNFqNcyx5/kaloaZvGx
hKWt41EarMVjhujLCDaARa+xWv7/B5oA8ZazOT1LdvllLwhuN0RoMq3sRtqco2Ae
c1Qs0s/zgvRwYoXXRgfMN+lRwrBwmCgKDsiXUDTV/zeRrTqhifNkKylRTrGaw6Jb
nLLigQTME119qbgIywpfcgkg99EoVP2A5cJ/27FbxQ/JKi4CkPRQ84PrnRTiUW2u
jKdRyv9j5vYBRHnYe+W7Edqhm64vrJ3f/R4QagE1SQB3QoqTN3vWohJ0vx3nLjEq
gOixt7cCmZH3YXQ8CBT6WQ53TeTLSvD4Fxk8leexU4K/3MHIZzrTBBOk612QoVr2
5JT6XGBvlzl+mAqpN6717BMJHVZ4M2cFraF0Eqdu0H8h8YsguwnDRQAikKcRhAhA
zlfteXSJ56aUHzIjC/t1huBWOMW7/0PWPzTYMD51slwrCvyAe+hIeKpkQ13/7Bxy
h7frcb+ao0yBMgjft9hBvcMhWDJSQVDGxWJGV1dvWHBXK5gnJ5b1urVpXpUhQ1cC
UfY17FTrZxJFYo3ZocoILuiq+AyI3AB/1MZIlLF+KtHpmMdxCplHtBT3YDQnqOXq
LcBo5grXGykIjjKfxl39yBOXU23ez7hQvw4EtJgrM6Ek3ysvHwP6n5yvg/hKCUS8
vzYYMvCaw98z+sM+V+1ZApB5fYX2T0Md36JaSNo8n6gypiYQ1uu0E4W9QQiPoBAs
NHnLodk3xZEpp4C1CtIX4+sOo/V5NY4FJRSnoS3RxVsxvOY5JPYO12zta4dZWBE0
D84zEzliPevyC7m2ohkzKIemeeYWGPPkYXkqRrccnHz8fm7Ri0uhONEYH4oKOA59
iDJPt5a2ixDBn8TMINPwfvx+h1SWYrpa72PSsxw8jhHVqSM7u1BoAEjDRnbc+BH3
awqNWFcYBZRD0ihh/+DV/cg/lrlfIFWEoOa+4wg5mldi4ZCI8EjZTVUhkLjIJvxD
ZbcKhAE3D8c8oP2YrTYWzWSsUXQRSyLwYGGMala4Tlln3t6Padmn1bbjOW8qsi4c
YAeG2zaMaSYxCGypjpjCz8pKAd/B64dShOzhrGyAnVBfGDWh2VNFIVPS1/gZTNWe
4+hiCTUiNK7J9rfwqPajMt6ch9GYVFCepLiSQSDVRhSPTMMKvUpwjg8zGQfAaD2V
z57gv0TyvgGeqahamhqBLZYT32DJwnVA0ijsb+Uf09WDgw7flRdbXJ4Oe51e+IX2
3D4jP7GUu0vW1NaGNHjsnW8VFO3lAoE5Ru7rqIY+kPQRne94XtJaWua4DDa66ypX
9/G/4WQOklHvR64o5uRg1vPXF02u7u1RDiaZ1M3kegOM/SMD0nSnxwhNdah9/gcm
H6byL417IUNWLqk9/515WRNQ3JaVCyX/6gwPtmTrIlxsTvK9mM2cZJqdcE3EGMr9
YFZcXUfdM++KdexN27QSkZRBtyjtuvawsawSclS4sNzwVMDfjhPjUJq+84tgrEIa
K6vcL/ykfufCToI0qZfAsNDVtPJQkBKj726w1HSmDuSe+ukhFhuK4g786/Iy9mhG
P7P2mfTURWLBQ6V4tP2C8HQOxV/aMU2dctsaGrM0qv+3id/o+SXbX18oantPrVwe
031Rck+rJ4n298wUr85n6scmEn9YHM3jZs1w2NhYgBYdcxm3TdAKKe5TNpDoJ4LH
FT4DCXlcCHE9VJ3FUyddB6AaFfUx2O+u65J/Mf+wx/j5tuGKR6Z5W61NBBSQ7CQP
8v4G9WBGVMeMOrd8T8nBovQR5lWeiqHTUuRzxHfDUj34pBNg9JE+qxPE4T1UKer5
1zYysTVAFEXUQXEMjpkUqS8hrUyvbSzuxrypBkmkfkzzX6dUBgiz9Cr70Lbin3Kl
gARB4jH9lbTP1uSG9BiL0kydm2nokmvBFfNN3/GuPpNdcK/f/iNK+LtABFVzl5bf
Bwnlj4k7BMbxHdu0Hd3VzTCx6NlF/QxVDQ4azMgnxP3O9FpyLg3s+64XyMf5QXQf
WnOs+KeKfvjWy+An7adzwXeHb6J1wGnMcunsCLS2aUGF3TKfSQhF/xLlA8lPfLq5
9NOO96NOzctz7X3sLsviVwsiP1LCe6EgmVpvaterS6Kc663AtA6vzNOYcQwTH1sx
9k6XLERydru90nRhZJ3em3Yw3nTosiwEJJabqE1ywNf/B8se1oBszGO3k4JTkVr/
rNS57es34mKl55IKgNdtU5Jvi6qoqYnxc/h2bpfyhZd3hZlfZeIWaxd1YgMvTCf3
82S8JbVK/GUJKJjSbBI1TkiECPebQu6mT8A4Sx2v9jZbYTEfEE6XcJeVtYE8YH7l
T6vUFfr4HqtqZAbARzr+PwaOAkuUnbSAaUutQM+dbSDpzbvVs7SWFSLoNGuzvcfZ
FPYSzESL8MIdrxqni14ElHse9OwpfrSBMdo9EaDMEP9SnrsW3nJjMByPrQFMuKYf
PoGP44G5VgXwTntErvPhNzijy++lC80YklsihKz66uq/AIuUdF+X+qje0XdYlK9R
82jTU0Ms4+Gpyjta+KIQT5Xa/pKrGC+0gLqRk5gn8VDYoMAHuJPQU7Vu0dXCTWRL
j5aNb4ujTkULL/au17/sZfsdM6agbLC2ldPBUyejNYL6dlk/ld8zmG6vgQvIVVdt
MZM75LgjlS5pFMhl29HFq/VqbYOIQs0y8Q++7TopND50FQFyUtEK3/oyUJb/TbI/
E9tVKRHemJBTNwRFaxMpzRex2Xi1p8SoOG9kYcgK5h7wTdFfqELB8Eeg7yI1xXCW
m0o6Yxa5hiMd9HgK5G/GFbxs+5TEauIEL0hyKVVCfBMzgfwvrkY2fZ2LDsBep9qt
8FU/KXxG0iUjIy+UXP1iDqh/6ZOzkQCDTWQ3I0JbxpWADg1RlT9QFwas3w3WMQ29
FVbF2MDrsUTaQTnSbvI0vzTNojMwFY4uCQSi0PJvTdgr71Eyex5PEQl7EgN0JI1P
9EyqfwCOfp8Y0zZiYqK5bP7S+p9InoEPTqdBf/hxWMlna9JWCFrfqLXBQo+zDzz3
NxgeEG6zRCzTGj04C1cqTUWHMuaN5cTPkQPSTLwlfvlZE6L1+83+XDPK4/MvEiWz
rsCccpNz6OnOcVrPgF8cEHwl42aOX8/DnhC5Hhc61RMmyx1eSFqVXifNVJQnOvQS
sdEr+svw1wm6Tbdsm0X1irD0BzqRBK5Nj4HWysoeWgWRZKo6PcPkAYhFTDsDahk0
Q72oxtYjyuc5L5VqzMxrD/SX/9mGkzFjYlDYnTsbasGtS/Ec4NBsN+Dd+EX+XPy8
lXYovll3m+DLEbhgTILXoIjADTTVpn3OkWC/f/1b/2Z/w7u47PRbvHkuZy5SFPbH
ucmt4ZEg3sMmQzsXTcWUkm00l4Jae32fXcRoqZphKkayZ0N6bqiX5K4TTG4CX1Y9
TZDMY5JdQS+JLEGGAw3Ws3EQNhyNkD3n8aDbIH4wWNJUv2PhHQN6CTEOKj/AFfie
gzn2v4K3z2ArMG8qTY6UPY7hQ9CR4JfM833OeEFw6kxvSjqAnHiqGGDDK0aqCtUG
Kk9aqTNL51D3ejYVzd46q/FSa9+9YFDUYkR3m4RZieQ/PEl3Qb3Jqc+B4tfbpJdw
DDKYqxkOChRP47QQWhUfK4/3cvLUwcLBAYjeWtLbH5gei8Ph3Dum39hpxpMJ6kJW
zYdt0iR02gWhQcGMedmiVvlo6mjSON9OPufb3TEwx5yJBOnMi3SruZghc3tkFay5
tcWK+vNX4BuRRtTjRujQnYMCmheNSwtagGOUVL9EJPoTHsRyAOP+717BKzCAl+/P
srR6d5LhEyIqK0RPiBDr6l1vYtkSTJ/IfgNUYq/pa7FLM6GdFfHbDBgv6W7UGqJ9
PW+DVgiMgNqjzFnU1zuaY0kH3DkDv9PyMi5SX1PqsJdc/Vi1mbkGsj6pwxMKmURQ
et9HP664kdKzXo8BHDhPz+78wgGvyJWsGeAfPJltbfmK8fT7M1L2Lo1tL8Lwk+gJ
UaAR7gnyvVqVwMZSt8lecjt0p+vA5lfDrApnvCW7tDtF9GOh9+H4XZJdFxia321r
uyz9/XjWPOFwtABVGlnmK3O/CNFMJo8j9RvPYJdbtvuz3EWukgOqSGPg6F5RkpzE
HwdQLl41Py+FHSZG/7aLqJpAEDDBgHg7AzjwJx6KCuN5mbyK/WOgon8Ccg4MlWTk
ae1FtPGoWLGHzHVL4E/7xaqqBlOHSTV/VuWTIt2TfTIcnl/zBOlilcHJkxUed6Qo
zbJs/ECf/sHBPmEl5gzRLAIqIfBiwvvRRz+MLZloDyNF5wHp7M6XFeNrgE9Gf7xH
3id99WETB//KA/9O/YblPgmG1RgVDNCMcSnl/EX7GJzxyWxqd3ijnYSn2JdASa2I
0KmsRNTlQfCQibDxUnGUWUnMq5/nFZ5IJNi3qoZ+3Uykltq7rULYhEqdvviqZ01a
h6Cfk2TVk4ZcCjkDhcHd40292YHXpwLHZi3pWOPu61mQYsiiT/0nbWYqTUfJomin
YZtFCDznd3fda1zD9oNQyFMDEC966CwUHvcEdbTDYtc+jk6f3hG7h7lHm4hRGwwv
7h1qiWo1QkBeG4RpZbapcf/GsBAeHcrqE2NV9WrEgUNKpkwOmgpwnB5rdqSklpIu
0RuPLbCMl4UJjcopEiXuQt7SFDj6TX/3ZUivOk3xbEQ6lsfXzK9PUc1ZX6KlKe4V
vrwsDl4XDFPx00nhEfIEVMdCKiPjFqxjHO2nKOa9RrdxLoguhmv4ReCz1NMO2k1Y
bm6iNTRKVVe0hKI+oqn/v637lSxbre72akEaG/YvV7+ZY50sW2K76+1b/F9yII6d
YV8V5LX5cn7f8eoOkgxP9u2FmqLAFt+UQgwFQIzFlD5qxGe7y03dBqlJ4aMdDyJE
pNycKDlbUu/ak8NMe3JhqEtHnUpYwrZ+JSsuiq20EHWl55T8hx5TZYnl5T6RnE99
EebM5ikTiK9cEUX7EGFH6n1MChSCqlrCZbSShSafeBt5aIvs6Qp2NiASuVeNSJ0i
wkafqZiuvlX9SwUBuQo+XdHTIOIC5ekW5kGe4LzSZfrPNdFwIhCFyqO+mqrUsb0Z
OLpybL7tsXliOxGECX7D0IVFLbltFcP1OdecbbXoYwUtTcRwDH8Pn+RlmwQFQ7d3
nPX2sj32ySzaUH+j/HHTRiVncDqnKKGStoBeW+Sy5nMQDYTsBSK42xsyRNSh7UZF
pe5Wll2PumI6nqI56Pfs9Ek7yy3ZxlCPQjL6LWW2QrScr08Cyxv4jsqs6l2vr/UW
nxxi3Yx6J7HBSiyTGpYoqnq4SLTcaW3GYBzDnrs2Ddn6W6pXkfvlG7XDtMRfW9oo
wFdEjZoDc83WFOiSS5j8tK2KJjP7HDvC6Hmj+mZBVR6gG0UkUzCMsegO8OmCJj0r
Ljzs2hYpP7l27ncAwnxAkK7j1oSHxxrBCZigrFulLZbyMN4gI8Mf5xDLtx55H2uW
qdxcoJmyYcZBF7RMxux4lxGOePtWT7eNkn70WdqAqjU/QZHiMCwDb7Wlde9BRDeO
ckaSaB92Wlm65vyzUSNjsxOOgT7PVmgaFJCyJRW3o+35ybWRZU4/2H/vLOtyh68l
UhT4qkt/U2I4KlQYgUig+xEOeZr1VJXNq/JCndNj35cGHbWHKb08864c4+9TMlc/
ezPgaHw5eAwaM//LJlO4wdL+md4kmXLmvuoRNSC1IMu5d8O84759AD6OoApxQz9C
Br7H3PZYQhelr2eov8DHAPjeydV6TBIH7q7in8DdANbIUF07RUXjSO0pZZ0rtRbT
6B7gcTd/PKpR6KF41M/qzy99yfF7Dngh2J4a9qpIZBmD+R4IOC4tcQKcOGMgJSYI
vX7UH+WhDIMEHFuaDFboops7H7KNXkeTMjYgc9GcNECnM7dBopBrTc0XWlbJoNWS
gTkdpdcHNIQv5BBORW4UCUPUCQplGxkGWE5Z5qgShDyKfTad1MxiCDSgSVgSRWuo
q8QQlptK4lV/tBfJiu8n/OcToJHRjuIbgNNgY6kxL1jb4IGiTsR5MXZbaDLEGwOl
UkBZIDdmaju7+JtMSWEotnaYzjnkV7R1hySCn9qwsMZAscIKZ5tK+BAk/wdy4dRJ
mg7Wk2d2r04/MgKbdEjFDLIp+ytlOSvDQJ25QyobG3u3XFWnDBmWyI2325aq1xKS
6Ol/HOKXElKhjqlBJ11aeGqqzN8Ys95DIBIQF9FuYkepiLBROCSZLouA19HWqAkM
e0FiFR4WyzY5vNJDHszxD+luUwX09c7AUK+UsJTR3C87xkwyycgbKs3He3TDiX5O
F2B7lwp9qRtXGasErNlCQcHbNGhStyY+NN07BGHeangduvAkt7hwmvVOf+2QH0rI
20XEt1AQA7gSL+Et9Rwk5kRcr+cqh7L0BPNbcYz+f7vdKBNm3kN+YNQKetir0Vdd
bLxKx8GCD4rcEEyPtZ/faYbXji9Zf/HudWFvDqczMY66HvKsSRwjBPIXcu5Ceq2T
PSQ3w443eScpqERPghwGDhYLCyFZU5ue/gKlw4NwjSl5+9Q7gZdsLNDpBCdUdmdR
fNWOiOXo16IiVjg28RWXcPyS00Q63sWJyPd71GGB0vRkePvbPGrALETlp26gyGVx
CEuRR0m7OCHeVAsWI+hVE2NwnNRUlDXV5V30hBMsiedbKxk3qjLojMIP1IscNr1+
8HKtdqqCuza6h5CkkTDC9mHBKdQ5A+sFqWUYV4+0yFRd5AwJ+m0p7jklPCZtwB93
xI8DmimSPRhF1TFxGh2jcCreWdOswk7DxUAheiQkbBQ2DXA0JvsX1EumOg2AEyp+
WZ0XI5yzXLFJAeCSvzp+v68cVtiDv111MB6WLmwi1c8JhU7Yb++CrcaWnVNft3Es
nkKb3FX+C+zPQOU58lXA4xdnHRkQuKkuUhDCHw2kiiAwJZ9TlGYfLXFosCShCwnZ
sQn9Ly1ovFh9SrQv4kN/NV6gkdjz1Z5BDD2YH4BAiBFKnAXJCv62Dy/y9F6ba/3j
T5z43M38ysacUGqUaf84IQBPCj6rp33bQJHr1uiePTBOy6QJxpufzgnBkBM8Zq4l
Fkh4deLJ3x7QBbOSvDWrkij1EB+rVWGo7zvtnr2Ngy7xqJBJL1TdXW6Qa85+w66h
3RbmySu3252Ym3wkog5qHfYHb70/TBCTQY1QHtwGBuvMmoWYL+A902NdDua+TcG/
GZfuGtUiaU61BttZtZMJNPpU8pGgyA+aVX0sHEfUTdVxyJZpMSA3h1uQCfzuvOHr
aUa49qKUPbHGo2CKQ3q1GVpJVPPZLcSA1jecs0BBgoRknqe72KXWQ2tMGnR0xf7v
t3MnXcQ9WnCDfW/kw2VxsgB3yMEmmDECCNEM9g95p/UhxOP3gK8aL/gv+AACKFRm
9YumJ2K8jNAKvwOUBUaMikeE8FwKpHIyIyu3xqX3qS79MIiAk7O1bfbIeBmk+fM0
C9dg9Vrwf/J7NV8ox94rF2XDcYWcJ0OU1ozdrZkWmdvIlrLXcuQpQDimQxcaZgLA
BY2bfiMICj+qzXa/t6V9U2kWjBReR+ODyeNayQP4eBXXjiM2CttqkHVxuNqQTqO9
hZwye//HexeCyfR8XR6qPAxj+giI8nI/OsQhdYkVOKaEqUEEIjJx8dY9nOHY9z78
SXIvEepPs6jun+nMw45ouGtw8w/yionP4hNgL6MTzcyVaRSHdJ7Ph6WI/duUz0YI
i6IXyAsbTXpuSS2KC2o/F5AsNWMCIBVRxkEdX9ce2QnppVLkJM75SchwK2AOC1Ds
Q94dzgnB7tbM2XjHsOpDn3KI7HyQniFRm1o1jgWjuY3RUOv0Al8OigDrbwH3WYkU
FwLkEEL9qemljdyvkuYc1QjN7FpRoX71eH8gvKAcFKafEa3LkN3eaFR4W9p5vT6l
oLKQAMnYVgjR1pqZ1WKtq9SysfaFJs+Er0R3LtHbrb0I6Y8BeEKsqSZkPo6mW1vP
HFLYLY5QnUioBfpWbgwtlr/ZHnTQVBuesVE5v6ky3pWtmgn4YN/08daihdsHhdfq
YmwrguGWe0txZZRP9ergDi3CfPkTtVJIfT6RspsdhlePP+Cpib9QZvoDqHOtF1eF
3xWhJsuJ2iFPC2/5PYOgxizX+Me5me+zw+me/TlDXx9HwUudqTZ1RUf+nhVZ0SfX
R5I8LGrjMVPRQHT78FExoefiRo6hSTJufYoOdbySnw15RP1su51ysRBpEMXhUnVn
vKeeivCHRIEM5fC+CvLRoOaYwqJG8QDyXFQIYpm5DKZWRiCB2jDh5wO/0fqCDro+
G2uylbgp7taFsEQoCaIs8nyY0GBGpOlXMFGGXV4D9gMh8f3nC8s1KVI9sNFzXaGE
/hLm6Tebjccaqu3v5oqEbFy/fe+n5Aywieob3A4rA+Q8obKL2AyzVjDx65z0suJy
qF5268ZaK4C0bQyi5AbRfg1kI5w0nMVk3gtrRdpofxL9kmJ6ZB1WX24HiEa8v2ts
hZNr7myngx7KkfQWJimiMHjlGHW/L9BhtO17gL8UuHNNcY3Ip3lBoshJQf3zMB/k
cRRZa2OLaBjokKmx3Aln3thzHj72PbhJ9E5YR+XZtG/7L5vbhHABW+WJgB0/3KGp
73Pcn6cDNomMjolgagjDTqvrN9RdMlvvZdMXp32ZgQ6OJ+Vzdikpgl2GL8yqJsYF
oYUzTR6s2Kx3M2j1QXB3AGl3gQGiYaqIDrsQaRZ+2ue9lJ23QaJ6OrVbQoI3zbvV
ahCBa/dk48adZM3lmcySf482Q5bTATzqLLAourCvrmVj2/teXPWFBD/0G7ftul4L
6uqbsWPqb6tGURdPt+k5/5WcoVZBwcDMXvNMNewIfKo5DfH/kNPnBV18z3CampwG
tjEHlxdvU5tEM/RJexOl7u/3wk4+GK0cdi5YJIXvRDLBDnZagsChZmHC/LDZ6yMe
gMjprvKxIkScXmTMLOY0OuzLLKQ06lRFuqBMiUSx6zGjZG85ML5WHwrny0CoLRdG
Eh5jx6JjSipBN1K8flvHC9QBVOQmMmxdoqtL1/WGZbnG4Z+da+6on/yUcqs846WY
YdhnKo+qmKHmGdpjL13mTiS8mw2b4wIcIS0wd6V/bg8pliw2VfYvRh18b+HyBIj5
4AYpG9y87FRePV11pDtz2gmRufZmqZ3tnzxH07hwe/WVza6VFJlossjSlm3Jzp91
ynDVIC/999rSrsHjbSAPEdrFzKq73/kn2WiK1rES2T/RaXJKvs3MykeVDPV3YKDO
KnqfVggbdptgv7u/noBGtB8CxEG/LcEmqLl/S1BbzspDvwphuJE81N6do2Lo1YkM
9T+mTT/N9gWeshBS8XL6y0vyA2cZkkS47rpp+YtAC49xN8YSULb/zsseHn9DQHDE
dEeUddxAy4go57+mIUPkjRWoQNXvCoXNQXfuEJunwZOHUietgFoMEeJl/PQRruxm
uihtZBpJ3UN5aSri8tEUs+2tSi8X/OsRwBdARrgPxKr7N9oLyrjXkAnRQAwoEq6R
aPTHeArw+j9LsRUgi2BCSTyaXbcJKhvz0/1gtCGSQDuprxEu61fqtw269v1oFjcO
rOntuok/uDxfaMRNmweNDzHvr4x6V/WClBL8eeUeY07syNiTJBfcf6bzA5KKP7lF
w1cQQZfpmhjTHjsNHynOX1AbCTLG7W5EVD6TfvggyB78khuH4EoT9GauNJTMTgMA
VBmDrFJ60OfPlxU8pu8rtn2b9QZetEVwzkEQjC/JFyt34eUEb+OQk1C++GofVWll
eXEHgvtn+sS61moBcJMk/1luUYLRoX8+VkkfhwEQgtGb6EkckHxW25wg+Hlr3iJj
puT2p45jbv7xWyCuq8ZFty+BzryHft/irlegRW47LtRiX3VVXOL8E6TarTnWjdV8
qmKfmP3eUz1P3K4DowVZNSMnvkaQRNc7I81TMEwt0VmS8lWx0jM7r5oAAkkO+I65
CsXEsfGvTIFryR0agnlynqZSD/mkP8b8FPZQI8w3pWtxjLjOKsIgpuYEP2ScURVM
E0rcVy6KTzK4Shd3gs33OB2K5uZ8KKBjM9zVCx/QrItuuHjZho4ztxMmg5JTM6r3
SxCuIjxrrXtWXQ8NX7UNNq8V8opcYor5tLEMnp2dZqao4sOrK/Ib/nynlzrrh6Y7
Ie9JwupCxsl7zU3VC8/yP3Uesq8DPdK3DgRk00eoBaaXXPtdCRtOp4f/34Gsr5ER
A+TG/NlwNnjneP7E2iim+TVcqfWo200X+/KmFBzbIncqX0wHZPYgse4qI1JEt2dX
whTqzckhh3jEDDbgesKQBS+bcWNSVu0VjppkQUQpDYxy5OafqmkbleqxnI7M4Aps
YgjLgGMTFF/3RTkd4nsORdVT3XdY05noWfVcDytT+8xzwrk4TA0Igz1OWk78R7F7
fK3gxgUBfyEvGNIjXsqn5bJ6wrC4794Yb4FVtpCHhavuGwrrvp3j1QjJEIv2euUD
BqBRZl7hGXLxFuvDVNFsAWge5v01oMYg8GP9zplfg5N9aMsKWX0yqpwgNr7AuoUm
Fp/3Uvwb9mxw8D8Nh7ouEU5If/KK7wpXZSI8m9R1873y4h6pFJc/KHVjfdpkUy+s
hus9uyFVLY07i5iSPTL+Qn8gdFSR8Uzzgb2+2efGvCFWvi+noh9dfEMWzSSz3WYk
mOMdeICdU6xi2R5RKf5X+m7SP6kL6mZKQlSfxSpCSWBr4ziQMpsqGNpczNeKkovF
rCSonrtYNYctRelFBFyrdPJyHjJw9OT074Qd0ZPdhBqln8k27db93szJx6OyBv3U
Simk1YNN+XrSOFRcmw31hPXDPxjMvV04LyabtHpcbALmEcVJL/oaQVvU7zIlOMpn
qJEkl/vEiFGjlXqSflf0VPgOvHfcEqM/zhP/k8DoSihRZ2SeRM352NAjXk2xVRi8
hkWhFS7pQ901shltE3SRZwSeBgexyfECr86H5lGpNSipremjx1G+isOvfpzWHYF6
kTxQilKgAgWTYWPx9pPmBbddZZzTv3kJEkMwkCIGCj62p7WxZGoqHzDeh6VZMgjY
i1pvuxyycpL4wHMCD/HMhgZqXzu51t1QPGDvJAZZC7WSxvzLxCmnpuKvJ4u0zpyd
zwcTwLZ8JbIis8PswgPdFF5mdTGzW1VgHVCCdVH1Sg2khq2+8zCdgUSrYFBFUQhO
d5ZmkzLQKD9EwF/XbNvuEN4so8AKI1EY3BrLRJrpbNgYaW+BEBXCttEKmJ0ZBy6V
8nEfrUOWlP+EDqHTMNLaQ7+x3ErBsZRzny7zSpo+zA7r4IU69DV0YXcMaiof4gim
wsMmH2MzfCkEhH/BYyP1yCJgxp5GDW0/mywYa72wx+EHPc6INH7BZP7xjXQ2xvmY
OcAfjs8GsutPlCgmGlR7Ijw+ZYXGZd52DmPv79k+24v4i+u+QUJsdBUPVaOPD1VB
bIvabYqmP5Sr31mi9sINs6elKVE84ii3JXQ8ho5nN2VusegTONdx6V3vtvBNRTCw
4k53NPXpcLa6xoCNW10aiTPqUIw/luD114h6N+8K7+Vibh41FtOqY/LO2BreWDQW
LNgx3Vg4rJx/v+o6lcbok5S0eZbwCTAam1WgiplahK2XUkm6HytLODfX/XuyASmX
5kmBdHDqb42ov8rebnVsrdFKShLqaMLLkywmYpZiTKGM6FIo6W0o1TBrg0FAdePg
v8IWrBxpxtWARZCOAWkCfu2NxaoCERoFotEdyG9Vl1Hdb6+LGBYqi3+Ln/GaCBSz
ykLKMI6Ogb/415U4p9EyTeCD84doGm1JCSiJGyRz1V+Ro5MZTyrmzXlYrvDalxoy
Ck9/CCC30+Dgg60lavuJOxS2TGh+bAKWheU4C+slashuByNMPGs42jNiUUbk0Iw+
aGrASkWym0SOY1ZR5yQ1lqjXil8Kuk2cuf/OXcGuBX9LAIx6BtmdO/WkxRONVyU9
CWLNOuP7G5C+ogwPXMt0xmNUo/t3Hmlll2p5OnI16FAZkOVJfEvkpmwuRcimgbQt
fgNFUZL/I+CW5SLjkIfKhemclbEDyQjzLngicXmAestc2XyzzXGMExwo7i5Cw5ep
6cPVb/GagdT+ILFLgs7TcyqIgzM21C4x9lOuKqwlK1dOz7OUf5iACKy8R9JWIXc4
eAFsuRg8vNB2G0tr+LDPIKYQJ62mAdkzgl2/VKcik6GTYh9YOxwRZeKs6FxWdb07
fJMKp+j3wnY2vXZ4LWaJR5jVcHvyCm6IED/DJLRzaHQxAXkECTiOUyaPx+/YjYtx
SuSK/3K6Of7AhT1wDuN+vUFIR/J+Bcu/RV4rAcH++6nhc9cWjX2hxDo8QM3O+h3a
KQUZXTmHaUokN4+WjAL+nw1S9OUdA6VriLOHb1b9ZR7PDhW3+x5e1hkIhxrWA9ve
yDwz9btHGGZTtjNa37XKGUtny/FTFpmGxHnb0EqwGp6+A9nzizWfBQYuWuyTVqc5
68+YklSkx7opkbgB6ZLoGoXM6vVhFwJggfhoFZ4bDN2G+w8JhFJ8D/emkyEnn022
PIgbR1ZBaesxHLb5+NnhYJ2kWB0EnHSCdDRtiINdc9dNMVZUn/euxOGsKOAzg9ma
lAwmT/r6J4u7EE0bVpYi49bPieeMuDbCHevurlpSJKuJcYkW423j/XuMzMY3uj+l
AVyACuv8guUn85T/7Ym+HiYnec7QY46GZGLoqUZpmhmqAuuSAigPSvD2LElEnZmm
WedCIl6XcPisERUgjswTB/gR78+0pjQmMn9KPVJd/zub4iBgNWNO+L3PQFVKuKdk
WvwIJmdgalQI+QnzWhGbxh04+7q2KIHXaNuchCdNNYJmRZqu1hR/grEnoYusG/RO
9nPrQmKtG2CBPOAGkBgVqgso5hk12g1nBpnfMhnCZnw4T5D4SiiimFEQq8G0v5Kf
bBT52s+TXKmT7T6PfYxadM9E821JocnDZDY7dBKthfzO/wtLKMbYLiY3kwNHRpYW
8tX9ChjT5nt4TgsoB65YeTnoM/hCv6AFs98xp1lbeqglrJX56hSSOW7TM9as6V0J
Q9FwdM4rCglc+X6ISAL99gIy4P+63Df0OwezC52uphn+LqO6fB2+Sb1Dh6j00Np6
ADzIkwuWhpTYKtaPkNcgF1WQrGsJtrwStCCgs3CTLoY4k19TwI8EfoW9SzLVZEjX
g5aO1BzE+wKhnBDiLep1z7P/1molLDeMmrJvr+Fa5FytRsgf/BjeXfUoLQ3v7Iam
W8daLTGfyebGfWRqDuMUztIdWkMbQky/IKOdD9nhDwKOlbh6Mdm/UdabNUoHh+mU
PkLEsyJjX2zjtIL+u1uaELgq6YrWYiCk1HingErnZAjwsU0moRRsIYPokGac2u/w
zdXawiGZfTxnGTdfoXuSgDCYh0jK1Vn2Vf+ZEeGhhG0LPpa4O9B8/JrqWGWIecvN
q6uWrrE62HgKNuyDo1aN0ybm41JbRriEEQ93OVvh0E8TZQLQrPdSTjp9+CfYkmZI
tINjHRm8nemCcfA462n1dV0P4xYVgBTAMJBIrUaXuugKvUpeRfDZwx3BOrsgDo+t
Ls+pvUxMEgBoBs+xxYt8mYAUkKICQ31UfQqm97Ql1gNSLK5AOpC8mu3lbUMF4qwh
oP1FgozowAcClmYT97egqzCJDJrxfIfHRbypVvmXcSUbjvH7iVn2G5Guek4tBaT0
B5Vm4LKkmEJa3sacOV9wd1geEY+Minz4zEwCOt6y7+IxfTtrExlv8tdpuCs1E2Xo
ut/y9xp/C53rU1QXH7Nea3Jxah7vz0zQ8tJOZ37ZRxEsJWsPDhJJpAqTGa0VtDpN
eOSdF5hyCm12p9y6Su6Ah2gULeDsxajton54t1FjMx9A9JeJiBe1LkKCpUc7ZHRt
uBhxnh6Okweo0QjLLUULhpOYHZETkRDm0iil7rg2OtA7cP+KLr+/TKAJ3A6HUfvp
ulZq4Lf6PpUefSEXzu12V5Fa7BG5cXJ4YDNfE9Rfcuqi3e6mfLcPZrV0UQxhfs2m
o+TsZKofHjWqkDftiy3iCsLy2X1nbU1BpLo3MZqRgmEt8WWvhq0ChkAzqgzEj98J
Ib96MgTOK1gTBQbvO7oyimPkX0ACVbUS7cjoP0vkeV75SZyhuCRuKT6Ry/1ijMGt
7blMBCwWPK93JQAMlnh0j3h/oK8JTtl1f46tgbWi46xbuIY30MbiFsZFbmIT4x46
2rIi4hocdZmo9OQPJzJ97a1WpVBs4FUBI+NTD6G7rThK0itV6Mgn73P+yW80s6UX
NREs1AmCrhQsgm83Ev5NfxK6mdSihE7s2TV1Z2mu/h8mZIdoapnIVgcA3GZCIb7Z
WkXY/Fqk7hcNEfWy3Ldw4VLeNaj2VeKk8MIqApCT5CElE4T/CZKtf0cPuoyJEpSr
6/8JRKmZlsPrpq7XbGUrr/9EhZ1xY+7M2FqelUwu/hbVoKFdjP6TPix/17TXvY11
CKsTzq2xt6IBCbK0pzHLGRX515Le0yHWnDuDHM0R0YqYT3KoalU4ZqvTtxPX1dVO
XJsWBu6bJBusnlHU9RWaV2a+/FLiyy+pyl1BMctqK7yBJLKcifY8oU0P03cyT+nY
W8ecnO5CjgCln7rhdEOEpiBrRGYNHF2RlPZAt+7GW8bqFcGWTlh6cssd78gxnL4p
tFOovGdpIDuEMJBBpsC3mhgNt8Bwfsvy7rWKAwl7oxf59YkRv4rfeOKWMxqb9NbX
vltRrB1uAwoTJZVDxgJG3BvorjykmJIpxex/HyVdw8SnkOfinA0O2k2HwylGm0br
4PPoM3fflEyKodZG+B21FoqoXYznBnJOKPW33e7ZXsxaQMK0idyWVNNxmyMafPSd
akbo4qhtLLoWx+Pc75WhEt6CuOymZVUGrCAALwVifbUUeP/ZzastB5vWu9xR6BNC
nrQ9JU1yDrTqFxExL0773gOxacdzhmrz3z0s5MqJT7pSoz3i0qYfSCSHaANayHri
AQUyayupIBDaSLNv4xF0lTzIh1UvPbivJRlu5UP9CdTjOZN80EMePtq4BMvb3wDF
+PXs0w5Y89PWwkPzIEtj9UFiOma0QGvKrvdVWuuFmmcWS3bTmAgK4hd7YZubx0Qo
lVFrEu8ba/1ab44Z3wJiVK3+HZLrcV1TSZ4bWePkOpPzR/XxKC5CFJT8w5V8Wd7G
yZZX+H4KmjPi7caMBp9bisLisjDjN4isIeUtzD9TpBs3cV0flp/2NusxgnAYGDYP
bOkWTggVjLG4NdAxIAKQHIYuOLBnHsRgG2a8Uklw2D1YuaxIzyZ2Z/Gb1nn6rUaF
nJK/t7oGZPV4LA/TY+bbLIVNGlmCx0ygeScGPWxqiw3gNCQ2MUH/IzCI3OVYoMa+
yWraQtuZg1gIk0K3LvFjEV/LPDim1xrrEJKTNaoGYPc/QnOWSQ8+ML3tXMIR03YW
5WXqLbIH0kKJoOUpiuIqdA3AtaiBL1QgUs0wwOLwg/kS9UMQIheKMqv34MsY33NN
YZTLmIU03nww76NmZI4W2FdTdnisxtwotFqF+4gBPKfLeHp6+3E16BGIz9kt+TQv
GX/7VsyPXfPSpLilcovjH0GWrtSd9ItSmVBnwmJbjI3urQKMIxSKmJrovzz5sDfs
z7Cb941zS2WrQJxDenGhkQmO49vRCrzOCZ8refwkjj18uHPyZ0h4FUV+4qO1X7xA
EH9EWevI2ETnmcq8W7JUGuZqJSTJU4dwcWIFFTYq4j8faq0xbJDFkrrM9Io8L4gV
/u/s7J3MBjbTfbrjlVmqJ0bWDiRJiiKMYQkit5ZxSFkhjZ6UaXMbnipHglXB8JrU
TBuD6+EsNY4Krlm4OJ2urKyGiu27V2GQJDJPI073KeU/Xrv7dYFds3p3gChDRHK4
V0GVM72hIEbPRt4605zI0Iqk8SfT0LhM4ORYSZlWRb0HXSosw+gG8oNfKaC4RG+l
U4V6C/PBjaIO2NYpNjkYG6hdbiugglqabXpPUsUIzSCNhqum39nkVmKvzOqcgJJN
kZIcJCA/tMmqv7r+ZzBevb+HDs78kO2rt5laoBT1B7HowAgd6JoEYpvGXKN+0f/E
JRilwItmf4uh4ON6qy+6qsZEbY1+TL/GBz0AOni3f7wwQuVpYJABQqC9DHMqpLJl
QIMuzyQyuLrBlgM2lNfj4LWcEAjEzdJ8G6GgXgOO7Ri1Fh+CXji2caAjZd2wZ+Fy
42rcC7TGhybCk7t1eyIbUtnGjdtxMGKXvzM5LuBBBXPsz61350kgUoF+y7r2HLVi
1S0QzVr/Pc6FX0+wnkUrhZlLJqNj6Jzhj1LIWRruoQv+1MSoyV8wiyLujCybzIHH
tjTtSYzp7DwpIl089I5CjfYxKA4/gPypyd0TbAUk6klqf4+5VMopQMomlHRkGKiM
NHt/pdQGPlmO34PGY5kqlo92KL1cuRH7IQWqnEubt/IKmvfQQE3nZXDZPksylnSt
4pGhcDyCkWJnlaEVbSwu8AXXKiR2JU5mF0ccJqpo4aag5S0bA4R3nKUJ3xx8IGcG
bntigqHu0qEveNvIbACBMP7MW1KtOVDuFO8Fnebn5zZhPIUAivB3n/TlTdJoEDnp
yXLbDigywOYodUJBRgAupVhE4AhSxonnz3AtP2DyQkJtSrPSD7KN+RvlDRaHlj7r
1Bq5VWnEEVXEL6ruHasu6nZAbrHS+lmWlxk70lUl18IeBWoswJI34ozabGj3Pw9Z
ckgPMRvhd8H2LrtahTbdBPp8/0hPqFDxnwfYDXKSjCK0sl43t7CzW113+q+CdFUE
GGC8z1kwooSXtYxBKCzDD5F7aJsQb8w8MXhA+d9eI0kZQfou7dByGushOcFXGxI0
MrPQRpvrypsuL7I+QY4SorcY545x2gGbv0yPp1M9IK1vd9lirH7L4UD1ce81g1kE
rcxCDk07cxd+VbJ0DW1r0X4bYDebYj3bIgFAB7qxq9jlsx5dLLhOpuzUMqGuD8wg
S2UjRdPct2F6auvyohSux4t9yMmqtWZ6MAKR8eKZEDqmK/JY9SMYWNAi8LqrV0VQ
SbaCxouB/z7QVnvNH5fhtvRK+Jf3Zhq5he3z24SmSghWL75CP8C/JGmAJI7MtEsE
0tDxLY2vBIh0UDrcHmhwgfmj142I0O0+9upWNe5Wkzk7h1DmlGJA/NXXCVKyugcN
Y/ACg4/nlwEe020UlBnezcI4WzEiPdHLCsJZAIAucpwWsHZkeFfUoTtRyrGgJZ+4
3IyY+biDT/VPl3WnHB5jSk10ss0H/V9q2daJlhHE7xeFfByJL0l/3i+ix/wc9ZI5
uA55MO4cGFuWgdUk2c/vIMoO7HO7uonR1qYhvdK6lkDUxNQLJnFpVibRJ43s+Pxp
7+r+CgsnAI0DXS8CnZaKDJPMeLVg9oWGlqlROMChKS94283svhF7bd4tQJyyd1d/
5WB9+RW+51rC5dzCk+jbrozigmce9rLq/N2rM/DnAoP/OEQ0I2sCDlrsbKTz2x02
EX8siHtgl+jSQP0s0QB843r7xgJKE4yv7dKNq9hI2kan4CpzvZeif3UhyNUVdVI/
se1L1oBs9qmo7M74u0hVbgbBDuU9TTH60xKXcmszzlfLJRRCop0g4PPCe4dPiFZQ
eNqeJ+1WSibD/HbJKC9hfUhs3+MD8PLZG7tWmeR8+U9xmkkl+aicQLT+SDwbkX4B
uOzsde91JnH8++D4vbqwoeYTKrdk32SuEYbfNnUxIzEBdAAZFmHQbaumqMmz66uR
QKWzOtqvle3rzvtIrjUdEhJHOv5+s4FFlgaISRRsBHnUNgBTjdm3CcDVK9ucz/Zn
1bHZXWTrButR6BWeUPsaUe1dys1qwkejhsuayAr0I9U0+nutT1oUAMw6lN/R79Ii
ValhBzBjNogs5YBm+WM+LTQfYX/vtFDgahIfzeTr0VSUIQlbJUqqDWTx8zxcWOe6
aYIRX107n/tHsM3mFvDsUZ0BFBN2vbG05aich+LiAEvNVCIAOFSKD9jDtpBJPrmj
eVq6XMwII0jb7OYFkhCTQNDlc0avTepMwCUU8uL2SUzd4rQgMOLqk/QwI1kMdkMv
bPnV/5C2ld4jbjbNuRBf03JaL7EeazDExgUXqGo8mUKFu5sonBYJqJH7T6UUP4wA
s+UkYUwFZmANn481RNbdpCHAs2RAQMVTiCAqPEmPqaxAsMgkPNUUEWRpkjGcI2I/
Q3Md1+kBnvHr+l3gK1gCmKBDEBLauI/5/YW655HPWsnHwARbUjY1wVbD8bQsWkQe
KOOOWZgdWmA5Psp0yy9sfxHrWLAIGvfayMb8qOZWpKy4e51xIgWLf27jMwcR2ie+
mrJlEfehRVLHoCK4E31QZNkG6hO7hBPWAkdiBzlpYKwJz6Tdq1mm7OKUc7hPR7pV
gTHQFURxHAwE0ZN7nStwScc6fJSSyui9Qy0Qv8epJN7p6jIlna4tE7KQVEzhgGQT
BNtnr5imM5OY8WP01RFvsuc5o8iIJBc9VCSoeRv2OedKvR8EYuH9TOsSH06gM/2u
/FiopeHUe8K3Ep0yP7NNP/BTV21UBuZyDODUmLm21lOoEFs5CJVXQDBW2TOeDfus
rLfSKKUW7308tFRhJLK2TWf3pYlXsrJI79FA5SSG/JywhtB6z1Kc4F/xfAUqsVTS
OtnkwSSGoshHxKixWVXFm0B2+h7ALflqc+gz/Ku/a9Md7huAu9qy0W0OZXsS5gCn
YsZAWUhykigBkRmY32FupV3q2hFQihdlEoF3g1TFolQzai8cblzZPbo59NC83sGC
5P5xMB4TXVifMn7KS3UuRru7Q9fDkoKH0soAU7BvIf/35dt+DOYixmKUq+r24K0/
sWOm8k/9SMq/W9F4nj0YGfRet9LEhTHmaKUDnJCbexcO+Otizwr7FPIXxu7tLyZ2
D1Ei3mrIK25ym4890+d6dhcGsGPCI+j0xMQc7aEuZbIUmOOvySB6E4UIjyENwuX8
EVlyBT+hfGi+XTdaNXQYgKT2rqe8K5lLNDurqLXAGIRo1VNcPeTz3ggR6YRUoGPq
NhJ2fldgyMWfk2+YZtwZPo2y4kVfXIM0ObwWkCfkCDSGOx85PmzEYPknx7y2iiEK
fJpjsMEndzRmEmmaxYj8B3bYHYitfdMSy3vID7HQbdt+2RA3v1fkoICkbQQsVbyp
XlOABS4DO00VDGip93t53IfGLoAkGvnNK3842nn7usjHupVyyRkaSvoNoX+0TeHx
S9Ub1lP3+34ccYSEdfDW9w/sA9hn8fO6ho9q2d5WCA+e2mvbgxH0YvCN7N1bZk+S
iqzk3iEtQoNfx8lHxy4hhHJDJzFefZE5qnFXCjN5pzkDdaILga7PX6NhM8iUz5qF
G7w1Si2Bg8PvYMBWYfFdatlFefGPGY8B/7IAME3lmzrWFTxqHYvPs9fjvwSQ8v/5
O8YYsmMkYOlIe6ifbM6lq2A2B1qIADOI9NORb8RG2Tvgr6662/M9XOUJw4dFiMbl
XTjJfNh5T5F5BqEyR3VWuU41XnSRgDpN3W/DKRZqHVngsUh89E6ph4fv2AH4XeDz
TIWRU3KSmJyZN6d9JPGTFQzalCYZeqgI4vhJXdFdqpDejfhMsmvV9ZhITafGB/tj
a3bKS4P5u5Hgxu/K3xOdIHceKUVVzn5OJcIbpre5jqwBBvXUKKDE4fRKc9FUOWEI
T9w5l478daTLbCrsNwXawPGaH9XrORP/9C6oQr2IDR2H4AMNZqfPqEpXM4N1PbkM
LT/K92P0TJs5wGyG2Tp+qFEmXuP++taS8eKudFc0VuQlMQPzDf7Ws/YwYim2rtq1
pjRWgORVWG44vYTNLeux278lQsUvnM/Xa7/p2o1hcua/FBwZS6CjspdeY0LsotKJ
G0DuufZN37+2U5ZgmUG0fMErAOiq2RBRFQNIjw0iVL5/lPsJbTkpRj44FXvDvQZ/
pF2koLzVYyZ6AblgnG2dL2BSoJ3UBFc2mEH+j2bEx7YwSPET4PxrTZitBlKuBOd1
xNci4YkswscK0RA+LZcjw9y2+hF5lF+h3fYR1VYKnV/YHl6FJEVPWCvWqbvNp6Ud
N+oRd6QOXmxf13VssIGVXONwz0H4WDjlY5Ybo3pmQWZM1gC2pkXtwiuyrvYF4v1d
/q7j6RjPbu04FQ8KHhaMBqNbqtgq7PiUknvClLCkwbSeQ3L1UQO5HEeKE/ZBVb7W
ALi05tqnuThBJ1EVw2U28mb2ZlbdjyDQ4ByERCLuc69lb+7wLbP9rl25pE1clua8
wcP+zDgQ41VwmOGpM9V/pTX+425T3fca16ae27HhHVwkJZqSQhqCXsYwtoailIpE
5Fz6QjfxwjfyLuDQK/w0rClMFlY1alfkB6+4Lj3P5RpuS0nHDt5Xbpvzrq68At80
F8DdO/qZSxp8lkHFHVCNT9QyU4YSdG+V3bI52h3k3rFLqJQ3qf3H7CbM1jVEF146
xXyOfh0V1lWTTJcZbCIwuFKTFGAj/yIHm8dEhSD4mZWrtbQmdccOhENAee5eXqwO
u4o+wN28JY2ne1J9juc7dXL8V+0RLYLT0LMXw+LCoUTjMJz4FQw+FujCXwvA6SED
nk5vsXSDAQroK3llZ0vihZor5CdwmwO0ylHN86YizaXLtfWeW/QtMkpt2P9kC6q9
3bIzR5nJ+eV0iFX7itUp8WNbC53r3umXbR//5mhp3oAVgd2dpbTGUzmnBLSlGtTD
8ZOuo+usNwAeOtHazo55NMXez11vMazdz/eXmeAHV/AZSHRmIPYrinrUC7gDreif
Ul2pMSp7E0Ci4qyxoj+vlel3nCo7Ljuz/D3wKSD0xbHEoS1gDwKcN7a9dqM3T+kP
3fexiSYRNuAhch1+bMjD7i9jkZV2+DEm/dfgPa6hE7bvCzgCZLrlMPDPXyQlH2Ec
wr0J+s6qTYB6bJbzYVe8s/4/qg85wjKbL9MwCx/XjxWw9JfpJRq07DW4dT5kcHVl
FPujZdB4CKep9X8RNsw22mUXaVHfqacz6Hz6DnEA+CjBuPHOtx6Q4fw4EDgoGRDA
DaMmrZcBrI1W3nCVTSVIpaFQmfoHjY70w9Ill4w6A3RDiEMjozB9pvCb4iMqBGRq
GWEYUSZVlSF9feyTvsqerlk8Yqk6CwxM/04+8txrHywxMdZeWThrgI2Zi4t6dpxl
uhhg2tsvo3CGqZOMzqLw4bX6EVLRCKQWldL1xl3C6rFqWTfFlgvYC60XJnM/wwTD
LddOVIXaNVJXvLFNOYfJwvtzFCEYIg5YSWjTRkoRS2xZ2NsSRwi17Ib2kAGBQ0Fy
QiF/52yhP7xxjpvG0r9QUfF6xcPe30hNSv8WiX68gUr5RwgMdqAcRRjOAgNCY6kx
dn+7hwlvP8M4qr7le8JLw0JUhLcnezPOiq9nbNitv7GouxnY739wJZA7Ez+35CgE
8aDsd7UpWyyxUyhn3tvql7xHiiBJsuHO44gK237osV9P5/TtkaCgq6sJ7n4BPvxe
xd6EzfyU5pWnYRHSFE+V8zSZ9qeeVBNjuhdFV/hSptXbuCfcpHSema5vHrzScDmp
X54cVZb2QDaVyySkSQ4yX8wDTnx5XJwndNUBWu0nC294/pC6WV0AyNu6SMTPW2GE
Ei/E5ZBnch87XtztgyPM/dJzb9XaiRYtUd4Mdn6Ia8SIvNETPldl8bqqQzZlCh/9
feVpl5EzfztCZa0aql/Jh1NzXNaMNbtGuvrYkd7pNkk1o+hwWnqHFXFlENPaZgOY
utsbj0jrGAYUuWHk9aJ4Ss1VVUH9TRu6HlC0oNbCQYfJeTRcGPbuXw8ntHfQ/2sz
F4HF8RLrJgwCWyuHF51YDXgQMrhfpl2PQI5C59SfgUs8wXTzcnDbwvA8kKfUyh5j
HzJPGeM4uePIOcrjLCD2/XUYYzHfO2uv/DLBPsYJymyj3Xozgwc8mjE0+zMrElus
wy/Slq+FyTrmPnGoDivLY5mjWHbHdGj0aLIAiJlO6/MalK4/O+bKkrmiZgiDgsUe
bZS68Fh9iDF5U8gzWRBiqpKvr8fhQ9ACwrBM1cK02bn77TPJZ59tyBc9RujRjnMY
uGct4VDJnDhL5V69rKiEqksEEXjloCVvr0Ir1i2fM4AkAizQq8js99zUtlqw4M/J
QiEO6lY0fbBwGIk1zDSfEUExxG7Ac27Ykv5atapQ8XzEXZaO7LdoRDFiaV6cVaQu
NWCWeNileleW8oF45vnUIh2pOeDiEjCsG1I4LP31v7WImjspCZK9w+4F+jHyKB1F
nHoKOoeiWIJEWcffXnCYJclIN6WiFgiWjGROOiG2Ge56d5nXKHg65+VHX7JTBtQG
pW0AyVJreO3svqZKFEApNPeWThUvQlMzHxa7kDLiAyxg9htkSi7TRraoUm0MZcLY
lT/ppAi6/46BdNQQCYjm6RkF8KGANxXjRCyzCK80r6ZcMZ/k6EkodYsiZDRVBRRi
+QsVpvSHHbN9iA7mmrBqGi/oVQldtQ/ystSsWSN1pvu+a6ZaaiYdv6wQYd6Qlb8y
YPLVRtMkJMsqiVEM3T9hwR/IxzxHSjB2I8LbYbF8dTHYA0PUdLrOGpswIx9zCLCi
1toSLa3z3J7jmmOD9of0felGaB+qIBKfm91lQpQlB0SyWnFDV6vNU5fjxFBycAwc
LivH7UsGi46D6GF/8V8GH0yWP82fEDyGnW9V09tvzEppg6ygq+t3TRaVpestb5PR
pSWb6OzWR+mJu0wvgC6ZwaoMaKTfkJl2vCAJhCXRIkHLO0WnUqPoJ7nvhUPMVbH8
79NCvNygNB9UwPsUcFcQlVCbCJUWOrPDYu6MCUGfeWNJkD+9q9KtUq6IaBm90cuE
BbLFz9mhDAMuNOoBgWHoCj9odTjDc/Hs+7cWuTtMbrftB8s3poGTgN7eJ9y8o0Ds
DiCyrVdmrmqstSfIHAvfBtixERtqNj5uhQfbAwzV5Qrhzh/1rMRg5xsVCINjQjlF
I6YS8tCqmYRvDFprc7B9B7cSxyjBkEXXaijhAakme2XzqF2vjIR6lF1ex4Qzhihc
6wh2HlsM1eg9RnpnigfuPaLVo4O4c4OYQvw7zj0w2NXUhWyID6zlivJeUSA8mFMc
ZtIGZWClpsYGOW3ypz88FzgTRhLWgRb+4XCsI862boN12Zs+0mswHan0kVC1k/fo
g1ilzScj/NDZ/Y3EBjQIWcKn1CFD59XeFJZznkbdnr3fDaiT3AN6mu82/4RWUuk5
JcmF2In/pF1DV9O8oXKn+9oE5y/nk6ll2QCa75Zbd0ilzhMoYyfjPa5PO60xM7bm
RNESWu1GOP1Wm77Gp/86HelOu8lkKeDQNrKWyBmyrLyrxe2QuTTsSy5zZyHs6MZV
aQl0Y8fnypR3kkx5n4Qnu1akWpZ9zcdCY+sf6FxB1xph+UCH9gCGV11+tiu86ADx
P10LHl1un+sPXIMyKvYnLpgeQSNNPWRB2+6kJztboAsfS/kI91NaAs26+PZs15PZ
ekS5SFE2GflgJtv5FklfkUXAjU4wODHVVz+DmlysAQ5KihTUrWPIZWSnhrXAeHvF
nQSIEWaGJ4FGTYzLvXvJePjhMxwfwNdxW1qKyt94lYRADYWvCkWr1v1ArsrRsHmH
XAyPE0hQMTDdfx9QTC2J6RuS6/qhowsgVVpgyvFPrRT8GkyuELliJoZNM6zeo1/E
brAOLeEGD2fe3HXzVGaGRI8A62AGSQoshqIj/lopG5eBSTw4lkcpW6pf2PQwe7Ua
1E7GC0UiQBn+ekndx3IeCMngfGgY8Jk9T0XzSgblwYf6mcYaIvd03Zud7sqrbLn+
OAFBhGKrXwV9dKZPfEdpDcPBf9VA5PMY9tFR/7OUnJpY2O/mTS3/nvR+WFtiUmLy
7zwOmDGq+QvSXAyB2uH+t/H4NwJ+HNgZutugCVTz8Xtx+e2EZK0BM46oOQ5XWPY8
CLZvwDN+E5pgD5J4oHyd9SraCgR4u9A8at6r6vNAhclzTYooTEdKDMoh8gs2FmW9
GG/nvcYgh4oL1YFbqHl1wX1xyqed9fjiDny8Ok+/m4oWMKWYOu47Irfh9RjdaHGk
I/DVMbRCeNtIz/d7ZvwU+93UthFxNn8ZJrc52QEEoQXTZEt2YK9G5hBiahouOzv+
lEIYeva/p5D8QX1dXavTdmqsSiKhVzgsgdfwXU1QttWOz96Ya4gy5uR/Annzc9Ia
oqPMBpiqq7HzLtPSJ5fcEdr8kqFWd0qSdoKiQRqIymxZMr40t9870C2D5qqjNbn2
CLmZOMNuiCdGxNIYwCYa7C8BTNhU3nGr44PVyJI9ukKGGg5HVttC4zdA3Owujoez
mhxHREztO4U4CoVpiJGP0k+JibPI2umZEGpDdjvht9MpgEP7qlQXnPaehQKx05wT
mRQX0v3VVDe2zCn8tYMQ4WBlm3SSNv7mtUFiaxNViveS//1GX0nLRZRyrQVRuyh5
eUrrnhTgDzOso0CX9og2FziPXM+8PqpFMYB4uIHzpKO7NQuZrVfqlZuzXZTh2FrB
m984ZFnVxpQJ0wMPQWHRSGgXxuv9zrM0rm5YqaYlcCITiE8wo3OoEOghsm+L++dG
y19P8YkvTot4piFVy9jXkfTGCDR1TJZul8luoSHMUZqXPwC7OGa/nyicrDLGXNtJ
uh2NIHhDz0kZDV+SbjEhumiwNeqCOB5JkC42sx83s2cUTU79BCwZbva6TjJQzUwT
f++3nlMPemKTIdMCiGyk3wxYYY1s7UI5BIKwjfNor478roNE7Sv1LcyxEGujWYlm
iKfOr4HrsWh00B4GY3+nbxR7BAn9vJrKNMMvky/n6a2tLD5Op3dWgxkMQ6u/Fg2r
8pGHLivZF7hxS9JfKVrbyDfTxTXLhSPS/xBAbKaG1nG69mDj4WTY8tYaOvmG/Djf
h9KbXly7ko9JEoBaIvrvrmuIMsf0lp1bIW1i4Z0GUxMiY0zqQHoDGQJ2ZQ+PCZtM
NeA9U23s1aomkAdXlqGCjfOFAld0KQyaVHUvRJHpmsZZu3Zm5kgXvC4Ptphp5wRO
kFcJJcNLkSnXvp6U26ksSLNrAUoN5yvjnVPJsmKyK70uJxeYY0mDJZTKwFYxEte2
Kifp4KZy7Kvof1iwpTtXtd28FaT1e+l1knNwbxvnR+gicE23dUegXYhFkvWAh2RY
JweTPTe6uLAu326lvdKsMMWhzf9iE8w1d8xjgeqWP8qFSftK7Fdxbqv5oyEGbOr6
x0eU2l3cI3HRcll/LU1gpWvdnzaMAYuDhD/4/Octsy5ZLQsR+FlDp9GBjTSc/XLY
rCKiBj+aOmreqT3b2y2rk4UsAbyVsR3UKAtjJ7EllOHAYQet/kHDWYwzOO7WXrqX
d7a5vOHnCu65GXMvsi+L42P6hjCzxdKKfTcLJqNfwVq9PapcQV3TjniNIQk/ZYUD
Kdsrj3cQpx+cRhkFaAi9MHvBNd+1m7ZUDjPx0Bzu1HfJOkKzcV2Asgy4/pd0DAZb
VEX05sw5CwEBcbJKWuyx53wXw0KYjawnUsFuwEaxMcXgda2gPkp4Y+/e3WZ2Jb+E
1y7XyF7k7N9rtH/b75S++sJZDkof8n69Pf1FmHDHtl96nuhz/ztsol7zQpqjIKma
2fa/0alCk6DJcGvlnh/qZt/zDt3VSWoMm2BYIVyzHduHTnU8EkO5kLZ6cjKbLLNU
hZd620NYYkvFkG/juFhayPA39gWrx1uw5nmCpoj88ME9RUjB01m+uWWneRyysDWo
Ncozi9LddTiiBkN1nDeBgEM/AVFQHxzUq8NjUUD/j4HJbM1RIjc63Vj4K9eh3E0h
aSyKdL3BBCp0x/qJuBOPAuuXxVBrUTpJbTvpSbZ6Wq5fDcjTAlNRklM+T66Y1OZ8
7bsbz8U1nmiUzZ1qUEqO10QK4G4TE0FSbIittcCyx0zh8Z/I2iFZ0hUKRgwpJHEK
V2hay5E8fmWkvTiQcW9skzWNl0h1giTIZOaod/3biMNGNGgYRJYwFphsXEWrJLe0
zGdiC3U7/nfQZLoEA0rwO9cjKrfCxv9DC+qYgEsEOAeDUqqbZm0uQVBMW8mvg9I9
zROTQAcrfBRaTnOTIwbs+8IIaMB/wnjDlvmg+KghEbvmELXDXiU8+Uo9ofqdMT73
47hiFjSbdDge5MaaiCSVVQr3ZfmO3s0rDxp4Azoe6r+LWKqWyJewLJ6oFbmMxPJL
UHWaFRvmPJuHYexn0V/KtYBp64xhvp3zfPO9dc/Dh3L0aiKRRcFvrSyHVMfYMEw5
4TB8VYJDsPhLfzLQjRCIoBsG5sx0ih/QmMG+3YN+XdiC/Kgw6eI+4gZi5+kHxted
drW+9d9QtYE33+h9VQJ1NvxyEfzfmJEDHyayokb5YuexuacZIlQgnxLYZ++tthd1
6f6hx6fSkOtJ90IYXIWAC+aHziIbr/2wEUX8vMr7cjCAX+UiYSnvnqfE6gTOyhw3
NNxG1KOYgzCnV7xhKhx1Mn0iZnxZkZyfXOBWiM+fqtAsZLcdZckvx2Q7v6vWYGTE
SqN7o+OsG0KwJr+eRSvM0rI+L4ttbWwMjg/jzTlg6ChyLqofa+azfiVIFT9qAo6A
b/mL6+QxOtcMigJRIUcbLjHEGI+IZYutOhjtlRr52Kr4/brBXH/EsILHA8fq9sIt
q7xIuv4YTYKZ/EcGnUKzDiCPGaGg645XC7zaAOD2gMsfEUSCRZFhwYkgQpOsufdn
+qW84020Zr0aIwX8l9E73D/SID7mBR+DW6grg10HkK2ym90+0YoPlJhaY0YvxBLO
1uTitXe64uvCtehOCGcDgiqk1QfW6j45I+/Z4EH0++pMG+qhlH8aWvrVqBP4dA3D
B/KOwOSp/DvmMwfRndOgDHfMewul1vlUv9YZ7y2jtTtGIOfwU09GET+aC6KwpaSH
cr91HI6XsXSp9DGwF1r71qiy9E4spB/QyXpxmTGOs3ZmZG/g9F6w4S3fSa/rtkOB
8jC7AEHnyllg9S5bVK2cfrnsJd/gY18WErYziUH5Kdml2cYTt2HzPmu4Ocx+qE2v
60/KFV8SOzZIR79aX/GsIj6cnnsByjHsfciA4sQL3R6qpNGMLsqY2O5Uk421SREo
vQU2I+vP4TLYEwlCd8U3bMc1MHgOPZ98xB4k4XJ728ynT4vxBg8+DJ3pgXlgquaX
IE2X3HGiUjtAvZZmhAJmOmjWbOw9x0aW3DZ9fk32N57fGnkE0vOvmcc1c3XAkcoH
ahGX8PYcAURHEXU85RJ05ZBc5mhaBXK5FetJ2rU8rWPCWYwcXSsXklkQNrbDut1+
5MYC5G9zElKDlR1540LK3VTN3srnNVvDP7Lb9kqxKRnpqnPYcehwhiEzCXG54n/Z
BKDGLJyFMq3uGeRWYr732m6aYD6MKLbDJfr3zjOxSusNdfzHci1PqcIH917Jsxhg
EZxQLBBPgE0QrGskXpN6gpbNjtO7KPTlDr+Ev6BJQOLYHlr38A/0zUhZCPemzTM4
az8Ye8t1eGaG26K6I0r96sJvPhk0MvEO+jJ+DhPPZnWpqRvlG0Jt5zAmzj4K++L5
m9PKZQ7Gh8wzFIBp7AysAaKileOtjet0gdX2gvoz93YQGe0RHOWhKHKJQQonWQkQ
Q8dGUe0jOK7xleHROG8yVBQ4FaExjJ9jZHEtd4gkbb5iomJx6pqifL4+cbPrZLNF
Svp5tSZdB+Pyk7CAHY+BcOxte3ZBWoW2Yc6ylC6gV6imWsUSvqkMfEBD8ITGpBI8
Nn5wy1wxPXVf+phH3OkYAMIXF0NZZ8VRBhQjelAKgaF/8QW7wFiphPW6/u9myz7o
6Z9yDuZtTcIyRaJAjM+pDVi0HFEmr7YIVGVeujFANu38l3eFlXyOtYVCxTPBs0i3
TGTRjLHkd6lUh5dfsLSH6tlaNwEG6I1yG6peOAToIxC7Z4Vh0nAqytAsBpmesuBh
Fp1B8WO5pwmt56dQAKo9pYHOCRT1EVIBkfM7KCg/5LnFSqQAr6NrE0PMp1OSRAeW
zaDNf+xnAtyu8iXsq8Ol7OQPSWVntyIiGR0vwiti5tgrDFH65WFWc7lPVl9jVKjZ
VdUeqPBcAZfc4vw/zdoZxA+1MO9DhoQ9yZEjHCbA34jpZSAMm7V7HUZbs13a4va7
nXYjHYAFmfsb5KOPDLwTKWrwCyxGWjRqOrJUECGoUItftdlClXkxvb/5ajLOb6GM
Ys9scQUHF6oZ6teDRa5meIx+NyeCjeolDU8NkCbjgg+13T1oe2VYEaI3WdvZaup1
p5YfGtFc691TEZCxDVc8ufhPa/SQf0fQNTHCKy9ZsvHgLBhGuO7xVSGOysjR8X+B
HgOVpzpI8UzIVkWFXfZz0HxNY/10/fn9UABKEglzx9Htxf9R2KUKX7ZlC8QZgPm/
P+paQq0CBxD58cM6kJVpeUdpIwHOIX3QF73xzfAEXdcQsQ9s9aesIcz1ZSS+fHfx
AOWKTjIF2Yf2UxTSXQy+OlbIL9yg4hithvHgpbIH/La3HOc9LT4J3F9V4vi79B/i
WhfrQ3j5cXWzPsGftqcrqbHDU1mc58ByRe3vx1cPyHd806K5To3r+JbSJdiEv4je
GzSJfyqtjREWckZYs1+4WehNp8x8rD4KxNnv8SWRSMin0OrMBoA3mHeHjQaZdWOv
KKB5WXmjRdpzGU6fXoFN2bNNo0hvORhACY1MA++s82VYEQNGF/jzjzpaqVVWoEAI
reINC+L+oAxNQ1wyuVbQABcPJYht8DQo/Ccuhah4o4y5gq7WWqyV76NZJ56E/uAd
78J2uen0giQioI+USzu6XmJURiw6ZOGJ+nDUDM2CCZoOJdOUFRMmOIx7Ta3vFTLW
6lvo9gjHyvqfnQiSITIAj/CQiBhXf5jrTdS3ojhqdTrH7FqOhcn0op6gegwLKMdr
6OVbKUV7Butiww6iItNRlHJ2XPiUC5trtYg7+X4GA2LtwGhekXAN0RF8IlfCF7Wd
tPjA3iIW+mc8HngA5YK0p5M8AXRI9Z/FbISJ7sEqwTWPs1TGWiXN1DvhMakPgRnC
gw6xchwGOdjXBqFu19+W9NJOsn6kp8jJwbEBhXIeuOsfnECL59HFuB7Wc0ruRqPy
7SE6kYcxPqEMjMkR6+5lu8k1X4T3AjhYFrftCrg85p9rvcEPsTug2zivBwn/LEog
Qfa9iQrzd4Yzn7F3Z5y0FYfy/i+vZvCoqEHsSmgx+Bwn+PQtmP8TXcxuafyfolFX
yND+1Lakov3gWFVkTLAd/yOmR1A1HSiae/6NfIcXNb/n9z8dtO0gJYBzNhIdnl+M
5ruE4AEctDnR7+JU2JoEXlYAoaYonyPbhVHLYkix2YhjPTS2Z7IpsPAjU8pvAdiU
yijZEvwxdarADWd0JkwIdAgeA6xh+ucb/o8hoFutJ8a1UGY2H7b4t7DnvkwrQO0S
8umHJKEypBJL6E3TVqupW5qkywCBSyT99aNjd7qM+UkiIejG1ajV/dafxpHRxwaD
YeuhgOJSP8UuuD/Fo5f8mlmaQMrPkastVSB+fNmcqbEwOIBbOVeY/3n059moXHDg
TD5e5WNW/Xp5FiH0TSg3vNAlHZghWgRdCEMtuwyiabH6zU11wO/HY2MyykaTSjMQ
v0ytjVf9MGVNi4Lx3z7H6UnembOh1JRrETo9HmWWEn8+Htpg1Ef53ImQhj9yD3yb
OJKBX4tu7czaDLGgKz6jURzYCGew11bEQ1VywMjM1GjNmgXYz37bzyzLAAYCjMX0
SwbfZ/AwDJW+Mh2vhsYBGAfwKce4H/axozIZyhjbn+luwyIUb+jDtpBUJSXST1Nv
Z7HXzRpFTO69gVOalrU3tLEY6SVALCutOI0xrwKUO2jdcD7dAWGMyram/7LXe2LV
uu5UdoEHuPHvXK0tUS6ReraQukTwk0tVRW7NhQq5R7pZO8/4cPiFtqRlAVCXJ28o
CPqQyzjB95xYtXTPwkM7vwcO5YubEDCBvXNwsQc0fayFib5O2+JvjIVHcEzqg5Gv
t6S9Equ151EGhE9SI98v2gJ9o+X/ngPzzXOn5p1osm5DJsbRKEIhZnp2t1BLlPCL
U8Lis93HWrUxKg1qaYK+NoivRjPmRxkj7Z5vqKi/vOirBk6S0N578O6959KsADny
/jGB5+K9CoGbR7eF5IMZJ0n6zzCQtsrCxw0wqEbl/bdhCg3iAnFZnuX3tVAGphNS
D1zp+MK0N3Tz9e+XIPqqeVTwHSSfss1CjPdEEqECahDQhsAbm182XCiIWYKqiwm+
sdmC8Mf1Mq3OCvMxgPa2QtmrGkzC2QWOW79Dv39s2TE63S/MqnQBdVuqK5ILOITt
cACNT5Op6OJcRuQlS7NuGUsZdk+M5ZoalIPkuDkzbY0iiUK5/na5Oq332lXnS+Gv
okgdt5y2OFGCz/jWZpwKV5pSrQWR6QAWM/sQii5qM5shK5yak2JkE/GZaM2jIcuY
t9RGtZ27iNmHJO2wwS423E38hg4GTc4bxiGfhx6apQ1jsFPaMH4q5DnT/IiTb5sH
hKxmbt8IfZ9i2mVBO58PBjyAseGiM68VHqqVOzTuoEWiCYEfTHyI0NBW3OkfBuxX
F+wIc5HgjT+btwBYrbZ8UQXNRPzqUkXrEkPnUMXXKkQiyR6crf0wVZ/sUf4uBCaC
R5RTw8r+6QlnHNKBwpCL8WrS8iwVV1gEQ9SPBXs34ObJifXmvUJ7HvMoU31T/jtf
TlLRhJPNFB4zLT1Zn3ZWrL3v8reakSku4NCvRowOVrZdLrXC4TmK+lXYbiD0GLeP
/jzFtUicDRIlrwAph8UH0Rp007o0knObspaRG9c4YQPsiRmx5/6tWPBn8hmhpFsz
AXWTJxp7IuwZgcYwAJOoaokvtkg2KgvbtMN6S71E0UApJhOcQk0M5brTnokSmnZ3
fzbSu2iMj09jYhR9RNBALXy9S+uit23Xegy8CKrgK9KPXGx/RNZPZCqDm/2BLIxM
Shbwje9zIN86TjShgAWt5XRVPq9lA2Ajoqj5ZPuKiPrz2hetPrx1cSutwAj0KpPa
vKV7Lzxv5GX7+indZuudaOT4OfeySNU3WQWNi+elxUiA+0j0odaIXJL8G1ZEpZ8D
39TC6+NAoK1sOIY/Tj5xLemb780svmfJ1qf1KuDo9C3WX5+dHImA8frOTuHGWW8B
mTEoc6nAkO+lvqyWONyCp01P3J9eJuVuGoWz2+lRxvSodstGAHfUOB+z16aP7sNx
fBje8HmaxCH+1/OHzIH1mN8+N3ZkouLmyvVbspp53Z2vSOrJi+2UgeIEtx5Jh1sO
Doncik6bD5blXU4uaj0ERowxOoMQZ9gPD1QT/s2ZqzukMiU4fzccoC+T3di8bgg+
VuI48at8OVgCzvsLuaZtc+YlaNt0RGKKTHBzUuam4fEt85uJzpFC7Ywe9rPkZNx4
N5veGnXJrhNmlj1ms9fj6agDkK93u7+eP3AdFZR57vk4aAEw9ZiC5WZhzCSHpHUL
P/MwP9EcTyqXY+3OHT/6qKhx9Yk2T521pqt62KzedQ9vMdptAP6w0NF9kRv+028U
7w9FAxKRLN4UcZTceAvFCta2V6kzvdMVQc3DfwWUA6ytUgkO4KJM8bemL104gMRV
3CwXU+iO18CVRZUKrzQDEyQCxaMvwKaH8MVfh8sqJc1BPsFIwfD5tx61ZNqHpn4s
pMsawxRi8fjG1EIIInuYqOPnGjVoFlxrIuMw3+2w3bHIPc2D3uLnVrWHucoBJxn8
LUpxJcdlex92A/EMRP1o4yMswdB/iTm12ZVsgdVb8Dh6l1Wif23GEZm4YQxNqmun
McfZDLTo94n7iNY8fnOpVuBATpxaW9HJKx382mEbpgsmEM6djpJQ2g9d2VSVegRX
wRgsdZk82mosxsSNDPYwXeZsVsXGFztU554RJ6bNTpMWjrc4HlMGBF6l1XWxgT8V
zgR1+k8D+YYxW1l5qzuCdn3ztf8G2e9oDvmTOkI3PSVZGnFER8KqJWkYxQx1EtvB
8PjwHv6DceIUwYe8u5kQ42nIprlfn/jX4fqTwjMKbAAWB8P2bwKsRZ3hVdhvXlgb
vq4gfMeLhngu0i7UqHjPMUVFspH2tCMi0LtlRXWJnUf0aKcxTHwmXyxaL6iXtZRZ
8xgKTC01mrXvZZl/Dpyh/7Za+I98dTQN8R0umAWt/G/r9mN9CLnZtKSCnpuUmIgi
9DGfwuCKUc1rR8eWs1uZKJQ88XStk8C05PZ7zTabgBfmmNAWYQIlfX5Nuu6WIKjo
NMOERbxMYfSrDELBEHc6MU8StDCJ+ia7aICHpdyRmoYQY+++Xk6MLv5zM8zc1t1F
LXbuDdIibMc5ryIBB40vydv9qa2yOAxbUlhi0eS1XbDHjBqLIoRtbVtuxecM/ozy
Dz8ozcIXkk0U+MFX5/xpsnXC2djc2LJEa3yrDdI6SA56MoNhIdzvTezH1T7MmW2+
AG8M1irsOTFBY1cTdmCcQSVTXdvptJjGNOT3sSWxu0ByKNqq948Qh1vJSR7AhBBD
qhs0Y982P54ssexthWYN3H1uSgRxsM0Rxja4EgcY4f4+Z3f60bSKaLEz8Grp29BV
3ypz2osmoOG7YPf/rkLA4iLsQNae+Qp6zjhVlIblYsFrGM+ptTf98aFBIQh80OL+
Az3eVoSH4XX0aODDABwrWK+OP+VZOH8lu8xQQQo0C3z/cFG2uxyNzERx0LOkPFk6
+Q45agegmp6qNg6lqSDvR/+hUIskXw4owVqbLoGWvmaYQQO83ps0lGiwaaqhPptB
7kswWu3ufpyGt8p4zduJMoWfCAFl4Komj+NZvNfdUlPAJ9QlU19go6Zp7JeDP1qL
sZzamoxdVkpU7WAv6U3svg87yOKFkjdXXtXZtF6mCc7OoH1uf2sQOme+DKrCYlSP
OlTPI0Y+og7zIg4V18O8TFgcf8vrvyj7iQB7mLmvcE5vhiWBexjpDY9NyLyJrncZ
UIhuHkP9DvNBwmv+W+D8H+mgnY6QeReHgILXT94KZl/pNNlyyVuI+T1fFYOJb+m0
VV06Pse29xn6YTEqLJdp3YIob18Pq8p8ZC5PHvToKe1Teq55q/ux0df/s31bK0D0
DBMla8OIMfz1TRgcCnZORHAvLjsI7LbUYDkwsijktZ9F5jjI5MgPCUizwRhaW8/4
Mdms5AvWRCuZnWwC5jwIpDLqrh/l2zUGYcxHEAF7RG6JWUBBYoZeYQZn7C1YjOp5
sF0LowwqvxnSxx2awAMO7SBN+k62c5gG9Nh2cXOAGrPjHR1l3Xwdf+fXc/O8J01i
9+kwdA5hW4tWActr+Mefikcy9dtZEUGp0O7DhIHxcZ1lbkImrLYb9Gtxap3PtxI5
lIgt9sZaFEpBChV6UjHgeqVdu0UwvI3L0ECawTRz5xDF0bQ67IiLTuo4pX3WoPQp
SWoPcowGQ0LScZMUlQ5CzV5QCAz2VIK75ZofPoVZdvG+q8/OmrzdRoa+NiJNOj+m
1F3D2S6FFVuuNwE5OUz7w6LwzSsNScR3iBR3LVizSVCTvW1b9CIFHPZZSXn0YsNa
AtaKj42fXfi3xZYs3PiXNfADwPFEGslRLe3xmoPu8Fvh95TCiB+Bx2sIuxpPhqGm
Nt9YWbN29FzQSuPqrkLnPLXhr+/sCSBrEl0i8PThJIVLjjoeTA1S1XKWYvEjUqSc
1AruTQaWoJYem/CDtpdgJOGO1Hk0PwQ9SQUb/jDEKVh6q1ftklO/4RfPxdpNbkzm
DxsePshDR4HI8FN3fq6497xEKTskxVasR1vk5kD0B2fszJ+vfKHfwx1kQIgDbv8i
rmL9hwlngCf500hMt3MIwvKrWAcdvKxbk4QKorZPf6gBZigUpJvbcWoKEv+sd97n
zPmkRmrKEZUgZ5WL2V1lQhVuJMApSERPZ4AcZqRIpZMK5IwJOyZde1ZD5u9IPHcB
2YEQ4W7ooQ/VL0skPcEnDVBarIhYtaLi06Aez1VXRn0/1aMS1ZcYneGh1Cm003VG
9LMVB0yDY8ufz9Tj/UEGsJ+rMFwGXYSC4iRhyZ9OCQxDqNWvUjUHRzQkNIYoQIVW
OMQQ0nfHasIy2hBx6st9o4AoOQJAmwZYk0m9zi2KKg8Ysdtae5tsKRCnrZOBjjA0
czhGNbhtNJxg0cHemBep2+GXhuecZP0UeESmcS5h+pBgJaSYPNrmB5bvQ8RtdoES
g86TUiqbMj9FPu7IlnjbSehOnIPfZay1swpjMzRhUIoK78i+ilQytgYTjMWZ+/ez
OYaO04uEjVQcE10y+NIZt7D+wlDgorgoa5+xzpXH96kkJrp5C7wKE4DSF/8rOwab
1MFf3SqQaxunvXXQsfD5F9N+OSpPYg+mjnjwYHcn+T4+f20oo2SQ00Di1vneTVkk
+NYeUY3Ewo73mKV9LFbHbP4ZDy/2chSQUfr/PR3GDN5zvF6G8BHap4eZ9h2A4Z+N
0tVxfsqzqw+OkUhJeuX/yA5fVNbEywmT1U8OqQlbnJu4f1nryWKacche10y3uZQW
EJsfc5zvFVOdM8zK+MAwkrgiFTnWfls9K0svUJkkZNeBrdfuTT3jXeoLT4/h5PoH
apUIAlqliI2Z16OHXXDfab7wOeeKbjNOeS0bE38etsfZM/XDzDRO8wYUxGZhprtS
BgIEyFiy+uoJw0CGTIVdcsyfpOrz6EOp8QINipGvOFRda2CFsoxhZfrhi/Kivf2G
DNsiIEo7au1XjuLVErguOzHr2s+dRti6HulXPdnUfVCC8yxEKlgcWMUpgIaCWPEe
ZkktBxmwQGmqV3Rq5Cj4RFHN7IXAO5pIU+qgfC9RXVOtaUzGtPvdqme6pUU4dEx4
EUzWyux4vxL+Y0z3oeukwY6/fSLRpQFTNhqKYgHA1xqclxuapk+s1/dCX5HbSoK6
3hwo7U5HW11Wvzi8ENyow/T/cHSECfLLWhGMFW31mDi+wf5Ci9kgspHaKh8wJQ81
tuoYMpZhZXn06muEycy/PfE19urXe5YGuyK33ka/F8yRmQ91Bkf7rIK0IQwrRPnO
aLkilr5myRzcHdzrsmBKHK2fbERJlRfi1/bTeLn9UY5BqSONsQjeGMqhQI/E26rq
IzAdbvA53gDz4POwAJZWQSYNvnG8EXopTRerz4JEYqWfP9qQb6/2qwwPaVaE97zI
R6Qq7m4CN9kbHL+M6+vZXIA/WEdDbFYJXIqPI4SCUmiKtsou8E71oJZvP3QdVRb/
vjYD7C1hVmIYHxU8PeXU5snItUh5Xyjwp/ZeUYN/1gaccLBFG8XN/w3xoKm+or++
ZhYgf3Qd063YVMAhaVdZeLPdDFmDbQvjhYaxTASKXHhSCB+IrEC41njGi9X8Y4If
U8O9p1ZSqRgZ+mIMcAXF3XwgFw7qjbpjmwM4M4RoaOxc6VfCYGvCj9FwQAAx98Qw
ux/i4KuATacgrNLU7K8iAIyjmvnWPJC5y5VCXEH3juy9hx4mO/3dx4fZqP24TGpb
m+QcVdVqMpvYPCR/SLTunUz15qeEUV2tjT6HrcmC4NoLP7pEBODbfBOhXBIDh6Vi
My5Ujyn3qDPzJEV/pcOtmKX1cHWv7nE5yPhHcxhJP837GGKZQPYBSyIQoDcfqjQU
9tBKie+qLgQ3AADF5AjHD34i9vXFkOH+Zp6ySeruTSSPNNysFtkrx+ytZAYrh2PC
McHdUSKfUnKQM7FloM0WbJynWGl/wk05zGCZMuwP0VZNIEB5T1dUbRYguVRWrf7O
/PaQDkffohMeyMWKKocr4aghNIfEOS/NOxB09suHo1l1+VddF/yNeTLM1Y1GYfCM
TWwXb+dkvHApK35MrDkH10sVx23t294NdR+YDi71ecXXR8T9NhsDBrGGNnPmYnM3
CUN6HIhglwoEYTRg67khgb9uWErknuURVV9BDFVdjHPZ9FMIV+IIpCWj3nLYpiP4
2Iif0KqNuoT8Jqoqmf354b+iNtDWoWobcpAtxQ2XcGFx3iQHlbnCb5M0g2Fz1hKg
YeerFo0LAJG/7+m0ccxTPKiTPIjx/Fc5JUJaVDc4kB+u99QJAPoQr0Mw726Cokap
F5pzDN4xGiaOnT3WmDXRvFaFUXG2uLz2/xBhJQs/TPcZmsEmrLdK8N8zuZuGrAT/
IQ01ZoIhEXHCEL4KEqDXJ/yIZjOxDM24R6D0U/YiWXPlpXYPl5GsMPLr5aLB6Uwz
fIsm4oD2jLVKCvkxiI7gp/5oinWUnssY01eLdNRhnt73pELYig3t6lOSXZCwpD4m
RU1txMIb5Ea4OaS9pkyUEoxRfkKdrvg3V6O8ygdadblbtlRs8Jmetk8nGohBm7MG
IWTwLQw3SQsPeUm5JQc93ZwfCPPbFz4yH4GVtGBnscZGctwzyDu7Ch4+dLybxpKg
JMQm5VkGA3k10DuULsoLboAjvzjAJfA8zCbetMYxya2gb4HLPRw8DSJI4hk6VtdS
/BuM4LZNhUGWwBjK+cOUGww/j8m2wnl+rD3hOUTMbHah31bU5U2NhSplxenXLa/9
7pz02/Z09xF225TvdhgF61dLbo0fCVzFZJLVvXwBQDQcLe4rf2l4JJvLGTrv2kfX
GoePceG5S74R/vcG9lq4HKSzQjBBEAnsCN3X2rZMSas95Nch57PT1Ol8RnOG4Ajr
dFjV3e9fy+556FXvtMESJQX3RsxYAPcLPpX+WzMQyKenan5KFPAUmBX1eBPTuCX+
tfxohDMKBv5aBMx8rMC8vQZOtjLlN5OPwiorsxV5H2a3xgPb0JsOHNB0COkciibK
e6yAbc2JRiovQXwdd8OqhQWVVR+FbRIhCpgFhrnR/gNwciaBkGXv9ZhGTMwK+zEX
oXKZaHa56vd2u+EqseehFKTdtWR+xxqIwFw2DBhUIqbniUqaiYEgXny+p4TQAMxN
ESbgoGxh39ZmHgU/FPxsXChu/2x39VdZbVhS3r2icdyc0wNg3QJOPOklr/ZFt2Qy
RTIWgxfMPbHTe4nK76Z18/4SAMQ6mlBplkS/MmrYsDAsMREPzl1q5mQ8EFTasZVl
HPERhTavt31wcwcD16EOJaSdemN5F+JZs25k2MBHygv8WebVDQbPrzk+HKixKIZr
o5BuSadQl99OJ7ppgIRf0tFCO7EyIKRAB7YsXu36hxehAPDXM1Yl+TOo5WwVooTH
qpESROVoWFt3wJUR1nWhHjyJvVKKB6P2qEijiItwCxEPgpg8vEJE1GQUXHkbUb9d
nMHS0LndQMRKPPk/BD9w0jQzjRm15b0bKHvaDhltRVFQgJlW9CfXB8v+lSoj/I0M
FiGNUyeDg9KPsnlDNgSlzUGKilhpMjmIG5L5GVVacnDrIhda+au8yAVfp02ropox
k/DC4E8VTkK4tkuZYRiGETxNtUSVBhIxOLAc6mxdDpYmTpEzIpdMak5pz+S3qLov
aoMhs+alBEsiVfyVlmZD6vPB0C7GEpLSBf5V3z6s67YMJHBwGMBrggPcBrck4oAr
XbiDHIuQRWO7sDysAooxyzyWh2GiqCaUNwt6P5aO1R/sAEA3rifEy6+zeZCQQLXA
UCrh16dxW6iXE+VJPwBH0kbo8khNFvJD5thmVmB+t6xBU7VU2M3OeRQxLdsRaTXk
M1OKTWZPooLJ4N1QyoQumo0hqLNx0/rPv3Yf/4LVPMNiPoNh364xIfY6T8PMGjWP
hulCgXYw1OsrKWH08s+T6oneIMMdLm8HKXr0LGlWrNZCshmrqcKoY1M+M6+X9q5a
Buwo5/dUkvI9+S3XHfukReAS8mQubj1l5Xkiu2Ta6OZj/XIReippneywnd2BS2d2
OvJPG6U3+qtA5tgarU7OB+JXYBVZ0lvEtGz2Pwq94hz4U0CRUK5i2qbu62WJIg5G
6QoVJmbrbxmUsX/2Oc3O1cAPXEfWHFU8sCUurYFjq78kI+KG2hTL5e4DxhZ7dbsb
TIZPyC+jViZQRJelgSczMgaMZV9Tg8VhZODgXKs2wbzsXgF7o1ssXfmob0jbsSV8
bCiVKAHAkH9hx3ljbYfjDLuV5kR/18ZVgN/kaJHMQ0wGBagwhl+k4KmzeSh6Gnal
fgrlyLYPigG398fB7+ZhSYmvUHgbo7WNFoiYxPJml2/z/dI4hpwmwP/12KWFJi3p
xTqzr1PvcIJah/lCTO9zwvlftbdX4Wnp3ZBL9VvQ1VjDdhgpYqmQTd3mR08EAGJs
dakjFj6cgYJKczR8sXSwIlOx8q+zVjKvRupNejJGrF9mPeYSkIY3qQBl2e+3Za6a
2AdVHJHjqSjpNMM0AZmUR9l3etuFayxgfcWfGqoTlvFwBrc92BRzXnasSsk4dCkY
jBcfrpUxmxwnWjSAjO5qZCKENmC+CRH4P5NXnSmvTXZtHIoZNsPKAuWgOWIMh72z
N2s3vr8VG64Vwo53rr76hRNd0glDSOs8WNoJiRZkSAPVCQWGzm+iJ9OeaA5gB9a5
EetlHbQXSYbk+8SbTSULbsYl8Icuo/LeIFRTWvlRdjLFvH3v11iUlIuTiPkvYFLC
nvghaDTy7fq9SUwmF1tXD4DKvhyF1lwffCh9bpXGdJhBSVzeH7l+xONX/Wdox/hQ
B2xZOjvrVpsd9QGiiBOWSM5J2Blm6WdQsDS4tVvJDlxZI9u1hZwPE8A9eTJYHSbh
wok+i1RRljZsYXj1D18rGLZFrmRTiEnH1EdmGKfjp8tMnYh97/DkOTqBYl3k8MHN
OZ6FnJkhyaBP4jBMPHwDIF2nUeJvlLKpNsE+kJnvaPbO49qGG5cgWJ+wcA/ZyzDO
sFHWIAjn3dyHzNmmYixOsaHJntvQqD+E6c+3aGHED+0AMkg0mfGlhyKATaoZ3P6B
JZNOMI4K+JYE3+qreVmqr+bkprem2+ofaCZdoGfKVWjSMX9jIs4D5gYoLsTQUsNN
kFYIy8I028kzEPwnuQL+48NMZeEjd1iYDgY/gobncjRpbe+pmDqZkrkzzmC9vl6j
QZ/5Oofn+HQ6HeZ9fbGdJucI4lBA48hIq29M1/oy4evLY62aPB2xSpPbuLP5fRZG
arTW6YooJQhDzD89fTqGMrhKZvyKoCZZQoEuaweiYRYWPInvANVxSRLX4ea6NbXs
RxE6+u/M4AIv6EZ7f4h6cemhRosdvF94s4d/Lu7uqMEr2FNX0lPDLCHR3xkf6lyf
3J9NrNkoqQndBme7ym8aBA8L/Sxw0GAjMdoNP+52yoB4NiD4eCub5hI5JmCtp6Gf
cjQ03JkRRxIklri7GNtORQhWiVMHQhF1OV5VNlkxIX+DUYU6xuANF+hB4QCVX3dA
/XFQ5taQHH90ojztFj0waxMF/ZJvRIyoj9mkGpwF9Re/V/eAfHFnX1hcAu7OMxJn
XwYUyNyHManaWkKBM2V6Xj+EtesXA9+lFEmIn2/K9U2midrDf0O12TihqTzbP897
g9ELcsfKSnFikh7MvGq2ODMkukluXvDYsHg3PT7Qcqlc8Ywup16N8HsdDSYj1UzF
wn7GbNZb/znmabawOwRocKU/CD/NGJvk1dzovV0H+S1tKP9wm5HkVHRulbzqNNOw
HAwlE/vk0bdwuVJ8DNu6ac2uHfdotygzC076DYwtGoBwTp8rcjK1XeJefxAXFmC9
3z9tit+bJoQFgLzg+pByLzS3j5w1csJOr2nYqG/rwt4KLkG/DZGZ1LtiJP29WUG5
JdYx/2GG9nU+Noon6lX5kTo5S06zqKtMOE3lxMOWWD7xbfwJ+cD6L02p/nnuU83Q
EjZTcYyiZKobRIzSm9r2HSgiE92d3PVB5hxNykE56uk0Nh/bXJKjaCdh2NTYKDfv
mU6vXFm2znEJ9xyrKFNWnuC/EBvdW4ZX1QVUTVTzxWg656RBG4StIzQd+ahuNc8k
9RVM1asfRin9nv6twSCztPXMqcSDZ0mlpJGoRdOXNgTOQUrMWhzd4nqZQhRM/6LA
94nG3dO6k+PYo7kGc8+vreqNBugxhg0gAI3S4kAQ3cL5OSGYvsA450IOBL+QCT1q
3uUnD3/6d1ueBwj3+og8vkJLF7U5nqepJ4WAtKOQ9KUUmRVNPsLGzks27P7MPOkb
hSETTXtAUVGqEQtyz3nNgTLW3fGtUG4cmjP83dqeqtDEGK15xL8Vht+9Pi3lAzwN
/6guV5nZn+jDVYhckrja7PT6TeXcUg1jAoWrWYOJQ5enknEzKCcEvZcmGu8HuiEQ
WTuurp4r8sJ4lVe939OVL+QfD/OFT/4SHQsDjDQtH81tfUkYFyuJjVZdwxeHG7aq
0ijt53GqE1bNWX5gjEXvg7aL7bUH675gsaiOX6S3AieIDSJ4XFNM46+HJXjORK5B
/D4GXU/q1N/p3Xv+rzmKOTKKPanM0pHcb3GiUhkGQuAZUL8RezXim4NoHjTCBtMC
S4sqJveEGleQd68aR7wG9xQNwp9msNe0XXDslnXTZc0/OFiMlDz2hfejlcI5U3lp
WvyxfQ7OJCHxtOvuHqoEYM+RJdKWXXDPPHR5ro9q/EVKESa+3pxGnhh8KQ5dAEXE
OwTNRgWDc0S7D7lo1d61A9mf9SShMDtm2lnPYCxayFAV6KlGiQR8mpg9N+/NsrAl
/HCPD/NxJz5mneHyGj0O/F858G0EnWeBS2sCAFGcAmFi7dW8BQsi5TXqPLUfbL3C
F2KrUDxC11zFeTopDsBANtagH2Wx5Ye2HufwAa2KfhQPjkATFVp9oiJBXbpmaRKr
49cyHaQSGNcD14+Or1iAJkpajfNeeMnCespee5hEOOyjhHqPXlToIM9iA4s7lbGC
85EOINDVcX0XHxg0ROj7o8dHVQx8OfSqE9+AVGh3KXtBiDMlP3iv0viAARJjCfQG
9MGgCtHkc+fKygBPt5qCmzn909sgWDOqlfqr7DjqdE5N2BXqma32EU3bVPTl5RZy
t8rzxpMWMAevV6NCoHMTCTajCHpLc+/c7WC2hV+a2LwApWHotRouFGYOl0DyRJFE
CuoUdpxIQE1gY6vSX4mRnbZHKsN89AyWgb75BaUzKvXnhxu990DujVJrJd+terXw
7lc8MFRJqeKJPqe2qc4TmySl/0eQU4PFtBNJvQAnYFom+Zxd4YcixyBCcEkBwHET
ZMrQwSPbiS2t+TE60OmvfOkRtW+Mu15Tl1lyTHLslC+YDYdbrht12cchcgo4c42a
IMZi2jwTSegdWumx9UOY9MK+GwBfonnqI8TNAQpRgHbDlcmo0XZ+1pHRZleH3mIt
3Rgt6PN/NTIhE/l0Pwwd6sgE5rcIuw9zqe3N5N6rbdXTyTdkIBD34OCllUHDNLIf
YM6JbODyOCuyYhavXkxWHdCkoONH5B6+y5F+i4OiAdKsXL5n1ccbAS1N2MbaXFzD
FeCwVUqhUUbuqzQ+gogBijUsUTcl5LaA511jPoFEsNXxRJOwC6Xlovdebk6gCtIA
h69/sFI3UlDuossz6iyTqmZEwtLmeqNYZMJonVs2A0prsXHorKaaA46WME2rZXC7
emcbIjGQE7YASLoSNJID93pI9TtQ/BzXMeo6lQzaxPeb4J4oGle8ZNEm9aMBviP7
3waz7Mhb5MHxH+L7bTRig2qBnR0ihg4nujZwCt9fU2iU5tlO0TY66BBdxFJVwW2a
iNUv0q5uKAr/7CLokxb9YqNln+g1OqnaL1uBeoWNTYMuE8ZYQxawnYoDuIJcLm6s
roeO6CcWFyEERspakszx+yb/aw8MagBrFFPp+RdDCW+6OKxnS0rAN5nd1/UU5Ex/
kHibBfmIODeVSzIn8VDokL1GiTfZqUDMjymtHGYBb35pTuipADF1Zq06HtcNawM0
35jCUY/JeifQmrjyYyDy3pkqbcLtY5MYV2DdkSwXoa9rU1p7nweYIqu8o4yWOrcP
+ptoBFlKMq2xhCf2MbrZLc/TTPe6ZLbUPn4NL+MhsvR5aJ26B+iS+pQ5hO2JijH8
on6Pik542BeRpcBTiNmsc9zMGGotXhjUrk8hjgw48CGfD9i3nz4ZLO6x+l5S8lJn
dhcoMlzHsAIx81hM6WSttQQvfwS869xXW2GWudxNPALTYJMc9gLUJ0k7lMSkw/uo
IS/WAPGdDf+Tf3QFsmwAMy+bvQhyLRN4fMqdCP8YAbev3QzNDJs4fDKZFffhNgKH
UFOVPw4/wzKZpZNZUxLlLL1iK+tV3M0CE0HOIMkJiRNjIjE9zv3tWAbwPKsKl+r+
Z1V46CNzXdPBjdQXi0iqOTuUlo5fh6MKgta39v3lvL+FpHwqhhtYSidJR1EBxKgF
TrT0WVNCgC4NAyInH/FP4NW4yQLg662EtOpdhQiKJ4r8TLTvGsARZfA+UzlVbKMn
qyyBmggMIvp1krVGMbycx6D8HND5jEUViX6RLjdtVc9awnlSxcU8xb6EvI0Jt1Wj
qWJ9/EBlmhFox0goPqCp/h0oBJ7b0Rruy7OglAgjRPDyzGNma+zv5pzoE+Zh0qg8
PIiAjDtKRlfsc9qkqsqwfrbSCCmFvCvgYm9t4CMf6NIFn3FQhH0PcWMTJlm7llN3
nr8e9spXYgZxAQnMdb0p9d/R2uW+BvRUZrAHeRvgjH2ysSDajrG32YineaC07T0G
JOd0WagEHVWkulSUK88mdFIMIzIqEor/I6sym3+jqrz7hJxwjIkuI5OF7Xs1vgz+
ATtuSaZ4F05IpC/w8zvLP+muVW3I515q3oRDmwG/V5wlLieO4azmCjnBaPC2YTyg
70jPkpGGFnh3vUW0GfU3UIKD5pmvLfre+wt/1kak0xb7DFbtUpxeEuEJ2in2PsBj
sTrnuExEDu2QCbnhHhQhiMFOKO6GhmEBsrwBsc8v4Uq8mlFZqgv9baeeMwKLjxyC
VuMRtHq+Pn9Dbajxw1MuMdyeOczVP8A7EiR3tGBs29BwXQn3hLX3OuRkzlIIeCWD
mlu1QjZ1t+SjsfVfLz8uHqCVyLXP8ibGOwzXC0YrL54VOxEmH6cUyZr3nU3AdQ4y
6xOWmBjiE0TZDQI1wMOOXMd641RAJsEqBrOjZCFROXyhLBPGHP5ZBveEIlfOtH0c
QBWJxexRUtu28e5yTwSCwoDaNl0bfBC12rgVqv4FRyreIyYU7O5bG4Na4jC747AZ
Af/ie9SiorJoFwzeJXyB7XFHHyCSS6fPccfp+Du4vs7F1XRk2UJmGskSP3jbiqMr
1THkyHxrtfKzCZC2XPiVr7P3HJvyFDaL2dwXqOmgiMXCbYiwxBL1gVBYXbvvOf2I
HK7flpqN4fFj50SQCKiQli47FeazLhEfv1TU9+II80Z2laiSHJChf9FLJEZIM8hm
j3beHajTbSYvdshoOE76jalrKZo5jvAn1s6oAcF9iWcHArLQvYvuW0jCxUj0bDoJ
rvCjmLNwCMLtbs8SZQ1SqqIJbOV5ycOTKKLz4cXTvjsE5Rkgsf/c8DAfD7NsgAtd
G2ysrzrmr61w7jhZgpF5nT9nA70IkvzgTCZcbnM9nqDpryroS2kFqBx431T/zAPW
lEmban5ypzlWRqCCJKPKQwSS3UROkiRkORq0mPukh42M9isOgYNVeyHa7YIpIMSC
WvAdU+6zLiHLsNtQMGqU/NwwYF/7gQP1XCKuYTymFqmIsdRxFa+Nsybyet5MxU1j
6lJewh0SZe0dpk6DlvzfecyIyPd3JRzQ5LdFKa27D0l+eUn7z/05DLUagO+orvv+
jfs4GiyyIgjPZs965kgqLM7AhGARrYg+THab4ZT+DkwWZMr7YMcSswV/aF9JW81r
LAFrMwRHQNwFs2eSzbqdYR/GEYHnO7sgNHyrpLHMmp/hJZxTOiQOUHNAT9T0PE9B
EN74n1iicuXs0e6q8DWtkVsHQoRvzkdt+4Ys0uTM7pLjYGJgAGNmpyuvTqLhZ3bJ
AbJnUSOgl+fy9tQXE7najdI/etCIUN9Th8kV5KHOkbugKUZJ9899UJwQ26UbOHQo
mQ8W+b8FylrfSzzdlgSVoC2KX8Ah3C2TGnJkpnzx4MwqIGQJa8hZLnmcDGRivr7G
i8gE/TxT1WO41dfhJ07arvcbq12oPx32W5MrlaTBz+M0rxiICn61i5RoNA9qtChG
/1wJPccUDiy0OzT3oo7/OjSp7jNOxwM03FDtEsyDIpM8oxgwOEA9jIhB7aEy3Xzl
krW5+Ih0AC5eyHC6hE/4M05erMYsrqxuuHXnLpua3TtCmtcOHe2naaTNjbm953M2
kr3YrT39anay5RzqfgdXHuw/1138QXXxZXnJIlLFdFFwVaAmUhTZKuTMlO1nV+Ut
O7qdNiHoPUYCzJ/+OrcRPTmCTFz8blr4f3pXrON3DycQvUWps1YSJiv3k7k1oLEW
g5qNzLceQ5NmLT66TyFPIovx8OS3E8HeVl0aOEfefhhUtE6s7s3t7/+PxgFME8C5
vooZg41FMX89wk4l7NHSrzr3QBtyV5ekdI5rONrm8WPHlBp4/SR1tUgQhBDND759
lciU9V36X2dj89pRKL3+tHVjvDTiDAG0oG8jblel2DTsvXYieXkDRZGdW8AXRlJo
B7wMBZFgwGM0ZVJfghVOFnV2VnfG+qbnAXIaL5TYU4iHJyPylUUJ/nOatPqU5rDq
zCaXckQudndXw/Cofd+r4g66puDm58w6jJiT75mzwFkwwr4JLP0mUdvnyg7Z3fh6
WjIq/lV7g8PzcXp9JelK0dUxuJ4S+wmn7gbUMndOuN4sCXuryaq6fa+grUb5t3IP
IQuyTHZDjK1cRTfpWXB+unHR9JHgI5VK3SwixSZUMM8DkXasSDrPfLWfZ8d7OOXn
IpgpOjHjVHQZuty2o2C7x/+9+0nAU4pTVlzgK5UegZ225Al/9yb2pduA1shYYdZp
LAl4V3GqavVhPTnjwmUgju0IIQcNQ27+I+gbX/XwXbaSN5YFTLT+sXFTCa2NCw9i
yJkMlu17W4gzeC3Z4eXDlWY+Vlp0FISpsHbIUS/2Cq2ouiptn0wDXDCWpSeLdrXS
97yE3sVixEN/JmdRcLWIUoMl6egWh0kKUr21hFfktFIijNxeJhQXsl0LlYIPZqdM
k+2DDk0rPOWGOI4v6xUOo5vL5GiN2kXSonAG+VbgqLkga13Noid6O6ywOOhhM37l
kZRjSq8ThCyA6NRv8/C+H8IElxZ/bnHnIdt1cb9ukctNu1c1Q51dVWH1v7R6a57m
6zfEPkufDKKMzq2t3xJ73SAwSXfkLne8KNjwKfa2csgzMWaCm/l0Fmkm1bZoDo0z
oq4dqDa+pOW8K7c3AQCrPfxS1vsBBH9c4wRKwXrdj6/aUNCgs+S5WmRvMrCk34pG
hwW+/IUUGWNGQHwFdScpjhM42VAXG8tDR56FFDCTpuIqh1YBGsqzEHTZB+25RO4x
68iGVe2d5jliOT+kXrItKRK7RCbpBO1qTN15xMJyvAaGaKpAPDE45wOZQowmdYCI
KG8GBxeZo7icj7rInzrq3vF+MiRhKtkfaFEJdP92b6nvyx9MJiBXJMJumtp4Lhph
T9DMDUw2KtIBjKrRuYR7C36H/OZcD791ucQvuH4paBTNYY73bk5m2zTmQsmL+vSu
CCHfAmJEBh/fSiKMrje2eLnev1AtK/L82/sW3JR17/xyKeVummcvK4IWqkebPsoT
PumpBa9oXm62OtOHTb5GMUVLyooIYTvAqnq4QDHaFtu7BL2+ET4ZlhduMIxzmICZ
Poa0PlVyt3Uiv9wuwcQ6SXRsKjckNQrk9YK38QINdnUd0rd4JJrqzslCNe5P/SdQ
4z71OehV89sQFv3D2GuPnuHdkdWZEPiTzxf4c+qpF5wvUC6wInyi0QWRxi/YoReR
AjU4D+GeZCo+f+qTJ5sgUYSlDY8Agob33SqBV8T0pC64KbG2kpb5OdUpb/ro6hTQ
m7/YqJIgD98H0Szt6q63ookPjV845Y0NHDzFZ+M40hilaoeMsTVJ9R//7H+arvkE
DgiIbDiaxnev2+6RCXmImFvju9NcnTYgXQ7Oar8PVexhSMc20lw/PGJVt4viBfRD
Jf5nKZ712P9kQyJbxXQ7hg5H8AadpxX12H6SEYXpYkCjB2GT3IJh131GqOoncy7a
tUBdLnX5nkrtucYY2YjB9jBWxsaVp71Z6/R2rJTykYCdjwWLmeSf/eG+TF1JyQQp
4yfo7SSnPgr9E23UNR45EM17+H8Y/OHX7mVYFrvDNlihIkKLUQSoUNflGdtk7qiR
fMjeic0Q4ey7EVBCTESSicJFwQuyCjNNfos/fIoeio6Y/4T+3w0Ijqjj9yutNmnI
JQmwlhUjOLTC59n247OHnzsHblV+0DUr6Sv+LXruvhlWJUIhUdPdJq/ldMDnthqg
IPZ/YtP/cXChxERjNClfwuOYbv0tlzoAouDeLg5c3VoT84WG9wRrub65FahnD9sr
9fZP5t2L3HOUChvokWTiAa1M4VuW7/TF7cBgC9NpyJtfFgvQUhP8Cz25C5ohQd70
eiWgfx6alef/UH+HQjajS66oyXDTL2PCVTy45cj9PGqAyzc47swQyTEyFbZXogIk
LLTQ/tl/MXr1DA72cCXJzzFtUwd4btZ6CQaPIPLFoFADV5I8tOfMRdJGve1ccux9
wtTy4+/EDh+t0h8rTwcRVKi+EFX/NMqvsEmn/RUvvi9hx0twZU+bXuETd29IFg0n
jXec4jn7AIEV19uqdIMpe+I6u6GuXNipenKovqHgeb+jySucJr3uesOZ5yR5LzV8
cx3m/ivY4VTBgYjjUHDij6NXj3/+KzlXxyB+b5Ed7lxEaa8fyGOdSBFW1zsWiNWP
ONJ6fVyvFDe1fsaBa1f4GnrH4LKHCNGmNZdrvpN5yvFrYqU6sCCX431J0HsZBMgK
UbTUiLa9fzhIbJ0fH4WBXpbsHIyboccCI/3DVK+e7dG2qnFBllP6pGZYbJcjxhLI
iHZAAZKY4unO+pa3FSIMKkj9M2RTsaEprdvRpN1LoYEttY3U/QW5ZDkGRsxnH78/
n0U9euL1M6NoOQENHhSbj99AQ9OnH+IRu3sm+P3lpqlB+3yyFcVszE6yyPQ8yWyX
XYmBmG3pI5CdW8BnmzFkzMdGULFXTKkd7lS+JCIFNiaunLo2ZdI0xWMYC+/H/ulD
naC/sEj2uthb1tn57Ubnfd3gg+2l4hbO8I+tYODQT6knuwlQxfWpFFpflClRTy35
ehRM0MN2AClXHTDzYcQ58llr0R/pAjsCAbpV+Pe//ua3aujdsYf2VS5njpNfk7nH
OqXTbVs/GA8U0omSgGRmJdW9aGBljySU3Rv0/Cf/dWXfkB3KHb2Wx0Axm1ga1Mrr
yr34VbMYs7hClKx0yhvZ0/e5U1TwXOA5Cuqq2Hle2EXwyVJ+kKOVwR5ackrVSz5i
8Nq8JrfJwvYn/t12+UrhrtigzXJ/KdgFGQO0JHzot9oahHMibTasZtrWQ/gTZJZ7
slfUC8AcOf9tjpM99xDtzFbAXKtL4k34no1crprLS7jVFX21rK6VMSAw0BodbRh2
HTrc0o452RmAq7Sq5cHeeYEYL/G80z++qVoTEZyFw1LRhYjiGzCmFX2XjXYVs7+h
2P1Sm3UyupEj+llOAqbyB5OlwrJnuTzJJ/kOAzAwa1K8xoWHx71QT0A+AKELhL6T
JCudyqOecucAjIljdjLdOie1o9u3jokbIv4uohuUyf5JspvApzNThdBOhvQqohDP
oi9t5PABzn6vzXJFbCCa+RQfR9x5MMqUegIGUTajb7b7JUyo9EZB34GtupJmNhCV
JVw2LUeiWfXuRIPGrvtoyPTsR2cPYyUtylybwBwDUTkP843zG96I9hDoc3Kh82l+
Vqml7NK090l9OXta1rZI4+XjQVobR7/hia+byycJeyjXCjUPKBQT66qvdaZRtbSB
JkjeTPh+LR6XQMHd+rPn3b3xgHeOOGPfZUKbKehkiEQli2yieFL3RBTGTrxihDE4
edlwwLBQP3FI43si3cpxJdymna793XpSk1kAI1TSAFg3hXo6clMxy6rwr0Y4E4i6
mL551NJl65IFX8sZN0Mr09r7HQ/h3lh8iRSESe3jH2mJC3WbpLOc7hQdVpyeZwX/
N8+JK+pkJaG86dsy5ltWRdjD8ls2l30PJ15uB/wy+Q9lfnaE8fJGTfyPMmHbHbkc
Jp2T/5T9Nqk0fp/o4ZWhI0NuFIPXVG7MHHMqbt/WP4yb/HO+rxH0WbzfRAL8sY4c
XIXM6ZPgGVKNcul5lvGqgQK+zra4pTKZJWfgLWAIi2Xp3mbvK9cZbz/OTBei1f25
LxuH6KFlbkIULrOrYzWFOOy8UXcKOpRqywaSSNp2hcemgEutmdbuhmRoPHGeE6TG
3xSKiS6FssXY2kx0e/Yq7WpUE872B56Gp55/mkBR1pnw7D+psbFoNmLk9e/FKD96
y6tpF4qBQRkuM7qnJXawH9Q6aOHtvtD4tIKfPR4S+0VUCajkkJIJcSO8jzG6qBPF
0chb8gTjnUuQfF109g9pEGP6Ky2bg9YSGZcirZwy3QvjARJkehUkytBIxdDNwmeS
ez+kZg6C8QMrNaFIGge8e7casXngZLIjT6+MvOVMO4zGOkB7HloS7Epr90NUc+0G
JH5fsMPR6uWFX9++eTD31JW8MI1lXy16HX9nA6t68y6HWr9wLbr+FXblPKyARDEE
Zwr2tm+IN33dulSo/xyrvW+WGVw8Tao1RkJtlqSiBJn6oJfveBPL890LDq2+ayRV
YpyVZLWyjlCYKdBPialqJ7JXmA/ekYfRzr+5kj0FlsqAU+UlaUxLd7vlTEm20ypA
u6E48xFFjQdnPpIJQfR0MNcoHdSF5kpsclBccVKIRd05U8GwDxeuf1zfnXUgo4bL
XmeZ5RaXp6TRg1NJEUwSgzHiuat7KzxhX8TpLYClRn+6gIzaAXn4iLvAIrNROkB1
i+NoTmnhtGh32o3A/8iKc53YJgvrjT14pkpXej1l/p/yggiHVMmIMPglSY9STiLP
HzFIyjmDz68S06PmO3/vjF2cnIiykXF9S3Z7A2K9h6LT2733u5zGgNFhcqYOlPT9
koilzJDa8XAvTbc7+sOmGQ+yttGd+vqDVQ5j2eNQPUCOQ0bKDUCruLhnyannixuw
05465g53Vu9nah/GXqx6Nm3mGmL6RSnmqQDdqg8fyrBbq2XUZyg/KSFp/0+YWe/9
moWUWQFfygZQE3Qba83DmhkZVueXS61Apsi+26i2a6HadeheXPzBq2kNfhptr7p0
Qr4mEmIw36jjKp730zUvQBJPQFg7XfxuN6lWEofiUyc9SlC6KRjen2MnMV/sS/22
+T98SsFqdjnzpL3RIFKk0AP+t1HlBpLrMmcbZwb5ELq0kL+V2fxDDHa/APXm/64N
N8B1wz9mfbh5sSxJsqf+eHWbbnaEstXha/nQYZcPHNN2pxFiVxqTFtD7LxCu5vcT
4ROuPK+JQOBmTr34Cg9NuIha0wT2xcN9Thhds98AMk3DRiJ6K09X9cMrHy0mS3vT
epHC8trxS0+9lAPH203xTwv8EDxnVk7M9TWkzfrsfvY9X2nXvHVSzS4T88UOsC8Y
B0ROgfLWHQXmwW/SRDUIANPkfGRNSCFnuZFE1GWO0ZQYmWFh8MqFNiKBUvG7Q4gV
PypuuwXrSdBV1MVbtfRbV1+K7ViOah9jkNtnoMf50PrkYAG0/nhz4fpo1Rs5Tzex
00qqBxUO4QytHRWG67qLJ9yMzCoI458GR4/Io7JiTqrufvkHcDjgyAvMa6ysPihq
fyRAHC8cz1N2N/PK6dq1RBLrHQ+HAkXWtRJyuknxcL/noANdFKkkKbJsLneOTSRC
5/pVGzHVK/bR1m2tThSq/1P3Kc4nr7JhMH7A1j5rqhCPNqm4gAD/YlkAC7oJkHTP
d5BuRYshpob5P5wWLMdQjyQpYmtUJucOSj+sY3Sh24QdRR1qAI/moWfEqexl5pk6
sO9lW1geb6gAsog4LAnhVTWJK+EA+HnZ0T+uudL0fbMnYZXDccc7T1FtJGub/n38
z/NFi0MWSQAHle1NDObFA68yfmH+WYEjFcvhEZxfxEANm+zeEHhheQ6yXTOVt6lW
UwPSLsgHq1doBDskc+UHU5fuEGawcAWCtHtqyoH4uu9i+GhBep0G0cG1g9Dd7F0F
pU3H4BLMoTo4dTZO1UqiYZTNfspZqlR/ZD0yhCDqNt4XMsL53kCEYAauu33Riyr1
c/BtvXj5xKPyE6h7oIh4f4CumPMqY6UBbuhhbl+lsc7ZFgIg8RnBXgJjl7WVHPZn
/B5r7arb6vcsYcaQQ5tbi72RaRoAkOH+W/3Gn/RysNfy9lzeT/ji7wmzgH0zhmlh
AghEIocmREkp3qrdv+jNzzPe3dJx3T4//9a6zZXjANwSJhhmBebfdu8YGEgEW19b
OMSUR4C7oPFmwXzh+qAnfBE7eyDqVgQBJ362WcQ9wz9v0pcOul17jmm2ZlN/yYX2
s8cY+Cyqu3ONS1IU/fprt0cp9wEwGKJ4F73WDJYMKhUFgubKOtRDDHr/cFzas4H1
Curry47VvxkerCrXB/sFVr+4ipO4Tc0hFqIcFoHHoIVT/EO3SXmrF0SR3xnUxLlu
Prm7nnP41ASN6Oh3qNNJrQWB/yWlaNnmr83N3aH8rTEDWcmSBlCJopthnVJ1Fa2K
/+o1PQdy0gRyBzJDWXtH+zO7TkrnMLE7NXjFhpcsZ7AwwjyDQbmTkfFVCE7W/ACU
VH5r0zWZ0VlWdU9OQJdI7E5QtGZZurRpHzv+gb1L9oMlJdZvuG9zUp+S5iusIOSZ
sI7e+YA8CdXhVgKtiuUoQU3u/gG3YFJLpUfGVHRU4sZDwc5s75aZPenyFKNPICOS
xP/xfBJ95wG4JuLYNT+9tSzLiynt/uI86mrgVrF2doWeV3ACq7czHV0BgitXmISC
DsEqThUkgbMjg7lnghNakkllFZR5jC4j0K4Rvaqm39lP4vw5Zr6LopbJ2Q5Rfyaz
w5ZG6QGG3UHOo58NM9bQz0f781i/iPssqinqsxGsIWnziY5uAjcajD9ApHf37VPM
P26xaqv5yXlOucWyxJWzCKXzGOl7FsSapG1YsuAsMMvFp8CDQvQBtkQNr3FglEvN
I8mwzaa5oJ8fzCDUM0w1UqrJtqjWTwJqCmLtvjCQO99VTZP3Vf1Kqjjlq5TrBXL2
pVF6Ob1spXZBpirCMIZ/+VVhda+l9xeOSEd/8U+sun+RhR0BoPN/m/p3ghy1S0Y9
GvSH3oBVJQf+fIICRaC18VEqGAASDlD0qBu/4htl+gRoO+eswfMlNvO/uqWiqHnH
UOWODlbaR13cCq+uTq7F7Nl+/jv3iB1ClVzGwlhoOAM9vLdEax5jROCHef8pkaRE
/RJzQHAmnKpn9/7ml343tqHUEsPepa3tCgbDNNS31TTNl/3dmwqmaNOs7wjEHvtf
fIurMMoOJTAtxgzIINL+ELHuVYgxv/r8i4BYKN77/AHbr76FOlBt0T8XcE0zOuen
uGxBz9XuaiCBq4CexevqV6j3McNzp7V84grCSqharbx9ydrM1ZX2wklVHpbE4Xz9
Xv6/UyIscB32cgnVpghwSRArt8XeWhRYWI4QgL3XEmcK9Vrd23xNybWXjKE1OGRg
LXbOJH3ub7jnSQj9J8W5lz4LmvAHIpX7SfCk7CSdyrL7+djsGkqv4ovNF5te01ho
gIkolHTEiIde1+NfmXqM8szPb+/3rlTX97DPjmAd0kmcKFCJcpcWTOyeqPoCMwrc
lbojv8j58EE+g084uS52C2VxmygD9328tXkLsJzhxglBife7Sx066HOn9TNeT46A
k6+F7AbOUHiyTNSTWl97e5EfJ3WehyTw5gkFaDlQfXSrBb3zf+GulTAhIfBYOO8G
MO251tBMglY3JEjChQySsL6hc+mIfm21bly7Jc5bmsvE8ZJ/MG+j8Usphbg6C09l
29XbTcnObvGzqNaNnLPS1LCG5wpoMznkKOCOiK6z3oqSdz/UmiRvQgAU3kFyIYDj
R10E3OBME8GwT2Yb6FsxCLFGYHMngUM27VgXNaqZ/almvDnp+aOu5sh1LQJWtab+
SQQQxACmljDRv5ax2U7v0He2iw7xLOq7/mcwyWUoQr7wtNEwZqXq2ONql/ug4XTx
L0MUxEPrzw3Ohz+EHk01MrQqp79eRf4MnOY9ZwiduV5x1bzBjAiMLjkMzgv//9dn
4MKblQIUbdegwzsUipLXHyHxqENisuNZZOoS0lblwd692S4aeIruDoCiHQD47Ni8
vfQE5rJTYq1eC2aTp4XhKUU4NohZqmSXv0p1bEhQrDD0Bo42pduakFLOnmdXpP8T
tgPvQJ2WMoKtr3zM15uHCvcCKiqJcJHCKPV52RNeMTk48as8hweOneyUdVjYbZxV
K8YErFRuEOtLFSTZ7n0Naxv9oRCFgDe/lZpFXV3Z2BcRs+EaKwQGdtgGV5nVBlyX
fOO/pEq+FyHzYwXpRsoNjPk6ICiLZ5m8+5O8TikfT63+T/Rmlq+9w5xoM/SavSpz
dLITBWXOZgrytlNnN7GZMbakZhFyIVvXDUebCtsb6oBvvgPIQDN1+tnjgePzxvXz
w+m/D97Yucjzsg/GfFUeT9vj9zjMmse3QjJ7Al17xOv0OWME8IJOxlW5cKYsMpgf
9F2vmli5APs+301WluEeEe2bX2e8hq5hhPFSIc3zV2SbbC6EZv669ruoqrQzzgME
fC0sHNQ58RIAE9UAxbreWX/cfMC5qyoD7lyJ+3HmzO+wmPAcleN2cf/0jw4tjf42
dETD8ZPZiSsDSV4zOS/Ynqr9QDbJRkRrA4Yf4qNWai1nFzW76iR0zH1vVhMgLQ+D
nVvIiW/8ckDdpLAvlVwzyF1PgFV6aZq9PDmxU/tdeZH5QtJveCmX+hzUoDpUkfO8
KLPgKQ2buyDycVlZ79dr7qZuaIaXXSRQSep3GaUP5hxWxxSVHyvjDsVbj+KMq49U
QSdaMkLEWAPrBgHpP5VapfmqkEKGXd3jU2QJIKm3SNYyg9xflvSdsz7uHG0WqTES
wuHlY1OH3w1TeoxXZwUjOplh8tEJDrPt5R5Y3dn2MILRENgyvLplUZrIyQWYekPv
QYrMm3GQ1kipWMJct4+UVQkljD1+UMff049h+XL2z9bv5YGucbVBn78QHao7vRVw
yHKw4NAR+bXylYtKERwU4nV7UOtRN7UbexFVHd4kh0vJAle8tO27qKuyd55u8uao
TpXMUPmitcsONDOAZ8Hm8is/0hRiE/ShzRMOgUbt8S9Zeqw5ypBrGzL/2qtGPMT5
qTdP5kgAsrlqkaT6a6gdNI256htb/LqEIzPjvsz7Lq/hPY1bwP6hqRAMjb4jj3Y4
70KSKoio3RcXhgDtja8XMJPi7ahm1kO3K50zpoiRmi9yZj0h6a8gjuEgWOQKHmSg
AnG1elXoHrhJtU6y0jpA1M2EAzdoUZZBzL4ObwJTjhOPPIndWnY7aiiBaPuk4TK0
BWjyl6pKiKLFagA6LVaGxlopsSnQy+e4LhxgiDVA58uiF8qdEtgdJhNzBz1lPEVo
43zYYbPZZ1Aa41xMMeMHR6qtfc5RyllwLSgQzrfh9IYU9BiKKEUZZ735ahaTb8WA
7H58BkQuJ8zARxnRKvZGLeKdv2iGMYw1NSnmcVezomz1OZMiGKKeiS3ynRkiJl93
TceIirHwvn1RizAIqCn2aHpu3nXXyUJF+3KwKqOGP0GtUWJTK6uVCuBnYraK6V1U
0W7Qt/pN/2YTPGpsMH3P4AjPQcU29gk+mSqz9gBALaSOzvegWT/qMpNb4Zz2y9NB
jkfaU9j9apdmiVvMdMMmLzO7XW47CYvyuVKfkukx/f8uc59W1nvwnUltuUhGRssX
L+74108P+iV3qrVcscl+1Oz8hUmsIlZm8QxUB0FO3039rqf5ZdfF0aQbRkMsb/eY
MjWPlv9w1SwHxg/Hq7V0M5DXeu0TT5HA00JAAipRiin/6XLgVn5UNBBom9KYwj2R
mjOtR4rBfkcOnJ8PgEZSV5zjxx4X+J0BxA2T5ijrp2EMk5QS9NY3+Hb4P0RvQCzU
z1VX2qT2s9RbPyWhUnd8ZG2po5Cs7lbjK/glmJv7uiLHQOPKLU9Zieh5LsK2TmZw
nfcLqralHKxu9KMJcPWRaQVwz1aYK1fD199hCcfFDczI3QgB2o+Sr55EBH8jwkQQ
OecfeRiJ9xeMmW/wupdTY5uyI+fTOQVwc6gnJ8InVwO5Zy0OnGqsO07WE1QEeAIJ
esF6tce4qPYPjGp9NfL00FDuP1T0mIQrcLL0yDLz6dBHU5cq2XE7fUZkx8KVT4s2
Pz9vT0yuHbdYuZ3TqTQ6LfScWwT50MABXb503JZzuqOGODCh8aSEtJN8XCIoNhJv
AEFJqlHWM7MspRMl5Oa7N0rA5QsWc/J7JfvvzNnxeMRErH/kSczd50zAXCxG2olJ
P9B0SD7Vv1WenPPiX/yFSZh9hFzh+uL3H8+i6P2vF9kLRShUIrGTyJM2PtSsw421
XbMjoR9A/xpSfCviXP9gD6iYkFouaNTUHPK2Nma4QOaq88jne68UMHXEieEumX5O
ouQswyQIA7WYlaq41j2NJ5BtdDqbXh91k9aEngD+9LsLu6o4qAt3LdYmmEhZA0Ys
zVXpHwOZDduuA/s0JN28RKoiAVxq1vNBRyah2GgfIMDPGEZHuT3ht29B1Bb0/xhn
R3V3xrquM9DYfxrtkwmYsvRRiXEjuhiseA4zEfFzLWVmZlMYbmeW8G4BenoQCpTu
RMlFQIoA2fDXAso0Emnur/0sxnttikagaRyxFfEqDcuFg4j5SCN+OBdMSKSE9J3V
rJ+wNQ8AQKEjzgGDdm/Zz+MPIRDyNMPT76eNbLVrRQoyBfobTllOD/u+ATX/mHqU
eoXZEpnOYoKqkavQF1JIxnK3GPOIzOkV53OovBg9Rvu8122A+TlrldyBHAAfQI52
1hnqzD3lp2dkcMM4dHTzQUEKUAlKobm7ZWBV1a24wx7wXyVIafxaMM5Ugr7mDgPb
upQTM9phzcFqa4RqyT05/lKFsp+VG3sFEQFNE92Qhxyx6fpkxc+cQbueqT8gLeDp
9RCk9a+9PTUWFOyMDXTrH3FMTiJR7SJmeunVyiUpmY1tk0iw6u8j+nWeArgn8qUH
kK0HME4GCjACUGMJUmkgs+JALEEjU6xC/rCcypi9tzzza7DDSDTIBhbzQA3i9hPA
ioi//vve3si0ui5lCRy1+3oha15C9fdHnqM4Ip2v+oOS17uZnAu4IrZiI0k/v82z
jiBUZhkq0yvtGWEnZdyPYAVTMLnm9hI4ZXbKvuzlRVP1+t5hgI/+LDWoDs07RwG3
cP/gMLjF5J18zjOeUU4mpOSnXeIcPmVwwmadFxDHPj1E3X1RQMAArBXYCDq5DGVd
PiIXhc9j0zOmzyoL3KHbaLDhCV0bqcOJpkVgjL8Hg8NLqns2AfDtiDZq+292xPZR
LVH9C4Mu14ZlL5xcXB6PA3v7NKExwG843SBukPHuPH+OtpTfUvtgMhdK5nDnIEu2
b9VHahFLLNDmnMmNItJ5ASJmnVrHvso7y8bc7jWb6cxWSpS/odhTacO4d0BZrqBd
W1yfJuEVw00BqBUAzUY4xAqDWPXVXplVl5RlC9gEsCN/FywcFQKcsl0GIqhcfh7c
JWWRKngN4ZtOYHD/NVevLXE/zA9FwD1uT2Grv3XkshwoTOH3OP64+JoPY5u01enH
yE7uMgKch4GJJWlXBvP0cF0ZOBiPkSrYqYWrYQw75mCgPh+H6HT9WjXV6XGLxKPm
UvZj/C+IiCT8Lnrci2ZSEXMfpB8eoqNCbyjeEx6vXRsSq9f5Z+zNdOy9rRJvLoP7
daQPjS0jXv+8/kPXYH1nMk0K7TiiAKR1GgZLBEPYWeNcWd2BO2WyjDdPt0G/JmX3
zys4VRJ303QdD7UaP6ckDCvBHzRl+EchwgELY5jnZRkBkQ5Ri/AVytGHzEJ89rcz
6zHLTyTD9uMYE5WfSeN9ZhULGM7NLRMBp2wL9lxFUSDJAg+LnvK4YeGIX6ZZs6EL
DWALcJAz2BA6juOByZG+tMw2KG59e22ctol5W86T0HFXb/BdhAzcOmiXZS0vTaSz
SGKBBcp/PdyuM+IX9pDh3pka3pLwCHvCylQZP1Hk3IOvZx8urHyafIo2OCXyuhgh
NimtDRSvszWcc6m8oFhSAGz1VsgYA+Lpb6M1tKlRBGpA6BZyoWQ0fmImLs8tOlOQ
CQLjPBI68hlOIvpkqQfOgVj5J2/SBNDEbzthsn6lUuwA0MFk9xj1KEFntceUWRgg
X/yXOCXWRy0/K5BWNeVV11WDMi4eM0wqGEpQwLnh6xgQKhYUDhmxGGc819xnAqBd
T6CZckB4kCxI0hGThsunBN0m3r15zqcyEYIYLmtW8GQd0+vQAEFVdumI9rSTLTcJ
apFH8cR7shqQwxUhKvY5mpP/c2+QL1UqEn6v5FhnzrXnfF88H1eqqxVSWBgq9ani
bO5X2nMvmfU5BU7K/7gicrl9l5gaQfH2n19jzF3l6zeqyWPwPMfLeUxAJagJsXWj
5cUFIB8r5CMYFFQdT4LwPgkHdjLAX+8Gq7mbo22rYiGLCj3vGxeOx0P/vW33VaMg
9lukoLhnIJ2HzlGgH8sCARzj2a0WUvegQV6KGeUOZFWOfv8z2s4JZoTbJU4xB9nA
HW6NfmESnX1I3wX4AG/deDk8CBmz2Xq0gBaSOMHpyg4kY1i5JqvQDyji5/3TGpXr
8MA/X8I+iHGo0ZbRwmg+7DcmIifLEply/xTM0x3A/TCdQAX9BuMdGzVhaCtONB1q
zx5LbTEpSohGsaGzVaJfP7LckzW4+WEw0r7WEh/usNj2LAapLu8cU1wf8eXjynAn
roZMBPyypEeFws9KxWpXFlQwx8l9zPe50GFobGRJ0HrSST9KlFk3jedgbCdt/3lm
YsjvoQewGlGWK4Q5mXoA+yjGa33dAZtFloSDEWPCddro9os8LJkAmprjjYm0Brd6
sXNHZg6KVEwuDTSQ4nX24kDjAaWUwYgkUw8ddQmIQdgcxxDSamJgSaIMRAF8GKvX
JF7L678TERcuFpPM/YipN9c4rmAbrUVjH+zvz8kR/NXEI9bHcaB9lnahwC8mhRkq
oZ+gNQSwCgruWjGpNq1TTKDTkhorGW6gFmsFMMOGVmqUnvj/cldREDl7MVHDD4DY
rRwdVZ5ajcOOztlm7PGlATMlqhwjHCvBfdyWAih+2k51xkTOn1SzxwTc1VGDUgK9
MyvxsU3/RVHtyIPFv3kdK6TUwyhgWdrYM6/fT49La2p5L6CWxmEt8ahYwDCyAeVh
fkkeUR4jFvXfwoErSfZSPmRqJeZREtgpL82HGa7nHNL98qpHjjdCvlFCAce4Wslg
o+TEpG+eSWsz9ryUttEf8ZdHbRvgDqibY6Svs72+vvuuO+VJ3TDBhNpaUpUG7zJc
0/hDpg6JDnvluoytZzjG32/rla83Z2i93EM9S67i/9EVW0EXqLmj0jLIKv/Cd5O5
tfCU3RtKjPspqgT6QPee1QgWqrOHJ+sdnLfD1Ch/BQOrU4bqgFOvQOma3+frhKZi
kIGHh1/x+f2KB7x7yltTCgypgWwO6K+hikSNLyaoGqEzfy0qkpfw8E0xgYRLnMIQ
nHL2bHn2X8IBrBp+W8/12fsac28YjqDzHXgu2tL41py2aMcbr4foy0qmHKQ6HRyF
RdFlOcPZM+KYbzUBotj8pAIApEAmVFEu90eY2mfW9Cj4bnB5F1donOTZRJ5tc6P0
FnTvRkgfuxmzHW1W4T5ojOrCVIyGlOuLeipQCLkFHaB4mUIby8cTVZdAUqomPKuf
LKa7T0I5JQ9nO+5MwPkGiRduNNAzSELrUuWkpDFHGclXmoB3tm9LsZKFR6iDFZi8
3PxEFPYT9bfvYhIRDYo41Aey8ZS+QmroS2TuFl2GMs8UqcFXnEHKW1eOr3ChjVEq
ndbyK47BwwAl+Bm+I/N3Ugl/DU9gEZ62E9yhSBHEBpiLM12tSwH2Z6PON74e4anj
HQKniUFo7hlJRUw0F937ehPCRX6CLlr9FPCXzGNc2v5tyu07xn0HMLhIS1lVXr7A
1VgOJxFMEtdL7EktdmRGRn8nY05IHY2HovZQ2tECVm4TErXovRKWvKiJfCKCh3il
50kTjzbY4LPUl+CJ1YJ+ACvzinZapviGA6ddXQjH3C6aoRHHqolURGQPgH7fb1C1
cTd8bVW05OccaKZKCn6PgTIzwkW800rPFBlQUW1x+GJzbLlz/JPVFTdbIaZG86Eu
Mweu1vNXj9MjntgpDv4w9TLeCUDoDS/W4g+jRXuHGLkr8O/KR4w41WSmfnD/x1Qa
NDda11LoLA221YEluUEwuhMlpU038MTQqNNRjOA6+u4SKoAjsHdxgfKYwRQ8IvDl
dEnS/ZMxicJlrIHX1kxmVQoM0/RJUpRpQjVtLK4rKJnoQLdtHQfthVyA0tGfZp+v
xKGm4/uP91aCFXm28tpvxE+TvKxHWZa+rby9uHLGSyjsRreET+w4g3dHrW3qImsN
b4PzbYiBStUB9uvFWG2SRq/JI0nd1I96sXZ+9CfVqDlrrdWRhTv3jDE6Q+LRvyFI
tmgp+VXiViBzfNn3WncAERjzinxQSpisA68g1PV127d/xzoIuMGcMGe4BwA+iRUZ
BLNfLlop9nIJpjIbEF4li9DYpsxbESsAFel9mmIcC+ssGXThm/R3cSDHJNQBdMNS
ufHkcCkP5CoxQsj7K67w3MJSPsZMNEolAgspSfL9rWgRTJ5JNeGITf3h2DgBbjlu
kMMwRZrfCqFVkXCoPvVKWPQDIlko+o3taljx+fkTpZ84uGhIzWBgurL3XYX+jUkn
S0ZXQI7EqOrk9u5ufhpDB+oiRRM6veHbwt4q/QChCCaYv5eBcF3dfNd2pMghZNQh
HxQB2ri0EnsFLhKXIV/LyE7ldrgIUS4pOxQLK9XmYsZ45t+sd4nai4qp5nIFDnTh
SaCYY3XR5s4hUh2i3p0D2yfqSF/gbc91VgMasOnEBxvggdoDhNOiZ+6VBY1SCn0u
I7gIN9VDroId9WPPuK045WlQvOdUDRZC09d5OUYMwyonZu9hJNTL8eywEtbjFdxS
tTynn8Zc5wCbMFr9C2vFx8RpoTXDiIUDtcbzxx25EFzXgwVB6+VcTj0w7fGJx8lM
0bKmHEJVumsQNu3AHd3lWgfXSM/3VhyHHZfHMNlWfNWpx6qZOrLJ9KhBOwZxG6J9
vXuoUhPLTbzE2OPqpQIlnmC0ZIjFkSnYxcq+8rPRFodJYR2BBYjIFCbi3kgnoSXg
JrH4iPVqmebdlgyxUi3yt2SkL9en/VMt0SoebYlRUeX5t/M2xKOAWVXrcPvyUHlM
8JllVtrwwrlVmElYhU5z+PDLSeAkzFfznDwsyFjr1hGuEwd779r7TiRTP4XIfsHp
qRXPML4amSVA3DFbbDP1mxUT6SXkmJk5FaJNhdFaV12lAdQUbDO14to6w4R+jVuo
13UwYrLtrv8rtLNvKmMcvg8Ai6y9ub1G9nfP7D2CPjBkc0yUn9HDzILPcZ8nbQ5z
THOEEsLp+YT5XTsH7Iki5g3jsH+WqdXZVP1i/Qb1B0QaV+cDJWCV7RgvO/Dtvl7p
/RkIEfX3l/NQDZVPgVPaG4d5WQit4lUrUw62FYBZDyy9vKMyquT5tw8NXo8PxXiz
qhNcVIW1ygAI6dn+Q3AvmS2CVMw+nCNgyfUMGIwo9ZiU6824xtt//pIb+MLcwTvV
sgaNIFl+z0I974mr8DaR1o/MPJgQCOn+05/1jk5Rp8/2d5NmPNfFzi0cBeWzkJCT
0XLtlyJFiHBJ3RntMxyIjN0knXy+NXia5fWmZfqH4sBMkCpPwwvogE16yxJx4r5H
nM9dRZ3cc6j51ltaB7lpnBWjXImiYoQ4pBs7CyDAXlKZbMPgAH8LZqFrKoMi5Aal
74ElffQCZc8tsU/ADT74X1n8WrAXV9f9sQ6vIOvpKySiclpWZQS/NNuTr0f+g33t
RAPnNLk6iGErN42RUEe2Eqk8eyQo9zpO15hm+k9EGvZPiE8TdoNaJN71MYySCdr6
aQXFhfmnz41cze6hZYnsxf7m0FN9KFda1TzTGTaSlO4gzwRuvK6S2XPSS8nyc7PH
gzaEhXFk++J61yT6x+WKCSBEtLCF79vz0/fglVMwKZRCZPI2hxJY4liVz4qZWubz
N1pFIOzc5Ic5yKBRz6hYtYZx5Ttyr5ZyaStMOl5cjm3J7iivcxkPz5+3kqOyPThq
oTZlF4ibYiufudo9oYB+9fZLpNM29sOR2wJio2tnQe7GU9rLo6A+bIcCUIsS7fP3
DTSvggYqx278LCHGvtHjJq6Gei7LR3A8ZGC9+fXdJZ9mept2qledSjt/QqjhPQ88
jPnGsW20urWTGBHuopZjNmxfuzdvCrOqrNgsBGk806ZQ1B8G/zMd7XCJ5HNkJr5y
j2TrXhm9b879rC7lR3Uig7Mrke3DucGe7i8WBW3zH8BunxtCKMuNku2DOc9mU4F+
iEA+kh/nRb7rYdcn1+R5VNor/q8redmVDGLdgAy0L1Ss5hG9L/Lhip/jsFLWGGeI
nSiC2eM61mOBmKQELxXlf1fYU/grP2aHsxkot/iuPpJJfJJtHLg6wZGNmjNp8ViM
iL78UJs+2NGVPW1udipKoKc/epY2qiLSkCJ9xAt6H2NehnbCVMbiZWh/g2nSYfXU
qmu1r3W8tP5sYhXCxulufPuC7wz//3DcTztJUEOEUPrcC05zEe6hHxWFcIbXGEgf
GJUN+91P1d55qgVoPrE8pgKXx3H6K0UDlwm9a6y1YZVJml2zUBKonq0mijxnXvPA
MRhpHkqgCBoTM2XCaES3JvYoa/n5drroW+q8wN+JjDksH12TvPGjVFAt3v/cy+yY
q8ZzvrSsSufeDLICMQ5ChsoQton45b6piXLBLMCVqFZxBoK2TrURJPEyQsljGTO0
rMoK2xCqrEjGwzQAIrQYztccKwri0MoDm5SlN1/tPl8IMbQWBIzMhENrskbyhxWa
ZQn/BXgAt/PiYuiEXEbydqZEsj5VpIWI591j4gsFFNkPR8SmZS4Ml6OHUVxbp3Vu
ADlO6YlAucjMuhPW8l0M4nce/JxFAt5SVEN0FfMsHEkCD2pIsAJgKDALjIAR4ezn
TSbEVkKqCK7hgJapu25UbRgILRLLG/jHmYJN1gJKmzLlEVs6BZ9P4m+uXnkY+vJc
XZKoyLXs76qpCw79be6pSpsIRntu2HezEer9t5lsv34FnK2W3ON4tD32aep87h+M
xt2I74is/gxbkJLQud8dL+v7KdX/F5JVS2TvIP6odtzNq3Wrai2pRSr+g5i/YmtM
ZqPhysUUOohTkKzUpx8lJqpLWNEOyh9e0l9iLdkCtUx1q9eyGXrda6SdWGVOvuCh
kqybc/jIuCdhXECd/NV+wLl5UzEhN7Pze1JfYPp+msn/FttL25tTy6acsIrw+cA+
pXX3LF70vvyjj6WsgqINsFLHdeS+Dgx8/pDKK99wWjtEHXGb1o65wfl2DauaJN/v
fCKs/IDWYlybOaa2zHO3Ir7Lr6++HfQfQvCeg4sMglUjby3OF1u2fwdlSBfd9qIe
8VWa0cwdLNgbCNCaFvWyKm39v/FXPgAOM10GjXkFab/PKf4oNWgAXlFj16y++3Bo
gU+lVbUFN0JNd75JNErAUJ3eZFAXoHmGzqEYyMsF59FHBQ/ElTsGX9OBduvzEGyl
+bs32Dl7Jn06WmQRWjwH+oIy4qJ1fdWHN21FKNs3C0FrBZ9mPoYu71Ty7zkORsWW
dh9qZ4d5Rlv9SPxveGqafTKNi+Fq9JDBfbgjJNE81fDdVsRDrFJba/eG9QpUfx7G
nHXgD/dnIzSVsXwbFbaOfakTwCXOQ2aZTQlu5sE+ICICObeA866AJToZYUDDXRua
ZN6pwFFcK4sTe1mlyFTj4JklOIKYuHsaNEezULHJAjsfn1Xx3w0cSLJZeva+D/3h
znMGrDbIJ0FgNQZ/k6H7O8FtJ+Ak90daoKEATwPgnjTyhk7FapGr2BOH/+cN5D2X
9cBK9nyUU4/YGAoK0pVAJO0oYYs43W6dprHHJOLZbu+MCH4L+9Z6ahUAG6uzncLk
i8P0R/QrvCyXikQGJH4Ua99f+eW7L1ehwPwL2AiorAb0plbpxoLjxEZLgM7bceyr
5Jo6C2H2M3fvD9YrG7poxY/mAYUq36uF5Q2ytJ1kRpfAXgcGyQo2UnWswa4L49M+
SkSBT1AOhCr9vcpokX4p0La0cy4GVzXho9NhCQMzcv7k0dQPeW1AAMgqlQQ/RYB8
FWMWPd49UyHjgTG3IeysCrsOl7gT2x66Cyh9L/PhVsswoPaZNfMh7uTwvRLeWpvH
ylrki4oAjyhNxgh/ioPxmVIxU3ceymoBRS6ptZ5PfwKINU563e2a8MXQvhOfveeO
QuqtTmnXV0TBjBz5aB2e6bmyQHvfb0dbLI3zV0OiYvTjTnDYzc4dd913D+rz8pwd
jDdn5dTVpMdICn5diW23e/xh0Jhu498mt6niNAMpN06FQqQxAER6Bx0XN6ywVixr
z+cUxmfgMlJFz4ZvgBOnPsR+AS2HQghBA3RnaFbs1Ot7pxtAAXCkak1VZ/udySSt
5sr7nDXtwkpBh5StJYepSRLoFD02OEFaO4kpelLExvGctUboRCg4KWjfSftDpPnk
ReiqYuWOzrW2bNOgq08XrwzBDzEiHV/b9zynhqsmwWLh+3uI4a3skblqm7rtdDgF
yCrS0eDAgRVN265zi1J+2Esyg7rrb7c/J9kqhA7skSfL5rvGSrP9R65ndVyR4+AU
A3zcbPhR0aL7F/tj5WG/r7kCswXcT+K1+5QpeDlERHH/jU1A3RNgpWvbKdJRfrTV
+HSQ5N7EXD7uBgIHRIOZ3X4zrFUw4yqIu2vNUpIgNDO/6Gv4RziioT/Lv8ObGLhd
I3l0KUaZ2R/mrrG0pspEfjaSqp1OqTaW++/7fRJZDEkjTweDtGHxZFASXowFiPMW
lc98f34FgHKv2CfIi8p5wrrYNNUSJSKxKCFMuSuaQb+Obr4EVZK6hLCsx/CidQYb
bZx+deRmuSTiYz7lwwg2BN+54Li5wvIg33ruwXQjyqmuH60mr3ZoW7SRylIPK7Zz
ZI0nwkcZVx9PB1K6ERtDwPvEyGwCQYbopyWVAsi/rRZR3Bg0xCnLmQ2zgLtirwG5
Xo91M7aTUgVYDFzUwEjWlENi50KNP2Kg64ji0H2i6gP27Qbvo/+sqkcX+yrsIu44
tVdX7qW0SINXHmz9ZGGM3QLfzIzMYtCjNT9Uwyclmapx+t+ms3fz0v4OsHI6dSWq
yNV+OFAo4BhRG9yFvzIcRQahqSyVVRnnwtspf8DuEiGZ2e0scfNhjk+JKfAH5HSM
iNuOO0ZPTOpQx0jYh0UEY1uBUolW5OlbjlR50/fTVDj/nCtRMrGtIncxKX8R6NN6
FLEOq378QqbXiZf/jnzn9iHs8ygkS5oaWxj0GMu2CJtmT3/WJfdvPMhXrptWXDSF
KOLBJ9CsTR+YJmljtC2mqrF69PremIaa8jHf2/34/w0mhsWWMMw1E26CeccNZ4nB
VTtzUkfzk+rA26BFziKrms492hzVnXod5n+ie8Pw03UGJYGsO2R0SDI8qX+dxgt2
01vxM8J34DWBaosWHcpm6bsLtN3CF+/Y5vS14+N5ks8i1s5alwuyalCeYjaesbZw
txH/kht8k/GSR64GFkJ9e3KTIWRr26J++apL4okVsrkUC4rqda9Tc4Gcfx18cJjW
Woz2pbAVqoqh42TefrE5zbTevdCcj48spIPX0fNskhtrBZh9mFD++MhTkzQO0ujd
Se4N3/xuhl2ezgGCRSUprj2pSDqtlGIF3Gbe1iO7Ffo7y8Qf1pLg8y1yOB1999DM
bikxW8uMDnRPv8/YUVi9+N/gwvxuviuyFw61BVZRGlQFHAwFKgLOyfuUZ+1bjPLv
2rWmCxs8dcTSoNtNxlfk+RlIxn5BdUduz3VxUkapxdQVBY0y0jovD/iV5Cs1PeZX
UiF7cO45IaP7j80GYh2wya64bXIy6e+sVU+XJ9zddD+k+FpvRp6MS03HQwE4Z9vn
DHNxUuuQwE61Oicpt7mi0ziEOE88Qi+R5DxZvQvSzkKeAclZChysesU0l+wr78BP
Km7EWB78KqTj2E949umw24tN7F9EiNv5JaqBq6Cl9SBJUKwQ0Q906k1kan4OVx0d
bsBtr0aeSm/erqehFTnA7jc+5uxIfsd0rs4ZsfZA87gGEtbXc1aj5gHTf0JI4DCT
NKtppXy5CuwbLBKCXLszqRXCDNLmY/SlCLyq2FQy2ivJLn/S7vuFz6Fg+9lmgr3H
TRRIywI2r0RkOaToskRvLMps7XvVj6GKiWJd0EJ30gH8PHun1c9cU3/FOEcoRJqI
BsZc0BG8Fq5L7qjmCRigzcGA1cubHXs6/YCg0uaYXIHP5ebdpEUAtKCkkxDQV3hB
r1709QAETR+pByV/4hwBDJRq9KgOiMA4D8RnTFLzieFatJj8WWXg5ImTrmeMpRya
5i2MNquB5a1o/bZJbX76HV6XgbtZY44W5U+VFxEqWeKEGGn59rEU2WgAWIAzwg+I
tMpe+c1AArGSFHr5J7g024lvBQQza6ZS3rbjikr0Bx00/vcCYWlI3jD87XaVUiI+
/oIOGEsD4gObMgrJ4oVo2lLcXbCb8yhRNEA+Rc2wHpyRMuhpvJvkQAA5jS0UHJi9
z1vsSBJDDakmiLyb4ujlH6lA41A7sBPzX+ahfcpETIT0xwxEY551wkAdG1FyVcjk
c3RacJO6gar6Dit46wrM5XkBxanYFEiPHS36gueDWr+rHz3nvndbPEx+AlGt4kxv
ds1zYxzLT79l1XI2PNIpnWnJUy+shYe+XAwbNVnYJQgX1OVaSdekaUb4agxocU5P
EcvYCAjjo4+1wG+HU/ayC05xcEChfz2m40aB42MXaubJe1zghDf8mhs/PNCaLSMC
M2EXndLJ7WV1XppT4PM2HXZOZYPnQw7vjgttxhC2RtIWNV33BK3hmcDgMiBU6E9J
ILd/voetE7xjdeH7bqJ2WayjHbHd4Y4T6P4AqgGNSvvWj2toumjFA9Wy23RRsAaf
/DikchBXys4JjoTrK7MoT+LCrUQ80iu1AMrL9Ot9s5vVmWVa9JuSQtez0lKs9bU8
Tq9K/6sRXjRA0zATEyaQYYrW027Sy/wJWjca9z5TIVCxIA9PnysSuoHbcu0Vib8+
2auGzNg+/n8u5bobVW6PVB8XEtkrNt0ioKdKQz/oDnQ9R+dFS4pUHf7T0C2ZefcW
fTuK0EQ1Zh0zEd/a7lKhRP3fem6MrKxSI8RnLXLW8fiAf4NGP6FBoZMwboGDy5tD
T/CKwp0gPnDvHLqWROGoWEGPigoRCuSTLdTbxxTsAyfoXC8fTKj09IW93EreDofu
UnHvRd22Y1YSakJlHNqsmJClZUHv9b1N0C4xvZO18hyQg22fmGZQpa8KslLOhO+e
gHyOc2Ua5Hg6q+PpMPitu9lJS3iZ296eoRZC0EI32LcCR4elFiNftkw5UtBX5WDc
fasytdIDBWOtIiKVYPXSJm2CDmhqAjuxyLWyhG9zqpLHv0RRxUDk81SrwGj4NN5u
/qXtO8/pPt34OK4UopR8Ng7OkjD8W1t4j4d81NkWLKcd4Ompi/3sdt02vaTr8Pfm
JBg3diDB6wp15Hohxm6vXJoHYJB0Se+4x5Z5G3XtBVoFv9mQq+pQEKPmBJWH+9pq
IxX9TnBfhMLJOuYscFm2J3onKJlSWrlbW1gcP3zhAunFoM2dYCasY00tbKGpu0EB
51NZXG0HH5GVN1CQU2K8u+OqTN+7nuakktgn0XP4DsYWWvRdVfS/vnnWoN/7eQVe
hB8CuC6JPPprEkh3c/2VO56e1mWTJw5eNhkYOdmuS7fG7emCNFlBG4PlFm3d0J9b
RcEbDGPfj0aGb396prp/PzlHyoA/wUwObDQI5kJsBFBSm3vqBYdDs4nnWJdbSv2s
5OfEUPIfRROWNOWxcb0XfvAoCBo1b8n1pULI9KOANJA3gsublso6AsP2WTBUhviF
m8GNONUR7SQ+aoMAAOBk3wZdYK0EQPiDz9XiDN1I6LC7Gid2v9v8IwdcNwOp6JCU
3AexblEDr/Sahj9oCCPY1xLUSe48PmzIEWzAJ7mowReC5yj3GPWbqoqzBFNtLqBm
S/NaGHT2K7hkScJrwmWynIvinxpte/+dgw6TImRKIS66lKNfb+8IWXrTsOoyNWte
vbJHXwa1irmVeNyKNxYdTotXRzyQvOU53YomGdCsHK/uBeAEYXccxm2F1mfMn9qZ
UBUa95srJcsce4goq1sNpDMBQorQm1ONfXq80qDozlYzWiCp/nE5vdF0pgduPGq4
15JFGNb7zatPrtlmnY2c1nK3M2eax8tx5Beymj/xth6V3p5tXRmHZotvtEaMe4ss
H8uzD/4TcNdPAkI8RZRik+vWe26a6DD/UM2ZLTm0BhV87a5QXRmDgg31vAqGDdyz
M3CAo2McDlPanJ29wbhUi+IBU8YdpGigjl2MwyvZboMUvWSdIXwnbpJ2LHllyhqO
FpH2MF2AbgNwNieLlxbXsFSv77qclWeLKSB4XgLwRTIpBov7gx3VDqT30/P1TfNF
zrjNm/qNwkWdNFQMsVi/RQ+SL2R+kTpiXC3igj8wsiQ2k0Tk+BNWhULvZ0wWcF2Q
HVYI90kE6OBKiKdlZxeTTo2g9+dJ3a28KNF7MlAmiPJwZfgQ05mD8z1LrgqO6hQF
/FDKx+moKmNfvwhViLiXMOeVujeDkstkillzEfx2IsrQCqnL6BqJkJmSqTCnRTlz
V/Vb/ScY4vLL9pDXhw7tsZSWzjApBZeymI4Etegtz38F1x6Dp5SSzQMPANicpkfC
U0d5pB3Hk9wI54wBLmGCVWqkFDHOtMG5uxzfzfj9ID5eHEY78oxQ/kYPRQEOqnVK
UNDRI5VS7Xie6D7lR57WC4hEXrchb1uYxVlnx37mUiUem/BGGe/xECSQ3ZXpUd3X
E9wUvm4nNHDz2OnhdBblvov7Xs5EH+Ct54eyq6M6F+zCVWjW/8QaU7kOIf7OBaBP
uDRW5l98rVr4oXWn2Q8Y57mJISkzyZV91bvvpSOtRUxqV0WmnreHhXtTUvpHQaZZ
mxvrVV5J1LBDl9b0mKBR2rIjblf4F1w/OGVnqWjW7MqIAPeqs74v5Xurhgd+CTZl
zz0Lk0XZKfp/6hGOL5XoKhMrHKZ0IEjSKC5ENMbIL9IEdRw7mHxxI1ELzZV3/aCv
CYD7onTHJNa3D43TSCCSjR0qau1JBAJp8h12xzTiNsCR4VLWhJs6WhBtP4gHUOad
C9uvk0vXU1gVsb8DkL+V9oBXEHFeHi1eBgqpuT70s7Q5AvvtYIQrBc4DcG2Kf7tJ
B8x84jEwteqqbCto9l8fycfv96drkH+GUSMb5igC4ltdNHuulRwZ1ZB3tbmgk19V
4qNhKW/+zjiSC4AdjeQK0e0dpgus5rpvxQfRmdmulTwJ6EmSvLEHxdfjKQOr7MCV
bndlwN4wJ+pDf+8mMgcK4+TB+HgMNoouzDi3q047ddECmFW1ZBiDY8r9D3QvMLsa
QJY1N5V8W18OQylo6+cSvqWE0goJrMV7u4llKwN/O0+elWX35FndfKIvt66YOxp/
XLoyDoHZz5dVkhSHz7mT3VSC3pJxrpY906Ib+yngaarMXpbxAgqjW9vLRwLRVk8e
tzx8uh3Eai7zyooDNVbu6OmIuvY9olTAWZgK3Qb8g6lKJ52Xh9/D6fP2aQ4vmJLD
rfJiCpxHAdtGAHzTPxl13tyLHeVyu/P+K1/y/iQ7XnAuoyWlK5LoFbOumE977vQW
UjFtc5E4OJTo0QyrzdWcxIcJ+k2osvmfWdSP5kbi4U5zFV/F0Noh6ep+TCkkIRsn
ahiYA93uYyuTKPXVv/fdm6UPmt1N+gEWgbMaW6Db1aVdseQ3pfvyt50REqvibDa6
rL+MoiE9FnE/RNkEU0lS+E1wcBST9vSBt4JBMdMbmWQJRzc+TwJYk9XAWhRa5U58
25xpc1BJcy01Qy5VVhhF7QH3O1NIeoNw2LpsQDW6AbKzYKlVtIEq/UfBsjofp7lf
rNLa1st5ekqmhWwh0bp89xzB7Ghm3PFbxK+701VLl/O6U5/I7TDnC3WsrfV9AIhN
k1fAKQw6Aj/zQV1gYBbDBMEpmHARUq5OQFNvLkqQqcogmt3dZiyRX453b8nD5Hka
cvwa7H2VfAD9YUXWufkeKMKG0ymI0+6Z+SGuEcmMhZsxMjq5JhfJrp8wwRApi+FL
r+eV19ZZ0Pg361xAoYyjo6ZF1VnY4rSyY8Lnlvs0yVZwMsdbyqa1jBdwk/avep23
s/Dr584JauZ0Wj92mpF+scYYFbvN+eCf/jK9MQGGX7i91JXuCZNoRKeELuKmayxz
rF5B63fO2DNwyw3r1jKN1ft3jWVnkCsTtxMtWFRCbVvhDQsScHm7vTpVq2ZaqpEm
hRrgoJ6J//c2PWfOHJpL1oWKAUiUSLmiUR+xrVCKaWiY400rre2DtVB22aoLP5LH
YUNkj/BzGeTTh9UsfZZ1vhdAViSmF6d1lMMgzwrUxhCzyN7e30tSJr6uAlhxr/7Q
lffrVb6A/MYFRVKhZojJv9oMqeKQMIrkS+yRKsV0dBIlFN7mAYUzTlD4I18hIaX4
km3pIuB/7U+rDNbS0wSyo+1ZtAkq23TzfpwnyM5yqXCUuzWpI8WhMaGqLmV3tJV4
Wj/nxTULnaoNayBn2hmhkOAmJlodTTwCmZzeXHbWN/eBJdnkWmAJ0gNbkZmxWNVz
L5PIMfS3gXCIkXXmudzrvc4+KJKxsWYT6tIEpnv1owx5BSv50Is8FlmZ/NY5NbGu
+0y2G9CEL3y2Mk0R7Q6wnIupYhkf37I091nm/FOVYOYpX5zwYMgy8BjFBPuIfOzQ
dMJ6WfdF7dl1MrXPU2YdezlhRtCdDIbA3bCBPcNnK31Zit90BnXIytTU9Z8QxX+i
d6RBLmHqAxL7w9/Cy3oA5UaJXqfA7mbGtUsHaflFLG6ivN9hFCBzDQ23FnNlCLl/
fUsP2oAKD2/ulc6NzZya8ielLP4fOTUgAP55CRswOBOYn03uNKcUOagcLJb4ti1y
EogtFupKhcE8lO/4c40Y1uuFPFQGyytOmtugMR8+rd0k9rH3lZHz4W2+//KlY7ND
gPiMCvX2PDMuScaboR4D90+au6IzoQyrqnL8CXlHDOhPrybKSVybOz09y6CBO4s2
Iiz4Y6KNvmJ3xd07ODwII8gdCnsulxoWEAR7SpSY51xOL6lZ4DjVwKsMTyiUrBjx
/MWrIOEBnZMsGCf5O3GFekruZK5YkglPf7h1fK8hoQJrOeGpPkeIKHhMb63TW5U2
snzLuw29Ic2qVCCwXPEn4kVupnQztK+Ttmed/3hZ7tSb74amytxtO/fWM06a/vbv
AGxgj5j8dxe76jQHg0lzUUbxJygGNB4jt9j3URXZSxcX7FrR7rngxUsaaNi8C3uC
JPDariumNH7aSG0569rYPyMIrDaF7TBKnPE5lmusVdQrNxAFFD5amf9JUFdSAx7F
kPAEtViUx1B/qn3FEWZUOoZxJWx6JWkP9KI2B/qpDHEfsr2GYl7RRdmsv08y9BB0
7O2c/E9KPmtkKXlpBH/+MIoccpK1XjXzltcLWrhzdB/HlDdqBCppKLCDaAMzgH4A
bEOuJljCGgAm8X2C9WI67AEwQzcziglR3PQtLWrc3ZJSS7fw79cba5p5UScPLV2U
hQ+qgxmExv4UFhJjy7PUr5QWKUTiclSDRFiOfjJPAT7qWsvSdBEOMSFo8jZYp+3z
uit3gLfksG9eUf3hqkk11JEl+c90BEUUBOjqigxZt1y2x2gzfY8/1I8TLq7sporB
Ib8Qv4vpX1fHdH/I6gfiquASTOAomDRobOjvCvmtmU/iPyScrB2u50ScGECoqCSv
x73PVBDZxJRqgoakza0lUw+wByNM3KP4mWtzQVmCTYwFxR6+FrufgOGuC1kJrHQI
R9c48l0SslybWAAg9S22cBiFE/OOWWOVrW9Hr3kFViwbs05QX8MHcOF5mvR2svAx
TqFWZ608nVYt2iqzg3q8IAy1jjsjZqVViPAJTn1qdg0Z0FsP6ZfOhjTGxPD2JdqP
B7tLsJMKFRCvOjzGaFfyYM/Cwzh9gTp/HaAgvJdXH0mZcZMYUQ0oJgPwv2ybZ8e8
TtdybzbFc7b9RxeugxWWBTBaxY9cqXiwL/nWff6FGHRuUU7kGh3HtAfWUATs0dPo
nbEJIHM5UQgIShLJwoMedmeDxOUYeGdKsHsJ3rJZvwHqsC435IiPF0v09miTNJG+
x9MXzVkaTMPlq4IgQZ6mEa94dp96lytWhIfvn/aNjSYzuHN6daOjzFLNOJOH9t9P
/Y4kzwv4oxhqZlvWmD6Ab5SgWaWxMdwqEnpL3JhZpRDHZxKwvDZc3TUMdWNETz6B
a+EbVV+uJw1tVxFn9mPsxfdFAhWpuEW3nYISu3tHP/lQwSE0RPXO6PucES6837XP
kQgkfIncclqDnHZYMxOGa4p8k9RlvrFlOSeLCmhZIklX9B1+xdoutswHpFSnx8gV
JSaO4vZaaM1oa0QRLWTQISx1RfplpXscFTmEcigBWqarkyQn4lzL7ZP7CmksdYEy
mW2tcaXIMXUI4EawtoqvnG96Olv8lvIoc3r3lI+Jc9yxHetQiQt/5SqrVI/csG5W
kWjfcZnuMRVIS0fY+OOzRP0MGx9YhuIJrG2JZV5qIJVVkbKi6sSf/VS15U5++fw/
GucXpxW3A30HTtcBFqpECXW1cCleVstD5usCY4ABaGhtlr1nNda9brjj5vvnEJIv
+m0eb5+p5cPEfnpZX1DJ2kwgXs5BPIjNm9mWqk7E4F4zozOiqnkr/IN+5bLCe6zC
RYfbfAyVtx4E68VClOvpbLcXjQVX9GvAH6mhc/B0SZKU/f8p0Yim4QIltuuNYRDk
cjVbOTnn5yEv2dSJXuPwvHwfYEFrU41u+c+9amH69HluImLWrcfit7FYJz1MrcXm
tsJaFlymGMb3y4b6XUhhir02BVAsmqP0zebm930U+ICpoZ183XChmO/8m/RO4560
NyxM3pnQVK8tnnOKp6yZ2cREyt6NF9n9eo8hWkRjNLUYPVlBswNv0X4HmCHz+fjN
UEo6e9CEFamauHLQeK4wqQ6mNWiR2g0JblxZxRrKjXiHVKotqURrt/3AX/lF49VF
y+6+K3nKILxyJcDPAofSSgdxbeTvgKJsraJyIdycQpsUjLMcYjZcTrR8E0Ea/PW+
cUl2EWr8GVXU4waEzf8jXtVOQL+2Us7uyytBRzAuy82Yj0oWQRTXRU0yFVSptVxV
5OYEV6v//IYSiYotoOuctsbuf7Tb2aty+KzQthwTKHLymtJGu3+DM73K0D7T9eBB
Kpc0EZojPlYvEy2Qu0U+Q+4CYYDYE8nZC8onfTdN10zZJmlDNK4mOV8t3va5hboS
gl82Wc5OTeZ3k423MUE4TT/7ohu4n2q9w4mc/0119896LLDq9Xv6uf64eiPiB3uJ
4vNidqr5WvjQZpEDjuKr9sz7EjSjb/lkvqGuC4mLt7tGTmSTHODPT91A/PEvF0OA
N4pX6N8z3juSoQQ65PzQjDp1Tskuvb51hFqJGtDbdNEWTaIvC4RWWXvLzR6Z4yd3
Kbfp0FrUmT44V759MRNAgkvoS+vIGaSvSrYSLUZ4Kqv7Xx/EB45M1CYmll7uGI+C
XHj8P9eDSzU6imz1FGDieW1LrO/c/ZmynF8eGGIYMzWwDDRXf+ise+cKsGNn0zGj
CVvkMMlmJMm8rmVxzQPUCb/Fxb2XLxtBdQuVZOKbIiLu9DFP1B+PVg/mkY5Iv6dD
cOMKPi/jy82QRhURY9NTGbdzdHVIJgW9+LE+XxgLJ7yUY0N9A1R1KSvmoz38gB9m
/yADiUWRiWatNcoKIABeOQFcsHRGUtG/x59la/BGKVBTgyH9L9RwFUHgoju0B8a9
qVqyeC7WL99tAo/3+qqSvTY4FneFK05LsOdPJMoa56AXEJTinISPkUDiKT8Kb01p
EtEdF15HD0k7ScFpf6rh3qtCoS6SACqAK9sFN2URG70FcgQ3BkBsenIGeEe+Y5Sm
kHluxMuKlLr4GL2F88tqni4/jp/zwXES7g4oxee5yG3L8Be2WdlPLyPquxW+whMx
rkftZoriKX3+9aSRu352MggGHXTVQ1kygAejPfAwLswaHvxqhjE06p2pW0aCb/mP
nl81Zr2E6y1IlH2/9i9Yk7GmmErpFUcN2U9oow2s2aKz2d1EnLWXv4cf4H176Yhb
eRa47bcnGy85+5hPWRVaQEc6NDhpQojuAiz8ylQXKluG809hbqTLvLaAs//1zIJ4
QgMwKDXEYUhr9tWKFrHJ69uRxbMq7/Qr4AARQie33beLW+8/fKQF4dtDrRenCkT6
nQMlO+HGnk9fnW2UILVJd/TZzPppwLFYlHQ3M+IeVud86pAaHwkoT6Xc4MS9u//x
peh1ps+cXmRq2eUKT/itbMtA7Sb/LzFSSzQ/wpB4pFyjdKwmphmFG52EzcgfdjAm
7j7RsZXUhqB9gWkw4ypCjpIZQRi6i/Ic+XLoLIWG3+UxCHOrnY7XxwkLW/t0KiiS
TlzcBpdN8v3bg7lhqBJej2oJzcEwyCrFofmSrCT1oB+xzG9eTJvFz5BHqqaimX8G
ede6pqarQOZyh+8r3M5VOs7iXH6Xc9J0Wf75Zd1qyBlCb4qjFPIkEpRnXR0CGDk7
5+X7/ADtlY5TGmp4JHHgwvq81GvP3ruGNqgGj3ZBthJxZjQgb8rSidwRK/3fff0y
kczb7P+mXZEn92q94Zen/WMf/jyFSvX6xxk6csqQcesezXkR79wI9K9pM9yNBZpv
4cO56AUK5PCej3Y0oWUIuiXuMkSKrPIglcelYC20QPrbB++jCfTRb/CtDrO0q92P
AA8baSP8IJhv8bvn2o2od5CyYcE4qJwIgEhAik35DnwY8z6bTK/s3fyV2JREoSEm
JclGPHLqTf/gR8HwH8wetxOdNTx+vj4cKWTbMO0jAwnSM+VHEK5PXxv8Q5nQGYdG
3sWoKtol0peU/eIKCig7ixkxY2vfGAUlt5W1otnYJULa2IzHDSluc532ledFeSMh
Mutz76F8yHEAMpXj+pOzQL6F3zHV0vOEhAhh2ah0xcFWsyzx5KG3wornaFxiyEYG
2ESJY5YOz1Cenp6NdS8YUO8zMj5YBnKdrcDuNzOA6ODeayQ16rjolEYZxHXEfoEK
wfXyk/xp5XV6gStLoQT7iaqQZfLBgc3zRWjubDh5jEcqn6SKKGwCLQhoHktYVvR/
UFYN11xTEvKDkt7KRyRjxXde03SKb1T4ABgM3F7lohi0OqejzTk+eukKLbylXGlr
fT4tuCd3O1/4l0j4bi9gu1SkL0YyFQK0WZ7yKYLg9M9xT2ulXucRT0ITGEJOoyC5
HWAo7LafSQkhwT/6ybmatsASepVziHg8WYFQEmNpXPY8ryBMRf3cWuguYsjax9rr
Oy2Qe7xRwk8B/j9pnweyq6jxCxZQ0aTIwPtcNhWK0C6LaXtw1x/HSA/oftAFswoF
EI/4Go0xkbRR9HTdfSRABmZ5/hx8Z+cpVyeU0Pwpbeg1puR+i2g42psNHCD+4On9
/VLRQs9fDxqCAV3xFQxMIuOjT8jOMRViNvodVKy/AbHZuHa5wIcaLRyPWydH5XZ7
n2ZKV9nY+PpETxHahI1IiIrNS0L/EGQVLLpki/p+3WpFDWxnbXUR6Y6niz5i2ezU
G8PA8DjvwnkcmE+9UY0hbnimSEDyucX8smaDMczQEg36LL6Q0ctkatrlPhjRGNx8
xBGoS+YWhsYoyZCEuRmdjGIZzlZG4uIKh32fCnis8MVlwtefCXc3JPI/srYrBwLP
1YdeiJc3NU7GDRIXkzugncKyMf0DDjyi5Ybu5nskqZz6c45ESk9/bKu0BA8X1V5A
oN05fXZA5TWLsjGDtv9EIP9iYGcSNsL0hot9cNSiAgCanvWo2GXjyBB+3yP+LfB7
zYn7aNkXJxSlkBJJKmT1T3FCdDbMHxWhaqg6AA65k9Qhje02ja6N8JPyFTmavqLC
IpH6KabVw5QDun9RFKyAxP+MxFaTzH/pOloA9g1C4pxPXuMjymefexY7NTf5s7xM
xgykLCMT1dnXV+4pCVcRwhQ75rJjzwAJpwyFkS6sFjgNktaqilOO4H2OR/oy3BK7
0oYL9TP/LAa6tZEldXwqaB3780ia70m4roDli3tf9UTGAae6BPksTJ7Y0r2dXz4g
kCBhGvIgniMFGlvjbeehoszdugpLPiz0ALEmb7BAkEQlYLY41SwuemH+5Eax58sB
acU2JzDEBd0mzDjChGk3OiJ8hx39zBzMz9PiKhJl7Oe3tIpcBSpuJJIncCPhS6kV
/5kut1hBd01reNi1tI4bfg/qfJyqis6+x9AJE+6SnLt78vFO0yD4oJpMes3fQhV1
WAErxrp+IVjahYEvGlYFQ8VWf897zdcejdX5OfZR1h/mqwI9R3zX7BikVJabusLG
sfAMye1v10pze3rmswSbdL6AitzsA3QbAqDliaR1srx3eC2+LPlUxSS7KTgevBCn
TA7LBX4CUescDkcpiY1DQRJnsAOlhpNRSQJEOkN9di7Jprnair5U1AU15OBStnrY
CmcYkHBhFbN7DI+lbF+tEvrepPPTox5iad+cl6R+wAotzKRtcN40CAn+vPQzYWZh
Lrrokv3LzvwNCneQohYPf6mZGN8LNZy8cxyVePAx3UtVLxod1miwv+5kSc5nDhA4
nawGQG1y/PYO7964PWcr6R8EIHRlX0CRPz6g7w3LeY4NuHWvOIEpV4DMZJXbf3Yf
TjzOsgeRmcdbKlnC7eUnAC7EIxZx8pxGhA2x9njAFJ2BLufIDwlo6WN2XWXMdDVI
fmXhBiJXVkponbz4upWIYhcnSOrQm0i9qgFTL6mJ1b00apHrBGrIhkHXkIFI058E
8uma8xzoMMmKb1qdhmTj+2vJEJEp5t0A9qdEnhxLzLmpXeT08hBZjEsOR0eEOKiL
GF7nhY7Wqr56TE7tldpN9J6B+QpHCmXL308U919nj/eMDpbv09ydSZegNYVjGeG8
Dido6uSrUPM4QodOSclDZKvQGfR614RkqEkB6+Sra7IXeVXMCy836AZ6Lr7DovRc
O42qcGUqqTJC/AWk2SzBeFfKbiFtY8LsDDg/gAHRA8dJt+qglQVwZohjsISQyLoA
maAuDJFeTiNQikBuY9q2I0vkaXFMA1CnzFe7QhivvIoRsplRMz6PX2oirOkhuPx+
BcdSsjzImyh67cLAvMGdnaH2e8mykJVuO1z6XrXhQITS9nsnb715A66p63Plk99u
DScNXcTa+Mc9tvWIkTET0zJxw8o9xX7eyavEtSZ5j6AT6oKf1xxQ5GOLhkPuKDz4
S3gbYGp5zw2xzlZmS146mVaN1tS9SCUHLb6Wfadu1aZupPVNtpQpBxLvg0dWpUK0
7UUrQb/lU9JpKcC+Yl75yCewWrY4CNpVu08ZIdSYhxmGzbIzSd6rK+Q9wIO2M0fG
ElAOpuaaxOqICqyksSGpMg5CDESM74efWa4A33ACueJEjvvxIyszl/Z+PePd/lKr
f8pRdI8D7vIIkSsOwbp9dMQzGiAqo36Qin10I9535lm/syCFBAUtLbaMpJ+LcENW
i3lXZN3dtFFV8YNOFQOVD11BI+jmKAR7WcZcLbeB/CLGwDhja1ivLHGAebHz6Cst
9WDyc9vDtaJXhp6c/Mp5UZADMSu8d0G0Z2ZqR7IgGhrk+nTVxAZ/8QOikjLoe/fw
kF4Wdfu63Ure90VZj2DhVnKaoGwYnpghXY2iOIsxiLDt0TdQWHVlbv4rTE0RjSC1
wn8GHfUP2347zxqf12Uqsbp5YEPvFM0safuDFP/eLTBtBtxgkCqvq1RugN4OSDlJ
QhuVCGP+BRml+372L2iP8ZfZsg+bKNe25Dv7PZYUvqJWaEEzKKCWWuQXEnRsINYY
bPVzn7nOpf6pHQqa0RIDsQ7OHqauFdc0RIvG7bpbbW4Ow89F0AnsgeRn6i0XraYg
+GmAjimXhWaEFNTic7d2+XGU8+x82eonRrVc0viH8eqAU03mGhQRS6Lfy/NadHrv
XFcW4vXS1yCG72mbIo8ZYfVIMwmpi04a3865Vti9r8UD/3Qpv7vWzWZrgq2QDADU
o9RIVlnSId+hj3TBWhOUJD8A99/wrJVt0E2+JeunJln5CbCS3EtXiczY/YseiMlt
xsHaKNvZhqjQ2jIj5D9GLYezG5WpXO2YIpqmswbbmJQHUUjO/O7fzKsKb+viR7Q4
ellwYH4k49UeLIeJBk06crdYHTW86v2jqun+lVYrLCgheHpKdB/aUyww24UZgBIN
10GPXbuCMlS6eL5jKoaBqRroek26ZT8a2PXLSws4UdY+rvCw9oT+XDmz9hKXWQ5i
7MOwQHYVy3fLrluxWEJBSBmmAIM1r1eeJr61gGzwOBAnyHeY3LQsKM9gDlZAq+W0
BEN3EQWJ1uZAeSt8fIsS2mImrL08hVrCk5SyqyKUJQy3+uJeeyUjIVXnJLk19SH4
bwNjmEUxKQ0L/gWMrlDJWFO4vhjwR4chxcgb9L/+5xaE0TqQs8EQDJ2JhECVxvX1
Bv307s3z8FfNZIQxVlHee1//fXHIDMsTRES5j6qblsXmTrYPGM0kxHE/3yBoq7DG
+7rslogLWgXCfIV/VFHXDvl875aKsBH/wyTx89NptkFPuyHI9NclZESyJTl6+w1O
+Z0bRnulWOCSnuDcRxIpojny4D7K/7d3X76ucV1jd+pIquNRF8k7QCQLlldA7/v7
INgWRu+gYQG26w7tltYaky5JQCcA3CVR6EoqsG2GfZsQFVn9xcuyinHyK4UIF9V+
uUVm+Z8cCf2mmhvYgQ5YKTpDoIV6JXASlbqalW+dLOS/K5VZUiL6ic5jNS9BsCvs
q0224dn8Vj/x7WbqiKWovg+ulo9h8QFQeM5iRCGDnt62McIq0R1rRYUIiyN0gA1L
tlOd6LKbyZfcZetapx0ygP4Bo7pG9JW1uFD0/JRRdPrh5/uQ3Pj29NuH86LMls8e
hWqYfG13YB/oWVUhL+7Osdm7on8y2Yx51IWBAOgOvx4tphb/URxkLJmshyxHZBXT
cIm2C3Jh36BDkPVt1GvX4W6XvTVvf8T4WjBgn+kgLUu6rtSUXDipbDNtZlZ6JZm/
1Ch6wO+5AkfVyPm8y2HkoQk9KVKLtSlphli9dgkx5jBMsLkyTV9NY33zAC+We30W
8BEVj5jV3B8mgsKNUWwsSNn6Okrq+dtqlSDKhTcXQ96//yDyf+cPwtRf98LcT+Mp
isoZCs+7zE977IUAKeqfDu9tF/6Nr2EXbXraiqoBEModzfwyQYacDqK9O8Aw8crf
bL1zyU4NKEVlqzFDfEKqI1hBeJ+nvR71oYYi6hHnBJT5nJ6o5LyeYADurHSe2F3o
isb40SNnRlHt3WKGrtN7JUFsM74s6SXWxlXwLiUST+IoKK8AU2WO0OEOlvbge0Cx
CpPTLcWFsrpEg8CZqHaOtBM+OIPntyiDJjjwbnb7zhcVEnerp+h6oaXyfQpSg8mq
RNl/cGaRn0XF2F7BH0o1JKDsP0TQK97w7DMPdDTQFxEgZr3UfWtk72u9q7OZ8GcQ
+klp1IdIQAwKsxRxIEypul5BihcjcWlu4xUoQU0x3dKRPaxTbIJ6ZW4o3833JWda
l2OZ1zlQWl1aWakVniUu+7zR5cY2MphDOAHuysmuphX2rwnbB3lqxrtINT+Tp9eE
KFE5NCONXDus221vfZKyHIoc/lUvKGGn9f42GnFV57+g5dRUj4Tu34UKdYh1Mta6
4JTuIgGS45t+viYTcql2ywGBXEwT4SKkUnc9UeIXRh0tH2NrFHucR2OfnMgmo13F
TwWHBlAFtq1Un1iZicCmn1BRYhfvjvsr5qZdbPTTIeDVzZ72Jw72laeEn8RQWnks
8xnCzdTwXqdhQpu7qZBoJJr9hivURlxkmnBIYaElEaknjjC7DSBhaYd+fOQ7Gwxh
LZaoa/15zFQvz9tNaIyiG+eig9WqQRy3VWJfbCgf/kZLzS/0oDJ/YMC0r4UK4A7B
O4fWNCcI1dVM5F6CCwCExyWRa7iz3kxd13BfGg106v7ygqU5prgO+nOL+iz0pf2D
KvrNwnJTWfRP+EzfUoeWTPI92k755OqYgbqCLpH/zqLMmmTEx0LyuPOIVnxBQMD3
OdHTDYD22404MBzsIds97Uv2ngJjY7ZMOzOFdx89S1p4b8kWi2UEpF+n+GF69kIT
urUhzG12io865QPUCKur+XmBRoKmH1GpPOwKBKxfeMJsc4albUIni6U7LXji1Ck4
LyB92YUc658y7EfAOpuTB9Ax31Xe3nflvUdZkMF6VwmQOkpzr7TKyZ8gitAkeqPx
pFlj3s2+zkAEyxTZHhpoyN0fqkhO2q+p2nq79e1BOWemG957QHtzi4/8esWJ0DJm
quEZkRjcm3cfzMmK5W7vhwMjKKVlAj6ZXg/hT9WeGrnsc35MfpsHCYPti13iNlpU
4K86lqPHENjYEwsjZ7nSbygrBhU5YnklJlCrhoTBIlwzbv0BPBoSaXpvpdkmQUzC
pola3I5vxORNqUZeH9/lgPlq5IB0/i7DPgIim1wR6j0i8RRVMb3Zus7V9ixIAKzP
qhQc3Yehgfiw9HtIO/m8glL0cZGXE5iS0TX4kGIfhg+aS8XbMttXbQ8PocjEKbDL
AQmeH2WH6Hw6B0kkPj1E5zQkhYJfer7dlFWdY28PQO+S+dfLlSLcWyIScCwx3tbW
R9xolpGl7omdg6yFeTQRYlkGQiAV2kLHK1Y6mJdCYC3+MJ/lckMcqnnTK3kNX5U0
R8nTd7V/Ze3GdklP6wxR30gntRGhYZg9GGK8YC3WHkH1WvuaAgof+FbJva57NG5q
wd8GcZNSxI23MV4KmwsvKSiwFPHNeaLAQf7LHvAWgKSrqINhC4ZIuKC/Hh56F/1U
Mdwy8y2jYJvrCcfArwAFmmIpgccvixIxk3fMWqkFyBlkYblI4m72balPgdzdfC+p
uYGK9sGhZinZBk/nPuN01lWaMYSk8Uz0cgSg/NdLqdXQQ3umynbCj5uRBGJQ3XFA
/1zmqJ2HmtogLqUG3L4dK1p91TfcV63bXj25CwoTQZSqnczpilxi1nfNorL7b/vA
HYqNicYU65GW9snbH6c7B77XLMHL+fMpwh6pnMyDhjcJBenWGyEU6FPhm91Y7RWO
hV6zhjTUuOE+EDUd3vTYaKgjmqNgu+fSefZZgQMf+m9s3V4bcbJ9A4kvcKPUab9h
4181UV6gU643N7nyWH6SJkGnfv2UBd6NxqjQ9VLVcanJxxDx4zCt2MyTb1nDAoKk
2y59caSaVrZDGGv9pTTFpwASFuxC4Y3sqi1etb650eSGc+eairsYJ+3Y8WTRNUz0
gIuJGwtpA8F+TQII39XgUgwSsEQncQTMGndiVRqGUy1L9ZatvvV/qiKa5uS/m5GE
OyoGUrTabJKqTgf1Tck0elfrveej8uE9/EJIxMJ3ID/I3qNcxrR7EVJbYQAEIXP8
sn/j9yj33JnbzHRVcTZEG51ZoYeOyY9kmpY7dfUQ0fhSPAP3OktwT+srlggzqIMA
UdlVkHlvEGb2PaleWHCrNi136FW4jRuPg2iiDaRDCWK0ibV0yxuRwzXaevBNviSG
/10sGyWW8hNrT9nvUxGF4FJdOQP5NG1Z5OPEmW09d5yDX+YHAk29bGP+H468nov5
tr/fUKlE+RzSs3FE4YOlARwaCvQCV/iyP5V+iQkvkC//ByoBya2t1yXev2hut5up
F32m3p+E/Dxp0Bq2dPJfKhzrysuBZ5mztrCPzjC+ZhAUKyldxDXIh3ZzhH8liA0i
M0rhItgOm180/tKKOfKmWgT91hG9Gw397fIuNGLtXNJyNscQ4WdyUB7mrS6euS+z
ux/DXVBZ2+RFXP9r/hPQD8hFSNYNyDJ2EpCKtpDJH2VrOTnPuXQ8o3yrpgSSApaB
x1cDzfX2qaRLROWjKFGIjY0SLGCsxzVdq0ybUbCnBc7fobHfdAA5i6ei0n/Zl9YZ
QEQnJFbqwk8tPvIhpwB7LpnohWXhangAl/CJduqTCC+J6YXYwaX45INPcv7sV/uT
8A9hkCgWaonceEH1UWyMktr023cUjaza+omIdrpZonDYy/jaDKkXTz2cJCsKImsE
7mWWnXck7jG0vSyxOmC0doPvNjIxulwtAa1OaIowB4HJicSYXLrB/I9ez6CVdHLB
TU1LyPGvy6yVAgieWcTFkuwPcfm0P/YoLOQGF9Kb1cJbdLyIgEIHeZjXVZ32wRK9
oVFLCDMlVsQ0Zy+7O7DNZNkijyc0ytAjXznpgzLuKGJUWms8XfXEWBr5n1ki0/Sb
fWImQHhdGIE8BQFo7YWjMKMBudXWzYns0qc90IAyR7kJ+tIjkWq1nJF/7UgKCLUi
gKEJRTATFmwjnSj2SFusWiFtRBvLqMW2S99ImFnmJTukmz47rVlvwseLVPfk+fhr
JAEYVioDUjs/18wBUd4ZPw63qqeVYhENu0jIM7U4acnIQaZc0EUlK3FHnxE8g9bw
bGcWYlEQYT/a1tLmndk/cvOeAWjownGf15p3OADtpS+uPdMSHKiezhz0KseMZ2EO
BdTjPQFZuQE2F4iJxs4S2pkmtkzYvkxUsigBlCh7VTV7qpf4CtdilmhIblxyDqA+
32D4QOjIqmRdWvwn0UfByLzLByMsWs8cGWcp77B9k4v2UECOhxnW9ggg3CHdPkiA
DHq5fNepJ5KzKDZoZG025AtPsctWhJo2z0FZqr8hmzWwIf+7bxwLS1VItDokwel7
Malsv6dm+Mje3Tx1FaaKNlQPc+nPMlksx9H71WD3/xNylLBAX7EzLUBXi6SC15u3
Cz7hWcorwpzXCUpDE5XMl1mud5cTz63A0nrlgXb8511cKXwcsumrURh327koGvvi
TwX0XNgpH90nOEH6lVnhwTaqa7GQfyk15n8L9nWc8/gKJ7wAdPcL+4bdOHNG8b5W
9OCwxen7Bsj0EMZSccpqRCRfhsXMzu8qsdH+0pi/415MW2C247Ju4zm1TFqlYKw+
EOnm4Osp7kv/zd4ECRX4AVCr+f4jOP2+yztdTmRjzh0phsI/kfhKQE+0RX6yzUxg
1kaL82jiMVNqzs9E7VYncYObfM69zFRiq8/DS64sRXU7vk1ZcPRac+T6kXP2/ld5
LN9vRs73mrSJDflTatD+5YTEdO54jATY1+VWE6RhpzbZ/K6M6K7pevR6/Zct1oy4
JKUO7+kCpvP4GnIqHzj0/HoSMY4pbdLocxUZ/qu8fzFbsCRX9GqLdRG4bTj2H4/r
crsf3zQKzQsNsZdXTWZejlGTZwoD1vK13Jv1PgqUQU9bUjtaXWpJmHsqdyTwqX7a
DbdFbOfBGUytuUVWw5KkLGwddBGCRJcXy3d7NwXrY4dMXP+CGGZht4CynTGh2Dqd
HB071GB+gtlYjbf5qrp4O15flHN+HE1J/97xbG3xy+qnnzvKc7eFidEZpv6qZJsV
He4PRKAG6z0GlE3mb+Sa3M62v4Zed3IKiX2cW9wqRsUHFKtjYanhUS1LvLzTCeI9
df/iSIgLYvRQrz+Dc/yQHFjQeOBauhHcmwSswaS1RJ6mdiyziH5uDOHgvrgQsj+u
vKVYZyWyNZ28s5m7fSVp6VSqGl1x6Ag1PQTVZD9IrxLroTFv7eKGpud+vz/77Tfs
NMeCIl8hMd2zqycCP1dhDw75stJvQyykpH19D3LBwBEAoMy/0vUd5DWZYcV2PzVB
biaqXT7ZslQJw4A5/lnsqq0hjGiHhd4HdNR/mwc13tzGQS70OZaqat/wBEKxhni/
AgqIodcMrTkY0KiHBC+P8CM6faBgFUah+4oP+zVtyiBETqyO3MAalRwEXu4D4pIk
iMppRJ5cELjQkRhGBgbFp43DM+Eeh0oKTVhZCFdM3ETD/9CPax2w25pMvFF+MBvb
HPwsfYB5p9uYj3aTFEFreFHPMa8aEvc63wn3QFA/KU1aOq+gfsoVH/kd3rPccM1D
dWSDOo3ommTCZhUK/imKrvXoMsXvJtlOv/Q1tSYv2Fus+jxZHLxkIPEBzW2ddk4S
3Tc6rZmuwZYv8SvGV3Pmy5eQ3CuqNUwrGwORkVQee+w9wUjaxmLW2wOG9eR3dnqT
xH8trkHQMF4rrXZnUKEkrSrhzj15LN9Z3Ja8ySouLW+Lynb3uqTAolTy+EKxG7Q5
xWXu1CQOMIGInJOk8fVdol58b+Ed7mq9j6smNxAQn4NpCWHkjrA+wn+cBWvNruUE
aQylfc0EIZztOZOeFjZgMrA9rNGZdEOFX6itmYZ3ebC8LWWj8t2Sv1/znxh7PfsS
EMyR/Hy1McWEJcaQ4znfQZp2ZVo3zXzbLZaN9SViIF63QGKfnYb8Y8XxMNliWHCb
ff2qBew5qXZIMa+F1NLsioteOVcLyaZK9KZT3GC5bRRIHSqaOXDrOHa9W1EwZOsz
NnRkpvX8fSkfVmsWun0RcJpQaIWtdk7F1wlt655FMLzrbj9pXF+Vl6gON8ItWyqH
jb8ylVAO3PKnWar2LyPbV08M8TC2LmlrEtXqVvbjyWJU4urH6h8RXd9SMZBdbzOn
IA1bU1C4gu+eXl7xYGqMkKv5Pf2LNx6Nu2W6GsVb/h0BI+2dCUBw/N59KqNnKakY
AJJJgnYttAyx6/edrLv0dH9r/T4jRaT93BDMfrEcNMZtq+Xsh5Ub6WSNG7FywVab
ynL52S7FFb9FbWkg3+z4gUiUmaNgxPjyRl0R7edfyYtbcLpcAVq5yA/iBzAT63Lx
lZ+jXGhjtYONr5RIyIZfd3D0rpNq9Sedo396GVbrxJloUs/nmaJnOp5iiXZ5qZLz
Pal/Xa/pHBIJsGlkGocxofsDPE4GjdemEMDt8nU0hJ8ixCmt7iO7UUOcnu/5zC0Z
mkfaUtIg704XlOBUDPp163PaAygTJirUZhVawa6r3ZKbK6n6xvd4pvuzomaq1Y6A
+RejmV67s8Ej7qY7rw7yyDkvR7jJhCWfOTjPGbhJ/t5Al3ggBe4qVbFtxBw5hrCi
XKG2VdqYX+KNB06LJNT2gVhyG1Kw7s1Vo6cvNDqiYlOwTAGxVet/jqm48rizDAj0
1alHSOMrZxw+FJ48SAe0fuNa3enfeEexlNdnU5ZNdssoaoH3x5wMJ778t6sexC8F
DiDKjuHpCWanId8KZ4hBChyO5EedoQ6AhF1zMCgZH46UHNfIe5Cwk02gHVFM5SAE
BtJU2l1PnDoce6NsEYB8xset2P/1MQKsYukRAM3hGsum8dk9sQp2l+l4aA17uawR
YmFFBg1gixCidvov5dd2nO0iMXrlTMRMUSg4sjk+pXo6zavwxEQCdftb8xPRDART
JNCQj/pDTW94jb+0PTT+FV2OxMq4zpsDhYQaMD8Cfz3GPavCKqFlzWERLbP/VN56
FvFv1YgkVTlMNRM1YkdQZMAF6P0dBhglzi5sJQ0bAWlSgSw4STkCnn/PKXt59Sin
VRLo7UN5CsJ+yls45PxyDKMleOgfr7/2DHUKTs7HBE9cEQY18R99gpcBz6ZvU0ps
MihoVQVXW3IaTvcjdT24YTC0GT3w1LUE4jW6A/M2MvdgxJOhuSJCbdkJzF8U3mcy
yoChsdz7yj90VEwWzFbb/U9laDEAWut/GlXeJVph+KhKs/3x16T8/4QLPDfjgVJO
aa+S6Zf9veS+yLFsqxXxWo9XGyX6kXByNnsRFNpHK+Ls1aHwL+qfGxKQ9GheIQje
R+5W+JJ10RjheQHJg6AvBpYn++TU9iBvacaxDgFOCTb5MPv6H69MiJ326YNtK1Ho
UzSpkxTwWAdolWS/RUiaJdG5x1POhthYpzblMCoRYJKNV3VVhGS8jj1yp66mvwBp
/Di8+t65VSXN5KfeHSBgJ/2lwjQ21gqT/zVLovwxXui2V+WiUPWJr4hNK7XdQriA
tePdaiLYEosQ4QfzeHM/ROp2ziU9m+9G57aifQWc/abLj0/uEYxt6cplNmpGzOXV
WfEWLmyqRwKA6qTjbvILE2phAIXpjZ/p2GvCxr3kkp58MTO1kTBmzt3UuV0OMip4
vXgBwpzBMlprFtBp8x+tW57lqPmMI0q/zMCK+36WDwCAI4k09TL4nP4W2otjH9NK
+9hcjHfrsjrP7d/LAF3Bq2LhJKVKsyO1ed06PzjM64/KTsxKVUFJISxSMAyTkser
XiKNT8kClpacX4kjDknHd26WSqxm9YtW0Ko2YDWyYQzYtIbntFRsPF7WyFbQVeHr
cy3zNpKRieYvUGrt3nOvKnBAxhjKfArIWbODkPp2KPT2RbcN0TKmZiU3C/e3bo2D
7aIwkODk+mI6d7mDEEU07bmPNiHyv7qVlhlGr2omS+fJSxNompebx0PFmBPRnHst
5q2YbAaJrMz79VbWJvoF6WRTe8apRxAXOlbJC0PuCDj2xpzFL1/BQPoWhN0+JiI4
1b/qM2b+JNJdFGVCCYKI/50RchLrQXFNCDtJ9UXtBL8xBynto6EaljCpPh0eWB4H
W1dTZQl/sTJgDOC/pTVwqf2FyH1a7BiRC2vYTV4bo4924hTXRxGOIdM6sw2eINyB
5PmTmLJnoKsDhxotMxZWPnatV+I9P8tvt1DLbEK7hIyeeOnKUlDP8FKlYGCbCGII
V1YfjB/zFgQMt/ZV5LQnD85rP0IxnObyxKgBhLZTeGSNFRK0fWpP/sKLr8WdBG6c
9qBTnzXJZecdQAGxA1iApIe3AWuBg7fbZoaEF8H4aJhs0uHLJmPV4ItX7ns25PWA
06Q2IyJBVK3+ilEzN/0MKNTlaKYAz2ayRastgPsXjNmb/sk/l6bQIul6YKSkyh/8
RJledUQwKCrtYFK29MGHbJNCLOJgY6G4euu8HEAz/MuJ89PPbOR9/ImomMh1Wqcf
uS+mvus1GcW7R4egdc6IQbQLEILSH2q6LsHXIYxrCtlncl/2Due9GLgqhQe5jb7M
qOgWLG05xEekB/rOHdtPZVW1wXmijlfXG6e4CAeFjdqO21JDHcTeQugrilFDfkns
kg8YxAt6xhGKYoDbJdsC2YztvESZezlArV1qvvN7NGhYKKKdQe39ab8Ey4/B9KlA
Qwcj98fasLYwvLORqBTrYPl4ThEV1E1J2ketKiXSQwpTfdLTAp84yKWmgBHIcKfX
ogUDRc2w/pEOvguskUzZ65EXGUFRdRqDbfYFv4yHnR0rYaFJx7kD0sy7PGn/oICJ
FYNZzWs+SEzC/R1HF0pd0qQdZpj0SoVX/JYyWDgkLvZwLYuWHVdQnwwcmUjRfiPo
JR7cri/DIBU+OBIZHeX29g5/UxKTqpK1XuxVHpaFA+BwLkWKA9VDs/TemzZ7fuM+
qVxaz3WeAY5Y9yi0DljxasnDjqBQb/DiodwTx2AWmN6ou7H8Sc1mEPdIBhW/hZDd
mDYCpD+HgD6XySeWtvtSiMFWIxVkbMcdftQIFitiBSKdIKDBBHC5Q7oDZNCTN0la
0cMSie6CmM1s0XxXZbHwCJ4Po1tLFV+UcfjKShSrvW99RswdVcDDgnwq+WEWakFA
AuWKDodJXomv/fcbgp54Ju0dhpuPbxA224NJgJ+29aTtUESHnhhBYfw2jka4FRK7
8JI2TrU2r0nef23kYenTo0KFx4Y8WiowOjyvINuOQsJ3Q7lNFV6hQBUwsIEV8mdU
kFKX951UdqGoBA4xhqPmv6IF+ycGwkIRQx+7SvFzZGQxoIwtngYdftYmfIBKnGlS
bbYYCZqiZjZKDYweBORSX/XWRIt3XXPV0zvWsSHYh2xCB9vMDbHuEpChSWYmNJCC
Ug4ctisZSlNKnL+erJDaalzNc8YtqiTU8tPGGzLZCb1nAdb/EZ+6nvCbduiBAeWp
/aHuLdP7VuwVtMP7OZeuXIaLpqsECe/WQcKbzt/757aobsb+hYv1RzIzAX9Vc3HH
hhzvIedylUpCHc1K0S6W+Mkdb/jEzFamOYQ4pmTLTuq9TYOb7bhUtYitK/xha1dS
IHuqzoFVfHofkPr4p+ygAFtvAo5AlKJgkyRIl26/urgIF2avd8OPyjmEFk1VR5oH
5y/P72WEtPelwrdOGdoDlxy2XLIcm5AjeFbUClOxAQR6KeDnFIm9QOivAL6pMx2S
Wr4mCl707W8TndYBxGPkqZRawStJSfce29dpl5ZIfjm2FVL6/U+YEcyBcVOD5ylP
3ftqQKQb3+l/vQEGMAb5F5VoJyf95pj6OUJS3Vz1PRaoGiNx1DXlwG9Uw7B3XdUP
I1B5QVE0i0931FcrLPWlIswn2QwR6wyzbbVodVd8ha/tWnqcVCUVSgOXZB8qRK37
p+9LebHiDmoYY0wA+m03fWLsrXrCbXHxCYdBW8YZ+ui9OwVaSuJFPPMuOzWPuLqX
FBFs+M5rluGlXWm546XoxHPhyr2QJhgqV5ldwErELjnvTdc2LMRnneJgstVEhxTj
S+nkx9m8jdwUFEJxOq327ELDwzVnO9whNYZnGq1CZKdxfOkLAvy7WPQJ7qRX2MM+
xYHYK8gleOIqIajNbK/dp2FPZhGYrh3b6GpQgvx1sB07OM+qFduXCPBYLqOFfXuB
tn2K2pWfUJso9/cBHVyBq3Gg8G1I2tcPin1mchGs9reinhaRblroNl2kk5Yw+6MD
6A7zHkPlbvrswZXeazAxCuMa2Gugeu5ar9GJNHveZoUXtGnN8atU9K/QZNjDSLio
PckcdC4EV8zmTZJup7kyle9QT+ftqR+9PVT+nOeAyI2EGIjAsh7Yu91zhM+Q5u1k
q3rvZzfD5jzHDwNGAOKl+hOEFs7TEuKJ8u5Hue1NSiz/drxBGTz4sGuLAnCIMD1v
ZQGe7ANI26UAjwggakUfRXZg+6iNlC2e7OBeWuqGyp//rUsiZiWwdW46TfHnSHdp
FAqTgYzKKz464rpERDGi2EwFWeXt72DPtBetAumxteRh2LH/E5f4ezvVJNAbA3wq
hOSgnPPno61yrWa7El4sb3Fo4d8DgmgppG3HFf/p0THQ2wjBbCwVfjCFDmuHFwpb
P7h4ACGBaPGiOuJWSrXdYL4ELWFZTWCvF2+viGCaEjlvGabfjFz+4QrU0LcpI+ab
9olrEOm/B4426H2qRz8LgSUywdQ20Lb+V4sz5fytJl2wpqviPBExabNwTiq2lZ29
pFNKkNkwsVc9f+DsByRViyCBlmvBWkw/UNW+A7KtKkdS1qVnx++U5Mq3kwTaD5hv
dhv3UOM5EbzhKWnjQ6SmuYpVP4Rw3VqUFbP0MBK4XhkbiMe+fqO01tTbci+t3X8l
ooXU3K1pGwU3vb4+qBG3jShFCv5ZYwwWkh1ds6gvDzuLprvllmKivELqwi8oCXCj
57aOS0sfw88d3Spp0eRo8xGSlnLxab6iWDY49BHfnWFEM+CocAumfmBfOVy+QKIz
13ElmJVmJA/rKWnf4aa0y1fUOuwk2r8sxvrkGPTZujxnWqTBF/4tVCLnMmLnQ/R2
Gqd+U5P1K8VMSLO1VKGamvwUbMx63H1Z1IDnIwSOIjNR0VkInyBnN4DyxO3WqGO8
4DlrhDewQhMgqC0NScLtJzlB1cmvdLKCrY3ZnG/NAIzgQoJ6l0S//8an5unNKzSk
FsfnXrL0pGciiUVlChfFm2hE4E/IlExyExe76grZpI3S19OC4tk7ctGMIggBvj8Z
DrFsa5GTwFAibBHVocGnvTpSWq9rwColzbU9Zh17rZ3WHqDZfjxmnZNo/SDnkxdX
UfwkQnZFHt2vnw51jQwekO5PLwpVPvt9NVBAi5a5PckX5BJwFkZetx3lbeWwf1mP
5l+IPPq5LJzVEttov8v+niJzXs5Wz8NnXk9qfLkoq/JpDW/6fbo9HOhoIjsQHP5u
T5HXEVFeGdsnNkZvsCmKvcB+q0+GKTGCfwJtlS9Vkf/2Q/Xti6COWr4FVpTj0P0B
T2Rh/GkREel8isjQnB11b6pU7Mw6kp5+QuKQDvu8F89WaXQe+VNFzoJFEMHkJfxA
I+0IQ+Cc2s3AEZYRulbZeDTOGyeQKgm36k00usFZgmZyHkBPnpKbOjheLS3LMmbp
AlXLvPTOsOoTjrPYJHujaCwK8zxuWN++g1WlA54CQISaTdDWHMH+91j3SQ/+xxna
5y4F95qxPAJUZzUtZvnm06MHUETERR5bM9E1LjVNPdfL6SZK3sMI9MjJo1PxxBgS
SjFhzf1E23M8CjH1Pep+/VzGsoDFGT7+XBpGCkvvkmDxnCTmC6tzORpvlFCHIXN1
xo5rhR/WTJ8+CpPt8fv/XM2hWBsJdo0FqQb2QB1EQNniDULcVtGg5uqf0s9OXpeG
UIpAtU+8osh8tkA0wH+xeZ+5Y587/VNEs9KWV79utJHDbGqnh5SbWM/lo3xhfCOf
+O3T6G1DWKvvLw3ATQiSDhDbcwGK7mIYwjJS16YKJgZqDmya2JwUObPp5u9b1h56
vAhKWEMULJKW2oRWLG66NlX6NekjQFbKW50PUI11PW1KeJUCeTAnmzDuPwciRz7U
/LXifUrPQYw48YVeO73aXyhiweKl4mCb4UvGk/JRop4/2kYMrzP6v3sYZrsqcSP+
eT/H75bibWRcioYjyNh0pVvvwT7yjiOTHLoDhPPBW5v4cyCR2A6zgNzJ4eWdLXKm
fISb3so9rB6NVFKzcbtuCu4L3bonFeY7ql2opEoOkwg3hAGtyH3vNWkkbiTFyJoJ
wAM/tsV/kKi4FtSS5CULnxtGJeZQuwAN0B9G9dfFSge1hhvuAUniAxj9tbfAdpqz
nABzl883lyMhpMNQnt/DsnDMviheZXBdtKNFL+ZcB7Ch4eyxmjKf+jVhUnuTBF7i
Gxba5+R444XA8AESWOfbR/M7A7IaIhO5+bdWB7xfeNqqKz2KDMSTTRXCdVNBYR1j
m5aLapABRR6mJXz1XwSYNk0qqwLZE3/ijgRm1ntYIEO6tSNNsO7hsKLejm3XIoQN
mlw7QSfUpTQ0SKAWCuBaAtMpg3C7RZWWKCsh2JKkFzSIkJoOiC6zwGb62KKGXDO8
aX7lRmxxNaycxuwfNyFnUFlV/mAOe7phLUxlEjO9+MbH3bLeugWw6dD0QiIPthqN
Y3+LKKBmzFt3zyLk6wz4rdyytNonNGAnUNXwnUQwpZkyaqyIRg2FPfM413i91MWk
iIUZTWQ+7CN/ZjkfOMQCRbKRHRoHRJDCkyBWiYQjMAAMJDx4aShCRt7QpXNPO80n
l77krPZMKuumtjM1D0wmHdf/jwIg5TICYmx0DCwn0N1r+7OSxlfJ88oUQrxOyikm
uXbdBw1KD4NA1YfA1Muc+v6wDCUmGcOQCaAvX4UgmZ/6qg8LvIb1fkTFCF1i7gin
6Mv+DmWNLDa6PoLHhcWP5LQn0GWmxTff7E1TY00ifNgqdrSo1gcwSQuF4nCf63qz
3aMnbY0zv6iWss+UZSFi0dXa6JYzuQhAnQmbH/wh6ceMOPZ+D5TIN11xIoI0hzFZ
+9tp3Ehj0zM/ef1ZIv0yvndgdHpvKpA/FD1B/AVFEYKN3nPfDicr/xoi18KmLhZC
HsD1Bxf5Ll5MHGnd38d7tBteVeCixHRRFZufQgN8drnKD2G3IlWOX0np1QvuNw5R
0ZZl5S4Yy2FAq/1SY9gM4c5pnWtX2wOI2VzTB2+RrxTLD4z1qYJXar80MeHwkZNG
+5xazkU6sLyj4lNbuGIZLj0g0UU0OUnjG6PFEG4RC2WR4Y3HhXpX1TJP348LMh/3
rtGN3LH5w0ljZ/EauX9VoBKt5/RieXgmZBvQBoxTln8exi1yW5BlCVBOXqGnQFp8
F0YHfOjEIqEfS+2IN+ovRbxsvoc0jZNud3gd7ddbiLSsBIB3CXYiE6n+ZdvMLJ5D
IN8AArt7cSmBojJHq+YJqq/ZdcEYBTGxvUQ/I8BJQ0Geube44s775+0cgUfEHrqe
4ANTV6Duw+++Dbmyb69xpiKIeFzjaKgqaOZ5OOtkeQk1jGyI8xJS4TVZQJXqHn7v
bVuup8c7LLL5vP/Nisv9SL0Kbf3ocm/P0v7J/j9eD4LF1lbbsmvO6WdCp8is0F1d
JausQXMkA5nsDkP1h3cyyj6ENU7uNPSUEtfVa6Bjp8xFWa5GzFwA7tSqE2PUGZXA
0bi5U8/jnU1Cg34ofQe2LtYakqs6o0qtweut7ALufyVHcja9/QvxNRVx48oq5Ojd
YiMTL2sf8QfynqLo7qRACdH9gOaCfXCFUVVSDw0AFhrQCbojQKEpoY3PY4GtabHi
mM+bjUcr4XmQB2duuuHyummnHjJCGEINgwSrWiSUyMe1fmzhHKd+2pP0o6ROQ6SE
xJP/lpqVOQ2Rf7jck5O6m6kZVljf95dRzLYLkTaE+szsrGCa+pUOZzDiSQUvKGbh
EIfbwca1iLVraOIhzyVopHe7osVeArK+U77Rpsagc19lezYnygKyInd9PRU1Xe8J
inCZ/A0WDNkh+edg6IvlFvMkHt8QZdpBa4ssXbKodkoEqbFcefXQOrLO+xJtD0hs
T8WI3IhvoOrPzc3MffKLiJN+fsESoCGB2X+m1gBuPPTOa7YSVsONQm7HJUHx+WP8
aHnapDwTgUbDa4E38xgxCLVGZToP92alEVcd5DYbBu8CWMbqt9cYGJoSxUQsJ+T5
/hG7f7L211ELXaQ2FHwPxc3+M2SeJEtmVW2KdgM9SyrgqtlzqMAx2m4aCyDwMbZr
NRUjgMPoa/ii2S2MiKudGRWCSP9EZvyvn31ZGUB7EgCvT9LzpqxP2qG3Q5/cKLHG
cA1N7/GSK1hcPSc3cOrrifVKjuZ9DFj1i73tQVD3IuuJHEvJEoMnxR6UGp/G9lyj
kH7fU8fZ+tcpGcpfxf9m+c39BW8hwp8vBtOTaewCE0W6p0KHtSV29o9h0UHdVo07
Atp3b5mQWCdjTeM8vwbsIIQY/ob6jCmJAisF8RjezGIg2yO7PL/0h8yTt2K7CHoI
jyJle72S9ZeOhUklC6eVEduubHzztQC1JAXWqvgrpsnoylIUbE2Alt4pEn/yAqcP
5PjhiQ6bCkue78wkwTqJ3pkgePopzFxn+i2hUp5GyBP9DoD46fytZwrwC/xczDb7
EjX2K8+YMD/HzoFmwEbFwE4LlxCqutcj/IeKrTR2bNcW3SpG0SWbHYITMFEJZhzy
3uLeo2ttrOQ4oXY+lJ1sRv21idw+1TCX0r2yVXee3tpz2O2KErwg06tb4L96/4cj
3Z8reuD3+ZKlDlopF0fwtLpLYjJjRFL/syYxsA5lXcUgcCl7T90gbGG+zQU+spG4
FZuWfeu/y551dYBhUFv77iBzjwAKRbKKJMDSxA9q49q+5L/fCThoqvRCnrK4jBLs
2j31Y6wltGZ4vSSK/7qTrmajYncrOIy9jyAmkbaV07Lh8cHwWwym0kpO2/icnRl4
IYaEbobcATmvLnUM3TQgbbWPTnV09mkwaUAoF9PsaAj+DPkGDhuKzNZ6k0AlhicN
LQLnEYw3Y9BndZTZMK1GU3kyDo9sqzDPTbNjBM8KjWPGauOnPxwRwoviujWRZZDZ
QiTQnDrUZEZyUssmXOfGGTHikc5/+JRdJDYq4Ge7cScrs8edaoZ91uuV8SAW7+TW
S7eNTvGxnCjR8odFp3nm2IQPaoGHe+Qz7BHRrOIE9hc24Os7kncl2lCiL/WKBmFV
kUvfnX96rZyJpjlzwis/hQEHqWlTmcP8fcQO0iU5s8yIMwU06y+e27ksT9P/lFG8
1zFLIBq6i6Cnlfmz/wNCgVFBB0+YPve5hst1gjuC2WtsfUMcyrL6RuHAxo9o2ORZ
HXryg0llpqQbIM5lGFYFnfJStAFvjgme8buZ8v1lsOstkyFg3mEa1ZlCLQXZTM1a
o7TF0njCbiECPFOKl8GkGa34eq93Ah6xt1huj/0Ut8wjAVPJKoVNd0dIy1oQNTKz
ZDkPNOgaXSdoRE+fnpxslrZ/mWyFfXszMaemg01RAyNqn++KdDMbPZP9YwKFRO4d
Mmb5qc4Rp99wy+QFRg/Uc9ONwgDrKOPuVanqno9R9EXNz4w6vYOup/fwvcK0fUVa
JpLqLflg9nm1uZqDS8+WUMxWNzI6Xy7ULHgehts6O1sHYYehqUFTwTYeCO6dcMHd
hEFjqlCoWNTR9ZiOLydUS1MpgOwIzkccwE7N/Mvmhp+b0qXPTvjW2IsXjkcJR31R
ubplMCtg7pAxCo36cZjl2FhwYUr0rklMdaBmpECeBOf61otI5wtl4jp/Vm7BurLU
iVYrLBaXzUJPfLfSN4w0WlheyCzbYr93r7gSxrXjGRWZp3zdeCJNodtLxF9hyHoy
JwTBzzGxozEnzYlZXOuKoanrm6rtVRjrIDMauQ3bySYBGZdY2ZMtucePyRZqqSEm
uRazDD62Br2f+s0GVVjLlwQ6sQSFtgwQSgbooU9uBQjcAFlF82NZ4UprXuzRoRMu
BIg/ZG4CjPqtuOsliQFFkhNlsuCZafpWETbecoGulhUP6bv7QvZ3l7hV5FKu9stl
bA5nQkpZtHFxyjvR8tiKsstE1S6e7o0xqTZWk/A6E7C8E8d9P9JrMK7W/uAGXQbQ
CPYJox8vJJdQ0DNUM1RE27Zpbi43nU+wGD5e/beME1GuGq8nV0V1wdakq9txZipj
uzc/Os7sQ47qbVA+VXZF6wmRnYxXM6LxPQ10BN5mjGMIQ5oQfYOyq80WI6DP7bJs
QZEhO18EA7EuHA4HDXkCsD0pBimh12UKcqM/WgfOvJOjLz6eF781vFa0EFXkwQs6
e9e90FkdyqXqzheqR0MTmzD54WlqGAvd52PtrkH/aFIhWGLV1p4c7UHnOBupu0eH
ny49wFkZiPnhI/fBMthloMG23ZomYrSDG2UTE1U0I0VdC7i9A2go1YTVB0QPplxb
6ocS/1Q+G1Sb1at9K7GVs2thKwSCwaqpAfvk2JQAIsW8CNKEt50bREE9jlBlkzy0
MO+BH3qT9xyhy4f82WZ+UPmmv1PUxVig7oJsnJiuv814KgB0sXSa6eg+6RpvVmq4
FVmtHbLksiYu6z4i4ZcxvT7YsJnyZXaXMrraHwyuVRsaQeZGPh0rzc9SQSpcYu1y
7BzDeu3SVA4NBHRg8JoMpaNLE8WpPAB+faChQUjj3ILmE8yVcnBsxAb0NrpBmS37
Uq9xKGLjopB417se875xmiaaGGj4urxHmDHrUtnwr/5oiTaUkJPqM2LljXMS+AE4
PVURoIRIGRDB7m5wktSCaomjWdqfStPG+6z6dHqYxX7wFU1CSmItwyvu204YM96g
R4v7N2G1xNvFNXH51Fs05Fjz9nb8+kSbmc6zP0mQIHlmGnAayo5SSSCUzynMUATS
rubvUdCVk3rx0sBIfllDIXOnBXkdBnp3h+89m2+zNvEeTbbs+4a767JNbUtQVfbC
trxu3pG0twcwMR19xq/RJ8L0URyoyubCBlSgCcDjar0DMHkTGaMTe5e6aFLbd5KD
hTucwehNnwV04+xSYRh+CjrL/YefrL4FDS2W+WQszyfnKqT9AhDWKmCdp2IYHbT6
1tHiTTga1KisYnl/DSIGxvk17Oa3KHMBe1ZCOWASxt6HCAMsZoZx5J0slQPJ2D1i
4HOAzouDbg4qgI4jHyFno9aqM00euIACRhcQDyxcvM78wimREYLv3pL8jsVkhHez
Q2PzhJW64QARNB0L8cYH86rpnAZsuG5hb3aXz7zWiutsBCHYnlGPZowSridjcUxK
gzfNmKMo3aAdFRrSUlZ9On0IEQ7mul0mSiJTPDL9sGsr83wVD3WO1QBrkOwqocC9
JeC5VZshWujzmLIZ0CQLJR6eO5J9sn2Zy8uu1IZmn1XKh0GP10oF5ttYZ0bKlAyt
oEvaUTHZJuXDN/34idDpLzZmGu1WGQ4dmACI/xquTLLfh+rUSRPVKYwLvt02+edc
YanZ2Q5X6hVRy7me6M2fpWifanLzuS+GDe0bBC/Z+q3OEjN45/dNmS14WDLsSb/u
OGLUczyUD7ldcHQLhKy4UB8K7lO2mxoZYaQZRT30l29gucxsouO5hx9lm/UQO5Na
BKcX6cI5y6ORSsjEgPtzsitDU56vnlG2Ud8lqmqPOSvERM46jauaP+lrS7kRW4QQ
tRyekUAuldG1yppT43JUj/psbBxjDLqo/VkgZFdHsDyPd5F7dcOE0X/vIeErvacl
y17tvYfXLkmmfMB3L/7tEtEo9VV59Q6M0yS0g/guI/LE4B2M4TPO94lexWFRtwzA
MLjajWeUumbxkiEEVo/M5DIA8aKEnMfKh6BfAKMvjun7UiB49dZnC2zso4fPrVLK
9Y5hOtP6hw/XvPi/34kZnD0cKuPNiLhTPezfgJl6w/nHCD0YMglp3HMJNXLoPIYr
RSXo6EnAkGMt7zDqdLbMKft9MMQa8lSDw0NccsF6qbDrSRnhj9wOODPMWViCj/tI
uVXYAKqkwtV1RmG9qiZP4ioik0YgYTLN8Icwtt7D25n3O8ZkBnu5LVu+F1o0XDwE
cNc6jpdX0UkfVFlSEJ5QXuR1TROWV4WaeH9KNN4xcL4cWkOxO1IE7bfHcvYsq+Sj
VFhaaEnSmCpZ07JFxiUwIQzjLM/xZ8Wd34zvS8gY/Pii7QtIVZWmslo4662bE4cp
V9GgUg9W4HOWTsA9aLKa6wCTQtHgCZ/0MBM5LrSDFqgeFuPlUeSHqy575mtBbn0w
U3Dn2MpotWuBV+w7x35wqWcPnJub83d/W4ZgJqzRVzE1b0rYT/frrVs+9FcxUAFD
VdFwuIy9p9E/YPbmpeEbniInuG70exnqfeA0bHWwN96g2MPk8AVFhZl4KHdeRrRi
j1DiL8pAsfwwkeLFmWPSJ5IMjAlhasNbjjOCq7DI0nXNpxT1fCDIxi44p/U5O+UD
Q3/07A10O5RfOj6qjFIPM89hCE5m/XYdqaEPNJBpiRcgUSErPfuiRjktTtE6DNus
Nd5zbXwCEPSchOahVBq95fIS14RUw4tMaQsCUc4lkvTSYy5TTmEVgezxan/e/ahL
FHi4MAFs5ZjNOmwyXIBgSffTiOJzpaP9buXLkQap29FtiMJu57WNc0yvafHULvOd
aOFxtLjUIEfUsuB1jGvit9xZ3WiyrLx9iu/Rp8czW8QqjXdFWjFlaHAa9wtDJa51
Pee6vE/fv/sYnXmw5ZYv5JAb5KHaxkAFHZnZjuwIDVZuOhXOE5EwDwbT2xgvoyFm
cZDS2r7GK1QBPqkzNH5aJxrPeQ2g8Y2qNsDKdmmrzmFVutGxUlifm9qwwmM5ziLC
73GOlcIK4pKO4ihw6ZB98lWXVMZQkGirU1cdoapMVYMD8hJW38B/BGJ6ZEM5vOxI
XoqyoTCGksfbyIf+sPBXNNxdL5wRcGacNNLmUy4mWwjQOrLfVvU9i06d5oc1ZqcH
0rBFF3mVkyPvPTVlOV3qbOMC3y0kfTPQVNM2Yud5uJMRtgIE9fg3RByPtiAqOJMM
ulw3pklhVXUwtCDaT3yHFkIOdOu9uxj5maJTbdPWbseRf4CgQg9aFdJJMng0NVZE
LbS4ZTjalQrjHBW+7dSqRcOkrMMI4+dDPmFXy8ot50+pZpHeqUxYyaW4JpUAM5wJ
Si149CnYOzf+weUpF9sg4iv8ZUfaC+CypGhUNd727mvwyXRKTMoMUSXBZ2GHDA6Z
JXgh4Hntma8E37P06hFeHbrng19br7KMsZg5CYa1YdNFd79KH0DkawAkdRYUY2Qh
+XbiP9qaGJveGmrckLnLcDrSDihbvNMcEIMZkYfMwUrEOFXH367jAGd7Cxvh1jAA
ey5vfOPb76WuKELz79XK6f/CVmimaOMY9/eN9Iu/liVJJqMqaIMZUmQPzW+jqdS3
A0AH9ceEhxI72mfmcioqt/BYwAb6AbEXdUFjZ9uNL5S9F3GVVRZaR7WiiN61F7q1
vtTS572BR2LNBYsva2I8OIEqzyub1w5Obz6pZCPASygxpUoNnbuD9BO0z5bXJRMz
URyPtRBw7a1CO1Ns7ytH7F+vm373SXNTcVV4QZQJq+LN/xF/IoG30EmSAUV02ide
nIB+NymXzFeJC/Rmi7ffwuhgd23Jf9rVvOOkl48yROKOf39EePPK4d+VWG+yVTe0
PzozjQb742S0MW6BMKtvHrJRell2gwKFhANmYGutzIOjJ60HYMwcLuTEkhC5zzHA
mpaEMnMvN0LHPXZMQtI0yWNjabnDG0jQ6U8d3YSILL+OyLk10yLA1LUmdDHvUZNe
oywdJMt0YGqSaZzKniG6yhr9475r+WVJ4fpXDd/1Ceje3L/pbkJ8J68Xle4Qj3ti
JouZ3/vcWVkpc31ugRMlm2HyU42M8f2RCwLkog+bIfuqzLG2/MPRdOoQXO6+1oTD
03rkvIhuTvWz6v+V1fzxTQGFldEXnengnbJbv0uNn3ZXJyHZSYWc2kkIJFLS08xB
1QA84MhCHIkMr5FW667PRYQCtsELMvZVLbXDjN1lOnr/d4KmynpY9jACpnmkRjFq
aQ+7pVYt7I5stjtFEnJ4QvImM2nytuz1U02KlniUxiqZ4/6CcyKE5mA+8XO28202
IhB7vMmpbZLbF1+ZIArZQIZFucZ5IA8kHaeQfcN+b3wl3MLaCYm3j+qE+jwV0kQd
AHPRYx04mVI5r537pIkhSpK2sKBa4QNLQhFflCg5c3bK8+ymnyMNnm3fydPE4SkC
tL5MDMXJqwRFkYCpz0kdHKLQ0Rpp3S6i/9bK0Qu8783okhGJ0eBNCts2u3FbO43S
Rl1giqbQI0x52uIO0E2H3spQFZf5AFqh6AscdWnFtZAkOUJyoCiiz4gP47n7n3Kf
W6WY+WXU8aIcELpFMCJcr34uHbqKHmPz8s5b/x2lM2m7LvNiRVlXMT4Gz9Lui0PN
JQptGf6IHstOgvhAdCZnmkU8P6JcTkC83walVBfd+U7slSnQByixf3djuq062gjw
FZc6jRgLg0q0u1gtIZPvkO1Siozx93SkVvLetFnHwHUl9qljU3bOLMt4wLzD+iPH
B63pxr9roBCQCsprJU0qVWFBtCq3hq6StC7xiA9JvFEWTpzhXZJYgffFUdK3L582
mXzKTcB48nxdkQUSAFkLjczIAkWV5R4gb8fn30LhDgq56otOLucdUkyY2D95jxbq
yCD6ZXMNT3XQxcdrRfG/dZaNLTuOXvAAfJni8RVABPZXkrQ33a8IX4KSMzb2bR8u
lbdynJ7K+B4L04Eq4S6wilE+5b3Su8XW2Dd8Ax8OGQ0jmF7zVRwT5x28yTWE6YEQ
thUx0qir5M3DdVGHCGxVk6OGb6iGU3ndNCYX7AvMRrnOL7vycCLOXgLH9s5mG6Xg
CSH6nqlqpU3mY0kIMU8AQgZTqS9Q1l7+wgxkCzNy+Eej9qksOmVaUsjhfn5MRJkw
zTd0xWLFxRpCy2ahxcAYi0woEww13JpEMV9fcTH/NcHbB1y2djhQKlhb7eL+v1lr
iSG2hkfuh0565m+tDdmeJlquk0AXWeXDDDH33NV0QvojafIgCCXlyxZWfQDqfcTS
A9hToGfSjWLV7h8j9onkebwfOS7DYqybETH/WNpQwDGkUBvSwWh2MLIDULGabD65
O34fl0I1ku6RoUgtUaFObqBoQbHhhFXIkVicc/xvSGvEaTGpUlCyGFanH0vXnd2p
+Tww4DdW+jMn+eaZI/gffw4d30mha8uiLPchwXVFD59LB+SvzdkTeOjRzg8b9uR2
rs/jIqMmtwqZzcoYjUo4pMfV3mSky30/HWouod9nk+E506KIs/OblP+TVNAgaBL/
7P7uYJJSO0AmMvVSpbwpsamGB+GsiKi6Npf0lyft0/JdFrDqwDFVge6IDMM5GEY2
v+DSFcmz2Txn0OQe5PpIOvSuMeQGyn0VqYnWaLEnI0MZ4oRS0ZifYHOVLMZcQ/VG
gS/2EatG3n+yYUKcCXcrrjJ8307W+ehOR4wh/vONcoyWDy7aDGraRXcqxHZZMBlr
hCKwseTHbR0d+1UsyAWNi/roiwbp4TqyC2SiE8dhFW9ldNFZnqofTuJdzOeZZw+Z
HNRuQh/CT8uyJ30E/srC5P624NdQTmcooK+06cZMEYfEcr1XZRk95Z9u9LiJ4r3m
wXjSLwsYuneBD+aiUlv3NdH7naPhZ/ZbM8hgoOx9k8K9cmRoNdLePqd9fLtNN3N8
33k0w6a1nY/ICVecIcTo+uuCVZRT837N8BwBbsBjjNEFOhllIrSY3D6YxAe2DnfG
CrLastza1TMWVV1XGFJdP4/3Rk7NG96ohrWJQk1YsfnSPc5zGW/n55RsnzoIHRIf
mIujuXdXlo9AH+hcN4gTCBrf2CHyEY6MSw4TJBIUyHPVB8NbcMJW5p7gdau9saIS
l9R/eCAWxc9cxadK3f3+tK2dfQGB1kiJgIBw5VGXSWZz7+iTIc00DHeaqTfuXZfU
Et8be76sa/00XUIwM+m5S6wizKrGcZ0Ak8xNIZ4aB8I5GXsuQdGMU2T5sgZm85xJ
bx4l92nTqfeS/vIu2qv2mimuYRjnAvs8X99p9Jkc8+L9h/X2sr/ebaJg7tgUREhQ
psI2Bn+/5jiCSOy5dREiTU76vIOLDptt8ETWaff0lGPMXEOu0wFYDdwjAkGzS3rc
Aaj988Dw78MX1mLfSj4M/BnZI14RAE+SvTmPEzDTmlz6+Hw15hg+7Qmx2KnUOuCN
yyzC2u7cnZLU3NVGO0tfH2h8jUHd5uHAZxZbNZYd5xmpcVGUuSM8tjnMWBISAy03
rXFYd8fAgWkcwerlQbpUxyRZGdg8FUF+eR2HyO1S54BBKSCiHA1h6jGCppx9q7Ay
Df/fbMxwgMVMKwTBQNpnMixfYit7S/DJemJmq+YKYnZLHpag15NplUJyZYlKf/+t
qO/aqUyeYmJYCSRSSnlKE25OEBV+mRGcNyciWY4mqs8jP5Wmzx68H6+F07C69DA2
0UtAGPINS4I1NEJ1Z527R2DDJrU5FqBbBkW4DBw4TeBstCWaPG1YenLyOTfEiSBE
/jK/IHsVBPiCPVpILy3i1gTUdjrA9lt+AqKXYiGvSmGKMRUmINNoUXbTsh9Tgix7
SJRezklvGJklXw2K6SYSon0lUGojzFDa1CAHh92UTYQZzccp0EeEoFxwaLJVUJWS
JtworGgkD9kzNp+92oLPQNdSOQsYM4kYwYGNk4k3wxnJUfjB3wH0PlgruUCTi7ZH
wMEb45Gznp58atP0L/xKAgANxHiBNzpTg5NdiHoLZil2G5P8YpF6OUklrzrYkZX8
92abFqO1tF/7lH3pqHr9NVMEmCB+jL6ggWhlowg1yRvK9w2s9s6rhe34cB5VZvxq
zk+UAwqsfFBSdTAud4HMj0Bcp17IZmDOP3GudR2j7Aqy80K8w8NwVUYwQomn349h
RKBjaACwAmmNRUxRGY6mBu90dQzYqM38H2B808iu1BhkDqPp4zYFZFJQJhcBwGnY
WckXmdwtp/SuDvm1EDQOSI0mi8drMXk6+ICEA4h3x9AqxvvqMxCEq6E4hfARfth0
VPa8eIxjUKmH4DR7newHfv3EhFYMG+pSKs9mTcf/Gyo3VwT9qQi5uPh9SasOpJWg
iaZkXmYAOGA4/2npMh7Hu5wzQYeCbf6kQV9aQJ5ElE2spqs6zwwqP3PFRvSjYICh
YG7GTCZ88t8Swon92vVTUne80zSuFK3BP1ronFJs/zwka5jFP/AQ97VGIaQbzWBt
0RBn9FJyQeCmjvXX04tqkJndk+cml31DVZKgMD0KNLLvSz3piFwAoH5/bD9vIrNl
0bzzwLxSBLEzaDS2b2iwyjarsOftSvIAUjg2IkocgpTBRPp0CQpDem+j2jOB4ael
WgK2hXJdO3TRssj2KxAiTvQOKs1awmPfiqD0QNooH/IlbjSoeCxtfZvjf7cHNdBt
h/MMQJi47X4uoZGMgeE7t4GhPBRNjM/8VlS1VKra6DsHggokgd8z36FmOOYbfjEj
Nl2nP+dqAYYRgvfbF7HKh56lvoAYnEXYDispWAFZAPWZV76K17CsUd9PM/UuOPdt
a1DBwDTMSCMEx5FlPnPh6jBGv2ihCPcd/RN5UvMPnrr0oM9B5rgOyc9sDWPx3bvJ
aTHWhGxAwVybzTeWjQrYSdY8C8zv3++FmrSCanlKk34d666knGN/grWKC6/kLgmn
4zMaOSBu6qvyZVkpoX2+cxI5z6oyIIJhqX9aRyVUDZ+kGuLisjvq0uUWlX4XBYPz
7OrfxONnkK8MT3xq/MLuuTANalEHv09dy6IcUjpkAMK1AkZB4nsN1ozM3BhOG4MV
YoZM3z81nsBUbGOh6AtVpIRwHDEr8TD5K7XYsnqqA9ABkvFcsPcSG7eGb/AEBnE1
WpHuFY6bQ/J0UkvTOyNBTrWkiPsewu6O2nK773lTGQDYib82OPc10C4ocwRZh8zt
w3sWe4+e/TBPqwYnI5j2VbmbjfVctlO9qvYacIs00RbxPCmDWHjwHxBFfcWkn236
3pHoZghf+3/ozFt+a2rwm8P2pmx0Ra+iO5UHQ4Ukb6ztlCMjkjNwxESdy0vOafid
T+v4zaGQ1jVYEYsA/YWRLyaveoWHTwyIsEvT6NpgA6/ycxWcclNongIP2e+jYN7t
GQ+ebF4QRvFgWxiypJuoOL8D5+aqykVqBOGfa4uLlSrn0wnJAxRyhEFpeho2wylH
vT3w/D03q6XXmItJDM/aJwnPr072ARaAgwuKrbeSo8YF4GRpkoecih0nOFGYzR7/
CGUfWgD1/aYBlfM9/z0WZ7Kw+6IGArZG4ZMKMQFg3HIgHKO8tyR3r8T/6BL7fdjF
Ir/tytyVCFyRqIScPRdhr2hzMvHOPonTQyHBS5X2oGoxRe6osQGRvzMUX59RLSLJ
d3AvgT3ejthnpWyBFTekZcCKe+A6LDRlvnSI/OTklA9Ct2Oyxf5lA1wBVvGeROoE
LapEtjEndGN0yW76v7bi6rkYCOxoePLcUCP/+9ftjjx1ZV7bC4wngo1KX8skiKzF
HVAnSvWj9JxW5u+4AM9AjF5z+aq9XzBXGXnhoC74IsG8EOnDmkW2qJHKHAzAwSkg
nO2k0lsYA5QyyJVv08l7quVfJvUHXPYr9dx1vsNlFoV9Zxc2D6aZp7bSFVOj6ojI
84jfC7si1JMEEwqj009/xdUT5GzCFm2Ss2MhDUTufkgQI9i4IeZ1Wh6vvvWHHU64
Z4OMRrCZGVXCiH6fnb5cXb8ygjCYlSG7/qlb3mPk55vkJi7RlKV4Kw1P6yM1J1zG
nypxgmv2WMmReq00Z3By6pRfF0co+hezl+xS3l/XFd0DRjQIH761mdQclNJw32hV
lYrq271n61jl57zK2Z0YZniEYUo1SyWz7xUDL0SxpK3KYPRTA5LZZfIdpjBhGhQU
v2hoyjzR3dS3/D8R97Mw9Wu3ZBQXwMeg6mGTNWXya9WX4EfiBkV/xVLjJD1lqhDV
64xBJEsc1hucnRbIQ5P80V5B7otMRggz8M4yqwmVpqBDCxS/WTc3GKsTyJh9x4ch
j88CRtv2meHlicULB+8yuG0Cyvr44Q1Jt+Jww4UipNVoQAZ+u6cuc4W83gOCTPmK
NqoW9QHB6mLxfQ7OX+3uVoFGRr+6uY75Ll8TEdAe+dT2seylhnkXJOPshzugOVRu
9iiGaUi2N1LRPnqJWJuJJe5l4+g1znPowWWOlB0U6x2svUVWP6me9FhcKi7zrgUH
Hs8B69By08kt6V+zTqJGv4RM+FeMp8ou4GNRLdkOWSGv0C3zhFf5dhEAmIbf3hGK
+MORtfhAoWcTanQ1tgBekTuNTAa5gus3mTBJCufFLGp3aOhP9BONcfgPqmkcQJGG
gs/ClEXuvOturu4a0lqIksUmHtqXsBOZthw0p0SMDo3CF9soJ7J2IclG/QY5O4Oq
VU2ey+el1X1rY0xpYbeEDNZN4yirdpXJGJXW/SHaH0VHvel6ASQQwyNUJCe/oL0C
ZMPxZV8HZRG6xld4BtZ2bNAwYIWdIB5Rv493ruZlgfRXqoaCqNZP0h/O78dO7jnl
KgG24EzTEWZVvIGcTcFc/gZqnklzYwrq6nWfMMXA+7RkgZ4KnPM6QDRVC/GBJ316
u2sE9CYOBnU/0CQsGKNkMGvpdyjhdGiEiWqqsuvrwaX4836vuyXegL8TeWlSaB5d
deCF75YalyZbsTAkz85iGA3+oOQu1QtcWzDwirwyJcUaYAgbjWnf0kF64M7zAFFA
5/dZyY778Z9xejjV3cXg1TU+GD9G1s8jqsLPMvyHXuNUlSGeZbtvvM2Y2+dLFvEJ
fn463bWfNhVM1FIB0dhyIV2ObKlX9zo61wOE5IHLk32QB1a6NDiI7/4jNiAP+x6F
xc9cmi4OufvL5/gOIwGVylSgQIXNRwSt74e+DUVjrrrsFjTL90epH4kgyl4lMPQ1
kZT5+AQ5n6U/0V87wC84KNYI8+wjn+n8pIG5NfNob5Jwx+iWinM42L2FcUXTIlOO
fp8qZG8cZ6mIvf2kXbxlDq0+gUUuSb1vrAqFR/0dLaYk5b2kkC5GZr6xG2wpVu/s
oZJMterF6G8ph4Fr6JFa5LUw5WIQZhH5eUlg8ZRqv327+ykLYXEzKQpnPjjOzuM1
zwHQtqqidzTlJgY8JAsMjtDvcKQOr/hr3SsF10PY0Fx4KZLtzevr5QRbirMLQRjz
5C7zXJu/yR0gVMOXUb+CeHciN9lB0q3cZYnPHZdFrK5nQKkz10R5YexgtkgvkLzx
L6Z9Iatbr9eZ+ZJmCtuoiST3ONamZrKA4d3nFi5/UvpGXeQnuUL/W5VwnNOZ0PVV
T88Db2zs92iOUuCuprWpVnW3BuJbYqArfchipK8uCkH0C6y8sCW2kfOb5INlgWGv
fyRKH6+bwVmgSKvmElnG2pJZx84xnQiyE5FapKLTkrYT+buCanDd5BqRr8xP2Us9
587M3H4IfaAzCFY/p1Weo2rqx6kpUA6VDrcabchRAL5q4zBJ59YHF0LlZbLH37Nh
Pk71X+i/+YBmeef/OrpY01u2TAOGje91gp2SthphTL46fmnZJiqqfahlcJopU57o
LgEpH0jY7d56dMxU94HG/1EdQ+sLswijP6dljf5LwoQeuQQJAZcsChabK9wEtuhy
vRCt+XlhdbMYcrkLauhp0FOtPTxQ81HAjZseQowQ/nZsCof4w8qTryEymMB9THVw
puKHCg8fGxVsGJqs7COrjl6PR/8R65plKAYdPRIgBUsj20UliI6PGFEetVnHdYSa
OiqgQVZFPHC1G3+LpELwSd38yKys+J4hd9hPioZp+h8I0DQZI0NyxLDpRuswS7Cs
PVAmhRk9ONIV0II9K3K0ePxVoT3EoHiJkclIbxqcRDHhLjPwip6IPi3aSdkkBF7T
oUPT2GIhL2iwVH9XQKkb9w6AABp/SP61UtytReGlKoAvm9Yqpg4v89K3OWxyqTvf
MpRc7iS+nXReCkBahQwcU5FHqTxB0mwxf+MJuQEiN3y8CLjCiIZN2Wk6ePW9hXdA
qx5XvslNJbE3Xf9IneoN1BpWWO/1t4R63ejxeAwK/JFQuWm1heBDq70IvB1eVN9J
QKjpZWV5JnFWDbONWAa2gZPdNdAOoFq38AgtFeJ/gUSz/Zpbh7/QtXRb/PYEDR9w
X1FkttGfxCiVFw4btosAvEVjmIEcczqE00fLzNO1ZzICXx1AEzZVrWeLcmpMwNwq
HVljw8BsBw0cnbTukinJGAKNl5HS09qRlLYlC84uM1TFUz2NcWNSpn1MGPQAwPOo
4VepBwgewAYyAbRgeirHHqxVuPsJdOZ1R+G2BzzOfx8U/XKO6hlNhub5USuQP5tZ
aQ4g49h44vC0z0kEN4bOJFy1GTK/lWbtFbtHRdSbDs0BgE8ujqjQNuOBl8N90u3h
qTPVLWH1J97amNhHnfglsG7h/a4oWVRKAvsABSeWq0ArfLx9q1KXPLOpA3shv7+h
XCGJJPs+S3shq52m5zNm1F58H83fpIY0lkiSX2yFGfaIiU9NocZgNIMM2iRpX6yp
OPR+oExb2hFN4DRPLEKbp9jvsPSWHuBvKh9R7w4R36QcAT4WiZ6BuUdY/M2eAbTK
nyFPUxH+syEjLzWZFr80UOHqhCcsb5WAD5uAWndAUsOM7/Zjigo7jRs59nN3tUPP
S9wku/Ayx7OtKiPmqiyT7Ya5IVvJysTScEN6gqFR2mfaGQXXJqeD9K9U1Dd+R0iE
yXL960D3YljlAydU+32norS9+QV7/c4PV/7kTBJwsAt+CeuzhQZlh6hr+DSBCr/+
kMTOrPezoAVN94tE1DXrgxazfYtBBgbHU5fHTpebUNGatu4kMUjP0VDZ1k6sZfEv
hrVVUvQufZwBXhP1b9rlfUzhi4HbDQ9xRDOfuVR/13L+oFOWGdhBFl7vbJIslVkU
/xnPMM15JrDKye8B/A+J7kQhSjXEkOaJ9njH4lCmKnHQqbTM6yUL+Fss5Cot4anZ
GGER5ST2ZWTf/lrIMlWj4zoSYCR/0DmrlNf3EdiEID3vBznawyoz6CerAjDu6ytX
7JWjio/+XU253+oCLuvOgFyy61nIH9la+MIjCXpVJ1Dpqq0WO2OtLj+7wO7Sk66c
YuabxRyXd+4vtyMEaT65ayr2E36KMRIg6phVfx6wyn+7b7FiaJDk4RIjkv1pCWHp
aBRmXN47BPqauSouFZiTD7jNJaOqxe+CtKYk3GMhPqU2L/MaX7JGumVQgA9g0Rtx
INQs4mNgiApseEbYCB9ECd1USPJQ4Q6biXQMbb3RCZO0LN+VRmGzKPS2SJnYkdSh
9en20XmMCOcgbQHYDpGNkFrXVfUbe8W5xFImtlygB1KnAgxLbQJvvohLs65mCxpA
0ck+SrQ7qL+THc2l9HURpgheRoXLeOE/k9NDBUKV29uBJ2+m5n+y+fmOsroEkYFS
Ejc2rDZHqAvSXdpBxDL47jcGy4WPNJtwi9H8vGpjgUh2DZ8tPVeJhLaCDfDJG9Qx
0SDbA/iT5ywjI7ZQ8HdAi+BUlslcvYeKO6ZdSQWmi4qSQjw37xzd6JctkrkJkxO7
xsDt88lEk5+9JOz1YOW6tRt0f0FnP9tjciXXWK8vl+N6k66LBo9EljwFFJUhlDrv
kGMLBmiMB8grgOQH4OWE1GIXBa66LVeI0PDrRTDRMqeBkkcJXyf5Gk/v9Cd6o6He
Ft7O2VF/2BhCGQ9/lyCeOGJ2Zw6R3rF5HvGi+HUAmPZgndFdX9vk5as0ZImUAOaK
015PeHTzLIRAs2Rg8NQDq/QqYSsal9vWbvPRNUB2pWGcdzuWX6WEzqLJ9feHv5IF
5+9G+lL1cFM50ukTPqmTMONnVswkJgqckTfzwubwPc8IPD05G+rR2npLqNGkBUwp
sNgNY9j5GoW3gkMARLysXzKY4EZZuPDVsTXnVaAC3BrQC01QJRz1UwEC7nCsOVtc
NtfXXw66mz9UcwbM5HZu/mYT33a/4S72OlGITbJ724oUFOTJcXlM11JF1MNLpjyA
4IeU08+Wo1DoJnOX0v1/oT4nG+BFya0Dtg8AyvXwldYtTWMe0Ik78reeCRvnjLuN
yBwzZTmyODrg9c9FlqurAHzqLxKPt5PMTnOdE+Y7iaDPtee0ZI/y06jqeJJo9Ps8
w6VX+9M/OHruBg+FLLkIHa60Mh9933kHu+8X4I8CfBBsC4oK8g6/dgkCyOgUrT9R
eO5OkEzI9X4HX/eoRnM5tJP8KfPd0kBI70wSnJuNUsi67NbfN8OnufHz0hX6SbPE
+Hh64EHG1+ZYj1YZgIy+R/h+JAWH4KP+rbBVbuzPtyr/hS0LVncIx8X9uBAHcISq
+9UkevjO5+LepxTgiTy0sWJvHMKTkcjXSJtvcoZOoEihl3lMluwKnHrCQxpVDvDs
V6qzl+k/KCtdGyQ1xKBtw8FQtFfAcP1bWaYcMwIKJ5AcT/P8YjKx06vRTExmrCdl
6V0/v4TTgmYdTdYzsqiDX7q/SdEDCmc/B69Qptl5jWSwgkPo7JQo9LdMyp1V1tUu
GHE2kT6B0tp8BfhHhstM0bfozTHb8cac+2ty7ZCnsdc6l330cn5xvXNDBhEUVdxg
NYkHTGjZNDEoiM9RRJzjSxEnWsmDeMwipkkcyA8AWmgmJhoVNcEQnUmZVEnAKJT9
cHG9OeFsmh+BDqm95tY+h8SAiv5ZytqOorfrYZsx7Sjv+h+knVSGdhXVWEVxSVJN
M65sO66aZsVULcVP9Zth26j4Iy4j8KuN7CqjHL8o50hgTCqL65np2zp5aB0q1/OJ
L+tmN9emSgfWMCZWBaFppS5U6BHKRpp6nD4jnUdFczGgZm/s4FYpphUQDApEBY90
/jXsw3HyGVNagqiTyhBlpboGfRtoy4XlMAzuZUn084N2zOm+7sHdSfvHDMpUq6xu
Y/44kQUgpVticFzvhyHXHxKnGlIv5ELEaW7LmbA7XUfimRjq4sYM7OpV9tcSHv1W
QkO4NLjdThzjiqKLjMEtJvJZJQamhrb025IZnEhPCqHQnzLM832KDhhbDQ52DCXg
Zb9t2QVrWlFRYxF/hk7W/kSC77wysAYt9ZXq7TcJ7m8CBnClWfUJe6hXD+InrcI7
YloCDbMX9qVJXZ+zwxZCZJeG+VSdZvXy+HVOrCv/Vh93/eWbWlP8mK/t1Gahoa3R
SDpGNo6EICY2rQt9mWkpIeR/89ftC/WO+i5P8d2kFUkq7wYl6xZqOZU50QBVqI2L
sVEZmNMYxaxMtOdEOaDP07zgQRuK/XhPb4zlB1IwAGbH0r8ELZ0C8sbb3Scsr0Ni
R8E7JGWZQu4PC2EsdqHkabevPwwHx095/MngpIzqxBdRpxFou9ZJdu4CLA01l0xH
z4zCjc46iiJz7cXzF2nkAzt5CLyYjgdWU5yhbw5q1Jgqzt1uo7kEN7T7QSwOHXj0
5De6VffwnQyowu/HFoefX7XuPMNoVLeSNumZzWnS8Yxd6THzEOqH1kAxXzaNjSNU
6wA4NWd+1GJm1J/L9oP6l/Sckq2is0KoNIosTDf7pVk+dpCQh3Zy4I8d5E6iWtH9
lhLIcYJhj0O3Cl6hYHOSJ83cP3FdvBwjLRLmN/SQ+WMWStx3o1IYPjZJ+a6WWZWo
kkDFX9WOXMyOOYSTjmaAE4Kbn73JH+VWxH1lj7BvZzMDFbnMHKI8sJqgQaJURbFN
nOSIBCIWXg8/YW+OuSfRQlNYymVNRUEJ9oC49HdsD/lpoXzzyGGmdtU9jxCN+Asj
kIQ/WiGMMB9Rr/S6Wh1zFnefBOXwlPxNoHwwudjVGh704PV0MDBg8bbqulx3q0OS
k+QhXmF5QdtpizznLTjqp9s1l4woScm2PUMIZFe9GTtxw6c66HPrzU6ShUDkG62y
5nk0Nb97/NrkYLi25eQLUaadz7Mc2tTCDWLUJhNfedkS6BopOXB05vp18eALJedw
ubVdRGIeJImZFm6NY72sxb8DQZmIjEKKdmIepq63l5GYt/rEu18ASPjAGGV6/S2N
rxTxIcEzffe7emFA+xnEBAw2D6RVwIs5NjGA+MwmcDymilhXpNdgWDnZbI4Pnl1v
zqr41wSWAq087FtH+qARcLYPNiwyPpZE5mWMBQ1NvvP9sLaXDsMOJpTtZBZ6FEs9
do5i20uaRXoAOF3OwPIx6ypVhixujSyYF7eMtVM20sh/r+r7ts4FnfgQ5De4sTYh
zxZ4qeJMEFh+tRbs0qbwnwvvS65Y4J2qHBoMhUuzQxF7XVIipjRrIoKINQCkKInY
/fb0N4MA4hHnsOu52EbQqRjdpEb176jITNIGCIqXUq3eyZci3KcfgzC8nLqTBww7
7tLy5Cq+thUd4j9POT09suzXFqEvUoEeAJkuizfpc4tNyI+p1I+lAhsBIUAjshRV
NnXLaWhu/N4crA/H+1isG2T34f6JkAPO1GG8aT9//TsilZPgrmjGdQUIuJyN2LPD
niRA1W5Hxh/Zcrnz4S6MfKStkd4Xo5x/sP1f2WCOuyOS8OVcgQG3yyCId34UynUg
+AE7Y/elWZVCjgxXWL+WFJiGDH/l01Jmhc1jyg2gPS9pITOYx1jThPyi4G3lCX8U
ytYskc4BgFuTtGsVW3zYa0DPnhOloUL7uxi3TqdREQIcIodFKjqLgvhHDpYSuOEP
GAU0puXoooZrGcRuAXj/URwKSzEDUkCnVcOOVf0aYsnCZi556YnvbgWqsEgpPty2
CYPXrLxbJW8jVFvde27ZYBrm8aP3xml8zVw85HvqiOB3v9/n842kA+hIWqjLj5fE
PdPH0/sGbaYvycRpbmZdXMqDQAl55JKxbMKv7KT4nBo31EsB84v0IqHGInK9Dfp0
LCXI4yQ84ndWqzy0kvG4Rr7e9pjprLTskkNh4YVC6t6KXBPGsfq3P/Y5k2xTNrAb
HuDuSlcMPQh4xY+2In/n5ZZirz2oFW97cX+iLvs6VwEYAkCFdF/cMXHd4DcAeJw/
9bcI3+wVo3Yh7kyt5+KLAdjwDt4jRiafuc3isGqXQ4Hj3q1XXgOYPD0Bc1bdaOtH
xH70sbb1QeqJi40ynwhZnkQRCRs65aw51fUIOglgMEt7QNjLotbcn0yNLX4Xb9Rq
j4ELBs3IRXP6MiWMFlh8SmLvHMsSafEUP96LAEGNTVRITTpOFhala7iMNWAMeWp3
BfyCsL/DV92+9Bi2k64f0Z0mNiu/uUyWfm1/wIbB9JxdKixZkJRBzLzrvFv2J7yZ
bKT0n56N/qwqjkzALXVnC/CPq855iBQMSr5MUqaO1qAdBpY/dmvvyE7P5bODPSJY
gwTRQEo7QH7eDzZdSFa6pidCRGVY/jlO+htQCYzTRKZEOMEPB+immyG8evJicMpB
ue7MP/vvo7xHzQtJogCPkmSm3eJ9Hu2I86J7PyNbad1pOQxSecEWI8NrVJV1so3T
hKK1cihpVo912ZJxJz+fz9sBwJ4fBKZHuPK+yy0hMl1EiW8mMZGzzc0vatsaW2wj
50J9u6KLTB1RcxkgQNOvuqyIqSEhtyf9gtdS3IbfvOjpkUNa0NRYJKTHFhdmkHIZ
xID0imwmSrCg6zO1/rSXjKA9f87mX50PdlIgAboGXRtsTPaxccJsedyebyh25wqn
mTcBn8FGg2BBJyArMCKuUOpke4/ttAAXdR/Xf/7f45eO1P8jCEh3scMIPQ9rbMGA
iQDb5Bln9WzEPUyZZvzZDQtYzWL/bkykcrNo0meyQ5IVdqL0F33C1BVmZdP44NGM
zn3gsfXshf+d+ahPJDc6O5Q/RKcUNk83TZB7YPWSpoIIZJD4AtClRp6/JVWBv9WF
UinWAYGagAQ9410QPfNT0A8KEIiVEXtP1qiQeGpUyVqv7OGnob0X4cAoMZS0Rabx
uRhP4ihnovdusXcwE/bNHEgYbXvUvtiQIDmFHXQgJZbRU7tpoqu3te2r2IYyMBeG
kO4Mvtg9HU/3pAu+HBXI17qp2yfmWKmm/64kfbbT6gPqfQ8ZVZ5LumTEX41cQ6Mx
aAEpE2tW9K91Qv6zNHK5+f281sXgs7TQFAN53SKZTWBbGRIjQp7TP3GVEyHMnLYR
LDm++7owLhuF3/uPnhoAetaT0U4M05NlNwo4Frnsrq156kQdVW9p+A0wbH0g4H9t
f4RcyQDNketosdUvo4BZHxkR0F2mX+L7F6ncPumEFqnhYhIGFhoZzgB5pEmFA6Gl
l2HFyQDVuGgDWzce52toss7rbFekQS1+NavfdhGVwxG4FnX1B3Ep0X3iQuIwohkI
wqLhZCQjmzl13Ve3kLVehFNUrMgQHEqqPDOVXsDKdQ9pJOdi9grcltT0tK6kPUWF
8tAXrRWlRpwKRyypTVEGLn+qe/H8CodOnwF3mTEsz1/NTdkeF6OHN1X/gf2Sahve
6IWvvtek4+GbHCdyVaEz3tQxZiBzcpVPdWpbHCDNvAFDyrClhafw1bdaocLXYH4F
7E0Py7vTaj/jP3gCp7wk+bjVuVn+VsBxmyK3haKovsEqQqpbBeM6EiQujmRQDYis
MF0+uk/CP80R9LRpLbuBxqqv98IwR5QZRTjHKGWMf0OE9pe/tU6sK0/j8qefgVkq
L/uhYYJU3ZMAHmGGKbUyaEfeHA+uPc0FbIWGn/ytQI75PWVqrCXJwepDBY2JAjYo
HcJdn15IpLjAcQGBZpb+yP8Cjg5GkNcGYBeqYmY/wnLYvCVoY5M2C7DGTMG83tBj
k5NYY1oVuh01sLuRJGSYWzCgQmaq7DiEFR+3khMXcraLvbbHrM5KoNXVcX9f4863
kRIKD5StHWMZf2R9TXgHTO8INRNBMjhKRJRK7X+d8XC5F7q0wxLLrEm8EQmCMTJp
+ywrOX/EAn4zWSFeR3PDjmXdG9UuuxOHgZMASdGQnJhhqk660BYPWgdRlhh1EJ6w
WDGYUtOp8pv/jU05ij3SxooRyJSUuunyQ02ECDjUqyqyd3jKY6lx9vcbwEgnEbZP
PJGYXCTDaKi04XpXysfl4P6lud+gbCI7ytZkHOKKems8zYCzTl6v9+zHgiHo4zAL
p7ALXCrDM4NNdwmjoz0JDX4prxBOlpi47ARIhJ1M4sHr+6o/lYHGuS5PF9QHpX8f
7c2ye8EUn74IgKyNs4DHvvsEvxjl8g50jUN49JUmKtG7Jr5O6aYeENR5+8HYUKGW
kxYMW4L2esEigLHwKM9QT+nZE7g6lMbsMoWoNs/56UT7QWUfToKLOQAwfk86iOrB
wJd7dWeMGSfD+Q2BsolzZ0JVhjbjMTpfwPfrZRfbxUWog1Sk20skQzk1UztHogic
wQWedIm1b3H3SPjSJGupNKsOORlC244Gn67NoccFc2tCe5YISdlYdYCAstSjI3cL
rS/n/C24J5XPGW57LHTeuDJa8kkrSJNDjI8jZpO4j7bldZbjPHrQ9ZH35AQnhTQN
sTlwTxzOQLHok13bgo+cif5Dgh80OSQ68AF1SBEMRjJAb3iqJzHdp/fKEsODwq01
9H0keiWkw5av0sFyvz2UGbHaEtD24fiFXEs/qO48ud9gkhamtY+cGa+4AaCjzq/G
ObA731n2Ub+61yEmLPA2/oH5+XcbBdEl1eyNmwj+Gb6vAZdf1yFCNjNLbrPAkClP
ZycnYt3sIFM9It9lD+S1z48oA97oj00QzVlkU1Ymg4pHDZgeduR69BfDZHZci1SS
6d1ZjNMi9+WP7r3n06UGlZIwvlDt+J+F1lKtbpki9N7JOC8icvAN7H+vp6XYA3Ia
UMJyNvGk1nTaudqNcc89A+7mUP8jziSuDQvBm9CC454rFzMxwWQN9xSSV4Jwpe8t
Vokwr6YbCT+OBHIqDN7CgI/3iHBSD6npEjrMQkzh8VoBODG7CmQGTylh1EO6qEqB
gTvBfBp1NNy81t6MfbVA/LYRFPO9JfGhXxk3yWgtaQ5cOa9/HCobTzgtNCDV9t0x
BRkyro47vUXcNaI5XTIavGCRLc4AATmfn/Ml2i8TcmyoNhdBH2AFPRYrGOY8osGY
qVlODGsdCnEFxnGKmxUg1KXUKtVMdyG3zLrQPEMwdtZ2bkfWRphDykvnKek2uCtk
Ogp3isYXZZbHMpkHEN50bkNsWuR/v8uOFTnAYrv9p7bTLIK86Am7Z5wtxxE6nc/f
ZBE67LutHjJfQrq7lcYMjDAeCjuXURriP67qf49xihXsko/X5TY9GL/+U4+NGEjo
q6Y2guog4gsMUi8GFk1NvGR4lTCAlcyRL1TusPhNm8IO/qiR8c5gU//lAcN+JqhK
3+2xg66vpx0moqLh4TPgbGbjw7e3sE4uOOggV3dPrLhAo7H+wMCv+ktaP6xRIbrO
14rbcIHlvbrcsluGPRTd12Rfv7igCj1+VXBsCmCQi1FCCt0eG2626Z5LQwWCxgfr
G2eImzg6bOIxDYsItHJCyAlApFC75zD+Q/WrBALNmDLXU5w5Jtfi4ogHpCIdrRTC
UTNKdX7I7T8r92wyofI7tFL18qG4ew6xygHIiBqhDgWco2EpPeDDZobLXzqw9j77
fpSP2GYNGEgObNJThnGTjVpwDooi+EOAzY/sQO26J9LOwJYKTuIxZwodPc0uBSc0
jKaivaIjh3kCchAT4HuH0dpJMHK+GQCWANofPRCMSHXC3GxMNC5q79FmvcRjKlMQ
9OFlJ7zzMIFUR9yBsqoQxeu+cBlXZW5KTdhL3wec51jcxwJFfKIpNbMASoHli8Gf
w9zQMWlBN8sQnDa+dl3S9o6AB7MG0XI870aCq0a8i0YPCDjCbPlVP3d26C3uGDNp
r7QjyCX34+POG8+eFBr7iqrHA0vaJi0sWzLe6as99T8jiQSxHUhOEMVkCI3gKscC
M9+pZk4UmmPWMnJyWx0GulW1zukobFj6gZyWuI9ifid/me1r8LFmdGA84s8kzNkO
xa5KU5IQzY0tMPEsaOrzRSEKUfI8rXDDaBZdFHbA2mHme0juofTpczNbYQgqxYVK
3U3r0QGWklxmFPi5wIMYZTL4RXZPFhjsBaYSg2KAhYmFwUYMDYhujGwoWnXdM5+x
eXvnQvhLLwO12NUhwfMETcEF09evY1lr+yjxrE7SQDKbgqA7QTChWOmkKvvwM7GD
u7tXVadEsP24OZoMrQpNA4LQY7uBh6tZiRZFaHcU16mSm2RbpjBpo2ENaGdn6MT4
bvBLAaH35/YVYr+I8nXuPEIt6eFQoXKhMTNwod56zaJpYetcusmfJt7dl95dyOi2
kYwh2QUvvqDnmH/QlEsIvLZYGFkdLzSK20CHL/lefidiyNQFFr7uezenTyV/Y/D7
peVjcf1Z+lyoFM/WDL6waatUPrQk+AjjkyKF28nBQZu7iOV7IeVc9Qn6WLfWTuAw
T0HXX02uztbYFT/B6+FRO7e0ZHgwijddc00lfLoDhVqE/bulIpUPoYicQD3uYDg/
aLZGZ9ohlpzos6j9nEteF6denun3qjnPq9JYD6MzKHRSURCFSxFa2czawgVuqJW7
HY1LsNvurPIQvjNkVcT48BNLj0tJr0vnOUzKFD5W7ADTEaZwv3RTOCseP5Fd1N0a
+XZ5QN6YH0vDlbCHyrj5StCLr6vGH6QJWsVlh47lzXjQd2P1UkFPpLMRrIkQOzoP
V97L/P4oqEDtuqlDU+T7IKQxgblSG5iRhdt+YlS6m35wV1dljzuDnuLOGCYJSIJF
tr2Btq3bgAw+B/9kxfYoQRsus95+X3VoOOFJQcdkd78i1AdwsPgVigWDcJ/qXj9g
PKTRyeT3LxcJiXJNlvdCjQj7xWVVnIOEJMizoYMgHicanW+ErHkIYIGLCjJsYO2d
Rdj+HoA9XrhpAbH2WiP4uu6kXNEeUrXuZwXQOwViEA0qogH0NkMmTb/lqRyFLGSW
kz1LYFJwHn6vbXNEXUmagYbEpjgeQ0DGDZk5aJu8zuJrUA/uqpELemJQ90hhzHBF
GcXNfGAQmG19eM/Bu8Zo7rh9XLR3TB1gazi2P9mByLsu0TfIMuK6EcPOZ8teqx5K
emdup965jTCltROAP6+O2zc/NBwlNmnbDnPO4pa25AEl9+ta0bRP3LtzAoE0jDz6
iMJHZHrkuSa6djfQv4GQw+8QSXiAcAj2mADJ2lzo0TKhrt95a9/lcDRoDa3Z8yxy
OmAASxc0gMeKq7yrIyjFtwPIuR4CqEkVhPBkVpaHukdyfgrE+Z+UH/mZ8/x30UGa
h7RbdqSOI9eyUz4b9Z81MMPDuYm58sEjue8hg19jzzMvgm8UOK7c3ayx44uN//fB
n/ghP2wDiRNGPJe/00PXDjnUZ0us2ruQf4D+tPw9UdAbNBAAvCjlGF+yNbwrCBBu
niJ4yeJ8Ku+gZRTfxDQsdut3BlfNixyAo12X/JSeTSY6fRPhvgnrgMrSPgjaAqvB
eJEHPN7nvYAXMzS1FSkE8VdZWBxRWrVTDKpzwxo+5GqwrHCULXD0ZsPRZ5nD9DkB
VZ6fy4ukxNHgW16tFxCpjfEMztF4ZPy4PgLYRE5i2pkAiVCHpo+qSs2mApch5y/L
4iukCWfMCTfLR2svxmN1NQS8/5eZPqlj2ZAX1EIbiI+FWSvjZoRe4tqtt5IJHmgb
YSUIubG97wMUI1JyE6aMvG1hGgSoWYCYKj/9HpN07y3YgIvB7zib7vLXB4ELZWp+
i2B0apdayw+iIeL6oTxtplfUIBbYDEqOPfkDux5AymJErOUBsRffF0t/yXOs4459
8ZEX3AlTqmK99vE7Qgrbfxomsw8GSRAksiIoZlW8n7vFy2CowjX/tIkzVLRI1sXy
tQf7Iiik6gJkOYxpQsIJbg3r4RmSc9egMH0QcXtfXy6ry201VDUMA6+C5OSmGseB
lElkreH8cJmWII9YAyyXclc82pA+L+A+baEk32gvlZJsm31RR3dHOeGQdiWIhHaB
5Uu1j7Yd7xX3qPDB8VPvl4ecwoFPmm+v/uf5RLhvkhUmxzjt/zFF77PIqfbwpW7J
tvA1BuExLn3pTQNsWCRJehkdHlfwAvxjgunNGJlG8LlM6wCfOT+Xba60IRAatEqm
hYSmHzVCNTKuo3vKW+vD6+7iUHlN2Ixuar9ceqF4Jc/wKFQWmORI6ubXXnZ1mWuj
EmH8o4Y+sE+4pa5gp7bLOW8AgMkfZO1pCAfCxljZxUsYJVxp5UeDIUND0GC9SsFF
IEVUehQnDiIs514c4ozqn7Du8Xnl2Ah5lZhXnydTxURr4pN+toU6oejdu6dE2o8C
qjEFUoVSnzr4CTtUlweqLjr82KhnhuM7fkiTUvm3pwSoxkp/GD7DR2ReHw2lcet/
xO1DOV9toFxXE008czMZNwfZYtQSCYx86AXfOIA7PmoObVI0zxuwIuPg+pvJ+hDR
PlJDvGRUem1QgpXQUZrdmdANLxg945isyTIjb/YlR7C+2V5qah419oW6Nrv/DcVA
9Wds679fISBUNETBU1J59Pe09EbTcT0/OiO01LaVj4AeZ9Ft28tQqQIdvJdzhFmM
e9YtAHhUid8l1kSzVF4N6k1453RjWm2XjpeuS/RsSOrPZF+quZOACAuwRR4qR/uD
khV4CTxT8n1l2+pJ4g4hbUAr2Ur+r6f6e+l1/B3GLG1hUXwFA4wuTOoihQCQpvnj
5MSBT5bmJ2/DakQC5LSY1XO6Axw2collC0sa1OmPg2DywHwMzyk5ZLmBfy8PZxDZ
kN4Jmp7tdj5t0ok62ogQKAzQNbyxdJp3sBONxBDqyf9t+aOYyJs1iRoOVdDdmDgw
rFaLJOjs1GTl9D5NrsCpbTmh6aebEbHPtKmRdOFAkVr8OgCsKzwDrrMLv/k28Ul9
iyvBaFb7XxWNMq1ShuwYWiEv8ysqtoGNPCywc3TayCHmryQwSq9WjRH2GB4ZObfQ
AlB6apfz9PN8dTGSjDFSAabH0OeW2/JGDjjR6InADRmPvi5zn4ey7EjHgFsyxpgo
HR/uXLkHllNdT0CviP/g9AwgR6Zd906O2Bk47cee5GCobcZi9cVCPAzs5+8VDu8R
H2Alzvcu3jDpgrhyvp+CnKwX7ynmhtTsj22IMnr+Um253RTHLi7TmXet+qafA7kh
Jhql7ZBg9iFrj4aCk1bjWwcYkxsQZcrZXtu5VpCUooY+1jegI1Pl8KhMFB+/1dOj
uAjY0ez1yaeTFS1BCfhg/woqRnZRF7z9+TZbe8AlELXm4YS7gI9gZ5iAZed59SVu
l+F4+lELTahZjURL+m3Gq61aOd8kJUKwHy7NyWkpVLeePKc+p7cdoQ6UGjd+yfug
rmlItFMo+45uefZD+QIZjVb0ElCC4r4uJ0YLPhHgz9vEPb0XZbUDBlEoHJib9+bj
dNFMvPJCm+CdflP9CYGokJlNhQeoatQslx6BTXLVPlWT4gb83vlhYHUL5xpAPq8W
ha2y11WyfoUR1+cEVZDSJvlcJ4ykAOXJprg6V4atYg7LB0wD4uGB4lbfXL/aTeY6
JW3J5L1+TtDeesM3DzD9ZXInobxYfyfC+z65QW0Wab/jymeeWnyuJydW2cRJ/gfP
xCj/GpCW1Eg3jMUXrb39ncmTveL8KH45Xip7KwTTa25a8t+/Jy6MDI1KgYKlAPxi
w/Z9lqxPBm36J5jKtn9JpGBeAazhwueBQHo1dnaJriH+O46KpiUQsNTkkZiJPGw6
npPDPae6dsRrF2AKutYHMyX0/LfjpWz8xkiU7XL+Zehf7b2GQSnNkCB+bELn1FAf
hDJ5YNdQJoHsZOy4T1/AAE1ZgJJNIDLmvXFqGd+3VRSrDC7ao9pkgs8uIhVCj2XY
2dyS9Kb7wlVt8Drx9gU5M7mVhOS96wr3t8WDdEmV9PfMKDfYnndQddmRtLdPvWcF
84cjQqNnYIMTwcy4/tK9QwwDDv4GRsWFOkFsmMvLttPzC1D9zA4DeWeTEljmzHqT
oHjpPxzwM4gMZvib/+iJWbYmRcZDiQlw9NDmanPxLkpIhZXQq3sbrep9FD8ynjto
p9JjFGO66DSy05ISwOG8ZP9Y1yRD4vt837L8aQlL+KzxJqXzRYCRYnnjatjAzrhg
J7R5TaSdQ/BP01x/w0VMo5Bv3DWvftarcGysM5N3oZ8JsZdyD1NPi+ZiAYfb1tL+
C6qz/CBzcAhc12YkMlbAweTAkMfwrL7ryamhiW09yVyudt7hrouv0JPhruKU5btD
TTzZWmjLfGqUDpVhDSq891cetzZVkat0UkbzmvLfG16/lc00zG5angXafbVo1heD
HtrIWu9+H+/Mv/kKz3oV5sSdzgwhLTTZtkPcrbITMXYbzPy5zMeYczgPEZK+2fo/
Xm4EpqF0JytHhbyT1/uTkDyJYR388/xwZ/cmQcXg/Yg5dpNiEFodKhLrwHFsXGgN
aXP/6Vgbkq6riT7GVex7x95kwClTwaBNAHgoMIWe5Xu0whg6rWUacL90NQrzRZq+
+jq1tpduyXaqFojJIEPZ53C/eOGWYCxMv7IicuKiv6xTu50LjDaTe50H31Hpp0dJ
AAEdRkwdjtCnB2iWGpB8uxnWpjhTKfNUya3Mlbg1H2ugIhReQJb/ALtto2uKfSRh
BbRAsuHxFZ7qDnKtBdF6pFjLrvS5cOkKOMqq9+YEG6/hvQXv9fa124x0JOXs8fkB
EltMqWeaqoW0VYU5YhCXgjmgc1Gv1EiVs0CjULFgDC5C16X0cnEGRI27QgFx1k3b
BFsRyQ6NWGQKvjhfpVgiQPvVWmwrVJENgyMkHMtuPvLiFN7Ao5D4Tsfpmp7VLPNP
LEO2vlUD18a68Cbx1dVSwP6gndkBPCJmTb1wIhLdLKWfGC9VdaqenQ9bGdmapVB/
G1C+avQOog7IfEuUBDF6eCQUmOxL0DGnghi1XpYF6yDj5d97zAhGzWVuxbmlUwU0
AlKTiIIDwsvrAP+Il+KATFVdWLE3f+ZABB5GmNbwJJ1/oFIzbLqaaG1tVxHq4+hj
t/1hlMTryzhWEPH/yZtrzPylfWDL6yd+7O20T8csNsqO+g+bNfQ1dBSmNK81eQjq
nGWQWJoybH1tV3Qjgenp/cJIll0SUFz8RKxTxTX+MXCQL3pbHFgO8/8axn1y+Wn4
F7fiMu5Lq3rfdKxIj/GUSVNM370T35mrCHHjKO/ASR5eEoQPrU+vq49mJ/q+FPOQ
J3oOG5thyt0SDfK0a9qXNJWD/t+GMcuhdymXC3angz21wSKdv0sEXh8rFE56L4g7
hgF7qcpAuw+DCYSsjHJxADNczWSh3rKeiFOcFCBLGugCPV3QkkBgw1FTW1Mie8+5
52RVnGx+9hufvTFC26uqF4gV3NNpr/ygALsbPqNAKQo2bCcUgeLLaLKs0LIAzvzf
CEe8twgW2sROKko5EShDQ8A3MxbMDXfJVcAvaOPNX6W2iKODv7v5qIKk+Jb4TPFp
0ld9WR4j47Diyi48xYmzQfzfBHAQAQiUh5E5SVX90jmxmBkOk4adwO6JEHNA2qDQ
MccbMR3N+PgWI1r1AREzwEQ15mGLJlGX2YnD3je3byfq33GVe83HMD2jJpJFlhEh
pHrFRSX+Y0IBOie432Yv91mrvbhfjY7MHnGgcwWHJI3a5Fv74BxeyuPOiFbakYua
ugjLIcX/dW6j01djnr5uTQfYsXTz6KL1FW1djZZAj1lQyO/ID1lzktRs+b/NVuG9
sjgjp69dTh3xycNOkkZQY+9UY/89dyKEHXM6rMHl8jTAcOMf+WIK254A6ilS211r
Xop3DZshC4xA0/UmI3KTPBis2rsrVZMdIqq0F9QagGQKtDtfPq2OWH9v97yQB331
3GUUItxSXzD5CkPfu9aZhklGButqhBlT1odUXK29dKUrjubeuuh5yrScBvfTs61i
sOQ20unkhlq6RrjXeWqKRgqunVlg+JeKGTaHDbmvdngHf7oOfXzhZJzzQEv2QlSr
YWbecFjXnzxBQ4EmF19hpy+ALn5MO/rpvTo7sUmfIG7puWqBucXjhCVeofYvbcJN
L/Y31/yfDaH6HCHTjwOeEzsbVr2DBD9sg5CFhiyKpzJGhliyFV7trIEkd9b38C+u
QDIEk9rNXoX2+GxS33RAQtkTPAz97++E39CGaISWV0OPGy/MVqLa3+t2qdBuhlTI
GcdTKdkf3sKtLCjnuMpQb/YrSm/AlBxpNJCPHil8bPFY7HmNrU7EWr3p63dvDUH0
b5VGeH+5+LgmyGiCMrKIUVpatC1EPb3zzt+DKwSlS9MS1mdTlWYE5pvg25x52j5M
ZRfzeU8+kQbOoLhaJIWZ3/6leETo48NXaEY47cICvFFyAu1LLdvQ+zwVxGtygIfJ
I60nOMDvP3ymmUSQHIzvJSPGtJtlJVfAT3/4OZbgZGjJ8H04AnH8KUR9NhhnQQE6
EcsahUkUp3P+3mFHtth59M4Dhi0ulLBRgCpwKeYu5X4vgdbDtFFX4+pPYx8zDa1L
TtIGOsoY0y9jWOBdS236A6QBmIN+wgGAINV1jFKfATF66IvwQvJcVjgwDxZ7jLre
sfE5wFdC5Wwh1/p6x4F7Az8/s72fU9W09ZfQxXUkVKI5tLMLhgBV8OFPye2ptylf
71Q0iY/3t0LLJx1i5xzOVeVPqkQDK2obCQo46U8xBzdVEkJC3n1TXlrPu6nBbq2W
H972I6MgYtMe8hDOUWFCW354fSqfCb83GPf60+iz91yGl8ep+5EKEwWY0zb7r0kp
WDLSiFKLdbtdRn0YBfmuR3XOBKx418FngE/nH2Umr3b9m7zqgxsrXUn6+mMFVNHf
lQ9QSgCNcSVeFErRwv2t6Zn3ugQuRaobwKcl0m/PA93/NmO1Q7rBWHxWl75A81/A
nNHyT/xKJ/nCeGp0LlxTGPkIsTmnwQwYbCFATJxTJ2ye/+42S94y3sOvCmdzsjjh
/DUR7+o4nClk87I4jtta80m2mgpMZWCparW1uq7M8VQaKIGBfQO//f+/U3sEUXa4
Bx1XK2bCw63oDO8dstK0whuFlLvfVzgQnNM0RAY5TPAYbZj6B+rfZTwgNcrByWz1
jMVzL0PaLWc+V9osAvuyhbqBYH51SoDi6s8wpxb2M0GDRMEQdJpng3YqDcmcDlap
bBn5g5Q8ZkH/RsNpovkGAdMclGmWfU2ELuuHCKrUm7Gn4MX/oAcgk/ZePzKrfG+o
c/yw9aBN+mHk4KMyckDIs2xk7rFnez16ZMaQhDWlsYgj1eJGsADOTKes8dxT7508
SWJxFgB43sVoT9SLWUyB+J2Zt48fZP7hmgxN8qYn2r1jJm3RCifQUM1/dF1WBI1K
nnpEeqX0n/gHXvm81m5IhqiN0fcANzwZKRrdskwo28qlBlEQjSkOayxLzJ0qmaM8
DFuD44b2LfOr64btRXIeg2mRhKr6/fnswCg3MteQL/Tpa9bE/yXxaSDEvssGGyx6
VGOAjE1a/bf08AEAnd905unSg+4OOpisIJaiHG68xnZfKN68xuFv2rGQM5U5N22w
FaUQjqPhYCeMRSzxqQ7Pc8exC3lDUZN948EMnOXLaiqqGnTnJf1tTqwWmAz3FTn+
LAj5KAZg40H1hNtAqI54E+Tt2BuQoEBACN+yFsEqn1ILtYADG98coYSPma5AaXEq
c3bFlCZSCMxngniZTAK6gTj/kSoHd1Gjrff7C87d4Ktw4QFW8PTPoe6Q5vClK04z
kKIRIGsAsJ0bokcEP4Iab+AVHnpRWLKNogUiOlZDJWbWdD7DJA3hvWJtXKe5gWhs
xeaLl+5rpgNMiLX2rZt6Rns44uDJbHsrKZTxy2+uSlE7Xwh8eFYRVUjI02zBEy4W
FiHTkV+PZUIBPUDq02jgzROrV9v8/nBLPEqyoLV5UyscZDX3b+JFebjQLdC0i0J0
hvVr1swkKh6bC/EZAfeVHNhop0uVJSfn8Fw/0zFMU67ln6Z/Vcb4kdMJ/aaOU7LI
r3MDpYymejciX/9RNinftvfnIhVEAjEdb79In3/FHm6+RLVB9xxVf38KvPG18pG8
uU2jX9sMLyLfu/S+Rx12WJW7YTIz7slTxpstFpHQQg6XBTT7tEtMEQO6rJ5FKWBH
59iGb0YiVg9VV3fAsdm63PxSNvRIMp5Dk0UIQGVKcIHhqy970WzFMDL33xlj6w0X
c2uv8T3JWBchmZR253eZ0gE73Knt0YH20GLmyris+45DGtFzbg96h443e8hX5U4x
Eif+AMMxlwsqVp68Jh8e8aHimL2ohYtLroBpBon74HKCXNleKAcyVetGAWmNeYIX
QNy+PZ4SCHHwVK6QIaTgoA3CWOuE5QK0xJpDetnoT+uFxONJlLkqOBJv9KX4EGJN
JA78DumpZ39w9Q53A+JjkhCoTuORnugJhrqPDIZrB1PFsqcWGRB70/TM3f9PIs9s
QjWznZO9bNpoEs4q9M/iqkaCg3Jb7Q/zW6E69s13a5OAZCAoA8NikVb9w7YMsFkI
Rhfc9+Eg6FGNlhH2lS7yCvaqskZJ8yK6JOULctErPWs0G4mNfl+FWFuX2fzHlMw/
VMFK1txMTsOu82H3iR9BMc/fUhZhoSNjRi5Gyv5VU2kM9fW4hMdFEgrpTcVcTXR7
snufXtRnpwbOqOLo7oEdTvJdw0HMYfY1UlBbk3IHi2VDTMcQpUabUNPXzWh8xXcw
Ci9wwqWaXSC5hRx8CCifY5nmRVIs5mIvHSd1W5HwPfhRqrQLsaBX+5zBMc+/eqm+
lFuJHNdVO7GxPUch9HpzRQMioLe/3ZQgrBQ/nIA+HGuwSlV/sHbXnYMy8k2Iw2c+
TmXKUo48a6LywcgNxYc0YONWIvCNITBbM1tTxqblGNw2npqW9lXHg0kWhtvxqX+a
aXx1XZARx2sTBfP4JuCcSzyQSxoXnilaqinUhRxhJRS1hkbuaccCNMLzjoB1EfTb
UgNdh+80UM5m0XOrGenEOX2tb/+i3qCEXu+/adTnXbbulw808PIyqm8aCrtjg4Iz
OJ4p+znuT/v1etUp8WBiXZp4eTzsZiKZGAdtNgH7vx7rCiZVuth+aTVuo5OplVP4
kdik67ufMO6SUWIBMhHnBUYsLMh/e3KmEu9tg2L442XkHi0h2uUOuPftEyjDDTJ6
EOMIeXrx2fS4c1vylRF3+6jb/a0PqqDvM0/U+WiQi2fe+srqgEU5Z52FBVr9YuEx
FlYzN7Rp1wVOhOH3qmkgOXXtpgsX7wC1jPrCTCvbd/5j+5+mzhj1PQKlhFQPUlEG
iNHDbjIWuKNnO+ItBisbJStaAeahRZq5nTwaor6PMI0YMvVbNqopOeR0UfQZz4Si
PB/VyMv3W7Ju1S4OOPxVwrpc5OCNj693RpTYsGB60mfHHLr6CswOnzs+u24MguGq
m7ipklhoKwMLgCrFCd80kWEod9qL92oaR8lWNWCZFrEhUE0ve4JReiFcNGCiNGHZ
BI0sTjC3RIWCHcEgRvPhRjbs1NbK5AbOohmobJnPtSL3zDVmEMKPFzzo388oM2BD
nnxWyIV70xzcqUAJyUyMCmhUCiFKa9E8fy27b56zYKrtstBwvfOPyyK5Py7TVMk0
VJ0boXGrs8qvjjfToW77GRsajqHbwtbfzStJNurpbns8/jU6pKpy7T11InMfvCch
Wf7FLBJWr3tkjC6UWA9NVUFYr1ZfKWP4S9k4P3V/UDmgjXTF6X49cS74W1CILixA
XH+9AAeIR6te3k3ALlEp9iHS6p9rAuPGZDrEu456Ckamy7wEhAY8S2dcoaWZY84A
qT14Dl3FveEaoc0but6QbgYVeu+OPY+HEx2sHpVSd4XXNB+hqo9O1opw3gMwJ268
KRA/fRNxsquZEc/jyP8LpFF1Ux1Ol82V+Rf8uduBTpJ9UTtNpCuY2x+pbPzduLNN
tY7rnumShJfE4sGl7h+zy9purHoGdrEkFbGzbLFCQeQmPQB2Hr8itK3ljTqsY/ts
fuzA+S9i1q2WbMb7+i9/jvCg27ss2DaDsFbX6WeXZRYjYLuZb55nOIc2Ghzv5ONq
rbKH1q7Utz4F0y2uHux1hfX8svjhisNyOUhMTXncn5pj4JrP09RWLBlj/yaExvZX
PhXF8/et4+2hCT1W/DLTODiwlteSC/gYry3dUUJA+xu9zxUqmTOD+48trYNev1SY
RkBVsx/eKOQ2HcnuBmnFDxhyMtEOqkp7JkIpx33ik0PG474lLR8IWptgzz91ATnN
kFqZGcBkWkBebcdf0eMmNDQsTmjLFmZCn7vVUU3BqTLAj5SkWSroW/fbIMuZ3LLK
4BBFfu6jgzNAy72h0JHLhdIVpLmyGui5/XFHYBmbeMJHIvimW1yXY/j3mOvb+a3l
9Mhe9Qiynf5aOrV0dsjUYEAmKCpns0mRCAzxXdeKuvqxagpOlEaD5+c6Gae/tJaL
+YJWty1hu3vq3fv6WdZ2t47Ht7QgTmqlI+3o/M7noKYYaX1V3gn0Y0/twBq972PT
DG/X7M8lro86zjPStXvTubaccA6OAaqDo1chkND6arEVAAdqM6KRbuuwhG8bbNfG
OiU6drfuZyzZHPILZGsy5uSMskAjl1bAAjbig2E8RelA0l1P9JUrfJMF4G3Zf0+c
ZWiwMIc4TsXYcI3tD8aTHhje5VQDhARDKAAPUl1arRb/v8PWY8vt+H0LGQ3WE3ga
GRC3d+zFnf8jZ5gXcHLKzqX2O9bsKEWpGT9DjQYK5k1SQAjGIxnO6iWv8GdbP1EQ
UFiAs8qMYtbl0bNha2aKSiiQrYrR0hPuq1mLJQIxxpW4PNI6olMcT18iXaICDg6P
Tr/PHzj+pXKHUA9sCiQbJHFEYZFSouPErad2t0OHfWX5f2TBMh/R7ybnRre9/Wkl
L0KnsFkh2U78KjyOt+2OoG0F87jcOmlycfzVUG9cXGFDkRUdBLz4AsGfCBDphS/D
BHgU8OdkDB/o0XJT9jALanaYUaD063Gt/e4ANXk9t1W1UGT2CQd/157gtdjTBk/y
cAUYeGdMlI4Q39u60eQGfeHzVplTBFi7G1r0OuiUo7C56pUDOx8UwF0Xs2BhCf7T
i+7xpxsA/dGVvlArJffU8+WRCYlSPZ7Me050yiAUwaPu4Btwl5wBFcDD/nJOCCId
1VwhSTTeVXTujnsBayxsOa6PVniSGAohE+UpN+6q3zSz8xlM+QZrs9uatxi/BjpU
li4aX6+eqRiuroiBawgsXk3nQmn+//D/myx57ID8UYmcSRttmP6AQgH5Wv3S8/vf
kQo05yV5LNZxkrJ0Ys+pcdW0uyepEiNVE19G2vJH41JofXqTxYBc5vyfsJst8Yu0
uIwUBT1SqmmcOdwtnXZeaobEH5YnlrrjsM9DH7LE5XXH7Z4G5LRq39QUHOxnCfOe
lQL7YgUD3f10fOrL9nNW1fYeCEQMieYV2FdRd4AyC6og55rBDpZv+gcuFU6z1pmU
8VZP0m96kp2p1SgnS1P1FR2d3+e2yEdHcjJPTOnnE8hR/v6sd4ZyFpQMzoYvIC4k
N5ceP+N/0iXKUo9gUPogeVwMfILeOuO/p41cY8bnTGf+OjxL4KaXF7RMzsIaBC6k
XD4nX0DQpWqNOENDmE7JY8miUeZ1pHJ6iYZJWV/Z+F18V37SybkUuVydQFgNGd6A
2CcML4kuWN+mrtlqWyMvw6Q9vUdCGNXqYLC9753knI/4ru4heEVN7mjHBtUn9DLx
PEFxYxQth/42SgftXnil7nZSv7aM3SPlvQN1vjS//wRRabWFLN58xNeYiDjYlUEa
eTi2FYr6i0ZXuYGenURBn1/kgb+2xhl+wEo9Awt3lHB3GnpcF0ELrXuJZaKBIeWG
GLrbYzl0tdyFBuwJECK3I00QDzWqt+cNvkZmtWEH0DPfpO1avpAvGtYuLC4NVsBb
7xw3D7UZOvrg6b8MDFTOYYkW9D3chrDzf4585fE9+AOFfVYd48B7HPF2kFi3psC3
WiFWmRb22Ulcyu5YY00hZZ+rt0a8FQ8T8lUEa4tcPoVYEk4IZfcrK9xnTUGV7sgp
BdcrF6DV0vu9iK4fe0joUihMlJIRRal/lCeEZdl/54sET9N24qDUh1fSa3kzPS7n
OstvhtuYohoy6QwJbbm23aLYTIKznBkJa53EXIMpLa+5HzFVRllIJdlRUEj+Kb8C
JqJro2kwunXN7B4aDpWiCERm1DVbW+aXTFddB4hkp5Ot5vtbFxukmwBzQbo4Vy+9
KpE8h9WSRXYeGECAhr9wqrHJXLoHgcSp64x90llRlFil6aFMuNkIT28IMS3mKvgE
8H83Gx7EsnHuK1a2gWi1f4/ZlJb8jL+dyJgrai+6w5rU1HPHFuaeN0GsvSKlDjAw
EZLrUppP0ETi68S26TioGdY5sUzGbgSzlauVdz3Oqw6IIGikLLhT3q7sv+krsmKo
x7kGYTePMffbmJ09AGps+2ad60m7xIKTFJul/BQ2X0iXOepXZUkNEORSGymbb2HS
64rK62m9kFawdIPN0zTfwj0Gj/iOu6OyTyt7pJYLV/0Cto6+DQlnKZK7WF0TssoB
PwHkQcDXjLKcjG7FFwrorvW9GqfnGmeDBn4cCaEFOpqpTcbe/KSIql1QC+CmoeHZ
6Dobu9wyaZUMDeoftgOpAWFDSALx6Qv+w8HiEC96OnY/eEknITalj56ey+/Are0p
NCfPIW279pphmvHwUIHMoWu3I0tqJJKajMpa1y8yF6rJQAeZJQnFIC3lThtoSJ7c
JaCnaU+5aDlRzwvl42lL3061ZDilnvihJsPNjKg3PCs6nfXvRKlX5SCzX6T9zYjf
air1n5tKPjsdkW4x6Akg8F/jDRJGD4hVoT3q+YeBwNxvO+OoCh6BacAb/7NSJnUS
mm4FlHQvCM+nMSZhZg7FxcowN6qWdBNu0+giBplohYBLDFPw6+c/OTFoK8WYQbqZ
JTTsla3iIIsOdCOM+TfaAGS2bVytRGIspwTC2iaJTp2WInAMALUADrWcUia1Xrfn
kO9J01K6UP0aeoauJ5YDF6cs7BOtF0ZqKpv1nx8CRqluIcnOSNgMjJYRBWEy66bN
lNjJlBIh9vaU3dfsP7GTmU3xBAgua5Eo5qDIfo0ij2CI3iib3KsaG6bo9RXElegM
CXuPJd7z7ugsgxFixpwn18yfelr45QT3yInSc+2GFGgKlvuxVXcZAu4Nd8QSsDBX
IgMWLovx1L3456emYKigVTH8rj05+lTno1m5jtHsSpggs7vQb1fQZ8PEqmG7O+Hv
lHjZV+N3/yFX9p9FCRX5+IUu6owlNRrPtVP6By6YTmZz7+yKmKurHYFOgMJxTRuS
sOcdnbEJMqbme8SRJhkF1D5lgKpYpIvHCxW5LKYGxNOL3wTBIJNUKfDQxyyg01Vy
2TgzmUwfL3i1/WJ0Q+I3iR9CrITx/sGEMSGP3CEhnS74PBXTleohx2iUtdGE6xcY
q7UXOE6fR205bBjulqTnvGFpJYoWMl2Uc5uA/EkChFOLl3zfktl/Ese3Y7ePecuQ
Jl8tymjUUKF48yWrth4c41Da7FM7u996AcfKSIGC0DVqDPq0a7N9sMCYW+vPyR7/
GRNz6XbQEqXajvmEwYgNC0rsplvKntq7w8vVR3vsYwgSqQS786tAtuAF/iQbWQLz
HQ3Yl1ntOae+bzcNHPy7pL/gF2Iru9QbsB8ueE3QKIF+XJOxmd+Iqs5MNvtqG2Im
g21Q85xh3MPidL+kjmDTKiZVzQjsnQ6kTti1cQ1XzPPuAP19O3z1iRkfylR1P79L
pzrSXzjou/BryVihwD8p4V+KULOMiLsMl4YrwQ+xKwrh8Q6qS7w/zmTIkL2CR+nP
rhylbQHKBjuXXnmq0hAP37Xj4jWVD/zHCmFNlq49J9TOT0fviO0io7D4JlQaJkNs
3TBPvvYFknM5Qfn9Lxi+ut57B0zHStHIZUCo1NUpLIAVm0J88zq6TsdNRCBSHsPk
RhO8hroorWnQ42HRjidi36tbWghhI7agKLpn2gDlFvwOM1Ak0NnvXFMa+HIvvvfL
cS4ChL9eBViVLpt8rZdAvHN1Ce27Sy/mBqDyvx5CVNawqQxl/M5pm6xdJbYxGEb4
QAw4kac6FhO76OTynuom9V54B/AbS3YRuOzeQ/JpUZsxGTavEp+Ji8+ZLdtKHrWw
9zjFRfuv/ql97YGmjvIq+mus86fRlK10q9bEiuotdUE3hEH9TCD+gPlzZsA8fkLl
SE0ZeF9pzPplz6SPoaKiqhJpR6HRkT1PYUeWnUdY9veRH7p371pkKv1/b/VLxqde
mYxF3CxVvYaIX47KBQJwJ3vxpBomzhrS4FqL+rsHn7NZQx6vpp4ckAxkgOXRDogf
SEVxAy8zYuK8ftZOh4CuKd4KcIf3FpeuTbbNOO0J/5jPdkE9ocZNlCKCnC+B3r0W
HCZMElGOhC/vaen9d5wmCdJqgPWPUF6DvFRdGM8ugAmrLCP1CdxVxKPmQLQdAGip
Oj8HPadGETEVCPbJnj1xhdVAOfsQyaWdf3An6f4eV3fdVhKYQzuNm2NKfKChBvh0
+3wJik77rDjE02xBrrky6Oybr3lZkndEuchXcZPrelVMPIdMAnX3G57jy7p0luTl
/8lDEJxvjXz7wdJ6mI4mFd+JFcDEcdRvtkdlddYGr0zU2pq3gzmE+CJ+0E3JvYOw
+nA75qkf00UWoV6QDUcTrhVSCbIU5+/hWYgZ2vf124rE5I4Q7uBYCZfRysxU+BKt
LPrwphgTP3aBGMZyTcdHeYGpK3J9Q4QFf+RoATp0uf4jv1q8x0J3euNnJcIW6UNS
1JGtDEuVpV+UI5uvVw1yWBliwJhA3M8tmp5X9D5bC/r/1laMrDseP4mbF5B3EyQP
3MpuXcUvwxOI4yLA1WNmSf6ozYSmKjTKjH7fm4XqRvj8EKSrfOrUAcO+2rvSWCd5
bEExi9kHuiFpdK4nz66wJJoNu/OtwF6kpxaOdRD9mcMOYxaHKKKk1bdIgv0Yb4yk
SwTKg6yb/ulLcqLAX2HKOK9iH/j0zmCjtW63i476Llupf56UkxbowitLbQ1vn9sS
CzAFekdJl1B4rGml3C2vOxFfcibEFeC7EWODb+PB63l2zCNuddNZ2r4JSmqJNHvq
ugl5OMj1CDsPt+ZGjvK9dd7BtQDaKLe1hmnvQHYzJq7TJLm8XVy1NZkdoagsmFb5
R92zSyz0dlLRWoBsDiFAYYTVGjfT12uUlvdJhnuQfVh45Ouy2p898W05Q5a8vkSR
0CGs8+0yWXryKulh+L25RLw7jdy2ID8J2+Br8iRk8BIaO4aZdI+dkEqJY4m6n5Oq
U1tD3CdaIHBEUvfUDIGI3Y4trZ97+txsRAafI0kASnvmP9O51q7WnmtTYedntjAu
Ublja85o+uHbSLB86PWzDWFHBYs61cSs9LlEk5ZPbSvZG7p+zsxFm6jizjOQi2IO
6ijCbuXgIYM1oqYbyW1X7ZhyE/pWtMmcNAvL+piWJQb0i9/DbdfK9Y+TEPCyBbRU
XnGkf3fQQGJ3SwHAjK8Cof9cTJC2FLvqnKakHo/kGBPYspRya5yASt/2ito5+Zii
lcTTLpF2w75sw5mAv1iw/cqP1VBiNKDbZIDxf8B7kGicx1VKK8ZKcBtrDJoNNJSb
+aOHqooerCH1UGZuzokGW/UPAU6iCvRUohoDqfGq5mw+i7n+fbhH3Doq01TKfM96
CtAIpUM4B3590HxSEq6osgTjH9G4ekb0XsJZcthd+suDrhpjlAQNGHd2yQMkxHEu
Eu3HSbV6ni7UAHTwPKEO3UGUhdUfIxZCQX+TOGzUYJnr8ld1GwWrZRDy/HlICJb9
2yedEx+kI9C0mFNqtbBWDDoKY9nbpD6bvC/JEDEVBnKgCARc/LOzSQqxC22/kVug
R6FmWCRyhKtsKsK31nFvnLqCiz33EJPRca/XX8zjYp3yMaoYxsYXkq18tojL/P9m
XaNgtd/kpPQ0nG8gPXdvwzPIz2xixiQ2LAqMBf3mEuzjyPZtX5VHZKDerNBgXZbL
sJNLFs5aO8o8j7Si8TAwJVQiWOZHGzzHBhM0JrpUKaOs6QIkI7KvZ8knrczDqYFf
x5Kh0QnHZIUvvACgHRijjkTa54sBE0yPi27lTJCpB9tOIvtbDPXlSV5GMs6UUr8Z
byX+vXdoskQzryE6+9cekDZuF4Xy52vhVZCykGtKxxATPfjaBNSi1gfS5edmHIgt
1ItKIZUrnRGqb8+pxYryloQePoGsvF5fwn/Glve69eq/Tgtcy/kRGdeSkvRm3I1A
CgBewT7XrW1GbBJCbQTFcGjM9FrFFHZ+L2c4QGtZCjI/I7x2/dMBq8jRaBQvdB98
VxoeHTTKuqpGXOPWw/gfky535AIYAe/geY/p6B8ibCgbmBO4FBp5PaZFnDl8lTcA
9Ev4kUHHS447Ymakh74yJbiHmnAkrBdXq68zjbdiPXn+tao57meqDUCD/pt3XHlc
qxtsg83F0h9XgWJ3Pk2aYupkwHi2vKkvY1F42F7cqZXQ+KEPGy0HO9rSfYokTP7/
rD1lHEXRXFzbNnDVp/T1DuXxuFwjoaj50y6+6pWOiL/wfsWEhpGWeoHEaz5YwVNE
VTcqmemy1t7K1gps/QDIQ+df4xgX9wyvsz4DWUpgxeekiaJRo+2C6r9/RJcgxyeE
iU4kXDaVRSHkFl8Mhn44GMEyIt3TkMoK4+sGhxKmTpPI8Ezne99hKfBDqWUyvzB/
rwO2yWAq3eJzN3vntvJu/YlTdg1XdNvbEEJb0J9HYG9AHlK2vsAXJaJccjnkfx14
yrrOijJwZvcaqw+uv6el49/medWSWfccTqWcAHU6LmEUm4RdNko+aqXiTLdnEj7/
HHZDpIrzsrQS2CLH5BJ7vgbCwgE2PssoJcAUA3plwm3mhlGa7K+4F6Y17Xdi6SO9
YcRSLZBm1+qemfk4tsqDQ4toh/KPM+DIHTGLwdSwFEodIM9uDZY1gl+j3xyC1ynl
jmV+uoeQC4EcLP6w+a2l6NX7nNZ5OEH2LY5r8PJq85EYYEjT10W5wNoQBN4xbbxx
gyixoWwdA7Onq9Tjuvj46Ek7qBJgr6a5I6x39httMbnAF43h3L0AeNH8EB7HkwNy
6b7VXrIG/Ni4YZm5eok9SWbPXqX/Q3X6zKQ8xtzHSDfw1wUIoXglHbDMowl4W03B
uUp/zk44fKe1uth3/zAKY4jOwTypimU23HAvq9u8EZMNDS9bH86wJvqpRL39NDxT
xTzElzrBnns96JEhYAPgdeuWoZqyIW4OXWjizJj/60mbY7KicRCNBkGOJDV/C59S
5zro0jhSWBntZSllXk+fXW1nUJQNgbi87OLXhvJ8wvDkJfS0a+Yfm4sdwQAetRMo
7E8dJCpcfkiN9xfU7DQne34y1nnvcdytDxfyM7YcQKEaokOwMCUJGYlyMXMVj3A4
+ISZFjRzqgwco0idUbeDdQFzqwN5+fTJnwQrtNNKZeXG1kosDXiJLcldADtLZvk+
xVxwULG0fQObSimbrcb30nctOr5MFaGsuKDWfbRK8m5X+6u4zbwpqa28lg02XSXH
edmU/ynD+GpTaeJmwW/deNlPKFvc7QfEEMlq58WNsrSJTmxnqW+eT023p/NfhYGN
3QTCvstUzq+CvyFUL6mvnSG4TlTkSMmHObfUQy09LuRN6Kcaak/afEA+3FIn4D+7
eFx8mEwcwH8duHhV85BRnSkAOab/9Qvmgo3LgDXJeHW939eWYgSE4H+l+ZwkzcPA
U6Bqtlyc8p9SsQw8oypvLRP3DVg7XqNNW3eV9gPrZpbqOZFU6htwxDWhr1q3deMY
3vCl+00342geuTHQHcE/ekWlha3r6jGinv7MvIl3dIfUZKPp1T0cNrvRAY+ybygm
CtOJ4gAwNqTVBzLktRgy62TH/R1G+CGLGRaqY69gbO6JXeSzdn3qpcvZUKq94o8B
PtJ9uazd6D+hetMkWph9fO1jJff3cN45akn2iCYEtYBSWlwqJWs46AkRpMcdxll9
vgtgdxk7V9pG25vIHVitBFcgWj14a3gqTGc1TpLxshMeARP0usDjANt/h0PfUisf
2FQJxCXrnIQQxzxnYGJsPpkrgmVYRIZIF0LuhNWx6jXoLY1m7eJn2Mz5ezsn/piV
YYRcyL8gKmnB8a+Yi2oLS88DInIwP4bFvcAd92aEdbP4d+bWZr6lMtObH796oJSx
3EUSPzJ1g68ohAoh0pWcaWemWgnICgLnDkTJGfOOh6kuBgZbahKuZz8qIld4TZ1f
DW6CAS2pT+b3oeuJcKCnGq2wH/SMvLMAaQaW9egaabE5FMR7sFw1HdKYsj1pHoQH
DQdbGBSYrN8NWL6oZKrVoRp9H4Wk2CsD5cdbRhkvwMSC+c1sILf4DojzysJoU/x7
D5wlEhadk7YVSDVHTLQsmyY4btnsyxG9ID4g6riCFi04hbSb/fWilOsrRVLvBC4l
gUQAD2GekG8cha6yb+5v/34TPMnvi/pAUjJglXEjWlBS2VMO7SHMzGR4bmz5KC6+
im6LhGFBYNXabgalkbN2RO+IbGgpMXEuT1rnSni0Lu+72UuYa3Rsoi8L+r+AzjgG
5v/JhONmqpbJIelAMPA4D/1JT904zea/a4v5Fr/QIuTRltLPm3opJjl10RBcdlUw
4e5hYZPgBnZ/G4gyvu+Ww4gtubAVPp4T1Rr0lTwMyldWHN/WwQsqm4qO/nVNvj3V
cUS7ER+I9ZzN+rt+COHFBhDGclNCGkxwkHKlTPVkq83a4tC+ySLsWInr9B5knpU5
Xhi4CnhTwAP1QMU0hPRjbg9F7lPQEo0a+7k5PwXF2V149H5b1LfzDmZ61sXgTiaV
8Oz5sJxpM43Db+N8yu96GcCQafPp7blqAOYo0dK7wLEBZLm4PR6z1/9+YVjs+gQl
rIgF15/VUvR6PItDYoN0Ez0R61z/T7Klh/DI35bgiF8wZGWqVqjfN2rsNystQZ/C
OVYFbU+A3+fvLWDshi/Z0ePyJvoPOVrMAJT9W2iBkcmFVuh/26S4pdcMSCNBTbZB
1GJx797qqDSyZk1w403asS17UGnl0j0abMB2Xtevtae7U6LS6teDX+5MXeo7tcGr
Iw+FiurrDHh7d9eFsXZa87ZsVJk8Z9QC6C76zes0qziOn+37FIY74qfxgtfQQ4a/
g3gMWf9NvkVHBA1wvlAlvqG55WltiIU9BIa1kax5R9dy3SHHxD5Ma8oinG7ftlDB
SF20VQCiugWl/l+TPU/GO/QFQxSy+hCYJw416Y8ZzY9Dlxr3yA5DJKIjlqvSNjHp
KT1ctU9eDj//p5PykvbVHiJyJkKilCnIa6kURHs2srTlqqmJy8bUCn7cJp9CC4nc
W+fKs0M793aiilSL8zE1bYeI+HOtL1DzyOGOI78muqUc1JVTndPeHWCKDGGXYfCz
cxXBE+ukOOpfgFwONF73RzhZBffOEpxALgkrnBD/ERI0ut4G5OyK6Zz9RAf/5asD
UJvN7GQwSqXT72FJ39XG27Ar6m/SB4w75FwnJLgzKqkVYJfzPv33SKC7T0PGUOyz
cdE8xP6R+CKtC4aDvG5k4QZfplB7mFDLddta9/mg0ERKFTNF88d1+rCD8couzjKt
jRFeEIl0ecRSusrpGy+Cn+ahvpl73zvK+aXAgXqanXCmYo5Ag9uy7YKSPEoRBdVj
8k0QW0uaSrL3ZtnF+GMpAMZs8QzLcSg+ArPo5REXPaumc/L7fEgJMISQia+2wbzK
+50X1or8CiODerpBCKQxE8HOPBT0LzMoECAoJnwm4m7GDDznN9M481vpzxJDbqji
ShWgiK+UEv4psrhdKKRtxLs1P4z8JxBBilu/qq6YRm/Td2dIK0LsA2oFhWQ/L1Mt
Ev0ynvki1aL1HPXEBc6KiJYn/wHlIYzLOR/nWINcqxXfGYs3mGoSm0F3usFOmf+W
VeUTsR8L8uQSXuH67f9y2egj0ErOhhNfOfkmRxWjIVo3D9NNc6QHIAXpt3wrVnPd
sndbLaMRVhsEZCP1LiEt+CmSX6L2VqaV4nStdBvkltOlW0uKGMzeh/AL9Df+KFwI
8eBsq8zSFS4vkMiHYz+6PhjyAJe38CnLWetRdGTVmyNRgdOgMyg6uYDmWrU24hzM
Mk6hgkQT55RZbrPWs93CcFSrW+nL7Dy3tinL0DW/DgZ53akl8Tl+LZRoetlWAvXz
+1+d8yPpuUaZ9RThPUe7kqXXEwQzvlhHgCMEfqXw1sivJSTE0ICkXU1g5rC258/G
TFUbR/6XsZuyFJwksz8qBrCwOfKPr0b9VYjmMos2Lh1rdsurapE2IZnxalYzsTEd
K550RoCMes6JySunmxisbxRO/xGJLABQ4sj6EgpWo9wDfbxLKLNv+O3QFS/OTMax
rGjOS9qeHJlFl9LTTvuRgbHEhOSFRe2wJ8eSrx2TCBGY+BJVVzLWk/KLbqh/YIu4
SGdBfFNBqBF1Fb5fCCUbj/8YvKqzzszq7FTNrh2lqEjmAkFqC1K++4U77eCh8A00
TMCligqVjJUeo6ZgVBE+DHVDzZD3ETbZ1yYRiOH9wjzTEdyZjjkaF8jG42fam6zp
riL85XMBT6PFs7hP8qOJHo6tlGxXCT+BP4HWZjD1XV/29m9ucRWepLEGoNqzYIja
55/mjRY/H0FeVANGGTKsQgelxKpAFTpCM9AQBPJWNTSSrXvLiNduEyAkgMwPwTjN
Ugxu2+CH+5s555nMb4UylvzsHoTuIizLmyegRvdulvGj1pXqFGaBXBqFuZb2u4iz
8Fp8CHFbgqIBnb9fsg/+f2jtrfZ9yKM2WsULibe1EEiRI8hyvlTLB2gJbjc9qwe2
HfXyx+QaC/wfDQ1H5+da9crkFfKQ8VjLZJqSp2l4nvXsgCp6uHa+s3Kx8CQkk2HF
9NVL2DD08nhCKj0p33SHRK+irb5N/JQMwVCUWcRP8/S3y5Hg5s1W7ZnU+6w1wJDa
y5vBAUQxEGlZSQ6aho2IJTxZVQMZwFAl2RG/grurSLt7rGuG85ZofhFa7KHQIiK/
3olHIQJSQmAAjrQy0Rc/7mBMC3wClpxl0RctCLPIhH+PCzRpZi525IqGnTpW/bW5
wwmVlSRCCpFQQ7a6ZPpUWobUzkcC4v6aWY7YAhLNiIeFT240t+k+qkA78lIwUwYt
gBNYGbr5bXwqx0KO9bPJ5vTUuMF1TxGuaTCxwGKMZgfHcF28bHhHw4GWJh6VZIFl
biCyxrE0Fe493HuZEeAbfNyRGhU0pUUDW/No4x80l+7d/+mifVSCj+ZzLVcgswAr
HxbSMuuCwLsXlMF/TWdGrQZtosR0k2tEkeZs7rS0Z05nQiH6XOAp5mjfT6a8ZDYa
M0I5QB9tKZCrkwcikdnt4WZA4khGBIT69R6ycVYEecXzyJY2d0qbSGUDjde0uZMI
nncQIrg5XA7eFlFF/m4FQQVEHe86WQ9jb+kwIileREs57qbNZraS5wdU4FMXpVLN
RZwnAmmUHgrUtazJCn2FJIqlR742W0gK7zjyI8ua5WxQEOI6mv953xuJkUkbxrzv
y4tT9WvsR1puGZIVLMKfhAx+CvnVojVaHf6rgBVmLWuLR78Bjc019GCjiSpDPWcC
aLDYHmjQckRBRugZmylAnyOVD4ZmceaAMSOtCW2r1UxsmSg4yX4//9k6D7SaILIb
ZEKmLV+bGwy4y9adsF4PSjv0e9Y6zrWADJgtsj4HQdB6YdTDJ5omCYixNuOMVEYj
Jy9ma4b/X8OBZuAfESUEZwQ7/6Ix8H7uq7MgmFRSAnxJM6lwvI85M8V40Rej5yTX
cgpJztr979VPhh1ynXnKw7spi7dEaaWFKy1oCdF/iu8wPgKOE/OESWZu7ud0wX2l
4FJ6wwKV8zvKdOoKdT1+NoqyeBZgm7gLtOMtSy15VO8wJJN7NL7ILNCKkzRBG12k
F9hQ1ergmM5Yg9yOE8r1hW/pwiJokx8+NBvlZoSn49Uo+64CyxR6sLr9U+vf4EkN
1kRu2w9vm7TL/cl05LdAQ9acfzm7vViiBE+WjO35qILFszOQof+kLa7BnNoxUf1J
lTKUdg8t9FW67ThuMAsoz3PL/+TQgcBmk0vRrG55F1mLDpPn1Gl7cqUlIKa5U/8J
jZKSYKWADo6ZTAG3HE+iIBZk64i6tdkSKj++z+e9L1sbu0Lxdbuz4bPdhiDZAkKR
tA8AwtmxaIsv80X+kGZ2wEa6CDWCj0SiMokK2sHLPDiqRTSu5O2ofkZEDLYL4GIn
GflUTT8KgEk9nM1x/GUt4VEEkrsF/FZyenqh/6FBYLiIYKiSMJWXEVdIhQRK82Nk
y+2ybjXPvmbDVavQJtXbfF4RcyUu8dzEJA/fg26xu1e8NrPa0Q0pp3W4PCpoOteV
ppQPfoR8MghuGJoZJyfYn/mHLJMc49rsvrTbSqiaN88lAxFOxMrfLptqyzqylqau
b/nBmXtaguyZR2Jy67dK2kumSLRa7Y0MDRqhcF9QdVlTteyDOJkyktJfypYUhzIt
qlpa20DuqJGpLw2pNsC0F3zFVHQjZIfefqRa0ggn2iQlRcLhmiAX0BNJz2QHwjIF
XGzZqNBR6r3EHBMzHD0f4rJBMM4Wy9w3NmK7mXWlq/0bXyZmTIZl2HLUFTNyPdWg
ypeL+sGLF8YOS6myMXGnUzjdXmJSbW+Lx9rFJlXwGctINEEtPSg484WwldYc9XmB
8Gv+7N0c+eIoWXUhvLLhkv69pGyEV76xO0o/aXvyaGdwaK9OltZE9eZnBKonmMlM
omqmunlyYuq5E74PQafHFJdcdMhGvW/0Tv7z8Fni1CFU3gWPQRRdZKPFpV10pP4M
u4xh+faGuxMXpSBXR8NI75abpxv6upiL2ebc9w9Na3V6d+W6Fk1EMPOM1gOtbie1
/3/QGwxnrGqlI/eKDtjxsLHIVqy2CCXmbTnzrHBairCzvFnA6/jFsI84XFK2ngF4
MB4BSl+0Yrhcqnqyz5f8ksIXM7mIG5JJg6BJmNFgkfHth+awR/z7NgUZsuaqi6p2
RiW4FSZhG/S/jE53MWxXtCwZaTtrAwWiHoL1AtWvlE8MF6OTM4JWXBMAAAB9VfiV
Kd2hY3roq5TGG/7qIxYiez4BR+NAnqAiRPCKfPQbQ75j4xUxxKUNTy20n+64VO6M
ToMnvICJvPkKYhab7YwV1JnNb+h0lvC4V09gW1cWp/VB1BfWV1FIiJh+yHCB5EuH
yJzhEKnxCXkWTBdvS6LywUKPIoBwyC+0Mmk4cV5EVRtL3YckExXaFlGvwBFrxVB4
XBh1akguTTD2gGqT80EJ9bfNEgqcWtbIyiwYdDqXaqby7TMsHyWh49GdkFCUitvu
PJwoYtQp5uAozkvdUoifnkmtkNVsqbI2Q7eCHw2IBFgN5NcIgzLnUCnFsfHYlPsU
KoQoot2XvYw2ImY4fi4HIPT289qJFdYkkwbpFJE9lKpv6cNBbIoyiK6bJCWmRHdi
alg9xaJUm/331MHyHP7GI7GUaO4+hKTlvtGZ9qkBLDWJ4fzOJJ8fx3Ewpg6QWkQ4
YsdUAui4akD3tmktgVT94W5i9pDC1ec8h5E8XFph1qO4ih3dTNn5oOGtYP6hQ4dI
Zrgfd5+WMo7/MtSozX2bbdcfx1pZwy0dYjKB1+x2ITQm+II0Sixg5jWGED30qdZs
slbp8f2ArvaGBdVJgUHRyn7WD5Sm2nGtkw1wGwEqB7qdWGphqcVPR3xE+khPDTOe
58TmU8SFAyaTiEuhqy2gheIDq8Qaz4YblkJSC5tiLL2nfp5JTQk0Nrxca3/IlCgl
mM+l4sVCwyv1Fi9o1m0GFKqNxQuoE7WChn6GT/Tb8nUJ7n3FV9YN6MQhZ/Xch0uR
1RL65/ZUukWhmP9zfZGg7vAjHxo3qazuWF6H2oJqryQvuoF9J7B2dqucRj1WXbjj
gGguhFwYKsr5SuhRWPgw9Jrd+HlCZAete6vn+xh9n/ttB7yrITB8XMRZFqnZRmaq
2S0XoAqUXx/8QpNrW7NuwkaQKwlLUhJmFKA5wc64FMeaM7a3gP8z7HhAOy5Ywjmg
kWki3U8WoM92mN9mB8y5Q82IoEiDAKGwuHjWbTFSE8oTp5xCmx4z6dEtKHOKp1ju
6JgPvHLTMkPeePnn2Q/EVPSmuTFsE6qAsXlhzj6vwAjXxvmkelBmHsma60qFZeb9
flDWPTVZnzgRGGMyUw7qGsARR/jrJ2FeGHzCcau8z25nINHzgNC3KKwvn5ORgRna
RfsKTcVe84kGwF77yUWewVZRl0XjEiCwPQoxe3Ep3PkpX/NmRaY9GFm5veuxvZui
jj+5zgoUmtY5E6Lv4+Q5ttXp000SmjpgWs0bxLVSnNGiblZ4P2JwO5sMtkYgtt4b
PlDtvVme6b/wwV6/u7O1JykqstHzCBLmE/zAkCHAK34f/dHFbQGhwozCZsDeJ8H8
VF9rtLyMPISO0ohlBlNu5cbZ8ZN1mLSsr6/IZklh4Ps5jlQqUFwH3V4xYAaNAwL0
qwtE4wPbCrQyS7fwVoITAY9rIBUFZBFo2jTKUqCTXM3drFbbEmf2qHn53C30qNUU
Ty8DHAsUOC0uPfL0JTOK+YVj4O/fFoZdNJPNjETWAgRp/ln8QHLTCBDoDFXru5Lp
N3m9VEcA7KisAVoE63vmgllFdGICxEKw+TK52jt98NQ8sm+gswHooPgqehfgLqu6
s4eFYIL4zLkzkeTiWOXo0Kyl/WpZIprR9fYRlcrEdqTZxThpBB2niFSYUm77JHoV
z1cnsGgFVwW4bJH4ZeU8PuILI1LkVmibOeS2OZP4SrTuv+t9U2UWVzA9CIi+0BOA
c6gayOmjaxMCkXMUQK/CwVXYC07Dat+UjsML3eZuy8Uk+HrkQHou+lv06vDD+3qz
ObKA7rny7Ec1hf5Haf6GegdYOTfXkWBDEVNBNDCYVAt2rgLrjPuYYKdD8kEm1PPD
qLDE31emB3DPTm+04dXP4k19e1Sd6pNxAEscikiFxmRWB+OnMXFje4Id8DZIOqlx
Tpiy5+c9pflZOowKgq1GsMwpSOnkNLFP3qfXbszDuOUS7HoLkgjL4pXouSoECoZP
YXOqAfeNOrcgpuqsQIOdXyG9BzIQ5Shkitho+g0Mx5odKAz2B6JnldnLYqVavXZm
TUOHSUEwW+JnMXWp0wySxiL0wBnXIgX8zU5lyon7SovMBFTLjwjmM4Ja64+xB4sn
F07AUEiWFZfPgEV9pL4iodqcpPUFtYSkRv0fepymVVXU9bqZEbLZ12P/Rru91xIv
45+Uhg7bnWFpNrnRJFKQDHF2xlBfA+1KbeXNT9EB2aUfcWtJLhWggi7BJOcDec44
Fv6wY/0Ltpv4ijwxeK9QA12z6HG8KyspH0CL/TZrKd6LlGXT4Kvu8x+reTi/Wq8J
YlTXHVtKrtzJge+fki29NUunbUUhSxyfC1xyXgIWUQEsPXuVnshkzX8A9J6dMTyz
cke6FUyzHFOwPNyMmxjrd5c5P2jOTFEc+ud+lR46UO4/Ld3/sYbFprURIUtGjjxO
Bz/pQ+XF/6karZ6r4qRBmpr84QmVPu5sfn6Rl4kKfzd9tIhqljKMw+mdkO4bqEna
WyCiSB1LTgwfJUX3AsDr2SYgK5MwD5oLdTuy8GGfXhR2V5IqMfllsxvgpOvbzXLT
1uqFEEemYruMlVq2xGrQZZqz+xXGnLKJO8pgNT9kVuFbPcNZlS/Y9mdJL+z/SwaN
tRq+msJNof/u7uPwQ6on4YpesyT7NH/Yt9JSnXX5zfFUoxpKVeYz/OKZnuH+SxiX
saXXsCbAVmM2TfFYEA/HPu3HJitU/bXwQq+dxIXa/XHjymiOcT85JMrFoWM+rA3k
IrE4emSh9wgio2LS6QM9fxZ4a2N546Z7Ct01t9yibGKP3Fb+ZTUiLgGR+HccLiiG
OCRQMdriNPPx/RwjUzHlo4qKj0Eb/cAuAYQpLe9izfBQaarMH6LLoYfg543JpAxv
eNQgBo52Smchj5zUwrMSJblhL2y0ybcXQJ8IT3ZS+KyE2WgoI3jaGaGtJdU/Nttg
fXU28U0rQtYVghovspMrpT8hlXWtvK2C25RB4C4V3QNruDKyX01G9XE0DP3O3VW5
GkRHCE3rNGugNz8x9aIMQc6jz0NZWt1s7EPvWmEsGuwyq+Ef887aNuWK9AG0OO9U
7LDo2GVErOWxYx+wQWmfWg1B9n3wwtSm+aGUiWcbne1/eLtLjHnD/3l6VYl628e1
IaN8VYqRqXDHO+NThZHngRcw95cL8KWeMjS+3uhOo2/Kb61Of64uqIxElO9eLBzg
sejFOAkKxrl+2xDkGgsAMO8X/qk+l3+AIxEuUsJNQvZtVqEQOgNAy0459/iP70oI
OUdHLeeSkZoIqYozk+KCvE++DcvwBCC/1x1vOpRt/VPaTMDWcVbgR8lX/qBdPxjq
B4RxrE0wLnHY6Eq6Z1CFsJOQZQMhTtbajkoCJjndm/YnRTLZtUsV5E7SiIqEVjyn
aqCKTTAew8aUfrAnnWADTP86aJe8cIG9d0i00j5hWVBkwwlrZsy3xO92d5R7bqKX
8nC/wTcOlEedU0Bqi2ZG6yRM0GXHHkUTuqtZRvUw8rdvmo6Bmj+gE7RgFM6afrND
mN7c8/oS4LtBszEgE2BMT/De+TfLkso1gELvXwfOyKzsyouEaSiyZDXp4Ht2MYKn
lR/YSnUDaiAcWUWqcRQ5WrfVdQk+ZwUAqpNtt7ghGS+GaGmhSuWZIme3H8EJ0VjA
q4Xzoo+fUtCUjwYiRoAyOhtC20qXs/XrLp5gibQaRLnqqROwUe1LbXT6THoFBzX9
z0TTXKxGq/u29qYnKZDwjrz+vS+C3W5vpSiPbLJTm7IGQFqgzMlGU88rg4Aupgu8
lG2wbUEX+ECTE+ESzHcL+Bm3gM+tCDQn8tZilXTKd34Wh52VjR0mYLI7sX+QyfHr
9T/iQP3Fr9LKGircPT2IJDXbPd7fdwtcUASS8CL9n6yRQV9B9zTny/Kz7BcXPEaI
aXx3g0kLI6/t5hiPpRS2vQE7qY8+scidPgs/UJrwh2TtHVDnEDiR210LrE3ijCyI
mVJpCxqtFCNFh6GxEg1fixRiTbsHA8n9HrEOUfkNHcKgtueY6I6Oqb1RAyofxG8i
+ci1iN9oTiQ3q4nw0HV6Qn22Oc02T08Ryu5D3A3jwl/8Rp42zR+xpaAkLibnm3W5
HK8CdqUuE3g6vtLV2/fNtdY/SG6oRvhoVx/ioplYSkhA3kldkCwqpO8W+DheaSps
GuxIoF9g0NHeZuMpCvpkmBt4XfUaz++DOA30/2s8NpEqhXjkXFPlpob/LRJ9M6p5
0Ptchascof/vnfB2bmafI06Q0N3AVzUfdkHRNeznCvKXPk8KyeUNb4vh0U1cUIfB
6Dg1WQe/N4HeA25fEzj1FzZRQZXFxRcJDh1MyPVencvVrx1i+2FSNe+h+o/LGgbn
YlCvwhquR+bDdk6ueFz3/ppuNMfkkf3R+M8S19a3ByVbjAnjz1IEawjEKT+ZEtn1
XaTw8g7FTPs+Lf9I7ffWPhetg0Q71ZocMOxLcL6Yk6o4mH1iRPoAk0jczbM9FwQj
F2H9XxmjwpfZi8x2c54Qr7FzZ9Vg4/99OI5OzwnI1hEilJSCnXzucXZ33O3tukxX
yvV8UZ/UXTEXtDA9jFOt98OxHTyCkIABSje0w5eXApJNW8BraHYA7qJvgbVYChZ/
7HPOXAfE0k2qmMzgV/1zjD7+v2JJ9aQKn4aVt3+/shPRWXfYuGlKNBQw69CZIL2S
9ecmfLJHo1ght55yTxhwUBoM4Bs56apj3f39sWw6qVgNsNcTGKvZupw3GiWYgxLO
k0uPd5PcFlExlcZoVk1j3ftlf7YjGfDkBwVqS2k7wExk34JGxw9oZa0xuAjUvRcF
gvOLOm1ExJIqeNUmSOziGKQ18ns96RF6I2WOE18pZfrm+YVVgHihQt0vE+WJ2AnC
/umSAUtKeuICzIEKjfBrfNP6hjVKhoin/rcTdgIyqyZu1WnQlQrXmnuKEUoX0cZQ
6DXm34gjulw/KoGeftpEsD4xKi8ez1pK43EDBBFxnADf/kyqhwCj6kG2D893Nn6W
ws0piipDNDgpQtz4Kj3pmlKELqLYHxwXqBd1IMEu/O4NTcB7UAtWIaqeJMSgKyK3
AUz4upo8KZtRd/KbH/gkEg0a2qms0PGOLUfMUlyLvnLwIH4Ci7JS/37hd5BzBH6G
49LwHxbeuwtDaXGtUdqTSOB0q9b1S7plsdkK4y7CyNpHKfdVuSOR0nibSxaIMpsX
GVTsuY61PxGCwiMwg7g7Mj6X/CZuLmVViyOhLdDC+dsSLaQxXNCTSWoryKQ4nD3M
/ctzLbtFyK+hp9xUdYRlITA7GT0xBw6OdQVV8JZkHHYqkoDlEi+TQgQbShEIbO/3
ZbF861HMc5mR/CfmcCwkOPtFZXy/YR02Ad1qPt4bvgBfv1wfaDSZjMqYgYuwBfU8
YxeaLoQcLMeajvDUe56bKFS2U1Xz1GOYaMQmOwLTWpckEJUoOAX7d/q3/d+ZlOhR
With7G6FDJPtquv3P9nt8tOaWYdF4BswuiBHvhlAUKYFD3sBOLWA5y0iFoYrR/70
ykuQorZv71OZWcyOXytgnmJUKHQvkuEosxjsqo5lcDijm8DJFmwE2teKkLNrrbhM
ES9qIovP7wn7U7Jbu2QE60JLKRQMr3NbtTL8zRxOempAKD/IrnnFQMdJkStiZWZb
BTqM6RU2aF9bCB0rQaGzQwm9t9dyP4jy3wNHwwpetnDPRxY7eDKbWl9aJ9UfD3fC
mqchxKkw/9GFpgH/u1kPzUbE6zscRq3DNvbynXi73EEXRNvp2pxXAbjnXHHffv4C
FzTUn7uB5LBEtARXiHRCCIFWWqbiN9jQfYYckQr3U5yAOmjA1J6cSezF3BRhWAjh
MRaEUtnZY5sSNPLRdHfcV2U1Q8aX+6iOQJuaZPPGCGuHKhD3Pr4P7kEy7U06zfmC
0NBxv0HUXlptRiThKgqwwFN5thugU524Sxz20h1RsqEwM5KJ4ctV7ByKk41ZQw56
9vEr1OIqcjhjileediYiu928isYYBbL4mfmdw+SSq5J8IrMwMa7017YvkrNdYFYS
6izuHgvijWTfm6CAOIFsZGDQeC3SUVTdmYxBG64PYnBwWHPNobl+DyCCwEY4nJRV
fdF1dYCUUPx7/y23Og5HCSONBr5XG8glJm67P/mVSEf4P1XcyDy8bfyXikdNxQBV
jTkRut+wna8SuD5i1Mb3R6GuIUIPq/EpVlksIQ6w4EftssaboO8aw8IlqS5ooB/+
mE0dBx/MBwDgZdUEdT9MHNwpz1LyEka2sYadEcFzP2rFiu3+vnZsRKxt4K3KLwgg
N/a3ojs1tyaqYog5r5cXy3HAFBmZ/0OlvlSoAmhvTcWp33AGvoUxZAF+HPQx2BkJ
1XtK+txDUEv1/nugfBYBhiuKAwxaDifIRakICHoLSg+GamWj4n6q5/ud9ZScz6MP
Evl69uzsPHiEB9Fwv6Tr12v+O1Xe6DZl2oi8OiMifcEFkKdRHobC9t1R6LD6Iawr
29Cd1fuhuDQtSnueoUOvP9wMot/TvDyNPyGI7SL/czKBGpZ3soCDN1kfYg2zP+BO
k2E/6aXzS/rTjNsaK/tQiRjLPNwP2rtZ87xt4Ph9Au3vMbxxZtdx0MD5gRxH23wm
FwoHzizDMpBc9xmkvX3gHuUURGyiOidA0MM/bXIGcjRFDI7itJx7mqky5gsGm51C
PBGQQBsGyODYW4stqVhB+l0fwcxTo6b9pjFVQPadBGgiTHHJTAPkShvmd/3vxBJg
C+SRcO+6EPu7KieHp1xWbOuT2J9dgF6AtDIRJBkW9RMLtDARnn76ScLZxZiT4xj6
aNFizQfOjqMaOSFX0guAscn1NkTMkN4PzzzFXYM0MTXVvuGkKvzbOmFG2XExACq9
hCAYzXaI6npUw2CfPwj5ZFv6Li3hNjSXAARqM+9UnT7rLPMBbmXPUFxOwYb+4l4x
t9AXb5DDvj4mWwc8fpIpv2JbyoBQELFodiOCS6pnxQOE8SGDL4Qd1QlOwbVGMiYk
WjpkovAj1zNXcr0JLNO4LwFkebFJlwVm6igu+UH9YR7QngPZcHb1inHcYh3QMqYc
YlIrd2+NPxO0/fgTrIxhkarr9KTpjG3ut7BnkWvFRUPRq+SZNY2qE+ig/xSz7X14
4bKWJhM5XxQx/HYSGotaiaER+0qKM781G4xm4Hqb638a5i2yHfrFFvnMYejptETf
YO7pzOPIYEcqHRRCVlZWYp6LW1/nIO7GFW5uB0K007DvdOUjTglq17oWGZ1Da/R/
jQyANsvWnjV8ljWreE26KGjXerq7/gjJ+53sOwfSC2t9PMbKPHSCmpj08A6/HVSe
GIG3E9o+QrjjEoueB2V/F+HuICCVBgjKo6xeeyjgk5Vg//amIX9vt7NsVsMNNUxj
mtIYEePuLLJnxEiqdYfSLgfzOs4zHDVHy8O5J57Ku4foP0oJ93cOBNqYd6Rv8t9N
9JFRmWEAEfzcGWF4YrP3Fc9GrhwQh8Z+Tj8ohb82euUD4crEQIAfO2V+dh9gFmgG
aPEh28s8cPAWgplB9jmjxxDAUOv6v9ovpOuePF5qZlqIM9pQKO53odGdUxfdghhH
fu9bcuMtCHHVXS+qAksaPhitvPaX1pr9VbUxEkIX760jB04vE5ir2Ix8SX47aMh/
hxPNr81vbrQAIr8hydvLJrSl6Gx54yhZzxI855tVzWqtsFxJEuibwAiFUvdPuxPB
uwjzUvIPZuYbdwAYI752TW+Q2Bx6wGBpq9HrHSs+fMqbqbu9nv0xs4hX8u6qqy5w
rbN5aa7RIiqEjxMJI7vZ0dugizshcWtQHTQ+2NwcLR63Hr8jLxZcMlNHIheDu8Is
AbzeOzY+Q0qBAkXQksKF2qrEHgapUqllI/CfO7evj17syXFvnBZ7cmd3opiZAguq
wgE80SdM/bnb4ySN5k5xi+W+mkCJvTEPxkZ6xgn+c1uZCjWoz0fcGn5JIRSuQ9nl
CJhVzpzFUvOWf3FnF70509bQO2wdqJxJrZrBm4toaQ7KzD1CJSg4X6FILLjQCyxa
KJ9LJe9t7jA12tC3+yC+FJRztFOkdsz+tsCOiogjYLMDgr2NWfDWXT2UtWzYmwNe
NxWCqUJhmj8b8ucRPMpXmSqqw2vjFFIcVadiM/qO/sVR2EmoiPvTCl1q+PPbufwG
iqf+pxwI+50kSvCAXEW5fFRrMopwlcOWfKI1Fvwge7AZIxeXVz28LrjDNr3pePTp
y47s8bHkW4IbjNRQPGHNc5Jc5LlfZBnkUhOlV5/lNRqxn5FSnlb7dSnzl4+hbIgO
3CeCQqSoXRSCkMnB8Zrb5DwldrG9ByO+bg3yZSjW8ra/AW8YxB+Ah+9sTVZ92Vjm
Zb+F80E0G6U9Tl0aQ7Wq1JzoUM0kETbkJ4GcPKwP1Be0cmewy5gWSYfy6mM8VdkM
75yeqTXoAibj1P6gIX/9yoZB9OQzwguBApv9Y5BxqXJ6NNylq20MxXV8Zh09BAwX
4C1iQUD+BBBMg3s+GPnGutl5kH4q+X5YvU23a+edZ+zjH7e/6ECqMtNaF6RqkZc6
RYlGhVs44RxlLzrk1vC2fAnOQ5OnrRFB21CEN+n0TcUB5hmqr4z75HT6NzdvnY2z
tK1iFW68kml5lmvVDEI40qBpmNbpeLdrDetf72lAk5oqqrLkrePfpTjpFhEtOBJG
BEs1F5l42QA/Km0LHURjSfnIUQA/GX1fpiCT8XrUjTZaGN0OCgS55OKc+CdTlFtO
8BmdHCDLMlpqBkzoVRSqeutobtTr6I8Q0pT06ihBw3y9PG9B2j4++22wqq5nA4zQ
jkRNDFsLTWLvrNiRgxLXA7ta7IimSyFTH4jT7aey5XRC414ym7EkJhIPImayZhWO
X9wsCZZEKK4tL183lC/kvfdL3EWXogLJVoj8/UNiPjEDMJ1ERRC/t5MYdx11lh65
G6sc20To3bkNZCPicAMlRakHzxcfwAfAAw+j8BNQMCvNJCNNwvOmPzvIZjAxRquq
czI0qMZ2n9fjtZ0iHRAXpNdAOYxx08uP+cTfnOabSpAKCnDlPoFIhZydxw9Q3FpA
nIZlIaCk98ayz+oRVgUjCoB26xG/csujGdnO7T+035AtJPP0ZUerftx/JSksCTET
giGAjurJIV0Q6CNAUrxBgD/CjDk3sFjmAa2yVU7V/rpx/BloSyZVHu9P8GZguWty
RU5drEnW13MX/MtBS7JwDzFomUB+ggXKXL75W+AGHU9f6tqt4o70hU4muQqLGyN4
5UhBsA513pPTcVEk8/3H0jOX8uMSNd0JOWzi/rOKGTszzLa3tMonMoqsx+KUqllb
79bCbIUqI0OzwRn6brNJMN0X/ttKmd160I5sxBcD0quflAGQaHDPsLwq+Z7oYaJs
ZRJuVBGLhYRmpD7ISu9ycxWxqjFFLNtC+b405N3U7rsi/USagIkW24SXLaPdCw0n
6L2E/wEEP1JbfTqxTOuRWy4mq4fwuTqwqK0JBM1TlDgCVoQW005Ql7m5+gJVcuaB
Sa39Iyrat3VNqisAFhF6QGz03bJa7f0iibUlrUwbD81fCYQB+SPKoYhATefiQwnh
kYnsYeSvRgR3PZJHbpWA8C+EOhuWnNmCWt6iZqvIeJs8PMPuOtBPza2am9AAhyPd
KHXpAUbHWeYwSSm/C7ZgsoQctYwDHQ57yk213HYlN++KSDGL1eh9Uld3xARvoNI0
1kyZ4ZCUlVdO5NzUYUzTP5bmw1SmjfJu9DKX5w0T2Z37YR93ZQhjWwA6QiYi9nnt
hIurhNqTkxdPKsCSyoW5LBs3r62AnMgkcIZEkPNYfOt9kXM+0fKyXA8WIZEe4y+S
lJ9Vj7nVf+jdKbkOwYAal3bU6c9buvxd2Tuc4jJqpcfqXVlGWcUSxns/0DZeTM6C
OigPw+FQOzJbLNzUgyvkKct/qAlXL1ttuJyG3eIi0Sj0tDXEkouusJdUByecO3ec
PVIyMImGF2y3SR6H7uk5mbRX0lxmgw6KxMgeLctMkOxC43hE/RFP9np+KiL0XInR
H6qOBt4x5I5z4NHzhaPKEqsu6jhsAr2gocWgFY8YPsFJcC8+95VOuSEaEW3E9Gw7
g2GJ6y8fP3tMPyqlyrMke/pCqzuFHTTZ43DCnt0xl+HX8mOebqvFTm6H6ixDNRQK
tNd5L1fctETHuk22qilKjuxedYkIn4RJeIuLt0FxCGc6VEai+JGmoZq0nin7LPKi
0eDd7QmUe7qadLxI0dN5dMQQbKKmnD2dDnVpycpS4x96ZK+Hnz3g/POq/G4OvKO1
/s+DXITeBq7W8TiN3b3POsKaiYnJCkLAhHKk8HqwKK5j1xfE4am6YfWr5awOT7fA
9E7TfZkXRdwv0NIKUgLOFLb5xpCtVzhJz2lePiivAae7YYp5rqVWd6dv1dKMiaSl
Ba/IAaJWmeIb4ExLdspJmeM4XZ0mcBTuuXRHWw6/vIl4YXSwvd161VP4IDyLlzZL
mRTnwwtcYnqNIosn9JILnb7yRuts3y+S0/MdgL4n9XfhVWYLiA+5shuQKohNH1Xw
OGeDYS/cbdl+oOjCIKOz5HykCpwxToLFvHkpLmEYFAT7ug4e34oWfMxiDmboARNW
lBXlM4Pgh3C7lIagMpEmdg6t4aLPSH5xb0FXh8u40mX19YLUCySSqj6CC3jJI8NP
6BJL5Dxr96R6d620yALlVNXGNR56J+Qk9VOdk5Tqhs0zYZeAo9SAEiLdS/xSTUxl
o65+LFhUSsv0hy0v2jxDam3SkhkqNAnlsF3afgMtI2FDLbsHAyK7K2Ew/l7Zim26
u4gaLXXlVvbkB/E+m+cLgxvMOBjQED8Xbwng1NZ2N2ZfcoA4cxbCal34czdYk2Y7
7kazEc8J4OsSZgr/6Pb1lx49TjZ7LIT2OPPUzi6GwGguDSgr7YKpXD4qOLvM60Rl
1aLRxCgCsoGwBthrFzCjoidMbp29SRpXHZfHQkiqBWcAo6oXoPC3x7PfCdnc++40
0pNlDHp6mfCXHAOh+h1M1Ag6zMupe5ROHnyec56JQlaJQWFrLysJ5O4lhia+5l5Q
I28Nzc3sS8hlJrhl+EucBt+52e0B5GsbMpWCkBEv/BTlgPxbcDGFPfp8+3wzwo/b
c5poFluMlMoTgvNzg2q3nYBq1hxKazYOvt9yBfzzJJJCuD5GIG7IBJO2yrXcvXD4
K/oaW6GlkFC8d44NKlOVE8wPmUO9so8A5QFQ7WCAwDMr433mG9VO9ePBH8vF1CiL
UN6l5VeKo/obAz+Ozqfor92DMcRbbVBMbCGecG6Ye17tkD7c88Qonh7qwY7skkTG
DXbz1Inor4aGALRhmsj8jyIJbigW2m80SqiidYY7siCIeB5Lu4drsDh4N052iGwA
5VT0uYjgcBtaijSiBEK1yp81rWZJOJckepg3ZZHh/YPUUxFl8FT/C81bMyBioZOL
5IUqsyrVxmvpfFrAdbeWKV38e+pJi88yRQ42STGcGZgxte2ct2aDeTbDWrrWsSSv
y5rytopldvl4PGnx7YOjxSl59vRWPLdsP6HkjrJtCX052u6VTkDIgoM7z/O3Hsq/
RLCYMydPrBMxHJCcjgnhy9tuKk/V9M3XH3e7O4NFgDYW5MoYab0lMOLko9LuCpr7
dIatPc7aCYPoOT93Ark/qGFFf5RqyzEESJJB6suSzwBtgacKgXGyRmMMAUa8sGZt
p61ZtEyJ7MiaUSuet5lQU7pdp7cOC+b4acN6F/H56oqZvXgsAirH9aaryhU27CeT
082pgQFZO3xfwTE2mXbdcIpoHcyheBkvm23PDXBXsQFIjg1fT3OwdCSkVQJC/v9/
wUpiiu3ZcmPg1+GFEy5MvkSnG4tgimNiULKZ1wx6eAW4FvvuWZ0TqZb0ZxjF1rxR
mlKBzzc+FAycTQDPY0lEBCaA3d+nkHYdHJZl/ID6POJyEDrBUxBFDgys5y2yR0Jk
l/Y78dBBljGjp3CBM/QwZ2rYtJ3unX8Rlyq54us4s+9A01kv9lIFKml4DGJLgP/y
SN0buw7P1Y28IQrZvcu1prXrhe0An2klXBAoFRujze8Yz8RoA4vjaNDJtpTHcjDz
JkzhKi0vDxNyfpb4NYm0ph98dxSB3Z7LXhb185P5igfVTZUq/kl8SbLVSOzTgZ5C
OvhvFUTRukk/9cwctlcDxUwOUCTcmLw0RuGBHjjYi946pYe+tz9v4i+ciTcW8Yds
3A6cKDbONbichbuYos5q5IB0B3brATub0yyKEw6QPvj3HuGFH2VaN6CkpR7lCORf
ehIBJx+7wiKyAmetp+NhsMkgWQoJqnqAkeikA9fyEr6y8UL0uhNwiRPb0e5R2hwr
/QyHNOVjlmweFTQ70PaU0cKs/FFr0VAA4pkt0B+bjlIqby9/UsCc2cS7cHTfA8xc
jku0k1YH1/a3uhP5qoIfz3YZHC8bax5+Axv52mJblXzPPvtG+LAW3aSQeELxnSTr
XRCowITGteE8CbjsBW1YYL7s4p9J32gGWLt5CQBWV22b0nXed28tM4qH+/3t7sbY
gyarGnC3yFgoYmSVXXhYjOZwPPKt0lbFOfM83t2d7Mk0QfNwZd9hxfBGFLX5I23j
iJR2iIbN7hDFEMfRmpnn3jUMRQ5hQsMwYbdNt0Mg/T78PUkw1N23H+PW5eFFZPZo
m1BuX8j4sOJ3oTgIwUm0M+TS7M19fZHuEN7rxKraUjslaQmOpGxMSwvykikFzPiC
cC9SqqwvBSUsC7S6142BHg1JIeem1mdWUtmzLwZV6dp0VizSF/Ec/x9vLodITLW2
M/0JD7uVGSobBbAQ/1ww6HvJHlYrIJePv9WiJ7CZ+o7kn1i9/vo/eMsFWfth6+lH
RsUrRP8PYVG7DV+j0KNbK4LSySvW8GhIA4vLTOjKk2XdCqnsuz9wYWOEoyOnIfET
LMBbKe+LiYYfhZj8WoQfCojhBCgFIBN+X6YEUhKv5dpsWvNenXx7Gsh3gow1bVYG
sjkUQD+noAwTl/k1PMYEQY8Ps/2Pbj4cMdM9PO9cLzTKR6BhfpAt04bmfFV/tWOw
VOwcNQCfY07nmCcKlulcpiTF5MfRZz385GiEJEfVoVcYJWuN61lwVWa9DWi/hqNu
gvRWNmf6mfgpMInaN9WnZgbvT1pFC9/HOkwr9aTGgckD+CL2HFmhiIqgYhmrv+k8
sNkqt1MiwsyokNctIrmcBbxqwQ3Xrsv+9homTuGWqRAl4CZ7V5GJalLDAi7Jvqxw
KbUSgRt+aDBXxQICuExZ1lLJQO3VNAX7mFZbf5fRbSKMqNtRV5s3kGwBxJwFS7TI
ytvt+uCkkoUvem1mN3snVBhZGssXDcaSpSxfhOJphZjI3CGcuX5LBIVkkaDDGFy+
uU2KQETxWnIGWnmzZwi5R8+m5m83YQ1PqV8cTCDp+c+ADOSuvmpCiLqReVRUKDk9
ZDMVh2lfYCAk5bT8AgTS2RLpLC0pMOO/itR3nUhFRo47frsks6lLqHExPSsjDo1e
Pm8DdUS+kPCLZTuYIBh5FKBX48vUxWsB6Y2or0xvvcJh93T9oiSjrqHOBcAyJo1V
2yt/ia0tISolH4IS2QR0SoECUr8Lkr/kSn93/lcnlRNVo3D89fXboni42HUssQ89
VR94hJLYvdnGJzPhEQJk810f9goc8QFTKphpXZOxVAVNJu9bvnfFcCusKK31HRak
PgX42WpqC4L6Mb+f+/gJMCSr/p+IHSdxaDJPdIGt+gmslcUAaJuLr2Ryie/u2S7H
h0n8VKNDUv/yQmMkOrf02xs/KbtXDO34sirUNna2vm0LV4Wf08mueXCWQvT5OmEO
3tk15IIgN4WcjBdycSIv6oT7PF7suP5YnwuD3+jEIRP86G/8dtMFHcnxkEAgBWUa
BfRmCIUae3pnEYizanidjmEvZCKN5Fvc+NB7RhwyUDAA2nY/YHxqrM8AhB+zFfp+
4K8NDojQJ+ujfxLq61aX1oH5HSfCg5r5u0RV4H4/L8XbCgXdqmQCRYJ5MJlI2ja6
K36j1LqAC9j/V2r8WgMVNwWtLMYsuWUMLoxmOtlRSmnqSfK/SNqESvO3khXTmJO/
QwBxxGFQBTYHsdDao3fq4TX0TLDCV9XbaWb75d39cy4jdX+7wXfBN76+UG0MxI3T
vttC6vVtkmlSxNSr/l9Ks7ZWMNrU42/4Pa5bJC2ydhI8N7KV0AvP/F+aMKYTznoR
F3Z6QOchX/7rPfW4yDR50OJPTziIQS+JqPIlyJys05PifrK/6e4UUvcphuteGH0N
zL/R4mhTISw2ZzwGpv+3iDPkAFgf1dBJl3wub6dleu0QxF1AssdzvOhGmD058je1
NJd9GLf2+QaZcOgb+Nj2fKj0JCI6seay+1xWs6g4xqg/s7SiSXIivTFC9C11vyNt
uBv7flahrIGrPvydxxBmhU4NK1GYA3fdjsyxCJzhm63MSufaDsSEfRBxO3ryVU8t
CnJfcb1ANIP+YR5ODGul5OnsKZSVYOxlqEub1P2mh4rDV5s55IogdhkGFW7IhKWZ
pX0Zb6eF6nZD/tvju8xpXBefuWXqZqZwpAYMCzmxvN9LwTKfX1D/yQmxizRg6cIh
op8aIcjfaSz/7hgrk/+F1DGWVdBFM3oQcGOl/UTEXn+i8zbNxdDoJqtOpCq7VaZt
dJAIQ/E11K4R/zP+VbTGws6PMMF+LRMpIwoiagGZzdk3xIqosyt15oII2VMfEJIM
fBkCjXPN5+0wZBTTegZ6i7RSjlltn0PC4Zncf5bm+caPS7py3zMD9X3ThvSCP3Kw
lgShrv1+8FYtnFBnSqB/NZr0yq77OZjtN9V/tHnP2mnkWlADc9Ff0nrAAsuzlGLr
t2tvv1dT+MsIAY6noNGLwihjbKf3nwYG+OGRZDv453Y4PAQZe5HGgg33UMT4OoJw
I/yRMtlJUC4KDZUMUtceSlX4to2PSBd081BS0GFa9I34WRltcDml41xakKmJA4Ja
emS0OAWvbO/Hs+/Z5di1vIlkK84Rr1b6hF9zOizF0nN54/S/3sLzO/fC4V+QfzNN
vCFB0sVahQstMdP0PMeaHueYWy5cO7VlyZxhMpuchQN3DPIayAnkQD0Fz9tTV57j
vwjVWRIyOA/fogP5qHuhGRP/glWRxN3L7myuta5eOCAGQVAc9lXWlheRR4EMoyyr
nDesRyg6kes/QPIAk0OWoY7np6SX4dbeaq89skhG37qJBWL/pHKwRCd6L1u/2f7T
9KPmA77XXHHSr5PZdXVdBrMc8RFTiXMfEfRnLoFSL4qh841xg8fvnpGHe/VpIim+
V/HUopT+ihzw9zTasH8Qmn+5/w5qLXIPU0PapBz+C9pYUN3LbtRrv4fndraqib/4
G9t2MH2QgjjgoT3WwPx0RME+mkWvy2KxMm1QVDqvvs2GtRyLjbqFf69U3FBvpsIA
ROeUfWlHognZzBx1RTR3SUZwpf3zslMfKp7gL2DPwKfW4AM7G5tvuk5UcxhsKprm
DX7yfLWZElEBStY4NSkLelu8LUT33w3VXFEbPmvyoasFJJntzLpsJAmSe+nmd5sc
V/IXYt32ne/VrJViU2hIlXAtP+WBr1P2+jsMhDFLk1X6PTkBK0LUwJO6tPBfzCFF
QT9M1CQDszJcWs53ZG7+R50q0E8kCHAxtpNrxXoNxc0LRjajd8TH7EAK/hY8/Vi7
tUFXaYbM8c6fVXQTLjzHn1vZA42COgk/Yc8CDeSKAroYZAE+bW4sDvvn2d9IO2vB
YT2NTLi3+n+uPuxqGvC6LSucLTBdE57RHquWmIPn0qNj0X3RCq4iclT8Z3ZYz/mZ
weLO42s/071UrWfZ/yQcSeNG+p7Q4fPuzmZeu6iZxJAvcBYe/3wcHqoUFFMmHxg0
9IxzhBDKuBAC4c/vBl4xD/qo1ZBKF1tlEgC02qkZ86ExEnhFcs/CEGOUP3RLoyAY
s6Rct5ZkdEiFVe65AeGTm8YTE5UEYKokYB+s7jBVSy8jOYzFR2kdcK0LLg91XGiw
eWbblKF3PumeZTSQU+/Ddf4JJf/AaoSOUtGRSK6tWbVPLAz1+wkzLqZFedxY5Qds
0Mtws+sKRZEkAEZIssuTsGEKtrG0rwUvjfa8o72gMOPe/BDxs8M+k8yPkESOgSOx
5RVUvSVGjvR1ctuSeAQDGG3hdSJSj3jCBJvVLngsRBAfnZzsutBv4GqO11IQ6z/e
EpBnoobVH3RI7ksjhQy614i1oPRGckL1jgN7kGnax0FeNkKXWcQfZc51zDA1yEfa
lag2M/LP18uBY7Y6kRoGJlZyUo3+V0Nx3EXMnh78uFHsi89QDIT+bfA5m66EWZ3V
kO3Nl+UJLbK858tm2Wj8lKpBpZK2THLnANQM4VRv1xjuw55SQgTnj9+S1tU2uteV
UGBoGEHFYDWh4UldUeCVPobe6NNM1mX95ampDR8cGI3CykkfxDkhwhsntj1UAMZu
7tUH/V+J8/NsLBDrv9+UuRU96UD1sAFDEj4tVLKaksV9jnGIQ9j+r+yz1qCUDeQS
Y1aw3g4MryGOQsFsP4TtSvZfZ9Lz6RO3ogrb70eOAEtxvhbCzA1VyMpDGPo2PCn9
BwPdAQ2Lz6Gfa9BrsyI/XKJMWcPzR7pwdmH5+9d7s9HIsb3wj7z+sF7eiJz/cmMj
IwqcL+b83u30Fx38UJmlImLAdjWvLgk3S7DDoGQtuaU6WvG+4M197SqH257s0F3j
UZXBC+Qh1xK/s+t2zE45DF1WUBsrkgjeN/roBRWtigW7QY+DZdtADl2ra5G4GwMn
kYewDPKUDEimHx6jD80wJWjbPcGncrOJD+vWcih8DsBEBEkyVIhcxw9ROOOJoCBi
f5I+C3majgFQQP1X92kCSoVcoGwcw844Hqlb2lL3YgPw4hGn3wAnZ4JmSHfyR4oD
CJBE/69xmQ+JV8oFFpnRTujneRKfPZcVQdz1iSvsuIdkolhZ+xaowvWwfP40cvbe
ZZ7J5SWVpXfRNh298k82S/Xw0ZGxE1C69m91awdpCKw/qMejSQQYQMdgQkJLTnuJ
CD7HVSxOBXfQUte5xfoBWYp9/4SwBMsXKu1JiLa1WDex1iuYaRlLmNSPYc7WHM82
tVfOH/OVCQQJqLozwFGBWQgGGMuWsaetxZ7msLhvr1JlS800kaQep/AWug+6cldm
7iBs+r8YxkEuYD7jZAkeW3jM0ceyoJQmQIL6i1ZsoxzOLhU/alyMAll++8hUdKuV
E6HE1PQnUv7qSKqqU9rVGtrIUH34LWonuz6RMRY0vXPCVqz/Dyu9YClRUfRVfXAB
+dKM98IxEMsrIGiF0yuc7/PDUC+KMWPV84QkF6hH8lFXMfraz1ye4/p9IZpmFWww
5+NAqCAONXDqRPx9HzLN0QQ3jm8mMNuq78zNQm7PhUUPI1RfGHmXhrgLYEOBuM9l
N22GSFcLKYHxUkiGz4muNaj0YPsbUCWr956KZikJjTwgLcCCQhkeRxkA1hVJBV0d
FX44SUa/2FnHbWE5294gDfipGhnSEEMeq3pf6wD/Q+XNjmCj2kl9h4hXssz/9iHV
pTECJSszHLF8cCNRMFBL0dvkjg0pJ/XRqpFVAgB6Aq0oDHS2B+B8FQ9n+rT9hijW
ootHCRw0NHJjHac65a7NTZM0yZHnp/djaTHTtDa1W5qdaLV9hvqVncbPnrcE9Gu2
YYdvAFrO8+Av6+fxei9VpJBMmdtzK6WV23kVYvxXAFSBnzGmhJ6w0Qx3sDqWHXLZ
42JC2RwSUYeWTaJJSiydPHWzXeB4nwgzpWEoAIHO/nS/q84a8abMZDODeLragj/4
kUPfnyHbAqqu1nfO+EYf0fF0gbjt59+WN0XMtU/zXOxFuoda9LuX2tv7rlHmW3v2
pnN8XGvuISAK/dIDhOE7lYZkUwO0qT9glNqPbuu9DNCAO2eC5Lt+9ImtH57pTMhx
cV0XT6n2eU4PY8gFGMD0TvTZ8ya0lvc+CcUdxtOs8p2RWCTuzbmDzuekGs8/dBmT
VopdkDWsymydyhI6pSc3BBkUAgD44S8EDCYZxizqlpz4uJuvRq6v433e4q9K4Hr5
80rd4Amyb1SJJ9+zmBX7VyluBM+da//Qfow3bMbiqxseuzcq2sr1whZa/0/OJ4XZ
YDNjtio2vRt10tg+O2GjZfO5/db0XDEDbkeUykTbMCK7AkWU3qWV5Fm8ubjNmWoK
V2Qro5ohQ5QnSQ3E6cjT5T2vt6vKF6vOACw7RuRqT3TeoNX/XXgHA6F+uWG5sblW
V8e2bPTzneoGI4cpuGP1j6lCQ7AwRPlFk7aRFtOg6V0/XkOiZ79D4c9yDHmRYFXx
dUAsalS1QMTDpv7H5uWLdUjAYwf3sGHe4+1b2eYNzx4lY+gGz4UG5UXYtB1MImHO
Y1xNSBTvFlcVbWCmUnHDFCzT8/oFg5J/kEX/is+eNUlMxZjQAsjUrPiGLd4U78It
wYr3ziCOLbpakeThTAaxF09ZfIpSKwRN3UHSfvSPB8QSycYNxTAMcRuNKyg4WxeZ
4W5z0w57ZWrmo0qK5SffO3ewg2Sc88njEw0xZVsqjIP/9wbIC7dFIMm0xxV/tDGb
wYQRBKaxkNlJbuS+tklWGPrXzdNzeZDIfVjBjLqXZ4Ycg2+8CmCMtpWGrN2nsDWT
jWH3TyLvU5LnGagVAFAle8FV2whtLtgcLdIQzZHvFwHnCA/D0xP01b0c+Qw2xLEO
Dwy6BHULi30PMEGx1UjgQ0b4FK1SNQfR4JOz3/qrI+qMw44Hmlr1wS5WomB68TD2
/yqnA7P+bh+s48yObFMlZ2yMUofkt02RuAfbv4SHtc6P+s6QxlmGiTGljYY+3K00
Kab9WAsxFWSqVGikDeFnQvwP6DscspWrZXhsQVu4NuNFN9C/pvOMMO5jo9+6+exm
HulKE5Y+OFmg6RBRFiLmH10kIO+orchI8Bv2M+pxa3Bh+JXRM+qQb/mg2qqpn0+C
p2U8ykc49dPCzzElwZiG6XNOmt3B2eKUSGkCwlF8UnOONcrul3gEJAlZ4ydV+fOU
axQrR6/QWM8gj+JWCNoVyy9se7Wm0VZHqPkltOgzujnxlMJY+9zQxUSJPMWb56vi
lwpwJ7T3uCTD0E1kIbMcqD377LFBsNORvGLGKAOsMeIhlBnEiAjqopXaACoeRl9+
zqflRp57s28ijIEnt1GBQwM9JeQPK3Otw/wWoIbJJEsfgxbtSc+fspTP9cJWCbNw
zyptGt0hFj/NdgQWY3K9ZZOc4E6K5aX4rIzzvR9QQOGpw7AWyTy9Oescxcs8de7U
Lx2bIsStPCt+fPyoCvMD2OpnqcYJ35hR3SYkuIBcn1MrkK/+FQseemh9/89O+gjE
Hf4xC866SeTT3IXBGJ1SsQVyTMz25d41rp1pPpvXk/tPlMbhssk44Obgbv8CpDnD
jm6jI3zXpACtj2Dh4HDBFiv+j50UCnWcl980R9os8tEIDUoBR/GeBeWweyHS5Y8m
+l4qEY7eT75iLLVY4d4Yx2faNXMHfqyh1l7dr4b/vCR67wwDqfJV4fP42sgcXPfj
yMVvRDcKSx3iSfJT1sDpXqJvmCEuuoolM1+7JMRytOrw5QZIl8PX2QykDWEiNTV/
oAb9qlMTwiKp1iPLqu49iQ5OY2llOekdqOZlZctmBxHRX74zFlacmI3NlwvhxfCd
Xh4bU2VPknU6wak7IVHdx/VVG8VA6SK5jbnrUaRdr5styK9maRoHoe2ckInYz8ar
1qIBhR43nPlcJMwhNcpyejb4ud3geORha7W5G7DUkc/dvM2JH0uAESmfpeNC09jX
Unm77zpVdatcKHm8PUg9sGQ74UGIT6CG7YwLFtGSKbPYAwgxyBVjC7PgYfmiE5/+
zBofnuXo9eQ3Dq1GlL/4uAN5RwmSgBY7FdgCpR6QZkVJ7kG+9/3om4Mi8q7ooOam
LKMeey5cXQGO8sofPOuWvH2/n5fpglaIvSFkxJ6gT6uv41nuciDgxN8PBWzB9XwU
4ui2ZXYTIru6RRzI8pC44XjRGNdiTmertFCC8sQw2Le+VAu1thMZpt7N6FH1f4t7
TrU/vJNI+qidOdfAuxDHU1LNqMxaGrnmayrCVGwcuTTSMyMmpKrm/1gDwZV2Pr2O
+zFe+GtDKzHoJ8JCPl6uQOLp46NwZR1s82b+ZLzkxCRybCTjXAw88VBjNltIuci5
fBsbvA/HYY+ou3Mml5D0RyJr5eyHXIJvTYOYrjN2jvbwl/ozPbmyADA0+KEOve99
y0b5nwkug9GAebXj6drGwJZw0K8h8Eh3gv/5hwrt79WSS6Z4xw50Vdi9cA/4n3sa
J3orkJBL2iUaPK0ktq9GFJaOtExiPbYoFAL9nXDJujj0YWL7O7ICcW7iR8vNozBA
c1riJ394Wfdii8NEngLn2SFqGBjvmCYzh/X9TIrJx6J4VzL3SVulOaVEcL1sXtUX
9nQDFlmBrVO8768sN44REfCGlfXkK9xDQ0AKOHCEqEGWJHkK1WkfTIcAcwBh0wRw
U/8Lpseh8gfzU3Y/UEhoSWd06T6i8eNZd75VwXly/dJMYTxofByWd9uYUziUQTOc
+67nGWtK665drpLZZw4vwXfXQG+cvR0dsTBqLSoVHgQbjSCbCZohtjL7DV0c4SPD
h40XH4tCD+dvVY+394/zFA/Qka3zJlVswXau6+cUfmXUFj/0BBuVShHPZe8PULJ9
sDO7QUs5XdOekLUcbJE0WkJxqfoisTIVo3P12ybiiaxT1g1UU3zz1wFLFzpT6H2J
egghszXs0bndmrm/fei6Y/pbuAaqfcCHhG+sduoAzoQL6xvhnJPKmTGmijj9b1zH
g2DcLhTtoBVWRp4Tqnzy7GqGAJQJ9QZEL51FMNcIJzAcUCY7A0b1KWv27xCZdHln
jmT6kbrtVakG8RXmltFGIipcwiOx6qBrhD82iL1k8ZXlff8P8D+VLtGGAgjsElMB
RJhueLQohTxc5QhteGFi4MPh1p3n/S55/M5mAvDJwxjgoLGDY2d2z0fp9rRL7CRx
xYADNBxy9JzMi2GtgMGRb6ZocVXi4fo5+meY7B5LAOOuPurmmknSzSX5hzzex4pR
bnrwxbWPyw3uYty1RZKou5PMuKaapEYlx66wJF3QqNX/aoMKDngGZrBpMfRi+inM
QYm3ymdolLPVvH+s0kSL2PnDmez+Pbmv+G1Ry+OX0wX2f2J4iWcgADUDKRwUWn53
t14PykO0ZFSihxSctyfjbfkWZAeNNMUd/xrWf+ImRZ9fZUtLQTBPAdaBx6nvLHmf
OfR88/bNjv0Yg/FpT6vcgU1qZ/tJkpbvSlzD6KHhHi1TCRDbnEjQ73SCgj1+70mk
qt+3iu0C5Kq/NLaMHYNcY2h/4X+q82rzr2y52DFSHz3x39uPRpumK15JKKoa9KgF
LSiQwkxNWo/405889HZNewjbI2QH8wqiGxokf54AiCvGnyu6aff4O6f6SIgXnS8/
VoFb5P8yart1oW0hQElkFcbm1OZClmuhZ080Vaczu3yZJ2rs4vF4jutkQPJdyvff
oiSekSeJyuyZ0/qWns2Jjq73Hz6KvDmNmE5WpiUvTkV591Nin2hb3dDk+S/8LSUz
OUCdpE1U4g8VLQANstU4ARjauhV8RuDcAUpQymrjRjcduKEhxoFM6Czkr+gysT2g
zvRmfR6NIAk9I26EdpGQkdiIx8KdehZt5DN0qfgjGY0BsL53TC9Grq6qnwC4zb4C
wCUzwBHvF1m3CdB4OW0qp3WY/jywoMuo1kSKMocrIEvN7kAAyNT3XyfbhUSF6Ndi
8p67ftlNQ6QiS715ft9oxAgJcpVVsYjDWrMS/x+EQjGAeA+FENDVrF+OQnUFux1g
XaZ6Y0LUuwMN6CkyHiKf0Yn79H1J6mQfcSeem8+MBJTNl0qaVpsORHGow2jhJSHb
G0Vs5i3+R2gq2lUKDIV9PQCWAr+pEXD2DCISvrwveXUYJnaPlwEgtbUzuw9C/idC
4Ir/ph2hhlrSoC3/KO3CxPydTvIxbYxCtzOM3PM7tEhAHiG1lNa/as9xdZ6e0+Ou
8+VMuvnTjkc40HtAN0B/wAfTSw4g+FqdPtZAFbS+IBgp6puOPsEWX1TjhitnrkGq
kFNVpPgXf+bCiqcfnfmQKg97szgINcsJ7jJYpvvEiuuWUC9YBVV13vt361r+Cz2r
NLMmtZ73v/kJ8mxbCn3eJe2tP/KKh/83cShmXXixtUa3VCm5NEGrAjLkxHHHv7Rl
0AlJa1UK6/xF9/3hk34hkpLT39WvYkNF8ex8WV0PUBoZAUBBRrLtYXYlgfj+moiJ
KnoYPqVO6P/NHdTG8fsh7SsApBR4gGrDLg9n/EJIieZ519We5jYwMkRuszuvwKzh
y2YEAUsyh3u42QLxBS2gLk1G8UALvFR/b5oT9LTIKW3go5Jk8kgCIMXHhIcOrd0u
nChARPAgdBVHnso84MCLJd1SrAu/N84M8Z2pMpQ9QRJCBmHxwDSJsDvZulRT6eHi
ViufKOxDIc2MjjbK24nfWn6G17PveiBFDJamGcB865nfHOM0qIxFYWFVGKgWY9rI
9/1pcte9ipDrINXKkzyndEHD7CHf3bN3BDvVqyMfxfUmmqtTWF0XSfr6oC55q/oK
J7oytfO8TvlNW7D2QPvYpbdqwaBXsqLkEZS3VKPb3BnaClAWIPswJPp0mam0T2kl
joyi3LwloS3UdA3TiPxa55epE9DpVSjjANTDZHK+E/Ky1+fCJ9fUoJUT6wLteO5l
Qcu/6Wp8uweL0jJWonHvBWTbXtBS8RAH35kBpFxZptbKLJ4UNho8u6hrT66ogIlm
BnKceaAuU4PoCpP/31zooDGmTg7a7N0aGFh2SbWIOcxLjJC+Z9NT7j5sXbTF6lvi
7bl+OAVHePvwde7F+PmC5DwoBZSx0CbNrmyC2/Hinyx5fuCeK8qOaV5ma/mNHJzc
6GiMtAHIXsHHTakXTUkPAjEAzdI/AIWTij+b1FOYuqeq3TMj8J8MK3qsFVsMAz8p
/GcB1nLqGcjwmuuzJq2LYLQqOgDfy2h1Xpa6JzhPPU3doPiII3ezOMdBFn/ybTFS
ivkr29SniBXVb15UiOTewqFciPDYwAg4RrABWPZYYtB6CQ+Vbz+FsTtnMu+A1EAR
KjHbQ6hRDj86YTASfqR2I/KC+0/XWmzSt0cQg70cnZbMPu+5XyKR0cYmp8Zlqw7U
XTv1Y4RN2ERyTaxw0RUxck+lU+DugID6s6Igzs3gBJeL2zHt0qHAyHcOwjZQGZhj
VEp7o3k2Ysw2g5N9iQoYfKVrSSSERypHwAEdtZBwlN0ActeGizddl40jMQ8Uty5g
u/gZLkIenxBQV4HIK4Q0u5lyqusS/Uu38lLc3FS//dG40lEOlvFtZEtgB75zXUvP
fs1Z5U+57y/oW8txLdCoa78UuHxCDHOjdh3+zOzm5JtZ6W+HtAdep3zR4sAx3aM6
K407X9NR5LeSkupycZG21mLHz70o/SpRLzfxnzbwBsF6TnqbuY4zHbXP63Xa3iSQ
c94t+8ZYRTuOA6eURQuF8xShGiRdBs7nQCkQRpEOiifAxQaUKXh1DOnPTRvFR3+n
YnzWsb5UxYeJV0RPIY7s8TSC43VUz147jAU00Ba3WSEhlruxguwWARDCNq7CDM79
Ks9mm6ZfqIcTBb4gAmrdWbMyMQeBsKHnJH0C0G4zgdALksWnYQiyC7T2K/yrT3f9
TVEq97SHsAvmWZ0eA/lytFB6IuVWlbPEJHQjlpOUP82rW+n59UYtpreV3oOYXhUS
MFWeXGOz5q6pxL+ZnydN1Sh8y7ShoYGm0GUN0ywZ33I8ZgJZVL1H3r2iZinxPmPz
PkKRG3uduiM46/7SEBsIT+7XSsz2EcQkWOJ9snMSMvKNxdLz+gNCcA5AXCJ5+5Cz
wfB6f4Ylfe86HN4Gmb/7LkJZhAP9GgggP/935Pym6SBfvCb2DC5HxVGEbTReN8ne
J8NLUsjwTpxVk0j4CAl/6VcoAOD0Cyqoe7oEHIvCJsg+REqGCTcEjXux0Ttd1np5
Fh0JdojhFi0CzfXY8g4SjHEKV6KfQbtVv0GQXSWz065gS3f9/OgDNzmAlmV9JSam
mdLzmkEbsov5xFSmul3Q201GR4/+i00Za+05/9DoBq4IWYCmMgCACufWXGkezWpV
lWqD17JbTmrsMkjP/HCEUkEIacSDqISEhv+2RKWlkGDCuLdGsWZNPv8GqNpHWOYR
PrKibfRiF/vBHDsaDLShjvUr8KuSHAZZrlobdrOKOlnqFC1dq8WV9PwmBQlWJPjA
6gvmMcUQ9gYXsReTcU1UQSdxNL7j220yBRKS4527xNf6lo2tvGxX5KmOAS/BCgvA
Qo6X727e9q9hwa8SnP/nw78kvGaYz0tmJa+e8dg2lRl9hbWd4Nzd0kZhzXbCR2qV
I5SKSXIQ6Rv92fd/n0hFlLiepraPvFmEDwfCo//0E5v44dndQziXe96su/RCkfOq
ytm/Vq7e7unLV/YzfcxsPxNbZWmEuQOjEJvjypzahe09XM47947WwcLHu91yL8Eg
BPV2Jm5bDMpq/XBS9XdPKrex6SpJEJZoEK5JAqndyRF1zUmW8kez+o5CSA03aUgZ
fi90F3xRwylC44/ULDntpTfJRA3gIbTzcrz+6jxMHH9vmW0HGK7CrkZMuclINyA3
aZ9f8fA2p3iFu20jKeWkyOKfkRP30hNdrcZbGjLznIt5aFmHz/BEOcOlxc6JU5/N
SV4h7xA6NwjZw8mEc11hEVJymOqlpZLH6SinwSjlo3oI6vDASd/o2cfNHQX4PmT7
Ul0TrlngF0Qa0PTeWCYK1xTaz/fikhJRCbzCVQc6ITIa9Q3CaCBeJGcM/tAFbI4Z
V8ivcl1dV5jGfb2WDcAW8PDtumtw71e1tOthj92HYYdbSCX/k3h2W2JDkSNqdqEg
K4+4jZ0DlJaO3I9oMS1sXkgTca+zf2P57M2t/hsrAb4Oa24SZZeWjrDC73CvfkOu
iJ892at5vmW3Xp5DeTPiLWrQqhjQWRGH90y4g4lSHJB8HCtdJQRLiN/EJrPD8XDE
/JGUCUql2G+fXr9CewAQBUHYFFACtu6C1ugKVAtwG7VPYf4hdAaUyDJufUsZTu5t
IQke3iet6N657pmv3u8St1uI1AsMp7ycvJYOTKQ1vfBVxbILf30yruImaK7RN4Sd
sMQZ3cG5u5KgZqELX71VKE77VN6DKQKwhEHMWOYKLsvYgPyJvtN3ql79IL0k8b6l
tAOHWCkXELhQnbB7GoEhC+Hstuww1mQZ/5YpbLOer0MSar2YUcPHleuOVPjk8FaN
crymGpi3Jz6cO5DhP6UiquURz5dQdEm9hGnZ5ttXKEsQood8G4D9ESeiacUDKlNX
Cr7rN3EsKhEN3F+opNp7iIgQx3pmgHyTCqiCO9gBnYiI/nxgirlG6v6w3lHdl29m
dzBbjKZm2h+Sz+K4Lxf8zRDMB4zbzTc7A5kCFRZCWvkZHlcA3G962K3rfw3Dj+iv
jcLtCZsuaZKUiWZSqjIQEydkhuSfikS/s5mrcBp8B4fUHmnE+FnLmHgYArHhkO1T
AeiS/5QEid5X/WJ2spI32a9E2MBB631q6ecBdHJ0FDAC/EFt0QLXvkJWYRmomMYV
6plUgQ5FZdgYcuqfFl1pQkxvCKZslGyaQtV7NbsDFBRBR4+Sihqo4uLIUxXf+pl/
EtP3sNgQ3ViodJ/oqfC5ZXu2PFlJnHuEAHCzRbiX3jCgf/S3Si9F+0+O/L5c2nYA
n/rZ1hESp+aWQCTfWjPQ2THF+0USNWZ+tNWMvDx6ZkvggGdbTtVjei1glijTyVY2
QxigZ5YfaUykAt6gQ5AFRLQamgbqbGEIzQmkjwJe+Ws6JJo5w6T22YY8nC26qOuJ
7U5ss3vDAu/aw0VfCDtI9MrPIr/t1Fc5PdDgLGHfuXPGRSOTrzF7usyl2wXXgSx1
Up9FR8jlleqOIRZTr4gP3Ji4vPxvZXsBDNwBMzW14eMw9Kkpvy26cdICQZDxFzcj
QQM8VFB8IC2tAfCypBILB9Ctw7XKaT0jm4PJ+FPErrcqQU1Ua6/0VsQ2oIk/D/nW
G0ci9UZEmfhOOjWmRubzPpC1qfrvSQrb1GvaddbEZ26W8veNh2+9IHNo8Mjbkbc9
7mfb+61/j5sV+xRI3h6tzdIaz1m3RfX7hAGNLYi/zo/csqdNywDOkrRAz5C5UC99
xSTFTqtXWcm44KyEOxfOagLxhjLYZv+go4qMp034qvO8Z+THIjk7R6Cs3W9GESIb
753PuhZO8/c75vC/Z3jcook2pmaMtji1VsG3g4OOeDm7/pRH5wDAMPD7laJNfZ0u
vz5cA1OKgPSoumlodkI0YDqJWGHmXdt/RKIs2Hwufhw/2/kHhQrBBpv4mm9dXq5a
Pax43S0KZxQraZmb/UaRFlz0G7Rebj9o6/YiD3WgOjV5jP1CKJMkuPknKiPb7BDL
b6+pRkbXFBCtuXgV/cXbF2E0UbwgYa1N5wy2gAIgIs5vNnM/hyERt3z9lNcBqeHA
31gVtsKqKO+lrPX3B7x/HnWDjFCsNKg3JaFTZ/SOsR/iewXpNig1eTsTh//9i37d
+68sgP8Kgm+JqHQgSesoBpYX+ukgkr5k54zVOLqeHVgJZFUMuqBVuUSeXh89oy1R
iyKAk8Y5/6pNJhEK258cpX19K6H9TRtIB5BzgFnDn6nwPMGKYgdg2tWyVMKZkRUk
rQ/MfOfHTW46+uZVyCQk8cEaCsyvVIsJD7c/nNVO2xdTmLphfJiNelfvpi+A/ko8
7Bwhgnf/yjjlRB2LRA+kEj0UBEL6L3QmXheTaER5HXtMafmw/PbQf6U+cry4FeCr
Jhc3Ebp6cDRlTw7nGIClnGvu9tmme/Vq3VbElvgEueQZpdIdNQFMEickHthTKCHg
/rmH74olLFCtk8uEmRiVuX8Rvvo4jy18dhAxEuhzS0ncgAXEXE+4K6ndoPzKgVQ0
x02GGvk0/SM1ylpaLJn/ERtdok8E48iHM2i3mOVeGhAIpPG7uvz62wCR1FxHCHIb
m8kgbPinrdCyxOc7cfrEumcFwJuPaDMXmoezErB2q7eOPEBGFXAwITJx99zhd3+f
kHEQrMo8Q4+oFzIF/3mrBkm13vRXoZ7yzHhhQbCLFsM/ZNetKSZNbM7SPuqVwu3/
sovh/ANR/ZPDipOzPH0vXr6yrRPQYFhNNu+h7YSxTyojnxmYTjHnqPEpDD+ivLRS
b5Wfqo4kwJcN8l17NqeT5CGrdgGRUCCf7kzSJKJcsxSG7SSZ2GdS31HT1pvc0YiU
QQNnUnCtzLOnE3K6TXzLgP2ta8wHDH10ksQgZReRmhp/PYCm9XgFSJIs9ZizWg/b
52yomZC78XQBhOzbjQ+0pmzefvQl9xZNgSBD05p9bUvi+2tt4+vmWoCT+Kw/i5bx
gs61TOmIEs8HC1xYIDr+IBY0LHaQq1CFIbjGgfSiJvB24VzjIdxZpQbu5pq1b7A6
c//LPAWWdTFCi6Vjze3QPHmB6v4bgCYrQ9yoehiYrk5aixmjYC3OJ4q5PFk1EZ/u
Pu49Q0WCRUkuiduA0Sjrx94AkYjBz8Miq+VBsO7w3S0UwfXaqRs4VHcHXWavgDlb
xdn8mEoP/aphv48Zu7owld/OBml3HBBQdoWfSftDGRLdAh1nzJP1pFXZv1O/CG5S
1yvrLPLgTJz6TSC6HMZcVDAEKqfY6aE2Pns1WlCnAHM0P3DmaOeqbVZdartfvzkS
Gl5zYtmic2bWfL8WxKs5LwAxk8U3ElQqmkxtfqhmTS5o/nis9oqUochAzeeuVg2/
D+reLTmufLSR82LjIdzQ1D5+h/w5B1EPkrGmD3pXL/36dejjNuahmpeH6ySaxQ0a
HrpvMqfEzfitRxFjp5Xh25TvM4S6oTuNCqVvlgQz3yf8UtatE1TvxsTH2CEQuVSO
I84DIGZYQvyAm0Gr8i5eXOq7X8H8yHd1qSjUU5908VOAtL4PksdHYBcMfhBPK5Iw
YM766sgIIdQJDPq0SFixoTVNW+T5FJEyWWB2RGLAHiU3NHw+czWHk0AOQAZsotL/
xc6EAtzLqtf79YCgxGLX+4Re1d9nDlYK7VagRVCuLFFiS9Ap/e2l3PiAcJldJvmZ
zOlY4GQj8YQL9kmRigC5FA4U1UygNFKwQrDqhE2DwMhauz4K3kt1fLaaKu93f3eT
+ZcD6kgnyXDERX8Db50HH02GCpThp7roS6xZFymlESkWB4j07v6jvG8W8o1aGVfd
dQXZXTzUnz4LAoUTR3sRp4H9qpOWnDEQ84EVm5NvAfgs6orKJ1VN/+qsK4wNHBYV
w7pvB8/v8JVtylkuuxDB5teqZKZjANIaYfNHszlcz6sjS9WRtGJpLH2OsXlbWb4N
pDKw1ZuV3qQSxxwxOoBVwmXwueul8SENvvmHAxS5jqmE+09me4z4wPrMmKfq1UZL
vuzsMhxVl5blkOAe8+Rt576wUAJMc+3ztLi7sbCJYZuvc38a30uPrSr/JkPVkgXu
RYzJLEuscE9I8F3lWj1I9al0ds/BU4RJt/5M0/Yg0GpBnM5xXjMOsRKIKqRkyXSD
JNaoU2ll5xrTSHqmHD4fcsjXKwBm1m/0kHJc93yvdii54y6gbinf6O2Zd+pEiw87
Z9YFHJJWsp6yv+rYGKYD49tsvvbfQQ8FpJu76tIe9Esl+a8AjjKuxgXJUTdRYFpZ
h5mts/j/UYioxy7gVbP1MnkWozelkOlgF4epJyEnPjaWHM//E47lI2wNX5LY1knB
1kCKaDgd+/Eovxc9qtVCl4wdnJW4vYqJm0wZDzCAI/yxMMDyFnZT3eTeFXrLgbS/
XP8f/jTth1YZwj0uqinI4LMJg8RPT+2/8rWSZj69r+QGfTkwUPyfV++OxAxlEZTJ
+MJBk+UB+wmrQfdIJO8wQkjxZ9hB84ou5PpyQQA/KptYnWhSZdWJksUvpMnBCDka
ziAR1l2MdNqkCAkQXRKhwJLRq2mHpBLXZxNa+ArDJfe/58wrgTmShcXAFzCB6Wyv
6fQSzhu6beeSYI3iNB7+cUr9FhEYw65QC+qiAVqHCBWOKzOkAmz06LQGxlg0YFa0
S/MnPeqF2wKRKa5mMJs1GnUoKDgFjmxkwIQe6EUGnDxfBjUa61wqjZUQ+NMKPsmD
zwIi+CRfrJYuqlyoSU1KpqUz4PmJqNbM4GJbXdXMHkwZMuN0nFc9Cpf7+MNQ3BC7
jv+wwayKiuVT11I1On4nWQCg+74lON8AxC9VXi/liQQY5t1Xl7XeixkCv9xhHQ0N
MuLnhpvDH7GumGns/hJK2avVTa9WyvkSjOwkQv6jp8hVqwUPaJ8FMR6R1XMj2mbR
xWjkQOa/NeQNpQt+KWuubJE1NgLr7/xaqo6MapoExOHpQ33oDWhETiyvoMeVaxEP
aw+msXBe0/QQ9JC+mybIfB3oGiHx+9yEK3MHo/QPrRwGZFZrtfAE9SBx4zxqvUWc
zv/d+1tVk5tR98aMpjPQZ380LTctCJ/+scgUuRW/iEJfS+l4ZSOG2jIgs/wBXy1v
iGcbvt55qo9Sdmzu6HmH9Maz4UI8qm1u/BScIjS/4i5pJfyOm8zkj8gfgf8Jyxlm
8v31v5LKBVkJ7L6UL+dIAxDCtfdrpQeVFqp5zPWRpIXpC6vWhBlJ0bOfVPwLYS1y
iYjBilBxPCztru/AdmFYPHkSUpcBYuV+zvdHvT+iSvmReLtAyHqCxB6LVhEWpP3s
gXTkXfst9aKJmD+1MFEuLD1EjV1Geu3NR7OxfJd5lGg8kwKyLI/Tyh4snc7SbaZ/
sa1i6UEcVWXa9alQ1L3yOWiM/VCLKmKmdbFNVy/MgN/+rtb8cLPDdhiIB+DdKICg
LIHp+WqQD+vIyayBYP8rv3gAPQymS/XFjHx+Ul6YgPOqSS6MC5ob0ftnh/HYIQ+r
X+2O3UPBgtdcGCYN9rIQs253yOFOXVzAOz0zBSsZPSTLSrL382XFN4+9cGmEK6c6
0OPn4CyuytBQ/rjif4ONjd0aZoc9o2N7kqYOfdJapA7+HR6D2Qoa1LifJuXaRMCL
O6SGACWMfhTtqFwEmuhKPNt1Y3mUpWzYOCqr5H3lnjhDKiVOvJrLBGUaExQJ1NPO
vBVtBDAuvXAbQC9dT1NVz31YflpOmONDIyq1vDmGPOjZRrV0lE0SwKrCpYQUHlzR
B1SwkFJJSxyStMOS0BZZ77Fz6FZg0zaAO61AbQXm28it9ZPwpb5gwK2uqe5FJeLV
yCHIrBoMRjvcTWTLALgCl0T98e1KHkFvUuA+AiLx7fNVp1QGbuF2CFBZHOyJ2dmt
5eQ8/kopiI2DwL3q05LY9H1gpICBA1MWxeIBFgWaUOzG7xd8loze5XHCwOSDAVya
LdWVWFulcZ4mMd9AHw1TfA0HN2tgrCFhS+1JyEF6hgoWMhBJtk+v1unXIHOa+plo
pyNdw3d9cGCpFO567aN2Ejy3D3qvQHyWAxKti3d6dbgLgWOhaF7O7zuQbyIJZjII
7+WeznCvEe3Zbvs0eQnaKHiE9BMI8ixEke60lK9ocXKUz24E+mQWHvoPO3hw4ft7
MugUvuYDbaSZ9CQgKqMXbJee9wQq+TEYjUvDRgd376P0O/RfTw1wvAn9PPaI2dDd
LH4dwmMqwowwtqTcMVRk7Tk5Xeqnks6KL3LVDg31k6OBtWpyH8CWFkwRiO5hbLGv
EmtZWfvtVWi4mF71BIzMOJVAdwYR1IQJYl4crmmDh/+8oDrUPdnSle7EN246xoF4
svC7oA446BcthvuYJ9BGKtK3XD3ZWPEtqDG6yHdylklZ5TFMqQqhJ30v9PAHAzHT
Lt3/iBsZ9iBBdeuBBFslZQphbtXChvpMeNcI2daKq7Dnm8FqQ5QmWemsHVrnwRIi
UX2A7armi7wj4ffBuXCJNYSWhulVKe0QvhLMF4b/lckpU12HDZzf2fgNb75LP4Z7
tQGZYj1A+gZ2Rug4BI84p9bjTqQRu+YkMgSXCPtLiDtoVBDbhT4tXREN0nawkgwH
24444tMQQbLMPB9So+4XWC4p2bn6O5mq8lQIVVOopl/ciKcvEr/2FCnztBS+X5YG
O2ybfvRrCfD2W496tNBZb+CaRmQ0zZn2y87wGofhheNXT3MI16byicxGUK37i5hI
XNU4MwrUfb1n9qIDv9bMIivh3Sf0ObYcqrYVzryGLq5G2FUwNgkjwhRfVMX00QUS
y+PFXf3mCdfG2pXCJFSAJurjWwcM65we1+0kBvBdYrdSqkl1rUIJdkgu+3viESNY
fcCcO0B9IlaMCO3IjCjGsBpaBQCFy4LMmJUOHOdcz2Jxzh9YIDDEVP7NPvZAX1Jq
YrDtT8CaHFuRUJZ+1Zcbwt3AZUjJlQg51ahAZkAxNCOQrRxzJ+saev2UmyO3WTVh
FSAImv0u9DSJasKxGJPikSU/fRE9DfWxS56Kju/ae4WvurCCKh0WJVQmuPhTnbzx
jhNjDSA6mtsSmme7gdlS/TCX7sU6IMFYyoQsD035uZyo791xrOn5SPMUdcwFAqvZ
6JSxk+YmYb8hpgCSscUDznRWZn337/pUC/BkrAyw3PiwkHjiE43KddjVWIpKiVMb
lWmPFBv8O7FlEeQdno8f0DjVy8/w0w3mXWPv7gYAmuZcODEgZsLALMLtmcVCKykR
Nac+JdAzjxX+XERIgrxLArvlqT6HjrH1a+h4SMzu+j7rGKEjQYaPFsKwxgnbNrHw
mp9REoF3X8OUPjWhJXRVm5hz76rXM1LfllBLldZ2YwYI8iDcBulnI+GjHOOq+At/
N0rOORhYq2z3bOHPjgpOA1fqYItCBFvunVMrGS3NQ9hfI9gkcOA/kOVJNgvQBk0j
s2eCz40fCLlzauqa/SACtk4IAknLbv/JW99Lgr2PmHKQ7OvfXfDnW8b5dOhvq9Df
s+TUFnsWvjfrCy/HxbE7RgThwFRe9cIxTyslI9oxqEtsIOlLfqGO7ZE5Ptxr8TP4
xnDmZTK8crCqGQr1bPNjtthxUXcuAIN1tyNctzXoae/RW0hWR5zO/mot8AQWeNe9
d52IrfY1oCNHliSDfHbKgwKDjgCROraqE0pqC/xedUvyZ7HTizFkbgrs68bqOcOA
mqmXllX6q/A7AYWOVYMTdVzDWjUTQ1Fp9BKZ1k8vZFdToQNExHubvpWgJS/qiuC+
iw6G8EzwGa7msxwiC7mYbBD6JDcXK5FC3AGsxKpj4Pl/z6OKzKA9g5ihCVFbeSHR
rPll+hSZmR+4LRvWnT6KOP1LIRWJsVRmjS9Z351EcG6KBoES3dqPax0zhj6R+6c4
nAFSfibvW4Cuw7vVCl1Q7VqdlAetHBN9uQ30RaULbKuXddZ1H8NXs+dEXMtV0OeE
2u7Ttq3BI47cdb7gJaSZB2YB2AnULFXCUCEFVUwRrFfmwBB7y+iyekMu5SCX3hKt
G70JsgVLMs7kH31gMgWNedDSaC+x7LIznZdysb2zj/FS6jyXwx6dpWybTjvmhXdc
5WHEhvelYATX/eZEa22bnF81I3S1G3QU1H7Y1NeXmBt9RNdmeM/wj3DZ6Q3RB0x1
B4S9EJD5vc538HYfBBdUZYiI4O48q64rvur9dtAShGcDU6nX+neq2i3+q4YQaeKL
IcCcQ4InXTv38BTm1njZFkyBfj57oZCaUOECmNd/+YK0JMW9BWXOzMiIMul5SkHl
U/rIEG+IS8250PcBx70Zt33HtIe+YQ0fe/odLuMbY7D2ZdytQpFKhX9d/3xHHAEB
xZBJbE9XkFrfpbaX/eNRhdpDhw0sMPC1mfYhO7FabNCJ8wQit5lbVxePi5FgTvK2
zNnmQugY76MKS5Voskhujt8Vv6eny1ws6R/1KsmF6KxxFSf/9geWwtaQa8afnXLQ
GypKd94qndNT2IlziRWUucCTmiC2MPfZo62uIZPkijVf7/Si65HZYUWRNa2g3UG+
Y9veMecf1oGonRomuEQae8A27KbzImsVX83B3zIMXa1VmG3ZcQVxB8z2mIxiO9oW
l1i9wNNJL62uXcsHQVHjCRnLIRwqZ1++1mItTKp26prLKUmvGLhTC06XGCWytPRF
XcRI5Qob0ElhG3dS33I5aoOW9bLSA7JQQ2XwH8hiwuf7P3z9Z/UCfnlsZpOo2qTI
W2diR5AtfG93RIyLXwpl5+Y46hJTWLfQ90G0OCBGgOGkqavm3KecSCLbaIIx3S+E
WhjB6KLYMqPM14m4jD4mbqPoprMqhpN6+ui1ErXt53j2xPn8nDCCWUScPCGsvYRH
dNp/sZvzt2x02r5jpj4IuBAVAYVwWk1o56BSk6kLSt62kOl7LNTNHC65sP3bmDi/
BinLShb7UtJPahyLi4WqzWyhM9ogtQzCB0btiQieAO4HiT79fnesy8589EQmGN1z
76oArARU/XTWBpQZ92wYAGz3mbbkmpZXg8fv/WR6QmpRlsLw2SGe3OjrKsR2eew0
lnyiYmzq3/v0oEwtTS2yYRVMJ5HneWFIBUAtECWqki1bUzwGUcMbhcrly/4UIj0y
11zxLwjeVa2lYfJq9ISfRZvp0fTGcU8NzJikE8JWldZSCwm54mxuOGY8OKXIHubY
1WTS9wWoOA+YvjgmCxvDw04pi6sj5I7OpE+lsxqnxSzhYxGosjkWCWpPcbTjxuuH
WcC5L9ePuRxnlAc8YofsPHsPSmrTo5U7tPaQZAwtijMhXwCnGEoPYQ7HfT8WxMZ7
/guZTjNtEXGtuTTBBQ1ATZrIgAu9ei5BBlYKimzZjLMfqXhlWpEWQN2KX2Fuho4l
IBn24/V7YD0LOo6E6ZzQ7Lsje7trX2NaHP7+YNzHmoooPSH2YrgecOPmBFDnELBN
kS2l7JuW2QVE0A+veXzheUYyuybHSDJCTfdp024UtZkbZBm6VEGbBzf/VdGOxRim
Wg0xSCITrwhOQ44E+p9JaIUsSYp7/wXYClpi9cgJuCNA98UFMuWR056gJRCII9ZZ
IqMu7Mqqh0GO+5TwKdmDHE7TOSVKdfPkN43+4jDIsxuaF2aa7KWMQWO8nXTv8L3r
HBJ9w983LIe59zmD8UkgzpwH5KQ7VZBjUSqJLSUAEwnAthcy9m1gJwy5v2kZRIrH
cUoYG1RIBoTiOhU/kdld/EVmeCerDAUx3LaQCk9JuugpoMU2wtjZKYpdwLH89zyx
NnuYbmVDEwPnGDWUnoE0TyZszOl9x3xtMjsR62iUssOfuDm687bUT152JPF1dqGW
mQg8J6QNwOqsRJ9JKDPvpajkSEMmPcGjkGlPa3hHMQPbNJNoo/EnxyRB21in075n
nqT2JpYrjHNZv4sEOxilkY2Oqebi8Fsx4J2ZPA6MXCBCL2Ebhl6Me8G73b3yr6CT
mq8HYU4FVcJ23abXEZea6A2m38ehQpNaqImRcPfI5LYtAJIwuqg/CLJgdxYl+zFS
ncjdHpGtXwQLuW5fBi8sG6YdNilfrG0BYyYtzjEuM6TJOiRsT0zwEiFyRwML5rh3
Qc+yhpddn2UK2Zo1MBeNXcmGh+Dwm2tJogmngKgSoSPk1gqyN7+OTI5vlgQliHaR
W4zjFTnB07d4pXpMWktIXHfWI1hTHDIc+DALciInbngq8xLSz3Hp6RZw3x0sGxWt
+uECFtTY1UKrlc9625diEk3yUg5GAkoUBJOh+qw1fPy4wK8bjy/sMsdcHzrnOwNa
lWZ2Y2NbzSY/CN2wZBzcMOB1AcKptutd0kyYdMcO/q0YXx9KRVOifJHRhYiPYRIT
dqLMEJnovb0v/lVdu5umzPKzuQ/5/cHdvKDpbbpOQRClyTkFNLRNQ6RoaTCb94Y+
UYB3Mtmy2J38ZGxOY19TNUe+RaBxXHJfJmDiyA+EtbAn+l48/7QHawUPRbEUL6Jo
NaS9S3lhNlMd0z2d2dscU7tF5+lSH6RKKyQHWu1pmtuaj5YZU/pTBzGFPv7+YNVP
WVuzyfykJn86HLayamoliPWhnNXYx9B/n/vp3y0MBOD5UEl5OTmFPZgF6SX2rvgr
fqZzmuEDEihGj9/XNEcTPslpFooAJAiG0C2LLACOrylz9iKmCJHDhVcN/hnF2pbQ
K7XtH5R4ChdxFIHnRSjE3lG5bIKQ6XamVai4J0zjdwuN5qXCmWf/7t6lrPViQqY0
yTJCmYd0nq78xKP1/YjXNPo11t1KBaiFCbUDouw2broXhw4tm6ktL0hApEyIViXX
4dmVgJBRUWZowicclNStAbSFN1dU0LeYBLk/YOdLRC+w4igmkrwJRgg2qdKwHpGp
lYs/U7KPbihuownt4nASRZ8jzNWhdA/pKV7YS3E1nh4/nyhSk/D38FGkpTkjOP74
B0ayIc95Px/TsIMbAH3oltknh/C64gWp8KO9q4HfB+H4iXxpyUk/rVDaMZGGpcGF
MnMGhRrMXjnnabPwKgTetmG6WYY6xp7pKvePQ/B9Kl7cpCUfpaEG3jG4075IzL8J
cC8xWtmYd5+0CFiQZ/yUbzR1bHscKIjZW88BUmkBq1tEdoyRDfED6YDBzUi4nBhK
Y/FhXokm+Q30sOssX4vr73BpKqM57zzmiyfEfjn/foa5mDyXyZeYDl4QYCtNQy1T
tjZn5g5q0cl3yPUy/frCDUiXXsNbibTXkcWaPEhnvbRdvdQaY4lMIi+fktYTEurJ
8E7F9S82cLYGUKhBmA6Bgyw76tjeAyeScijOHZj6H9I228i7TUcDZ199UrTUb0nP
tQpgxV2kYqu1WU4OpwCkPZrs95bm0nke4moA/gwMPTnpCyInbagOw5CKF0LQSIuP
ho1vkhOjqPa+Z7sDYcwiMieR4lgBDPHSQf/jaDvM1KJe2EqocxmEH7eGWvHB5UCQ
BmXUkucnfGfPRq0GNmLlEOtIMvx187FanaQG/TU4BPUFedlFvPL/FwxgBl94UwX+
0vvAbX+lMhvTlLHgmqHCZu2Cq3oNey4v2RVGaNV/EyQbRZcSx6HNLD98JWAik2HN
11Sk2YNoGupHntXGl0ASpgpfjkrVOb75/fgPoy2Qu2O1op0/xR/qZzDDwkQJtoLl
qfjDXGw890qyOimQzo2styNosukym7BLOL2YpnqvELvCdlRBudLHHib0ipDByOhq
HIv6QaI7ZEFnr8sr/jEFHuYCtHNrEJ/GJiSGavj6a3LsEzYCBraQol1oeKj/k3Hx
h/5U3c+lqV2oSUL64/DVvKwWrHUGLYZY2UV1Tm6xKfhaI14sn9Rm4z1MWMQo8SFq
IESaKzw+lZac64SjFvv39xJndJK163ZWRHwNY2ssHHwvpX166ugn9QqJ7jcXLYDx
/UrFp0qnP8NgBAGW+Uhilm+8utMN0vTDI8uARqz6ZJBmtZJ3dWFiSw93sC52G+pl
dBeKJrYPDcx7teUoSVpDl7lMTUjVRahFlRJlRzqaLWOGZd1FAenj9fdCbz9ZZaWC
XXMpwJ6JacWfYlJXQQJtzbwSKd4EGzOyA+Nv86bBfvXX4ZOYRNiYd0iA0cR2GdDH
p4LvCSmi9jpeC7zOIyTxUYIIfJTY6DKe6PZA6CCpK0e9/hnOa0R0K0oA1tnlmLVk
BvwmPnI7aN00wXepo0kP04GtsIz7k+04jQhsNgY5pfMCkjI/79ADpc0IhZ4YQ/QS
AjKHbNO9VxoJfOftoE+uLrlLKqf93q3V+xwgIr1azKnBcfY4TzFLDvYyzsekS85F
pVDMOi4/QXFxP37/nCsdC9g8hktZD6C6ufRztFY6s/hKd8EslGmckxvIgjFRJC7p
hQzEbr8mkG93ibxLgj4If/vKyR2jQkDEohs4rbWAkMnkmMi7pcInjhGjXyy+/NHM
EKaLZu4xZKYjqly5wIX0f+1shiMRV4W4RcsuDT0470WbdoUoXZJ5V4IAto3/yLdN
6riX7a1HykTH4AUP/Kp2N/9MKIjzKbd3ADYqHR/q93w46VYOcOKuZy50LoHeyhtB
lVgTu2BkrmIsg1yVa2vWsD1QQsdGoRJVIZY8ftjQmFQXaB2q7Aa8PC4HxwemBD3G
Ssyu5KUmEViqJNH48MSRvQXnB49pBqnWp8UGocGmxrLRy3JyYX7gJVKaJdUmonLv
ocfryNOPJnuRhEHxa2Af4YLZ+F2u75/RCO2ZfQiESXn6Q4osWdhwiB9A6x0gwZ9Z
JDuOsY48bgIW2PvK/Durj/y9De3JwrB3SY3e/d/0doGlhwozsn7ua3ZmrYRvKu3G
/p7+0r9+E8A08x3MqeKal9plwUwiz2itbWLjEb+F63LMb/H8VuWQjEn1A2rudN39
lAygkOvNqp9cJK7kyg0YFgV9x8VQYNEm5Vn/p0rwXzMsjC/167TqReTh6FnQz5ga
uU6uG5IftYDE1qJfCRZI9lB/smkxu/ZfGvDDFsv6R52jYBb0giEAvnj6Gcqr7YDa
KIBDHn/qjOGDxmv4hgz7l/MrmBTsTyQItVg0ZA/2WXcpZMCoc0Q8ABJ60BmqmAUo
/q9dLrv0YrmLTGLjQpgsyK88kOY5LqUxxnzGyz3XD4iJrftEa3A9zRcrByTvc9DJ
/oO0gycafsnn+2Y43x7ytM+BaJ69oADX/hzbQYI86VFZFT81kZg6PlayXO+bC/kL
OsU1rsK9PJ2jlvUzwKrngMb9f0gHdS9+GiPq+uqNl2MlkjtzlGD+NQyjVL9haQqb
cAI3PYivzSRAPUfK8oXtCtKYqFH4rNGSi3+kq8TBzPbVoy695dWmoSZJvb7xwlyW
6pbnlZIbOKtP6t+grA8kJIuqz+E7KdB0g0TWMMF81qYGtE/mQgeXG9WWzF21slSm
uYBmFIsreT3+tq3gh1oSjYzJEmuhPES2zg9SLGJKO4SfpFHtAzgw9bUneeD4+Z+w
fMu0sVaeeIM49ML1dWDYUkdVs1B+c/w5kbmtyvnnvGrnYOqSOOMudhvhM3pIl0Lc
CNNVfxSMUXy01rGG1xWcLu2vvGGYZ9jFvbx2K0liKFd2tk49EgT6wFfWJen8KBu5
J9T8HqhI9KeQgwoPpR589ZkNlMLJ9wQgCWEEKD5O3bX8ZYBpCl1RdI1gPddb7LbT
GwN/Vw5c8fKDUxh33XC8dODP5ueeimMD9A8fne3tyPL1BlvvZNKs9Sn0m2aQVoFJ
d5rb3M9L2bMM6fcz9gTJYayBUEj3GirrNzYQ+/36JrPt9iglnsK9aV8+n3zdxlvL
hB7WDfps5jI6+EwslM38fpPqN0k8sNd1Ev4zYrcpnt21g8TZf0181UdeZhaxkNPj
6uUP3qFJAEqL35WjxamoPNEihmE85qqISO9EnHfuT1hWRrQ7xMX6EUHI+HVKFrdC
twt/pAK39nl14jCcFZpzJ5370jzDfdHBZpM8IfL8nRNAM976Xb/ipQvEVMwvKbi5
1ac6Gt7gQyFmYrniSNbdZz/XRPeIgcnapBshgr3Nk5vclKmQj9By6p48DnHGBDni
uvqqWz0sNXIwG1W91eqVW7x0guknlmmce5N0TbYL41kSzAUkkwPWjvYG81JO/ETd
9n44XMCfpxv1yiMWUS6ceqLmjhymcehWch3bFl+4eFBsmXiCo8WyzvjmfWiM3yGZ
ofy7eQM7EhcxJhij4aUgDdQPs3juqay5jLPnIPQsy14s0kKP/CyomqCGuA6VbYjO
ha2v+bMN0aJzb10//oi+VumoLZqMoZRqJT2eNF8bP5KH3Ji5uZC8xBY82S3u4vF4
7NGkVAW8HV+HCAIqe7BZQalCuYB0exqRYL/woetzN7MvEAYtNYrEaDZeBZzo0MIm
xJbzlGJkrygwVMQcWkumC4k8WLkhIRMHDqciKQUIMEBps4tVQXZf+2nSmWIbx/YK
5oUG6VGfXQUcvdYfVHqnvoRMAmiiTA4iIayYn0+2FFNkOJhlH9vNqf0pcSoesvJm
wzYVbUUOQDP6zaUsUrm3Z5lBHLMrYOj717KWnL8Ij+0QY275e8ORlX4+RC7O0n0H
PMf40bcO/6oabBwhw8Hcjj1nTONWYclRY80libilpIeegVx3XieeHeNHcPAZ/ViL
3xE4JtxEowCd1bXlDDH9YwKGrjmvOconwJVfxtJr3d+4+pZIXwIhfwyCkV2EqMIy
Up0nhg9YsQfKX6E2uvtcQ3Jd6hUHN/Sjp+cDYjeNZxw9hLtPvDk4+C+J74CaFWY9
5xghyiogxMivEG+1Nrdxd58yEpj8DXq8n3aaV/FAEvfzQYdi0XXb/nGCKSoliQhB
BERaat7t6NvBDSrhE/PvWdtV0h50LYF0Z6W738QJWUeBUTnR2fd0L5e87yrop6Bm
LutvuKMXjcbPt6RulTukJkAcLXKuWP6v7Z/cvprxPTwZDokvVjWZeZ3LV7Q2Wc6L
cznCcWosRx2oALE8s05s3YEAlqE9QhjHoJ4ZNaLSfIb8oCzwSoYT93ucn8Dm9vU/
D7Jct79OMkbGFNQAtEep48/TR0X3SYwwDIPLVIcUCxmEAzPU90f4/y8wPahIx0Uu
o6gXhrJjhvRd6ZClg4faNViaoqMGZj0tEviuK0knhLvMRoau5ryCs/mep4LQR2Wb
61PvpmC6wRQNN9e9mN8yO1ujz8OulBgeTokQIN4kgNNGY4BIh+OkCNnykrirKZDQ
6WakrtCYOuPiYpD5ebC4s4c+LwSIhdQn7VOcgEsmw8/id4W1scvsfjOvM04EvroP
J3YdoENANJWF5bZcHQbOlH7GmMO0jbpXdwY8rwoMLyXgcgeiAVWSAwmGlxqzNQBM
3R0kHgRovI0KSH/SkLRsxHpeI4f+T9kuUlyn8AvNHfH+nbEhm1GpygmNmdKYssS+
xMUuSpty7cgF+m7OF89cU6aUSLov8PVy30rfAXW15xL8IlqIeurujCifWmw1GMAg
sri4f7U6kMqm5CrrIMWT1tAHd4FTcvQg1Ncwchho84Tbt8WxO0wDvyyYGKSFPFgZ
FXscFlYMyXcJ6mnKtprykf98+IX7OMhoCzXIlLhFxYQfXXzW2i78AaibVa7W/eJS
o3NfQM+dDnsEc6RCHWZqUd7gSB2Fu1rXsvCJq2HZUID2YD6Cfb9tKHAD3lo7iRj7
r0X5FBY6ewljoRRoVaDCpit8pnjp1di46SBLfM/q4gxYKLvU8nseIRIKBiGLGe96
Tk3s/FQvAgD/eJel95eIMx+X6j0WCHAdDSlqdkuOc8aJgouStMK+Byg1pb++euuC
zRZls0Rxf9zueMSlwGsIkDMCS8rOtNEP3kEBthd0ckNbp9y823x6FxMQ3TTbGNee
vEZMtYcbmaIfBsJRf1b9K7TLHb/1Z815QzSVz7tTyTkeOgIO1Qlo+RYObE7ilGN2
UlVrlAURC2FpIxN0kgiOb7wvZOOjdLeawPo8Gyb5sLvi/KouOlLdrc00CdA2Al4J
ok1QTsp4GYpZYEX+4iPPzE2lTfwJl2310iU0dBZl18uPZOnqgXRDBPxSuEWKOO2A
GZLl8MBsuqMRYP3EHuPXNxA54x8gDWQ7K7hJfgBeyd58OqNSZ0e5YMjhdCe+4jMn
51c0Coi91zRVMICDS7ANAd6EScLQcNRk4QAyWzxlOtlZIZ/IewM+2xRkzHjUluUE
3E+tXi5nx6KsEWHFvOaDV2yHni9Yn6nvqNa8wYWx9D2kkYLiz3J9UVq5IVxM2hGo
NXsLT9LHHLjzv5AbfPfSO0+X9ybGd6CWqBMHpHs+e7ugDVLOMo+EytutxVBRMi26
qdJB8UGv4j/JB7uwmkcc2Uo3eeoYQreLsi1yYwmEVLklTJy57IoH0/7b8IqSzw8s
3L1JIU+ygLenIgAIeF214DKllncwZf5FOv8SAz5CBu+h68wjHuPWYbq1PLgKhBo9
v4Jnz8RbtwpBP+IUBgcBS3qBPnqJtOCLdTeYGVBFStGwX6h4KtIpWo5IDwsUO4lA
rqdfXPtMn/8FKuiXR3d56EiyliMoyeN9m05snpMt6f1H51TiR+PNHkN6YDyef521
bHRgTyWUJDE/+Z5PzXSJ5RG0apmQy7HIz9lDoA2IlUgSzSko8qTL9EweszrtZn7+
pzfDc0JUGtkfqdix/etBbx0Eryb47gbN0yU0uWMsgv9jXQ3qsRp/wJJVEeNIFAHE
4VHltFYbka5hWMkhdDdLp7nOZsctwzZGjP8Vz3BsthVPT4TJP7G489Tl6QO85CvQ
uPjU2TAifSb7jA6UmDO0Ih7Gc5OiqIRJe0DGgGiLvYgMnM+e304dwBu7WRLUknQm
BUZiSyAeNFI4ViboxobiPiBo+ztE0MYt2ixeuAV48aD85OHrsP8836W2o9a22iKs
2WCv9oK7aug52VWkRt3oMis2fuJVsNQF6SNP7D8hcM3eDdQv0xGnqSHXoWDlEvrj
eehsV2Ymwg4eXMLAkiuPHJMejrRrdtOGnmxy3NaQTpHbq6z/Ll5gOGu6fNk6YATn
Uge6W2CdiS+GYf957YYsriy/uJltOU3XBfbdnDsm2BlNEpoZMralOHHmmmTTAys6
fbAU39zm2wHQ41oah3LHdrjzaq//yizJTO5B+fZLyTm63GNuz/HwhSLg2llxFjuz
hut0OY1vXpOa80i1FrMwqes2AMLYs30mq4qp2aScS//wq3GlU+svuwC3WEa+nRC6
UtbCp9HwYxUCWUFcE4hew6CEqQAgeT4eZY/oa73oait+osXXAuZ9P9XaEd88ENcJ
keH+E/UjmoWfHrh9OthgJjog7dExXUhHg03vhIixjtqEP9cEaMehN406AFb/U7Ey
DdKaioGf7bJO+2kcMtM2IA1RxYyaNiYq+xTsdzLz7W4WgaJ1NjHovX74IJNK3jJE
artjwZtbYsI1j5n1c+08ZuBXR0k4ExPtlXKZc8xqJfLiR/KPVW7VEg+zBAuNfG2Y
NmG+Oe18dXxHPKx7xxoERjPeGNeg9H6It5dUq4iGzZYDcfo9JYEhkavwvfDIuLsj
994C0pTtAOx8KaIM+f4FBRIDN5Mokgs/ixEvMknqHWN3EVTGfQg5/EsO0paOnF56
sBqKuPSl/YvdIC7/H7p5epYMgd/gFuqzkLdfexI5A4WIZHRpO7uiiqls8eOmF+CO
u8DGFoYv9cpIwq4HvnbK6G+SqnVxjagvg3IAjykbWXOkmi8OHpP9I3wQk/RPZFc3
XeTNgax1VZSw8C19fV2saD7vISu+L1x0SCNsM4UoiyH5GRFOlvuRo5G148a6shzM
Vd1OoW808a7AVdvykEGMeTy2zZZ7E6kyW2NYaOuMuFLYHMS4eAVqqN1wPXjvhjX4
lUqUToJaX7gaN1ItqBtUeGg8CTuSisntJ0PF0ed0ynfKMUb8cTZr5Sxz8snN78Ct
cXXsENyZpSfim2QjQfbOMoLWwsz3iej2vLNAsoUcjiJfDSOsufc/GDU9IEnbCoAV
XGXyWPjgAhrmEDZJU8A2MSkFwUQ2NKp9NwSnA2T5t11jxgd0KnQ6qSjXc7Cw9v32
mqy+od3bWQDFuJnk4bVteixh+BfS511EQ+WNghPVej45fwY38aP6Xv5isFQ95liL
M8g96eJBehp/+O6Li9bFptDrcDPAcxtA2nZbGlsOui2kCHV3VFR8iXVsng/LkXK8
iPNFyKrdPy/z1fvjaHD8hhoQVrUgTi5L2YSmPSjZVCTTsmFKGgPbMqWDQAfCYz8s
R/UMSwzNGm2LVjXeFFRSk6PMb9dyt2RTwnjB90lfn+QcVCLuEm7Y/FtJ+0nwMjdb
X1yzd3o/iIT5Ui2aPOZnP/8wIYO0DaDu6z5eibVitB3XS9AVs7e45lBxBMxe7xuS
W2c1x4F6osBwMGsdrRoA2YUm4E2PSkVX71kP1XvQT+u3wcjmmESsR8YuasMPJrya
/CNsIbabCxYJmFJfkkMHcUgWERZpPj9EM4RxhCz2L2v5O6CiwJm1agi2IBbYWWQX
TkvMS6GW2eYSyNIGagnz0RKys1SkAk3R8t5dYOHq5Twb21SA8thZZea2rhyCXVeY
A4cPWd+YcezmntOqg9VEdQvlnb+a2+jYYjwbi2FumlrSdZr3HawgUHL9O7P+UkUT
KDFLHmBPbW1GZWToDJpVK/tAHU/ZMZunJ4LguUbwGGjknY654FTk4W14fp/1gaGS
nWnGu6rNOnBxv7rMJUbTc3SLSOOOM9OhpkaEaSjNLTlmWsn3RdWNHvAoNnj4zc26
9UVPagGML686haMtRUqz7fZvcon8YiVPlxpx74RlSIu9SpO7V+q+siRIScfkzpsv
5E0G8G2mNCUt92U5zrefIZyJBOzc208SB/lK88M/x5aglnlm/bIPw1ijVLA814qD
6w2HPcaZKBdY18reCw83uN6r/I3l7xEDYVMCFa0wDLcuuJsFHsed8PucRuH39m8z
AoF2WR7Gwwh1c7ViOLcI8GAjg0xCRCFkFs2zZocEcj3s1YB2dIUGDxccKxBlDujG
K6fhsQln3yRxPV4TO9p2QM2jdd9WJEDybo8n2HLunFjYZR6MVFya8f4daPuoMItX
2dxKMS4DKNTGyJbCnAV3fjLVdiDGL3+lS0tqaTiFUv//jVemaFW6WwkIFGkmYxHQ
1yWvDlpUg2F6hDhJXQxCCh9DsJMtVcz+RxeUSSAkM6qPj2kd3yb0P2f7txgcr2ZR
dJIfRomokW9/AslQepkD/GE05J9MX7eHUee7rZyXd7uK62PN9dHmJcOGAFJhYK3L
ujIxOHlkUaPB6J00OfbZiBpkPhRTVVjEo29q7XMLgyS57AnUh6IYp4RIzFUOQZOq
QkyFe0Vv4DGaXd2CSEQoiO3AJi7ShARqiya3pXAsLMZ0Ald6cb9RcbN5CcuzLuTp
myOntUFUCm/bGgKIhsN90tp5s53MQ57a9zHmWw8wPuQJB/8RkVHAfoyrDlFS0SoA
kfaT/TttuTwXTME3DMKQM/Ksj0lu5Ijh6sfCwWo+xiVe3u515p0Uyd+UN8HS4reJ
bhNKov0wMNO6RS6ronf8Y4HITRnK4w1AQg5wPxyG4jB5WN95CEzUlOGRN55bWe0o
GmJ7GJndDItY2ja9dMzE4rWtynVyO7ry/JXyq/X/1BSwcl7pE5feqSFp/BRzZSgG
/N1NPNVckdYo3hHWoqEGKN34o7h3SHCgrKsAAQHUGt5i2eNA8/NybBtdrqRUnSQT
cFRz7ZGVV3PoDRpPonYnzoku3ESgYbN7e/divIe3BI5ICDHnP4UY/fNRFpeSxoYl
lSNu9iEhpXpOgT6+9Nkfvx5Xo5a+ujZvisvOSRu3p1jCRalm2VT7oP6JTkRO/AGW
Rf+UnjIcYXYfzoUnbR2vk3i1nmFazkunGS6027E3CuhIIXBR1l9MktP3Nq04IM8J
zqL/eBb6kVK05sHmREddv8AMbNMe3OMtWfJKV80sSmf6mVG848UqnijoXu/jWkW7
K1cWRWfWf8aew6iISCP71+Dfdj1N5aokCQUmB9xS+g9ZCy6J9beFRYwNYC1HGqZ2
okssIDeGXe+TSoEMtrT+0GowmqlZg3uWnYxMINV63HPoTJ3f+uBPv3yTV0UbfYzQ
Ja+04PXeLOQCNBZSrExV9rBv5DgKvTLz8Lf1iDpTA6tFR4kpYADucxD8R3pUC6+L
vmPJA1h+WltFk78OIbDTfUMvudeRXepyjoPB70gBkaRQkNBdqM4BmJ1lq+FFzDO/
8QKbHi/PutU290NKXIQkIgiaiKI/pGggo7x7LwajTEoHZpg6OhDJnKNQKpTWo+gS
kCi91IergOqkdbs9s9AQeIXA3kKjdGjgQy8bI7WLdLXZPEoQsSR8gj4ZD7ePiEML
5FG1LgKVNzesN8fABlEdZ4fIyhdSG7Ok7j8WcjynmfFu2BUaS5u44maUscyIMniv
DV9rrX2Afs1KdWACA3Gi6wswbg7elMeeF7S9tF6up/IH35nPP8b3cHuP9XI6jKeJ
UypwZ7vHnqAgvaARkJCsi1unBC/6Q1GSgmlHlhaQEIJLihdtsTbJRcFad16jmG7k
xYxLX26oClFdbwSD9z/8evwuhKMsXl8fmOHo2X/fK7QKE0mVnEaRKZWpAzAZNULo
VObURcB4pXzDGEwjYpYVDeDaBxZsYsJlTT6fdNzujIjjPx+v1BWzbzlfCy+UzmzN
k0DX1ffV8aEG6v7dQW2Mgwfo0QIawInRghukAjux1ycPDWZ/yet6RQKwc57LoUXM
tf9yt0i9giIcMBLOdqt3gGPrbR+Vl3yzBB0R2Yc8fw2LVpl07I7V8DlFKiDAhSHW
7l7HQsKd7+emefwUhAOOP+Eg/3caTKLd2+u9BQsNN41jBlPuuqK6bWYOdrBuYQSn
BfwjcawunfeArnsmdI/Eq226BoEM1pHBzdxqWcbt6dH5O/r8+j1/5UMfL6GwoVQg
ZmxGvVWLIIiVgA7E7vSI5akzq359Ch9lg8q2ayUzdmtuSkDUiuApdoWjl4lAU65J
I78v/foL16EkzYzrSH7XX45gZmGT5Qe9QrPhAqu1dPMjegDQltnTXDGrHLbv7mL8
k6WFkjf2QvLgTMLOUFWvdtuMpgj19xeoXQLaVJ/Kk4knOr75PM5VPyYxQOH93NnH
wERBC2XX1HXqOHBnphVkMb46SPe2eB9SvRMQ+Rs5vHdpL8667l+3IucUP88yN3GL
qDGSoyN541lwLpjg2dyNEh72AVkdDo/5UDjO9FjxeyCLyU2hY1I8c+PUA3JMtGo5
dF/BBrbTpAbP3OJ/64hVO5yF8RoZU2JgGfNSJe9N6VG3HZJiiH4luNTA47PN4t1w
g0ShwWWqcskka50oLQ/8m6pDGFSzrcToG8LOy7PZG/G/kUqX2/vHel6H0ApYE35C
PPBvFk00kXd6z4XF/C1uBw0lsRz43Uy6K1TTVXKcMp/0BM8YNsLcSVLAwKORH6en
mBasrXPy4ivrE8v5XYsZaw3OW6IO3Kz/QRfEh+siJmvxhERTmEfv9ehXzR8FX7+1
KLn3cUwgD/38ixhLOhyPV0IcNxNdDNwqXCO6wyqEAJi153YvfztlBbuNZatOu2r9
3ylJWny3oVySCW3HMN1Fsuc7KZ6r93ppDD7FBoZurrdIF3E0E5bIeeqpsk9w22vM
Xaobt0aiRhf7rByrgoiMvtXT7nOFu0LRiNDKVryUbUV2/oJGE4SQ3BRNHSC+qRqR
m2kv5Cy0ZG+mGM2A9uZcG8JTwKjVdcVypDZ5P4d53mw7yne+wU/QNTGqcIJ5fayU
L/08YGPHwAxC1QpvrPDhx6Hl6LSsuXM2LvO8/Q3af32DDLXGcA+HLRqA7ed3Kjr5
gi5L24Iu9Z63lnhQGVo4mhgsD7FHhChF0LTaFKBpPcJfjMmQ5pOyMlYRsJto5/SG
zhsv46W7PpOM4fbpcVHnNpSvprDkXL9+hbiMc6GtYY/KyOBV3GwQcQOw031YiOsv
OJJCw9BJ/6Sfpk/lUrHvK6NempJ6OzHYcScQErONx1WfdoQ32ZpnjDdP5EmijTBy
FXqS1hbbZf5425kt0DPnstDvGlNKJ1z+cDCYbabybZdFP9gB/NyZWnFVUA8I/+rx
mqdA96D1MfMw4QteThZaIaD6PdKbHOxwfutcRJB46B9pPWMkb9UGoJwKt551/SGU
QKjwJ898bXDm1r89WTb22b0fa/KVzBcqhd9OO5vSaYchLkXWR88Udu9Acf7pCjQa
mabk5bRZRJs2t04DIbfrZ0lAJeCBqaNGZjpEZMDsxW/CkEbLUn45JlX0cgJa+z1a
ZkqTKQK8ZG9iHjisjviGdQZyXd1JbB3JTEmGVuTg1gAbzUx7dWilDzZqTkf9HBTC
lSTdr+c2q0LA/PsiXhpSJbFBY7kR4+kEl4Z3FitbW35i6nRno7FTZu7gEt5368An
3/0UvG0NGyjsi9VKhaWL6sMh1FMLJsploJ11FAGNzru6CZ6457OUcUpJNf2sSgp2
nSHM/rXB3tS5YyAWJcS8qYVaMzm9BFVngAWUMaiVYY1H0kONtpYWUwWHzamHaLxq
BMvdAB9Ja2jCbnaD0XtvUiU6Zsp32oj+78aW4a6JQz+X9e3o1oIFxIGAMdTOTlVM
XF0/0AYHv3IslDPmfn/Hb5eUh3XiI1V1tOTMWXhOEopEh+Ck6oIk2tbAz62OxpG7
ZvtBjhlLMdzKRfOFepVZ0OYd/fotgLnHWwslM5i+SqsQ5Jr7qtGl3IKljPpC8lNz
C/EE/NrfmURBXCsnHU0HqCWL4lbFZe8U2/JeoiyHGJB+Qb2+HtWY2/Xmarsvsyen
3Edf4BuvAV4JHjA05xjaSVWZ7hQ2ahmcMJswuamhWfvNiKqTZMJfZLmkHvIeFtaf
mp9KTYK8TSjzezlKBz89n2ZvsQvEBIGTzUxB1XEfMgAoeI9SYa1tQlON3YN99oNU
aV1kxMGgfXV7gTdelyKtuF9zjXN28Wn6WOrOz62a3FP8+HOBPS5Z/KvN3OBdOeKZ
FhX/yCiaN5AuhTabKGDRFC5+0GcbsOFELeIyt1iTQ6ZGbJnTZauYuQTCItMOSH2x
NkIx3z9Mkh65n7cAvYq8X9MMLx+3Nh9nt4MydPkX8zWKDZqn1fDZw2AqAJfeqblY
LXEeU1ilkWPrxS97aZs/CodSWUHKMbrCX7ogMCDUKUVIcnuknNCJgIPZFVCLwoXR
8CpN99YP370BAAQr7AUH7gqnKxqec4/Ao0oIrSWbebsTqf4daq/08JrZmQVjTzDS
g5O1gAdXXtoJpF/XK9RH145fZZFK4BMtJZ5aJlDcDfwOWTCOzUZMUmPz9MyW79NN
eAlujQcPOk4RZqwmy8EBnI+BF8t46odiJPb+Gft395k8Yw/1eMyy2Ct6Lb2vut2x
zaDRPCUxbcAASdRSIpxRjPG3+3SNY3P4OcTv20Sgvk9AtjIrikATzdgYPp1sJzaE
lz18R6B1w1k9GDye3gbx3rYWf02DxAx7qlWMdrrLXF99/F3Q51+ZH4gIff0SHAwq
MbuJlcAtyGFo29M8llVnMse8yNx5mrC1x9vmxpDjjVV/mlCBepG47W7S3NeB26yq
COcgma0JKk6bqz1Q0kbh0HX6ZjKj5LtM1LvlS/k74UT/WqtNOmqp92yxBtc22etq
RmK3oTQipHdHagbUjA+uIUWMTN9SuU0PKJhrDD0AHIIiYgH9KR1RGexon2c/tiyU
3VotjcjiQ9Xjggp7xYGRTFupaBeVhLWNRirQ4bJOFRcc2Oulk76Osz9pMQufKCZ0
FNrDhvkrKOSRoA0SxfSZfe5BdZdGzcdW4lgeec+80b6RNKSyat83t473Fwhz/u20
FTt49aqBKJXkORuqbnBRihSevNUgVcSj+8dnGEaiCbd3dNwsqptVsjFhXBlXn+q4
unAL7tyAc5xRuwpQz1MfrieCo9BYGI9IaLeSnTNevvhvTWo1LMWI/VWLocxjlvhk
Lkvu1+Gjm9faW9yFDPtQIGrkOyL2u6wV0LEk4C+S5tq9sf2Reet/oRCEPh72HcsU
sXo7kAriPsXTid557xIoYBPubKr4gvHTsquC9vlTIedXwFaMiql2xrw35VYlFWEL
W1v8zzPQDTB8ImvO2GOc7u8/JdnrwkhCnRrlcgXPyi7y9KFO2fWSPaUUjslbCogA
SOaxAHm8lv781DGWKZN6rfBMo9+lj61i6LZNUOcuRCR617b70Ae/uG0JVvDHzjo7
jJEXPEGpLC4EXHzsGbPNRu8hNFDxg+rNxzGz72/cXHoL0NZDY6Sr0A4DZbHxJPqX
trwuDZ2m3VF2uLHrWA/Hd7ODpR5W5m+aVJmoEjz0KY2so8Ky9VKKv2QzRm9qo4zC
pbMBDu4pPXiW1RgyQaTh/eSRN/oJGSuEwcvHkUtVCWdMZ4AF8bua+gT+GBeNoQ4k
ytPQuA1L+elN6QFROWgVlMZlu/vMd3GN1cgrS4NwT/aAKl1y8Di/xGI9nZqhUAX4
aqHaAVkyMOY/siDWsX4CEgcmOT+95K73elSNP5XsXwYC6Iq6lYS+I0XGmu9gv1kc
Y0VzQCGNvPOGXOZtzbJ+k81bSVjC1zrcFFeCwFdoXWwyAWIglVk9T0u2zonqujnY
x824/Jl28FqW2iiec1CoO1lYM6ilp5vMiYxI1eKcRXVKKlWho1S3w2jM94q5wcLW
7rjMDgMU8IztMe9AVMGC2ZqchUxi0LtsO2QzWUuLrSHQl4RGM72HTiWnYTPbomr8
6Oh0cB5xoxvhcOvbg9OdVbzGxWxOUBtG/k84T8JaHgTr4AUxI6m1chWpa6nt1BPX
nBf4r8DD+4sfNYzGQToXSymmkH+am+mpijGPwVo5UDMgxnJ3THvK0/WF/NuvR1qK
1wHomKCEhpxmxD94hbVm5WApqNh5oJ6AOtL459QdDLgCkNt3r2SE4NSIrnFoykjh
rcO67JPqiaF3mbSZITqjE7dhGULiS8RrCngXcPm9/hdoNwq5Ji8tBWG/TL5GYCHj
iC4zMs/tVJ8gqa/wNW8R3yKP7jnHWmkZufy9SUyuIGclen7YCPrqJR8hbCCgQvSF
cfvSo9R0Pq+mSQM8+mtp/m5UWLHPOrXUf6wI+ddKRd81EU8//z3YmvGTHkJSmn9l
nuOcKPnbEvyZB3tLJXWjC4ocqzLeFGrTJNHaducB7upefoc/OtQqwbAt/vzIPP3l
rShz2s0MffegwOI3XRZtvE0R3E7/8fl2JwA4p/45ZSr3U9kydGfJUaIiCbI5jtod
va6FwnAqzbOjte+mdadRsaacWSvBy6zVEQyEjTSsLoJ+au/Ri7QN7I0xc6J4DJRn
PP8JSdS4W7za2fShqHAYFr94YmcdE6Ose+KKnKdl+df8MOa7dfbv95oRN1780f4y
zoKPepoUYe/liEbIDVjlFekx1jz38hTv0dDS19Y20ZKZrZwZ/VpCtBWR4G6NK5vA
oVFDggcDtz95z/THm2mPDT/O9Ek5+8Gh2z98HIKivSdldf5Y9BalIG2gOleJKZjR
v9TfVYVbOiWiV8Ze8x1A+p3r812kdF1KSOT+cXjkIHHFjEyse1q+YKW0EXCqgX+W
nkAKCATeA/jS2bPRbKcBcdsC/BiqrrlY03ZGOSoYXpxniVrIvD6EP2zaxFA/63nJ
aB+glhjWFXB8N80Z1L3Fy6T+eL29WdBk/b03fr15Qb/UCBHCw7n8HvDkyCM9NK23
MWCcOJdZVHqRgCeFmMZxLgYhAqkqDMTo2PYoILpfpjOnAlOOVwqFBnVRgd6r9xaJ
Q0ac2xaOgocwilbADqx0mPyZlkrS+ddozyb/drGlXktobvoeLMCgTqkBo8ePcr14
hVbJyekLcrpRNzmAsNwHwlj6xOHHD64mh6O2Dv+k+ycCnbs/TvnjFXLRbTR8NzAs
jAbbVUtfCQ1Mwtwvl27xijQU7nvXu4c7Vwc++5wrFXeMKBFBMWmKZ9LmL824qE6F
lllRFrDK3cojUKm9wy/E1bIyqAFMuLIvSKTEaRNE+ep1tAxtrRIJ8wYMXMblCUQA
uCoIZsyGb9jZrab9POK+om//eOx6DquZIjeilymfNYxkMnmJnvtiTDZu6Kt5qWGg
HVUNgrxMsSyBDbLwzwK4WC9uW2jyyRIqmn+QDCtXMzqfDTi5WkGWVsQjjTYSywDo
NQ4h16ZW7MPp+dN8Rps+SA2H8lmwzjxDtPg0jXkyvTljaVgqJ5gN/4TBz0YBavj+
oQ0kW4CJSatZ+nBc9W9IPMYT2GjwbK9YNBqhNOkdEiLXbQmsmfIgh6Hnv5IxUA0L
FVQzIHn9GqcZEVAV0b1spRNVw8KVUmSR3+DpL1bc439u1QMABT7dBMnKWHNAcrac
NAm6wB0IrHjLTdcFBv4mE8YVwFOEtZHFdhix8LPda22KMyV6YvmUkh9Z42U7ztcV
596NIESOZK00LhTb8KQOncofkFansOE7hENgN1Xg+xmdxuXG/O4+bI7JdutOe0T9
4Ik4ZLi7qlSUMBqye+JxrkLx0qh8SLCGgjmgkWecLl4yw2i05CnYKMVdh/K96kxC
4LcGrSAvmOoEKK8sWi+jOfSHjiDZI95bDrp7d2vUja4EPLqcX2Ow+TBwNXBGms0+
sn846Qwd4l4pJ94B0Dim7tlmgtKfZe+k+NRFe1K/uXLo7EGnVZ+tvEggjlvR2/Zd
+kfN0m7n8NXdMnko8oOdWlmfBAbF1WTwwZ9MQ2XZMKaej7Yfv+aXVP0/QP24k/Hq
MWqpEamG1Ru0fCltlQWcyC204v54duGDpksAmufju40VEtxNAeDt506H8aqmk4IO
IDjkAfCt56Nvhg5a/RcyjxwfO8fh4f/isUNLCaGSb7KOT7tV5Am8kvYYAjyhh+NF
bm4cHcCDIOrhfwp0XcOiqFWV5t5eB/Nk3gng4G6IxXQFAWXpWVa1Wohj+luRXLJL
LosE6RLaJHX3Rh3YhRmtlJ5cYJWOZ2pGuwhC95LIeDAeYVtfp5TWPK92ByqfWqYH
hLJqqMiU8hrY/OvzO08c7QPZTONE61e/WRWgrroUkhJ1xOK41nmVjRS/0SfqRk4u
73Nju0nk/8kSlavFzSXKPQwynFS5VEw4Gqh4HvZ5/XXhtEVtgXP7/uiuEv5VmnJG
SNkKUNjjj22GUysyNGZ+bHn0GG/eMdlldgdf/xIIiTYV7aoZ+K0xoosrUeh5Ll/2
nxahCtHUUlgSxEtXpPwxbGGfVmMYWoSJPbagCQ5eqi+BAHJMc+vEX0l0vILA8n/g
a9SpAIwqSLcI9wJdTfmDk1az+QTlosz8Pru30TdUplVtXtp+7ixFBgMOZlHvYZ9L
V4+DmM1H5/VtsAGE5gvz8kIvFibKo/mcGJ5GRg62wlfOv+fJphTfCaUEE/eSUBT4
1lJMgQV9EpADaO+AwuTubWOoPNSFRhznhpkYb1LqxIJyraMs9ovmnQviq0uaq6Fm
hsqp4hYkP8D11UDF6Kv0o3DNp4K1JkhlAJfqyYl2OSDYkuHLL8TUOdouztCIufa+
xEAzNt/K1mXq8leDt27fNk4su2ziiukPf2lGU3KbEUtMGHHsCH7VaoNhHPm3cdd9
Zc7WIUKA53dav2nPkP5yOGL5C7ztBzj3SC5Eeb4hA/Oy0MMf7cuhQMV/eqnp43HM
z01NoaEsil/De2U1BWD0Nt4D5EQeD0GLDV3pYMgs74lERumvGTTjIPGm3XuD2Ntk
Unc+b2WNOKCKjbRFEFReOC4R/QDCk82dozEIjoHXjjya8vr5AG1oLFIpjumBPSR1
lALiSmtNEEGg5q64SrTVj17FF2ZAAPFaFkcIFz0yhDo339A7o4d3Ft7OBS3zwBCr
aw9dZmgP/Rq1gUnfjd2ACCu4za2mcOi30qg70WLgQfQNWuFvn6gDrlPW3hWnNbsv
sQ+XRnjL0mqqQdw0LGJgnkh0KSh8DjYuZOx1Z9tZ8uAjnMLP9te8/fP6GaumblIk
o36PI4GHF78n414KtovEV6WK0ExvrI+20JGKb1Fy29BRbjZA8UEABZ9pIjJxlQnS
bPE6xnmGLpgrxSih2i5pOqTavua0KTuQWgBunxftT7+NOTGwBOORU31GU1nxYf4s
0EXmVdkfHogFNz2q9Eo51meYxJv7RTTD5Jy9aoWCR+iwdaZjMKTDjfb0QZnFKOzK
ztKE78YlWzQi6huihA4saohSnDnKSmXDypfTw05qvu/NGToHsyOAOGGkFVQg927o
LfHJN8Lei01UDisWEXdvXlFmjsmZXaqrBIThF5TVU7XWr5weqpZQeuehNk38dJoa
pn+pVOhpmwLJ83xfGIbMPyETKfvGqh9y/AwqGBvyhuVOkjZgv8DUJBRZgD/jlK81
yXCsJisvAAD9w0pL9FPM/ABsiJjG4WHlZ+JPscItep5RSMW0dMcDu+vwTXTFqrvX
yec0M4x5K9p66e5Rqa3oZI1vx4aopZUi6G9Svgzf20szPGrBOSNUgo1dni3AXw0e
I6ekPtJW8mIPKUzxE7CwNR1hfQA9yB9US8G0A5qO9KFG37Wox6T2PgKiTGz6yKpv
JU0G7I9U+C0z+l3MsDCZ/GiymKN1O7DIwtatd9plGdtOiZzOtITc6e2fH6ykOcEU
PM2g3zRpVpO6hEDMpU+Cs4Zb8zBnwClaiLGKlulWk2mrWGmFyDbno00obXigX0TZ
iL9/NELoR/IvbmAaCX5nDixzHRlIPXp4aVovwhWsmQUZ+KAmpolzk6IDrPAdLhMV
h3W0BALSPITNgswXnx3k2PZIC7ALO/efWymt3t8uzSE/q9rg3YLZJq2yGPdlUrKY
fMIzGRQ/yf3mJ3qqkKCGyD8u2fA5UorPsNOXeKjb4M+lsnR0/f+iaHN5VLb1u2J5
ASRg3YqyJJJThG0IU9/sWItnPx/T+VXnL7VJM5/mDWLDnILdmChMhhrAAXKtIsQe
+0yu8nGtQ6OnLmxeJGG40BAD4V0Y7A0TveS6P38AQCWpgHxNg8IR0bfnBDvuJHk6
YwGK1QrcORKeVrdy7A0u8QQQBvlf63czeJdU5YfSgfpt+rrUHqb0zAxNT5c07UwX
p/gUBtvYCJndrNKjd9UqErved1DevRuChXtg9tg8YyO4f55IDDwPHZAS/67gxznr
bYgEjhvHuZd36/kkVRbSU/OrEjz41Sn943XwnjxdIaApNjoNhiTA3T++EhGWc/V7
9eAQDz4ORkECekdp2P81iUb9KyXjzb9o3o3l+EA9z7jDsXOxuC7sJos6x/HY6aAJ
oj3Sa6H84rOEeVfGrAWkl/wMu+Tl+uKAqfwhYcnThrWqmAaJlv5P30pMsLhGKtrS
arj7Al2+HkoSySrExG41zGuOHo3Jo90oBBovdIGAQbT1n1kXPJADzIUq47w0n5xT
Au9BxMeae5/gSXK5zLpJGUXIaVPDf+LvY4/zrj6VvgfFLu6xP1a0RgPoAqU1Hxfc
JQT/SosDaw9ZELwYMAFpRHqPdBs9YCWJ7o0+phFBzwtmW3stzIg14aHuxV52pZoV
C9DoiD2eNc1nnA9EACM0DwjoJ4VfiQOXkpUf3+bUxM8XxHKLU4FgJxbEoD3zzSlg
JysN3CQuwWAyB0fHGDKr9OydAGBoRnJxFkFub0RH2dpwd7onk1TEfwEtpWXrWEcK
YCRkN9y82kI11h1+oWMb8cKQSaz5XPUb4gsjSas1BfqNVVeGD3IgEWQNQHTvi0R5
RBRJEk1J61uapDDsMJ5XoKR/QVK61EsNHehZ1fCYrIwO7nYQjZLe1+HJ/JdIH0GR
VPPXL8rcY8hvbY1zrc1aRriXxP63OmsMRswOYvINTrdHbrKhyUoc4OMN7uV5v8YL
jHqy8yRy+jxQrd0lreL4mBla3XZ87eya+Pki2dUG1J+Dnc4sbEkExILly9hphDkl
8xQ/Udy8zAoZF2zPMm2dB4gz0axIFLGZrLA5n3+XMB994R8kIB849EVN/kfC0bnN
3SxTQsCyJDhjSZ6ybbStKd/31wvB5hQ0Jbtl35P2qpkkbky/Ptk+rltNGnsABN+v
Og6LNJhcHHPDjVwdjomTGursr1dOXQeABxFd/b7/LHOU7Ht+n9BebKPKF+dnZoKW
ckvwfrPMSWVhV+zYcGdj5zIugvO+xN0OZUHAA31CrblMW/4zXHw1ydk/lLhGWOFv
Pq52LDc8aIgVs+v5HQl0H5vpVig/CTzRZ/4H/W8Ba+rdriTEdBNg+dNO+s/tzPvs
m/DNHoFG8m0HNoQC0zWaH17Y0S4RW29F800VcoDSIjLcLrWbrRf2TYffcFPjbXEz
ElqCcbKtA/FTVzps/BOiylRyf3Uo4NHYiIb+Ws5tLxgB9aU/3dgL8wnGQwC+ky7b
SlfdtoZZn9xrM2pkyjnmSelibqBLcJHtLJIjVr2BAkVflTXrtfd3iWW2FEoSrqJ3
8LqwDhYFgbCxovZOYPvYsiYn7mw5ICD6jrDQeWaCwZaqBylvzHtaYR6X+70mH8nw
r9YCSTet+Mg5S7Hw2u4kBLbEpgMb//WtZSVrMN70tqygA/oQnBT3kGxcww8blRXr
Cv0Ty5+WPpYNzstaGdMAOqUDg/pD9DAvdzD4LjxE12CNmEve2GPIxRmSy3W2YLJG
xw7YYhI7nTkwH8J52FWwpENyJd5HfyBo/X4/dpsxurOl8FgTXxW3r4e/G7Dv5lWJ
hi3wTqUk3dXIGQDuoLmBgyrkjoZw8RuVNTgoeGYhMw7tvfcciAMMyUo+y3YgDKPv
IXRQNeJS6hzVjmStXtDT517zdsiK6l85WzhUIVa0dspKvj5n4vIRIKPSHF0BIlBj
slhAEFKx1HpnDva7cF2L8eCQ78cEl6fgfeh9vyb5MbqioS8l1y7d/psEpCtt/Pyr
0r4qpBJQ+e8DMx8h6RsBrqARxQa/ZS3zhsCHPbyH+2UPJqb3O3J/gs7RoSLrFZAQ
F88VMH+nPU0AI1hs2s6CugnprPhycWzH/hVpVQRBiEoLKgQovTpG/OM8RXlRp4WI
RiAkMPXgGsHlbT7Wb7WXVjWjUCm0swml17mbJxauYu6ziG83SdoNLOe3kjcwjTUB
43nGkAt2UqE3gM/e3XAxHz6m8MRVfLhRPbK2bSUci0t1aiLk9UqjdU4HcmTA+qoZ
ajiwiJNKwoTNWaCP1os/ZiFd97PHRkjeG/y3Ta7OiCs3z3dc9HBajI/HSFRlIZV6
9RkAwmUUeJ+2dqK9J1UPuIoSczaCAbFWtqtfrmwGBL8LTJLFFc3fbGUmG13oRqcl
g/sklFExmS9WIaA8G4F/KTRU8+k7BkgB9XfSRfB2zwQbBmRTkW3nno39JFSXzzTq
uePndgK8UxkAlTNJZGzvUZ2Gnck1hgtty3fggKzJSpAI8J62g58m9P6v+hXIkGkC
wSplD0stNHoVgCsFRHoEo4wNFEJ50tkpadQlx42+z+STCGkuQqqKX+SH++YPkibp
0yhexbUhe+YQ6O9LZrzQITYxzlrwDLM4ke8+uiyLe75axJlTixDH8bmS3ki8NzIg
gDaakPp7V5+wxjRkqKhVVs5wK4p6F3R7mQOm9+f0lV1Y4EesFBz8oYTrqkjd0O1v
W9sr0SoWtI4YQ4Jo5FJvS48Y7Z+oY2SyrhS4RJ+9ixnmkxNNUeeFQ6r1qd9PmxW5
9W6X6ObL1eTcWXXIRNmFgAmZlKpkKoMCeMNK7NAPcnUfmW4mT1ASVxjzee/oQVl7
gbUqm2IkQhFtGlBxFJIBdHEFxHLNB0I7lsT3qW6+x7vc9uHFObcmeXBPqO4FeG4q
S2jZJjWGuqYkfTp6yVihwA9RhndKd4eV2gpL9Pg2VTYYyGrqmpr3XixWfRCbajJa
SnWxevLj/Fs9VXLidYQZD6lDEtvEk5HWTDkESMjKHwiHZA6Xdrjuo13U03LYAkPq
f4ZZpHIiLEo2XQffQF37qw1EKikh1YI9rpTX2BVfe2iGfE2qTK+ugBgu6XB3gCW+
uOLaEI08dzMYhnC9xvP/QLeYoyEqWOUZdoFOZG4XFtbeYEL9MBvhF/jaaD4B46hc
le2wJL4dGRhuTzI3Xb9JF8uPAfJ5Dkczi7yMtoK9xG4RkIoN611fT1HKi1Mmqqzh
aeV9H1edv+St50J5HECD9LlMA5Nh6QZYVHG8/1kBOLWAttZOXV7/sqfHpeR9CvxJ
3QJqi7kTj28Q6xOVN+q5bovIVku/yAyfivLErVgtwJ3UfxelrAyY7QlTO7eOhE52
UJKvnio9Kp90fb55zVBH8fqxbJl2VtkUGGZR3LIxAA9QQDKU6Ud8thjZlRAxQKrU
1M6Z3os/lo4ufx7R7/K5u0z3wW7yd5+SIgePyPQ9yAmdA9WcZx2RhcJ0XVNyFT+W
c2K2ELswoGmo/RwBdOVRCQn0hzo20TQVQMRoTYRJUAHOMT+Mh0jrZHwN/uBPMGng
QLQ8OmKRZIaGgHqDVhfcleoR4sHFg0ngYa11vptUmn3QDZaJL6UQ9qNlPBaN3LcH
ZBZrQgME0k/VZR/NGSmo1oeTU0RBonvDC11E/IKTsUjk9MwOUNvI4KOkHJ0RD6Zo
gi/HGr9o1QGFTTSzdi+pf5brq+E/bCB7J+kGYPdHpgo1/o4GzyAVDZEBivG1zP4q
iPgqIh2a6EvdN+x92+UAALQb5iP4LtR9L2x2POw3srE4/b7LXzNCD3+JFAFdRgub
aLnYGK+a16/JVVPQZlOpf8y0tKjDUhKQbNnS9OybdowidTWFhIaB9bHHb3O/dQyT
nZRDMsg+Al8ZC222NBibMOjv5CMH6wcii2pTT/Ui/xU78RZW6+pJIIyYaVwApzl7
+dG9mwwrOPzkF5yp16tdle+LzdZOPH+Dy7fKuDb/GJnjh+aivYFolIJgcCBiQNy+
d90h6izX+BJk7IlUBWoGjfSQfYw8UkMNFuqqBgAv8z0vWJ40iN3PlmwmkYQgATYW
ZZjBE14PkpIeS3N3lhpiadcyFluv+tFKxJsglk+OeFG0lfD/rbxBfio4OZcPBFPW
/2dCvgupmNSl2Rd2vAbRCmcL2OtCAXjlxr6uNdMFZ7EjW4SZzoMuAlqpMHoKtyCd
vC2+hNnZsdzk8GgtzxTzXgabbBQH4sRaTzQeq/PA8NDzdGMUwxEorerWZDqHXk+v
73H0tmi+/8bsW5VAxn5prucO/g6xwcuV/IqY00YT7RNEbMJTAsSBavja7GMo9WYs
FVqdb80asDGs+2hd05rIh9rNcJOaKlPGl+mS/0RL35tBLYZvOpktddwcwJ7fM5hc
Tkz5wf2pIvPFyStKpG0krbnZd1aYTVYakTcooGh6TbMLfN4FqOnDT1yGwC1mSUK4
KPumh8v9B9k0X4F99C8e2JbzQofel12XZ0M/kxK57CKDDJnRmvihHzP+oh6o6Jzu
PHvLnxwxTzMMN2jNiajtDV2HjGbF7cP0eUf+fw8d9X5C33surcpBBPPYukqVspgx
XOpqnyIRHhd79Ej734TAOrnxgyYf4gppMmAZlne9mHIl6n1kEORsFly2hkeMbm/R
xVPr1pD7MW6+5c6l/lurR6dF8s9u5K+b8nNNsXJA3gCOnl5pQ+oka+I9rSRTZvT+
aJbF6Igzx6YQuQ8iMBqalFyuBq8I0/r9A4q0JA1b7gBIkxWLyj8q4MmeL+3GLohn
rcDejPzBmN2/rLH4bwM0okjX1e9S2Ve86huC3zqpMpRksEQeSAJAZ6qIRpK4ez8v
YE8UKqgc34o87mJb2IYe9h5/X+fGH88oTsFr3Ida028mdCDKHUhHPHSsr3XjdiBn
4oYZ2c9QiIzTGh47tVwuRxLEC37dNBoDpg7UNxi+ZKhgrPENCQ22vISMIrYpWlgV
Gg1RiEjQgtKqPAUyJcp+Wko6Wn3f6Y2EGgo3kDFBz2JiJ9OrJX3aQZcmS6aHA4Z4
pPh4vo15H2JaDT+m1PMWN7YZ9zZxBhEmdSCBqmQ3j3gKwenVxzKFVG08ZVuD/nZj
cM61VjuOeg5Oh5fcrYQt/yQf3y9Hk2it9kklN3Uk+DQKqlDmxLS/QmA47Hh1RXhx
0LJ/YRcYIp1yJ0wVpNJm9orFdmrGYoQi/F7v1TLpPoJK1/3lz6Y3r5hkZNkdWM4C
JdaYdos90bKz03SRFoY+QjweuBYHSYxSsCG1zzG0NuMlAtpQChxQHcz8w5X3mLEX
XtuaXDsxVpu+jRCjc0xKLYWq2GLjIOf3wUYT+gnrfWXzRXdlEqTAy9+MDXMxc7x0
/KCBBFLzZJYZNbWRbifXcWrNDL3KnYdTzg8wlhVbd6nCyfERe6N8S+2VC2JEictL
zPZfxeDgZwMMDxQSH3tGnbqTBGuRmC+tXztOGtHJz0NV72w16trwFxUEb7WcFq67
YkTmTXKX3dcGMq4BKJTstOKyphQk9LCaGBXyDytGo8BmY5QkCrhseIwuWTYv/3mc
KN8OJG2dH0Cd3eGOLlpyOweEVHL+n0ZmIT2NHpOGPfTKVOHGooX9EhXa5Nr3oMZN
VA/+sLWCPlVS4oY1W6x3xiw/Y+8qPILpHsLiBptrvgV3HTv3qSuC1f0sqk2QjXYn
4wpdum6/twx0rNqPx78ITpg3HvrxLWAkro7nRbzymIODbAxJHaAsMpjS7yWd9zXe
BYoveMLhK1eM+XKjJB/sISDp87b3BpqHSNBykV/QnwSKt3/bR8mtzPgMRTQcgRR7
1yXYYY53yGAGP31ex5PLiO+VgAfMgNq6b7l+sYIiKgz+xE5wsnVh57/stn5rXrn1
YzmQ/5+F3+otfL/yMkLrfajdBrU2tis0pO4t3pZFmE9jWPxEZvD0EyTIUrHLersB
lpjACy5HpP9KrbHpOIksD6z52vq020J1NiGYv4UApPUDl7nRVIoxHX2x6xH/vBqq
X894t47kAZaRMYd5qvP4fHpriZH7cbxv3ROxpbNPzfeWq1TrRY6Aj+yC4R65FYV8
4JbMu4Q6tpAdoJpD2qCp1Q67VbB4miaXrtgdkLr/ZM7Ieyc43qEfZlkXWIiugTAK
F0e+c6DueEbS5Ni67PPxbiMSwoi59HR/XyzqvPa3BwigvdrIDh7WZawwbrUFM581
+F5Yj3k4sPKW+UILWJCzgOxuTfcxQ+SfbR3IkAVHoTIeEvQPyTqilu8es8j7qiEg
kiRVVCrH7svC4jmN+rrjs83AdY2oeFH90wLe9CYZJhLygSas7I5xcczzyzZeSb0m
IjkXEdt3b5w9y5lkrZ+lxumZz7KOu2aKEWgbAByBB6acGW3Qszq8zKOqzspsUbXm
aELTIbrQkoJ668LnVgJwn0LH2DUYkab0LMy3FeCADKTCkaBvoIXBM3dFwH4r6gd4
PP56zpVMDjURm1ohhVP9BDKadHydUAHdtJV5O248WLcHgcOcbbpN7bDIHIDtmHQY
tqdigzNii37gaFZVIqvvFQdpkJp0MZxh0LVnHC9r+3njDarKmxLZjRpfH4+L7IUy
jeOGYFOIAUIDDia6LxKzJkkEyAVVFJUS+zPjhIFCAGoH59DkEEsQZj/O9k4g0+iF
dNMBQLnqb1FxieRiDvXFGK2UQQY1AZ/9iKlEnPlQgyl5V/hq/rcrWY/0hIl/p8LN
tVrpix1Z6gy9IlCjSA9mv36uQeHntv1T1/xc/uGDFHXrufrrDJ665YncEkDZ/E2M
SFoHFMyMqoyyHI5xsc1k4Lg7C/PL/hlg2BTFl9OrLMJnWu9ynIqFX8HjjLuj8H98
lipatZgA3/GWZ+SlRaPJ800yOgDHQJKPbNvcnmVYIYZVIgeS5D7C9TGBJVByFrh7
6/QQQuIkuj7DS7fJbgbBGIluvDh6lFpTZMGEjAvqWeBHlasgK7UqDXMb7udMlUpf
ECMhJ7GteCai22TViqxM20oCzwvi7kSvgASi5lEeL7/m6WZ2cOzPsSxO+dKahqYi
BkNlkzu8AZncUqLHaUJsB8RW0ZuaK2rslJ7T9jnVRPJCIlPHUqk3XUt9SkTd1UYj
0cLYkkYtFwV7Gc8le6sJtECuhaMNPt4u7nMFCtdu1akhNijWFLOVLBoafIJ3F0NQ
eYQxKaeLJs98ddz/2OX+O4kGO+37SKu/pqH3+Pf2HU3P/BT7tH5L0vARHqan3/po
YwCXripugD94QB8h3L7XNiVEpo6YUJyWyAYiY/lukArHwJIxKBSC+K5ti3hbBG0g
hfVodFv2wkTXpLGrfi5eYfbsf5gYAv1j7F/WO+WgUdaJ98FVVC5ONdruHveuAyU+
JH/Rh+uWloPDM4ZFfE13OXlQIK5Gu3iHUgdJfPSzy7Wxg49Yu2fEPoNZ+OAxB0lz
/GPApvT+mkLulYKjYTddSsdK3/xKdOM2eoA02Lm3yoOEgveNXdZgSPEH9MedSWnd
/s4m87G9uCBmK31UR7NNwMuknqezVznq+VqLVxqUUgzdD+v3zasp5Q/e4e1ZV1s+
bmROVD4hiia2q2A3lFinRpLU387a22RGlKgBnQHcm6BYfhQPUqLDlMRD3mactKRg
QjevKrJYTfWMKOmkigVinriL6a8tlCuRTSKLyzINQHzLj2NvYFOxAhpXw6rKBOCZ
59OkOljpx0HDVHp9jJY8BcX446n4olBRet4G2Dz62FfM8eXqSPUH6UkkCdkFy4Gs
m1DNK06IQXG5vloWdAWuAVw35F8Kmi0TioxrghYYAzrlicov7mKGwdVjh36HM5Zo
G3Tv9MM2HFPPw2uQQhVc0T8oQMjBjWDLvilrwsaVnUijW4BSl+sN5/CBpfM7Mvt7
BzdyiJWyqhIy9X+wLiqRELVBHN74ZA2bzVciFk6dfcnvZEXsIgPYTAH0p7XfM1UV
Jmx91LxPFvuQMkr0iY8dF8Ye5K9rNALGXHk812d72VDPyyqbOhWedDxJKhe96Rhm
L1/4FcYkOr2ltZfmQJVeqa66G3Y+wUUSxAQw01fQXazftC5r05So3N1S7kkoJO0A
YZQuyLq5SP6xnKm1pFczorpfvWQe0xqPQL0IcTdJjEXfMT04Fj3mMvmyl+EiGvIr
W3YV+B+Udzolz7sl0k8JQsqurFsFKzHRGuyj+shZoGxrgimpgHJpZ247bv8VCVa1
qQwYp7KNerrlrJBhbUoKOH6om6nDBMENzGF2RQKJbx01HXLfy7L5i/OogGVp+DJ8
J8hZOI630SvyAjwvRcB3nLylZDfaGyQCWnCNEZTOKxF7rsUE5RPRJh8ldCtpCp1F
JI2tLyYF0+30NT6+nhtiCY6HWmiIz3/kIOfw8R3mNz+CmIeGyAArvkXRM2CajzQp
0tjtH5RTIsMLYtdgSurWq/Cxc61c6w8dPMHiHXfXdlD0DWwzwCBl3VVoEpmq0tVG
bDzAXjGSvs/UC++KRGR3HcmkPbNFg68NWPCpK4i6R9ZXAiviN5+BHT62azuAue24
j00iy98iuffe1K7j1jPKWA9z5jELMniccTxjseGBIEVPyGZSmcyV67whTZX5A3WJ
IRgUxCIOwew2Y3/tIk1QOLfXM87g+B6WQPiwjf8CF4oYdpik7oIiTkTlXVdndENZ
fRFzfzV9otEztVyy7IHEOt4Ja4owUwgELepJ1F2l4BOf+tAJgKnTNOy58S8f18hf
KWd3L+OaULn4bIq/2WpuD29Y9DIBBf1xc/cxcWDWETiyw/fhmdF3WECWwmGny5Ww
K0E4aHqexmkZd8m9NWMkIC4NuXY+hLC7qUqYV83rJcwZbviSzMutRiiDs/IWOzwW
T231Dk1Ir15VgOM8NiP4WHeWDZZLbdIX5JZ7TB56rXs7mT0d7rEA0BYE3L8q26Gb
ODz3gNRCawPBVrvW7aP1li61htkYTbiUKBdzObdYUGL4uDJp9qYYVMz2CN24Lmgx
KlEWrhLw9A5vBRrKGv3ejR+o1vmfFvamET5pPzczxkONLvamtqb1pdunvwA1kp/e
vQNoNxNUTU7LEvnBEMNCEQr63eIf2PVRAnrZnA9FSuxLo7FEViQgcV76XyADt4Qa
p9tcalaQ9Xkw125rW3K63q3zQUI5FlFA1n/TznAoTiZwZwM6HDs0Azh0EI8UOMj0
wADWIlqRxp1PjQDobnQmswNZnYJz1dtlplUuBXCCtt7h/iC7rm628TTDPD1H0iTv
XPbRSkBljnRit49VhRa9TdQOpqr3PBrLspxTahvOGJPN/4P4HWNpYXq0VO/wuELi
anjl58IV6zA2Nr180y0vQyo22HPNwlKwGzAOq5vtsyKcv1zWlhi2XQYbdLmU4pHV
29/qjoLV3dTqYJtzmJh6E/1HC78OYC1aTH0P2Rotrj05CtE5AwbAqevtaUk16qPd
efb0YnEz8J1pia587C9OmL7aIMI9a05XhsTZMEuWC5e7jGvvMqzeytUl10FRCQYM
nlkw5887Qb2koPDjI56U/TH/XxKklo48TMiqgeG4E+nyfEX1ElVjMRebcDiIRSju
ttQ2y5lsnEKLT1htw8QKET/DjgkNPTKUxdU1BAYEezqNHM0i6fT+CLtTlk+uIVaL
HxAePBCUYWvzvrLE/px1iNkuGVTuWZIFXtpuLW9MKUYJsnGF3eo9ZS9VtS+xExaH
NIIqBfILT2OrfinYpZxWYsN4IpIXjEile/KSrKWhT4tIhejfGzfsb6JaYngOaoXk
dh3pBCihCQVtt4712lePzk4rSx+eP5XQMQElBN5FH3vmG5hsCtWZnaby96iw44Xh
dQjzPlBt8i0XazZ7mumOpxtTu3EqxglJesYwxuteNrWASHbeZ0j8nl0a0rBAeNYC
1b5lGXxDOQEWRMc5C33JjGTIWdy4NDG7dO5HpK92HSEn4H2J8xwUFh7MGpDFPg29
igm0nSrSS+Dzr5MBR7MK5pG1edAhrd3AFg9uJ3yETUiosmBqEJLaLC05PgS+Mn/8
4J445ueNJl2hzLK8i1qtAX9dIv64GYrtWsnpeayGU7fLpKILR24Bm6ZuGELK5f7h
w91Ps8j6CxDJQ+Xv/jCdVsoVaLCfmKAnXzPeqD73lyTIkqISYyRnSOZVwMH0Q7Kj
h7AShjpmjubg71gCx3tvRj6Zxi4XvYZO6WgGM1bB/ddYI13Vx+lm13AM8yQOxNnA
hPO4qPgn2wBwrG/ybhiZgvOTsUpZ9XPwQFTL8m8MGa5C2wVBCKGjoWeB71jOPbWh
mcALKPDWkUdUZd8cNyJglzjq4e1awrmHYuz4XiRe5AJGc+jDCsDwmLZ8EUBV0muH
Ahkj9VDQLBLxsZvP19qX0RsKbM+x7Fj5y/H6Skf1Mxui55jXnRi5An62RG2uuAnz
JRhceAML8zKMAx9Yf3DNw4WxK6pTexzQ5yWC/+xtczQdeAVoc+W5NRO8cC+P/jCi
AVnqPWgAIes5BChxK0f9iS+YfnyHWd4cARXvN2ASrlMMq0Apg3/hefacuOBNeiPJ
wZjsQYBrk3l6GWiqDDySchYCZvSnncBJI92Dses3t3ywm6rn73hbx5pbZM7MrmB1
Xv0mE82vNpVLX0623DnQpI5gpYRCNHL7QuFKIxn1WfYEMcM/OZR4fr0K8T0j39qB
LpWsd5m2emefuHhhHWnDDIxwLzFGVEGj9+6c4WJVfH+HL77uLGtIvcKuoA2cYbla
Zsjaweam7y1oH5pr5Jy/oJOfNQ4gFljYCTDt6TIMTCNy+y2qQYQntXt1elkVnziS
GmzMqqXp+ucmaJjZqMds0wFBrmEHtDcxieCQix/BIDlRza94k5+phwoGuai37wwZ
D3IPl1vVkyYNDkk81oMBSLGSqis+vIs662Rdru2kVo/sIr90aqJosOUvCCkeZv0Z
1uHJmoZIhQJy9rW3rZXdy/69Mtnpi45xUfMUGxaB+DhlEwLSB0ul67joCT0LR/UO
1gtoMGnx8LuU+lLLa1nNJbaP9AYVzQbrwvvH6I+YJQylOwscEodOJAics09G8W22
wEqJRPq+/Ux103j/kP1BtXxaroFzojm7MQAADCr/YzPm4Y1i15CVrIaGfHAvKjGe
9Pwz4zpyyKA8HVasmZqmZxntqOOL9hbwI1Pm8E6Lomp8PqAwLjcMhjsTPkfbVDYc
8ch0EACXxd48QWew9nEQbIQCTBJ/5FeEN8jZsFnYal7SZ1w/X19oTXwfVxd8Yu6Q
zJX1YExlCgIin4BK5jTZnZB+jbMzPzqjZAo86vmzTsRLYJXg67B30TdHIUJk9edD
ho29ox4NmPe9jRTtsBYvl44rIRTbwlqqp7kwJRITX+XJ/EceeDJDIUmh+3JtLYfs
LpiAdR7F7jTHu0/YgLValpRl1FMF4bKhu2ClMf4IuwMOM+TuR0dKNwvZneJYt6ur
BDBw/rpAoQf3+n+x/txZEiLww0hdDGeOQaQRPAOlL2WyDQid50t1rt0p34dbLuec
bDYrVryFd5Hi2x1hDQbCPWR12JEFRzSr1LiSSdWWkGJo+Q/KWUMV0cM/z39xXDSP
JI3wRsc6o1Wj6gWdara35zCY3hoBqqw54BqUlix6zYRUEbfLJo9Hdg5VIm6/1xtT
N0ZVO0AqyJc02IwyoINezXRXWtMPy1YVUAHkEt/3TqJYa69MaQAhmWTjSXSGWsjh
LuAJwKYB+UEf+Ye/x+XkJ5bwIWazQfGPfBTqkoUn3wc2GXxd61XQD2KP5jgLJylR
6Ukr6RcgCixN2EehVO68Nr/KsutHqOZMJMu8ZA4UFtY9opuiB3dogYlqpPdYaBZq
etS4HzehJaiBBAy/7yFVWlzXDOvdRvNYHkm2daG3oKwPPHH/7zrKDIk5MZfNfZ23
w/4qTU1N3v+bMhaE95IMuxEiKIyJdZ6hRWQWSL7zkW/iZ8gGZzniFQtEVlNwASr1
1NuOqk/f18t7mrzDxejazuHPyqvxY1ovzUB7IXYNAPF9reqhGy8v0a9EiH9H6BSa
QJrWztiMBOh4xuQp8CYwGz0AQxCoPLCcjdSwiM9A8CPbUifV/XKzImY0+UeOk2S4
Ds3Hf5502jrGPRYJtujkRXrR2gYGTIFcXObessSGPbT7v8PkMVC7yg9jnuI2bct1
24Ua8GsUGN5ry2tciJTyI05Pmnr3L0Nn3XhgllAorigMb2FNXnAcL/Ys5KP3SJk3
idbhB6zABWZvEJxPtblLtYcz5mWP4RrhFGFhe+xqmBHFRABMet8lM8tF6LQAQUsK
jaNb5UFVHG7RfhYtkbJn/GsSoY2+BHWFUEF1FI1aSmoviUKcgCm1aFxXn1ExqIYx
UDuEGeFTlMep0bC0G2ko7nawGP+Ym60wgVRy9avca4lxko1pdWnLwBeBS2bMQNmX
q/MJl6GrMWoJG9NOTXAjGh9vu9Gl8aipGe0ITRZLlPNEuOG51kcZt6snW4fI+iF5
J7s16+JESEkKEv/Z6zcPbPMPbQG9rmDPmzDtbTfrqTrXHEcDKucXTDDSTIifCv4Y
asFTtnHTo2tNNhacCGl6fCesd1lB11a90q/9YrjGUi3EMlGS5WWoURDloy5JAoX9
D89/oVtcIPoRw++xYdI6Gd/FPM6a7aNhqWkCJhmHgeyF6U5SLN0Xs4Hfl8++BUzP
umb4lp+by0mZair6ntf6yONuwsisNVyX25mROnTLwqPJlvuKysbWPSj+ZSytM3W5
7tNqDz9uhd5T52KG+B42qHlCNDHfqYmIgNRpd3KNXe68J7l8H0Nl3drgrVKr7EE1
EZDQFavUF/3ObY4yxsIJmvC5DrLnsGTQIB432nVXl3vyZV+QMBWQAKgdmmn61zSI
9d2f9tRQWkMe9GMY7pC/lubKnqkNRCxkAOaI/KXrHq9AVnsoCT6hKpvw1jt/qlgj
919IwVGMmtmKA9nkBR6pV0s/9q+Sg9kEvJfblRfEHVka1vCA/X1rf6ScTSy+LYC+
R/qsG07reSHkvmAeCOP3++zJu6wE3RKCuHe2+F7tk3vxmlN5J/WHSxT/Ry7P1l1v
bbsaDq6YgFO7Y+WKrNCy8Yo4eoAnYa1EqWQxnQtaRE8OiDFafkabKAmaLZ4G/dW7
bHPdQ56hkWIpomAcBmuh2G7jSbZ4/GmJvk5f3ZxbfO01XfKffMe7ZLV3+iemktPJ
AJwNHZraBtjfYraS7MQFeQC3NnGk+oIT3d7dQs4mKbAeAnSGHIYXbIh+a7uoapcW
mk/o2Xk7oUcquthdFItnQDWWZA7NVe5eiV+TiOIjPzoVSTArhyqt55LrwN+lj7MR
q5jtXZzF5ygt7pnx9G8IJjLom1Vr4N6KWckGXCT9zw11iKoH+FBNyMGB0FUTcpf0
nya70wYxgJhjgDWDOhoOdx/+ZWkcg0T+BdodDPiXd5EX53amiSS4TWVUJm8jr9L+
Rc1P7pv5DP7TjHEI2Iiwu2mQBf4fmwqw+Ni/SohnAGRFVCxlp2fxelG1J1IQQH6N
mXSNdyEOkuYrvOD82YtJKv7cYZfqrH6OqLrcqgNrkut6t2SeawhCUJ/RDDOA7hu8
vnY7NKv0xdy0xvAowwWxNrMsrrjoDzx1paf+CAy4CyQeA5h1PGIhQwLKmyGt5U/X
/RP9RNAkqlkTWnpREPdqVqsXhjrhYvkQ2WVIsrdOLXF2xLkT2flVzEHyPY7Wsl/J
rBKNoTzcpVpvfkikuP6eiBsW09LMa1Evvf923iFBS1YXsL+tFcDTWVR6UCb92z7u
i0NQv04/qFQX6dueXnLt/oA4kUxzwQQB9EKtWejr2qwz3vi4cDXikOvD/D/+ZllA
57U9SMXzhx/49SxdRzeiGJtbKGi2iQSad4fUak6a4HUmIDYXrbWXI4C3iOLlJrqI
MwL2PGBf8cU/KZNZcoLlOU6AJgF40DMagedGa4/Fqks8Qy2KQi6AmZFp2Z65lhsB
x8JAyNCEM2RKxemfaqLU2WG5xR8+Idq7ZcaptnTjXxTFzS2iGvkl6j5FD4+NOA0F
jFOXNZU3mBXAKgcwQ48BNj3XMNTS/e5evhlTnURGqmhXvUsVBkjbXD3QG/hbmein
oqfiOlNE5SeYFr9Td/7LMVhoZBpUKZHS54egDOcsc7nQjyUrW9w8CCfQJ9I8AgEa
A7PnTWNeaAFOL6kOR30ElA1pzFKbtnYBhml49P0hy6yiQMgr9pz9bXFKk5aNUsu4
d3uxPFiOCYjxVyjEDUwczB/g4JctKhFyn8YPe8kJhvz794D3PlYlH5zRfeFWgZJV
QwPDKwVuJlAYHD1cgmsgRuFokFrCORBSwBTT4P+2LBqLsw1hKOfY3ZP8W9TTRbIk
yJTSSF+oollqdWSVbfNwoEF+FxXtHBbCmy9wxry8hz0SHZl2O6IaNYhEGuoU3uUW
V5VtDtWR4qtN3Idsl621XcUn1ZpwiKD0EASAYVDCqqhZIuzX++Qs1WsxJZN/FUBA
TzjwJ6I04Ej07esk1bHKZ29ivLY1IKML727FjrjsOAapagyULqseLBqJd0P+3aKd
gxC/ctTPN2M7f42BNKOeb9jgbTmKqOf44EwJp/TYt6XiCCo70kP2MS3u0NoRGaw3
boDKOBkQEztoHNnOZS4mwRilWplsaia4C+90dhnWK9ANYYaLHtI8paNZRY6+sF4i
xf3SkDiN2LhzUX4Eb71xP4LJj5uWIhUOP/RG6+JjtnAWfe2I49YW8iM0uFCFNEAn
Ih8ha6bdlKK85qYUNC+4chdKHsqxlUburDwzVMgqPEnc4kQcXwS4LXgylzzUHJTs
Lfbxw1jWIzxYXmA8+hOFXxtOtx+av0MgiHXMpsSDqx3yRo1/IETWR4s2ryQxUeHa
IlPTT1LMpWnJsrqC5eh8CCwaFGJTNVUJL8mK/pUBjYOuguaYvRojmbXI7EX3GE+U
fDx4iLt5HQUSxp74euY7uFN01XYgPCisi8vroEZsdBi3aN+Utlbks0v1rkRvT379
RzBZ9KbE4ehK6X0S5LDgRFIfEBF/mBZ4jVCQFEnImQkViRUkWoO0W/6hmLb/mhME
Fo+sFdtZ9lUHW3XWjYGv6fLxbuGM7SqzajM06pKFjGycuKd6YjSMy1/ve4U7+kZr
UDT18Vc2LLVSe6F5Q3icnxEUI8AS1HZ1eE13jVU94CzR9rZj8bES9GB+hm4+/dt2
eM84A0ZH3zOgELdQmVR5s9BvVnJ5auaajPfoSakAKH8PTookcjoQ2Qm88Loex+E/
OFtCLW2TshM9BSCPq+mCCLanZ7ZoNIgTVysvfX9+6+Va16hfS45Ff/ROpKrlHmeT
4Uzcj2Kla7jTbSwLjUazqkqFl1b1qQANUF3MJQw5Q4/2cQlrF4g6Fn4x/ZlhUTVD
NAfwcHmyKgIU+F7JjO53pmAHnQJ1hU8/wgnTRwEWWs3GVs257j2HntgfBBgJ4Gom
jQF45El24lPqf9SHjUptLJ+/LV9iu6Mvp9uua3jFmd0m+X71O09bnHsBhGHCNhAS
Z2Gzs0fisDk3IVqdcgBc1PHpZpWygwrpw/SM09zpJMQUJqehBdgR6P3DZqhJxmS3
hKDk3/T6ap//27MEPJWRwULpaYF5ndLNGapRuqyHq9eSLdZpkSlj6Jy20kplqiaE
HECP1Awz2aLVpt4dCRtp672lk5tZkUb7VUvW/c26tKaeDkPrOZqu1Aug34PMwa/0
zUbJWwfpTSMCktnkuxA+l5OMkNLBTn455PQP7RNjukIqvHGABCxn7CFqeW0M0GJg
bdxvvAkWcowOlT5JzPTEqzuJeB9ACbJBpp3kHT1HzkxQ5J8JSyXufCRmXZYeStsA
qHc9agseStssyRNg+RDhv/W+wigU/OZNSmw0jNW3uca/fcktIe7NfQpsrJg7hhFI
LtCwJn5QStPigokvoi7PCiwDbYboTiQwCLMYQRySS3k6MesS2WZCdzy0FfPUq3FP
qmsWK4CJ7f00ERfuszjavekY/wxE6xDxxpq21pEXPhlXyd8ld3GVzyPBRDHduzwf
lyTqvYzteZduwups8ZThYpGJo57GZLXp+8mw2NuuxYFlkBaBhc+HFXy3xP5C+09D
j7meis6naKJiBgnJssHPEWpKPASDqh2w21lYWUOTkR/ie6DbRd1cgBvbAGJJ2+ZE
y3jBazeQq0HCRCCLdJnnllQ3LJXu7WCT3GOHYRo3jOF9OW17muYyYODoGwAlnrOm
zMX/r4at+y784wfw2hTdLD/jcb3mFlefBqnZjO8lLe0taMS8MlGJjURsVMzO6doD
+lbhi4E/SeLoGZzTZukDR9LaRUnt4+JF8yErlWKesaIJ24O3sJBTW/zpP9cCytl0
dfWztUlgBRA12Nqggzo0IzqHCqTmajSi9aE/bmxmN0IqacEfLAlV+e+ftRJbdWLP
ukOn8lIqgM4OhjE2Z7puZgKulKM0Gwyo4Kduv3YIMyvyoAXl2Z5fmy6I4PoVZ9vL
Op2VQaPM2n2m4gcPQS/JCiU+nWX1/G8U5MR78g+y6L2eKsxgbF5elDXFiGMfF8Gi
CGMLBJbPvLc2zJYKBU4c/E52P73GesDnwJjzbAxfOkN4ewJ1n8cfseCaU41dXdMY
1qC+0CSui+llV8CXhCBlXmc7o7dbKjGPSi81aQ7+NMfj/EYbzX/DgLnbaTPGw7PO
m015A250u7CQHFig3S1dXYWJXH88fwQ8lcPE3Nma31XI5AwEnDjqKTeCg7mjCJy4
Fma7SdioyAqKErY50v2zKNW9sJJDUNh5uqytUkvtIvlzMf+fzIYouCJ/rYLXKk7w
zgd4kOY053ddMh74AA3e8h1+bxWlcRjvmL5Et4xJ0cnoE4bGhBokqi6md51i02mz
Nt6ivRJ6F1dKiT2nLPmQIOteIJbU6hlVEeh2+upiTh4WBqafGadx5jgUc0LBvD+R
Zgp2bEFzh+GxUlrbCrfYMF/6OOTu2HUnNoR1IZnhmEYUfBxnvOBUqEha87fNCFr+
E7IK5+ksoeK0iyv2LpNo6kS4+tcAv4JRy074YRjpRhCLetrvo4VHMJoRNj6W8Sp8
LdDwaM/TCRIU0pAvhPwvHDRZ2AKMS3YGqjUL9ygdCA+zAh/Kd33wBHO3f0FtQu7Y
b0gvOxCyaBZa9ZbZV3qtn8ghXFvE0g5/9Wlv4dIW55T9udUR6sPUuu1kbeJknQj9
12bPmOVRYO4cAS/BOJL5RhEaOoImYOuODKI9sY15txZoQm9y2SupI2rqMGZszR8L
8qXAMY4na1ETCfdDVK60H3ZHcmNDKSg3eUTa8v2MubQOp+gi65A74565ohSTBzmR
HE+XTj34vGpiQJuOz0+k4gS9NtmaviPJOlIvL9a72ehvFDX9Xxfx4diE/bLnwnJy
z1W/f59+1WPhH3zkPTfpP4ajuu05zZ9gSc9CjV7TkIOfTcXuGlkM89fn1EfCbHDp
r00wl6tS/Yo5aiCvUtxvA3Ia8fQKYMGp1CGDYv72MvaY2ZixjmljLJruFCB2dIvP
kGFEKTY+2W1MYHA4H99MT68C1t3PKE0zvZXrVb8I9SmZYEwO5NZsAQ6QnOylpwiF
zg9137t2QwPhNLjjKRyZLdggdTIcH3DwlUFYNgJEX+pJxMDizGg+O4eunnflXJ+a
0lzlH6xN4uEmip2SvsnA4lUa5dJ3xme75y29o82x6Z4Ln0qcDWCO/+27wJ5QRX2V
S42mhsqV9YBbtpzpPOc8X8XFVoo+JNI2nJd3I2tGnwPCDP/V6rjSclIUuSimxPY8
XuKTCSvuObXk5O3Yf65RHqco+Qtmx70HjqhOrcM5DljJThOKqlL95CkYtDo85E6B
loMDjGdPwU6dSv2Id7paRY/3RnmJCNJenaHtCtwEwblCvcBNy6d27ufCjZwAidaV
PljVm7wS9pwloGdUnMmkb4GXkV/OFt3zrXHK0dX4D1c8dEVzFZvu6IzAf5DFi55n
8G7HLhQH5h+uVeDnMHkyRThzD8ClTDBk+V73f/ytTvy6g8/F3jrAwV+vYLZEg9GR
cTW3KaePm9PqsGlc60B3GTfA3D5dTLinjc/SRCr4yYGFnGxgNJbTKZU9c7JtoKwn
dQ+4ct3qezKihXbQEmkjfwmpY5bm72Qk2KkUj0dR9WXJ5RGEGd7gK3XrTtZUQrd1
8lrZpfshSoEIUF3xcSLRBwlWxvm5J/sk4s3k/Y6iz5yoIkM2SUx9ZuuAipLd8wWT
CbPAHCZ9AnhnlIWp//lgi/+In49LrazSLI4wTpQGBINuPUggi2QBvPh5DGq4jM5W
vDLMOoeMyXgb+Y4UidVugSzWW5ihyHiEQLFmhw1w7wDTYYAAASNF253lcYFUsGn0
QyKWzM4pgdfbOk+vjD9ykGyFiWYzmu8ZiVRLsZmYOo2ZE2KvYaCmpW+aw9FNfF8b
reRj2vRNWmQ2dRPzqzDGXsooScHhrB+es7v2FCaPvc+vrRU4wTcRq/50lpuI+bin
AsM5yjR2TJnQrrsMpfwQaFcqErk7Q7t0gU15fDYL2b2jbWFM+01OKdRps34gx+av
KypMmVyKbH3sdA/Ma6GX/CKWJ9FRsKhP0birP4ocD8sX72DJUWvR3VDxia1loulY
RNlO7ioZE5qEM6dXoDKnQgniypYw7359tJ9YncRH3jxveA0+HMo/BF+4EUUSYdN5
iaQXLUNxVf/PmvRQTOxfIHSATmF8q3EqbKsegGad2AS2Qesm5jpXiY7aIbxgmGjj
vzWtijgXkuiR+eZzabIbVGp5xBPLp1UfOX99bbdAPiYS0cD3Cja43ck5OJublFOk
RxIXwWBpsFaCa0BP1gu3FSTPZPAL7eGwbdcZonaWMB8cDTZsgbhL6uj1rlRp79HZ
850sjOBfn5XeOFN8+VLIb2YwZYu7lDo8tF240+LoFF7IF0qvg/Si+zQS5n7t3lX3
aCAxf3NCtmWfStEZ5lm3LTKnnukwOQWfAyn+9FTB2yqjkKrNFC01TnNL0/Ch3xcI
rxtO1kcl2AE8KnEVR/24Zrn9xsE6Fa/V1qtQXXI/M+Ql0mUbJ8FMbcJXkQBtzFXs
HI33KgqinqLomWm/jeoDN57FOh/SS4/2UDEsN/EwiomZvJrrVcpEQG2FggYBNMlA
Y/1OmJAoWV9WNkFluUbmSUGMjUhk0M+Yhlv0kR6oDNSuNtgqAoWcFLXltNsoV1/R
dRE6pOlyDEXtUSozqnaf3603ew3Z6ZXBIzxadMU80wJ6tAyHa7dWqaOaeHnoIPtB
BXgMvhsrLCdJ2qaeikaBgpShtcYTOu2d/P//N1MoRpv5hSHyU0TohZMnDQOD8gwZ
CPIOzc5ipMK1cvLBr/WRMJAf9fyv8mttT3WAXJ4p0v42IN+CTRT5dB0IDFaItW1x
ptVBM1FB0QrPyRt5/FaQ79ObP3rRi0ZUjQgpsZedYp+G/VXGFtJqb6RAE2dJP5Oh
uw18yZxn1b2u1gcpz+r2HCvUKhZWbCGnbYRoiMCoRpS4C0RlMSXnfb03mQ1fC+VX
ms3N7x50ahGu3PHNG43nzTh/9Ztg3fbSPQSkmPgKiMs5j9Kd41Hh4G4Nm3F79015
6706ocC1OoH4hKAtbK3NqS74OIOS7iGJgyiQ264O0wqU/ObK7iSmrAga8BwXNqCn
vmKK9MI5l+n4InBPpqryAaZYi6a31hAVhTh3b8oMA2q+kbJ6Czawk1xJw4DRs3Wf
wfzef8b5c9Ewm6RSUqgFMjlt4E3chOqtY6YemtuRKIGm3copC7Npwr2ptVc3TDXz
LoWDZYPDOZ3FwhTp4d68Ko/aH8B/WgakbnL8sacU5k00cS9LHLG2g6/Dhjis8Xjt
bIqwqAZ3B0uI7Dy12iGuxdNOd4qA5bWokGs6EHPPYUZBr9tENuv5zKx5SUbxpbd4
x9uuDP4Wxdjb5F8s+toFstKkwvZgoi8ECx5BqKJvrJMKVSfh7KwhqTeTqUl+RdgH
wmljVcT7+9LOgZoY1LAp18lWjG0vfUOFg04Vcjfd0Uweknm95a6r8j9NkJr/9wLe
Pf3WQEDwIoWbtREJ662ShSp+LPM+3AxhOMFrj/b6iIMgMey11MhlF8rrOpyP5mnv
X76wyhC/01XIZBny4JoBy+KQ39via/VsAxPGnEK16zSGG7YRdUKgnrbw3o0AQl6/
UhM2d6q3ysj9B4H+DBaGE0+XUtmBSTw1mOwVRGW0BxhTf7FDLCO3q5QOxqFVhcLr
G1f6jxCLBQy+uqo6h2v21tIEHgjD3MZ0nEWxu6UPB+WuuUrWMXbaDojoeJXd80ey
P70wIIFkeFo4pZCZd4nkgynQJMIz/vcfcOI8bQb2KNDgMXFK4w28vcUvba/1tAt2
BZbdLa4tIGF6EZkMdYweRSbGY4N9yBCy4oChkVPvLWYdHuiKmP6zcbVunCXoGHfp
GhX1tpODQL3UwzXEgh30U7VUXW3YKi52Hk1tsAt6QH1rbq5yJ0Jju3Rwmj/cXvO/
Ucddz4SFYYHe/lkF4GpCzzZ64u0Iwal3uD3wVH5cL+6Z3ik2Fvry5Dz2WbNpw01w
TrwSjd5Tcpin3L0b7mWEwSXlnVaLaeVm1D3sWKrDo5qZMVqAcVG6u4buHVa0WHeI
2n/iWoSxawPch6S5CwfiW/xQkO/m+h45JeRuptVtYuXDXRsXCZyG00jz3WGWXXcQ
tZflM+DYDb4ORiEXKpm/Zo3rrL8fsuGPSqq5TSRxMyOn5edw4mVnxymWNI8jYWZ7
8uBmPO+Ev1A42nmcuvluGPSN6nbHz8HZoMwxx9dI6/QymiG5j5cOITnLi8Ep1GHR
T0IBnk/8fmq6HwxONrJ2L77OBHCyNDGdF/r0/VeDHHndUL5rGFTLBa7MLNfebO0k
y8TBfDV1RN2/mj0yBGYEUAd/ETeDY3nkuAac8N0SxY3aiRAOEEwlJA/JS7Y4FeG7
dfJZ8pMDAVRVbj7oAJuZBc//4OztePMmEBCwSoIIis77b7b5MGX6JMAUiQrXmml+
pj5vS6SLnOcnDuHV5JgdM7m3xObwH8o0Mkced9oT+R7cTNe8TzJ5afWfaLM+6s6p
9AKfjzr60QMyQGq/RHlZI4vqeDNi9U++RT77kl2umlzntsGSWGNexvc9y9JFkDpx
1rExvzsPEInf8f7Vec0pScSkrtYIlRFPCjHy9orOQhzh2uC0R3Y84suz3ncEmD73
O1UsdiOkhU2lwia2j/M3EexdLmiB6WgK48ynA5CPE8dZtl3zB51ditaFeeiYl4E5
LB3a+g7wSJqniw990o5FoYOdbb8kGgWL0lmnc/xsLDkkBB6dWZVDyRjcwo6Fc7b6
8QL9sBI1rBjhD/pPrXjBvG9LqmXeBhZ8EHfpFaRgWNbb/5YsA+p0PQNQDtyZv/Ah
9Ymm9JQzyZXm9x1ZsbIq96KVQVVk6n08q9fSvqKgSKuSy692IilUgUanbGv11Yxe
ocMVMLyaoch84JN4U9X0ndCN1SgEboLQQfKJOXG5fg5tzSYyAcQkFdhKgF7H75uV
DRidu6hqJQ+q5QQQLvWuAVwbiVAaCKGZc8Q+X+p0zvuuy9h2CNZRKQQz+eAmVz6B
1Jt4/sYw/KkD6QqzEAkaHCaUw43qDI3LFiUih9zq2rW+O5Dl60NVF4i5wznurgG7
YS2Zp89BmcwMm5/2fi+mYg3Ep1vZ3zyU4GgciipoyM/hhetv4MYdYHk559VczEzB
mI2uFLgx35aFpFFdFuB+HcN6NokREgOpYcz4tZSPTaKZZAMAqnxXOhhpGvFfSbxb
A2blNyLbbXpqnEyymOXD62SMPMwN5UCRiHyr46ynY7KyDeJ+Pwd48ALgk1upMmbv
V3N/uuuabzn8xsqZOmGRgrbzgOhNomPcBhVfJUAaYjL39YLLH20C02ohbFc5qKX6
rTzDLv4lXN8RPE1PkkDil3Jaa2XgdA3aODSR9hseU0WGpA2cOIf/X/vEjKotks4V
YgIdvb3wOh/3gBDxMOKLSVhBMD4d32Ykbh438wnNvFwkJ8GP+iNqwmKeWak0vRv0
vBh8ej/jj27k/vmJorTMC3hCEPCd099QLoYlDwfxWiMTAjfPNGoD+kqzy268uQGj
ZpxPJ6WXIpCqX9FWQ3E/EYldJJNWeF/UHtWLXCuP7iMiK94TiDqvm45XuHAIeO7C
2XNe9AGhxlMh/nwTEZZ4BlEoGIn5X+L1IiqJtO9cXaveKhw1aSy8CRJlDIxNHzBB
fhTBzlZHxLjmURqUMzt2BCSVvUTBXwWZgxoMKYpeIO3On0VH4tokTR4zWa8Vudbd
W+WgmTEhKb/mkz9e0eKsMW/2vDJPQornYItN1E4MldrX8yT+B5KEvhmicyyfjy4C
53aNUkLzwCet7ctUuRuJ/5AP4py6M7EMFW2+SfJ3YWjllh4eN64i6ww3KQT78/Gd
dgXvLDHwVMxHpr4eNonul2fGpTO03TBGs10gdq+gHH1Mivb/VCGoY7rSJq2o2P7T
pIu6NWfJJAB2ghZBeNBI5WsLlBO06TIbeXkx0r+8QxgdxlYKlTDfd7fAXwjldXVB
x0LsheVwZz75Hcj6gq1LWy5VRMc5gYVRarbsZ1ZCDf+cpjDn2/rcFWPCnb/E7qUB
96vAs0VJBosDwN9/+yyLBgQQXVsPnBIOfgwTPwRH+HsD6q6tYqXE/lXpDjB87ybV
uAAwT11x5nxjIVYaJCnGEYbWOnrmw08V+uNqgSNUO9WTOzHhD49EUJGyZ1R5lxvH
YxrP9TSNBmMcY8an2LaVxHgQhPTlEPbETlnl5kZoat1F+FNsBiIqPdeg1CJwABKy
+zlQ0OsU6T7aEZLSCdXvNIBfPY/6NI06HLteOF1cE9/M87PZY9J1VfEWiuroXUsN
6PtbA6BQkBsF6ITZUr9JlHI2sFeANeVHSGLTMCP3g1rGdyPggtZUOA/G/oK07B7G
gZ8jd5Bnj5nQlg0mvnzxS1MRT60FKTF+QeP+v//cCLbDO/v6ZnB3Kh0Giz0lcRyo
Wql1AwCBzIAgo3LFhjzlpEba0gm4T1378VqAuiXQ3lBlcKOX11W8JZEhjael8Idc
8hdhgREYXoxXcwzgKKp+vQU6TFpH14yFGYNCz3nzcPPw28QSjQwRfvcDm5Z8iWAR
CwZO/XVV+U08pxlUgIJxfVoNUgvPIA9qlkIxycIhoeh+ICM0cyj1QaPqFZWv6VCv
ZC9fds7SUtXHLVyLWgd/E1JD+lqlj0tiev5cYtUPwcfiqA8gz6WT2+M1KJ84hUfG
vI7ONpRlHqXn8KnQ3Ghd+Cv0db4dimzlZTHXLctmRChu+SybXSNEJbJptGNpM2Sy
A/9J9bTqm0HNVuUWGSzr9bHh4FkpYODTfObJNtrhXYciizpbfP1ukx/ZqrEczKVw
x8hMQeEXAn8YyeoIUstw9oH96DUM2plGwkgL8fgNL5Bz7z+IlJ5kM8NoJXWh0dNe
fm+ghKKhlPcP77XTvbkyb2y73ZfxceJ7xiRZPQe4o5k8KTbOsNTEO+zGaoqE/htt
mzEt8lTwj/qQARFKmIAQDoNQWadOQzpUw7bHUqxwWrcQGN6w9au3jS+dFeDpCBl8
RbhUncr9attah/K82t2TyxG+/VNifYjHeP0gBPkxFMOh6e45tU2d6Jc+wJNTmnqw
4DBylZvcX/9aIrdhszyUyfQ4xoS7HNNYNAkgtktefqOyDy6WomRmalgYP1WiXhsh
SGlZvnM8nQnq0jzzIkKsz5jcvf7eVU1Q/EfLmLXKuv9sbVxPVeTzz1x1bqdD3NDu
mmKi1IMaX7f0b+CpLYh5oS91ftBD5ga4WPhJpBNwha9HcXbF5a6WVj2Mi4Z/0Ant
yr5ZdTFZLJuyp07Hbxd6DkKMHEd24hVDRuD0fIL8dXMqFFAVd0iGkEmTWyHquCUR
LylBdtHaZwvBLOgmPE+Uj9qkjlSpX8GDVRUq87v0MfOQRtNFbWSBCFyQ01VLb3CM
LjVLyD/Megtx/an/Gvc//PmfOdz7SPFHYPz0hsVkHj/TmJlIoUrHmJm1M7UhuLYQ
TpkLClCKVpd58419TMHVU2G6RssZorOoZ9PAL1AL/b8zUoqUh3i43eeMiV+xO2Xy
/F/7W8x0IvJhls9VZ6LjquznPyIpTsx2CQNvzOhjOYnTp8VdOB91Bxrx8ydZNPBe
HuhvFhmiIKZSi9SJAr0e3PpggXGQjn9TkbOUzFxF2aR2PP1tCpcF5lm6S7m1He+V
WkEXef6OBJ8IodXdPFl5BNnLeApEwZ695Ps7fXGZPxw46eYJ30XJc3mvDuWXgLkn
jKkinrCgqquceKaSOvzVs+mzsnLY0vSK1x0xYKYPQ1F2z2NyEQJ4GCG5+B35NCHO
hRHK3WHt96YjTEEvTyVqGqVeJ6xhpk4YNGIohrD+wSu3LHhFEeQ/dWh7ZjmU5cK3
TL7XVxZv4CA68KecSUtArfVTq4OsZN3j1LQAm4Y//7BnGhJxacgDPiOIn3HEYKcA
K+gPzG+WUgFOCBBJ+pPGIpYO9nFdbH4b35hl4g5KoS9FoIcVR0YQyRyn+Yh7C+f9
N5KnJ6prLdVlVYHsUeu5sRymf1bkSKMgITGRRjQNf37Lq943L535YHn03CtLsB7u
1wISK3u0m+wAvsaORCDELP1Ti0Gzr54oxAZKjZbEwAaKvT0TryIqElYOwY6cvaZo
v/VNJ3xzvk47JGmuYpjs9QQJHJePMZKZk3JeA24AegE3Rjme0vpc7/6GUhGtCFp8
YZ1PEb/n4BJs2/v3dH+75laRZrFxHJhL3q0WKSXReFrL09lsvD55n5/cjcu6kzU0
1ej29TLmHav+kMia0mPwvR9JQJ+VGUrR+sGpZmbIoVnh1OUmD/7yuAns7ShbxJpM
vKSV4FFgyULkRHhgv+YeKEebG1yBSD/TJLFSnSdds7/vAezJFffLrrW5YopoDvG4
eysayLw1IM3Oam4nOCXU5aDrD2AbtbDg2ddCBV2PA/FD1OhdhKQbJw7kkCZShut+
WdDBacF/KAONleAemmEdVT9Jo6l1xSSD5qjIs1FB32moOWPfdN6TR8yp2uFFAV2t
EuEr8BEqfw9fbA6jxRFTHWiBfajg/miLI9J0OEMugJI+jEJ2ClW5Rt1pmGU8QC2b
7UNg8b5Rbls/Gr2hLyBE6/i8+o4w73EjKD6qCQi4XrQ+2rwXqCGIZ6VuhHIOCe6t
M3qxyN2pFhwN37C5k6eR4nsjlPo0urdKdDjPRS6xX4c3Uy45U0J1RxgEaws/T0PM
FMsDJ+/SM9pQx1YSoLvJn2aa9eppMvptZvlhhiY8XnonAwUQ1BI1r8ep+MLKzUoK
GHkqXKdqaHGQcJI7FkpjqKBwbdVumeCiZzEDYVGHWYuBIm2Nbb2gcSwZMLoAFClP
2kh+bkUWdIZzqjH35AaZavZ9ieFXCM8nQdcGONgj1QuoITpZTc7ZPcXHht0vb7NK
iwBtAIl7a38ygXj8ijK//SQFxloVUZQeF76YGNCF5e9KfG3A/66PNYO3N/vrK2Pe
cBgTQDNQeHNbLp7DVoOKEIz+OsZvuqbLg0agE45jvYSa1HFGAK8bxNuiQxQJrLEG
FGEPWBmqLGpbSkGxIexanXWn1NWgm1zTJUM+pSknia2wF4YPEzgq8pilWpYMFfOt
FXZCHwntJmXe13kCIVzfYVPNp5Ce88fW8gyn1AdMPAYgCZwymhtaGEGsCb8JtWUd
oFr22vdFVKjXkiwWmuYnjBjrj+PNsn6KnfZkE6qpjQQUCN2voYD3cb6Pr6L1Wh+9
l5sYOoeVUqExgZk29TQYTeB8Byeby/Ypk3ZFC7LjX9MYbh6z1x59naxxgDEyWCdk
KTO8osmidPuuATGXZn/f+A+KZGbUz7TvNK+ZuI1pOThSRp2s5hb2+ReJbBIlbQ1f
fHTZxG2dCgO7x+IvKGXfvxGkXWcYFK35KGuVKwUawTHehESu4yU2KaFq1Fwbu6VR
OaC6seB5FGxorNypegdLEq37Yyntgy/w3g1Uaq8aGkEMDJwijpNRUlG5/x1bj8VO
+/dfHLjUF8BGPIorHi4saZPGMliEgqzg60keVt5NtXpbfFE0RkW1BZhmdUUBKMvt
8a+POybaT3cNkqBeyjtng5xdfKp7NxM4TBNzjra5iCrL1tcfo79Pk96NxF5byqpq
vd8ZboRoiz4+a+Q3zUdl4a+j1de3Fef4NBMnz+5lhKBhgO6E7UNVNxArGbhlaqBV
iCx7OFZyNjhnTvOYbgZDBa2beUQQMMdrUD5ocCqA66BOIeFjmYGptEMo35KMv9oO
go+VXVxEakqZhbi0Kuy/GG0LZnbbCzegRXS7dVJU4fMgx0naD3arBg8A4B8f4iep
qR54nL34ythfTOHARepgRkMH18gzIQOt0rnachRvEo9JRN9wfJYP1xHUZJdPwYUS
woNp/r4O1kNrwaBabJ9D6EmXDoSOUUJuEaK0wtBDbRV3NgsZIyEMHM8tlsSe+gRE
v+H2uAYmopRKybbH2AlROonl7d/O/e4iRMmWdcuThJ2tQbgRZH/dt/F9gv9bHzBJ
7srTp39R5aB+biEbmpIlU3cVdBmJSTAFh+JsLWGL1zFTYymRX0zJcqaRJREr83O9
RxvrxmGs4KFHMlQcWfj/zmQJuW51eFBgMTIoF1ArdnuUd/eRB9GMqqvoDIJStVrd
uwBIGqDqw1ByeHURulz4tw7Tx5PwLsAzb3I5rSkPqxTY+j4Hv/baqELqUglGoQWR
M4AYXkzVj1sF7EirvE4YgMT9VNn96Eu7NT8LanAOqWhpqDH+nOG8fO9HrZWAsle9
bIWkzfJQbTk52zd1XwBR6AvwxkO7l/VhPSGvHOurqQHddTnGTdKHF/j7m1Y1K1PU
ct6Pw5QKrww7By9joxWDzre8CBNTa7e2CJaZWGi7YgTgdbrPHdr2gacRFRD7RBcr
q4vzV3vOrbObD2uT0KTDCHyQxUd4/yM1FM4IwUk/HnSKeLrmJPByL5f2m/CJ2ygJ
GLqGEAsBRHBQwvC3mHeZKFwIRa7es6go0G3jQ7vATOhcxoz7/ycpUQS72rPcTyEx
5EqD4a9YyUfgM2jKVXrCb6zkY7qrN5bYDkDi+E3x0cCCFNZvpy2tKpKQHfCqMI4q
S885Xn/uN3f3k7+lop5ejFRboW4mFcaS2FLWpUjWwOTtnhYi+U4eGvnwlZ5ECMLt
Jq0KRPn8TlZ4cetNcZYRwbApyXflHGfdRebugNxfJs4s5Xgtw5c+gsJINtp2T9Va
ralVl18Oyp5l7we7E+icvIrwOQ4sxhePOj/JxLB1KeqrTqhYDbqrvxj9QKGAX1Yg
njv+Xz+Mn4GTolkS+y6GTiK2RWUYQmKxg/Zr55tOVYs2XQzYTGXakchE5VBvDCml
Rfw4UhwPaWdwZTEoYMo8lJ2fINdG61D1YTB8w6n1x25Cl6MnU7SYHZ0ly/s4YgHJ
JrYuxC3W3Z6r9zz90Dp2XYKhQT125JQ7e55t+B/jx++30mc9NhgmIhsNdyvsT924
x7VA5n6cx94N7xgh0UZ2T/DhqJyyFCzTjfZwX9shUhF+kgeFQOO/WIasjaG020tW
euP2J2mxy55lS7b/2cG2aIlVAhDN2toXLRgiQdLI7lqHzZUfUQ7PnWO7lrsYR1BC
dB3tzRoVZQ1LnSavIR2C1l5m2ZHK4/Pow9Bhv0zBkFYXOdCaLatPs3kLUZH/fUfl
+516V+UTkHtXVT95HCYj79ur7DfVQvN7xupJsQXJ1FRw6CsOR43tqQXQr33mUwPf
k+MAluo8jm1155kQKsmrC5h0dwQfwV6jWhn2JjcTYPQIBr5Wla7wfUlaQnGaXlgL
PR84NQ7o83c57VCSxWZ6YG2xKasnpeuB/1AMprIz7hi7S5S/YpvwZCzS1+0M7qqT
M++4Q4NrTID0AOlvmMT7+Inst/CXpVusJ/VUw9h7osJ2ur9p72Yk9A3c2TO7TuFU
rrKBy07E05Oe0CIFCqRy3ea8X9+fJqxsdLkfPhxORpC4crbqXedlk8wHrHtmV+Bw
cTgeAY095dy3t4A3zOZj3iMUH4E8hzT5u2VvmAeKEdo/Uw7/w9D6J0DIt1y7fmq9
sqRo+XoKpuUQzTWW4SzGXIwQ7h9DsQGC1cUUQzZXDyzhB+oA1niZeVygVAnxidve
QBjULj7wLyKi94qz60rjnrQvfJ5/r0cuwpgyy6pOxvNF/xAyiRlKzfBxIp1XatTl
3e6/mwQ0yqQxoMrUMiI9coMrAxqcbkWC/tXPhkbtGSfCo5ohT/n+7Xu8uBxwtQqd
1S7VWGLWUgMp8KoyL4KY2AUzWbBiywEhaEF5APQZKO6HUAfw87h+2Q9OfnBNxn/m
O4kCJAvN4xI2BuQD5+RWKSSXtxfzZXxGjMmYmBFzOV6tH6dZxmb9x1cQHRijUjh9
D7FElwHRr8Odtpvh7jl7g6sDAeEAyF3rOzaAkkiZggxR5K0viqi7j9t++lj1fKTc
x5kGmW6o9u/T809Xp9SKNiR9dVU9QK2QnCmaMq3jO91pz++0CO97zGM9XVwu4Ly2
YKwnkpyHDRBpcUh0y/KJ310+e01S1w2onVG/Sk/gvVsCK+m7eg7w/YLUZNsrc68Z
AQ+XTO+qGCUvRFj1302Ri4DF+D2NV3eILS0JuRv/G4agt4v1L8tKjNvHVYJ1rH+p
4VZNwPA3eB1CQFNvvjzgIADe8EJy715fsERnjR/K7ujTBAWlolSi4C5CblycJV46
oIEllrhoZL2KUmG282p/Uv/0qssMBDJS4UtE5oAKR5vA5L2abKbTRb2Zxyn/MhLJ
EpSB3Ab4aiUl96wgGjLkplWi8B6J6HlX/xpvRTZEhJcyPRWzRqb7sOgL60TnsF9q
Cqi/SIiX3ZeRftZorXOau7YfuFkAqCZjwf84dsykt8Zw2r0uWokH3Jx/azbDScUn
RrAupt52QfhAaIQzfwmZmgk3O+DVYWba9mLc4e0zNGPKrgSz1zImvOcuh4vODIod
AaCMjCdurBqayXpGkOh/Yb5urJIzaO7qvF5XfuAKPmngbu2XdDfn3rs1t+WNf0YQ
+ppHlh0elGJeP783bw6eoNvnqa+lOKdRbvsLb386cLNKvoEH735dkcv4ahGLE0H5
ISgx1NuA2H13dOO47PJ5GMDtf+IeYNX9lz8llXYvJ0thFR5uBGsbA6zxwUgUxoo/
QavLGdIq1tnu5RQoREnoqoXRraOq9aprLGQGbXUqfvM2GYR2zy/20RYM9jwzKEvz
tKWQdnIDzpzcDwR1vCZ+KxBhgQOGDT47WfI2MxbR1IwktYXk44ydr1yJVEJqO4Rt
l4LJJb/XzA+LM67kg2ede7iUsbTQSo+K9e/l8X+mY9zgVZCWPWL/L/zS4dCqPJbC
2UDXUoes5S5O5mHxLa9+3JFYrRIqSTNRSGp0Z7y5OWVXaYmMen7Z8VeUf2F4Z348
9C9ZSEpj2PwpWL3KuTv6RI/l7gkZF9rHblnWV7X8S1VKRfas0txY2935Xq/SsFVb
CRq8gONrBrw5mBdVEBgDTsuLfPrKf4DPaDIpNchjTL12YJzlICc7bidY/vrqzbBy
MSapM7Y1OwBpJMVIW9M1iN87/zFNcCCHGSV+rWrXo5cBe7zJxAQTvYnds/zVBjMD
4NvNV+SlwpIChtmu+I2sTJ87RSycURsZgcOE3LX+rFoFwjUOFrzZbBNVXZ17JDof
Jkbo5XC01y/bbRMDYsQqJv2sPf/IXuxRzGi5cZLcZJGjxbvAaBsLtJ0dvYY0anjV
IEB8dprzZioGDM6JNYB7sllkSXvvntKwwbC1Ia7fa8mu3Z6oILgpozTTNKz7a5qR
LdvLy42kOe2EQpCpNwl53MPwFYhiW6P4fAEjUBelf2HQlSwNQanTKP74pnpYSw3w
TDsYucnBI67LGsxS6o3wYhAHLCYoaibYxgzEN+E510g50TKlRh89U2Yxdk10eKYS
zgDVdgSVNXt0T5ZZn4JxQyHFLwtLw5D8n7Hen/nBVc6wQPElq2EA7ycL5hD+dx4s
P7V/PJwbwOkWGEOVLtFyxjBLO4B0eNmzS9/VpkxOvp0dNx+gTV8QOXIDHCMzQF0k
NTWQ0BXKk/IfjcsNrBdHHUI+mFCIvVkAJZcl9RKwz1+SUQk0pP182lOUTcq3x7u+
EmD3udyCVoPyo7PtPAMLOhQcWPIYqW7GEcJheTV6C0bu77YjQ4WcPMK/zM98cdkK
zzylo5ULycuBGCIM9J95OtGD72j6tSywPPOjwAgGIefrrZpk9FrqZrkfTUJpaPWl
jBf3TOagjzEeoJZ23G/jF47PafflAs+R6+/xfkPxtOOdCwFzG7fS4/+f5RqIGrL1
ifeWS9D/31jSWQ75ojD57hOZ8TC5FjdZiXLBBRtJkw6ab1/EsBnuxAEX92hPMT+7
H6W9JUAZEp9G7+SKCRXLfTlWhadOQrDndOql1qYl2qoq25MRpOl7ksc+lfrLn++a
zaviITmbYR1j+3fGXKxIdX+2ITJWlANv1hcMKZ0go/4MPrYHyzTj0L64WSKiPnOp
KfsL+jnr5kdtOyAddTnVenBj3Ed7unRnmW34blsBSojhbac+W/khhTnvtOvY5Tp8
/ZQ47Aahtbuu2wS4lt8zQUKFUl3aqRA7kRfhAqSNVjmG0pFVmBZbraIux/SvO5Cb
tiBl94prttS9ogiRaPklf2wX4py+cVR/huAXk1kD23GnyT6DWcVnsLInwcstg+CN
pcIYl2oG4W9Ept2vZXLh6+1UrUj2sRINrrTTzjh2cA98BbVz2fkyB+M1OgdN/ePg
kejxDacxiiAORfYAlzo/Azh40fQSOiYB9OAKSl65bvAjsvxUlGpdEq+nhndpamDU
fZWaWliCDzVwpjBCEU7APpU/AcOJkZXA7XcYdPurOPJ1l8nf1exCRchFexk9eO3T
Z5oGWVpu00dEsp3OHP4mvh0tG3sHM+ScEGji6fNGOlgIvDHpvnVNCgHhAkIrUPcc
DFYsAk7Y1I9Hiw1rn1LQJX3KIhZwRmyiot4bH+kninQzur+kUbYNP8pIxLWm0Vpb
x8e1HluQGAFRrdBArksEe3nWRSTJEXkYLifC/549a9Zz0KnjqQ+fv4AXUXojf8rm
rBhjgUr3btbwNJ42OSwtoERIhsfkj7ugUDSnhVb7Hqss/E+WDrWlZ/0dp/Xb1pxe
gdXD1vhRkZTnqXd2lzRftp83gTifLHhNKVdQ6YS33+1NPDUWT4fBZymVkMKcw86h
qwab7U+ALYZfS7hyjhWqw0REUaXQLvodR8q4Fh2o6CIqqvLJteGLwAKvXtDGo1sq
Bt3LzYJSy+sYJmG9YYPw5Q/8tVcdOX47Eqwsf67jtYDCFCtgzhkpCEgVOuFQOQdJ
Y8rsXvpANiNyhJqzT4XV64ZjLyCqHzW0KMivSX7ol5+jhGMNb89PBgklv6srYkHy
bOXJqGwocvt2tCuRh1IB75adLmdJaxshjzGugoSyB7qtKzomyLS4bx1IurWeht+7
mgPQWd12qdr/K6z/Pz0Kt7HJUZV6BQg6KnlyoHLhMv4Lj7do0GcG9vnWjU7oV36+
A44E92Dtu/54/D5C3h21Qi/953BFmt2R0/Lpywj26qPX2YKamrAEG52VA1FjEgim
V1e7MSIZJYGqonGKOZt+l34EZjSJEPZpB7v0iv2gklaTmi/ttZ2U9DcCdO7ajfPj
uSNPkCDl/809Hb2MphDUuHwlxqKfa7HZapl3gD/FUWxp2llZfn4gaTXiEsTxwKMY
Ha1yXXMGg0ZgOmo+6pMKPlYbJmcjBEISM8PjCa5dfBwu6uO/pNT5vXGWPGL8VLpV
Mi4kjt8r04PSxLQGXAsMJFdcfAfks2QIcl6sD12G8ea6aY8ZuhVn6HlRFwZ5Kf3A
R2nb+lmwdwgsWWXmPmXskkZOLTsmHLcoEtg+gYVkHC4ExOcuNt450G3jWc3xP0az
C2lRxFHysY1v2UTILfxHTtkj0hcbjtnUNvKhgym0xp5wfUq7zkWqgXnBmKXnvvPW
Lxc6Ymt/So/pi5B3VeFWpNRpKnVUfJQ+e++7AeSr4Buco5sjhU+m3MYZzKIKO6Oo
olby06FqUYhjfDPUBUfznQ5APeTAZhZ+HiLrmM0oBjOatyABlpNqlHZELMFQtE7o
Bjf9YH85CyP1MrnLFUOTNIeEaeqtGgvhrpsLbo52V8ziqxlzdGYnUakU/J0uXEyX
N4K9lZSlncSuodieizoAI0SwGm7F7vHyt/sMxyL0SqN9jegthBEtM0GgkBkXnjd4
qTAXzsMvsK+Y877fxwrYc+Q/TK/9+XyiYWPoRWTkbu8hpNZfT0zO2VvkeeRu5rmk
jiGcq0X4rlZ/il1TChfTaKT+XuISytXnYdrGI0XrjFfwOSxjZelbixdunKUwA4VV
3qqME90GMbzY8pVRruKvgj+dDesXo+L5gAuEG8A61BIeWB5gjHJV7MCTuo8h+ddl
8MIK2gwU/LZt1Dn1K0ZIKd0Uwb/HXvNgQLS7XHp0xTimMCrRCljSEo7jXrxIQSJH
6Pfrq/cYIBnOUH6nLhSUmn42r5W4gYVycLp/nUZwQRGtQcO7RWBGapOV6oYXwgjY
mMuXjrohsp3PZ3xVA4+qqIw4Ywa9dH+N52S3aHVr5jVgdfsZVsN/wH9N7m1v5PFt
ihOFzJZfU8fnpBMZZDqHopE6pSTGSPYluko5Gb/NZUtqQOv2XWgjWNxOFP9oTIA3
V3GxLpcoLbmNqR7nXb+jcuaOq201hkiIG34/1sFb6wW+zGIS4M0mWmWlhxAKA/1k
+1s9qQOCFPZ98CScUJxqjq/iYqaKvXytA5kjw63K1n7QvgYqFjZXvZwTlmA7UpDS
CBNLXUu2fcesbwjiCNnQ12QMFbz8tsbAgl6OC8Wpd/JepzFhupP29PHTgAANp/e3
VtnKJjpm9ooGZhVQ6ZNbMncznC31gGMBNrV19Nk7XEGhEr35VVCMWYQw/u9I88U+
6Fu0A5OL9Lk/ius/SVRuXoyjSYh2dVZqq38v4sWO0ebG5jmo6b6f/F/ILeGBAZOV
69mX2LLipNJZnVuJAL+Ka8sqpACoCBclyVyeeIrPsERJ1UK87CDGFq/499VmMNgS
5Kl+Orpyuu2/4C0brZEwr2MK7N5mXErMD9dEwhSyjxUshlPhTaZBsym3pJe8Gu66
yL+IHX6r0mKqdEcN68+UwDkoQwmUdexBmu0vcIcV8f/NT+AifvgK6ITQCr1G1SfU
qKSxSxyofVe9Ai19r1YMnyohqiviCqQqh/ThpnDDnoOqj2j0S0Wg/yIwm4T2AhTm
Zff73dhFyIdYIPmNVYvURwwVpzK7Z9P6HFhFOiiytDss/kxrAiLf62Krodau1Cht
FkXrQ4NzZKuHwnKT6RxRNHkBftG2rfr/RD8LD6zz4ApNunLKmCxC+fusRpLdgOlf
fYHCLga+hc3bxaJA/27gdS8tg4sj1NBhXwnUZ3Zwvt+Buio5+qtj40U2hy24wzVS
BgILITwjyvVLJnWHHTjc65w/Gg3PP/u4jw5eSy1MWj/ChbfjzSTN6cDjlpoUxp1F
8vTfd6gcoh/mraELvbb7XXIolEzFlNgoo+hvDN+n27cbhegGx7Qe9Vgw6x6kFUsD
HSTFlfSlgoFLoxsOzZg5TFfl9ipJMYsjdMEZcF/4rIpekD1AT/AZaEzdTho8lm6x
B2vEy7zxXYT/f6AFmuSvMfZq8py6UIQSyWclfHIA0aDgwkJIfWZmJu3BkyZVMzqs
Qxk5g4ldERtEQAzNNXUIOYvFEP/yvEbdpYQ96bQY7oet+lCX75khWh4Q//jG+Od8
qkmQ6qVWFyj13mt491aRRev33iGzwqb7qt7AJioKCz84Hcg0yhMZA1wLwhtE8NMy
+4ImjSLP2X32GnnBlmPklrnPfqEx4KBDrUhZI+mCo7En4TnMbFJ2KswLM3OXWX9V
4BHCh58hQweQfJst8APw1MpNHrQuZm+tGzqIcU2SeMyboOR1txIyax0QtpUeBKxF
jPs5S1WtKuupmj3WTuSVw6leaO2PsQWkcHXhTpW87/ETeZHa3JIMHMKeAXvsjG+f
cd10piyWq5J64BECQ+NssC0qVZf4XzRbhmeuDzlEEu4qEGl5P749EUEjwpLhTUxN
6PRMNp01YGANGwe1jz+Plg8f0ZoR4Etfl9b7dYsj5DFZz6ZZ/WClEljowtiL+myS
t2R1gGOD0p3g6IOH0bNWvspS4AwEmOO9uXJxhyRcszsUIluRmjsuQaITLxQcgQwo
PH1cibCaVHJN/nrii9vvBjkKS5FtaclNUiLjkdfOhi0jd8kMPsIWXpY032mpiSKy
gy0s75OupQfcFDhl4135XCpOPmyCzSCLUAns/gbZa6/eK5Q5EqVvPys9iA307ZBc
+JD+FZvmg0J4SwAyiYMWvf6AxtqrTpuzC3OhRGN5lKa3g6GQuelPdzil7l1H1Fia
2tFZvRNhaEB3mIFDgNMoEpfsmOcRb7QYp6ZxSTjOdr60ITkbVrL9A7s7VCUXvK1g
E1zbNcPjJhBzVLHUJ1nktV6O4PNf3XUNydRyILE01ujWO3lXyJm84c3TFVZP9xx5
MUcLm9PpLMfj2/1zqQkc6JTNsFeiSJ9vC2fTLnr6lUyWGLIRfQ/XK0Ygq1boZbYL
w6FLlKFQf8iegVqD4CmS8aed/PtyXZqg3sbjO6aQoootDuCwHuU//01t754kqNb6
vY4gNGM7uDsJc8c5ccGt7RqW9rb2rhOFg6h7c3gNw65eYIUKyn2LiezxkpBKSxjE
/VdTK2dOal1gGvzhnzz3L1mWVDVJ4HImtTbSlQkuZxyRkN0AtNv63qnMa7uPn+tD
I8uqTP96qQDAOdOXTNFu6EH1btYd3tGygkrQQBgAGT2f6wwFPKPj7uZPHt14D+7C
df3KAOnEXKnDmpMofIOpvWz2kMkD4KFq6SN4RNE8TQlRt1pqyyz1GJDixX9bg2Oh
Ldiy3EKxTqxgU0wjGfpp4hkPsHU17pWC6DWNIQR30kmLaRV3W3jvl2viirzIqNJB
PSULSJZ2JVno9WTNwoRGiaoZFyxTrrXGS2ZL15QRfQ9DDVsGrXhlkBEKegrzHjzi
QibYJd2zeausaQB3fbyuseRv5q1R7Nho/k9ADApM29ZMZOJmhNrhyf11SfEVZh7z
J+tpQLTjKAemIjvm9gsGN2qcJnA11qDrAsKZHJOfiSc2Jcx7x4cKMg2LrT7UgRWe
JDzbDqeMKw+ehg7QEHg39f2xDHYXj3nnhwS7Ha43g5i81yoTRkrR/YUeRZrrh62j
fWrRpmUF8SGnZe3OuPW9zgYdB+K+sWROpSngg7bP8I4bMfd45YxTtnNvkOdXPJaD
lmMh5CiZfWe3bLkPmEKPYRH+FPvUvHr2gVd5etjdDfla02GOVK3vhvnzyFEjDyRz
171rKxMr1GpxApYrDc8A0FcKUOe35xgAe0jgen/tkh9UFmosavAvSzVmlDdWGyXm
03/L2VRRil6AzLR/cDbBG18ZcVlHq88NZkv045a7pvgv3wAmkMSpNVro6gls5+jA
d/bI1xE5r6SQMVdY8+D/vfNBl/6a5VnGdL4Og8O9bu6un7cYM3tu5G1tf0gMpMKN
czMk5saPB/kecZLlfnidFFv9IJt6TaY4/ThCUy11zvaVTa97TrELqztePdNh3E6j
boOrbPY/FkJWJ+YDI7X6bZqswpeKCGIlq8vjTcK/zgqlROEGfabKf3iuc2EG62ja
DGbN2QP2isjOE+WTwyL1ZHTRMXI2dWUXKH8LD2U2741kaPJijCz3I8qWnlYEdLzC
w1y1S6bulHIRYPDr2yitqlo6zw9AQvgA0XNPgkf+hPQkGwMixF7VDrzau4mI/Q/N
BZUh33o0/G7QEjFOYtyHlXRKUMIFQ9gpR1RnJvihng5m3pyhfQhPvK089q5dfFxT
XYpCMs99Ni3ayUrEn/0ssJbvZf+OxEPzmYzlfOvosXZ4du18HchcS0i+0AVhIj7s
bDIFxnM6jlYrw6YJUgwnz4eOr51wg0w04FPPgX13ABQ+cDXE/LYR1glsD/X0nRwu
UbU/18rWFdhb005+1s3pGHsTcbaXf9UYjZHY6kxY8F1eMGPZVrtl6qYvKQ61vyAa
dsdEC1yOBH/0QHaY0xnUXcUoFwEd4XFsnXV5h0GLWI+gn86AUJ8RNnOg/PfWu4aj
HCyCndTKRujTdJna4cnOPLTF6ShrKn+CGxhIi/kcbE2+kWQlXGRLHBrKrtz0xNHQ
w+eZK2ccdks/xsHg8MmMoyYm/AqoTpNCnsMsTd2KU+zC7F9MHY1YY22CAOZ+5oBM
94xxVTYtsKxHsJ8L02NXgikpdGtKtw0+me2dz3qaZ3LIgPILnR1OZxFWjrUcyVja
OalOZrvlHpGQvakGn7UviBzAgaZQf1WNoohv3OwSL/waU5vwxwZeYAkxefJ2NzTA
mfIUEBRTrVBLiub6L3UalHpVOsyk9VqP/qWEVPKHLCL3TnT3+hI7vIYtma4ODHff
vtTlgkcUDbXkX8pZS+E+MeWRnswhIgqBqDQFaF1hn/hLiu5ZKe3g6teTHs2LJKVa
cCPYgXURhoHnjhCoaq+O8Uy1PaFWdadB8PlMGRs9mun9Oq1oB/N/B+ChOeu8V6Eh
3rFPyHvvR4H7T6PQN2Teo/VTi8Y7J/EHWRJND2tKFJ5qgLQSkG7XLpL2Jk3MmYoB
kj+pTBUCaDf2lfFgKoSxZeQBbF09j+iuAlv9Uvp7Q9CcQr9j32/METG8QgRvWjAF
Ki61ETkyfqt3vIKPUFt5iVG2OW54aV3iTNtE3UX9VKLfFlfteFOJ/VwlzYDRhk+R
Zs2HB1jDh/gfAsIE11i5qWS+qVZO/nV9N5Ura3L/JC6+RcUvPdE9vD0RRIaVB9lz
4JBNCyGmUu4WUMvcjcvkQdl0o0eeP5K679zUTofnM5nbmEBLYOTrYdF8qGBPxaZL
XoBiWph+bAGkKXU+SoatKqokpV2PCdxo89eqeTfpO8osGDEdl6HVu0hnwf91vxxi
FHpbE9+0+LIkUbKqfpa83ihHeS0pDDZheBGrvpMRl01ibOmFJi4KHg8ndz23O6Ph
Q+94fFmgelzEMDHx9nIduxqqKeuFqZjNtsGR1gv1WG83WTQFv2h3NQtyvB3Kh6PW
39Ax82S4icqovOxgw6GpksY1B5oXE9wbB4b9qfIJQcpMQa9j6NWaNb34LP9ShrwA
5dR0iT+QqPyOO/siJkpR4H6YMeuYpoFNEMs5+3YSCj5cf6HE3IACSFjSCQRNIhGR
Js4S6aZG86GlSthUct3HE5aAdE3t0jq7XcmW5IzBxdyk4dLPf78oG+c5Yy20xjke
mxJdcMQm68jnuC+E7o+7M98rJnpwMJk+RrvI5Zh74PcyfLoMx+bkH/S5FmNPdFPU
WibznHbzsIrGa0p9Kn8RYWlzOQT6qzEQ49VwV68F1IOCuHZ/xHfw1J40wpjw5kiX
8L/xqrEwtsF9oPFUnlYL0HuMrnAxmxnjX59mdNQy8c2y0BlOx/3eufQdWqJL45eL
lBxnG1BYDH7SOaoKgs6tSWfVFUsDVhNeDaF03cQ3J18+pcS1Pk1ASHY1elHcmehb
DftmB0NGcyVwZyGax0ys2NBz1sPOhwcpZOc8jpGlVT1Q2OF4Xdhic5+mOyEdILQF
UBOba99zxfDMESNSYBoC4UiRzwVg0QGKk40/Gg2xKcjDJcmHNG9JPHWHxZo4tVCx
Xouai7tu12SVX26W7iSQB5dGr3bV26ss1+B0HlAjmTF9EktxBqK7IJYq1NCmAxqf
FlXmKWBPtlzDl6jLv2/2bB8Eoz8B9yT0tDqHxeyDHR69FSxh8UwCVjJFzgdK3UE/
+dqWwBLi0XsezJzBe++QBGwHpIsn0CIlDA0NZmvkE21FdiKmzXuq1FYUwhh3zKMN
XwxDREBZJ9q8FYyM5ADyJlhQ00edXRpCOsQecoFW0PCmLd6l9ykDFtyoU+pXAH2Q
NzDkG4wwMdqD/S7PmrutFWLVCnazbRRLnLnuXjxXEKxg7WSyn/q4t7oeLKLEzoZw
KV+rnPG2j4WGQ7C5ETHYK7xVSbCLd+fGyN4WC463glFt2SsLZSyDHSFyoQdC8USd
OzmIOI41omXJ2JX8VS52vrjgs23YkcLTKsxJZi45ZKgXr5EeEXlh7TrLeRQXcg+i
0LAM+Xzw8C4DmFgA4WJSrwNo79eVWXUfKOp+hgCjwOlL0YRI1/+WOtOtpl8KiuZk
t2RoQveDeph0/oJNbouL7xCCs25L+EB1RFfptImWxi84MD809Oz/gTLT+L5AT+/C
UH5x+5rd/4sN15JMoTUj353hqW9qN3GcdTbPq9PaeT58IH+D8UznGDQXqi/GW2Iw
xOgmJ02ohGiFiEEWvjCtaTikSusYQuEUr33aBCvzXXGS5lrTu++51ZevKVX9Knkk
Z3iYYe1yeIIk2JaaAYdVA5l6VMvX7+eQQri3WCnI/NQLkovz55aZFW6bmQGVN2JB
SJBLSf3I48/5yzHWbrIa50ijO+F3tq/QWBdlwf3sOXr1q2OQc8dWV0IgRLwQtovN
Vtpfgw0ir6fmVVRe8wm0pOaJgin3kIgR8/s87ISRhGIj8RBGedeid0KqX5w/nM8I
KzhfAkdYLYB7u5zRgT5O8/2E8lLDVofztBWNiK1TLKL7+7AA1CEh60hWmPQXd5nC
ThLl6UeW5S2teWXG9GLxZkRuU4dv7V2egofPgrvr+dpNDVdXBhBFfP2KntNq/Ny7
DCCrePezcWYZccA2ZS9XALA5eGf1YI4tGJzVuTRPxS8pknuWf+7YPS1xNkhCgo8T
t09EZH4KzV4KcbIIVyMJ9GAyAK5n8zZPOfRN7plWFW3Gh/Ra2/SeDthbeCVxliuI
d567qqweimjZcVJzFva7LQ6hW2CGPQzarOiOGeimGtum8uB0bWHaW/VTNko0bWuy
4LywOxW4kdZ3pEBqtzuFfpK/Fjv2jYtxsxfgRei8OudmYlGoMfyfpWBiCKdAmMOR
JChUAl+YLVvwPKWDt1jpt4FT1R8mEqmcnEML8q5MsMHUXTn9PH+ftl3pmPO3wu30
rl9i4pPYuYYF8qMN/gjHQbSDG/v9v8XpibPgqT1kbjiW7VqCQySJqbdilahDc6xj
o72Rbnm7l0pXy29OdFcGD/r3BJ2XAtJA72iz3ffU16Mr/bGodK2osIZCawpmshBS
htGYy3Rr5tp+0S/Qo8jbblc/nZ2FsADh9UmfuKqF5W7UALECkDTz4hIVhVvz2CGy
RmNvwkmJwolLGMJs/7MvTHPzD9v+PLTH2lBCqejVeGa6+sQQ9DxbtNxq3y0dDMFn
qu2+KNcxsVA39uD8w6ZYmGOoAVfRfEdKBJmO+94ClNP3BYXjkJt8L0tooKoH57j/
zgOIetRV9PU6UiEQs0rJmonkGIYnY+U3dJl1FODVL2INeofCDTVGxdEm2wEo+4FK
Hse92aY1wdtHXmO6KBbk4hSf6zm92ToTiun6dNj2JMmPbqMl06oSFZ3Gpxn+6ysI
TS9WbMkd8tnGws2ra48TisTXjltqi1IqzBndbxYXF6LtcomkEWSkrbPzyUp5r4eI
/iOho5CX0isgpRpBFET6JysPmkRny2GHjLPm9vpkpSHTb1agyT3PlHvm7hzF9Kff
po/YavEzsLeINQWyYJsD1lcre5YT+G0MiaJFtLslLFgpt/w1S7u+zc5xTzOOsk2E
tRuYjBnGx5Z94/Pg/FW3zTk2nPEtr+RCs6jh3iwawvlP0+7k0QjjFBs7RUpOgGfC
bfrdqF0lQ7obLc6hVoYggJtltG48uhdWqTcV5on+wr2dKxjVHgI4P95VMgtpZ7Jo
f+IRnl25S2K3uKdpj5qmkvXfdMuYfuMboraGpkjYrxZeUduNcHMkBO5XupvrEdgm
RC1W6JSiifXtiz/iZsur8PqnA9/wjiHvDKiX4Bb66i4shH+XfzivwPZvX4BDOUJo
kwcbM2NGzGZBIThDgt6a/F1e9zNJ+X89P8aTSshtNtj0jEputtZSpvE1mCKlC36h
V5ERV1uIO810KUAjh7WSfbY8/rA+JEI8QBgigsIuH99D85prr8wN+q6lKlx6EZEr
BD6F/Gq3gSnwqrVQKeltyyYvVu5mGJIpmgEURTPAi7XE+HOEPrYXZ/baWJ5FnxCM
QuMEj36VcIo2uSW4KM1gGsjz1YPLE6UPUEU/7MIAF+7PEpWR5JOHBBbzIi5uNkvD
cLuWmQGWPb/uWK58/a4fcTt/LU2ML4mXSeLnwumBzjPYrIITAffc7k+e+xnLBidO
DkXKsZm0mxhHiawzH30JdSy/QBS1D8eKY3Qcb5F+IEHWfcP5FD1gmjCnC9BP4I+v
D5qBrQXrE+/XDEjXtCX2Dq5AqHh52Q5m2agUm5LjNV8Sx5lsPG+OBEaCYq6GGDyr
GXV6fApM21xdEtdtmL+z/B+RK8WOdtzcORM1ZoIdguWG3WbGN/6DvaT7tHIcMqLr
b7zUEVG7b4ZHpa3FZY1UsHYmhx1PGgbZGoMd5uW1gvmIPMVa7WesEuVGjq8RYWHN
JmiBtwTQCF1vOLrhkiHsZ9AMgsFl7eJopHMdHqJkosXx1Z/R+3gSppgEIwWiUCnm
JGJVto00fOCZYq8VTxustiv4mrKYpH7+9I4fhLKIzVerMXvfH7zVkZYtdAgMqo20
81L/8GJIyrDeQRQiZcLOoCp1+gmZBjasd3qx2vry0iSpSJ1QVY23HaBT/WmE98El
DbAumjFlYo5dhr8tnEXudALLQlvNW9CaPXdreFBeqtENWwFuSQHpo6Ypt2RErot6
gtVC4HqnVfZAYFPNJlBRT6rs14+NgmoowF0986wBYySDzdtQrXc9z94PHP9dcuTX
Vlx3aiZ2JdPGfBEkzwQFgou4WAFn/LgO/+xZntPM3xlmX7VHAkgU4eL4RHu6uFem
QkSDW4D0kzbLJ+IXQqRDf/LZwgGuC5TYZRcHcFAYVJ3GbNEDxrpLwXvHJbpUFiuI
oK+Ola8wgULYWW82uXEcWG9ujPCV7D69YPkbWYJWPAqDRFGPfKEWeERrMpcypoTW
9pdbJliY/zjAXwAtnbtYfE/QmG5vvQF/QaI9SJq7fRtkvTQn1UhbTZp4oo26h13G
f7N5B1mg6A85trtm+euhinQe8OJY5jtzZR/uH5maOVvRSyYCSIMnZaiIUIuNnZTG
VqaCmPpEb4muW8l+0G4LAnctaN+neItZS5K7Q0s41RPbigaTF9tMFfm8uglOM7t6
aMKDamK6Ivg4RoKsJSIul/bTRjcjN0aQk7hpZctPhNkctORWkru/qRcvF8utTkYQ
0bfklDvGN11Z8hjYLo+tckSopX+ZqwoQYAg5RtxPl8xebvNRKljlMPD7NPZVdZfY
kvlfyONbd5LwoWmjkFJTE92vOIPCnMafAiU9ibhXl1MDa1MrPKqZ10EpOAcliOEu
QfEZQGH0Q8DNRos8r8tw8NwCZgwHEamizWI1yDuN1kADufybVkhLyajY2ZXVVX+3
3LqUF3YkwCrA1+R1MFJOCQ/aqPjLu9LngKjrTAfkSvWJyCm9EQ3i/y8JiEdDfyhO
V7/eVV2NxG66OF/lg01/bqAtH1Xycx3OSKEbiA2W8rGCI+7rZ73FBAU1RZUjrq5T
CDq1To/s7PEY9o+n07mW/ZmiSRu5ccmTZ5c9paOuVHcwa8EOOy5fbjhK2BzH88KE
0b2zpN4U80ETZrz606r1/FdOZCdnc7kTIHKbvpuYuFk9oY3ksQIx1CtU9ccwJohX
Mwg/2e7EdkxHFSDhiFFqcsls/azKrhZ/TMK3Q+/nbrP0k/Ir2yqpyPl6tYRYcn3y
eE+D35rIhhvm79Yvbf2Rilg3lXMO5Q0h2B7VnvI3FA4Vqs9akSrIOYOoyjEkF1g2
jBR0Hh07qasU+K5l8fmZH3ZIRpU4WANA2uVkZ2KYSltaOPuPlUxHbVGrc+Ci8gbP
fCupPBhS3OnZKUNDvFTRe+tfcMbrJfst8e1fIPck/vG8D53ehMmEIrlhCKCubZXJ
4dMA/nqsghQqyexmYh5taYgzZfA2hKhcURXIEGaLRXy/c0yYlFGtJaxu5qN9txy3
gt63aUJX3TYgl5f3vIUOAuGQj8/6eix8qLc1wSBbIn3ylUpjbIkbR3cVNOQ+6LfU
mWw7To6O9vCtFjtqQtp+TuyPE4O2tWmSuBHJD/G1JW7eD+nEXEeKsX4eDX5xsegp
NSmQEx5R4OIsAhYqdn9ITjHTT/Oq5gl+qu7vaicO1wpY3FzYuMRc3z0n7RDtaTcI
QHQiiNrp1GkRmUfKtkYpipHHdNzb6qgYR1MgxpL35Gkkw5yxqF+sr1BiZXbSiZIp
OY7x/TH0cnmVzhMEWhjmsQO9P1C33huOC/OULHH+n5xc/4QJc/iElNjtX9IIeHaR
bzcn6qgp779LANR9JVkGpYuooovG8VWTE3myDUScQzvgfnnsH7fmbPmQ5RVwDNFS
xE+0COm10XOdwCVsj2NDI+Ct7T21b0dkd+jcfxwxS2D6it7Js3/Bo/YSSOY7k42n
y6hf6cI0cWD7T0SjafCvqnQ+p8PQwaNJj1TIiuOjQr4OI5nGkdSYmixOQ2AGeTAg
0Qz0PmdLgTJb+34Ex7GZdZk8RMwKAydLPmiDIT3RlXt+lMhlguYvnXyK9vLwPtkY
y/xlxT8itHtb5zWDAKim/l2cUQeJAV8QSupqOz3abv1Lx7qDAge1EGQnFznRks7a
IAAt3Q/6YaigXvrnPhw1nOu0ZHBOLPC7fzoLR4s6qlNEcVwBeQ0HhMupprmFk9NI
TR4O03bJlyzAQEG5g18nf83asT6XA5j6Gf82/ZRqnVoNVOM8OKhHWfw3F5EtZ6bt
napNrtgyBDSMLkRY4gfqA6CY9AxpRvN0f1+szN7ICcEINJgxQnadDY/Mta1h43OB
OgAoYlAkiuyrXnehsPuYSJG78Rd/u8LVVQY1AXMC8hlt2IqLkf51f6f+olUT1og1
do4EQ2Je2I1nPVxE+DqOSmEpyaYasz9sqRHrNEbNxpgGXEW5NOgbHzdhBvD2u5/R
jvPigs1ls3NovSQmeaJsTCsViRzWutncvl8TtpvYp6zvbl5K4PgwC8b+uykHXMPw
LO7HrFCQy8UmG0bXE4EjbHDiFivIRvzo/TcEZmwgkfNYqNi3XrTsze3GtdBoy5uQ
kPdHm71otXLGe+glc45ftpir13IfzuNcwINIosQRYj2/7E1hoBKiey4oph3B285P
/r/+ESue7NeKF9b+SsAqi2LJSHoRN2cTxf4KrRHPSG6HwuzEmjT8lapSRJmTC0+L
JSVRjMofM+ZRuL40sSb7fJFsVDkEFv7u5HjhSQDu+nUSo+NgiVI/lEvtM9K5LGIQ
32YrH8Hq3tQFK3k6lwwVHs8VCkrVtAmc9KvoIM9Kdef8EJhALd5mgKgTjT9NFpga
y1nuCV/fFUmz+mSlgnMjjXslQkPkupCvMUwLrKec1Ldc3HNMkz49KHAUfQlyfh4X
IB66ZzPq13DqTmtGG5wvf+tgxrDgVvB4IVXIjjviLnGvoLmA/SAvZq8T6iPSyS78
gAtMX/qL6+pDo+pA8wlWfWn0cISHpw2vaz/nNoAP8V6MkBECyc9XD/SdmFZX9yax
Fjd2iUciGvlsR8iBHMNVrZBH5x+H2xyoCYQdYI6w3QlVWmZ7biQtdx3q4884Pr89
/H/Nhmk7qrdH6AA0dZ9V5wS4kOxm6CmwR7+uge1jQdLJbxwBgTs7wqZtmW4/Gt9v
nPFqqDP/0CVee4A1MXfqOYxc0wNgsngp7vy5OLIN8yKWiS3qKTjsTFCoFAbEhoZM
apMKdHDFVIP4yEHvVv78wQEHkr00X9bNv2t9VIbc9UxJZi0VPJcs+g8EelLKBj5b
4HTBHrh629bMgWoqwwIZwsl5lhNDzyYEF5/WoemPubFHWJdV3fvzgfkde4JMkvfe
ckTKZYPpkXzwCdPNThsNKjv4+8ZeyZ/Ent6mMMYEHHNGhnIcTOM1p93lki9QBRHw
6u4uRfOZLktAmXLVo3DpvAi/ETlZI30DclpZXKJV+sS0gseREd78O0t06aYR9gWA
mpS/6eq3sCcVLImzkcMlFXXU3RvSQA+juqxx3UlGnid5U/5mBKrW/z+W2LOZZfxl
5MiyCnRemhyCtGVn0R3jS1ym9uGnNks3HK85b0yiuWUcAhzSVuyvXRdct7Gs+cki
38kx1r0l9OvvhfOwanGJBCJiSnzZJCWtums4D7+3K/AIP2i333Mqhx3bm2Za1ZNv
J1tsFQxvwX62eK5uFQlxjkORFUeKOlt2VTB14/+uLWZkQ5+iojqZ4OO9w10twaIC
tm48GsM/KC93FR7t7YtwfxEKRxFhOXaqcYofuFGx8r+zN3LJyonhvG2cqMrRySBo
o555VUIB2SP7/2k34RX6UtWb6Zo/LxDxL0TLaLJYcQ81+keXhfo0dBI+0VxLddve
++lB601uXivd+NdYsm23hHkRI7dV2h6gAsXRJ10PmRB9MnyZLska/CTM/4GBt9wv
xCeecSOBm3tpg6vuOs6x2VKW2HBHZE6A75dAFKGlzfq3jDZhK8SRiF0atx/Qqnsj
qj2hbmJsmrWDLUDpQRx/TxJYmDH1XhyKz0k4QWa++Yipf0DJzWBxe7sxijFNJD1H
N5PzK3vFp+svM0LMnDOYsbI9HROdhbkjZBsbkQkyHYSYZ6Oe8ncK4G0c3SitvoOp
bQmU86Ie3sbX6mxQGKRfWB0/XjeWHwnGzbFlpe3QWPz7AFkwchO+GR/hhVLYnP7d
yg5DQQuGG/nS2KpSXtF/Kjv3cYdAuvChAwtuPN1dMecmzygq8I38TZXKjRQxNHbD
my0Ljgtvz/1X82mW6rp0A6A0G6hpqn47eRK7mqjTEMloSg/uaiFnfxoanPfZ9oPE
jgwlXG52S76ozEiOa06Yhou6Nqm2sC5X9Pd6A9mRF4oTdT6GmYbYeazyddLZLW14
KPSVzU0XmeA1qiePro7EB6/n3YW+CSjDx3BAZN+STNhCgMx4KzukWAsxIF9Yhn5K
AEGuSz7C17so7qnue89P8FNprQDadNDr6gMAFdRbPCPtQ7q4OyzYyd/dQKxqe/nf
9q1ZcOdnr58nmPmTpDDh8v5fH3OQonzvxYJhoFAFtDN87WtDb7jeNcPF0jtYhlR9
hRpjeN4RUeDrLiRYQDLVxxHt161Jg3DHP4Gm5mwb0xHltOLLVVqF6duMH3Bkzibw
xCRJ5QC0YiPqKMhZkAqjQl0vtxvfDYOYmTRDCtRWneD24goc/LtWcyP6DqYiNFXw
yNTp/c/l5FuRUyD+VG59M8mYM/t1K69p8BLnFOs2zRxLatIOOeE8mFGhQKlk2z9x
vXU+MfcGslKNdakp5Ogo07TQZanLcPSEp03nxTcsLrd9ABXaV+CNyoOkidU4a5hR
n0PEqtOiO9IlcQh5k0LUQ/jhe2RvaEVwI7HPy00XNTL5oM2pEXLGZeaU9tcICQ23
O+N+Q7QqWNme5bHs+J497gSyJAvCTrLK4itz2lzi+s1hTmoXceaNCDCJkNfqJzAc
ZeO/Lq2p1Lq8f5H3N6CmoTJb3bqoTJvUq+5La/LnHa2P8RUgcNX0X44wf/TfwyFP
c+/CfW8ezWXcfgU12KYuIR8uVVKa8Yt4gd6BBz5+abva/rRaQqO/nJq1V7UauCLL
z3G06Znx2wl3cqHDTubLQSK3Ifp+tIj0anHCwDzii4WPITjkBGNhX1QGW4jOx6Ru
OZ07J8iAaosauV4XW9t5BopyxC+FWzfFfj2KGdXiPhwFyMFoLmFNoatsWNSxPbVJ
s06Lw6ZY6u9t5lnx3NGjGxCanbnDPDEjt9ogZE7b4p23FImFFHIra9AukuHVY0Op
IPdwkgZoELhcOVp8Du79kbghC6TrkpuekQ6lIGnbMEZRGMxPjh4naHi5gHkw1i07
qZkftYUijva8nGbW0hfeD+YxoYEcWf4PhorX9qTgvdM9m4eb7viHqZheXxJXYmRA
++mKhehFDMnVVL3O3uSgZ+z3uRugJAm4U+ffZLtGqB3WLJUiuEJ3TaYr7ydrFZln
BZ9NlM7jVc3DCFm3GPoD+LzBJTPIGCRU5liQPpbMdga5Iyq3cq7mI7uviwJ6KJwQ
aoV4nE4XPD3RbSoH9UPH+XBUSKvyOsErQRAkrY0I+lewIvXL0EwA0NJw4wyVxDPt
YURGNL2PDxnwgF7HnC/jL0dMpQmbCk2F7xzyUwhN77hFnT36ufzvHILDc8hWE3Ev
ugkNyVd2dlYXgyRYrhsHubcGjSKjGKQRabo4jBVkVtnEdHa95k83MnY5sWOrCyz9
3EPj+OxwYjvmmyytRErFsZJMQmeO933JiUXIYK1/3nD1j7y9qE2RNTc5cMOD0oux
5lClTK448tks9vnDM69gZyLDs+0UzQ+8/8bxpuH2zKEtZqtVzq3IMks2oPDdwu2a
0g506dCwoNuhX+h+cnxwXt2YD1naC/dEKn7OhAMKnriuFjwv5hqh/KyZkqw+nbNg
FR3nG2A5IhTYnM43I48+UWwbVoXu25bM4xamYUrhlooTtgCwFOqtDEDubrpmEY7K
yww8up/7T35q7iTs2t4X/X1siYDujqGTHBCkKer+rZeAX3/UnhVAUd9rBn7FfzdD
fqeS5fJUtOffqqyZSvhgGJkn7cMUTO2fLPPv4MEUvhYLuhkupxeEUrWoJLLVnUDj
9KwzKaDDlN2i4frRubIWIGbAfZySY/umQ3D3mcOtV4ebxoQelXwnREXLjjzy3YEb
BA+HJBOZCqlWL4bCTxehmQNbmJjDMepMeEBszmCZLulIsId+7/Z9yMXX26rbMNCr
vQaBay33TbbWRvX9LR8C6tzrCKNDwkVdyFGQQNV1AlCSgUmxIZbAipLKbSuZVtTq
Yl4qltQRiftd9wLvZeZxUQAmIod6CZGzRJgscWa3zzIP9hhxXWQmlOcsRy6pPj46
osGb2Cx7TMx0GgXTukOjz12ziAYjBMmU7m97hcIuhMI/NSXfxOx25o0heVagF1nQ
mIsfz+DvjKw/aayuLxFSfgq3WXrXO7Vm6fMaN4hQSnxjqsDiWOsZtI1e3WvSoY5+
PNTC7Nc7iZOZa+uPNAt7FCComLagGBQhcW/Y2nfMgsVpeoZk/KTEVYe2bd9wYBG+
L3A///Tc1sz8KFmOiWV4nKfBy6ldtmN09EqWFXh8MVmVWmGuHymjLE3KAtKWc3eZ
5o6K+7O3cizV87bCQ8bn0zpv+ad1ygwR25xJjtlQ0xTtssoKbFh4eBOi9XOw/aLX
nDFBK1xBN+qAr9mJ+30zMQrvzOX2IyocofgWmNLtjy4zVeb/DKYOn+C9kmbfk30H
oQj4/+zTNpymLBM/5Z+eBIa8qYvYQI9sC3MzSGoq+9SzbIFYYHivwLO+qY5Bcwz1
AEsLRKS7VPu4JakzzrPKvSbdUHkFzchL7FW3yf1wI40k6FVdXJzDz+KvrsDn4g2E
bBxA8LwxCFHLLAI02J0GY2DWCccrpvG5oYlthJlZzIHOMsSD971u2YIq3vc2zSWm
smc64tRJ2DvPol2A/Dg6RRegusbTTsJAcZ5WQBTeNY4Wph9vizVC933lpth4Xj8Z
gDHkEF0QR13ghaPOOB0TudzPilCojgXsfkdRh8YPBoSPzlxusq56AHA19jHFF11u
y9od/vkdSvteNGB2UXGKGCgNbBhw6gV7Kkpb2ppYXNDTDxUShZAf9MdTEV63ag38
e/tRzHqHZLfSu5c5m4ix7g/1cSyVZQgPDlf0aGSKR8DUu4ccP4b3A2iM++c3tgw5
fYqDU0TxyE1gKJVLQDiV01wYSa7kosrAyP3+hYVn/d9TLLUVx6DRi5eR0YfhSJlI
vl5h4ECpMrNzEK1H7Fm5bMk2ttBWjHkbU+ZzUouE3MgINUS3MmU0PUJ25LYyN5k6
qZn/lUHFavXKYL6Hf1Qb1NvjwN0atY4pqLv1GNrXxsduEJ4lWqfV2OS7N6HG5Q1p
WgYCJ36MK+IC9J5H+zibLA4v4Le1h99N6WRm4FhPNqm+SJMLeUcmSzxOeCOIeIXA
zo2yHtR4TjExbfXR1/Dts0IJ9G7n+X3x4l8XEHtKbvkQJALZcQrGrUXwy3pV4ZF1
fdob++eHhKCJPaBY7shD9CXbXoDMPz2t0N28WZfnYatFgLElKWP5B0ggx7cao5bh
a/ah6M0pI1YvdqABKpZQx7X+ltccxPQeGpO+69dfLi+KDOPRWdPYf+t+GqHPC0GN
y1t1yIiauiWnRf6rqTjLXQnwU9Rktuq45AS5vGLq+0Y96/FU31j1wWOQcQqn5eXH
7WKN9XkAWclQJg8qKDbcSCQBikgpkimELyqONulVivRX3Zo+xGlLr1EFqtVcjWTn
JVcEnFDXUpt4WNh5Gr/gHheS/JkF5yyiA2h5HmTyre6G7c2wXg3pI5XuKtvyXWP+
enCo1blj1sC4GYpsH9SIxmkiyqhJq6AEgrZIAr1K8t7CgEGbx+wvhpbsKusq+WmR
f3FgA4fn5OQ765ZKmpMn/EzVLB0X+CdPwSd3qx0tXYAFqRYX3T3OPjMTaaBdLrUE
WUAAkUf1BrVb4cI7jnYjZy8r0gO1cJwv+aVw62WebVFS43FpAf6VTBWY+aZx9FID
23NrEJvJw9bePjxwA5rfo81/lGPMyx3ophTGbJhn98OoutkAhSSywlsyfvTXXaQG
a7KXaZW3CBx22d0F5GdUjdr+HC5SZ/c3KNf9bEJdkH8W9ws9eocZUTZ87dNQlrP4
WATfkXAR3ESRlOGWHR9FZzMsG20S1ePQkRdrH8lffYZZHDZxsdnp/NTXy3485LLn
7SVGqMqkyUqz+7CTZW1pgAI/Df41HuJ3S696V8BtUHAtcPEtCVkcAWltRDEIEKOQ
VvDgT6JqW9xy2b0qif4M+BrueCgLPUAMP59LU0vPgBhfprTkHUusIf2OP/869Y16
JDsSQbQosCVZUOMAUqcoEJ10ma3HrkAHwBjEOPqtWlyPWHcbuzbE+NQmJ+Tda1Yj
7p4PsN+jyGoSQckvyoFwgxT/ACENL/qvo64kkxAB0gPwbADE1bXRihYh4wFarIrj
d035e8xtvhT9PQxEAUN6505eq1S+pny6PQ19XeyUfjCBxEL8SRLQvgqHyHXx86BQ
4ydsqr+Ck9jR2l5phOrW27UcIPoAFBm2ZuVKIhXmov9ABvtZeZV1zoYnI7708QGu
lKmS59gAJbQ42kcrapFcmjtii12T92J+iMKGtiz4yKZgif2LI9oT6U2Vkf4l0Gff
yW5AJD1t4EPXrb6MnHZsLszl5nDxq4mFbtGLJap+KqbZ4CODN41fMjEGM28IFfZm
A3oznCBMtZi6mFaz7S6rWOUbNu4w9swpACDgr2WnLdzxns62o0zKSS9I7OMr2IFd
1GYfIyqYgmJZfaIMU/aYWGty3Ha65hhRz+iUobYgsDBccIZEHnJvPm/aUW2LWXDX
F4ighTFz7eFr8mWEhwNy6kA2pHuBHalemYT0DECDQL2UE3zJoX8bDKRGZRPhdPJN
261EJvomq7VnVGssTQf7VQiVc8xdsat7xscxulq7ikbwtbUfPPqulRRb18kXB4yE
ThViakZheb2ZnuLnTOZL0yUotr9tBb1glrdTsbJHjFShazn5YPXcfJtwSJmgYeUd
y2EAg2sg7g32B0Z1uGxL1EMfBah+c9yjGLfHXi/KFNQesBRycXlSzTSqNnoxl4Ju
42t7KHRwxVQVyZJTmnCQ248eRfb3fNuP11O6GM9TlxHC5dEawCdGpJEWv05msAeC
KV/30TtFD3Z1Ec0IcJ1Oy/sVVsm2UAWQoapEdtddutvILTx3i8Dqy5JjQPHuZCi9
9DRco34m9Iue9jsw/AZk6aOD36exgDZFCE0pwnazH+jpS333qc4S2asWw81d4b3r
fmtCEmXvISu7FanQ9upIA7X4s5BR/hj7vB9xQUXG/QuXWSMW5N7BtH04J6yawZjP
xZDGThk/ymik9voV01ihActeuNzeGC/UHJr/G+8yu6GdbonUy2swnbJ0kRyFPwRI
vEJsMANoSFUXjP3xU1EsNoMgQkMIOpG8+W7oajWA5pmCifIBBT5nsKYAJvscdyho
5fB4IsJpigl4CTHAJ3vhJOWMb2cdX1i34vafNmc9atx9xQ3RR1OvkBqlq45ezaV1
5N9ejuJZqHixVSnolbqChit1DJFshvtCIzvvFASAQqsa2KdtELx8G1cgFrOmdo6b
kKsZt1R0bNt3Kh+3KxXatJZK9BSZrO4yIVyufWq95A+hmVjHZPUcQFA7tF+F7yEg
cIJ/pAs0PIkmaq3BkQbg0um+AHdpbMALMaaa9OwAo7c52NsmD4ZoVv0vBwAZIMFT
kYDXhHKsjEmSb2mOadNT3Kq3JV1sysnOMENPMAavNLZk41SXsHCwLmfitoL/+UFq
BZTM3+onrlScLEg1hzWD2yDPWiuiHUlRDROYFkd8vSx/kiH/5cjml4jthqPQ8ax1
WOwUg1RxbUP8VOkZKWAhm9dcBsbDLgKL2SXTkSw1WkIJ6YeGC8r4cOzTCmi8NlAE
dzNpb4iy74SUbe3wgB9EQtbevzyJfmTUw5DwYBU/sPm5JXrjXImWF3o0DJQhPa8M
MShqoPqmg5SI7BJHLImp0bYYdJPOS9YZ3n5LyAi9uHecEGzfX3+g61s8CMuXbXw5
zbS/lXKenicwPOT8tyYPzvqiUaphLnSmRuM0QtY90kVPM62NC3c8eIoHxkJzEIuy
7NsK708JRSgrwuyf35eLUVDuUVrWAb6pqm6SOM4N4aIHDSs2vSCkhutMlzgVVoFd
7s6U0WQbhUzebevRjP6L+uTHMPQ+LP7q1Bcqk79bUqsrXeAD1XGeGgmlk2Wzu3cM
jUkwfFTas5MB3zQnpHIZqW8Vw7lMrveloLDNX7knOSiVDcqI64n35KXKUhxCFGiH
NGcqXrWV5+DYts+sspzmRFJd8gV80jknUstnxUduwp+0SSNAFlEOcH776ZRIJEaR
I7ukJz0HFrgmnj0edUpSLAIWZuTw2sMd5JocjG/h9D+mEFqxml4CwjFoEOpH2BHZ
EOsApXhj9DU+VVPDsSdZ1fAfljKiaMgIS9qlBVL4XcPugXT2uCuSbcRvUzarw2ZV
za9KdYp0bXcC39sjx8FCfwyN5adSSSUWzYcU3ApWZHTt624kRiqpm4FIwyjFtIoz
uV8WKCmKcVKoSWTWTJbX+8YaE2tXRM69Ij6DgsPKexLuroElqy9hkwcRzkO8xGas
r23xF+BAepz5bii+XIoG2uW+FU+X9TRQ6QJQYuKou0irQeQ7GL5FW7Tk8066TKwi
h/GIOHDwrQHhTF/6obYuMglaaMnlmRoyoOyMQM0vN2Q1Q4neNcs8Tyec5qCiMhgU
5Ut2CbOtkBJAM0mi1veE8Fty/1t4y9rTfJXUAUdl6JiP/YodODMwyvG2sz9k3dcL
6YiTX65QUrf8nTRkj+y6X7AYHZIKhXZdpj7YJLq5dCExPHGClLHGfgx695AuBvVX
MKaAyCgdvFb/6naXbBSLUGenFt2oFS1/8RqVBv2sUaH73Wl8WNtP36GIy4vsQ25m
HPHsLrrnf4OqlSYXqjbp85IprqO3NduNcACZI5/VFNHYX7cRPq1wSaJOcIBDRGUj
mmgh1xYotzwknQ6z1lwSKqjglc8M0UqLg+vzBGEwklLjtK1t8BDyU9XDd3aGhTSk
B0OLoOvTZqzKsrb5nyslolOpnV3/RhbU/cm4TrtU416wgmnknnqGFQ8sNVFl7FI2
WpBgN7CCZ5uWndFZPrzTbIMHaECBWBbQ5HFaWh+bONePFeeOSqb7pa5PwMgZd4dP
wh3uOmprrJuSwJsOLOROmlUql0jvNb9jnrpUWFEoPEqsyDdQU9QoLcI3EQ9T/9H+
Ptw4DACCO4LriipaZjXJ0i/vU2NtqyzE8FIh2RHOaamV4iruno4yJNHKIUlRVM/9
xMA18OC+7mUJ3dDdWLbAwl0801OVPM8gblShXv5rHXxhWhP9jY2TusezGnpSAsO2
FyF+lVMYMLYdVZZtc72X4cXeEm/zJK95J55AzNkdMVdH5pXc7DZeUzc/sJkDCru/
AoIeWEW8+vSj4Kh7myNY1t/4ydkajgIog18Vy9X2C4xe3D3+gHCDBKjECil5FJsZ
4oQaLvlofiuy1gCcnh5ycPRnFrh5NP9ZXPPalVxL3veb+Yv9KPfLeWSYmmEwlM68
W2vEJynZFM29Xbbiz/Pwr8SD5DoMRGTNjcwvB/eHEs8z66cCyk4qWuXuMMI+Gjce
zesbRs63PbF+jDk/9y3v5POTOHvlyU5iUEn2mwcwNLoqKtMhvoxF0VhTDTQIqPeu
tH2MSUumleoVYAiwR4l5t5YPPgzMr+rXrdodWNNm3sfg2M+BL9Yp+BYvUfc/Z7iO
fDqJBq1owK7HZ+itA0pVzwbqvt9LV29TC4Y6ALde5po+CDSBYowQZI7lYamYbzT7
HrAxX/FCGR1gtCgoRHcrYLPNC7ZpLt3TTC5w0gPv08VNQQutkpsH0IoaL5epVar2
7GWG1OQWqQlWTQYsiKJnr+Y3SX+J4fK8tHa95uGAFXmTgfJ0wMtsQPONoA+Lep4K
G+xza1r25RgMN9KgiWL1VQSqFYRUx1NU2pwNP2J5u/CozgLLUbM24LnWAA+GX6Pp
hjN04B3mRXVYqVcXIW0bi/dLcB5rBV1DK/FyrlBToPopjq41e9ryVpZR7AokTrwX
1Xsm7zp7tw8IPdlHJa76Vt3rio0m77iSIF2dwCn/xEr6jBIGans8hH7Uz4CtLtVB
ezfX3DID9Sv19XCaTpcjA1neehip7X3PqF+U+w98+Gjb+0UtnYfYvAY+9rZizst/
2Ks+0fzy+qFJeph0QamalDZmqpiUrPH89TlSsEomxIm484yu1W6Oh+UsZ1x9mw3f
OdOCe1vecYAbPgKvkRJubRbhjpNOq+6Vhm5ebFcBuqc2jaTS2z2LhdvA+3i+VFOd
G3egofHUrOIzZGcNLq8NesVs4eJyZs5VImqCbbqkqA2B8hqXnO//oDRcWedSRWEw
yjFt0BlT8U2DT7DNpl1uPmJMoNnCzD+wYSrUUwlWD2rswbpOlMAH+5pnCYydnnd5
rF2dRZvCcCGtaZTyiSf3AIejbv5dBL27u16KfDhJUiqzbvTyZrNtnd/bVKxekCvQ
jYoduG+agfmiamYYnczXTLhzsGWDguUAUf53yfNpcyaBqKXX0G0oHtWXvhZFhW53
PT1dP9Z2Dt/btgTR3iYR6KJkltsjNAdqzVX06bjMhsfHghyEvGuIIIF6sEPSY/MO
SxLq0rALme1ewXSkUanx9dgN6ddysr0V8rsmsdoAvcMFyT6t7Aa19h29qiFrOEkG
3ZY4F9JmoTCeQRIzlXtByvz5+aVy1yhsy6wZ+wZVwmggkim+TBlrrDmQtzClV7jg
3X+RDoZ7R+NY7Kc18WCRBk7kf4TZNLVx5pDGKdhQ6DTYQc9itqOxX9nvZwc5/jBt
ZU3B6wWjgEZh72WMX2dCFIiNYNmh/Uaed9x/Md/wH+J8OKhGrIfQOHIMCmIdYGqu
zlBm0CTGWxrZRVsN9HjW8ZPqblpAHZg/GpLdjFhv+mqwFsDJ/GYmSeVLbC1OyLqx
+4+NnwFySjUix4gy5rBRYfSiGaEgfR+GF0OwuF5VPSNH+fohaEGYaR/43NI5AM4L
T2BCfb+YCB74oFwfB/zVYymCKK2CRBu4S5DuRaJgOWxN0fx4UtkV2reAlubcsYfO
YpY+E23JLDKhBWoJGsZbhBopDgswsNTyMHALgi8HeBJg42gKg8vxOIiIBwn1vhwO
DkCH2u32guCh6VLGI4vJ/VVMZogfbbPYHuSkrn6aLOuzaD0eu3yz4bbW0hj85e8w
UNXGM8zwjCLH4gkUznbnkyRn+RlfWqxIstaFmqhEhpg3jJgWD9nlEdwGcSFDBlvj
2NYx8QrXxz3Vb3dMu0/EFgRFoWio2mYD9UxpoXbKtglfRngMxVubGAb9tqb0bXu+
s1WJXzfpzkf8SARr7AJahQ/6j2J3iLKpXk3YZtqjRDtWZBCVpy0niM05lDMPJR1z
ECttC+lLQjucI5fQObDUTxtH60AjbgH+nJFe6Fd4ym6cGvWhELCrzI4MzzbZooIc
XHxKSN5rxysMrpMx3nKqd5ubn0KvyTi0V4CKrOkDUjUyt+BKfsbrdEHQivI/qfWs
WEkxo8DUM9P7Orlf2y7DtsjX+0w9T3G5jsQG9P/DQ55r1E8NpYM0sR8Nxf2MrF5E
KYxMyoQzeofwxbyjH+ThA3u7kujybIu78Ea5QENlTn5QPhryBl+vQ280CWj9g2sE
CN5a5sCGtyTrO02n+jgcbP8XYwgvJexOHoRzUPbMM/EI1snVxHNLEJWrx8wPGNQ/
nICjAYTKvYIsgr2eQXSSObRKmE8Zu7e6cUBlJYlez+l4OEAgwAg0a976n2UkKsPF
Yd+rpmGEjjwOb/ZdZF/rqpy6gFU8Dpl3+ehRSkb2kckSlklRx2S3yp/exEaCfgwJ
BedcyREvoPZUcpdVVeNxxCFngINkb598I2XrelCXYaZCn/HUMCFdhEj4a5fOvNHR
6Fs56VQOhLp2DoPOHc/BBb6m8dedoUeTk1r2oPkmQ6g6ZW0QjCKavnubMz8/iwVV
nrgHprK8H4einSx2lnON68pl3juRBbwmB0VFeoz06sPJsgJU+oHhataHtL05GTjT
bZCvg77Ttlp+pD5+NxlQ1hJKtbCk0cY8t3f99Vmk/ylEExSZr6zfKQCVbNHcPdsE
ePZtmakOrdTN1c8JWd/nMyonczAg7LRenVSWa7nWV/P9p3D5vqx8HWldm3njNv1H
2PCM8CEupmI/7M+xjjWQblz/Pfmn560YBEN3BQrGH5vm/M6fvfJQdFV/HSkUWQCy
FaXv+eKFnJMZS7rGtgxvHUbQQcBtOrzJeffINpXyfXzpDrB1rwXnttxrEUkjKjMX
GEMgU2GBQAwgd95aLqSjOoM9WNuTpB4brcYMve8/3soWudP3gjsMVlNSOzrU7h+0
USiko0pJs5xfgldv8FiykvjoDFhZSer0fksXGinSoKjBrVpD9lak1LI7l6vNukRH
SJyDt4Jt+UC1a6Z9E1f2ky+Mt4uUL96tHKNYheuZSLyx4UWGc1+BDNp72NbiInA9
8/OTLgW/r2pQvAIEq4KykE6h77jhQWc5eFyKYnfmHtAsxyq6AX6L55B3lLdln31M
neAadWHwCnQ2eLvSWl8URz17IpntvyfZGlUmKRCrv/5SkiH21uBrwpWX7xpHYpf7
1TNV9FisOVIfCQ/nJ6us2fpiVhUUXBouv2ulfuYCMtEEP6re/Ya0owLmS8vmMeoJ
7ZE/dOR3Rj8UAJRKrfXehlA4fZ9PyAzFz2HzhWXxChIFvyewADtHIHzInCzGUCUB
6vutETC9jP7mnzWM4wLtdCN5eduvVNLiB5jwE9F+0wbP/KV7T/KhkpRgHVw3sYcD
bX85IZDouITkBM9vGy6GZ37hHZwlcL7wpm0n6BEZDvmFg6t2mFUMxNcN+1fbUj8/
6FjfFUYdqqBacD9fm8gQDBB40tRQBl8enl13Fgs9VIjErLQHk90U4J3kPrjKHN/4
gFGSM5IYQatxhGUVWrv94dwHjOeArhcRs2+cqSwRCKF3FrFrLU3/VAdrAYG7LfDC
s4msDxvWrOb0UXbNHXuY+UyimNIrooJqTb5NyUgIZRSvvhOMQTWJiclQfU6E41uK
K9HJtfKtOdj9pL8184PivOiY6uzaAuNI20X1SMq+elMj0pWW178qZB2Sw8meI/cs
f99U5K1vuJh6X4YQb0yrflFwoECKN785JPKyhV/7oDdlqogD4ZkHM4lD/h4AKwPo
dwDBmoUo+OlxpoYhflt3JD9z9dgJ/dqp/j14VZfLTp/gTw8TL4D7PoxpGjqeiwlB
0w4HcS5kdWlOBbLFq9UfVanT68DrS2AJa3gAuuBnmZvV2/ycwJEeSsdGFcHQ3c6x
TjfOityMXDm1NAdFBXVgW8oWA1/EwshPPJcmx5JPVrTRE5GCstjw4+nKpcQo3cMb
e1vjg/NEgtg9rhUTtyZ8DiA0kB+xRjvt4qrNjX0QmTfAkOJ9mmaw1WCv9PigFafR
VatIbcULt3l7yc4pl2wmG2w0RaaPIRbcgSip9l9eqEFZZL5ndO0Gyp+0XjaWSgNy
5fdkUXgwF0ofvwbqDtT6VBL1LXZFm5nXigDVgUCxVtiuDMa6ghskN29ggrq/+pRQ
R9E2bUVmaceSD3PXN7vKnX75Z2GXlCfoVS1w58mghqtVSD4H8lD0jplMNnZBn9Kq
KCvStRLLRzS5JFvyPokUTXfIjYo5sFDBvQKh0uU1ohamKy679H87AyFXdfpCF7o6
X1N2Jl5r+GoT1e16IupXoc1gIcVLgJO00RTokhktRJkLEFVPPaqNs0XFRhQDIB6i
BmYRlGiOh72ex/z7pxDyJDhSAOahlvQE4fg0ymchKEo/x6E4MMQbPbaT94nKPUIP
vaZmfPWLXoQydwKv5NjIxdQL663cW3/lzCv9pgRaKI06UI0BmU7Ipxni4t5gcp4R
dmn8Xot3VcgNKMrslnozO6s2n9yBCQgD2Bnw5XfbVrpHnlAWsrRwtv0MJj+K20G7
mBBdc+PtXmsT9c19QqrbXl4q3B9R8g05mFLG0G07pZezlSrgB6VOh2qhKV4AqcB0
NO3/OiFlB53MnD7z5YWmV6dsWK6OhhXHpe8BYaTQsgcOk7Ha6/toH+LTED7Fvi+c
u78wgKoViuuOYdw5vNIPS3ki8ikmuQtJW/Du5fORU8buJxAT719iipZ/8arfyaZU
maH7cULuhoJAiOiQou7AWlMwdygcCoJuHuLt8XsMHXwGpuGFEGaWcYqXOXVniw+X
MeMN9AGKOg35KNdtpNR5PrfXessOY/BLFG/G38whGnxtjgUZVInLBNftm1eriW16
xwaT6Mn4mXL12EUSdBlx23jGr/Y4MOYj0UCb7rcTzjZDXM/XQlaL2iTZADcjyI7c
jakl/ScmrlcHs9bBFr3arLFFS5cRjfxv1a/sRLBQDmKPMMIgSDb/xJA4CwPuG6in
Nbexh7mNvRx19Tsb6WeHRB3khzg8zulQlFsNBa464qjiP31B5zm3ny9lyAyQJh/s
MWCouCrHXHZeD+M24kWL+E2LDFUZY0ay+5LyuK9tsxSU8C+rek2J5TBntic3h7Xt
qxmEuEBMzaMoayUsOyWVY4En4CZBOUVRP0fZusyDXIOzLbNyhVTI7tmBWSzZbpeT
0jF1aTkHmQWbJgOwS0w+soGr7l9iUWm5rhbT/wWHQi7ZCPfvMcAmtSwW/vfCcCq2
RK3649nOkPoonqbSNi7aeDQNI5+kw5JpoD1YsvYvCUsfcrn1oHO9Jnj0Jl9ql0Pz
1yaohPCJ8zzXx2EQ9oDGZ7smggz0+XCx8iwPHknTJLdJqXkg3PDJoJEjFwsbomiu
fQhxYbgugeJ5sFE8KtSXMc6XRQ39rkjQZw/tZXff7dz6L7nSrlVgIC/I7TnaqxjA
R6NYxXrN+QqyxGerGF7IxHytNK7bH90Y61pdmWYY3xnqmgPvSp1cD/Sdj7W8NFxo
HSwsCwTa9QDsCuToQicpCsB6Q8DU/tvVCYsRawWrz2FUOHveescmzoClSzGYQeMP
OPEs+GoFMKp1i5aaUAaRjvp2H3IfhZV1bxOnNcAAbQyYjemhehywQuk1RMTe3+4m
57FRn1fSbUnFWu04P8lg5smRlzHdF6txGlbuDhw638wQ1vlSRFphTsmhshRuL3h1
grSj/FSMgPG+AmcujY6mAIsa+rpus7ZP7F5YFgooiI4RKubQkO3vzzYhMuI5Snbc
VJkb75XrMsasoQNCo1wYsiFGDv+B7p5lZRMcyD8JTa5NDDX0u2b/m3cLlXO9tOcw
HdHXmyxqrbmhGTphpsK+AtivrAR8tVK4oNu6/trYeF4FHFKBjBxrWAwmc5FS0lec
cQnb0uE/44LBgndFIVMVE2eCZKUI0hLX0qHFTsMT+enhgiWfvBlouPi3E+BQkwX6
qt6aFvEhFtLPjqus9rYJlEycRYBjUvaJn7R6V+g67ytY6B5wAou/PfAHHXYAC2X1
HAvJO2hQdkMrBVebsc8Te418CwimuKLLHxKav16vEWJsH9aHstP8ZyzNoq0VLaQg
Fk9R0+nuLfclxYMUDSf48LL2tXUFeIFHFDO30QsdL3SdfMbS+IrA7sH71Vyi0C60
26NlUp/tIRlJFsCOg4QIu0RyGiKfz2QmCGwHyomIUk1c/pHn/m6IayNaNvJRPJIW
IfzdoBsF2LpnLsn/aftu4UU+t2M61zShbnf64S+50MUqmWhAlvXzUaA4nyEmO9zo
sFVHPBZcRKtkvaTy87mBO2OS/SK3ANuPWpDcoT9PVmjGXcqYhTOkskDJ70RZn8bR
nZxdn9XtrbqP5vi2jlHWihqnY2bTX1hvkEMBtO1BOqTxvGKImkAnNddCbImwhxQD
Z9q3enitMk3FbFpTmg3iLYdkV07/r/vT4TFKgdvT40xKBKy0irSFY+sj7Gy2VLga
onHjx6JDxHtKlvOPJL4Hlz1KNkwRW5UaWOJt7GCaj95ZO9zNmZarJEIHFDUTbtZw
FeCI1XZVWvgkgGhyENvMU+UbgCgKzE0vg2otpbtlmpOUVKNQr8jFulSUzBTjyd9s
0Hr9fPDgNWsAwINnffReXluAe0miEueZQ7mwpgpVRzFClTqhfgDNWfwBdKiFvNvj
sbmZBu/8yZ4JEwqgbwtnQmgsSJqmrrie0Z/0hEW+F8QFJ40Roi9w8qFq6NKqtyxi
e5HVwi7KCxpqsJZJi0ogSP6AzMUKn5JUgwVsOfLzRT96oMfSngqr4BXuegSIgBk3
ZQb/b/xSRjOOq7ppmoD41ekfkb4rLbKrUTNhvBRCHIB34ZvAu9UVyx/WDMyb4WRm
3RzlAefG3IelChvCbWgbW6znOI2qYJL6dfxvKSu/ecUoOLM4ul+hC2qSqKGlChlo
iGlAc5MZ1QAUaqnR1VU8iQVDkn9kEk+T5B8i5BxA7CUmflmreb5qL7NT41XjONbC
WQTFNma+v0iyKL3AGcXyRSOw2qT948l9pksVA9pPuQGbiuMLSAM6PbkjCo8yajAP
lRZLMN5CgtFqJO+30QcWokloWaq9rwOO0s5CtJsQ6MXtQjlFJwYWCBT8OdhoF8hA
+isFzx/klGDi1wGkpSI2FynR3P79MJlit6Nt3SpaJu4wbGEUIcTnwgSVxCvoKSlm
GxPAGdz11xG+r8AP5+zYfG4DmvdfPo1RnqMxs3uNwuT2LgyYsxE4V5Ly7oG2aONn
cKtXLZ3BaZiuBghKnGAEeEjuGStzW14kJsI5gDN8fon0m/j0O8dwpiSeuaaCIjVd
Nk//aHJ8uNsoTT8Xtn+7WFyZ7YVtwUiqyBdh7KpWDeVUTGdo9XWH2vL3Qfrn3BGk
ksw6qRFocB70TdmCiIJxdJhlDL4UA9P7hfI1PIgxg1/J2uVwr5lUvEf7teQ8y7Tz
6K6fuiCcd/5wb+jYgaiPSTGtKUmYa0ymDnNLS745R0VVSpE/oZCef51xyd3GzMWM
wV6bdQ4sSGClEbkvoACOm4/o7RxS7WWLSLqsOffiUGxtqOUuz498pSO9Mh99MP7T
AdJobljB1EMU2O6e5K8qKwKMtDE4G84QmuTlulICRLs9tyDHMJNo3E34cT/JX3Fh
PK3aRNbhNvmj4lEvUZuGYSUFbVEg7neZrqxe8BU2+Pw+YkAvwAtUS79yXyb0s1FC
SRvvPRehGN+Yz+b+MO3eXfxV+FCEBHY4aHkth9jEKTMJtaHupGYIDwmUftVxoRVV
f1lSsGR6dAPG1xMvoLkFK03AENvLnsfduL0QgE0nijrlNVtouGZXgqNKhyY7Vacc
jOBsutVVOdPBhiUlb3XEP9GGSPir1dVFKgFmdzgg1b1MbxhLoUR6qhfPZ7cqHYHx
dBNnKvXivVngL4pC3TSmCXyuri4gAlALwzEecPhNka390sqMyu1RNrDG5rXUro9Z
lryXKDYXk83uamUpDvHjPTkgth9Z5IPk9b77n7/QcqP80hYHc29137TKJ56+UCGi
APaKKRxgRXzsgeLHivJlm22c49OwwFj+MRz+PqlpyiGWLdUZtR5wxE/+R/wOjdKp
ZAzM/Pa7gf2KVjR7hoV993rBp0vUNDyqROaZDcn1VzPnLI8Ms/jXI0Ck4jInNOMO
2fWfH7Ro4HASW6Y2/3Qvrq/9zWqWaNireiRakaAXq+hWWV1uvqWXEz/btXeJx/k0
ETkFrYm+M47Oa8UdXCLuIcZ0MNyrDHT59ifArrUTTDOXoQVfITCVrAVHG66Zitet
i1Bt8x2BZ9gfZ/usW6+0Yqsutc5DqBdx4YFJipQCteGRUhsDRFCOG7/nOYwLtmnG
k0Qf+E7InWgL9apde0E2yfypq3ftBG9NFk0PohSNks9+JyEsRQakdSoFimXV3xx6
VRjJRxNHeTk0FQYs9jDotZz7z/lEnAWxTa1z7lrHDmPtuFR75DxV5ljZFQzvJ9Tx
+DSzcnEblYBDsn/GwS4AjreEVaiAWF/uWKtGtKUvSdH6Pd7KlOFWSOVsdhM1bH4V
xW8ggDRUiigx/3Er9FrDMRrYwvtKM+bBOrlPcxZpQZ+cX3T8t9mRwuHKsfHGKyp7
d/YtNqaaxUPn6NVBxg2giC5TZZKwXbGCs9pqN31eIZAUYTPtdZgIOatImwm+Ecv4
Gz/uCZsNksscRPULdAiS4JL5Rn6CvDD2IDTLGJfQUEAm6HK+yLQNMe/A9o20d7OG
iyMe2rLsmRNRGm6S0u0aAEIF8ioXuPfzAsgYv3wtP6K+7fVbQ/O62+8SD35Bixub
NGEsxaHzWfrbmzOciMu4bSUgJXRv0Y0MVsK/b2pIglLkcmoG2yUy+BYcEwzJ5hIP
EM+xO42giZv6M/ZYou0Iolf8d9B5IwpYZQlsBcRC6dgWHOsy7D+GPBX2Y8A4BreO
yR5QqDTB75fRVvtIQMYGKIMFPA+LRjbH6MqECllo7s38OnXIq863Q6U0VuRc73Gz
IHfaXPAx8n4H3I2DTMKvS7L+1R2I66m9l9A/J2lA71sFFe+D92CtTJYI0jxzu8Cq
HonNZxzqGfvkIGExGLLH+qZDUVBQKxUEHCcp9Jndt4YHbmW299Dkx8UQBfeB/ZXf
zi8bjoOhkz0Z9laygSLKRNGqZu/0bD0CWO5uaeOSuJJnmUAjAk6L6rXpITo3hKap
sw+w1uirPMR3+MZKeGB2K/xjrTHsxTzWcLxrHLl9SAouNStxbbFzdYT9iKqFC6sW
mgr9b928DlMBdcgKH2sLPzrX4FIuDZ3qWJ0XrZj0vCcoupx/bUMMeN9TKOTL5fxN
/2vDmsWZlo38nrDTq3sJcp2HvTnVI9UeI68gyLlAkX5DwtidnsZ3HHJSBcgwEDYm
tXpHGJi1TbAN9OfHrqaAsF8sYQa96XwVtYyMYf5Y7gyAt+BOS58+0e2yTUX2pyMh
O8AdiKuwOqGk6HJd87mtFaFzccc08Oa1xDAMNN4ta1DKNEp6E5QQXn+lHJfVL0l7
q1P82DqVGvjDnRlTF7RBeDCHvpMi+En/zazpMh+DlvW57BG5hiEAP9Kl8BaJdnyk
foV7K9kj/E8qQ3WkhbV3C3MBJIiKkPrSVnLI7+muxeohMrOtUPGmhTTZfLF75dmu
PRP9nXjaJxFDMlQLXk+ZADRgiJEzxCBHzrDvqCYe/yM7++uz7XXSr4VVyOOzHPd6
shzJYOvXNapQ0NXXnnChwIIxImXaxSrCqnwSsM5z9vUKnA0eonsiEL/pi0PwPxNm
AhjNh84OOtc66i7os+iLSvd6fQEh/diRjFxrAHSM/g/bzS6nEDyLWEzCUuHf8Jqz
0bwZSykuiEJfdmMEeXqs4i8mZT4QG75xvc8/BZ/1RhVHIdKMk6JOR3jYN8Sl983J
9i0/O3yY6rrlc+yoYweOWR77HjRdBcQwBk0TGQJ5v/FtJcOr2FE2HQ/USN9PzvfV
fdqsBHNO0fSELaJIJTi8lfzhqFuU08t1ZgaKWRt9jarGsHdaGfv9clglHML6/GOs
GiH5uLhQQXFte1xnowBO4iS321I2j0O6fVd1AQ7wC1od3fRJoF60WG8iWSBKj2CX
n9Fu8lojbKK840urIUAuhtd5CvJnxfKgn1uoI3TsrtkHV5JCqj/UmMYOI8ZNL86/
htJLpTQbUVx0+kSyp6nmYSxxqvyw0PPZTV35KITjkoI5gJyAcLom6cS7+sLrdyTn
Zt+kzhJZRG/OdnKKogz2v9TUzJydXvkBQX2bw3eIZw3pPqkdwMScbNRm4WNRYf/G
or79oukQNk4DJuV9TlzEDn7Jj4n9zb9qSC4hKH0N9RSEFCJQC8/RKpeccxgLx1js
ZQiN4I5OfTgj+BI0AO4AqiMZCQWyJgbC3K23PdD3C2JRAAaSHZDjNgI+F7rplbpV
R4p3Vi37RByJSsTPs6xy4BxXzV0wAcwLzpOJ7nQHRkCnjoktqkRs/aq3hkTT0hu4
XgRFv2xGy88R5S/XUvQd1IzLWft0vkuEXPz2Sn0NXSfhDH7EP+8eeUElybgvMkmQ
F7QPdQTuAXF6D1TLt9kbmiyWiXTcJ9eslB9u4+jo9WiY30ncViLD2dLMow0X/R69
Rz0BlJip7XDO1m23Y8+wc5756o9X9KqnJO6dc2ANk3E3q4ESzWwK68reELUTrYz2
ejfD51gwt8lSeShkAjN8OuugusxOAvvr4lYkvPG01kGTip153nzP/mO9ON5kWuTi
wv/U9U2h7KVIwgbtBDvMzu0JjqPqQzTyQpVN8bcpa1WPfC/1zWD/qGZdN3W4KYAw
V+OnSHKiTKgWqgYyUi8bYT1SQBSVhf9tjVdyba4zPturDUZ6WTv0UQa4BjH+RI9K
2VI4lh++QKR+R+V7/4gZfeNzRYJmAkLlJ5Tgub7fkkluk/vzdjR3k812+vhd48sn
YnEoJfjCDmBVolEGKlEEVsI1ewORLimMOk/Exh2EXt/ppWmTm3QN+pVItnbclLiw
P5KfdLYKrMQoZ4fBmCjaZyZLKpDL411lkHtRNCFjBGQz/CkHgEkWE9sOSQIPpyMl
m+VGq8S19bzQ6LzrqbreTyu+KUHpnaV9FVbu4IqLPlobupeM67q2Hf8eHpHx8K7L
Xeww2Qeb2VWA0sQ4dO2tAOleSt2U6lUWQeu2jAkS848P0s+FwJmNIws4NwBLl0gI
QgLnYBO0yixyQT02Bc/St4WkCjK5c5qGpAplijj9QmXLfgMzIPVDv47gQblcdFVy
BXLjCpFyht9yERCpnCIQk0/GLnDiTnPppospnvMzVjOnskqucsDHPfTHbhqFsJZM
+7F2t9QxY1g6ptXowdVWlizKmbpWU3/pNPRzcOsZJHDDH7XDpvF1Wss72CQLj4i/
pYCjg85S848V8+HLm//moF6Ri953lkBBn7d3rrFkn89mj0hP8eyaL8sxw7bJqIc2
Ed5BdqadgnO5kiw8h0weUthfKOPZshmjTz9EkW0kx3lS8CtM2e6Jf+SeoshjhOtl
gziZvyoKCV9Y26+wbZJSgc96e7LVFKasJmHRp+juKw/juNfTcWdVIgUIqWnLwAzi
rNXNbzLK3nJNLXDlwPu3z1ZNh53RiAiqrz04xkpcpxjyzFWpnZbDD/4i+lIIm8Te
ITvGUpW8unQCpzLsDgoiRiWLqE3qTbfqyLITDEsntfXUXr0FZbLXz2NyfagAWpMq
l6mxUy7uKEfD/sesHwZWPioKRjcL56vwG17JAhQW51b6Hux/VZyo0WMMvodUK9+e
nVhKgejIRPFOEYiLyoegYqvUcHulO2d1WkDXSPUO/JMJohE2misdOxL5a/x5h42W
b+8CCUF9VdDeQ/89LJSQPFnuvfUrRTuNC9haigF1yFNPR3DHtDwWF2DbEJ8tgrey
0FzL56Z5Zle7/RJ0Dz6brW7J7PkVr22ZDTNE0L28K2ng7tB8Rsu05YQG574Vc+EX
LXqAZRhMuq1fkFGiUfE1lDrB6NoFjXTPp1nd5X6t8I+nce4BbdFSGJGZjus2UJ2q
YcVAvuMdMa0EuqmiriDlPTcysfQfl97K/DizIQn9OlgKm0esVLxLB1VDG1Kwc07F
aRq414vpK//irCEgw8+VFvI39jR0MKeIIVGMpVpa9BsZCpKPehpZMjd8vyJLXHHb
fa3QkszIcsUMgjPdn6mx5rX1B30UHRLdbBgm3YtAF2VrKWtWYodQOWyTS+yoKU9L
xTy7jq+9zw+BIVRoFXEmxJk8hnwcLoIFFvnw08qrQrhUoHD6M7TRssuxU5ghyBvJ
KcooxRFndFbz1dgbWfjPQ6rAoO+UTFZvZfCy031som8DXGRR/tPddDvkTll+pzrv
4oKO+5zu/8f+uztzpXZ2POTHouySObUIvviPEcWUf8tDDkw8+NnXjb9zFw0O3l8k
VeIZbzCvCBVVgP6vvIecMvcTrRXDIQey2dB0hjW6+rJCnECy2lYXdEcPGrf2dhml
QixRZRrADa7T2ciQszUdgOsCl9rMnjXCNv3rBVZapR3yyvwoSl5CzgMO4nX9Xgpx
DTDQUFousi7NBLYIy7nhDycMH7MLuBlZUIByYjdJSdhJhjaYI1mRuH/Ic4D3f2M4
DLXnDBinXyhCT2xL40Eu+RVU0F1PssxnRUm7s/0k7p7+AnGzujzq12ho59zC5fmw
/el5/KeL+MjGCXBnlgyAKv5j/zf2CMZn0yA4+kVOyIoazcOi/ehj/zaqMhQg690J
dcj4IcjD1ET6W7oocth6TFi7stxEuFS/2VMtCUL1R8cGc5lr0RGb3WPjwgtrp+/D
vHkzfK3UdIcM50eLmBkE8hrK2pV+qaFK8/o6kF7HztzWITP/gp/EohK8nkqxdBU6
oDj2S9nf44fh1JmYniJKwJKnL06EowqqxPoq7r3ktOXeO7YtVLQhqcoC3tSuq+n6
lNE/YBrCHyANhKmHcQ6u3MmXkNPnGrgtM5fDGDL/O+yT6aQn4rO87RabEkOCABww
US5Ayup8IYYV3b+fgpQUIZzqavcRoF+NBqpvBp8rst85QBAOf4xNrm2/uqF5n/Zh
JKVpSEwvLeFhT+G1IfwCwjuhLQpv3erEdQq1e7b4GVzYj6hpcP4JOteup7Y5MHAi
alROQXAdkyAAHlQga32aCrEhB1dtxmjZy7QV9CXE0fOrEXiXj3rB3eipk33LLkDQ
vB+ASevvQfyHEySYZC4hq1a3aEsj1J9fR/3s5aKGZE7f9LKY1keL9eX1/uBdi5G/
LRAN2gFq1sxIcDSG3sAqkVLXUr9NnzWk9XrqPn3Y+NcRljSjlRue4wljrARkPF+o
ANnITxf/1smF6J8iW9XNTgVfqOc3Y5bnTC/Rf+QrS8RcYC6cimQ72MLcKZ61EaPS
MItnbqg4rHV+4jm43F036UzgsbDMdxnuKgMggNjn6VfyCepNs2YE/38tyYEvuYfa
7vfzG37uSZeTvKsoFyXjzKNcf0TB8nVjpI/595vu3lZzX7rspbIMvtA2oN9AM4/l
YWKIoMhhHE0UpdM8GYkp3uU3eN5NWpgedebGvb4yxgO3dUeWPxc9kcGLMSCkaSUd
vYCuw4GYRtX5qIU6IOQCanVgK40Dl5k9yfXST7OQvpVJTmdPAo1saH/gOTKsIiGO
CeJvdCejJ9X0m8O6Fov2x7x5EWY8PgtBoA3JVYhmU6klwH2uSOm0FuxlhFIbqHuo
w5aKvh3pQz44PdEaVghc+5LO1mG0xD5mJlXS5N+3PR+i5a9H3+3o2cmb5oCqZ9Yd
wY6EyRmqsRMefjSdjNdlxKPAvYZ+JrO7OU2M59NoE7mQkRL32WyUGNxF4XQAMbKc
Pw8thT+bnel4RnzbRYsMO1OPTWqkPgfIzS3nLcSFlU3UOihGJPn9wdMB6LtGwKlZ
Gfzp3JWSz7tPNMGnF0GtYM1vsIWdH7K3oKrcd7/65UH/qCisIKjF8Sp2u7h4I3bG
F1BRBXuvI5gXJ/5SbpTOUm39vFEjzNEh6X1cmuQA/q7gHYXPrPpHDZTBzEh/EUg3
w0yGmtqqXruCGhZEuXt5LRwyNjbb1kqVkyH1PQqyGcfzFFX3CK5wNlOynfhREver
xptNmXEopzR1xQyswFU1wAx57h0BO7vZwX/uhnzyGxnf2MgAn+xPHnAq1MxteEnD
nqXaFIYwzZp8TAwTi2csBjhAu4bB8VZHVI4Y8whBln/72FrqvJfJCwzq5Fut/etO
90kDHmHYtH8iULIbCucVchdGFmJ1cTKKoqCrnDyIB5LRW/9k5/Y9/4uRG5gGGQI0
yoLaOU3+RpbLZaDDcWv7FtoOE5bX2q4lvdau7XQx4GJNfzmTQWwk1OfJjVs3IYrK
OyHkwtsNc9UIxgXGXiAWJfh1XMftnQ+Kx78eb0DtNtJnfepUsRGvzdkORb7mEZ6O
mNyFENOu4JT1f3mwVeTMXAAfopBuOn2tR0SkwsrxGK1iMwjFPDWi+JMA1eJJQsFZ
dmJ/6VaqYSo4n1vIlLq8eS1Moiablc1TsPCpPGj868SqbJh13+VRJkC8m5XkM9Nu
gZTolGznCuoy96Eg+OJT2R8+vF1xaGlV5bDNcN/nxz4S3FH3TpvjbxQYnEYOvvrC
Oj82YrlJcJwg2VKvOLe7T42HYKJYe7cAsPg5ObRjjEoPaRIWSiuY85YuSTA5Zxay
SZR0osWJ3t6bZsxq5/UF/PIgSQ9C3fgT1MgrnL1k6CfmddHMN5jwGAEQR0Z+3L9n
S8DE9VXpSHmqcemZoGFmOlhw8lpSTtKSHOqDoxp5e7uXFJHxMqXLJ0y/aXYF9HvN
mN2z4dI3HF96vdogz2+bOIBFNK8/4TMUXeuyl9ih+BNr4FbGO3j3yCunFlndSB/u
YSEe6AA5PPb8Kxd9D3gvcRDhwWIxViMnwIjShjx+NI/bF8iyRknOLc5YKry3OeKT
NbTxT0z1FB4hLOGjSUn2oHvsHaSP7u456izkWt8GBTp855hyKZpqkulDMelGiSFz
IMquOtHKyzznHTG+JeHs3DNq9FNjpEm1Y1Cpj+geJo5Zeldk4j9v4+Tx/nGynCB9
cPAzizN12bYWF84bqnJnOYNlxqpOieLAxRHUltyfVe4GKdxbM9d0eLAkoewGWFFN
Ikh7sedrHZ541jmW48hFAd5ZCaxHmcIVdsSOANGCNgvfqHJ3NhQuHkyeARnNMlu9
fzNTwiujIzwUDk3nhK7GkCp1KIVBuWyGgv4Y2tgBe9eZLg0mJYfv0SJC5trYHAAg
5GHkfLSwEPBt3KnI87fUN3Hc/eQH/byLzrdSG6WGkgiCC568j9uwbO1oUsOQ+u3F
edoNCaBCZJ7fdaXKgv2Dj0LCGTBf6w/PWCCzbweW0BdUaS8RDzuMeuBKeojk9qtJ
uUqr3LgtwVqVa7Mc8ZA3+AFCUxl18IUqSIq0wlhXtMyAi8na3SdLAmnEN4SGmTT8
wZ45OsaJJGuxCx9uZYHqw4xZwQuyM6bRPzXk8zA/SFMHCbhBns/GncCBC4cpdVc0
3cO5xcGh9WauqLcPfcJ0A6845KkQp7mRew0CwTwv4zUjFrNMlO21Bfk+y61nhVyS
fDkU8t5OlxH6RxpZuNzlKxKgBwnASzED6KbNtBF/TVILx/5ZeRGVoScWLHuOMNjW
ONt1/Fn3EgMlDGhy8/TaVx1ox1uNZHyM1FQk8pkm+sxeCe8RmtwS/++IDqZ+OE8x
UvYelby7+gxNwLfJeWa1W4ddg55CjKWHJyc0+OoUe3vqykTWLRo4CywA+1zrvWiI
PX03jh1MA5cu+P5vWWmazHWPXlOm5Bnr3zD0r/4jw+IjML8vVopxtzADm4C0AIn+
0DZiUadSZFYdB7rrlzNfUBbETteIEcnFm0cOOXa0ARNvj7m7w/7ntuRCymviWyPt
nmx9N5ewqTLT3+7q3pfP1sc/Mkw8uSoulOLLbjh31AiSle7ZHE+75sE7DANWj4mr
lPuhTEghNpLY2FyozXqpJXk+LaXKS4dnwWjrmO3050YqyEfx9oywfNlQqdfiJnb2
iWsM16+/Tc6mvc5GGV/D9Q3roJW35LJOSUNq3O/GmfPCY34qYph95EABtHTEUQFp
w5IPAsViwA52X1k8Bw/NrNWwqeJRF+EGoV+JgQ8IDwQDkvtmJvhk52fasY8UaVFB
XPG+ZmX+ZG68FoYLZMVy1LdU4jMHBc/STknnyAgd8hQ1Wp7qaZ6nnNdukwKp7rfT
JY52zmeSdRtGQBTBIfz3eI/TpvSio2788PyGPYz6bdofgAuS11WJjwkNFBuyv5y8
5mR1DeVsy915OULVR3RLp4oa+T2rbd2dNG6O/uwS/rSFKbhOJ1ft8TIOSYmAmsp4
rS/FcmaQP8SjM0ZKEVa+OBxe5K+ZBjdJZluNGmMukFQ+wcg/M7BEGdRAwD9PxMb9
hH2h4uyKet5lQhVaHURYsAK2mWVTw+IQxlgOm+iQ44DKfquQpPjsFYQp2lTLUiGi
1GvXFtYUSGo4WVimzOKeysX7gbclQY+7QesXX+SKux2dnwcnNT8m1GrK7xzIP57G
E1CoLBL8WWcKEcYaq+qAzgGJOgINOdBE8r5Hm0npDxR34bIKC9dtWLiUfFXe7Lz2
bsOwYeJAYrFTPpgwcbQajm7feh0oHF2T/A9f62qReq549/uWps9ARPYvs8pMRcou
3/ZsXbFgzdBeQFe7a7y0TbalgYHjol8X7ux3usOfrRADg9IuHZ0JN9+3n19cYptE
i7OXEwncgNIgsv5sOVIWL456I/tZZKdi1MQtmU2M7GPZGcLlDRl7VXqnOOG9MwDV
tKml0RfR2y/iBnSkT4gXAjTKTNjHfpk3RVzueJSUodEI+GDHU4kUV82asSGFmb5N
/2Q7UAzenK9KiZ9RMmZfAafETyxENb+ygOqUngWIcbJ7U1LxnXG/TzzdHX4cfEMg
Wrn74CNAf3cl6p8U9Rm0hp+aiM+CVruD6QhT6r1dKh8xLb9UB/6s9HahsQQ0wUo3
165XqZzT/FowJ4IiqMT9xl7HSNXDREyqoV77Vpy4T1GGja4o+ozz8kkxrR7G3VjP
R93WbA0f6q3HVdkfxUQJYD51uA+cvixcyt48L9thwsLUi0HNAm49EzfgH6aWE2XP
unQ54woh1hz6GbLZIDoBdhqD8tFOJJLFarA0p458B9a7+1x+MVpnp7c7ij3YtvxS
pvlP+UP2bJZpw3f2NuXDHrlu3qlUF2BnM3fkQMeaCSuKGfnKkXUJIryHLlktxepn
602df7PFQIubS4CVpdZ0KSd/bt6EqTokHheUIc2ReMfOnMa2hplXwJZYVvpGRVm8
u3af3Xc7ww/vDTfPoAlXAO8iO7JLV1XHHpO/zafuTAuhhFB9WOtoAbETzxgwZGCT
RccNRUX4wgUmwPUeZmSCaxrZREr+W/5YKf5vB8LMmxaEAmkQ4v6FvXh/kvXHsqb1
yWR30CW3i6z3cww0LfybVmsgnTLUI2XkriXCGpy549yM8K+vdwOX+O+WLGyjSjvx
UCUJjNu0LiOzuw18zcISAx8wv1nxJE8uPm8Pyujy8jI+yOaIOHTZevu12QP7Y+vo
Lej+5ByzGKDHJgWoLnsvswrD3XOyK6O4CEu/GaTBYcqH2UMmrgdZkRlqPcOhnUqp
T5DIPIRm6YYMDn1ZKcDf8tPNn6hqKAoY1SJze88CQsKPgBFhGZ764eqqtYvYTxiq
posqgZYxJ8yaBAjE1VwNcZV1nnwb8ppopp0DJdeh/DLfHCPfNoJ1VKcvB+sLulRD
j4ipQVj/fdLlTtlxkivfV89rXVm5Z6m8X5ijHdLjhW3D+2sFMADtR/PggyDQxSUe
k9EhhM3PqR1jUbT2dVRcvgZx1RFr7+pY7X5Bz+E793sE0EW7CJrR+DpmhiZMjbrv
+w9Ni7EJq9bANSh5ci1NrtGP2nZ7+hKqUcc5Kx4Fs8vjcV6841i+i8dQNgnIQ/nL
xAMj60arbOddayKRNNlITai8Fw/f08SiizZRMvVE3EsFDcP2NNQGk9Rmq0QCMeSk
Jk3yWGI+7dXvUFvK8KCGRTDR1GE0RgToN6UgNhG2NZCEAJOxChjpoce4en7fUs5W
+4iWNjA8ypZAZE0HODpvEwCYqeqs1h16GGwQ1BaP76eujF2PmLEYxV9k+Ah8ekER
dynrEa5Tt57Qy6rWrJkTy+JJvRmSxQ/f9nPc8FBQxapyIX+Y6jr5fh44JBBnKeBr
uXYFIHCc+rManej78j/vjcrTAVihMFEX0N6/HtDcKzK1qKU2CBHtakAmerROedGO
9B4H8pGGFpAerjkqvpyVeMejZeuGdBIMzoFOm9ENBgdSwm6S7XCK+wjYh+l57yxP
of18ujWzyerg47JygGO00VRux3JD7aTJ5Ax2CUcTYDwLwsUnlhR156xGnG2D+y/8
+OE8rPrV5k28d01BmXq8fX/VDPbi3UynmEPyaV2dp7ybQQe3dVnAYSGfjfkScn71
Mig60LAYnees95XUWmz+V2Ieo8AVuKC8EZwbRb4OsXvyZhdIb9aS2uEo79LazAra
SvDKMs2PgfdI+fI+NsVRSl/Jte8wmSaB7g2F5Pd0tcKySU8q9fl0HJXDJ4sWWNuC
P+qS3A1+WVaneN3uTyW7akdjw/0DVRyYdHoD2NxYE4G+B1bYUTqrKf5WjFnPsZf7
QSc0niyM24yrJYsTkUgVIINr7hhUC6RZJewMIN7B4DAPoxuZ3biBR4c/04hS0Y52
QR5tmhowPE3O+37PHsCmi5IaNmg04dzwIe15XsJm0LgGGHCovTt4tRltwv8ZHj0x
KmtDZgjkuTYqlHsrypS2/VAxfu0ws2t9ThQO4CRvzk9Eigslezg4KuXoucNiXoGM
4BRddztv0q6mheCQ8Bmqm4Jisetoi5Tt7mWS9pSVArBchZ2eB4SmGcsBDzpD2aPc
LnX26MHVr/8Xn6/AfzYVLIIkaRKJZRL98xfLIgtQpAXzvNHb2102pdcL9l5SrICa
udcIC2aeuKyb/ti6JyrQ9NVa+BVUAuquMQoXDAapIHqJnv1nMGVm2jG3fF4LkEV7
at443omIUqoADhfQ84UNl93r1iwzQT79OZNeNzDEUK7qvwW0Ns3YqULTLsmahnQG
MezaOm0w5aszO1bLt2K8jaLL2i7ZXMQhO2MInHSTAp9g9MwH2ohzAp+e5DG6NDPT
C+4H6+OW/0RUMS1gMJnG5qkTbPOrNCUwCzhnoUeY113tePkU/YXAJ9n3BXNlZPuO
3U7YTz99k1f8N+b3rPyoC+7tDoCfUkhznO8y55yS49XduCp9NKoe+3wsPLRGRY3j
JlhFSpfiF/kncbvXQbcdstGUvVIu4Vs48ZAoldycOB3FTkv7Tn0WGBFGVZ9kdeGl
SEyNDqAn0zwAqnF+rC+IxhAE+bH4mukO0OKSmg9dkbqUV7kr0Y4UobXppi9na6CD
AZgC3OFX+Vy7UBKDYTgw9UlEGYK2n3sOnLxE+pCHBf2/ih84BIbqHDeUpzYFaY9+
TkRved8KgIBgt47RnO3mOhRaQCFdluo4OFn1v2TBN/3O7GrnWWxx6s6o01kiiLsR
K5NaTIgrGul8T0p9nfbcQUNZBnxvZGlQaDUmOfQmue9zmmpvRjQEr9YriOKXBDVc
oCvixMyp9rmfSL+djI31qYThE9zgYo9uWYWSvwC1k2tX2BXPyS1qYg4kBTsmd9I0
DqEDDaJmimPRImvgX0iJedLRmdNOsSZpLnAEqS/DenIf1bAsDKepkIq/F/VwgJiO
WtoSpbHd5TClFeViw4HpsJIUdxGf2wHaU+/zolymBRwTF9N9mQShEaXXOjeOp5us
5Qz7avyhS2ygbnnQFg6Ceaj9wYV8aL3/dIM0d+mjJIdgShDehWzPmh+qMzziCG4j
1LNTbpxARSx11NRn0o3mXW3wwgqRUy36FRnpa3+lUft5WgMU5fa/xtf2kl45/50e
nTokqLk7hbNdjKRCJpRpF7bbP6/XG0R2h6sMkf/OpFyHFtLqFSAbbeSWITtUgICG
Jf1yTp9mA9xe6l94hjRcpRiNvsvYzHL9GKTSrZzpfoVvnub1nbL6oJVDnbKwOFJ1
talAjM4tDBd0xL3t9uaUD+f+LJEj5fIIv3lVcD+sGoTysFBFwK3YbvWMqW/beBQJ
gn9Szpr9ygX5JsyjzZRs4hI8mB9G2xyiy32plesq5DTuqDNnFnwpqzEPDyDNhOkZ
pWvPveJXHcLGOKlp6i/jfPboVxtr6H2znVxp45uUH31LHl+MM71n2OT1DQWgoruQ
o9ptyN3z8Rjn7Of55PNn+FbOKF7mm3vQ/Fbr0+eQDQ1+E9u8N7ZQD+eIl/u1Ujoq
eZzdBVwFIa0je9Sa+gHQ2qVks9ET6u1UWBsgnjlC0M2Ji/DR9aLldCqX9dJ2NjOM
p88LiC0nyA0G2hj0NC3dwyCygHYNoHSsFoQXl/MEJ11pvodi1fSlkumXqmBvmM90
AZiUM3pZc/euoeKTmImhXxjHBv4s/F0P3zOCJ0b8KJJw6Wp4+ebDwaCs2fIkXm33
vXwodqNQUcuDOYkAIDdE1iQeDAEFxKVPBEn0GvZhJkdMJhFY/V6XIeKxnI0gsBOD
NDOo90OKh27JwgT5Jemj158XapqN+b4eGKEOP1vJEM+P8d10D+UvAmH6L5v9x6Te
J2AtPrwDTQ3DZM9sqaTMmAJvlYycNPUJ1LnfghAxR706HPmjZFnjeIf9CEbS5irt
+6O1v3Cx7TD/qONoWZDbj9ZbUJED+peHabKEQfYmoQLNvqLceSbnJdxjA58PwqfB
gmOcIbBzjDWNL0YN3jI4QpBBX3budjk4oBXtneezj9mxfHZve/OdK0iYI/6p4OQI
7e+i5kIGRkm+wdn9TzvlbdG2bxv9lvF8gz+7fWhMD3zYwWgjSDPy3p5q29HcmIT8
Ys2REx1Xx4IsGxK9/ialSH26V3ios8BPnw/q7MbUvC8ugTtBbulbKyDSyh2u+QjS
xVxep7dZ/5QWeWW6nvF+IG7Ogqu/IvMeo1KSWqYlxnQvS+utISn47I3BmwJSz1Oj
Pn33vhDNMSQatI7SejwnxtAwwDTUTVoIBAnscSjztJ6W1FgEO79jUYMz5GQvkCtY
M2TcXJSoSZVtn8n3y2tm+i7UpP3htwg5VjPVNfAkNC3knBdAmvAnIXCbLwlsOpIc
saz6pzucYbc4Jzq5qyqH7WbrbdLHfsT50mlIUs9XjKAdWaBIYtMLz4FqhDf3lDwg
4sx9BTGIo9J61VpUy2AdD7jdklpeBSR3nI5uoB5Ab0pfnN42Wq9Uzq61QUMTnCP6
cdtk9m1CBN5NSS9W1+5Qd+Bubfyf9UR/+OyVF3xSgLwfNDIN0Zrkb3N7gHNOsEPz
Xt7a3jh3cwtpvcEdmxtEsDQEuQehQONXYjvN593u9K/qoAgsqFM70QF5R1/plUG+
eeb56gBF8E7by5/oi7UT4oUeokUdGnvkDx3s1MQ64txmeWhJVGvPhLBbz0T2ro3U
SJzAl05tWBfgxPuFUi1Kgy7BmwEf76aZy+X+Txs+ASUs0+IgRgKbBXd5dye5T+Pa
6cinfd9JiMuW8ZvjeayBXt0K8UChpClYgtCcaUzTFA0Qv+aJUAob+WspnRDcbOHM
QWP27DrNmhY6E83pfGWlRyoWuDo9H1DQibuBa5p7eEvN7aOd7UMzHokK98l1FhY4
rLUBc04THwleuGVkU7cWftqz5gZVlK31LvxwkxqbGlOTAHVIrUG0GvLZnblcNfl5
JNa4wZQ3+cqbYmyhCN/i5eRBuQjxqiEVbn2ncS6xI0TLJrAbzossbmsnCylukhe4
1ECj9N7VBUMEtI9mPTS5KRmrfpydbFBy7dDhlEy8SrXcqVCNRqf7pgnFgYHR7qcx
Q9cVNT42AFYfb0nFC3BmQFxtmsFpugqIkxxCzVi2dpeZJK62FKqDiuLi6+thb/ON
5+VAhXyeOIwNd1+npjwn/WFkD8M7kmArhm2LM2hYZj1x4l5+B1UJDbKHs2FuFPb9
hUoMjGS0wo/GclM4kMZmD8FeGQnOHvvOqLIk43g9RLqYXY84mtgrffRhdrldNxsk
a30RS/AXc9KjgDcUOEZeCZ2sbCN/8WKS+47EjZzLXapWlIrZtfe0TdkOuTitXsM6
XgkiByEvbXclzrPVhoc2XlJINgUOdMysZvy0Xd2zIrV1Vn/F4kc5uW9LStWwFH3a
LS8kLBSOq8Cd4wR3S2wXJfMZ+sOz3wdqVw6uTWoB/rgB5WDuW4yLCbi1K/7Gu6GZ
9vSjiQY/9hYQxh5wDdnxT5k3qtTxYSr+76NzFQaHkRBIou5G1C5HtbadC2b6y+v+
wJ0qW49Dh/MJjccCOZHTH5s2yOiwOt86OcA63dc2PYLsf3D7PQNh36xzYqjftUtu
ZTmaQwBZyOTgf/Rh38Sz8Jd3Jv7Xv7Q9kZur047bDAJp2xK6oe5t9xHSmKw3hnkA
ojBicaNZVBVLLK86Dm6h/2KgqeBLE5pe9A09PGOsZGSCufBUWNTF2EXfwIqVebcL
NoCAH/lCNSiTprHZHdMqjDbFcGEy0dWu2XZYToOGEUkULepBtw1oYiM63bGqipxx
cWhNoSmWZY4IcWkN1kJ66D3RpIyaGyEx6cd6Rs2iPM+OynhgRNDiEKVMWzJQpCu+
6dzX423aSYet5E5bj9uhby6XzOquqtmsnNBZ32iRCD1D9+t5Iq4vTULJo9wTol2Z
RNfX9T3amB7bUhAkvR4vDvPvUMvejvbMDuEn3MpB8PKetDQFbLSbgGFpHH92DiJi
BEOskApBgBRuQod6tqTLq/d3N3xOXjR2WoO1XGDJh0/IXSnv5ibEFzETzra4xnNw
bNX2uZB9UIC1VPUwVEcxiEjbVboDXXimTn+4d5tMhM7IaVTZY+B6d7aPxMJGpG04
IKXgUIjM4IEaQK44PjvhHkmM0TjJZtxAkVCfSz/GBwd4Nd5FYJaN/vDKV7pHHjq3
vEFtfDtrwSCHt4S5iCAt+ZdyoBqhJr0Z4l/rZszFYXPRBz83OfvanX7/LqVxdl2Q
6xHqcadANdpOKhDZB4cFOoayaAKnWZvhXrwe/NSMPKkCcorQY/erH3Uw5XVevfD8
uhRTHUABota7rl24WMNveo0CB4NVfFpvqwFChcT9eNNGRkz/djaJ2RRO316i7/Jk
yJx09nVgP8y+x9A35e7GFwS9/4oL7B21NT1jc6ep30u/6ET/JwRTkLCIRv5o0eal
UDQtDR4UfCwqdcbyhSsXUo3aWAEYPS7NmKI5zkDA/fgC/gyw8wctMT2htYEAN2vg
de4YJLvIyw+ym7gXvAEIlMsS+x8PziuB/Pnr2x3za2i+ihjuEF6+nisg4uAz2vcs
8bwXFneREBeFlcnfb6g0ovSXRmn6b9ciEfGOO+p4CC7/UYQfciz6+qyE3lPXHjxE
Eiov8ud5l7Abq6Ehbz0AhBZdx9J8H4T+RltFow/rp7bnqQmBzR8Q15mOZ9O45XPH
5agzPLvJFzaEcOZCmMjhA6WEW4lEJgQ6Yvxw7mQz6vvQ6XOvRBoNrn5/ufYilZy5
XiineSv3IuPr9LGMP3uLbcAEjJy5aqqPJSPmcUfpD4fDBL/EEDRN8AOeXU8OjkiQ
BvIPsA0uojDWTPsdPehYHFHx4hFXioHdn/1qoinwcbfwHzt/H5xCftxx37uALF1O
O+OjEg1ZszmBQm7C7MTIPxZu6AB+8F/iqaKmB16p1xsmDHMzLcxyamYpi0dRIm6u
A7mdXuJxqgFcKh8ket6GryrgULxwlrysbeWk0ccCcAbp44WuFe5G6bqXggO/zVSd
C5QYqcnGZrzwJdyN/cZK7fD3LgNShfeeyUhXABJpTZ5ZRZNWvyvfhYFNWoQW2jAU
EhfBnh15GJ2gxT6k3xgrxZ1tSunsltulDuBn4zjb7mBS1YktzgFMwI1Rt6TITaRW
KldIiQMP9hClRRGhjAgAb8ajHXK+PfDELglKhEpTnlozRgJvLW6Zs8dHXBXtyJBJ
D8onQ+9Wb1GjD1+L21lfxOrCBgNiwLdyAKmR8iFnSUOe6wQVaxf1fekqcx1PtKlW
h7Tcn8VGRbY6Lm2J/tkLITt30q2pbVqcSNm6gAu+nT2+X8a2Mh3nyKPvYVcaU/NK
aIsSZ0KTpsLtQoengRop6PdvAaa4b14H2QH3K8CEC3SGJ82kpwvyo6wvEasuJuEq
E1V4WCo9sgucRW1ImdnjoAu0s6DRbkoPHW05/8G/Xorg1oUngfIwsxlkK13EELfP
j8+QBI71SI4Dq3DI4mboTbLdgdVy4ShPGOyeeU78X3c/NIV3z452qtN7KOEYZcto
8hPUPxlGjzN3AlRSs93Qz9HGfqfSJy7SPywOuZFmDc9cikgLgrusc/GR8ErBYDQo
XM7PN7646Kffsg636jvvnmUGChWjRrDSCfr9WDiHaXxELwPe2T+C5hn74Bu3i7fj
Q9EyabrgwG/fcvZF8mF/IJ6NffHSUb+OUwLtovB4REtYSCH1xtqHYHarAf+fX722
5EF1smV/pq8We0mXAi2rxmJ71gycO9fYwKp+fTOkM7O4WpN1AV3sMSfJ3M48EOhC
yF6NmIbR0S4Xt6DKs64Tjwl0KZ/Xs0WaQz8MyOhq6AiOcHskwCS13t4M9AGmGbg1
JrPCxQ9gb2IjXd/3ZaDS6YXPoSQiKi6DAQNYdgj6nXWAA9hOUzUTv2MxdkLhLvnw
hwp/wwmOmr71C3DdwlCWht0fG55uy4n2c7SUtgNcHndtVTTDFHBEZChQQKHFF5Gh
3gSzPQm95rr2c7noqG8yLIFg+ChKQlc1pDN6V+x60F4ND1pgLEMC/ch5QC+9qK8w
t0vWYtNqtUqWdhlM4gVa5nYXSpVrWV/1Gt1ukcJ8KUeaX1HyaerdjTwAlPOwcgpc
COTdED859YDe7NN4HVtzF2yV95uAz+yTpB1A3hvJqjFWejMehgc5rsOo/F5UQq9Q
QDsuz2aNQs1inBvcAcznHlNJ0SJxM2MX2klKw1veGVIp5jtp/fu/hkWEEpEelWEs
/1kiRmsEJw5g+peWhYUHpmvYdpyMmwZPinzlaTNs3Dn14er7AaYZoqs73EwebHP7
nWm+5JgX9KOrTO9/YyuJ7BSeyflTxbwPJUKz0StluyKCcyJzvkyAYcCyBE+SPqWt
+0nzoYRNTUvL5JtAwo3ZuoNpT6eU39sOjGNLfDEaNy3rFKtamJvw2cb42IJ16pdJ
IaDUk9ouA1G9HLjxecT/6t+Jl22N1O5buyYdTymvtoruTd21M45e2t51lihdSUkI
RPyO8XK0AERqeZzsoIdw7bNWxSMSYcSf7ZgUx6ubXVR8lgh9ZsXXJaLKgmGqnk/S
MNDNkJOgNTBb8fbnOJ9MA32ceYSBe2/kT0MTcYF5cYdOIJsMY9s42rZCJE0HnYJs
rAG/qQImMBTjCK1lxDYxGYjgsOwa1WPJInZvESoXzWPTwZ3fLpGk/wsTlfsfjbKG
1gPoXrOiuMJFXgG+HViza66pMy0MH609fwT1Vun9sCcrsuY+1ln7JhcPl14RwRkE
Q5zfxbmoMUmwzFRyDIo4r5Gti2bFxBnUZj5f5gxgAo0rrTp3bBXmIEzSu0uKIYeC
Lve50pAlssbVy/kApzYE1Vr88hexoNLiZD1V3x0bV+lHINDlbhv5F+vPypPByrJl
vAknwtWhBT4nzc1ZGsCsvRgRtiOhluQeAfPVXbeLE1FM7jwBQlfqD3GYB8axfHV/
8VVLiHI9XRRFhCjRmvrUj6/wCl98to1NjSK4sY1kx7wFTg6mwJs7pjTlSZucxPul
9bLcEfNcTDjNRQkmWKQUHphUqPis4GdSMEXw25eEy1Mb/SSMYp1GUy7KPYt7BYNt
iZRbx21Um2ezCt9rEZfBe0WIDeB7AZz5km6IpAoSw0wmhQn98Z0YxYIA/2RPuzKP
gC3Cxae5mwRiHjitvA+GJU3z1I5aQsFFqfC4iERyMqNVqaYnzTpevLcFbIx2HhKb
O/QfB8/OwgqrjPxhTidih3I11yDeEqg4fKq4jgYBw4pbRe9odna8/BNZx8Fqg+qm
PEZsX4gbJ2ieydCxtjAh+U/9i4+aCH1ZiuUHe1v0wLzhr+iA8DpifH+KpZBMlh/D
EJBU8KoidJvMXdVU+ne7eS+bVw1YkYNas08HxlGXLSiClbx4zJmpK+EjCIIY+rvG
/YlWBJlaMEamWXQGhvorq2WxchdJhfOC27rlJho+nLewhY65GOqlFUbIY2JcKhrh
RsHUhMS8AeYsBp/V5p7+ZzbZFtpVbMaSPIgRiG5Fx4PcPf8arh1VeITPCzd7I6iy
bi/UJE5Iw1qoS6n2ZURT2yLqZiwiu5cWkGzzz+P0GwAegslOwxIQ3X7jXTQLgoLd
CIN13FxFwf8hHk2+jNTJsPXnlQANGNf11Rbp58+t/l8Be719iyuE0ntXn3EUSl0w
+nO8zsz6ClfrMWyZ37Bgpd+cCRXquwQiOCPOBTcdKCCsc/7ORLO07BfIb18LA2+2
PYp/KOJreRF/764pSc8wVU8K/1XWhWQY89YmXqnSqruuVrxnuxzON81dMQjAGqBo
xlTRy8ZI8yvCkPSABbK5Tg5OZZSNpSKA46o9Y5FuAg7iHo4vAJocITA8Ux3MoR2+
udWse7SWvyuu8E8+l0AgHBMaDSanc60aKgfkRua5w/0xx5cz3hoqBHO5fYHjFKGN
4DKTdqM2mBmSz9qyI49I/jEMsNZZQ/eWbxMH5OGgkH3UWRpHxBj6mYBmSd+GrstY
NLq7AYfxiHy+OqTOvBjtGQXWUMKXv12aGSDp64ZrD6YTc68HKOMLhjBpVOtX1nv7
a6nQ6gcDx3dMe2T50my8iEYQVJ4EUqDk0t+LGJFH3nsCwG5JKTZOqGkVk6JVryBf
lr8j0FNlfOkQ2lnl0t+j3BdnLazbz6wYufu5inMX8qdDCYf1c4X25iZNZXsNRFdP
Nc4/qCzQrXBecpUeYx0WMP1dDsBgDo6HYpU/njtrRg6r7+TFjxvyWr9Bd1aXV10O
uwqIC4o7+HVw1gsKjYsNwpPUiuhgbEJZQGo/OUB4gSbfYPGCYxNoOPmNAEDMXqzd
ENCHvPhtSE/YI+ASbwIdAH9CT3k08aRDSV6HRVSAEBK7x9FULOLWbKm/eslDlb9E
ttfy1z0Ig6QnSjpXn2V/NYVayYlaXeVdAVP/0TFNX/wwmc4GpxV1Df98/ma5xBiM
X/PaMJx3LJ1b/9Yi14Pysd06T4ZvZ7bfnZ1jTZMpCbA5xhvQv/Wib1DeNa38iJVV
qrO5GuFqzTF5rcAx1Vo5p9tvcf24srSL2Lzs5lNLx8y2FuZdBVGWJZdDtisKs3Qe
pJmM6UT6wqMLXMqPlQ9HAPmlZKiKW5qxkjqXEZmpJRw25nsJnU9J/PopsWOcXOmF
7zI9sZhqWECvT8F+z26OlDNq8usL0si7ZX1tREFvi1OxuZtaBsYiYqplZ/cc35aA
Y8rx8sTQFaDhABvdv/D4CEo+QGpHlVKium+wcg7g0aUFpWnJF+aGzS09D9Aq5WH8
UUenk+FF7QjXs9IYUlD3yaMByLuc7TGsn+zskSmzHgNDOtAAHbVLic5FpBHlYeMF
cic34QFTErYgYM+AN8syDg2Ml1T8gXBRE6XkOuUKETSoz0XI1co7lFuVs60upssU
H4Jwo7l3CuqJLsfnHZzKYP4MxaOAL1/je0b84rbn/pD0+khcYrYReckzVzp+imqy
GgybjLykZXM2idjjCtfLDDb/I1t+wwuxIe3qaOqjIa3oMrcIXfIrdIRCh5ej5m7L
KExdC8f5tihy8ZIu4vhRHi2Nl9g/3KMPdUoFLR/ie+dW5OW2to9tB+UWqLRTy/6y
YcfDbNXo5gX0jkdTYobewfP33h4UrnA+fqahb0HfRus3zDVPO0orrc5GwwCnrrGL
BqNxWFtqXxcgBDsTWZx2avmeP8On1qE9dZlz/P3IqGzqWy3yahbKgbiOtpGJrPYB
yIbXtbwJCfMJX6gGimQU4/dwNgVRMXb/oEimiMfEEBdtXBebiOWx8Cjz8FzBllOa
9MbaU1y60iKEHFg/nd9/kFhs7KbAMZfPEqCP0YYp9fTd74WofwuGLR6UGiJO85K2
9jsp/s/kYRgGKf+Zd29LlgEqagl+QS+M/huZJFxbFNhnSeH2umiDnRb/hka9tXzk
XAZamdbX/Czyt313cj7Vya80rw+f0/vaV0C3DTPHABQkP9f7XBhnJEQ7/ex5EkfY
dPzloTgrk5LuwHYc/R/p8HQOPJCedmWyapHQMw2IS1t8D3UY2YgyMUMp8xwrGJDD
5U8Mxi2C1fNaNiYkaGspplR0qod+fLWtRblO/M2Zade1SNdG9l0q7qX21dWpNL5M
vsN7zkAktQ5x+blViqjvSraNce4EgEXeM3ygg/vt+13XOKmTeNN87toXVcdXpl3N
iYdeavGnyLjSwtwNbP0BvY4ja4KSS/cZIqRwinwvKfEaEqKssAs1sQ87+tzG9JAt
pThv3Hym/XiKCiJHI/SYJU5hcpSo+1i/zSnhFL3Gfnm95w+4hyHNRp8zbHoJAaC8
/ytwQBftZfuPgq+A4eBU7f/eSeyLgXQWdrQIHZaaICWJXSV5DIFuc5435bFO894l
4is1P5f6yCk9POAX129nYQeKDcI2NhghAWOK+KMYRvV0KvCd9StzE4BDsibD2YeN
BLWeeS5LEZsz6sZO+8EUriaavTQrCqocaJl0N//z8CfNQNu301cQQrlOMKBeDkXx
vCbvQ6wU9hfSyenDHrf3HCoaJRaoIl+BGKVT+R8UNjdnLy6NDHaYzcVHKgC/06a1
wrR9V5hNhj+pv4HC+z5w4X/sz59hbvrRJZ6AJFauG8bOspBy3FQXMddat1svHlOI
xi13DO9LTFKONCfoWZMr3hz+zuR7q+2T9ypAXvYc+cP8KaneVzJRZ6E+BgMDZf8e
lDr9YeybWY/0xu/O8RLHsbCjHTbaEDtzjaLoDNHofCXbeghjmaset88MqL3U23KP
nb8gOpw0YLyjkkaPWXneYL8j4OTY6xKfVIVPGED/Zpsr6XlmbR9fjCEzQwrdWm5j
6+axc2jM8P/l5I5uWLdhKuRIBKFxKIO+RKRJlwibksp429njjZNN9GtCPW5vdtPP
pp6O+dLKBY6sB93fF9BEDSUOt0gOO+BzXObnF0Of7o4yP3NNiqjYWL3G31+PxEI4
S2arQrzHTTFQAne56bbB3ZNwA/mTusRhkm02jZj2F0zgBsZe2zpGAC38iA9bnojC
BdcyseNNHb8XWEbkX9BbFjTVaLL/turi32akf4ncP1agVQZCgTmFRDlnh66vDRwq
vNVOPPL2V0+LySi2Eb1L1RCvM9R+/GI2TxgS5meo677nQ0v58ff28oDCa6V7j+b1
dPbs8f7jlCygAp4goLqxOpKg/SlBJD7pWtJx1ECptQ7NH1xmxt6lF+fYcmpff7D7
v1/5Xpe/0r3devNpVfPjyLB7skusDMyEwvzpt+qJI49az895Ww37aVlf2hlqO7qx
gTCLDN6eYd2qWuBgseorhDQ7UoUEDca2wdC8TNMYbRsrkv1U7qJvMoNP2tM4EVTR
sZx8X/NdJQTfyrC5dprGGExKisKeV/6CKDUqIiw6ydijCGYRDAkmGJAw1n/ci6MF
jS04iOhx9VZ9fBLF+a8//5GnCQKLJ32KUGo4YoOzHwn2ToUMX9aPytWBuLqFXK3x
8NflcMGcT0vMd56DIYwAYQ2G+mO0qNDAQoYXaEM7vz5vmolm/8NSqW73hM+pJk6o
9JILzvRNpMzOLzgP/AaD27GS+gGlehpS1WkVno/rhfSXn7g7GmHoVt+zLI7f5OaG
LsXoZGaFpVblNMRB6Rfpqo+XkbkPkEXK1CyG5PMn2q56bl7C2UlRMSkWWxIcBl98
C/ox+8FNzs+QNUgxrFP31zKKWrzujeYJSreYt80G3MzcNY0tV4mVF/KmAWGqeuge
kkNuvOMOu3o+QXoREsBO+qwaHMUgmjI10VpRU6HBFUAOsYWQOOpsLo8MPz+tewwT
uUA3EdC3Qat6NjbZa9A+rWOEP6UCcIyORTW/r+xI+P/4AJB786GsswyG0iwWd8tE
xhQRAkgWqNwoO1RGMTtSP8ksuWCqPJSGFAINzCaYEFiBrI/zeM5Ck5WYl10Nlldx
JSq4pHIBGPFzIiInpbPxVvv2uLkEwfcQfo968EkVWe+tW3KcwVRpG9pxTne90LRW
xfHDFUv3vVfw9Rd8DrOsU+XJ0hN1ngz7R3lAb9tn13ibmTlcEZCE+6Hg7rOHAKUy
TzwuHseanolH39JVj5jI8AHkcNsdqhO8JAlNQizGnk7fydXiF/ct/EHF+a5/8Zr8
mL8Pe+ok44964hshqhKUdWV0y6zfqHSWCtfik3Ow9/AsnTegVaQI9WiQUekyFnJV
XlwZPuk7SGV8X8jW0VPh+lb3DIvbg3tN9bC0Up3gwgS+NTZlO1cey/fX0M0+bAzc
Vr6+GChEUg/U2FADFgtfuxtVX2yoiThtYs69oTPptQ+S9BkBGbflBcujbMOLv3KC
VTk8J7j3motB8GsJlh5B+sJFv1l/VfIr1RgXHo0QPpoAKAFV1YamQqISXW+JQgZo
lNxJS5HeOYWf4Sj2QvsTUZjkwu7ZKb3T7sWumWJtdAaGtAshXD5/3I7LP+Sg40lR
MA/fjWCN7FaGiQ43G7xtP/TDwL5bkjLhUTGvlBHpDPEoR7HgUlsAyCn8XqWhf/X/
gNdjOYdegFeSKl4G66fDX3Eb2TpYpZ50y+wgsSsFo55Kgq6UW60SW7Le+4AYu3x4
uRyxMIlQKOv78asl0m4OhIFbjvuezagoOSvUsnr6BfNyb4nuSlnapGSvc7xEkY+o
HZ8RoEWLeW8K5nfQDGkOlKN0ke+euSqL5TTVBDOWuIfLK27LuGtP89nNowdcYHc0
JOz0cT3eyyWOz4HXAn6mkm1u35pn9c09ilqGLjEdc0wcN/0ALNe4UhkFouHufBbg
/y1wgtbRQMaw/1UVyqniEn2UTrdvT8tYsRguQatBCmyLCup3VJK2nT114hIwnVw/
imzT2wqDxNMg/2aXwlHxxJZ57c/Nz5CLDR18pJucKArGhxkPhO8dujEOSMLwM3fH
99U7ZHcotCvacYfnTdVJJoOxdBEaEXhr1l2PlQyGupO5GfrL3+4knztKQOL/LIdw
a9vmdg07FlZDC9YvFP/ohGyrrseuk4axZbTVK4Y8jyz62yvX6mXSkJTAun/c1LbL
dFQgstn7fXG93hec121FsGK8li2ZbUwnz1MgtZmuuErmuIe05amT3e2C+ydHLVtb
iMZCbefCABsw0K83FcC9qIBXQX7ZXJXrnHgTLyURykEn9Awk3jJYt5tMUIXFAcMB
il3hJOm4DMWfQiuecLHdOUFkS+PSrUpmHQL2uNch+pfaHKdZvErX8uHBRzwQf/7x
7MqGdvtJr/HLR/W8cQgkdpTlJlF9oy0EAqvlrQjLSTMEuN/6y/Vw1KDimg1qpjeY
EfMh0puhJfORXuLJR6HiMyj+yIlWzmbAB+bo5rmP2pKB5tC8rgsBgAcp9YVGXTFv
szBW+2JzzyFFlZBFtJkLJcS3Xlro0iqt6umMXljTVGwcJdrEZZkgR5EHrI4eKrtz
sFSeO6pxlzWTJ23WBYI2++5UrxyRmWVCA0JS05BRFzTNzHyTVDgp0BdICV/47Udu
zwUN8/2iOoJmKOSpg8SJg2FypZPXdTJ8lSsWVuMzVgzYZmzChbNCodKrSrrycbgh
Su6PogR8o9//Px6ws5Ee2JU50M4gHJ520hCGhmP8GSIUqDYIFNuhYGKvigqoUyEy
9xAuzqSOn5p1COLU5iVakAUMVpEHCYE2oI4WnwIJNlUTCIimL+LN78+u3AH4Xv5/
yLns20QEjssmgaTKqI4v+ZxmL7GGPrC2KD1XwyoGMSS3SZpvtTC3oU6aM/gYbxqM
OhYAPVB5xHrABdDDV5sQ5IEJwR6CB/SiA8XuQ/PAqpgD37/LrGJpDizK2hO9vyn0
X2LH+CVG4itNItPKUMalAhyjnvGpcBJfVHEjYODmi+f5n32xQDK/nYhYqJl211Gy
URHysBS7S9qpXmFCe5EBxapVbfLqWVQRWF6+PEcaXYawxVb63zkBRx9ljNejk1Ev
jxomUEXDVGpzV/IsV97PyPh+XoXlY3i1SVhe+q9GSOwJl7dDk1LXtdLJOKsPVWIi
vre8v2kXAN8NQZyC2/ZiXGQ1NtQFPydlSuLM4Kcv5hSaFFR/ABdFR405hYmgenVk
MX3H3AaP8VvRGN056kCn/sYbqmmSInrBPBvaXs+JztkmRohvAUrT0/OgjFhu0wre
s6pq1f4y2IWZtwB3i3d/KwmDCxHLZuCuZPDUmaqyJN7HI44N4O5RKkfJzf2VgYPa
5d2e713kIyVYDM50GZGVRfBI/WuarGAt7nf2eBDGML09e3Ucqrd7/bi5nDd9QVtx
O0992q/gUBQ/xo0yOZhVStjIUacgHw0VQ4cmAePAW8EB/i+fnsV9MbpBXdwXn3tc
+ZW+wuYnZJ+W+wNedx5Gz1Sfo9Pw9j0iPudqS1KPwyKNIhH5djCsypYywj7dcEpG
HVJoSY2k9c+VcM0pnjB7U0Mu9Zu2tjYS/Jb0q1jRmLwExK4tPFb5HbhJfmFCUi/+
+2t5QWpeFIwzN39JwRPWHwecHGAKGalumxbY4IoRnBXcxhTm6Mk1QZRJbhsJP5pd
jKDed5ufbMYghzM9HQrSh3aCB4xhpRYX9zv1+QNAOC/6iWP6C3lqYswOqlk8Irzt
UyJUaxbBNNEq+EBTO9lJXSNB6kS+v9zpmA8oun/izBcVTnA762YsyqYqw4OJTAt9
918rdijsE6ihMPP+o7gEOFrd+QAvN97K4nCCktgfZuKc2dWu6H9loDQLFD72BG/t
wJEE31RHg1kfwr7jTss7Jr19vlHwMIqLMbmOSbj6KMJQaV9obfULjGZya0Nhvbm3
VX5efNB1GV5jLVBvKic+Vo1xRpiqZE2TvxXeaYakos5hw/GYr//Q8DFHAut+j1qG
dOB6v44V71AHFd8o+Fmi+f+k/qfJGNr962DyBJAVwJv2QY39wOqzYA/xSylS/rZL
oZpFtceSNOEuc2INwbnwqohJ7tlhGzmD2dMdpKK1ta+6ZUbo+ia132GkYNufj/ac
nrush/X5YHDupaYhKG8XpMSllw0ohclY8aaLkOq3R0QLZkHUAB1zuRffQmvebGO4
+ChwWITFLEkEZ2h7NJHXkuL5pe6eddEL9DJzrQETRsW6TwdlZzB/HGObPjSZ0vSX
uwg4fiS0ZqeTnTyeX5mMcOJ2H+tX2mKG5nUqUXd5lUedQDjQU+4G8CWElJXvp1l3
lxUdJUNA6/xFY8k8vG3YwqqmZsaLGJuhMcmM/6uZJQkmRgCVs4L1QUF5Jtg8cgqP
aruDe7nh27l1eiQtH7sPOzjtFl2hCIMiBUNCrKX/BD7JTOTp//ba6zbMGM649TdZ
Z66bmElWlVPbnFTjv260KfVupD98tcUjTdjtAyk+spgZTCP8WuSFbM1mRvVZ/Njk
0kxKO6w+k9Luq7rYOtHIUVhrxRfzjTo3w/cjG+zcSXK6m55TI8LLC9a7xCTh77+B
BfMPxcQVOh2hFE0vN0yu1ppKvXrKf5xYBzWB+XDymt2lBM8bkgL3wbFZidL5b1U3
OWBDLgk6DmnQd8dqcBwXMhUMVt7lDcZIZ/+GsOVNSwDm6ms2UGekRZFMvxV5weNu
txOloicCse8zSyC67HCtts3n321SStQpZeuLC8peEDX7nUNdCLs95g7vvCeRAS2e
kU5TK1sPehCbShFEy8I7x1yxI+LvtTtwn5CrrlSs0n2MNbhVxm7tNbRSICFCC6+F
GibwclP/G/J0Fp0N0B8CB0HONrlP5GdtIR32l6xfUOmgO779AHvLU+/08IDevfuy
kFk+UwsQ2BoRh3BZw7DplXmS07EO4zvtM5HwYr8x6K5nJ9dXBrhtSfyids7C6Wna
lV6Kcj2rJ37Dqgi9SZE9F58OFmTBYH+pGGWiQt/ewms63pzXLXXLm8Fl6gswUArZ
G5rfjHRz/qAOHMwAx7WmlUzCpDHR3w7hFhWl8+/hRAPdvMb8Kj9o7SIxbfydvI9T
28gU8P2YYHqpEcMckW/jGGz1H6m2bEfZuTFNvHAkKbfLNc5Lev/Nnd4iDE3jGjTF
ntlQ3eIAGrSLCpdbnMtFdAGNJClgazQGnAeubypKBqxyKwUdpoAgN3R4BiKHiTaz
FCT4nvtAwW5lwpHRYZzHTjUjGEGUYDo8Lck2boaskpk59XhLXRufQkTJt1YlbDw/
pFxhYWfDJxV73CgLnh2pgLUa383GZ68NkKaBw9wPbKCwcIymp1RKQITu4fvHMIwY
8RrWpSqcGxlVmqvw72/DyvkrTAVtY/KsqkoM/uFjxEuAUmvYfFjuUJZVOJCLt0/J
Gja/UnN4Z98QZr7ZguyI/0HjV+si+6TRFUKlnicxiXPTE4OeNhlA5DQkufDGyHyk
qe3XVXcC5deztNHd2Krccr7Cw06amLRwB5XzAa+NTV6e2lRsZreq4mX4IBTCmK3C
btan9fZU4uuEa6vOycBVSGHMIQufZEBKr8ldKH0oaazX7ffSOrS55MkOpLTgx+RV
ML+Fqfu7YPiz0y6ZL08V6oN9YxViIUtgcNc6+O604lkaMSrIFshHHAWjIbtL9ab7
O/GkDW8PGyoA8tHFTiWnJhWHQS2m5jWlTSZru8vzo/cRvpuQX+HAP58N6waj3Lhh
31SKdLTzy4cugZy4Ma7usE0eQ/u/Z7r6smv71ju8BvAcDl222ml9ahBdqJrnUTdz
f1k2B2d10PFqqAhFygZuLkw2CjtvRYlp5Uy1K434+B//i+E/IP+x7Rt6AOdjMLI4
oHx2+NryX7jvzz9sVFDbhbhXAtXn0OnxlQlBueiPzF6uRKcqqwTjgskaUcHM8Zbh
TufCvUeV5Oh9sdGvcrJOjJGQqF6oXS5eCx57DNtd5OUmxFLPrQNOF/HtsZou77Z3
P7HX+STX4xvSJab4Xk2znJPE5eayL+7J5CqPSZ7lO8CS0nJwEf2PfTzXvrPJc14F
6OcqI2wTfppJ40ERgYF9GQk+8WtajNHkQ/youzO3nQKjGcYinygEny9rGg36LooA
5nqK6Ov1UvclIaXfYFXGDHFQCJHgaZ2OWsU6PuzynrFBfXC6iCMErW3qzW8qug48
esMAHc2doUCee7PbPTM2F4pWyecx3Lg3SLF6/Zr4Ti0lCDKKCaPUcRWnhes8NWKG
xVpytA9amLjlHyCxFY3j1d8yzrxUMgIqmcgwsSeZRwJ4UNgEsXy9Zl/ncrODTihw
VPpPyNn+Khbd5ddycoCUFXvmLoKHTUubHtiyS3HL9+e/58lXT5XOW99kFv4KTqiN
4fGurQfxYaIhaA3Rt6o8hYM1ntj/2cPZ9q+qs0FTc6OF8cnNfDhGvo96GHTngeyd
bo7bbYy7hPg6Ja9ovnp5PdKUqc5goGS/Z79wscURzZ5XwVxw7t8OFSttNyHr4tOb
HHXa3i163n2x18FRayJ5n+CyYsLaeSPln/VnOmJSug6Mk84sXQc4asD6lwR5KZdT
v/t9FOZHseqE5yhfJN3acGYYYxbkeLkXuUlvoUJTYil8+Z3WS1F47123rH4KdSPa
FhjSYEgG5ovfG30rxPghklXIigVVKzKgN8L3ZIjsang4iAWEZXGP4nUyoGncb+Aa
7/Pc0Pu1HhjJ7Nulk4uPMxMSrbcFhOYIGAzqkPUmC2ZB6Wcr9Ud03+18l2n8qjCN
VCZMZA7heFq6vtypD0/A5RFJ7xX5w0OIarW8mGCflbDoRgZt2ci4xXO0pHll0DNl
NSAP8SwEk/PDWBw1B4mN+puYU5fvnEF61WhwcPq9nmxDfGW79hwQ62td0hXUPuta
ELLMpXoUlcn/MNMrhV1dpEmHb4tiw+n774TzMiKUIP5tkLSW4Dgv2g6bDwQCLRVO
PMLUyqACQFF5Eo1r98I/0aU2l0EC8mYCoQFllPZ3csaWXrN3Jvg6pOLYE9myM2rC
7YA/H11s7kCKZWiGE57xv26KYVCcI8FAneEvyyff3wsSBQ7cMlHLY1eDCYl21sEb
nhxwfawFMYNfRxbrtjZ9eWA2djPO7GuE/1fSN5YU9Dk5vR2yt3IxWafaehdmVLKD
G26Xyib4kH5NnYZjk+wRKGvUiiaSWbI17ob0c+uL4OvOrne9NBNGKVenALW9puLU
kEanGPTNA+m5gUIw18PMmKyfxir1wxuNWVRodikWR87JruBzqZygV0nZCbPuNsze
F+Hwpfybpj1m2356GSjyirE8VE8rGWK2gHlfCdJXhakR4/DavJ9Uh9fIk3ssjxsn
PR1NdDxBw7Pe5uVXDDN9T2iPnNOarG0aRDud8uCHVgZKAaKHAoAOiK46ihNDQ26v
hqtNGRngKPj3wSG/5144Po+SNobpFpTUs1yAfId+cL40XugVf5Xzhtx3N6tp0Lpy
kRw996rblJ5HL5x6seo68x5ssiP9F3hIuwkIW4V7P01UYlZt5pAiDByaJh3eo6f7
W5UAlpKc/SG3jeZbZMHzJYXncr0eujV6Tu9u4RiLiep1NLTTM2Rx1a5P5vRmaNMs
8Jzl+Bc62R8tpYJLAylKSAIWwvjBKgrjaRpYnphWIO8ePuncd0h4LptVKwQow19k
lq2RNpvU5B5IDAthg5ydH6vC+UoxuBpcv6fGGG4txyRgnjewa0N7Z5uK+OfGTLc4
CEy0+hPdbaQu3jqZb9zvllaqmEZ/wU/Uc+wtb+vducIlakDjhelZNBRvxFaa+QOL
4opaD0ke1edKvA2mpAWlGMkC0R3iuB21yMlLhdOSOLJ0Oai4YEG7ISuFaMrwnqVG
K/2vclrcQfOt0SbOSGEhBgwbOb0yql+zqXoCJ5TCuQyUavdiVTFmJsKGYBNh2b4c
2BRUJLOHa3X3BXUN5B4A6Q1+l8lipNXee21jKIkHhT3H+TUtot6oTsbNny9cc2xg
1E3Qzm3+SARWJZ0bDfxyy7olUIo3jMSOimmt2k2zwTniFUijb7WvRpzuOxTIRGDN
2hvwO9PIKvxmlsDI56NG84qah3m/AzWAa7nCAQ6yxXA7p4NKOhHNHH6roEXTSv9a
N69D909InKB/yzCAm1Te4Y6GooCVf6qGEVC/gLA343ASTeIVUhM0Nuy6mw5Na8Is
f5OmUPtjy9OugJ356WBWT81qkNmJJmKUmThEeSiacqRZNnaUoEKGLpcT2Z2Z2WZy
QWnCYiT4OJ2wnqMagrdzQLmI+wEbo0o5VdLuyf4J2qVsAWKLsb9/Dw57HOWnqEQL
rtxaLfidw+/KoOW1J0HX973czXVBpcT9nVx3IErsdZl3BWJNhUh+NZ0i23Zb9kXN
0TxIKe08usDcuaIOa+AHUdPS+HyE4Zl4oKI9OYvO05blo9XXWSTCI7p/d2RoD8iU
wO0LbAOvnJ5l2uzdWRLdYbe5kBH/xKoAB2YcPpPFB5D54y8GZ0DBftCoGFLVK52+
XyuzTaTvdxlVqRVqpQkKSkFMZ+pfc+yRbqw5env3R8uUpKGwnodXJ8HAotVSgNXH
qoOmUjUZCpaiBAiWvrwjYiDMWPJPokaU0cj7zXJRIw9Jq3S0ELL1hr8Kd07NR/iu
vVdOte7hexNbwSVLluhXjotgj9p34RgeujNglSLgK3sobn5m6c56abGWM/4zmG6V
v1pxCq6Loe8AuM96Yh+02TKKKvDyk+Pxmza7spkj4bnxye2aVw+fMglle1J91tcd
QVx8g3DGf0cx95tLs8GajRaQb1jWL7+iidq6Lth9ffbDZm/s7bHeeET54EPH7RBj
bkksHepqDCPzHU4iG3ZRZE88RAj3v9Hp6A1RQfqzgy/aNqNDHWTJYVEN6lmSnFvr
vjXdTblmOuZTrbM/yyV+C7B2XkB70GcH5Baaobo30tX5AbwcNIH+NVxC5dB9C9dc
WaesOP2xVzErsA60YZy3lCTXSARj01dWiGhS+F6dNyRUnbx8HTjoEG5gQ4UKpS6w
+XnLR8/ZTLUR+eJtXQU6lSkbhyiNms0ymMU55VsTikyebIYb95EdeENR8esZ4QxF
hrLvboNTrD2k3joohI1kRwFDbWAxp3F+tpCKGl1BQzzVBe0TuvWncxQepZnAY31y
cSblsRP1eLdsCDu/VANzJgz2nKcXjPNo+Vodh+xzen3ptoFJQpUcsteIbwIZCFJJ
FuoUj6jQZ7G5sx5bFOHyzulVZmrjR1vgPVTERoRp8kduQSjD3Fx/H/2xkSS/8Nge
dMypH525D+Hoz+GO3iAyeBAl/5yv0n40p44S1twcYsobkfjFHRZUWXG1mCxUpeP0
Hy96Q/6UOEBG2UDo27bQ9oqA0UDPsQ6VxxugtUqh8kFN3MViTPWLNJg76LogejQQ
sUHKeNNLf5WKTQeKhXmAvOxfzkyMaiRg1Eq0ea50VYvONXIlDj1A4+rQ4mLTkWS9
lc9QNxbsS94p1dhZzhstEb0KBvRCilHC2FsNjr+w0gDAf5yyajZ4QnrC+yyI6uHR
geifYDDJYDH2P6FPdrIJ8fRR0/8hekL7V4NHQiv6xPF/neCGTQXZw1IQGO7q45yB
FrDH3XBrleBJcAj8bVgTFA8mxWj6C7tQzfn5inKHcfmR9l3xzfO72L2ULOyiEoq6
CUObJUKkfwuqPWpqC52MlR33P34Xu7I2nSCXvQ3IPvvTz3FE2zEn0jKYKogFZWSW
qIMCaroyLl3+dqy3GBAViheSOloSSO2aZ8q7F+VUX5rP3UmcjjY8G2ngPk5vWTyH
t0NKeazZmZH5lDmFwz/uvoES4HvmKyViYOdWzC4LslvlICrgYEb5JClSB+/6qFI9
rGiOP4w7/cdWE9vzKgik8+/HJKJvbzoJoQZRtxKbur4t4NsV9HYhT2Dwxxo0Kcxl
+GlU/YWI6CDpmHJgTPVEuhIGM/vzRYY6kyxcKLtLO6avUOcy0wShW7do2GJx7pYs
DNbaZ/gGpSESWToEOsrlC5v6gqSGraC5OI42fqyo/2RCdtdOGXRsi94uF53Mycih
Ak/DhBle4+AHIhoLopXmN8v1NE5IJZ0ovP6Edt3tLrxM174g5v80sfhtRTlB3Vk/
nShFh9VLV1igx2uBqTj0J9MT5t2ksvMADHMQ87SsF9o8/QI4f2DNgh46Cw80HATQ
vqTx0d+tg1Vx//7rTTIF+31+qdPvj6zbbnNk12+VMj/mHFBnP1vXgiwO69WVuGuK
0bcsnBnAlTA/GG7/luidT+MX5ZYsrOdwBJAZ73cKL3pTFcVx4uPeXqMAOiVTNULz
YWUDdqaEj3u+Sm211OrwrIG2bVdfsjhvUD6fL/C1MtkC5Q1ExkPg40hTiUubop4x
ipUvFWRcByczU8Pp7hARF4tMWSaU6qwqEPoY9pVFlZmN7k1rFae9Vw5OHfW6gD6F
mPREEwslbCxCCplivbOe7HM/dbSM2DZNTJ1mUYpOGcpbjih/DH+SJS3xVaw+Bz2h
zWCYesNhjyqOodp+zPfuttGNdZFPBamO6u4HK7+43RteCRNuFzPvZb2zd9QmtT9l
78YIARZ+0FBbNdgu+sgahQjD623Y+ExCqnA0SwQCadAUYK2+dYayUQnm6J9GKsb6
dUq4rtfQnYn7zwuPEF4yxyg8LtexRh+bJqoSYpy4/S6lZJM6f+l80ukzlUmqLGIW
+dO2m3gyYt7EC3jKmEsvneT9n9RW4xJXRL8L6p3flo5AyLT6gH496AenXZGnkbCs
kVauFytL2TL+KobNaRSzxMvE++1K9VdjxtPqKL0ECSWHm6gFmwIC651XFwv5+JPL
oGM/8jwfRVBIJPaAynZGjz7sGgOO2NQwZSWagwtmdoXm9RGTahZQbfoFpkrZ8n+x
P/EaXT0rQQI/T5BVDF9VXmZSaJv24U+PgCw76DFMmvlrNDnzazl80Rlz2oubqPFO
mnDbFQmB+Zh4nWHjRltPS4GbaoSqqzPUfZAoQGqNs7V2h5yyCSP5k/aHfsYrhpQJ
ZR3pV9Bl9Jj4prqvsQ3Il8QJZrNTLwHo8ia5H6FaXgMSl3OVOkGOppIEmQ5kDuFR
WopHSSe4k5a7e2ggXE6kVRreL5xiembkFargR2eoRPbFne+LvPmoosBmN6hmg7Ta
uCUYuLDHpOCXMsxlWZx05sZXl10rarwO9gdHT/6D8fBi7rP0sf79weXP8NBXcjhL
NpUaPu/xza+e8sogfFXFrtjtgiHXVqaqHUBfrikMAr/4SSMNgjOKb/qtwafUhZ0w
BZmN+PYlJiWlnqJxwGuqXb2VIyHr/3JqgZlsdprZLA27kTO+mgcGI9rpRzlUOLfW
qN3KxeURPz+55cgZ+KCK7IWEoDeqiDUQQCaRAxh2yd289xVeKBk47IXVusSGsXer
NUmY2pkXO7af3j0zp4Olwqp+Vx6ZW9lUdUYID8uX5Fh0TemGWnZt3f/S77T2xfPW
T68q4T2iT3BBA2otNlQvhNsuMMhsmAM3LuXdjbL0Q78GYOWaWU8b2uva+f7C1K5t
zd7eGbkZDlFcbtN7DChUANroVnwcMGmIvnUiarg2a0XZTGjhKm+5TnWcn2pCL0gy
+jWYFbArE6ulxTiqXIiReNzE2GruW4t0qK6jTMLpqovVVCTO+4yin/PXmWistsvJ
6BPYZHyQPZPIcmVfbA3JUn8zgvPeqhuUYQra1aK0khL1FxHL5LvGTfg3R4n8IfRR
vy2uhAxewqNvIYZcXvC4dg1iI/Mf8gzzmKM0lWpC6Dt67J7sdq5KTY0lWjhXTg4O
GYZ4d0yL/MFuZmAFr4/EuMwgtpIQpgbEpGTmHsUCgvjYBuNX0OYQ3O/c93ocMpaR
MGUm7FhSqw4Q/u1Tg7wL0dOTyYUgE+hRjdUy5ddrj8W2hUg39kxZqHLYMNEukF9g
ihoDicp3BDbQhirYvDmqBnanfFAHIJDH8xVn9w78NFiD4sYGry4UCeuqHoo0n42y
W26utmAxJHhNEmaNfikMF0HX0/HXa2zY3f7Rqkoo93WwwKUsbqXzsmTrdmQNc8zo
+14zpFPAkU9V9Hx5bqwSN7x9z2KT/CQHwPA8UwoXqTsMecJ2AX2+MB05WG3mdums
8TrA5ZPQh1JS8a982EglEiAHF1pMhYoL5Lb6Mc6Ty1WuU5VFXPSajqd7/hAKzqGY
OrTwFeOjjvGBtf1JhOnu+4OLOJz3e+qm8Xs4O+1NP6voSrhSDF3k6THdcIWVtWYY
oW7KdYpNIXidh8ROpsgK3StsuhJVUwlZdZ0ibNoTHP56i3lyrc8hVsdoYj/B2nrU
0L5QswFiVqK/W2c07/Ax9EuRAKYwuHfALBUkIKNKpzVa0DjesNUlfqO9R31Vxvcv
KenQaebe7/YcXCmkpKNNRG9A0ZS+2DgZ8bVxLdzXKi2iJlYGzKYmtKerVicnG97E
LkMmmRvi6SERxRml9auNRrLtSLZHkz2SVpwZy1NN+gPs3rPrYybUOtsIKuaXAVSD
kKnlHKmxd/Nc58BmEiDBg6wZih/SnqWv2nCdfXlhcKSA+Hu+zrWcXJAmxM4reQL5
uCVe0/yK/z2eXV9ASUxHm6g14N1oRBqMRw1DFUTarirjRsUn6MEQcBFFBpNzizvU
d8F16QxmjtUqTHRXbg5px9f0GJax13rARfe70C2EjjrwneZEd9cDxywg7Ytk7676
nAj4nt/kHo4+FPF13q9P/5JEVmRPNx4XWOpDsBdLAm6EEPy68MwIgWO0IsY7iMnf
K+0EqBzJgCjDhB4L9pEl2avMB8OVwU69rdn6VJsH9vNBayg593JZC2d2sTSLiAa5
vtL08hlO/gJ4B/goLNTzRJouZZGa67AtBA/nnyDedStaclWKOsbAz76bvRjgSv/w
oG6mhmjPYSlBWfRYeeegIM8E0RNPKTrOVogpw7tF6xYcFKTeMT6Y4lqVXg7HS5Q8
e4gqleZF9o/RGfeIiwf56wymM7UqoVBEQE4ODQK8Adfj+LuxAG4cyTLOKOdznuhb
FOoFdnL1spVnG9W0boFyfEcPXskuEtwQ0UEUcSF0pKv18x/zCBEW3DjFK2XJec/u
PvbK2uHXs78YKrtJI7lgGkFX+N5UFkpHJKDlWw6BQw4NizuhYo9NZDExd2AiJ4oy
JjoU4YI3qBs3XAfOIc0j5K+ngfoBer7J0mOu18a4DJCKWkMkLp2tBHCwfEd24Gsk
gNSUhUfUQQP/R/rYlsRrepNc/uSVIHY8JzI5Wdoj+u3eQzfr1c3rx4l4uX1V9rqb
oT6BT7nM0FISBsNzqC+DnBAkIQn49RBnqSBfyu/iA1gi0h5ncD3GpGrfRWqaW9D1
qixgp5obJ2+J4VGhuRAAc69nZz6AGYgsU4lOI9TGi1Rq8soP8dTMrHB9xwoc6ysq
ZNVgRAcV4+xWSvBfWQodVbE+toQG71278oDiY9v6DnX7bKXw24Qut6Tt+zgh3Fsz
NrlqqdJ82HPujI9mMfyIPoNfLQlkr1TiSszjUtF8wGK1kNu/fKyHTR8B6BSsCg95
A8c9ngs/VcjU2hrxnw9wIODe6dhJUeya+X5r8zIEw2VA/R2odDNJp9sL9tABAVPk
W5EQeb3BjRPFc9+494KRB4dhqtp7j6denyd/GoI6FHLqF/L7QDCY1LbkMGbaAOs5
YVQ8TazLUlPYNXbwYJjHbZDE3npkXUgs+DPnlATcAhItjSqoA0s7XgA8uMZrIA/T
XTxm3WqQ6yZmyAMgfx7s3qse7kwJa4xtZtwvGorwPW3Zb5DwVwQM97jj2Y+OKcPL
y4hnC+ua6xNlNTGkvd9/9mbOzTVtRcF5ZXAalI76EyZWu3YqfNc2MWpts07WGUbT
+HkznEOb+NrZRjPjcLLyypISMXrO3A/q00rKZPV/GQmDdhfk5gwV8WLXNqsXeF8U
4d9e2Bp0/CfUVq6jQ6QFygjsODlT99iRdPNflaiT0enIwKhF/lL+lcuuMo5ej9C9
tUSg4lM6417B2QRoygT0taPfBvI496WoFLn/uysNxVStDptobn5nOFeztl+B1el5
TZI2meOMu1WBxszY4FMD/hkbah57wi78VA3evgsVtOz7x70uu1MJbSPnDWsfjcIE
1bivLRHHgFtdtyvm7c09EvTXgtcZlp/2U0Fk8kJSe0BbL/tsuNM86JH4vO5olyIi
mLpEHqwx8kGX3makPNGqjEvCudebHJ6lnKJauQ+2Mcr0erbs0WHxdoS6oV2cerrh
2UF6Ta4AlFmzjhfZt6Wu/MVeYkcpouFJ3q6N8PJ1VZGF0SbZEI5DngkuTXc7ZKCr
tvJ5NnVfEWlQpaunckATZvW1TwrNZ5gm0XFMdgDSsBlOuOfCIqbng1OEAl8Gk0p5
q4Lm+UR1l7b7Hiz/x6eC0l5S5z6R79BgkOxH/rsmqHX3PaAXsHAHIXTFyu1YhFt0
omO3ThSbL3IGLWJgRUhJesE3GyvHN7bs67DB+GxtxnA6iQW5wQmzQRbFZBB6Uqvf
5zfW1stzCCTS0oJarayiwcZzeWeiq+ZTklZiszx6UpU0CeRNVd7bj25yj+/MS7wS
im6ueJ8w+7/4B7EYuibVQszsxKRRJIGvZhJK7ejgvdeWCfof16yOC77juaU/fxPs
oBuYmshn9xX9y0Iu/H22DzjJ92DjyyUXgkxFNhlJvenkoc26BXwVI/zK3N0Lrn7w
Nn+0l7p3r91+5SgnqMDVhpeovIfgbLIr7qsWM2TlLbNlAI5njj/ggBvGTOf27bW4
UJI7olmvjEg2xcpG4XKKfvTbpyFRu2ufN0tkVmQJrkMiQCnjX4cnj0KljmgAmMTM
Rqr3dqgRSZVwk2oh5AnuIvfZfoZF96WSrvzKAvTfVV4WUFO6W/iNW7S1kZNQpG+n
7KZ7WiPpK4CvzN0Un8HLOdM+ao5FsXvEM/rOA88voz3f00YLSdNtzwoBWhE7XtPG
MwhRaAVYR49+ta6wJitPda9gkmzqd4GKLqmsy3zK+PnW64kq7ZgxOJuhsl2TZaJE
S979OTrOu7aFIavj6RLd7BGsYAAKC+a/v/p3k12NtGFiCqqOWpW+4Yp+mnm+EBJr
RNAd4xGEqyEXFwwCN1+VeW9JykH8+0+rk7XF3oYbKsE04t6A2p7znC/w/9sqhX3+
zcySQhJPs3V7JcCZkkBBnCUE6ACfHWHOQpzZC66Jss7+hw38nvUpK0JS5D8tZjOg
WhByKUxiPIVE+iHCc5eJhTECCfyGPZSQ77Zmjbse5vHmPNRs8s9QcJ5QwkJd1ak+
N0z2iLiGYdhgQS7K5TmDSUlznOi0uYPK9yFeQufnGItg8NGa7ozUlw4XhnoIx5O/
vjhfn2KM3SPyfjPmtWCfA6qDyphMUpS5eJ3Ykrusr78FfsBkFGYBiPHeiwLybI08
nFKeJA2sp8DP4WnW9dQILXx8Ap6/V5sIPI17HxN6EHsJaFz2DWEWX2KbJwzhe72v
nHZtvIt7NzxQrSUbnNDfiyCOcxlSoE8QAEPFzSCRXmGRWsmvmGbkrql0uQl2Y+i7
sf87NIT9IshmNLUXcqLIy+Q9aTAKGwYqBqek1j5PVBwKYjygCht+/MBhDxNp3Bd6
KPQFkxgScoh1Fvqhkei+GSPzuyjXEvLEeC3zgRSBOp1XanvuzcrzTzmf/hoytpfn
jYRUfFo9WwrpWtUNJB0qqOy5lIJBFXXiKAFnl8LAI0EV6l04LtAo2pPRhJnnEdoD
vs3D+gzsKUwyWwItTtQaFE9cmk0Aqs7lMP/9AehhyIxXYlZEwDO5i7Pgh4iq6WiV
dvhN1VQCIkPF+uEtswJybrxJjkOWlTdsfXhBDN2sD6PVR0kqOwEFRuSvz8akCRlh
FYKpnpsw3h2JVWY7ZcYeYGhg+2ALHlwdD5EyAw1k0cNJ3XoEAswgv9aqQhKP2sVm
cpTk+2xcd5ipLAvaoheqw/Nfvi0x383aa/82RS84r5DPUYk4sTEPKV+RfgFzL0ru
Sorpc8Ajx/ZJVh22p9JR872KY6XVxqUpAACag+SnVux6GjN4ic31oYgBfW05mA8P
8cpF6Qi//u6V4YBufFgiiZ62i+lcU+CVQe2KMHptJyNJqKSkOn7Vq57/PUxySIR5
kQpRx6oFpR4QUXgkeot1GQu2Bxw2yv+E1WMoFewzVegpgqoywMg+x5CI/LznyffX
RW8bzi90BD8+emijj42LcT4UeNtVs1pGnF0VGpDkrkwU4ffvSlV+l6aWXJkULz6Y
0uI8/BDgqKltWBxI3lOGEeOhlTQX60pIvc9wspb0/qrRKngW9YoDxdUul44kVPCA
qobOJqFA808SlJy6OiSf9pDMT5k9StiTs8XqrjbJHu8GOnUm+sX1rjUYPItOt1eq
xAyXSIJf8KTsL3AnFKtflWejrJszAJliVVhj1k1z+BPumouWZhUpY2EEE7gIQ45E
VnYsmvEqxNVu4XWeU73ot2b4OUwB0oPfhEUXt6rU7Vm19hlgDZNs8+Hnlxcr3XU2
RrYc78WOhUO7jOaWYYta5wKQPdOVl/U2L5OjB6QQgPxp3YsBTd4QiUosfhb8Vu9V
eGqGwsfS0Q/XGdOX4YgX/wqzeZ5U3YmuQVLsIeYRS4RUal3wVhucvv42SIC6oMD+
xOkNSYAZx3Ia+rW8db4beww5hFFHy2jWtsDw7CAPQ8p0WcmDdKhgc2z81d7OXQfU
Xw9F8Wb7Bn8rgzEchCkjwVvkfFsC4AQxbJX2fAVw0J2bBVk6iDPSezGTw/frMrQ/
rzmoUeDhsS153ra5T3xLkYp/p83U54aqCCVvj0lJs/uh+mp24HBo7WGzEb7aIGqf
mdLnBxPpI4hrqByUECVQRN0q4bVbHzo2iyoLsTPNMFSUP+jiKw23/3wskUiiiMXW
CR+Qtx4gDogQ004pz3qKiAmITwn5GiuAnI73EOD1awJeHeHmN3Yx9hZD3l4QAQCN
q63J5uypo+6xTB38aAGxYtf7HK6eMf7sJHtbX1ZYy5A8zNU74cd8oM3wYwmfShb8
vOcV7do87zzbhmiJ5d8uOEF8js9fea86Ty0VbPQbW8Iha9sh166s7RQXA00+xzU9
UKoHUqOzeqhvIuuBMl0HQF5aZ2pDYH6VBxHWQs4Dednip+MHgrCfWSXpbeEt5ufJ
Zsxx57ucfX0t0+KkIk7yzYFprmJ0mypdr/S9xbOnAz4ueWR9yAOL1CjiOBqH2s5N
+Yn0Tw6yIhss1CEkuUIXDW3BADbqJ2rK19pklk6pXhULcnSIJ+Q4JQbhyz9cunGl
7dhp9+ppL5M4WIqW9ZLdzbCMspJqUUSPBUdY8tkoMCk5H/4rfnMHLpBv2iKx2aEt
8Tp5BDkSa7OfY9J4EBosQ4zenMa/UDF0K1SmmyAA1HzjDSJpPIGpRykEleJfUC1y
c2DWttwCzWJBrOniC1mpgvV5BmK4osEev4jCG8M8sa+yKJy/jbi676ngXYVC/aVh
/qWzvXxi1Cfs5dtmw/R3ktd1ExnxkFXsEMJ+NOXZPpsDaQQwiH/jnheSEWXXYJij
Y/ctEBF5I6vCm6yiu2+Etfym2FLVp1p/ksrpHDbBfr8CAOKXItnHuf5Bh6HXxPlX
Y63HDDrPftEC23n2dmV7ojIExBt6DrHJnIRxs21Z+CAznMY+14tnoM5e6i2+ZvqG
cSD1pMl6c5PmQKedWSz/Fcg9+XwFT8pbp57mjz1m9/9RwgAfQhRyeAAQPwKzHgvs
q82h/QQE7xBdHuRCi8V+nIG8Y7I0cF0YfykPDzJP1PDHJDDKz2i/s8Xck5fAdGVu
gAYTfsFRRekyr0Lc+bdfLMM6+wVarNb2E9j8ihnDkqLw+6i3bgRwZXtwKIWGGSYa
9CRcKAvD0hzSnp9INmwnYGTfGeiEsc1+zjioTaJYbUyZUyzLlCPwn7EIAUZzQ+/c
flL5Hw4EHM31CNgEjF3uiur1AtxuUqtF1tFvywrqTX1Huz+R+uXQmzXWC9QIbgX6
3uO0aWKVo5z3wYz5tgItAj15WasWtl50fjmWUExlcORtVfrljMNS5DNaDi6cVCrQ
1sd7plzIjDMigiJbThpw2XOTbayVUaiHdKaDPEsq4iN07GWDL19ibpgZEyEBLTiQ
vcBw3/OavUzLPinAxxCuWsIfbW0skoFVfwJcXo90ZNbu98A8JZoKyd1EynvVDC86
KAjljW7p92NYLb1gHxBI65ZSTPMOPh31cl1/9Zb7Q+RY52VzliwhHzOihHMoU866
dzH3eu0ubOwaEX0J7hos2McAs3ACPlaUHzaOHLpIlE7pFJah2s3peO+bYD65dMqV
i2TkbMXq2quv2rxmfSf0aXH8C4Ib34w1De5aiEj0biP2USGawjCF+jHHrPEGM5V5
maKMQ5tb2OvVapomhiX52g/9kE74CWmXpnQY06GSHuCdG04IuwF5O3kkxxoIpxVV
ZwR/05CQfM3J0T8F4zDbbRrK1VmDFbaL8jH4IIQkxW4UHLK4CuJCQc+weijOP6I4
Xfbmv3eL2J/vuw/HoI/6LDV4gI2GnusexEi88dT33IJIcYE4ibd/Ku05u3e2YWqL
s6iyaZl1WMbUTU8vwYrpMCLlXwzWLCxlVoiNpni4xSBrsnXM7pt/AH9jRIbwUrxX
8YKN7pcun2yrjPDQNuOAfuEQc1euNQRi3z/MjXx2/tWy9lCymm0uJPr/kG/xwj/t
qhilenrR6NGShwaWmJn12A1nBHGH8G173X280p5uCHwJDTMBUcUW9b6TnkresvfU
LDK2L+impiQGxrcDDFsy+rMD9l4orCUoAyQUU5ro0TXv6OiPKjBMf0LeSkwEVHyH
2y5cci+sxkVwKhaaCmOZ55uFbkeRtexVbyRcqpN8JM/2dBqvTzyV/eHA9aOKsaY+
5pIxlRiii81lPu8lIHGzovTvgWJuIllgrp0D1kQ6RWN9IYUy57GRvJzXD55gVoRe
JzpqbztpI6OLGjNWteV29SduJdkCYGH5VyroH6UPq7Umtkl11CFP+F+rFE+BpgVZ
N2X8s6l4xftRCYZ3s2Y7w/UUMs/x8HPMPlNc+KKgz39jjfCBEBz3TrlCwgHwej7p
M4VO5FuDXR5+MBncl1LjooIYaV23t++rVKLXf0T2u79ITz5JnLOex1n3WIMOIltU
kIrZc8xcgO9vvBGXb8q/4YTwVGKCScRlzO7LG+S18PFFPfCuZjryx/r+J10isqMu
gjG3uPMGDu0mNF50durmbpxnVDhupTLddyrnDCcS1h8turRXGqnuXKxk/hq+Cnb8
+w4huCx5+XSxxOOkTNXcfPbaJ+HcuGXRLMvHunLyqDjUyAfNaKFgO+4eqJIPKIF5
zLuA2DlvAy1bTRh5cbpO4MgA07HapuwVWp4mDLfC7jOWXxtu4xJHyWnvlfXlsgQP
h8e29M4gqpIIQLh82wLyeaB/UqBxNAwlDUGkg/l/mGSSZdZV3/IPcULfiXQeRLuR
j7Suz3fF60NmqMSJt2PY0jGQxfXbfQIfwz72HeHEHDmTPA0H8vbUFACsy1lL02ad
VWDAU929Yvv8ARZEjyzrZcw0jFSDfyjKHAzSAkG1XjxT0O9x8Ho89o5zeSGqovFP
wo0cbR5Cv3QKqfQQLf+P+cD4GfVacFAiJYG+HdGud327/AJPLZwCO/FWU1RpuewF
eBnPVMeEm7YsIWPZ9CdJx9VWMyyqz11C+cMY8ovTobrswpLDJCwH3JIuJDYtvzE0
QKlcp35u5I3FhcUgwJpVbDqIT4McTL/TVJR5YohZCqc/mPhXNjxJfJTQFuDqR+qk
37a4Nk9LkU85UUzDK1tlPXkymnKuHXIqMwqFu9AyfVOGipoCC/bW6z+YmsGPL/1/
6ETR8arMoxuK+sGLNIP18LWhPnuyY9LypmyuRXdR9DGY6Wg5XZdc2K/PEzy/kcc5
2khXP6RJYhmfJltMMwqtvxLiJrkY1ZmuJeNkfbICIx1hsbBY+8ODC7ywgP1dmD0O
geLsvSnVTtkzEriSpQFN/VJawRRxEoKXzb3W1Ev49XWaFrOmfVVuxH6tFOjOUfpz
hQ0+kifwBN5a3Qt4LbBG/sd5oH34Stn+PiwyRpTHhUX4VS346kBLbofuesZ33HeV
NPKj8yKgljpiZvc3exLlL6KKiIcwOdmw2SamFzC7wHQxjh21W2sGgr/7rc4al2Eu
v0i3qt2oCQhsCvqjY2aGT78SN8dYciHfhGF0O9LIZEOyf4LJoMM1jgH9aHDVWgAm
ZmfyprRV907zgaWwmvvSNsRm7DnSlxupldqQ25eefSvDSqrkdkAZGbvWnhb2F/a9
tES9HCf/wLiKCAKsdOFGeCRIPcVsnqYJch0HlsX5cW3GHM8lORhOhNeD3kMkvz7q
Qyy9+sE3HZN2jpk1M0cCBbUiyX8zB0CHRmfwvWq+BDGiVT229bddmALtRUrZHfnT
5AcVCA/E35KVMZVYc8Si+kCxfMM3g4xO0pvEwgO5ONO/9CnRUJ4AewmCML5NVvKd
oSPtn1c9xgFAxYQKEHzNs//nKJ6sSa/EoUas2TJROvzNaH7Q5McaiL3Ppoq5FouZ
6f6JBfyP8lCmtRk9G8zBv21qoI00OjRMM5WMjcEUGswN7CdMzKgaxHKx8l9npvMv
h/BFtlfVPNZNGTvctOJR/LDy4YQ7NpWANnnnTjpGDDPzrsalAg0MOJ97dpxrrI9m
URnWny8yLQ2dxN6Q7Qd6Irabm6l+ob/Slqw5ZZGqniASg7+YQDNTbvZp/x/klLpP
bj8NsDpWYtH9ESMLVkAiFl0DT8UEMa1S2UX50i4ap+uOX5g+myqEUXP2SuL+icaP
oIvgySG8e7V1Y78hYV7ekLajREriV4+YCTinoNljQU4/C+LHJ1tKMeyUTHhdD5pj
JDEA26q3mvZuPbgg6TBICjnS08IuO5GzTiDnbfdwf9vi+lGvujWAB7IIQsXJK7Gq
+C8OTWKw5Jxq90yzivBJaVy7+2tpnV8r+2stRw0XRniQrWp18A7f+FC8/OuqKHHG
X2sLdrDZqf7sGTEWzkB1aVSC6cFLfTuudvWDzygAbyFMil8eoSqjASFVT/sQ7iIk
yjSnsEQQomdeRbKMSRoSkxwSepwN358Wuqewm4VqORQUo6MvNwv0bNH0UKDHsuXP
s0cHaMBbpEtU/MezWLD0Z8Yv3RsYJAD5Q7l4wfulxvnETxAMh/7x4Vk2cNATnSXg
0ck/WSAj0NfLGHjL/nm6rnGEc38b8CgHH/ndjVR0cm/rb2YKZcJ2wqXVKGTHVzkA
hmO5sVVNd213MFborGMKu+jSku5gKTboNf/MZCnm2ClTTzttfTasPHgJA3dcotrF
CXXU48gqQ+OhsZT7dLQ3fUZr5kYarRMiMQudbeslzN2xC6j1J/DTMexWVGk3c10C
HrxObk4FDjmg7OVv+yeuZGgGXQKmr7I5K3lZrn6T32A9vK557VdOkRQqO9K0UUqE
Olb+6UIeSwclc/24Ljm+Tk3Ltz651PxmMlRZ/lOHOx3JO05qIgSsDEwy1rHvRojs
kRtANIvh6PDxF7a3bItmZs9Wwc37cW2WTfl/6qOeXnMAM3jheLx9xQq8dkxXOVo+
Fpljrojb+rjDvKp1V+GoPosjo3ITO1RkuN55USm1WwhSl8CXJsUP4KnWzAc+CBRl
rooTfcfoM0lm/EeFe8SOd6tq0qFMhu4CJ/cnL9Ah/ro8Bu62c+aLFPTucKJVRw8L
0xulyiPO8U9oXfo35EoaNWslKVB8Z8w0/cbpEVhyc3mt/lrCZCxUwUA4F6g6u18B
FwoAx8XqMJjs4fIT3DBRdS6bawpXO/XpJCgFTEbbnPf0qV4x2c1fQkr19aGcpoiV
HxVMDeS24GOPN9U5oiyejUwWHvVvfw3imAhXkNKVBix7p3IH+9KosNem6CQG862r
QBMUTmHxV3PZX2n801EmyPbm3Kp+x+rE6IwRQcLOrZJrCvjesRUficX2LMXnWHDV
w8hflGxkPmjGUPS/PqpNpUITBdh+QC6ACclZn3orKQgW9ttCckRCmdV4lO7QkAGG
1j2qgSpGYmdNqVsfdYp7oCwms3djTHZY9wSOOzci8FG+qBwjDlNgZvBI2zIiM8OP
5LmS+xP9LoTtIAp7nWckYzTg5l+7kLUXQxpxLVtaxWWbzXcCrVx2AtlLYbSxYEwF
uAq2vmoRT2hGr+RX2fW/1WkhruAC7x9NeUv8jrZUM26RWxeBIvCwVGZ0GaV8X9OO
X0/sS2t7yijD7tBfhCSByk0rgdt26rWEXkAbmrafdEElkm8oxpCqltnlggBsxaCq
Upyzn8hs3DOjIPZ/onkTTViy+Q43+03sVr0oIpH/ZjqTBtXRttzw3W78sbmNJ2kp
NXRkIOQIv9dUSgWeHH25sAOyOoHHIlIbSl6fnm/IdeJq8NovrJVH4RKqqdPm5KJ7
baornD7PD3YIjShhB/NvYDA6NZvDaAAhWaeFQNCDCneZ734eQXdhLcEyJmHSsYQn
59reNgKi/05tAfNgrQFrmBQhVyfe3bT/tacbM99l50xsJWnuZUXB+o6e+TDXmbcM
TOQxsND7N4MdT4MWIKgf+gIDzD+JTNMUDvDwmWBZ+MgP9XNBreWgSBydKZe4Sk0y
PrWTlBHAfdfmzBZHCo4qX9FHupIqmpFToA2WxF4c1JgFAcDExTjDkaKgCbhMEC8Z
v/eveLqp6w4lhzgwD4N5LYxRTCth8KcrnHk6V5PKC/drpJkAuO3Fc3XuSxsn+V5U
66G9w0oW85FTAOn4BDg+vyYntkgJW8kA6O10fYAsp4JvgdH2zdipFd8RW3vxpEWC
njTAX7sAZwAd6i6ogd5mlWpYk0pEhKn/bYK/VOL6IrC4GBkPrtb9yyQFWwbAYwpl
BDS57lKNg0j7WjeGoXNhV7RIUFmtS9GAmCdqKP4IhEgQ1D5Sx6jfkOQoXJd1AcUg
FPb9xK7sFzEtUzEBT9LhyZwxZ+Mk9yGisa+ILyPrPqctxlkCt3lnmIxhHP4U9n16
XaKS8r7gTl1gdxFgysX9KxPqrCfNRiHxebiG5DSUH2iNH7Kic4nXQ7QWb4ukE87e
xXgDa9pHy0MP6f6ZKzFmazHNC07+3YlypVn+QPQmBQ2utbQK13Y9rewcMOyyyQXU
CXgPADycMQjB6XVHnN41RJ7utY/8sGvu+VUHvBoXz/JQeMPoyvpJO6lJ17+Zq3qn
8h0ZUJ33CYuBjEXQJIuo+Qs8ERfPbnmjLhOj8w5sHKOpL0jMQbHNdyIKehuabDTj
Z53P10o9QsqL4j6HzXp3b3cspOfVnTrDJqQDB2eO9i+2LzltyJyDvE1jQFoW1BKA
GnD6BoAZdLmYyDRKBkGLl4JZmven/4ts4jtbB/EmrCfclUIoCOq3mYvpsrpzNyHN
7VApdPrURtf+k4a8ijukyx+1zn/dpTqhO9aupVTBT3PrGWAGyIEask4PCO4UDVcq
UTSKyH6HTz3iAfKF/GIKQAe5ZXBq0ksvht4272Y462M+g/D+EhkL7lKYdKZzPbeU
TAPrcBE4D1j8qxp3KFpkBzjbc8f+pZXGcxFZwbf8CyfLPb3v5TyDibGNr5Vht1gJ
F1bdZ91gpw9BXq9SOwFRFDbRQG5HMLhED7LUt7vC5MV6471P+4Q1ietOaFWHlOTT
yK27GHhHIWyIm84DsAsA8fVgfgY0Ea1OQPje59HGHGZ/a+xhr0WkzymSID9jaDNF
HDRsRN9qzpdtMXLoUfFx0IgKWVzRx4E8l2JKYYMh6ri+kunsPKIdUrwJct7sHlUV
7wj5ddzFQHrnfWYqR73iFJvgXP0y1dFz5S7CmFpmtShUN8LiYrbgfk4YrCE7lhSE
tR/H+CymlyRMSvFJFrfEwQUWAHU5njucSW0Q2Q+h6ZYqztwMNaGtHrjICet5tiRA
cauw+nW7Lj4STGytMw1c0t9aUaNSu1JiX6xro5pvGAZvl2SiST8qyYPBBvbvrdy6
nATxXsAj7zrBOBn0HPGWEp6U/SIjLG4R5vFunAA3FXzzGI0Vxd7EBn4EN36colpJ
ApbapG1AQF2jvtQe2MjEDmhAuJ1jahzKi+7866JuPSwnln3I3bTOhp4CWKxqnkm5
C5M/HJckiKle1FBxuTCmtFSTitvu0Js2/+OCNaeYSJ96KTVvb0KWedgciQP2AMZC
9viVc/wBVJbqXlZgtGgeUyUl0i/r1uFANIWovF3l30rPQRiW4mRcpsQGxbd9SA2R
m/r55LlQoSLnG38YjeMh2nn6QOLF/+jmhpNx6hN0se8OTtEZ2UZbFGGBOhlf3h+s
OCVV5Jd2XObe0mD2MeKX1hcj+H/nlIwKNzroMK0y588Y/Op0TCwXu4dXUupvDYac
FqZbmzTQ2AQuvPfhN83bM+2Tk9GAKghvM3EfC0q7uzyrcPpsfRJZ5j+aTf6k3AjZ
RBbmmnPDcKu/Pq+k0G6JuUNFG6R2rmT/EX2y3kpciVaUqPewsYVXIW/nWnsuifRE
0LODGy0GY25hEMt64PCvPm5695asnW/s+p85S+xzn2wrqbhe92YsaUQmBzRXB/Z5
AgaIZUsWRTQW9WXYOlnwfJA4HftwBeXNZSnKDm+LI1V0cY2w4WTdR9/AMW25+FLN
6I0gTJhUEfpz9FId5sQmuADSTQPhru9tfxu1ifMdDUZF93PLamoO3kWoSHdTHuAU
QZiOxaMX4AbBsqG93s92hjQs3savT80LyrF2U6jdDCcLZIn5O38BORrqUlpjiTRh
wWdBJFaHqvQce84SSbwQFXo4MfIBKEwFAKOdfB1fNEaRdoKWlIZOTSZBcTRiilii
nHy2zwfzHe7mA/D5J+gbunuQuG2vcLJMQ+paY6r4XymEfdj5QHYavLJPR6tRm/6F
zA0jIaJBVDKamexGVydjsVpR1jirHyApC+Z2vHnFGTCy7V7GmYHALN/8f161leib
3+81FcspLu3XYL8eKoydSan6oit0RRjqwydm6bJIdP35zHZAyqcsefb6ZeG/wKNr
huzoCw8JdoygbbsyckRnxQ/d8xCpJpA70oeCwHvTPDHCRz+aZ4kQweGe1wkNggvI
VHNel7d9xIMGi1e/lx1IYtQbOQVOt7kUbrQLs0KZcvnvopJ1GjQ1fKQOlfCpCKW1
nbYBvyJSIJoVEFRM+y8UknR9ZQx36OB1FtKL8L0xT1MV2MRzWjiwcV9/feCi3039
wfuOZKYNu5e9wM7ohapglY3NuN7q/Izun/MbZJSqlA1ldkLw2sDghawoi5VO+Soe
c6G0YYxor/LWfIe+D9S4oF5ZO4x+0AOvWhaYvLIYTYRi71aI3iIZVzGTMwvlegOA
BG/678jqefSFwO7/oRbc2jeK4UTtO4AJELbtd2nNvDfL88n9LKcnOy176Wbg/G15
9LnP5OzFJTuqRL0m2IgkLauClRBEgcUh1tXqElMLBsUuKToP+FsoiwkufwwxmugJ
1mQqb/CemY2a4GWSWLMHh4T11+YfMjE23kof360x61xDBVxqUFlLW0K+AmCSdKV4
gTCX8DDIi+lFwbYHxfad/7Ac4ZNx9PiWwkCmRY7fssdVPiqt41ZVmF6Sc2+6wU02
kS6wWiIHKTKERiQPn3jEme2FH36Bcoxf8WfUpSk4pARKNOxL58KdXa/9gqrv554a
4I3VlTRja6BqXYdY7mwS7UgbchkFj8lBCjQP8QUEPDfVHZPSxGRaNdlnRdv+TnOy
1jeBlHwgwB4RzarhyseFXKafJbtaNJBe9YDYKv75I8/HhRfABYhjZ38LZGCeZM9s
ts9MMaUMy2RD0jrvLcbBNde89hdvSA23ErwAcosAYHFK4z3X9/+gd1O1KAO+k8Af
E9UyN7VmkjF+NaDnc1NoONUxLA23bcyCndjtGkTEw7GD0BLov0TWJgFgjrTnQ/Wp
w/ICWokx05C0BZYWo/FAjJf3bSRlA56T0nJq+28JcPw1xPWvXiMyvOTFO0zgVJq7
rYuihWUsrWintcMIon2y0RbBVmB38hpWn1fiFASeHaXfUdf3fY7Cjxc5XTAsMSvj
ERc7OZfcQOdHVwHynJbfGG6Nh6mRd+a0WvIlaGCDWqab+nBxknwYYHjNGGBOf8R1
ZZehvty5V3VvZbCCQvHydGhHHMEvl9zlGlgbPGvOS3wDiv1kN0hQvG7eJ78puzkv
7dvmRe9SRPE5ZfRqAC88bBWRpxKmKzxLJ/rc8hk0RqvI2P6Os/EBifOPGCO4QqFk
67Zlk8BxgDDhL41OuWrrpXBEKOtJ9vuryYKTs2l8IpgWB/LD0V2vpAXoA95LBTjm
A4riZDTgUej/roG6CJ46z5fCrPb/PdPa2EBPQZg9f1QVTYhsa3kimp3jRYlzEJxV
CltborhWnzq++UuksEq7Yml1Ksc6JNew32GryUaiUR7UKoItz6xxnd/0QC2r+mZr
OOesLddBpkgHFqYDNSOP5Y+bqwfjFUqVfiJMvZff54U76L0mmtYFURlUoHpLe+HR
fK06E6XHid0AR29Fl0HdM1akfSR3qCctjKXvJvB3s63JYV7LQD3p6YZCZXrsFWYZ
f0AanTjvJdLl0/OZn+MhFu5VMXcNr/drtQfE8OoRcs7+c5XLjFjfqRmoo5fDqxoR
xdyAnKU88GRbzODdZNg1nJA6ryVylFjQUsufcSWlpbfcppk0O/cQcYJsFqKVuBQ7
0lF1rUgwyQDfz3mrcC9J1OpBFpwiMJwt0SMw4GgsJwiliZOnFIBgOdcq8SJ/znkx
ua7vp5TFIuFDNC90XRISHPDnL9jc2N4WocVFVf7FiYCtAChbMXj8EjnARouHRnb3
G+j+bQDy+lVfN4tZl42SDFTEmRR/gPrgM3AlgyYPvYPcrMV/nb693F73mEDnygG5
zpQXAqWCmMLWGHV1jcn4aSC/b7jeAfGFAHgWPcIVVCjrihe2TR7KJ2jHymi11cC2
MrBJQuBe0R3DPOOuzK6gQPjmxdn18Y/zh+DdTiW5wNcYr1Ie8BoaggC8ibZ5a3H9
gua9WW3GQCeGzwBTFf4M1uiRwrawKJqSskzUtad3lyueTMODz3GpgpMPL67u+98z
TrXkdCoJh9XW8K/q4MFjRUt4QIn9U17/a1ynzFcKxvR8LbN8TZT3/HhIhiESlOAq
9KEf22bfR+zMyHhpcaXrssEBAcnxPPlx/obG9btE2rAQ/b/faB5/GVfDo2jZWuNu
uT32Ht2XXcVVqIudbOBR9vNRP417fJwJUWr/KSIAWuO3pfLc8osequMQUfBwV0gu
5J626oR4vrYF01789Q9V52sd/FLgaZMxRaXkJvYuGsOPSAoMXUwlfqYX1EVsgX7w
3YrktQU9S3QaszvXhiOjogftOa3mywNHWTGIjhXjaVzRbIrRLyQKoyKcxfatQN3P
BRF8w40AfKHpDtQR8WFmCaxszzk/v8D3aEvTHLqr2sevzuMxf5R9QtxMLss6Uubs
LsdCX+0vH++D/ZJcCGsJfKFAVmoNJ0VPieuhBgd5fxhXHk/28uBLNyOQLX7CrgIi
8YHLDyEG7WP+d9A5rIC0u+AyGMtp2cBtJVHLLZ71GGBn2JuC5ZPjZddLh3tCY4f7
+BiIklGWcbDvnRPQuh6ea1XXmEMyHI/9x1DsmzWXOM8AYhz4KP/A/1ssu27e643X
pJCgyH/PC5pVb0IgjB6vY7F/R3JB50n+HhneXJhhvNnBU+a1SBe0i6YQjUIQUYmB
PP3cCYtJaJph18CN9inD6KshlIVntvYyglRNt+c+LkjwG0z+y08LosEj9ER5knoB
TKSlFGtxdPfO5xr1DxRSc2CauKC7kfTnque4hq19QohpzbJ3PzoPpUB9S76r0l5M
Bc7AYnfxhtBF/UqK4/xqIgZyYRGFmsZxdAhF+fhnIXvyNqidLpvOFLof2qD+WTFG
UZIPQX0MJCQAXICRpVyabsL05s7D+3eHgIZNrcfaByNAru+ApWkIOW36onOAizpm
br9jLaGL2kNsXyOAaNYO7GvESuA2oagZuORvAhUlk1dMKRVWc0STjOFCTCQ8GtCR
5iufzghcww69y+gupzcH7/EdFGHFHU+SsDO/OxGLYnssw+1P1qUiPiWP4JJPYPhH
3IKNHmfxG8fNaKhBe4b1CD7br2+TlwopKdDfWfIuv0qrgXUNBF4dnsqWbUk+fh94
2vCfB++IhsYYNU0h6tb4r8do8M1COFs8bCqAzrm5WQLpwns7PKjj34qhDyZjyHcC
AcX3MBPZ8dopySWy6hMi176rutd4uhU533bYtm1e4Rit9PIJIEuUXevBMaiOSMyY
Gn64VxKznerzdWISI6dX6dMO6XPpyU+VrOPKWyxyUitkjMSn6gGJg3AG7jiKmd+m
XxWy9PERhrjwHTkftI5FYlarGvOuhD984bkqTfPnmpisP4xX8rryo4wf4HmLkH0R
kZmlCJ/oA3GASdBmR9wYP0wVQd1qpP+Xq/9JtuWI5gKj6GT5lPW0Hn247kQ5F3og
A01cCX4K6M96TDCv5B37+Dfd+h0XEFJIuQT/Zm0cUGv1Zvh1rq7VIgxH4CA7LdfU
Yg+9H03QbK4bMn6cUklcJRYw6vcJ0+VHWzwI5a13L+bxez7vthKQBWIFAXfmPxeJ
3eN2neOTf2KOnuWnBz5FyUAb3PuW+MMhPi3S0dDgGy/0S5rjqDhMMNRSXrDUC5W7
2ANRRfnkCRWzXkQT8FzkhXoChoLu02kDZAiN1mMbVwMY8TO72w4UFj0qTuDlHrwz
JgslN8cXWxerZczKY21OCFueNwSdcDOip94lZDOIsmo+g6ZEuYxho8eCTgOM5oyI
cuqewJBLWe5dkzh/6Zj62GA9kAw/qrE2B1jCRyTAKM/r/qe7aFPZ8NbYrk1qc432
K99oi9hJXLQj/WJMrhafSv5TQTICAJGcVt3T/ORWKg6p5JDTFXO1UMwEjaN/eOrP
cBdXwes5wtBPbeV0Ov0m4KjWEYcUFPjtkJoLUp2R3deQm3+j/nFjkZlqMnon1zC+
knQk+8Tp6LpS39Zjrd9z4qoc3zrtyLylhEsvuCTB44ZRRfyqFFbucwX2HaErbxjG
miEtf78gP24lA3hAJyljp/KOxIEKnY5LVQHDd9mI1pLvzhSMeG136IojF8O4vrws
HVpPVpkj1VXt2UqBePUb/wUX7+At5kmljm5wQNEr0CL6xTwR0LEUORLI6didIncY
4pr8P5ADeAXafzOZgew48iWCbc3FJj7TMEqarnu7/890oykHUwe2idyOXo9JOLsH
a2D0vvBIaTHFayoaWiSeYJRoohz5QVjnmq6uxlN15sAGg6cOoNAoCvz1tCi5luVY
fuKjrIEzU8+K5rEih5LqKVLSpAENcMh1BZz0hH884OhxbPv4JsNksymfLTW2dZ7e
J7sBbedDeSaPf9cHhUYcHMaTku6HDJFIjfuk00lViEWIuGN2pncRRd7VRaH38yKG
iacuCVF1sBnP1gvYAFMH5fHRonhtZM3C+nRABZcqITVf7g0YwKJZXfHUgEfqp6VI
8fhjIzX51Yrlltsb4k746RKbh2tB48fNoFV43orlcfRuhSd44Wed09MCtRKFJWTz
MyX6+s43Hgq0cHCxhJTr7j7wedumJReUhrXAyoDTdvc2iz03u389+bwoBpePH3Jp
BIw3pPQzxHElLk7JP9ODP73PtgtjQLF+tLxziNYaamg4wom7dWCM0DZq4snl7BWM
8KHg36HlxBY5pHcKNQHOjWxNdh4i2E8iCxRDjs6Z13tcsAiKGzqnhC8f7lpdD/qX
N4SahSZbBQo5jjmXMGzxbPiwJN1acEj0OULCgahyZsd3LpwGPcus61PpLmbuExAH
GQOpWTdQ06+4plG+QQh2r3HLwiYq6X3AdFnSK7LqegaEUWTxKGhMdJKLgs2nEtZs
9YEWICwTYgFr00PN6t2VhQ5fYKuXppmQVodeisdIFuEecY3QYMUgd9+oRz1OVRU+
fSivRz1dUuZ5Dwt8VHc38ZpUT2wvwbm5cCb/nECWLG+BjzJO81Pzjnc6yckmCCiJ
q46Re/aIEQ1KPv9YHdfBQ7LWqQ705H6LPHPl3CAa0VXXkEWNB+XyuVsugduv4kdT
8VPP/5ADgieuYEFH7YyXfieBso1mJ3quTQitpkor0m6/PmFjxCwX86M/LEUTlcR0
GN+LEG36NAvkkPeidV6273B3WLSDZP3svUf2JUmbN27GXLOnO645qSwWpMQEQUCs
whWcT6ImTHiqb9vz5y14mbw0e9q3Xw0z+r/xQvGJFiD9WxqXRmyejyWYRf+DMCZD
om0eszih0/S+A33H8Nobpl0tmTkN2pP2+FGj4FB8ESS5GnJ5kYj55VsH6u4My99b
c0yq2EqaCo/XSInw9gwP0zMv0jlXA2JgOoa1zwEwjEQESDvk973gO5xXretCiJAW
aBiOwZ+f/LTX2EQYOPtxb6geIaCS/Y/eEoC9/bx2whRaknKxjnz3kguyGZ610N6v
Yxo76Zp7HmkSADJPG+w0+6jqMkBovGWnAcjdcmN98mWoZRu8CTRhzVnVJos9/Mn6
nMf7CD2M1gwWAwlsPqepMINVVTiBCG7jguj7wcbhvAtHPofjLYtAcIkWM7rZZKI9
+rVeE/g7aj+Wbgqd/InH/fP9ZW3sY64Xb0uVqKAF+sCHclrHhxhUXJWDxYWZNB2x
Z+gNFGEczmLQwZKuL9hVxj+iWnkOgH++VjJ4/HapCgpIa3E+Zansnh8KfJGQ5bOh
AWi+qxtnM9dZUjGS/FgoTzmyxF01v7fdpBdebdURSq94pyXf1gRQpW1o4a2xDvpz
qTptpIZHRSOPOPv927NAVXyUN6L7+5dguew6TeePTOiCCFAcrYsFEIaKfMYnsUdZ
dFCPQqMZ3DeAYyzn21eyfRrs7sjt08cM0fWlLevw250eWTmE5LoJbyBIH+ALCDrP
jWVflorWwjsi9jvkZSuhLEUaZhwcL+NVjh731UDWkDN5d7wxtrsITlFjHpqHXtWg
4RkELw6UWo1cUKm285OL3k1ArWEKSXYkNCklSZs0GKN9glJBDXYUqtqMpA9Lc/10
t5zEMRB9EGYEqcnj5+hlLtHvrXar5B5CIYW9V5UWI/Lc4BNG275lKQF6WEoUsS0Z
TLZRIUvKBp4pcuDCBtzE4h9fZzoa/G9x4XoLUIJGKQrZI1t+qjXPJXI8z/lSQ54T
gvmxgDyHgDupma5TzZkhte7flLMpUImhKTSS/UqsfwfzrHyBcDzi8xTcKUytEzXT
AtZ632DTfmHJLrWWKsbmJfZvJ4dbK/N83/+RWXh6/gX0z5bLnV6JK/2sZg0FaoVu
NhTzoLB28tZw9PV2AhODGoXU32nbIjfK4rx/UGI666t4HyEBAE+j7OrAARDI7TNN
Qy5jFhp5Fp6cYz8SxI29V06moE3PME9RYlQOXfVUNpZrt498TqP5fmokru8U9URx
COQKu4o1QQIG3+jypvXRhNPbZRCvVaaeW4YJvhz4rSMNUeN84CBvRoQ8Qz68secy
s1+cqjQEV2WzoBtlraN23lL1PsIceyk6AI12l0kuZwwJcfuyEWqo54RGZh/0PIgO
rCTIzKdFsV9NHkVqxGp/JvBcN6ahgQbtDsT85Fs0Dt1XorNoZSao6PYMOJnazrqM
h+7LlQRfSzXkqllUQZTYy5krq5yWTROW9UxsUBP6dMR+xYYKSk5SsjOtSxpYQ5Gq
bU2OyNYxybCv4RRPzARsB1amHdyAYGBMNqwvQvgjWJXROqiVDrN0yEBrpucJV+3S
4mBhors6AKqoeBFTco+WYpPehkLWhtswKfqO1yoY2L5IGG8cT79jHAgAkibhX0IE
24rHQCe/8QbM5iJyvaltG37nKBCQejkB68c37dw2kAf7tj/61aoJUxDbxL8MPjNR
vWb+0y8vhjFUxfNmbQ2Dhn4LFS6MfdmS9BUIsKB+U2optgSU9F9K1dpeg0rvKxIx
ugUwWsYNddgFNbRn/hfEU4KHKltwt4P3KuupkIMweHBqWFYO6xZzTgiEYMQNrS/F
dC7yR5b6vI7vRRvubfBHCOaA5zDvaZPx+sMDiFcyTCG19c7QwqlKk03iMDKOxVg7
ES1VBeG1d4m2LXY1MicEO0eHdCVl2dHUGm5NnLWQYCzrM6gLHLVptI0BUMamEnkL
d/rJY5VZoiMrCR0po+eu8MYuLUuhnCIGegEJrsAW0+x9hip/LqrLFKva5GcdjC50
UaWJKxos4HjWGrceSa+pzPSMXG5IrFxRD5ojqxX5StcXp2Zvh+o7xrFGpKZ2u6In
x473NlERwU973GNVvR5p8eKQKD9XauBLLa6gocY0gTG4olu2lfF0b3QvcYCnK8KQ
37AAuRwQ+6uOUTfJnBgc7AAzJD/hkkvjuRPD/uW4dabz3/DM9NLtPEmy29vFl4dB
GhXwmBgM3k0PjfTeGIwSq7cNrlEYWIIgnga2bPeZtEDzFlmIQAGQ5ewpV8ee6r7D
T0e0o+fHrKt4NIhPH22IEpUjO4Fhhegmp50MYl4mMNGJAeyKFY0rHf+RfyqTJhTq
W7FfgVWzVyFB6ClEV2JJHWyXbI5Fx1xWCraKVQyvw65kPTFOEpwMfY7mNz3RRITC
JoPwtt+Nca6daQ77hrjjipTn+6z630w1EATSR7NI5I1/OStA9uVL5eRzRbu7BX6p
KYBKpOd6Kl18ovkhYQjcWEqyg3Ydk4GVxM5GChAeUKQwdcMhh6F9/pCp1sgMLIA+
m34B3gu2pr2S2xpDD6T3ZtvzVi049RbE+HnclrOG0W+eAFZm/VDjB7BMF6rm8z9p
bRkMzCcAxCGrQgUFnG5CLHwOsyTQ119NqxCpZdnRdg9fxiR9wjJd/kxWzCKm67Uq
BnU2kRCesAAmyeChlbFUcWZhNdiy54z/KNYZOwId7/vaLG3jg+q9UyEh8MGR13kR
1ZDFvXiq8aCrvObBcTkHVhLkwNfrys3IZ4C8jvTQBwvuMxZcIMPj4GmL5AGbKBcb
+RBqRTGbbuWwhGr54vM5PwCYnZubeFIDZpTFE/ppCYi0EaU+DZ/7anYjgwhkkCNq
VaIjHaP2mmOU6O+vT/lLBMvNIaFDvrEL5QNXoLAbRJpVscVk9KtBoM/z5SdmD5B8
FgcCVXRqyQ9QtnWgEviZinuUgeeOSX7cVwDF+Cf1159VMkw9HOUEN7ML87ODhQu4
TyPc3AaydYNj9gRc2DyI/j5F2rOlt/qYg1rDnbFjaUALaNZgv3i8XDvvDKRJV5xN
/ryL7DiYi70N0azJMkAiqPjsfAx8vPwhqCulxKBQpP5vn8J6rutgMlaKVtpAkAa5
iZg9oCnbbM+loRetT951LhWkgTUV0sFUjyDq1G3pJOFsf+I55qqs4x0rVhpHyzQ8
QhqC+e4BkRQAlkM/8sycGQk1aNHpV4bJA26WsD3FaDBCYuRvW7tIbGmsHUr1Z6tX
1UaeTEgzK9KigOV/4VItkyit5jvDfAOp34uIos+aMwKUsRFDhQjlY7adr+jWJmu2
aRmqBgfDdVypIKAuw+S4Uc2nWpIT5D9AHhY1ffSsQihp0Bwh3r9SNPxXxPevE9dd
+z6Kk7IQFGhbhx4HAGmINulia0e3/4ndKFVPOhAMMTBko1FUfFqyFWolSUqxgcya
CX41kzKJmP2nwm2TRCUUvmzJzLgNkkbiCggyt6vWpl0V2xAhpPHHc49uAtlntfJA
Sg5pG453P/wwwplLB6m2Pqs0NNw2wQaQezPwL3fzAq7gPKRF0hmm7srfBMVSBAR5
tMT+3iXWGmiHPOYLpnPLs//IgRrucpPIAAkAgG7fBg0CuHK7MWnb7ejrJCbAB8vi
aHY7YJnfw/v/vc7Ret88ZM4xRnhFc7DSp73iA4wSpcBCGMG2hfE00Yw+pdZieIVE
ICmuCyoZbvWjdVDtcE/cyQUpQts5YcqxM/OENwa9xqWvo+ez06ufLOVWplc5UiM4
/cYw2ZBK6tRe7j1b+SGTTBxx6Lu1n1A/qbMJgleJVZwO0zkE3kn9Kkq8U8dsWQ41
vDcSJC16/2MajeCe9IxYYh0ABS7yaJgABK885FfqSrQ26B7rx23uiGq8e6VRpqPR
+mvAl6mXLldWPQpZlnSxW86sTbyi/cazfKxfkgOKxWqWlBWpZN7M+qKgfl9004cu
ocqqMzjWG/x2uOfp2zoRDl78nmy2zFtakUTllsV3XR3sKMW0rterGaTb0xl75S4L
yC6fLv/tyf0AnqxfJ3do60agV9dlMnK1JmgSSBaIGGILfzHA5NF+3F9W7SZ2SKny
3eYLjlfuNFeU0L0SfzIGCFfvRJX/J+RgasY1KQ7thWm3+2IMbJ26QDy2eTCUMons
dK4D1HqBDZFjMb3uh2EDuBtHK7X2/v92PvP5r0Sg9QSvwkWS+PIk1bUpYz01UmVy
c0q3sGmqz5OUuwqGSnYUbkqyOxMISraKNpsED1LNI+I2kwcgvDHu9UV6l75mneHS
ZhDKEcgooYk6BeeKhw8nveUzlfoErXAI3MCn4fVoEVyinPnCyFV51satkIGb3T0W
+VLtAyJf9Cf7njvR/e1UJFDZQ0CkQq+WK/AHXNPaNPFF4lC3D+LMiewrp/okY427
AIZDWhnDHoGA1xfERpoMFYck76zGu2dhi9DAS8XIlJpKk/ssc1PzPtTO3ISKemOf
8rIf7FNQtzM6dOXs/nPIaCmq41b9YcY5DHq3b261IjyVPQA/E8YADERbnreNE+Oa
6EgkLRkgZ4F0pJlinq2vydQEftvpqLili91jkcJkaodOLdJD3Z8/u8E/L8EaA9ti
ynp5awgjkS0pv21FFlCAxndo+jKd6ljZnBv424ekbiMMkXacotdUhqwHWDR7iy23
4S440Ujb+hPAXWjr1fsnoz3FavT/JqCjaKcOlkxCJJTUUTAZZzCB39OTpu96LP4p
kG/t0u5ofzQdIFPrVl+NyYsx2vyfk0GLe++oTaCwpGQMU9vJ9XXun5bRGvbEwiq8
DbePGrumu5tBZ+qBp63mMI8CeaXoBzCZDi7hdWQmTR5tTqC6CjxmdZsf+Ke1zT6k
/NxRn9DvvulCmiqjfamrSPzbQH63T0LzxO+yDcQyZevaNx+iUMB8YEnL3TXk5Y4Y
j8teIMdMIc9l2d44vtewVoVTkdq9j+cV1TZC3iRH/8gzz+YigHDthgs9w3hDn/D8
74863WpoLvqGmUbF7qyAzvoWHdZB7nq7lvWc20b9+eGpxSfdtHSjfDxbhPCS40Fx
Q8CDWt/k2dOlJaGn+lBKInarnLX3BLWsshSFmHIIg3phxgETyEVx0SOM+MBLI0xZ
UJtwwzGF8guVNLJxuYurax4nhrEDOr3fAKjdEJOx14ShXAXlCHi7dGYW2jAVZHRq
JW7HQofcX1l3AxY1KzrBoFWV7qTWC6Ifo6lq09YmG6FYGv1X0qtvI+DE9SGxrTTi
5ZjOIBbTdRwikoqAw8LSOu95cpxB0N4JY5pUqt9xrK/hSADsgxyqTNgVBiDmFFVb
O6B0cL6hI5loZ6Fbp+1o/oIlI8yVJ83MCKQVH2N6qLM4zwrKZF3E+ahnVZ/7qFF2
AnunDye7QyZkx07X6YDFfoeG1kFo3yrLLoxvRz3xCn6QbHQ0ageDwy5dIZmJDd4T
PCh1WbvFEu9jYDR+v4uBQA99wMSMAZNs/PEmPTFN+kvVQIv/BjdBMlw8Q9ZjMqsf
1wtt+v+brPbFEI12dPI6LZIkzZ1OlcDHQqy029dqx8Wya6oBevlByRRH/V+LCpPc
o+7eIE4Uy3nJWbRibFKhSICb/Hd6z4KJi7MqsOLmR4an5jbQcXRQcJTZ2t9LR/jL
KngkXv2wy5JRmzlhZJS3IbtTgC0z3r0pgbY2PBOp/mn6TbUuRJdi9wr+TfsieRQo
yTkXwWCe+vuXEqOdRihf2BobuwsmarQMo0FSN5OOrCwJiam/k4Hm+I0we+lKwezS
kOuMeUW0nS/LbHas+u0+LEyA5zWXKEPKeEpEXk0zvTvVfgFSFHhxB6nIckh5Hl1a
R6rS0Doohl5+p/Z72frHVQ7Wgwv1LHaH4tcoesmksy/u87NLatRj0cYmVC68QVAW
prgRnLpLlNfiS0Cgi/iOtHZXgARAfcQgdDj3vr4+bbjR99KFkm/Ta0l7BT2XfV8E
+rYHTMuzeB2tIJze2+r5TR2lPOsajkOBPiPIwPFW+vBJtFt8w4fP68HBenm/reO5
ZfuRSRcMZoIW5F/tv1SOzCNorqr/FkJiUPebFwVy2fS9hE8yZTLsx1Yz+1LihhKe
nQYxSFGpGw4AM7Gcdkw7SEtoxe9fvT+4OdPT3d2Jf/SwtdHMtA/BKsyKgOU+OOgg
9Ha8NyR514ZrEs/47hFk/BvlxZJ7s8A7lUdia88Ghzjz2tzek3b7Izbp9wKALEIX
Mb9Xolstz/6f0jCQt1ZGTY4vpunx3nAu5MsSlmvIwvUturW/Z0LEqZQWVCN+WTlr
EPa8XvTIFe1v0xryUOAgYCsn7dumyeEbdgPCczUcdruZR0ZWDYWpI3t89OQLsXLv
VwCtBth9OGFpbZvVM+kT/Sze2gKJvmGNAs2mCoB9xRU/pBnGtZ8TFR1B4iR8nWAK
CsZ0ZPaIpawugECByh6jsf0PTbZRN4fzZxy9tCyOlybqEGvIkQbocOcMrSliFCof
5SJ0us03EXJYiQNvVLtQ32ilve5GBNaAY6YXi8PK9X9OTDo1UjDstkgNUUbppgfd
jCU2BPyU5+eo6bY6TIOOvo1WheN5rwx61bbueKSKXOp4PNxlvQfGAswd6oRRie+w
8fhZKMFMC+agGE1kbpnG9zpDp5LpxTPFAYWKfx+vYe9aKVTdZ8dO8sNB3nq6g/fH
oXsfu6G0hDwZtzGu2CVe7hxi1SgBNzlgG2GULfmsqrGBXJD3LAnbGIal2T7l0SGF
Xist5DiuB9gelpqv4NvR99L6ipLIIH/ODjfAHn9BYDz4DdF3vpjnWGjO8I3J6iWe
FhdmYGxGfIA6s+6Cw4AiXmrs7B1qGd7gctP91ysKv0d+dLgLlrkToCa90Xx9k1GA
3ijLos180UDLiLcjn9wcTObum6CQgv2DolJLBgi8x0gSDmQzymUpr6OHiit+Bop5
CENsHOnUcLbcXEHrtKJfsUHyfTo6DkpLuQpY38XlFaSZWB7nN82TkXNnn2E9N1ld
u/KDP23eZXIY3QqsToOrhkmFl8sGSZRnc6NYtm/ZxUBkp664944iMs5QnySnwu3g
6IncZPQ98XcYseTU5t0ySsTLA+w1F2REV6qtkPdD2xeSL/WpsGdMKHkpg8i6OFES
XiWxRZK4m8PEj/doOdPCkZtIjjjsKE5Lj75LfabgmSf+CdNANzM/lKfF2dIZK6cb
rWgWyJ19mOXqUgpcOvuXp/15dP9WkHYI1eeb4Sk33YN9YucMx67BFBON1696dZAW
X9xPakd6GU8cRszkK5lYBLNi9cK44Xz9QHwu/j4sybIEBcaNq/kQoEL7XKnqct+E
gC/wH1vPeLSvr0xrQ/a+1z5eDDybbotsrjSPRngF7TG1TMKOVHbL7B6nzXHw5T/0
fGcRxE/GIR2Q1GFnymbrvj/hQYS1FZjaQJktie/5OvkYKN21iPxcD6YM/QvwTe/a
6qYapabUyuZNdrqhYdzRrCqOtjfOK9zH47t1Ie3mpsHDlsBFJmSS+rDRXWGzF+F6
eSI8+3mz5eMKFLfP74c1PEosZ4D7atzFnavXj9f173u+3f4xlt1tLZh/WPwyd7xl
YWz8u8jKhd6hI0ph1OK94mOt5XVgEPeLCDPpDOqTm/4tGOwsyehYiOj+n2SqhVWi
7EogYfdOfDB9zzMwbu/NL4Hp1jvzaVJ6wV8ZribcBLf1P5aN2dQ0zJ7oZrnqKfr3
2dNxz4zumUlnJsr4e8LX/Hc6shZPXMolgb4+kEVgA1CmFBdcIBQ3anXcEEabvxQX
hiRt39XWr+uSUR7PGaAynWqj5aV2OjzY0exEdpDZxIZg868CbpLITeT3375Y6ey+
BT4jYZwYRBkz+6klu80qlzvwbZ1hsh3k9xKto71Sei+HWd/ahlE8vShz9SFTLlr+
+Wss4wyOmjaXXbx6UscNcMTLjHaTpM0cCNldIgSJ4WSkdFKSV31bBKF032ulcZYL
RMz7/+ZPuB7ztYBTF4o84/SAbpLM10FMnHp+vlflrBtaCX1O33kpifkk9JEXi263
ZNEbQy4PKhJ6XiiEjacYNKF9XDQJCZF+FM6vIa4Bdwx1vq5SJ9pLVxq+Ln0i8aCi
PGx9thkUPAOk78DrLNpA2JL5+S49BHEMsh3EJbG++GHRgUOX6M0Bpr15JYP1qLKM
bsWEySYDCqZ0/rCBTZhcQmsr4Xx7J6uRrl7DN6Sqo893GyiGy+tMAX6nmPFm+tvP
o7ZlVFLlTvgJUZtOMXDMmlq9XX9TnaQHp8qD+DnfA4ZNzzSgULL7zP8HGbD3FMCO
8hegY5oZ4wHKGnjbMxOigJxOGIXQnOgcs4SyzuyMxhedPY2x5EbXE787SkI2Fj5N
exw8WgC3dTjHEBOokkBwu2GlOHMwt6lIcdZoUks3wS20vWwf16lgac/C+BjQJVOB
FjoN4IYfxeo2GrTK3c7mxe6Enr5X28YJW6cLbdcfWuegDUnbzD6ryH3pCHXy6JuW
ShknJAett20l9EDd6KaR4QfWlIKmVJQhgIdRptES2LqArRmaBpxYwAR7WEA0We6Y
pCej8+kUugQdHIWooUwGdSkBXXJxCuqhYZEWgzJ00tJAshyyvJCIF6kDDkwOb8lq
+xuy8siSyTxettfSrd9twxaKoh4WVVp8UY1Svt2ztjCe7ujo4P/n/+5RR0zKShHp
Vs4g6oZFQBt2OKQEiKqCS+X50cJPvVfl/NWUVJt0kLdWxel3RFeXl3jeoAnmhqLR
mwjdX0Zxt4eTbtHTyBBXZ8DuB9tnTFFO/REtX/AL76Q93Mshxhbng6gxIJDKRopg
t7zep5p+ETeN2WbESzjj0WVC6QoX+AtGZQpHugvedF3WGa/lcansUItc0FDQOS9H
WEsDUTIUD35slbgjQzWLFhJA9bbwxIu2hX0NcTs4zPFTqfVorzPK0lJ/S2NNjgRS
mc5pp6r2jl1PoZFxhVXnWnaNjsofnLdO0F2fCcRA8mApUst0qbEc1TzP/DezUKrI
e3dzkVO4zPtMrgzQG/L0Gwn3xkoMAOMvJrMq3FTmRyUMvXiKDlqujHzET1vwIOC3
CKy18T8fcRzrZuG40Vcj9E5neV+5CeykZBcvMl9as0EI9OYNdAqkLbP4e1TklLks
M7zDRc2CX5da2qQv2LLW0t08c7XNap4T7nT+LtR1mWJ2mkQDEgyVUUwyxqUW4RLc
A7KTgC2blP/Qoko9hSE/y8asqXcZqIL+WMV9N5jVPXRpqwhQthKIJ+DqyWR0M7eJ
8xDjDXI4g5fzU8ufgGRgF5jDc1ixPV1EdJl6rVXDJMYtyTaTxQhzwKjBj7mFx12y
pc9w7Mc8dyBaNbrrVxLQZell1AGjPlA9r+PBbmS65w1xM+xY8Nwwge++y03shUAh
b0l+ll45AHFL0cp4EEmjaTNeFdt2lYcGJHyLtfMM19f9ChCnp8a+tHLxE/a6ysbE
ikZSZRYPfFH9FCgxua/X5x7JtsjbfkB9AO/XCcK9ZO4ytq+rGorraBUtaVmHPR9w
3QD1WzHS8ySHK/cZdzG/quu7fbWi9ULJwG64n9Bc74HyrERUe+3fiMO6YLYdUOCy
0sjNOqb2FH0hdnT7iQ2/NrRQJD8rYWRLaTdk7M1ipgjqEXNyoSNvqFGA5rz197DP
qUdA+Gpz+mtLWMGQhhGS7oZUcj9FD8ntzcB5Lxu7UtZk/sqC4H1FhD5/pTUGx8Al
UUQNz60PUm4NEqOBQrOmNw/eRypVc+5dxNiKRrnLywTCrhgYAFDdu2eKI0d1epgP
Q7jbO6PZR/qy2Wcw8xTTfAr/znWT47qgarLYYg7rrytwneublc8ZfvuMYa4cDslz
5v2+dFTD2M/u0B41ASw1jzuN50YIaSWv79Gz130MTSrWR0Nj1uTJjWRrRwM9Jtja
nFjJ1w1uSTzXoEKlXcx/y6jkWZ7vZwwWgMSo4Wy5Ic2ckhONzd8VM7k94uNrW4iA
wb4zfIycIClP4i6cM2XZdFIvExIu4OrcbyNkz0yPMmlw/XFMEawbMvZ/Qi39JqIN
cKCWPE+RTQgonR//vo8plas7VKPMJXINRuQUO+na2nnHggbyYFVtf/did9e7d7aK
og8HRfjU4hTFDb9R1bGvj+MUjWOksSdbxDQsWny8061E/7yfS4RSbaS66ya+5RMa
Ci5iM/HLqFaVTqxb/rcEBlxIAKDpgl2EHq0vjZeoLGkdDG6J/+5jUQdvSORhHwMJ
S264ikTLR3w0Pfc9aWeCgzqXhYetmvegkQPvhOlW88tXBE2clZCf/+qbM7QNRlrA
5ruFcBxiESIOi6/NsMpX76X0Mf7JONAWhkL8Sweq8wTUAM3are7XsBSj5Isa01ZP
p0jaWOUqCjcDO8R7lZtmeZKB+xNISqZapDMw4s7CdHSyTZgVAahtHQcgjnUIgqeE
hg+45HLyg3+PTdoyUwUnwMj/qhhV0+TSzEy5RT/oEKJ7HwvS2PYLWRoIgOAONwUB
h+SKSJLfCanXQ1kkq+ADtFO4T0pYlWwHt26ls3Cxfklk1gXetihMGcTroVOFpXBo
fEJOKnetYaioWNj+GQE+vsdkbXvHoCpV7aCbWlNrrGvOGhxtn3eKCa+S99a0VlNe
+ngHiq1KGPmaItrbt5438WQe3qR6YRyRD7xVHxtznnM/ncV59FsoxL4Zao4+Ossc
NBk9IeQ+3crdayISgGR5Qr2CGjyKaWaIaaJxypiq1qdT4oxjL3YkSrjWHNQI/rIA
zZmlhUYS4f1ug6Ebb1O+fEwh9gawxziFDb76Z8Uc+Mcy+tgBWRJ/FxHggEh5cbwL
ZKYcINi6Q9LFmQLkesu9oO9VuDsOPhkehOEYujfU+RdxSL2kYXNfH9qxOd0qZeSC
XktNl5FM3N2jO/VsoaXUG6srYz7f1XrC28Dh8zpAaye+Q/cHXnq3T6A58lw22Zag
oMMLS3wk2bl4n5GmpS5sRymW0YhSbeZry0TExPBe0fbRsATBWq79NkTZFBHywguA
gPtjDQnlJb4Y2Fcv5fDfCZ9X4+jc+wm2eNCdkZbkCMGGVzgJYXvO2NJdZY0B2ngb
31sCVu6QMjDQ6loUYLKN4R5TBQYhHPfaReR6BEENpcJuiq5VK/aoo2SbvMAZ6SgZ
UQUAv9G3apvuHkAUOUZgdXRZgNAmh3TLXWvEYWQF/k+JxA8yI3gszHn3sYtwAtzR
PjubuhqU12Y/ZTf0a3QkHakwTmXgBfBCWGO1BV1Dc7+U+g8OCMYoeo/jr6CkcIg/
S3pdJVsvwDnTQ9xKCUZZ0sdjbvDTzzNvhadny53fdeWgWS8pXcctm1zDJ4i6uVGS
axveGoSDggk1PduWsrZvzhZMjV43mGW1IsXwNqXcUAMr163uJ23nOp/tQlY9K39H
2VHtF5gDGifeVySf6f3bjK+Ln4wzZWoouLX3N9W70zvIh49SkAUb3ppb4RcH76fe
M7+6NssLomAqHXeZCfxd58IDt0iVTd7E+X4m1HAEGT/ErTYmdEyC7AvqdJS2AbAX
w1+MdJOugZ0OgM0NwK0+EX5BUP8K3nc9QM/D2ORe3ZZwZFifWCsit6qjiSA7wUGZ
7qvHL0kYbq1eDBFLv/lophae0iEwhBp5ZRTSMt/9q69rU4Va6qLaDSSdAW8MxNhA
SgNIaxiKnHeJkHAceOAja0ZeawmZ6HQIlaPijcWm7q8NIXXCCIpodYBITV8jmYF9
cRLEenSnCAeosBtaGxGGQV5yNs7QGiDsD26c7zNfL7d0HkMHIC+Sb1YI0tt+Dr3w
WgiZRlXG7/ZxassBZCFm088VyXoCB9g9zbMrG8KuIZ53NRyWVl1uX/KSCuNCp1Bo
WtufJDoOT22RgdLDBi3RoXFsY4vCcJpAzaYkCrwCrmoLv4Xt+ZByDqGDkMo28tNm
ftrN1c5xHOCl91aa7wiA2LGX/CGKyaxZ0TA2ppUHp4zuBNR26HxjsIod35/lnBqt
rGO8RGwfzJbdtHJ19ks/YYkqMKl3AWT+jrM9N0NmWBkK9tVFb9AZ+hKct+4ius+Q
fTANH4bKHuvs7Bgq/ykq3Q+FunC2EMB+l9WD2A1VOR61Q9dXzaqoWAkH6bVQEJ3/
3cMkRqM0pkrYtfVXNlfEhe6/yDqllNvqGTnGU3u+gwxLFBNeP61dmAPZu+O23+Ax
7AL+LQNrysxGABI6Hp1LJYHi4ZIc/t0ttaCpq7eapwjKdExTqT/w1s5cApjE1OWB
HK9unN8L+RolZRUFhp0Qbypidnq0/COi1DkX8JTVgdsR7Bs2tcTrVfkORbFA27sO
RpK998AHzNSRmvaiXHpe+xOgKbW+6jucs7Osx4shkb0nVu/zs5Tsvfge2yy4R0iD
rJh2KmBGIdBt8EtOQArYpcCvBFKDiNs5koRDs3o2DlvUiuvz0APHvX8pk16OJgkp
v2QdabwdaA0QdjznUA4lOlUz823cuFule+pD/2qhpX1I7n1np3faDC7VbbVxXr7c
fsn2f/Nmd83471ZRx1is+C4ZVdygCwsUE6d59e76FNDEdmLyu++1Cjx1ZxfwJNSz
vy0dSSrM7ESiPosjvDz8nOvsJmAxHUvNBqhYE52cix5I0LChoVmvRwpl3ZbS7gGF
phBJnSnC7lD2y2brtY7yj0P7xiYf7p+88L8qIID+zQdWMvSvGZao7nRJ7RLSov7e
peNG73idLPC3fbv1WMwWmTclIa8uMV4cIlxr4lCzY7fvMaEPeUHgWKhgkix8w1Z7
p8sM4HFaj+n7vQ9tkz7lFGP8YXQw6sHcXPatGskMysxmf0ys+C7dUVNcFLS5AKBx
3ff5/4Xc25FU38KeCQ9klLT7lXh+bIxqkOCVToLYKnmL50VUIKFnLzHHqbFi32Ls
MEh0hbGok0T7huB0WEsArWRRohJ7+XQXpfXllsoAVdtAtcNdb9ODohQxGmiMAtWh
wjLBO05CH0U9fSprL2nh3NlpOrIQZTLkwerLPiE+PZ0ze3Vit9kZmNYZPFP8QplY
uTSiTf2+VSGZiUBzwc77Coh+PBzXSc0AhAt9v4zHJMk6hvX/LSGZovmehBcLjqNC
J6x0FRH5PLkH7PO1AvWJaArqZmyKVunYuGYgh22QOjIYdT0YlMnJgvVRWpxqSRyr
d+V58FTGFMIJjCkVw0EYTlnDuSIE1e3vkinosmnu3S98zTWfi4DijGtIMzQkd59Q
921j8wGjORCztKcrh7x8eCkzFvAbk4uSQ+a2nQfVjVodMsOSnAdoB7mf4n9t7P70
lVJbEKdVyT18RJDTm86wKmKDIml2BoOhOthd5N8mgwz7IgQ65eU+6WRWlLMSv5L/
HDmnznjpc9bQZtHbPyseEikQiZ/pf8hwciKMTW8SkSdUIykD29apALajYo5ZXhbc
KK59wBOu2rhVtviyovVMYMghfLe7OldSFKBKz8kCGBnSgQy6wsOrkDPSd/dharg6
hVtD50AbKNmUpz0QC8VPwC2dYBS1mwfjmpQ/Vq1cUW+h4YcO2VHSdOXTOjAReTh3
tRSpGCRy2PblLeEk3ARCDSeeM3PZw4B8RCsV4kPUnla00SsLiV7og7POJa/RSglL
SclwVZmZWGSY/UXJ7TgKxgBVk/NCnd9ObJwvAcpswjsnx0zYokrUbMhDkzjnbruD
RoTq4MgfI/3OC/0ftT7/YrzZCepXmZQ0BzbEF7XZa5A7Fed3APUjhKdnXM/f4lOv
VxS0284sbWw9T/3KgNMKj98F28aNLoVP2NgGzS+YGCTyBaOSJemzrQC5A98xb/Ui
q0nUBabqLy5bD0dukbmiqtZMToornE0OHKpdfyQGSVFlmscREantm5I1NxIXY2DH
aY44gwk+BDP9F2vsrs4lbwc90nfW6SMgQhLhYk+qrtOSQfaAF1pQwkJ/f0P84gXD
TO5PMcaU8aZ7822q83g2FXHGzC430v3KSHgLw7CBetzP8cDSfYpwosDrmaJithCX
Y9y/Lq0OyDA0YaZ7r4/axYdER/ATtfd4pJMgEXFoIFz6pLglIywXUDhOAPQ0pEDS
Y226n06Qibf42Iz1aztxSjxOv4skyU9QROQIp8E7w65EBdaqJ1VPRol6TocX4slF
Yt5iE9VTvGr3VeyCTYK43he51Vju/F5x9eEAunL9HKTksfJeJD/97D7NXhXart7p
bO5x3J5yUgFyyFD1ejvGrhh9qCwH/sUbZoppa8sBUFuvbj5gGVNVYyiN80hSEvH9
y21fwmZ1+gPNgpvoxg8DG7nethPoWkEiLp0PNTncnVDrjuKT/70ErHMKXV2MLKrg
zSaGyOC36OqCuzTS4N0mlzEVXJxR6EsktrC4wBcYhfWRiYZNjJROtLgn++PXooSa
jl+V4pflMyhuqNWEj2sJw6BOyvd2um10Wc0MTT+YR2RDpQCpgbpi46VnStegYBrA
MXn1+eOP4ZcFZdH0TnPz8zH9OsjRvZgu9nYXzaCPU5s4ee0HGFGgFrz/n8qgqiWn
X/gFHz3ZLS/YbY82mNyuCEXr0Aj6IGgp6r9dqAgyf4bfV9ejPpdgNomcqcROgAMv
APqEf7uVyHgwsnQv45p+GYB8LbREiQDjP10T1h4stk5yvdyIBCMyZ9bAD5ZXc2kB
JmslH3KqzrqHc0F4RBBw309+I7KhyoUO8qymzMP/zLrcJ4OcGtzMPghkO9ZQ00wH
YAlm0ESxJRJuIbmFK9HLTLYwXKlT3xwmM50fte/ybeXQxA+QoFzHngY/jpKlVMXp
lDAPxToUiV00DxMRKysGCDCLL3kAMBZYW1xCYeM0L4Dqnt1aW2mALbom3tJkjJQm
0QNYArAJCScIrHeyesn625t8L1mX9+2RB7VptdpR3wlxe0aFKOKPR5jkDlWdBq69
Q+eRZeBzxzvphzRB452iSG0mgR9InNh3m73f9VGBiUt6ha0L7og2a+z3LR3FLJ4k
YEtDpNDGL5cagTurPdGFAS4oMTEkhhQ8NMkP+ejnDGkEyF1zLgtSJjo2BEhNk+f9
aYMwr2lGkor2NWty2Zv9Sul8v7jOKf3r+dFIq5AGswQ/aWcglSf5fSmPGGK0cgOr
oDuFchBaFVMErmppQDNrPeOG4sjRkV5dfcArquD9Ich3VK4OdCPSbTyivDtx9Qp6
9ojMUjjsxjGI9K8DpEt0HSFerVsR1m9yd5h6WgD90/+qJX8cm0OQ2RWjJxwwIDfm
FhYqUiJ/ITVu6YLiZZa1A0Lsvh1EXdOVq3/xbLcg+jz+ZqBz0XuDRqPF3OSV3TL5
XxWqvqpAjjf7IvkOI16swTYjn1HHZzZTKLAtmJGQN6+YspPhViTxmi3bumLvwVbq
Zb1mm3AjdmBcRE7ZuWzCixTgZAHqik4EumY3/hufW2pikap2ToajlfU6g0Qw1Os0
PN5h4xSLsu0qSHcoClHp/dw2eaukLYujrVhExAT/ZL5SCgVy86x/dg6dXn7N13gS
P5DUn0pfvq4s8I6k3Ndh+QA86s+TpE5nzAiAxLCyeK8At2p2brvsEQC6idbFozdp
I4Vx9usbL/R3LWBVWTl70TC+dyo6GOLlXTulxgTWcFxYbB4orPsEVgnu8Krp3jP+
LKmLtkFhssUcUkmHsftoxRk216BR4LvpzfBQX+P87oM70oSfZuxq5iZa2bVCp0FS
D7aT2D+YD/VN500nLMelfcvlY6rzP+2Y/PAUXP96bp/uLJxosCqOvHCX872bR9dY
qRhT4z+ahrv+vU70cicKgnr4xugWSe9l3O73mE9jBgPXYy/Xx4HuLUf85F6tOmAZ
CCtp3+qx7sDP4lrTFTXXPibMYpLvzBBU0C7fc60lzbk1uAEgf0cDFwp7QQGZnpsd
LLgFCTzsjhAL1fzA3fMQr/76myA6dvP+6kMtpS8r3CYzojvEzix1Ep5ggOae3Ige
YML2tl9IQi4LaDZchPW/esc2WyCOlCtDHNEJpkBHjUYxwfDhxnq5R1zsewyZYQWI
1qPXLjMOnLYxQSE4BPcHluQO2yy7INR5lKipu0ElU2+XkKzwvxptw3joRODOltk6
tOnBdChR/c3RFY4aFHojUAiz24tljWL1N0B9vBZJp88unUj+UmNdE2T7lEyug1z9
BhnMGgZRZvQkzT2LpL7xPIhAbVNWhpR8valypw0xjYq66LQxYUgPUpZhiHk5fLIG
VlS8u9omiHmk8VftQ02OeiXJzk3of2blKHQ57O2ippSU1Dn5PeMMS2JopN1Vo87o
Su9a+3//m0ienEI7VG5X/bPOcXuf9OPGnij17qAiS2WtJ2YLs/n5XdnrvqfcvOSn
B9ipLZPHnD2ohaNeGE93suc3qxz1UYO7I+WeoIierGNEMhp57ODQ6u629hWYIYWd
mu2o6IxyAI3VxDVQDxsDld5SASgxlH4FjqIDWyjEyEvsVDwqvI6ud4oyy6hSvlAz
KC25h0pRF55dTTw9RTBG2MUn1GUJ+6dHHkiIqJvwO24qBuef8jDymHlQXbkYwRoi
qylBowNQNbjFF1MLfURjpvBOpb4I8BJ0ZGSj/raVcRj6+nSPgf4380nw5qBphCcl
P7NGz+lnbiHW1PspvMaKFhGji4Cysf0vhSWKCqHvYQsFF1IpI78Za2Gxh8yg43Ep
rW0cD7yutZXtTnfwnE5d8EbNVkOLj2So76tkCGyMv+g+Abc/W2qWOaHgUkQKeuE4
C3Lwk9n7R99hSLgmnt4N9prOzFr9A9VxhiHS/ZhxUjXigo+xkJQ+m2lkljw4qt5o
pBMAF5VDe2kVZ9b8D+7Hmkm2cxET2Rzw71zoDqAelHwKoVA5bXIQ9FMb503ZUbpO
lENN1cwBYbb+6vFekdK7b28tDvbj8gaCfKECeWvmXi0YsOvLKj+lSe9M6dDUasEq
c6RK6leBelpm7uD9+0S4XGQ9hAgMgOtwSKFVLmup6w5+OgTX7NMHCGohUL8fT/SI
UFiqiX5/NyIuRpzfAIGsKefNT75U/jwgtzH/1bAzlQMK/Dn9vzNEP67I5CqU73x4
W0NH5IyDqkFvjWPcQXRNi038jt+0Gx1WWKiouD9gKsKyHGVBIDayEutrfUiUh+7j
s1lbU/m1O93YRwnFd1HAEUAvf90oSCIxLOS0NGDJKDzx8DIqoGDdGKKW1Fgm2xW6
EIF2S26Zv3vcxp0OIDRnglOdJNAODR4IGO1TVeAHZDznFUBjjuefEkoQD17dDlYs
eRbkFI0wuMHRWZ0gvfK3YsK4nv5ElRkaugDlmgTyxPN77iYHyl+lsNcpIUYQ1f35
TKaMS2QQ4xl2T83qEewbSB+tIC6BRMOCvDqXlqjw/BnpE+3wREe/CXGBNZC5VgUc
q/J/NbOzDHhDnH7Ry9Sfg1f8EfN9YN36UmWHwZ2Eeav2g0NV/eaMgnf6EGyEU58O
147jx3cCO9nxNCUkhvCVJsUnVJpK93kI1GM2OXvxmN58cz1Ih5o+Qg4ejX1zctcb
YdqidKfEyBc9u6OKF9X/mJxB5HyuTkqN7OXqMwcVcdRq+dgNnXF6suCckXY03Mgx
9H452v4WEd9GvXH09NqKxR6XsJJn4+i8avuzvxaLXBJn6TrsU5KjSV4+Nn7Czn97
N7PZOKA7DAwNl9E5zk54MJrFIb4TSBJpVUUtoBBIFcMIEt/XRqzMcxVlOH27BzuO
ZtGJUqqLW7kyY5wnYLJ1R/PRgixPuqkgBcdRR0kacKRcA3YtlTPlcJAIEr8C7r8a
pw3ukpFHwL673A8GDT4cq8BP3E+ztiniHWJbp5XbWJp16JrlYGbGn+TM0OpCmsnR
YKIF93qbwb/he6fURbG5KX8/x6NTRvzaXSlDtvEGuGebtytpGIL4yvXY5BL/nknD
fggAwwfzimoW0ReSpQnkwQqHVzhKKmMR/80Y+qjZZ19nkpnIsP9b6a6iQE8msTx3
3omUc4yh0fptten7kteFaqqELOwQDX2tLhGHvUHmdRdLb4tkDFL0xl86prgrQVwB
cSNp4Qc5DixICwHQoH0Qp1Th89THpmKU+sxR7+06UxRbwTWoJi8NuffetHccKWzw
94sWpP14NGuWvwYT3qRymcLRnsIVHwhnj9OcyIFVywAzWXiQUYqgFmjFGzO4QjCm
o9SLJydiEyD0siFv7kMff5ehKZV5Qzm1ZB8nDT7CDwFXyNmReqY7Bj0r+mlkh+kA
Tx/hCS35n6iWPov6mtjGetH2//jrX0HrxrAfkWKynV5PgIgUlZNfPe25PVecJ0Lr
gZP0/y33mZ1TurxOaIVW2QaQUHR6nV4/z/n2XTtT9bjvy5qa4jgjtUBwflUdzIYb
b4OASd4p2e05loI7iJ5jAOKWkQX6MNukdCQ9yzdC2VsV84G0tdpBMgCvJpT/WdVF
21IzvWk7jTcrmIpqETuQN5A6PPjCTxcJCCxmFqovC2aP14ZLMO7OP5BS0xexgHZ+
I8l6YVYGWwtgVYfKxLR/HDtEpw2oJRaHg5/bbo3aYdgaKvbLZerRdJXe4O5ChcrE
N3qbA+56IBpyr4GDmGeSLli6eULKb2W88ISgOwJORmLHqHMvvM+CVNiiB7PPZ78a
KmR616B84jBbddyRyUIO1kusoR3GJuVt+GOdljaBaitxkuwplaOTY92b9XRW1NRl
QAJ/o3PhxfGc4eC2Q3u2aSJGTpUf2nN5e6zvhJWJBWvGD1PmLGk37blQ3omm98Cw
2dnMiyF8oU5vL8rCyfP4sVXpIo3vcETxTlzR5jl2usfrT11DUWCatc4bi0tCmWtD
sz0ZNn4WPuj7SL/0toQbblSTkVgJdS2rDsT7NkGqYh/IOTJl8fvsBgPDZcowwHHN
TZmk6ENI46ie6KLjROJD32Osonhe/Rlr2t+y8ivUAiEIjh+oYueuuaU0zlChvR7g
Hude28IrfU+IShw4xaRUyseU7kUPZYXV2RNsbmxHKIQU9Iq5B5rT4TRX3dFEknjg
57zjkEw+S57OEWSWXDbuqGwQS8TQ+yYsBs4AhdYlq6J6esw1jOutkU0OdcC9PQv4
wE4C7MA9NAkqWycRLEHbAZ3aCVz7ySG27joR7AYca30+9ogmz7AASrx00/e6qLyF
ZMcpmHK9luDu6u0ieEDxKID0GXY5kCTOte8ue5UEok97mCLPsIwdA7L47eVWhOpK
PGaXgoXrWI26tKd5IdA1GxVxd+QFVzWh9/RT75KIuhU9iXa+lkxNN6jXkuaWXN5z
XhBsFEMamrpniNkhVHDAJCL25GdPT2fifcl0up6VKyYgm9HfFpdBIhSc0NXtscVa
NZqlre/d8YwHB8tBAOWrFexVKziQQWtPitBheJevGhs7t/fLwGa32NeJmEUWv0QD
0YKFJ6twX4+tYYLejBDobARiuHMeF3w6U9w32VgkKIEc/eKgUV/ZNDj19WyYMrSR
iL3zpcnriLUB2xyY17dJYFSs5ZGywOGmCjgnJbNvWaBpWTpxcAZPbpisTK1GkelN
fkzd+N5p2XZ0BQmfFfS9r9gJEQB3Xh8LbYI4yTJ+b6zueorzCTYHmlsjEoE6UfNl
597nHUtctVk4sriv/olFNN7JS0HDtqK2wEV8l35YEReFGTCmOh0gedZUtdQsKlbf
ascbBX1vp9i9Gz+94CBi6XPptJVK0HuIXziV0X4PzfpP1cuok4ygH7BC5X9f5eEx
YjFQSzA4hIgk4P8pojq/40eVE11GfiUQRkfqvF1A7Fq+CapvD0fY55tBQWb4usUU
lpZsZK+Xyd2OMPFEuk31raNFwzy3lkk8e0cR+3va5y40yI4+Sw5z1sqvEnsJ0JSy
hBQqNbd7POoLAy1Z0d5TElmU/OhFCUTlPQN1tNvnDPAvI+xgKprw2MA8KnI22R14
wcODUbycCDWqLFRWE8JEMH9Z6N/DQFnPoIC9lAcgctqDNPQ9NSAhjGaZDqL+NWSI
seG9fv6vTg0V5vsu6+FeEe4rs9BXTFKmoiPOKi3Gf6pi3vxENUk61VTl7MNyrUD3
jHjQeDPvmROX8kVKKCGg8wDCeSD1ty2XFaZhNTma129bK9EvEyC6GSvQrZ6OJ8QS
Id1+TqZMFDklRLHjApq2R30pcB5z6RQ33k92FNrNXFxbT67IW/90yHNQjDCB3fxC
KS3Bwl17H+KbZJ8TBxgs1LM5AXo3lxlFPVOoV2CBg7PM3oJCqZXBdSlIBKjDj6S9
o0dx5Re6Z0OURNe9af837z3cgBJU3UpyhK6Ko/XPLrcC6TnsxpNPqk4ijCHACbK4
0Mdj3ncEmQi6opaBZIIgG9fgJBNwJrDfq+n1PyGHOpeQrIzwN49+AhNeO3bFlFdr
koFvGXnMA00JxLSDwIBxmHeHrGkXQaIKAUjfCKvsqD0UQ1Vdifj5AjpS3AL4U2JT
RPjYTzh97sY5iuxrI2u3KmlBVFRzDkRqV/duRLsjXYJ4mzKxWLGRla3NtNrjsHr9
Y+N+I1q/3KCK49AWaR31haC2ydHnzvzIrIeAaxTvX6rqfTKzJfd2/YUgHf4wS2uD
nOPGulVM9H4fNFSQCAPaejSKuoCgKfYVQKf0E0X3Q6Qcr2TbSXPEAVrjnxL7QvR+
HAeINkcEI83VE9bDLEu9KF9inNcbfDVfJ7zZwtDWsI34JtO6sQABU9Vt9cbX2qAZ
G9Qqo6pxwPLqSvO/MLuIRG/17hoICoHPCKBtPk+wKqoG6npwVb6D84uXbkLXZ7wl
zeY2scsS8NWwKlD7olLiHpvPIRgCbbbvn5gajymFGcc+mrBlIEP9HtnJ7+Z/9lkr
gGrxK72yak9ilHsNyhSDbCSJsBnuiJHJvf6LiMyql3trTX+C9tzl7XXBwc07csI1
uJ0+ZCuG5ztr9Sd8Gn67dghLXuruvuENHfJf9yJc9WUeZ+1GK1bM+D6OnbkIhtmV
bs1emUkNXH7HodYZjl/gSDJhENFEDvaF/Qx+YvvQMX1RN7jnVY/BbuWjtNfiMQcA
kjJTz+y/6oEBSRTyUU8oX8l9Ahk/Rjv+odAXvrAtszwDwk/AH9mqKb66klObaCGc
A/JWifa56L9z++9+WwaON5EzALSfEzhhk1noe7VGGTJ5lAz8K4ML1fgv9IxpPL36
85CFLWAhfvKobWL2THnZ7kAAeUZrlWLP9ejy7zHzNR2MD+2wF/PCDuj2VO1XKFjr
4NPrwd4Wdl5Y2qG9f3fiQvQvIh3s3N9oqBbUw3XrPeDb6dJszUlMSpyLtHFOdenc
HIrjXraPcBLtbENrPuB32uyRhyaf5KUh8Fh+MM3wTj9dH09EsOcs2hzJMKu88rVW
aLfmgOx8jZB1YGSRLkC5n9C1UfjvmkllZOVYk8c5YK+lWER4nnqDXQyrCCrU5R9N
AjLGbNpQnVJ3KZ/l1S7cZ2Ttx/9xq8vQ8cxIBvCB4yLi7+qvuhiHjfi2DzfA+sNN
pi+mOz+dRYGPfCvOmRaJM7MDO/gCGpx1JQDjSsRPZ1oA9v1HSyA5lRY7Fl6QMOjZ
VJRzRpBB0WD9pWzH5hA+97tsv2LJOqJnTu4ucd+BiGP6L8PMdi05pIugf8ab3JgW
pb+ih3rnJXGLOC7WQmjMO7HeUzvGyphjueH2vgN1Ef+A+1QbYd8ldIdCRxp7GcIZ
mM08MmbtKw61izoihO0IECxUkNnzSEQq1AvRJmJ0xdcO657gKTUp+zhPnRNEitR5
CyrokDnVlnibO6er46NoEvM7mVN2yfBTHefF508fDR3nH0KixuwdwH0iLsVl/7wc
qPBKiq6d9cjCGEvVpU+AX5t6Ph69f99q97ZFXOCKWwvtapKm+cOSVJhknJMNaoUb
0uZSBAZWMXKW6JoYrRnMf25BSmy3Z/2Zv9UPyO/msi9zoGGgKcvElUO4Ylw9lhMl
ce+O/Hj8nIY7hFunx1mV7eE9Rgm2Vh9XZXhsw+ZyOkiXTE5a8oLTwuYPo1L30uOP
tonXGAI5/KHIpxiSwD/iQORRIL5XGIsut/hjmymF0ifC13pFDiaIaHt/T9vRFNxY
4uM08SXnrkc9RzXAoI+26nQm7j8bTa2KGLRM4OQt3x/g04+zDHbmmycbZ2XDgJfO
PeMSwqJuCxMwbiLJfVx3AmDf6enSY4ubghSrUS8LgKsBELlAXzjEt5w9bBfSSQpl
xXLwlLU2KHFXQFtx40yNznmgDyL5DQuxoqZ78Ha8UmcA1Se/fgExp7FrxHUPPB5i
miOCZDWEJMzGSTqhkLoMiXtFMO/b4uplyJ0XEhPkfhhpwYlT9XIHmTvr0T0Ll+sa
jpuV9M4vzEy2YizABdQkgx9WInB3T+0hygqff355Vjl/nM9x+Y7MsB7/1YPGyqlP
0Ex+vrZceA/LhMpUlBjlDqbmQyAeU5Qc/ZT+xf8fEM9mb9eTtbPNhYLwuZYOvowP
c4nwkEJXJ1qcWfyShm8W3L51kriuvPrPcQUjgmmx7c3T99vlm0VF+w5ZJQS8lPPp
OlsP790lXdzjZKOaWNkT8WIsFNgIYU5D9W6ZVAz5+5+tGBVOSQMwlWGKUbqBeXMd
s0J531Ee2Gjf+mYC61YmoP6iQK1KAYOjuJFTE62qc6DZy2CmG1vaAJkriTp0mXk/
VuYkBObcKjJEsCmuMYkv6hX/vn2cVyAtLgZ++GLAXvzuZZoH15cR4oPAU3vv8uF+
XYIPa8VSEeNRm7DEBLfIzuLYD7gh5qE8ZT5Q9mnB8yij91Nf9y+lfWhZyqDsXRq5
BsHE07kXFao1Yva/LTpaUM+T2NnbCnvl/ViBJaZlCsL8hyTo+XPulmaLMnfZCBNX
OtfsOJLg3lTzxtwMoLiddyeklGt9Twfq0flLhrwPn2jMSjCCjezfF1ltsmS12JaT
rbXT1fr6nSN7OdQGT2lmD2o5fmFI4pwLMC54sVnVI6+T9by4zwNCeeob+JofQoag
8IBePB1LajFJGP8zCfsRV3h9wgrMyiZ7gsI8uYOnICCLM5NuXdhHymzd+jWFOoX2
dd+a2EY3s4ZhdRsvqaJlxaeqMS6aRfCXn82aj90cRnOtdrIOl1g848hAlB6Ue18S
AbUx+JbEOVxzeFJs970OZ2kpxPQMGbbxjzAqhgtkVvKgcU3wOJgYX/tLpmjVkpJ4
HWquVVS002TE9xwNt0aRZPzTXipqhu/WQCyUor2YntClIySu2hTdcdINjOiYuKOb
VhB/DvW1Gnk2YeBhktX1ZDSgbh1LJo3PgOh1EC9MOz6uMOw3vXwawxmeKj5k3vya
PloPmXcOH6R3Q+JwHE6sN8a7ryDggkcEwUwiEU315RFi8X6CuXROZv0A1mBZaDaR
ggvH2yikbNOwYK5qbcElN/1xpcwkV7R6QMSx4EfBW/28oMckK1Fp5e2ejInL5lsz
8V3o9iAnZ+bKeabQmBqNJWAc3AQn0oh9ddS76pq7EN9h2QKxl2oAIjkzGx0x0PcD
eqZTigJEbvgtKY5GvAX0dXT+Eejt2UYH1ZG9Ja7VSHDdV+n5ovG6gMgV7oGV7w8O
JFcieVcwnMNaMdf9BLj7nxjbmpEiZNfWkS8Owc+FNKl31776id6n60MPA2i40J99
6+b1r0HqHd6rFlOkXFCigB5nOW8AO0OnN3E43JpFm0k3l/nVpf+WfT/KsFhKKcem
5qDKIRfJz+cainK0ECau8I2abAZnM3it5dYNungCzi0+9VLf/n+wVR1mbF/6IAhf
MEqkJuSPhWee0OliUdS7spzSzjmcv9cO+NQG1nLTV+ot0McIqI5oMca/yYFNth1Z
bjEsgcrYPqPB/9dxIJaAn1xTSolcvjxUzTBf2g3V829GumFCXWUe2TDBZscmhPzG
ZsOvFpqOovvJXfBNAgLTVOcda88ai6UIrEal+oBoqosjxZRLyJ6jN2vlvQ/VyuIj
qdAlvD9GIQ3YKCtkgZZfXCGUuWbDgeSf24Hq1qGat6FADCQbFQ6WhA4Q5CVWZsA5
ESEyQE4oCCrx6giu7wwum+5sJlWIn0nZJIFQglotYqVbqwyJQpUSxW0/NhFtlcvj
fiMznm6nTCm4Z8qOZ69av6oOpBgMKYML4SYzM00/71GSVeL4fjvdGIBtCvkFMqee
x5lcV42f0HhnAMHQN32kJb1tEtSTPMZgY1At2GCKlUD6Wii55tieCnKzhP34u9dB
O8eveTQEfJDDp140KEZ5PsNd2jQXYuV2aagx+JvZ7a+ZK235PwE9RF4Cmgs7mn9r
RkL1sBVEzZ5kJ7YIdjx5G8nkI5XDZY22glzMYtFQs8zXK0MnHoNgfAZi9P8gJNhw
qjSm9mrRQNh0vp2HqsseF2bI37uPhRIeLg7DPjK60KflIxf/xn6VyjQDnPh0EIs6
+nJh5sV7vezLKiGsjEIuFjErL56NMlvouknwLtxSfYkwuVRG0964yWw/Yc1JsV+3
5muEwqzw1HFLPzIAxg6YLwKhD5+M08N6uvcibrj6IxCMByVNeEfNGY5RhzEB4vBp
kIzg1TsBHPNWNOer+4gpO1au1EZtSf5HEOtpg8Uc7DG5K9EHvqqHV7rqg8yaiaQt
C10iCH099JKYrr0lNcgj1hbtQRf7pqhMMEcg+IAz2qagSkkEacKWwKwAO0aG6RoK
ogEs1JvNrAzavmUtXEbZ2RbCU8Q/71DDIZgAXQelkN3SImmLHL88VCXqXJYOeb0X
DqfSll0mAZo1ZnlZ09d0S14Zu/7OF7ShI/b+7GWlL2AqAPd/fGfhq/dOIW6gyLuA
geOA86TzDF2e9GM1WyksrqzTR9wgwhE3rdGKrsUULw1G8GMzwGPFUVNP0IK5ItIx
JlO7vH4BgUnzwHICui3vZCI0Qi8sszeqErUDh2nmbPT8YcsWuIKhx3qnJpeTjiGX
PMQdyxddvWC2InSkhmIylQ4WFer3iwF8okhCF9PYShGCNs6qvXxJa4gJMTpaMssh
3/oGC8L36H4MzzO2B0qvwm7vKc2lMUcHBfa0thknn0UXaqRqiageYNggKeM+4N2p
JOIYQLev/BEYA3r3QzBMlwle+Z7WHSX6nHuzCZwwVjoKYi2z8HydgaFz+M1Qezwo
qpiTG8Q4g3hdTY0GkmOLmF6/0DI2H88FNwSl9221w2M7w60aKDsU6a2c+JCFRilE
pIFD3V0nScVMKx9RGb1A3xzm9Pf/t1mYSPArfrsmE0sW0NHEOEXFFYKjRTNRtNTx
7JOOld3yIeZuXNQ79rQwv7mOb2lSsXcwFW6H80ZTEqxIPRsKAENrm+DRhayBZ5rv
si/aQOsKEUKhH2JF9KZ7WMNyCxGxHfYfvAJWEmGHqMlUCsKSUg5VVNAoq93M4R5j
IAEXbgdL84zhsv2xTopCIh+D468uL7SqjpnGIXb7WsPwpjiQ0jD6ft+XVKH9+lQZ
kHFmjb1M8jqwzAlDBHCVIxVSudXJ98oSAOah3Iv94Ix1jJ8CSkzz/0QQ0hpC2Chy
v/IAFBqITvi+p3jNGG3jrxEE6Hs+njBB9TL7lxQO6zlDcKN2Gj+yRQsbLAlqbMYn
k2xQROSDK2yWqigbd5MeqYtLQPCnAlLDGOvFZxhoFfX+vjXZcVu65X5Z0aVi5p41
C4tzBKHCJwKv9tEGzeYsiKmNDlzGRvNgtvcL/NF2Ml/0gWzo6mDEx8vkQWDMWJ/J
z0LgpcTMZWCDZcESOEifwwcT+JKExldHBnsxqbQGGOCJWbC+D+DvJ7TnYKoDsgoY
lu176czUzE8KwDBW+Eoy1142EoydoNhScYJATXf/MYbg792xriGuxOdd7p9iGSpV
IpXufB3p6lHXi44d34fo2IGBSiOx+/rt17itt8o/lmSJWr1mIp1DQNoiYMkb4eCv
Lwsaz2JIupXyLq5UYA+4lilRck7JtZpKpb1seOLoQ1QB+LQqn/PWgJ2qfrOXebHB
DgBZQViGHNbD1sogSZGFRZzk3jbk+Rd7+W6DZp9HEr8C/jciMCEVvy7dZpDUO1EM
mSCZA80ucHwblzCDeFEnZ7c3a2fVxU3OARWWNxBvozoD2KmYlzuUqaHqb3QbASy+
tNpD/3ZmKoEY2Vh8VifZzaaD3UuFwOfpVt682z/okxRohC2ro07kChZqkNkPepOV
EnvPMjgBRcLcVQTZEJGkviptnusjQtDXX2SYk5GrXqzq3HrOsi6AKSX1EZfB8nC5
9yi2sUPFqiueq7Q1V9VBKFbcMOvJM9JvM6EzVQYUxteEXYs0AhAwXdrQcmkUCJhq
idqVv4ToXsoPIs1wcZZezXH+Wt6IMJaZj7PN2uQZ16lcOM05iThEneen8XHerrKE
WBYhzxQt1LhoR2qCRdxJW6d3yDla6bDap5s1/NQQgPJZmrrUaj5Y+JJ3PYJjxeFB
cnJcKaBBMJk+ifowSWdHgpbNQipLFhNeHy7b6QOz9sf2TyNHrcobQWFI+kwmzpJk
JcdlGByLMNMIYAEcpl8aWwnYupw1YcjJQ6LQlQb+cjqgVSk+Rj3VBDoOfm2wg+15
xo4GgzWBprhlbRQInoHTIqKlHZzQnREGH1pCLa5xYbJanFuaVqd1dc6+R5c+dw4Y
3CWxl6dm9ItiNMcCuzW6mowIc/c8FrGwLNiHst1RxBc7zb5TDfOaLysfZVePOB/t
vCHpLPVV+Pu381h86ov5r2+kX2vmrLjd1HW6def3Pwjp38p29Lx1R+CjWCKJEkrJ
MBChWhjrjfdiOA3w0Erjpzu4DF0JwegTniIv1wAzUIcRMaBsIk+qfDZ9RyutjHdn
mGQimdJc7gFe+jXehqYwnJs4YdR+SoRhzOWUkxCPTPOjs0GyKyWB6mfnDTFbSUXr
xDEBfK18q9ItPlx2TC5s84iuxt1gbJZ80sT9fHkOQGwwyb4pEzyedYP36ew7jhMA
U6cxOjueIq89R1/3Z1gauiSoceid1EFi5lP7P16gP0XEzGwXjpJjZSIAyTVu8K7+
pIa0PEvVgvS8Hcm5qXf2Dz7xTfKetcLVk+HHcI5GdeFLXyXQAAP11BQ9Gaqze6FM
HAVlahZ81SA8a9TESmrI4kZBL8EA9V+EBr9UCiiV56EyJYZ+G1IxnOhniigIG9OK
2GbI5Ph9OcHHInaxdSFV/y8qt0CzQEbAOfNhJ8pf3RG3lDRO0MgO0RZ4L5BMfNkB
2efexQhUJ+gsT/KCi0UViZ/i2ujB4GiHzFtpI1H/tp9t5ztdQRFtdzGQ+4QEjIeS
Zp2ePICAn95HMIv60BXYVVKAEcSEdGSNB5OTKIvXW6tisxxI5QKztMTwCgFI+Smd
ChAsZdS5di79kd46Yclwq8RZczEPs+KSpsqvCZR5vdRCqc9lcgxQbKWn9KWLva4K
cl6uOT02UcaeZugfm+NQD4sX19wmR0G99iMhUN/wf7NniIw5DIQzwZoZNkRktwNB
xpBKbc5DYubeeF9Hkcks+QWnQtPEVgGVDA8uPSFPomg0sCKcOUXqpjV23vWwtB9J
TcAEQXwsfw4PBDCOu4qJ7jr10PsFGFnNa1AsSfn7nFylhGhbx+t2UfVADnG1a8Tk
PMRN+n9ilsgWWGZKQwvY6vrNTsUQkJSnTsnziIhTjIE1Ne7kz6Wjb9csxL/i/NXJ
hY/8OKY1KGKASDt0AtGgLBFSo+b0LQ/JI6kCMNFH7TfamlrhLAepkHSEk4hMlYKw
7P6bxAW8+eW19bOmGbtct5meZqwrNsIlcRE9zmfVpUKmxzEP0D4qxOL2PeJILXUk
3QOwCMe+hAiaKfyqIigiKV6cj4rtRJD3Q5Q1ZSfETp7vrcVe6JEeBvCO3icMYNY5
+pdeIA3cK0+kxbKSwBrrqNI3URFWkuqTHuz6oxBIrM45YwGPanSu9nthMpatIEgI
8NMmY5QvHnrDf0pIUwReb/esQOpg2uZTvZH6Zq8FJoFCqWoJ1TtT7kOK9+IBka5n
5w7Wke8wnXy1D42NvRTB85oLajaZEeu/ZzIc/LjhI6kPFTa5jL/W3ewkTp5+gi0z
QQbSAEXK3WjWOCTL2S1LRXCfNu5kXJBdxZiROPa+X8Y00v5R9q5ysmKwvu3SUgBF
MsS6G2cfTDzafhQrQbNQSw6nCHntnzrpN/9NsunC2+Vgpx7X8mdz0QvEskQmekPG
fxUcs5YRhW8O+nFHipMjFBIkWR8aCoYoLbdq9FGodQfazWl69jctVwNPZAhC484g
fAfqjsszsWwKzpfwWWyfhWT2inbfrT1ke+Q5oVfF+ojib9TL8MP5xT+Lairmgouj
h+OjOxEAjUxCfZO64WCFr6030KDSa9RFMNQv0eVXxweW7aUYwU9tjtLpsIIv0cq2
FfkCkwAL4Pz/Rd8ZIkK1dKOYU+5RtcJElInR9XYkxRY121WQB0iPGQD/zydtbwfD
rU12dTk20ZygXc4MoLIVNHefcj/5AMkk4ykNyXxCylkVKXZRS5JHZW9uTJnlD8uh
2GUlDBf+gLXcp1R96jNB96TKjwZkWyGVefSaPs1U34WcatqNvh1n9ndwaF9yTBp2
XJ/pk0ycyevROhkDRizf3xjVUJfkxOrja6lOkFW02J/1MXMIQFay12JuQpamUJca
bqXt+IE8lF1W5jKo8g1UnjSK9iSWsanqrX6PBJyZMd7XY5QoAYOXwVYucVmngBh3
+0/Uu5M7KfE1WnnYs2BPyjCekPjI5YRyC3+msYSecI5RlSAjJTOsbijfGEiZRFSZ
9ILj9QndZIe76n1Q/pz9d9Ue/jQ8niwIZMoHbpSJU0OX6nfIbPMDfH9tBEv3pVHv
kVKgowuSqC1+XigSX/lEsgw4+t+iCRgXApNCcmJCmmOGAMqf18hbmvv4JD9RnQMA
iFITITSJV0qaXPdgoMaIrKkG8jvxTlwb11RoFFP6cizX+ikJyRrQyXkXhvz3DJr+
EbmehzrQkbYgZ5BKw0RnYr2zir3mr3lSi8rH4pZWs2yaymfogcvO+F9J9UFtifvz
cY9DbWlNsqTs2IuC8EATKvwZJX1WLBbcau+Hcdxw/6mxBLTVDQkbVbymHNeb4BHF
gH6Vbb8+2wcaklTYmYdwIp/5rPGgGPtk8bT1fLXG3cygf3E3PIIR+IMmlhSCmaBG
msVpHPycImNOP0/eTiP08cgMaUoKTUGfE990WtVjUvRssKj/MsUWV8pyPASlX/Zx
C4C7h0kzRcvETyEyXkWPSBFogTaG71IrWvomcsznt0UQvFpy8/B2S7pz/ml3KPId
ZMJIazCo94j6C2VHVvkdlyLnr1l8YVdFyUlIHgUkFbw0u5hGKscmzq6MDSXnUsUh
pysRRXbSWcGRRg9z476S553d/FHhGcAPkGD19fIgQcnO7Whk+ez5dIsOaDg6VcGr
cGJqjUIS1eNxNw9PmrmKTHc83iS0KQfuoxLGAhmgaoFKFN72zo9MxUUYSaBCOz0/
Lq3OXx/D6lDk/3ZQPF2YzZ2RsO9xK5+r94KbMAW9zqsjRagsp24+Kg0XxKWLUtqB
bNyMIb+5UsdCfmY+RHBj97qV2rjO2Duy5Vv9ilB99gPTiY9yWGHAGpU+C13Musxr
MoMqz5JSCJwSmnes4wQiJV2PIqE2PHWhFH2croDZ9rOYtKTI9dDEqhSYM6EERVpr
yXbgj4QSJfeYEqBD1gs3TXm4QyOrTSvs39rZlZJt+JZ7EvdHGROuOfMZ7N+7c0ep
9/h/A86R1gQVDZRGWFxif0fuXMn+Aj8LRemvSfv/5s5c2uUEW5rfNZjtFLFj5PX2
kmFYoKQD6p5qekEoWf98YGi6crvJuqKInDqw2j6Jn+AOUm4rsnjNN9CeZhpNZ+xl
zAf4es9ottyZw8qgMq/0U/sYZ9mDeOf4uZlVv2o4OvAkVIiTkp6yRHDNrUC9WKp8
w6eYx7P/UNCZj2wsideSImLLv+5BtTpzB5YW23PVDkJ5etAg/Y5qee0S364xjqMn
EmSoBeB2zNoq68sajBjWysOAjwnY+7UT7k3mzQP/QsNNiZPxL+yLu7tp5DW3BAMM
seUEbI5384imTS7M21NcDpyEy94zcIg/MXLmLqzfWAxr71URMBXm/a0p1op1zwTb
9TxNCbqiY0AcHzpcasFus06zGtKBzgGUCxQv+h7ENtcoaTBhbx65ueZLLJO0lMIW
JHeE4xub9DP+d4pPAaB1UhGpsX2aW8UytslTxbvtCYhIOtn9Z2fb7GUoBWvTI5j8
yO/4eKFE7uuQ78KCwp4BmH3mvBqbImOmTVAdblrPuS6f5Chqv9pjU6Spj3mFYow1
zHrjdaZnfahElGl9VEIiktzdUAsJVieS5/rP2kOFo7c5mxs9pwIn3vsI0WDu48P7
HtyML80iYo+kfaPFja/9/4tAEVyjQV+B2idwsLN9pHKlKbjRBePnFuQE/V4I/kqj
+8Gp812bqTtr5E6t++yZGtjgf3djFNgGq6Mh5K4lP5qoNposqkRj55LYrvZQz6as
S8FNQe+5KnbHiaxae7Sk4PiqsfhU/MxO/B/crtfryajFRgiWPjowiXPY6M6668dp
fNpUWeWhG/5hI8NEcIwfZAficRGAyggc7AWjLY/DOJgg//JP9DkDEoryZzMIrEkz
oRacktb0iL2LSXNVDUDgxi4gWEPJ8Jdg74AdtR3zsOsOBXRJGmWutDqpvq4h9v03
Bz9s9IwANarjUFuNg+yCG8xDYLK6RGSLlNuDhCoh16jT7wuGDTkZHg2oIKlMjeoI
AxNoL9THGE58qI+2oZM+Fm44BQoMJwv/kk1dg1FNApvwkHI3iecRKcjbDHvsBLrT
TC1Vyz4vuJ1vimwsyubmhQtQLP2PqbFup4qdcSJCFfimIHlvQyOusTKC/2Z/I2Xi
GnGL6eV/+oTR8XkUg6ZmdFgRRYoPPrSEUkoM/Whji+72Pje6ET1s2C9loJpp1WAb
6D6nyFoSmTYYWKWlBPHJv41wfdjih1l/S4uxugC4ew6BGOsDvNx40ymz3I0xN1K/
ck/aClrKjcMhjmaKZCI8NwdDPHq3gTZqatjIIeWgvYE3MgHtk3LBhiCR00GXV63T
bJRCb2OVyv/elordoGMh5QJ210x1b/wYlXeW99jB+q/5z4sbaaNJ5LSl/1YSTwOv
1xvgGxUDqFUUlaUjCzr86VE9u6rnuaTQG0vIJ4utJT9oBoaax8PI/cyoOUtCBsLW
aIj5Pw1jmtEWHFEV8dfCg6nbpnXKZmrXTvFzGV132RXnpDAHpFCO9sw8WFkC25va
8grHOOYC1GDihaaj4hM/iHgC88XA/N1KVjP8JTlb2AcxZGsm+O7x6dHXu7vlZZdm
OC9WPVof7092GezScP2yrVtTfmY7ZQrusdNdmGmhe6Z+JYCL0BQQUNAUfwmQ1R/i
6pxPLubNynY4+Mv+lOkoJpDmEMt5Ps+Nr8ngO0z1UHdbzJGmB7yvhmPBqEsc53Zs
qp2ozemfaPm2UfbyyzSVEU1N3hgPzAKdpQn5NG1wftmVIJkzzQGMzrZVZUa6xYcx
GsjK8I74+XODSzpBSdJPpdKXCi5yDD7d+Yt94CeH/V3kaW9p0BHff/5IHF3WFfnS
41lD7nFxUarFCNzVP+bJJmlpUhO58gbVF+YAnsDoRCa5QCyTRTldktjtRfuUH8zQ
7pt8Uow68abIteL88Ya/2oG9ALunTI3ZJqngKBWJMvbgCVRBoORwGVcz9Uy7EMtU
UUvsGkwGDTHA5X70BCz2wB8b7L8QEUONBitsBMRENsSYALmG5yhP7CHH6RB/pceo
M8tfM8klhVvrX0pQ1vtwe11sHFS9vb6aW+ETW1aMVf/zRDKUa6SMCaFCK0XN+DYU
dGrFv6IyH2rZOY/Tr4gON9rgLnd/5DcdAa+G2GxyZ7VdOw92fSFtav+GnTQyC3z5
ul+6EIDspYIbG7S9o5K47aCq6puM+1sf0CW1C6/mi8383SZ05sIZWrjdtbHWcAKJ
zVEgT+4YnG4dlXjedOvZTi8WDa3j1GeLizBWX4pwNtCmsFxp6+TKkwLDHmjX6l2r
xZoTsFyqcn/CGRuFHaH90oOQkNhqBdrBATK92uFTrm45UThZ+L+l2Ea8OxjO5/9w
qljjTMASeiRcC5rVOWqUGCUTPFuAMYC7DGdKb/gSqkUMtlVrjvAzDzQ5V1YTN0QK
M58HY5yo/4pbzCFROlwwb0U5rIbeJF1lxQgTujUV18MbXh5Yz2ER0vc4DooMY9NT
MkZRmBwzUl0cnpdjmBTopkpvLfjK/DWMAwiBP4/NW++wmF4eexiTDH/9SxM0Urxw
zWTPwjqU3Xx69ccKRyneY6sO3oNtH1U7HjYDlEeh8InyrFOZhGeMFJ5sIdhI9ivT
TnVoA80CFnQQ89LMRlaYXcLbRo1tdQUcY6dI85EHTYFUKBD6Rc4w4LYemd4MRCq4
SdXjxksDcLYD9vLHMB2l9TrEQ/AfhQhVGsP1iMcP1hjgwdCUskOmRPb5LdERtuw+
ffrxLbl8T1OKC1w4DdMroJP1SQRd8vDgcjlMWpztsIZQaQEuKT9PkBUyBzxjU0xX
1N5c8LHb86hrp2QLiADxDL3QGOLg0oLmXnpZZmU+xEOHS/6uHeCDqPdHvsB87bEl
zBl6YhmOvQKaO0PkDY41w+g3PosBjGkToEqvO8Wgw+vKSudUaIKZHzUyyCc/wybY
d/Id59hIoK4vgFLJXJO99xI+PgzbfTkRd8g24UOdI1YBJtkUyD27FRnyTY81SynB
yjUlWUOBbc8w6C+Id4ViTIIocfXoVXM4tFEDoses4y8QLsNlKTuw7teypZ52M+dT
QEZ9WlvpJm1zAyXDlZCixzYhNLDMC7wq0gh0p88gadkyC7+552XQdmGp3FNQZB7e
yn6caR1T7ym7GxD/jyOccEJBPt/A4FoasI7Q8MBuNLBkImo1SU0Gm45Q9SBy+ckK
6LGK5gpJkC5S1p/POrDy/Ongur7Z9FrCSfq3g6rFY6hrunzBi1KdMSKlAsqnN7l4
mzXGr9FWAtesG68sN13aYiVK8qgfJgrJ6Cr5NfLigCcxiWySNUud5Ljms6Z4zIiB
DT4QPret3dajAiyzaHQGj6RQ9XIuaKw1w8X8oNDGc7Es1xzR9hqxUhGx0apQsy4x
9xCva8I9jxLOArP1gQkEKdGN1cHInGUcPKL7xZD3PXQ88KOSFWGYtkD7ZFWbOD55
aC2eE9VozcYdqt69/JRREfBNHs42hkoQxwb4WBqLrq8qRjxILTtT9J6LlkMaaOA3
myXMl+lt2zhCM34yXxynlYhySl2s/WOj69TOQ5hqflghOK/g2boG1gdXoFy4XQJt
qrlk8J36NEgkMHjiPOyiEdTvIEwI2brbP6A68OeRFlvOX4diQ4WAr3BkAeLyJBlt
hOUBDgrV1EMFAkenz3+n4S3gkj5RZkT798di8e1nW2OEOM/9zR8mW6Amqbw0+2/p
6OcMTIRidVMLF6ZxNvU2wsfSuVSgbrCADviivIsuiZJy7KWwugKK0YrgnX40OBzN
+LhTGaHM6jmRp2CGghH894BZHP5+K52ClvYsU3EqQFWl8k64S84oX4vG7JD1l/fc
cxuAOseDeGXh4ASoCcdJnidBFmLV7j2P07Y1498PpJbG5gcX9Az5z19WbE8Ikyk3
Fz7umwpb2AL2aYuq5ANWBzyKt4Ob0JX2pwDuZe9bDNGi78e5V25D1K4PaN8DfD02
Y83X1oXyy5ho+DFduY+XAoPmqQW9aozHdNSliIcYA1+JoEYW56ZWCf33UlX6jfsE
69c7V7EMWATG8qnzdc4/WdYcfykDwgpuJSLfw4QxSQufWfKtDUTaUVIHiXRM6m6v
hRhdx+1C1LXMTZB9MMbjRjSicgdJvbfuZUwb7y76sbzgZltLInntf206Ja/a2OYa
QDo3J9UHwRIBp3TRP9jKxY9x2OaMRUeyn5B47s9RTNXdSii4YZHQRs2Aoq9leOtM
10dxeMvP4esjKSDSoXlHJ3FdchtKoM7o5YZYr7zw9pEtLJVlv7muzXsAfzlXWLjR
3RfDYHS0hac/pFzowMcX5/MUlQH4akFyfIlxJz1tkLB677xIIS4o2JixJQ68Gbdr
NclkLCYwzvz6RVlD7uQNIiKhm0oHvoHL1d9VL/eM55hJ7mNyPm5AnhU6ep66RmYS
OtiCKwz4aWWaUiet0yF6txmXYT/Aq0rGXfZ/xG6wGGc0jOv84JVnZqW69rMWSQVM
+ayzcGomBrPiLC+9TO/h5Mv+YdRdxjQ1jjGZozmDDcEXGEQ0twag7ajwkJKdorkT
AawTyeap2C7o4PWqSZpV4BW5W/jZ3wFsu/HdPvcJkeZkUbTbFFdtBVWGdCDm3wLu
E5mu3fFiE8IW799htTAIY/yezHdtrm/U9ofn/zmzQm0c1Jp0RnWGTEaSuOHtlrjI
AiJa3qd2WRTH2kvlbd+MUBwA+Q1GR+xbCDis9QkhVNFaVH2hxfXKWyHBp4IrWloX
LfcbLmacu+tpYq4avPeanvhwWBqUW5CADP1/hfyF82sl/EWUA/WMnlYmGArQxEj3
N+hfKb24GEbVJAF0HNhfeDnbAUWvRjZqe3/pMPXpVB3I+G5ib8wiRAr96ty5fZSM
IgxAqaBXmIqJDPj6iH8kJkI4ETTxRtlZkbESdjzEUAGPQFhVC/0+6qODnr5iPnYX
PgtmOc4Lt2Z5z+Ala3/6UMjJkRATevZSlmDCy1qA8zQCTUSYzq+cuoahkYgDAZbz
/3CflZBqdBfLBvuPQpkw3x0sXomkpdeLBwhjs7jY8WQ0J3la9T2Fm5aGMT+foU2s
gWYXaHo7AWIyWPoNK79RgGMJ30nh800ZqdDoP18t2ThF/LMRm6v3vTaMKkB4hhT2
nd1Cd6n1f4vBQij51CJ9GQ04LY2AUrVJmgW3O/Lrdekdc0lnLRNfAUm3deM1xC15
cmMP1LkMq/dfm1+DuGNdCWh7xfpPOyTzNB/K7XxTExirdfoIW7aKjMV6zsPcxVeK
S6z5zhWbtya0/yr58yIAkczeS5/rK91JIZYBfpI7yPeKZbj8kaD3TwBUI4Tvfg38
2It9kvc+VuAu4q3rf5rneNyjeoxx6mvZlIln3AGX9dPQHA+k0arBmFLzg/veRlv6
m8VHsTqzKI+uVInmti7AaR2HJNBBo1M2ylZJxfWnDycKrTLfIzDJDmyTmfHmsSoa
MzAI27U2hp9SoyuW79CkO7UGPjyzEv4gI6nCr+mhyJs0owzUAQeloDqu0YkFfrLp
4Dz85g1uPqvTEjL55pxWFzphkB7wwKnFPwuS24MzyGkzfGzrdkCL8k/rXrq64hQv
OxFhlBL+357xUkUbtZmfyjoPmoQt9CqSKYTClISEUMyft9WCSo0ewSvRqqU/puA2
Jr/TsIlaSxrbS0v9nyEmuyTFd4tAg7ttCMsuP+U8gLtMhzlkSm+LgBYzvJ9om4ym
z0bGQQctNuZ838TIMFQDw/9Q8s88KVFncMwxqqTcgXXraWdOyhLbKcn+ckoH6Zm/
SBfxTie727lLBNxazeGwZKerICJdOSY0EmtfQeNz113VT3Cqmkt/VjthWU+/S+HW
OJ+56SDZQ9vL6d1saXuRjoh7KPqp50bU5FV7LBVKQK7R962mlfk3ypyx+XRkbRxH
uifTGJd1kO3q3NgOI8FDEd8XRB8H3RE4g778TmlkHelQCVF+tSfuEFuVYhzMK45A
jOsrggJC7aIEevat6wLepsBomVWuosaxJHa1QjDu2kQDV6KMyCaono/pfJqPdggR
YMOTf3n5n7lhd6iycVMjlwS1i0cKOuETDLvub1VL8jKKSDhfuitx4QYRFOMhXmJR
Xk6ewgYGDbpke7gNOLVlRZnUzQzWmO5qiYDranvogMeJyfRMOXeJE1oSLq11Gkc9
A27wk3XnKzdGHpBuU54jPq9HRNO5qb9mUV3CYRH1xS3tJJxOJQn9f/dDEQz6czJt
qo9cuExbFYhVLisRfHcp9QTkB2GV1c70+F1jRWN9/bgh4OtX8TQINpvZ9finJR/v
e5FbEtq7sH6sQ4y8oAQyiPT+92j64U4bMFVfq8DseaZq8/0Lu7AfohGF8da91iSi
bVyd263CQVY+irtTmZwq1gnMuoo8wOPRfSI5g74nfR9JnJYx1nEXaTF2nSJlU/wT
/nwfjU3I5iq3jvfm/sSV3oPkNMO3Z3EoKPZ3wqttqhgro/U7DLh9L9scULy0u+OV
ptmPz9sXGx9pr0MAx/QCTEX3nEID/4Fzl9cxk6zW9nzH+rhjMdtBhAypx30nbtUh
dS7EuXFS3s8ooOmWW2gY6jvWDQDnAVlbvnrC2uPVAWVUojWg3PsJT5UKpHDRQOZh
2aw+cXxOiN/wbGEPqu7T5WzpPbcvCYuzH3g9hD2PjAHIrELSFBU71SEtmhq1h13I
JnYorg6yAwg/UymJsu35LfeWlbgdzwieV+ohJJ3DmQTh4p2JU1kWxzUeYAtHWdAV
xz3Ez6k4rVOwoqoOWC1fuvM/x2YzWSLtbSWSjo9LVkVhlNDvIHQpnxbLUb7dunNi
5+mGk9tW6UnIHZZMydtsw6FSAXB0WqKJve7NKh3k2Hnc3SWthTvQ9CuYgiYp1Bu+
TzibDEa3CUsyOUIq6/yIBOLWYdYhuLQgDRAB7kBdX0ev5ZP5veBcLz2lUME4n2AD
T+rCwW7Af8oW/qSKaUphkxHHd91km4qPvyAe3I+KQ4XYAzqVE8gUAuQ8gZLXs6AB
BT+fX1gEEZ6iPOM0u0HmZAQSP7oYpYoLAyGXWpuD1WDzyR+jDIEBsj7N1BedZQqg
ZVvhxcjcCyQFq/caqZEo5OPM5c5ubKbzkQfL6sPAfp1ODqQGz58ffGYksTVuO6KZ
6qRy3fdz2Qi0bfKk2C3YbE9TT1P/2iupL9A5OWrqpsjeS5jLqIFXCgaiNzKc4YWs
IOjJDocjFFi1IH/nplLlTn4qveQiZPZnRS/j/OnjtkF9b3eq4OaMaApx7GctRqoQ
LOmk36JuHgyMf757tXzA9OrhYOPjb8ynjicFv6+VIpZH76kNvMT1V4ZRxSJGpP2e
NZVUkFlQ3ia7QCShW1u613jWCE85PscH5Spd5KrnZchZv2LoZLtWkGdcE1B1C12O
whcJl7OPA7+SCKJvM7fVDDZwTH2Ip/TU4AghAsZTf4pTzCx1HTgD95M4ZU7q+5XG
DDzkNYA7UrlqRWx019zA9VgZ6GBBXPXydsiYskZ3DeUyc9OG825EfS+Bv0UCX+dm
mWVVUKp6rAFxEcXzghQXfpWGX4TX9C7nJR/J3ReNGtPJbj7DWIBSDu1PnnG+85W1
vD/OS7cbGyB6EVnW9FrkRBN0HrWaxBRMrboEpvRUrqP9x054tgWuPYw+msLm1Ilv
o6+1QrCGFBMkrRs6hf1PrCsHGgbNpZy9Jg/GGQ5zbMhS0OY6Pk5YkxuYhJeQYLdp
UH5DNMThk6jc/WoCiYtEGQstY7rQxrot3q+VoUtevmqrEgXMY25vEUxIA2pLt/7H
RbO1hM8Vop6Lz6pxZLgHJ8ljT1Rf2Z4zqAOjjSY3SmlIp6TWIDhI/cg6+VbCty7P
Ut9ZLMA+UV5x1P3MiiKgT72Mr/vFD7Gx4AV+pegQhsj3SNfGIbZNz5iprOjdb4O2
TDT3A+0TatMmV1mUg5THxZdPe1bsWYWXZRtDF+3rmnAdteDmm6ph1pKPMIDYtewO
fYEj9GtqvxOvBLhOnynS2TtYtbyVnm8nebJ4Kqlb5ssn0zY5nUo9Lrpy2EZIw/J1
+/3aVK9lIqZ7vX+zMMuY3rZ+W++9H+8QiZK4M5xw2Z4fsLcfGHrpWTGBWG6YGe1J
57rd0DekBYYNc5ELvxSQFREVCpe+ujhMn4bvmE97jY0mzeLLJvK5AJaAZEOloSNK
NM+rrpWDavXE65F8DPhUPc5Neerw2iPK+W93OJPouEy2NQSemdCJaaoGO8kGAlg8
He4DtwBUYMP/C3IgoN3LQbmqTWGj1ouUlRWQtFne9IHthMutAdpAUaRRtdCrsYqf
ZtlfGqNFckxjtinZbqXW93WJij8Z+eupLhfQYqisJPfFt94wUkXCWN4yARKtpF0v
FHPKU+AeRHChL5VWnlvKzlc+A4t2avOYEXk1HGmY1FOoW5jmcivZ3swCE7NBH6bZ
giIEwqtT6BaOBTcESAUeR8UG1iFoYeZB7UXoOytNl89VJLqK3w/DXrVB79tQsNMj
PRTrdP0pqljdNxf7mGEFxUlKF6Wzc50AUoKTaqSJTBjSZrMQcAwu59UQ6YuR0V7S
KP1W3xMkYj7WklPEBVQ5YcGnAZlMVJWeien4HkaP3I/AuKvzlRuXOl34O6WYtmJT
Fv7WgalITObsqMtqQuZTBIKDCt8VL7ua0YUeQQGC5B0rNNiea/zZLv+Qw69k8b+n
3tl69EPy7vZZC9mqbzC09ickpNfkHA/u+79jOj9LMmcjfxqnEIhK0yXo4SHNCCfA
P7T32GUDe3S8OW79ds5HDblj7A4Te9KvSaoiJRqXycMe7pe74fi8vFHDRTr5VVtO
7Kt1ECO97HaiUM5yj1ORpygyQZ0zVzhOkIGKsFaLQXruEvQYslw2dJ3MRnG+P3aM
SBT1uW+cIuAb/l43qYCx5EpVHcOK3jgunU+Eb/qCWY5EOOVGmbpBJF44kMGkLM0d
HJgPtaI08u8emgF7fmel1wSsGXfgf7g2jyRZ7bkwYGDMm7yCnA5xbLsCIfCI/jdf
2lXTKyNUVs16j7DRGO39l1JrL8Ypdy62hc6A4Vu2Qmnac3uAKVO0nNCEjsuz3LbR
CEa2QNVljMXwkj3FmVkC/ilC6qx1i5hhZ+O0PcZLOhAoHbUq9pd1QrvcipKWq0BW
rG1nZ5T9Bqvc6k6XjkwhkcUzzBnY8JAH41GkPVXV9qnFsvMhLvpXWzBC1DaE4J26
5ERdHCWjPMgmMFq6/qzuFJ1NYG4zUKQdwnIDi6qYFK0o9kKeIMJLTfWnBSpHVO2X
IOWq8WoCTl8ufobS9AYFXZ3D6QM2o3bIcXChGCLonRAqHUls4spukBtvWYVUSVv6
OkFL1SXdGO/afkSY5C62N1W+JSSuB7FvIsFwpW1WwEhWPD+XWDk7Y8trdA+69iky
7mwAx7bGxq8JGil3Mq7pzmL83dGE2YQ3VOk6Y01G6xbNoCBq97ZrWeVpCP/hz1Wf
0M2OMAaYMi2DJWC5YL4imMQMl2ZodifNROTcaVPJB+OA89kNtbMYWXj5g2i0JIG8
96DiQS+5I4GHouO9zG6WsKU5FST7FAl4pG5gqDDAJ2rckjmDFWBOCsE4113lkhS0
XsFjSbfTXKIAyPpcmruxxlxG0o0zxYmt4a10F2tOm18MJh97zP0gCwQf6shUi++6
mJpcoGZRuEZ8ltkBTVG4bgLWH7R0GNnm4I8svO7/qjQUWnZUtQQIItNI7JS5NHKK
H+NB4YKod1fD+7P19BxFythBlP0ln4T6qx2DeeCfTmkkzUeYhMVzQx8ufNHGsO0Z
FOck2IoxPA9fRcOckGz1/2L/b1ePu/Oy+NZxx9ID/JAArXPihfhMAmnqjf9CFF+j
WWV1gWcBb23A580ej73Lp7KgH4LYWJ84JuIq9yBimcDVeBap2Q3AuCQwo4UUYpQg
eWS7Fbixy96C0X+fzCbWZU4Zo/EA5USyYh6zhRn5K2lu3kj2lh0ARDmIi7AKHoRB
6hATz6pkAlagWGf9c2adVcJv6HEBVR8WeXhGPlGAvv4NwlGCqHmxl7Hwnwt+wD0+
FC1CsYNMyPlT2e/Gd3nE8fi0IMCKyUJ/KAC5pgRNnin+VAY9JPxan/haoSorYIuq
T4oTSRZ3rdoEseYRScUkvi+DsjfDx9c64zDkNY8jywHtxHT5vVmLkEBPtFw36qjF
rqbt5sp6EaMNKzulCSbcCyDjIqvlJoVt2BBQF6PHjGBJDKth6KHeS+s7T+iqDhqx
MY2Q7TuAWkNAjg7njYD6xBtqQ1RHCSR6HM32LJ7DNAW6a96dcRazcPE1iEqx4erU
dcrzf0P7hgqFLZ62CY9jkRplhVuWN/zz2zideefqV7Tw5SiauQlrzXCdvJx6+qMF
N3Ig7sbkbQMcW2HJoNLIeX7/NEHUBC8GjSZC3MHB+ih+LUz6BKNmRuwBK5rmbrqK
ozplNZMjFO08WZZbNmRYX3ENuZsNy0hoSHuTrxlhEGjSQZ/rWOs1Q8eCLHNwZ8JM
1xvxK80KXfWBEs/ugzw2k3ppiL66xKBwTP0DTjqcGD5evo51zKrM6NWZ04u0dpk+
SjpB/iPsxMGloeXSmVxxJxyLy7zyszGoV/w3M7HazoDbfu9KMe6EeoRhXe7MXCMf
+/ZqTlSUmnMlMYwg4ixsmbtf+i4uNaIVz041lkEXTyrZrD78d1B6oyEuXg64nF+n
qn8BhpoQhyFirbMxF8Ivi3l0OR7ekck1fjhDBXChPNfYPCesCkg3ZwfBXuvIQE4K
tDzJ39awtFRqsqi0JMb0nTrRZkkSL0zzFo9wCTQ/pwueW9/MAg9laXPXEZ0dWYYJ
lp0R7t6wfa0SGb1JEFCsctGxGeEj41tIs7LfymwFqUZtIeSv0vEDmyUjOYEBxPMy
/Kkkm3Bje5rDK4MOamf+XMIvlCQnwGeYkfNYFGX3lSQk1R0cbrmEgdAVDGvVqaDl
4puPw5Bk3uo7HnydH3rWz+M2nhhsPq7KL1lkP1L/KeM5a9IXGmWwHunrcrze+hyf
xdlNoU3zrFZUi2/5qBDlQjjVzkHXA8kFGKg9DjplldkbuF6yid3eJeXZnubXfxCc
lU2JOjVH+e6n1r01Am/ubdqzAfRnxQttzNoWWFPm+1uvVb4QBcnoE28jT4chLK8h
he1wUt1x8PFaVzNyrjFE2yHY2QaPkyUxTgGRMzifFNMoCMYw0hA+yrcHlA/noXIQ
7id2AVIuM5SwDpbp2bfwunlL3NYCQgfZA6Cn0O02HwiZ26p4hjElPlINXy+vO/hM
7Am9UyhFOEEdFnHYtrGPYfli8WI+O/bgK4c+GuD/cHMDrHHJWAGhKISiOkTPFrF6
nCk+N+xPJCWSl+euDjxx7FEWxZiIIuxprrTLG6xvgyygZZs63Qp6SIbACPSt0k/r
MVqnvrkYmxPKGrBWH6rCHZ7hgrnIGw7clDSfrP3zQx7YeXcnnNOSq1qnFZYS9gsX
3GVmhtKI8kMFzOo07QScw7oilB2jRd7Y/9N8NJA5cCO/9NSWaNlEE9bRMr7G/bNK
AgdQOX1pmVF7rkNwrQzCjpyNRRwByq+SLZYSmhfkTaw9yJShcZT6ACDZO78Vae4C
YgakE4OJ+5cQ2fJRREGJb7NwdTlM90hmJA5po6jdqgwjJRJ0S6imJoPMNxmVFbJl
9Xc+vUIjYlFV1J1QbvYQIhYATYvB6/jYpCbi8q2Z4bu5ere22Kmh6m/Fz5CkoUNZ
m1KzCdrrP3Bsyt5NHrQGxz5oOKbSRtz/asNZUPJN2+7Alwozf+oRvNvsYLWdMZQN
Rxe/fqe+9tCsVsUUXjfM8mdmQEmcxAGnqkiQhyB/B+/F5nN/T19IHsLWP6dyPIji
BFiE77D1Osl+roNTu0nSTwDbIJStY/cmdflFtJ6kV4W9emQp6Ps2gWzk5rEMGGCq
OnZ+/SjRNQxpnXxPZyqyy+5X5dGsEgRw+crsm8hOu2+OJzRpA7uM0APGMzeBZf9o
6IumZHQxwkvuj13XR+vP/xiMeKnHVb+GFZ9/HCWqj7R+e7U2gypCuaqS2Wkcajco
5+6Ew6YeOY/XKJoggum0Kq92Pys0aadoaZQZVAHij8MY66PDY1p2QnMAn/OpcdpX
AglCa6R08Ex43sgySC2SX3hRUomVlsD5o8JPMpMz3Jb0mae/BDNMoHIbUlgvOVc8
H+8m4p9qaGerKlqk21D/k+JFhlF9Sr8DWa0qhFAgUk+GPBPgzRsYc6SW4gpLKAk0
yZzw4qqo3+TAuHJfL5DMGDtvaO/0U8sUzgQLLQXrqClz49DCY6Yb8cPNvHLTwZnh
yc8Fa5+Ee5WQ1V4tzgWwLb5ZXj6Fd1HxGYD4QHtEfPTp+JcEf8nAh1nMuemJZFWj
5oj20BolSTm52j1cj1FP6bDb7n/R+xqfsTcxQ9JeH62hamIcIfdxWzi1ExyzrV0N
NxQeYwNc9wwyk3y9P5UPpXQ61DpXh7ium4OxSx0xy+38oF7N0BnPKfjHCclnOOzd
dSOYFajn88s0Wu0ZDWtyfgsrb9huO1GIjImZ5MipzE8JO6RH1S7QJBFIQSyDF5Su
RhU3m3thETw+HLmn2dCJw0IPr9jM/cuC2vufgBv2RgUd6OvcnbAjNnG6U7e+BqXl
84hfekslIkv05AXloB+m7vmqnhr0ZATLkIGydJuPYQoERTPjWUIjtL/4ddabFWji
W14b15AhM7cgs7yYNf+VBigy0vJuLrnVtpgX1Ki1bSJG/vX+TFX/bL2OeD/j6t49
6knQQeo3FNAm8bk8ScEJaoDU3Z+mf29CWIbQZtB9M7CM+n56gDhowRDamWMAWRw7
na+6UDJU3eLBXWBJXpKHX6EKFQ67aLmZgZunttdt126xNPjHOiXqGZVhQTSJ6O3X
tT3dVxhVsJx7F7LXCDTjDiIRA5yfETFqRv6uJOKQ1dqoSK02+nGXZ4uI7A5gcjz9
fuEIrzfElT5VTQo8PRjs/Xrv81WzmLtc6FLDFIbQEM10sHe4teo9DaA++09IQjcF
Ig/maqdGJfpQgcghe4jJi/ZmryrfHJhbBoIGbVjOITLHxfJukGFH9aJeIvmgRTU9
eJ7MhPm4RAj8kQDbwGW312OZx2M3SLr8qDO9pX5/yq6/lF5bULnIVsc7yxdYlwRs
qyaTQ2PQOpXevxQrY2y7qjuNLD/7Q02M8te6eUW2ZyvV+0gWWrQm0bBtGnvpxvKZ
VfOCQyGaM6kHtD8S+79fb1UDn2I6FkVy1YjU1LlhR7SiNuTn2GoGgCgvOL49Ycux
AmxlFLrVJOS4U4tw+hkcZ2S1eXzHqXeT421VKJN+GFcGOZFYbIWdQOUQalacS6nS
OTVDjewMc/r9MBczPk/zwMbfhU3j6xItKlyABKM2mKcxY6BO3vTTzgdrkinlfFTn
x00IrQdOMbHmPCjvFTt5y6rrg4A6N/GM7vk6MfLQPrkU3xu2LULKONNOaSHZ82v1
+T6oaE/PKfeHH6DBTT5ghtK1ASyrWuiIugFYNxbtqOIDv1iSCv7T6wWmZtc7QFVG
8sToirBrHprPCHSrflmTtmnxNHrmFz6im78KgNM8IZw984TZnz63R4yATAibo+wt
SzjHIFSiGQDG73TW74VdgoNBE8Z80kaOB533U04u5667YWmSbfwqVOH0bPjJKP74
bqm10mgaiQKWHr7Gp1x77BXZUz/PoDD4dDnAAS3nZLsl2Tq1t83h542O1c3F8Sjq
J0ahZLfojE9/Hhg0OR8tyex0EqQxiURnTlNUcWLuuD+paIeKN9xY7kJ5/xHSowIn
n3jZz6p+ywgbByRVFAgsOiGXTzeLIqsycEp1S+DRcsS09lGaDQBz06GZHLYxnjhT
fVnLkTcssFYKd2wyqKYnYQSrl/HWWfsjYFgt9D908jxPZ5B3D6ifBx2hLbvfmlYO
C2dptDnPd4DdQuJHSSDYLZRaArAJZ/xitt3QxttL7TCF8Tvm2Z7Hx75p+NK48RhE
U+P+gn08LN8uumcE4w4R2rsW2pCqcIo4sCV383dUWSekCzG1rQZdZhy5UvWa5x8Y
4K2iVAJR/yK++1pzrkjX/YbY8K/ocqzcAPKZn/UIAB2MAGjBjbauaOauQz/BdkGs
sxL+0z381qw1hJjRK8pgda8L3RH0PAmUSoaOmSXG36Y8rgOSCACJA2bcQfWcoNpr
MhtGF/L+Q8XiUtzTB5gWVFUCQqMASyYL3kbcpnYTlL7ln0b2ERDFdZePhUezNR0R
NtBBMpayS8LgqUbGggi36nXCmEQbmMYEdhk8Z7eQhH1+dnrJM6ay5NeWW67Sg5eU
FBpq5751TfnwqTc54gAg6IY1VUgPE86l7L2/BTzOUVHMTCk/O008yKfQsMMGmkwt
NPyKjsiV5ku110VW8UId/OzH3JcEQTQZEQh/35qPmwwWVIHLTEtQhCPIjqOyH3Mh
tp87GPKa9YcumS08zOw11vDEJGUTpOsTUp+QYhUcszIYGSc2DTMUugwudZV/zx8F
qOmxRTf2WqRETxuxB+BJOzCsKmuFvyq+3vZHyqqjZ5WmlnlQNy4WwewAmgRUL7b2
PtQ78nOP27kkMIOylJYFxBgKClYMwmobByQmmHPVVjSUmInWJU+IQ0Ti3ZeZAn3p
N9gucQ2lI2cOucbODw02ls1AZcexn3hc52nDT8UBQFPpEXNlej+zIzvv9UrK1uSz
4EPUY4oawph/SiRNPRSwrWBOLkc/yKz3G8jqKikqbTjKPdUwni9asPCvvn9e7gOg
FzPD4GjUwslA6kqHmzTO17naT+FcY7cji2TkEWhK6wVIiAA2M3wfnImBWuEWyHL8
Pg0Hp68iE5ngwAA0/9oYxE36T36hsuZ63/hoKpfgC1e6djXnLdWFmJZG75IrGX0H
bZTaO7JoGmr731j3uK4BZCZCsVHlhw0+d6wBuxxG0vQE+GV5H8pbLigEVAR7+eXQ
TUjwYeB0aTp1gRbOzP1PkleVc3VciaywwrWLJjRLXEkQPeg/4pwtqTMg9CJFz/XJ
2eh6cjiP0BPY97aevQGHmGycX4xHP9A4KifBDYkJU0IsfSqSg2cBCgdUFbsp4ppx
rfirhIqCxHVYTK2ilCrl8kbkkNsILrq4VQp6LGl0GhOrShEI7dblohTtYVmbat05
K2c1WL1sJVHiURGAo97iybC925NRc6F3YuSO54lHy1k9xQg+nN1qJ19psC4N1r6X
pebQO6Tc7sESCENTqauZmCXrrm71DNz9C/Yv/chWJ/mcsJM+L1299aJ8B6pLsduo
Rc8BCo1qavzEJaOuFJTMGSqoHl1E/+QVOWoXyX+O436voC4evorpGvYDumj/GoQr
O9TEmVO6CWJcpVN2V9p8vaR/7dfkmfiTzw82V4W3Fiu5bGRSb74cLXgwcieIgrUt
2iASeXMXD7+VEYquMRwJouchwE0TCXQN8/pCBatCGb/yfmFmOYAB3QmJKPmXXpY3
YE5UTgN/8/rK1xitP4gpu4tQhSY8W77VDMSZ2QDt+TibAHoLVgekoupxotVDQ3fO
rGsjJKEhdvm0sneb8iL3HXFOt5cB6+hM1mzkY+xZDQRzriHzfjj8T11RgnKQJFGI
4FQ5xv3EUOWFt8eZ2aL+vZlpZqKRbbnktcXefAMMf+Vl1lwbDA7yGUbIEWtmD6mU
T5eGXK7+w4ZKF2B0MdrzcpK7CXmoBlydWsCcBnmdwfPJu5Xv3iNFKZlzX0SlTNfx
bWxpz112DnRaAyuv4ShFa4opP6FeapN6M8FwY5t2QKEo7xnLKmfUsPJpbLbGgTWU
LxrOngnvNT78/sW/dtd3Jj0pcMmYI6CwgbEVyiBKTyJQ6hqZ/KKVxpyY2mpRAIva
3vbL5qDWTct86LiOd54ktSUo6PC7bbbvb1r6K5VX9ny+/Enm89YYi+cJ8CoQJtBR
M5k/A2Y3tfrGvAk8C8r48n0ZyVTmbDUooz24B1if1cQ2Mg2PE6UebyDEnTZcrImI
LjkvPkYvGLiN+d0n7EoQR8Ho6UvkhQ50y0aW+EWwHlQaOdQnHuRNuN9jRBegudOi
0EP+JpmpLnYalr7BZHIRU8g9ubAlbLR6tVwmD+5vVyh0OU5vUX8I8ekkyijr4Obc
lu5ZzmoYSZKa/rzHgO0AOZU9syGSY75Ywh5hVpMngQ8k1Ajo7gjHVArh0+Zz3nNA
pE6hJCGLUE8lTs02SKfvdiaQAF/YuSjkKsH6iBhDMijiJzdBYpxWSd+gAU47tx+O
tsu3KhXULkuZcqrBE2ULY63H4fU1PSCt1TBGEMfbRrMbxkPxFyGOYC1R/rljq6aE
wgLQXkeAi8vwCSAJx7wEygEVyt6l3RvNjnJ16IDp2TRejUA3ktPvA4zEo6L57XG4
IEaZNDcfn3mnPcj/JRfNgXrzjeIn1HLgRSXm9GbfxPtelbr3q5hOa56V74zgYVTX
P64AJbWXZ/Ck0mtT9T486TyKMpgc5E298M1Ut3r4/XoOLQWh7poXZDcZxL/gOTm2
8T0zg3209hCiAj6kl3MBZ9UpLnuW1gawx5+p9Cdir+40bHHj3QsO9Z2fI69HBwrV
4ahAy69hm9qj3hs0qzq24xsDfFdFjJbpeCGaRpsOBv4poMlTORQ0CnuhY4WPPFtB
9+O68cbUt7mXQCH0Z0r/6vKCzolmpCu1iTvVspyaRHm0BOKR+vgTbMUBrDfDd7jY
oc1rkYjJIvEewmsLLyL7xwTIn8F5zJTxfLC97x7SBOtn5tKv6bI51ADcK63K2auM
I+/clwoMxoq1NPC4ClyA0osU97Mor2gDwX4YoRvhgdPbBSTSrx26XrybPpSLon6k
8h8eZIl9tRBKmvG284xzk3WHdZZBsa5O/D0xJNq8MSuSMd8WZKex1VdGybJDRvnU
FPCCOPQ+sftFOFPkE48ALxMej0PKgrepZzKbHN1VMBAqZC2NlKnI1F47SgtGTYFw
7D8hCx0z+5d7SfKCM8nhCo4Wcs9Xu2LN8TQ+aNNoFaOudJETSJWRUm/mxKjb/ZLo
e7R0l0k8NeoLGzMLT7F4k+b7X5NvZTX7ebSStWnpIBnYypsTxkoBplM2fuNkWCcQ
WY5t6wEtFySzraobs93L60GBQ368nKgb2Sd8AqROTc3A6MA+kw8RVt5Ikp5LwReo
J94segH9cztZNQtEpwNXDN8aKr59JoyKRtakm60+Gqr2LBbYTHcPZ5UYGwCMr1g7
Di7qeXCCdfUmtibuiNcG4PSVLr0jxHwy7oSpyzkMADa/u9bXJww8u1o8Tq8UisMc
m4tzVmcWkk3xm+TVEQg61YITESPAA255Kh6qRteEElrAWR5Wt6WzhG1LqrEUDomn
U0c1XlqmdzY1rj/D0HqR8LVi5NDFB0LRNntLxtyeGVCWdz9rLnbw21Ac2ukj/xM9
0hphc5AYqJDfz9OLmzFN4EzmN88i6clHzjUQzLaLgagRvi/sFksB7Y3dnzYYnBy6
8Ll4Qt4Rm3wYkSNu6ct34WbB40clUzs+P2egXmkkBfvCEHpO9AjgBFk5J4lxjfG+
0p5ZjCSifs0LZvtu4hV5IlZgrLJDNCUuJ8j1thn/kfILi7FaJDofTS8gYrlOebQJ
dlN8w3HCNyBumTqBbtpW++m92kWBJTf9DlfNDKg7SlM1W9XQmC8/EnxU37/0ttCY
Sm0NRNkhLl5gg2G4N31cJW0z31UGZ5cjyOx2S9AfTQbpS0Q3UqGayUv7HY7/STSJ
H9bOervUwa5c8F+cN2Vm6tJTkHU+0BDFX+aF5j42JqzmiP289z98PUmm+mP8KhDX
Vy1P5fuNpOSNv9D7OQd/8QL9idOQSSLcYQsoQD/1zLyxLFk8MkyAkjDSZPrPC7F7
tE9PVw8817G13RWFvJu5SkVmy30SqQGqbLfz1nZcJhrIO3UqhvV+/yoBCxApreHc
CUmuxDro2w/rss69YfswpEzn3j8tUYJ+SdH7YCN/S6M7TxFEPokM8TuyEARaR6jD
fEYqvhjgiqk1VlWz/I6stwhO0tr/txpwlbveTBf5MM5uvcpspiUZhb+k6I7zPYm4
RF5eSiSIRxRsWl6nAfEqNEhemoW8+7/BwPzlzkkUoviT10zMz++PqhgjrFyDNsIH
BsDqs8H5+dsNaEdqwYG43ikCFgYsb37JCwv1/OBVvv1ak5eKJ2AKHQT48brww3/I
ab3dVTbqHlc1hktzze+PaAhWEFBvBXh4zrXXHEwUgQtAoG7QLvRpllDEnI5QjGle
0z39rddy4PTZuIbsl2YuyQODY7Cpdiyfo3GUiqgZQx2LzMI81P5iN9ID9yoaXe0d
2Aq+88CEF8wIiZIEe8/fIDa2m/I2a1nTmQbmKR2m2vG32NVOTBjlKAfyYF9amdn5
UppjN9r+x5R0nXHhrZ8ubcSFiz0WTng6TrVNAevsWN6w9ENyeyC0r+EUxjX/p7sV
d+HUzxMmhPA0zdbNIxEDLqETkOpojwxxfHy4xvGh1nk8mHG+HSflgZx8GT3vIGsB
yDLLL76xAspYZ4sIGxRk3/Jx6WsGXnX2o7Q8JQU45ov0dU/ykLLaCpGXFW7MYZqh
MnUA/O1fa1l+DPnbTl1Fqz8GtJWEhOmBNlbwFhVACty55+qXpMetY3X9RVA2Z8gC
LHoJ7Qc4Qx9mW3kydy7L9A7rv8UQQ6Wab70I3sEtXFw9vuYhx1VWExPpSE9lX/ws
cXAfMBTQXKHbHOnRlLV0Tz9M3dXWfiR+vKkm6IHiUIbZxAER8CKDm0eoeLmgIyFM
nR8B2h3Sa+4R3VSek08wRHKI39eYUUF482CIPeVvpV+Y6rhm9DrXUIrejAO6CcTz
bDZv1PLoyH0m9hjefGD6Ij5eBapZ8JY8uLbI6ALpmb2d48Tart3u9pT/BhGr39Xg
VDgcm0mCBl7jvMGeR9IOk75vIN0oa42OV9ZjJJe+N3PSKPHcDFNrziT/C8wal/YD
2FXlhdBqKugxmV/ahR2k1cNKrr4QrFQhEjEg9g5yzDBH0OFJlsYYw+DROmW8G2X5
xNPsm1vtgHYLbwmSNhwpE0mvlBcOWxcRVDVCLgDRCLah4E5xS+OxorL6p1ydfV57
9fg9DVCXQ6gT1FRFgmYsySxlvdmOCBfAJlLxHxX1DYv2wiI4gGHbLIpPAunsdzJf
syZJ1lVNcTVFovc8DF8pW8SbTpIV1KsaK2cdqxz4M5Odjb3OLfeVL5YH2G+c7j9q
UNLFs7rwuxuKZTfcIFVpRJOH+Ur3dzUEzu8RbdpCC1GDb0EOBiPg/14rE/qcuf60
NiEk6GaEnGGrUD8klzz0wz1mkXdfVXjrcXUMP/sMmmKzOpSRtj2i4TYizkISXSJ/
aNMipjm5irBllbYd3EZuULKc+NIqkJmBRtDdQp3goa9DtDTLzSgaEx4ndfhqkPsK
LyFoMZJfgv5SjLrxfh2FZ3cbQw4tGP6jOL9e2mhYuzkHPiOFYSc4QKP7g74vSsCw
n7V4kcNh77MsTyTZZK531Mk6F2IfuL0odMF5O1psaD9cetp4zIywuNXvtKrxB0yN
qIa1TgpS7C00o9rFZJzzIg2u5mOub4WYntYhbO5ISaXE1tFbK9nhvoP0SKURh4Rb
I5VSKz7/EqMooLbYE//8nPHqnC70mZmToFNCm1vIfmcS/CIfACoD5hsTluEaKDOC
3/KANOskqlR9mWl3DNqQf+gY82bT70HqWzUGZlnutERssrWnB+RpKxy9vZgyC5K9
d9t3pXFUS3tMha3y+jL4LR5Jtyy1mLT2yscs+tlgs08WGRbxY93X+OqHml5gTL04
A2kcsBcqF47WBHfJwoxoRTNoVxVxoFDC9KbtOOs6xM8ZobOnK2Lavxzv97MEMRGC
cljKzXoNaJg1Ziwx/dVZTfx/xFsxNk+M7PWq9m7vYuZbsHxsGuQ/+g7HVqSZ0o8V
kjqTEtn97rTaHHA8/po+kJq/4sJewvMLgV+IuvYYCj7W3XsTUrwT+LAwrOkxQ67B
/QIn31gxw9VVdrXSMrszoCZ5ZdeE/67+TkAbSFOkK42u0CyvHXBMVQwJZeNyclb7
3c9CzIpxygCZoOAOVDkekU5Fxbu1UIz3phTH0pwqmRuxtEe1JNb++f1K6wmLyfzq
ERMIWOsJ2rRI5hu3s+RMVMcyxYwyPlYQPHUcjk4dq10sk7TE2O9d9FlFCeVOb7P9
IkiostnFzD3zGbYe8VcIiZJ8IsYSlzoe702rDURvbnyhETEAWBee9lVTLBrgDNAf
EN24IBlY08pxccW3TwXrYIvVWnapnZ96Bijhmt9PPUi0R1nwnKPQt7RyfFHDPUDo
XKZd0VFpJPHCKkTNmnCE01MvB4NKieoqMMFTDCBfy7bfcXa4hHvBv09ts3oMFWqm
+hv2L/hlfU6mnaD2ZwJdzkmlzYLa/Rs+MlEW+M7w/ywYvSgxfbiSxiBDxnusw9fp
WpBD1nRGuaNnoImj8s3RUbbTR3uXyKH8dhFeNjq2iZa4yFpTbYXrB2LZoLuw3gNV
1cS6cpLOOy1mqn9HD1r06lw3nUAJWoQSTmO7pFrOehXmQxudwlz308Zd/6rPQqqr
GB4zWU2fQ+egvyfYdNW9PbIbG+1IoIsoXy6/xbnY9Qr92vPvQOhtEiz6dylWfr/9
0Am7y8ntc+mLwOQCEYUQocIewSP4I+C4rTBfncGltJew1UuxJKO0PWnCSp5vNYw+
70zLy034aSSzVTRqUYuTbFhl6C2B+B5v5lyurLsGB1KAY9Wvz7GcbMnhRfu9udGt
ttUuOovBAjtG98J8RWF3N99R7uIjfk+jAuLq7HjUf5WDFjOi4keLXk/X9GdOJZ3+
Tjrd8mws9/c6VPXEA73d9i6fXseBfV58+73Q2DJXRhoerl3RMCnmCaqu0D/ogV6X
4PU45wM1agoMejY44oXk40bDsxznJKIWoBEGMcW28BtXl0nNZVhLZL2WY/IGVwgI
YALqI9301iErDSLbGiA9TxY2mQMW79sE5QqNqwWegpunPMZlSAZ8PRzLEwplfPjb
ylw0RpQj4nm3MzptelF27MuuLEr4VwsMtqcEpXffai0xNwIGLfCcfvW9hu1uA+N/
W7yS7RL9Aj7tpQiwsEvyx2Ola1s8RRb0VUkju1/f5v82+xHcaNZ3ob+qixU3Tpcg
50j22s0lNOBXdEH2JPQgJwRAx0utE/uEAjiRpJUTsAeTd1QvQqvQXZ7gTjqA0hiU
P8lxfWLhRo2AQQ7U3gWe7AUxXsTuWPqHARY7XNgXNizaMb95ZrFF0Cp761MfRfvs
475iPX4pMMFqobYMcO4ycmU1nC+2FXlf+xckcEx9Ed4ofu8+ra2DhO8CJv5+ydDC
+RQquirHUCUqM2G+JCojGCTh7g/ulxpGa5IsR6z5f41jRGBLNz2PFGg4P2na762e
v7c/YMEPsxbpW7WKgBq527FU17tAA4yAcVf8VgeKmamAKy/DOEEQjdtADUktIl/T
XjSA1Jkzc2tlfMXdehXqtCcBIv73hE1vQQ1ljzJPlSAZUHwwQPRfY2FMaVrFCm+q
5/bVIw+vLTjtt0MOmf8TqihJPscSZc4gG0p/EksjMDhuHDpprpAHYrvQJQtSUk63
ypCOPV1eshnrNdU27Pcsx2nzFnRx/gkuKRT+6kzYHbDBBtbS5riipAyLX1iexjBw
b2BXfC/31ML5VGcboZgc4iViC3XO7TrGo6TnMs0xpQHpzhjld94yTR6l459GG/Fw
XOtnJIxBSztufqt2MLjYO5qWLXRFyseU6sHFeXKzbZLlOZSbT458/ugX9W6izj4G
NFtxm0UMIV03qNVqvfFqjubm+iSFbIXMb6rV4TH2T70gtC75KfMIMxU018/f8vgP
AfQLIR76GecYQ1NistFWLAWW6TGly8MaeL6/IJ4Uowg55Yn672xB4JJFYxpViaM+
hSNodBxNnvic+A7t77pAaEyuVDXhYz57SKiJsErRM8aCO/0QxydV7ObIURS4/tye
gJsdHwZtOlAANcxLAcx2MGg+zqMX88jjfbfMfyAsVGZAr1by5ZjRO1JsWfCQcmeH
R4Agb6Sc8geJdBIkhSeFPQ5uKoARnr1YnIGb+/ngs2rmErVGCOF9Lhza2n7paztj
ZoS/z+tpDMyccXlFMzuLaD2n8pb2yMi9D7UQhhS0LEbT6iDmDJjDziBXfgNgWlpf
ifsjg8EeSDXvcXECpqTek2S/Dw8N6AE6xqnQsGNYCaNywhgOxEPcB6IZY7Lr5kb3
TnEIK13xPwHMlnhltNbn91TW/oyOVAEgokRx0zyVTxWiDAwATlR9YMnRHP+NiyoX
wRKTaNrF4GEojhdqNJ72G9RrGru8dtD5J3pOz5aD3kAOwIn8MZkr0I1nzgj9bIp/
lRKehLj68cWEmREcDdseE6mLe+4RUGzRiaXAo/blN+2O/xhBCZACnGI8zic17FWe
itqZqaFELYxuayf+4VCF8hWLe1cI3XX9WbSbSgJQ3K0sr7uda3UNePKaO+ZBR2z1
ETroGDnujw7RjAdgNJjCum3ZGV4OojAjtEv+kTdp6wa7WAYleAIXMv7bkX9Hy0GA
j+MkAA4RCUDMj8f5Xj6H+Z9DlQRgG6w/a94FZBJja3m0ThzbFLpfQzLGxiuZmxPp
HTeJGwmxj/maHEMYLoAbOIYEkwUILZG2nfNG/OXva5IC5sh/SHKha/ncN8Dr6y/n
eDAFPPecy0st2mOvxsUNZbtc0BS0/3zgi84r8hBpE1rRon7BF0qjL6isbPZf/Mfz
cGohBBvurqRHmaWNW1JyuVDfGLXfhJhebZY1AjmskmRehmxvGFj6/abHo8Aq/DYG
AHK/W7iVVrhuO6qa8mUrX1GLcwQk4EH7XlHmSAih+qjWuUNbUKOJpQqu2AN8quPQ
RJInsM6PSijsuqeHJqcDm7BZHNj3KEfSexKY6X70EA5pxVQ/pof4kszW+nPy9SVj
8k91BvIimcLv8sDEaiMPnttMORJhPgb0zpYFflfa01sjLOwvxebzCrh2cZC0VByP
OMlm/HOx1Dxh6Nk8ZPfzJdGK5tExUV/2TJsYXWISzE8ZHzuSqFY9p9IhxOEkpClb
rSoJMIme7YF9GzAdPdgj279o7wurusm77COHLW6cHq+daXjxMDH4dBbjPVg/mVrJ
2RcuJQqcfp2woyriGQfSf9ajlky9zKBb6mbdYz3AZ5VRSDUA/geslfrVrTOFQoBT
wBJHyADTRNqN0dZMxsQGTAVYcnLQQCVl7xLiycuD0ZLjuNR1haH43sYljNy6vv9Z
j4t7u5vY3RJ43t7PBiUf5cZI7t8rm5LhBaLWKUMkOHgeulClDnQHCXRAjfEVq0Es
W5VaiKQw614TeGMd9Ta6/vv0a9iLi+zWs5EsepA3zXN3X7uyTfWIWuFX87R9Z9TJ
55GOnG1PoDG+EuPY3Jpt421kkO4izbQoVMPMmQzDDJ6Rd1FD4u+yyVA5QfawHha/
bzLQOlXLwDt4Qks1ICB6nVxTfwKKTBJ8pQSpGEdpouMq98KGtWjW59kh5NDNZG5w
8/gfRLq+qEwMnqRKfWhQ7+mhbxTVG0AOzBJXHyHBCHnjSDUNc+6sG8T5xj3QlZe5
aD4rgTA39ReAFkax987qG0BYxtiHzh0Eo86rif+1B+0AjOsawtHBsw2QNN+5SX8f
ZW8St8O5ddWIV1QdhGCowUzrqTRsffhwFAOog0LWHSvQABSnvNWx5k5Y8DBGDCL1
Ap9szxm2UGbwcIv+PO479cJnxGBAlkSDOtGTPXXAY1YhKhSIoO86OddCrVUtu/cm
OdM3yvA1vfbUGsCgWOZyBXcIZKekl13lVPqCEMtPnJMmqPkBS8koUQZtFbzrNKz/
KdXs2BTtwQ9ooc69brHc10YcVVINqtZ59NduOMPF6GoBweLJ1SjijpIuusM0KaEa
PV2/SJgbDC3edSicIu/BrN8MIIkcUc9EbSNmMdWVPIE7ECrIocJyuOXJiZNuEP1Z
bpZewQ67M9pCIAFaS14UxKWzfwHFvr6/01n5xE5sPbhjNYG2qp9uBn7HuXjfxmgC
tYhwNafEQYqlTZW9Sg0VtQZc4tlG9HNbI9ge5OE5mEoJ4TpvLSaBAgqVkBFZpKk4
uHPRrU50xDgGxm35gSDeu6Y2Qnya4QgKSGx42Abyn3sYVsUFgyBcpMXn2Fn8h9y2
uFjn2/a2AcbMzPGGxzTA0KvhG7YDDmtuGIY+8uX8yqb/r0yHgp1vKqzCnyXRm7PP
jSYKiNsjvxPniIlIqBZBK/Tm17IUCEvoK0X6PIA5QTZ8c9+Nd1BDW6JStjIJjjeN
pUvNKJXh0roHMX//hAS//is+bswv+iDPgZf7QA6YFOaGFydv+ABGAgvxmtvzJKRj
eGzFJUp6zPdEzA7L2v9WnamDIud1ywEuEZgX45fPKS4XL9JrHDEya7r8ibCdDBWY
hEYqhlqAaEqOqnm8YReqMOfOixUQoA3GpAnRSFGB9E2mlU2Z1c/C6zsOrJfgSIZY
GM5u0dqGD8nrcOygtyZtW1KatNT820S++sXug+OtYlsiRp2nXO7KnNuZjuTVHL1w
6n1K7flEDGi6dSFSF6QYSLuBdQhdjKt45sQj80EalD5j8Fxf8VKi8gev7rUE6ZQ6
FlOl3tqdX9zlfiXOyN893meuMctA52LrHaLW0ov6NhL6tznvntYjTbe2sw93swHg
z3D6K6TuEk9Qo3nJcn4mCHIyNjV8vLbRDZxqNc2t5JhtpvQ6/Ot+K5+BgTVFCUSg
6aU1tK+FrtEU/gxb/z7tbQDFjekQXZJzk+ztbQsNYvZ4OpOZRRWkFryQanznmte8
DX/W0OF/8mkGCW/NXkNM24u/wscAB0mrnyVWFwjHQ/wAIqn6AjhXAsMZMzQTezwi
t4rS8TX6vV9bnEcib+B1YvgLD47petU1cxnz8FpOQRXUNijeqCQxALlbTz+bs6Ib
MVtcc043Xq5+3szwYxNBBpb80ziE4GDgaRZx9g0i3rD7G/D/RcmFgDf6494WzNU5
CKILuq8zZ49PYpNgT+6CMYFHZaWBZGaASBMzrFGGZezCPFJoFBGm/psAbDLLeoNS
1dOdMZuGmRjrLN0rofFTN25BI7XZtmNKMjDXd8gAcACG8FCphky+kshSa0XC9xyX
0LvZdhNIKgqGAqHG1tXHLgRxrpzzjU2r+qPhBnAOotiFWbPogk7Pyi/AH41rxMgg
gMa3whrClyrM7kAJRrDKEvMozrIAietqmr9/4pJoX7fYYo5R5CW5RhkYw/p+3y5o
pgLxI5RiuFMfSCXy2cwFvDhDnpjOIj3gZfuqhMZqXf3cTOqG31LbIJoMgDaxmJnt
28iw27BsduIBRV+rYiCyyHD35Pq3vaQD+WmEf+vSYIfNl05VPZeiK6h+T7ZQIrM+
gYRz/W0at7WsMSIal2DApu7g3dTDTUshZQjd7EPTiKdoMZZWc6acEi4p5vAevLFo
d98YY/JE+E503t9kZ08oZvhPOvZMNMcdySd8fGZwHITo9TnkQ52xCxWheH/F7f9q
NZev+0KSE0JycLDqo65gXEnAM/WWpNx+qbyGUtUy2a8gEGglAsT39qLHjJMsMPGR
6JDtYun4QaK2RjPjOuo0Wgf2NzxCDHnJQOUAFU+rdFYPThX2Hs2opzJaUdHJ3T4G
eR/oOBoCrBlSER9Wm0cR0JdCDPjNpBAMmzVMP93fbmqz4q5rG5liwtitOijOq8WI
fWcwuRN3TcxvnTurU3ji6f53zHMw74M2vKgvlquxivw2x22CXFM0o4r/Om1YqKQi
dQvimwojxLMEu0Xx6VcPeK6e7etDWgTjnWKfg/p+RxzGYBPxIla3I2yu4V62nofE
Z6wD+/ZAIkJdnWH03ZtwXmeMAdmBlSR/Yaj33DlUiFZeks2nudqN479+BpJNKjj/
ovh9JM9cK0dJ4OdBUyMHZH3eC7rKl9WFscIgE2jI8Y9VH12r5SjRX7cbj2qTenuH
ioovOh8puN23bU4SDtmzKDwnyjvqJfJKYCOy6vEJxHXo4X29tLVsrlgKiXdvxcO4
PKOHwIpmMTYy1JI6nj+hfyH0Ve0rPYLmi4vJm2iw4tZar6OiohPmxPnlCNxiWEaO
gVmIKK/b1VTFHaSu/U/+MXPM6lYHcx/u4kDxc+o+E3jd6+YrfJDFbDuQHoPOpVtT
gRelCJKkp8LFTnCcL9to5PfjDRszQJgWJguuY9HqqT1wWR1X75lc7Nvnstmq73vg
THCeiOzBiR2BDN1+AKpAMRDzJkAtEf20+V2FRj2oZCkqwrBDofagHlAyOxIy3J9n
cdH91xa+loUkS/Hn8HxyFbMbfF1o9MoN798RTx9etbHWVLYmH6JnMIkUjKKqjKS2
JCn+BmrdNNUNkBllzLTVgdOGvzTnKKbLYo5GtDXskywy3axzT5hAN0v94ib1rZw6
voy13rhWpk+jxDSU8talEac8C0wzUiwl1Fmc2eZ2gpH1GI8SAPpDt09HdxqjVi4M
kwqvr+JCRvOWKA0/A5edd5hnvCpR3eg8mUXIwAM8qXmkPy2sGOzC0aSjfq2pofqA
reBcm/e2gHYChHbZbeW8kk7zi3trSSIXrgWo+vAFKCY2iPAOIqK/OGZ0JpbY31AQ
TI/znpGiQTvH6U3X1CdZCDewtP27OuWuHW37SYvnBgi2Ms36sB3VkT0ZzcL2rroa
9D4vJUKfRhyOwHexmFJctli8OiPiKlLxssduOnaQtlR/7973y1rQjpIetsrJBXJ4
c39K4rlb1uZKRXwGuV6uD7FqVHh2NvBYkcH2qyzuksnsDCxBuBsQpu0SBiA/yH5G
Vi/qbUWyMtzdw+cLPEbcyw/Y2HtIMoHAJEFKon/6N+yBLHc66p3Esvptes1Derbf
PhVeeg2AX/Ux4IFkCV5Jj9CnaLa/+MiftcTBsGeiiQxklr7h7fREBn4A5lw4UlMF
MIbWoIfbOtiVNZYUpQjcl/bGIW1/r1K9NlSV3fY31TyFO1ne8TwlA6sS7pqSq5ii
xG5Nk760t2Tapgk4SHtzL1Svy4DChJTTac4epyjYk8JUX6Ec70/AoF0kGh3/hH9z
4SKiqzMcZmtFUYxwm/HwrX15FOr/uXMf+ry1u9tHJSNKW7qLTF6xVfj9TSszEDrP
D6KOk1+v2cdij95w/dfhb44iOwbffuUZlVQYbz4T7624dqz6x67gxWScAfbWiew7
UFYuC/3CGRhPJs5Ocj67ngTDCY8SIYHi309OFPHIDVxrrmZmHaD6/8omfrqwYlh2
RROY4M+PC6pBDOiEis8wnDyVzRM8opxOUhUXyP99iGTl18+TwyiDaaHFLXydyh3n
TzT/nZhwbEWBrsn9DMCT4ehAS8W7Fp7KTaitzv4NIi8zQ51LRj6jrsjDNDDbV6Zf
lpRKWTsRc4IGrCWrvFmxxH0vScFgJ9wIlN+ZsGA7C6CgbJMRXmorkTd+8uZEMIPo
iaRtohyFDj3TTITe2K0335jTzaiVKDg2CoKLSlLO1N9T/rUJUr1r+Ud/3xOlFg2A
C8Ve5lzmGQV4nSl/ebie6WF4lKM0gulxKeXRnViAjxtjEg4IJZIRBlYeiV0dFImw
zGFRtRC5gBPuRP/idemPjFQ/ZLKh64wxBi1iVr+YwIsPRSEOrAomDyV/L6narQkE
eFdAIgg/o3pcJF7uaT8Z/4I2xjKW9HF2Gz/OIxV0YdbS45u3GT5UwVIopBKPUoOe
9vyH4r6X+TkSOuqv2LVz25ANI19pfrb1HOqHvXn+koKc29wiPt6kHKeyOg/1BhUg
PyeMxOEhCa4GaFoYjYxDWbe0sHQ2xPnaoqrgK5lCd7n+e0SCGjEYjHsWUAjpDrZp
+FKiTqflVal78d5iyJbnwcO8y8gv2NqZ/pRCjefA0eZDeP5kFR7dpF6j/vX8z+9Y
KNGyhx0n0w3sktM2ItT+vXsPb5BqWrX65Uz5nvODwCM7i6s8wKALHLwoBQdMhBKY
l91wwghQ1y1wDmRbo6ihyuBHVr+pFuafS5QvayOlEYkY/K0J3og0Qa9S4gJmlsE5
f9VUmyElJsQB3RsGai2gR2OopAeU63SnsRUElXOKMt8mabnBGgQQ0Q0EMUwTSQyR
lMkQDrCd+k6q3PloZd/IoDAFnxuHbIbtjd6jZTtobW66+Ot5tg2zdG/TEoAeIyF4
YjIvigC+whqzYdTxp/c5sc79kV6aKyw2YxYuUw5znk3JiecSnKZU1Z0IyeS+fGYC
9rY1KgFL49cIVKtE6VMGwhVIRy+Nb7yXxBnWm969lIYxMk0G1L/qxsynC+ztJ0Pr
GhDSdJcNC0+yGK4fkmL2XY1Wg+5cYeuWrszfxzgl3irobicjeAl65FpOkgYqjZZY
+ZKgys5y/D7dxKSZAxWDdAZ9gW4pM7XAdeqgMOq3PS2VNK5L1qJHoncVrFRRb/PP
PAgAvQCe+FxMGx0maTOfBFQ2igvkSGyxwGin5p3lm4b2pM6c7Chzr7Y7uV5ZOo4g
PBhyxB/4zJcwaF4llDf4c+TF4joF1v17KnDXmvrGNSWoz/8dl773V16GrbciFNiY
SpKOXp1taXIcQWmeprKTa0CELAcbmsQ3q3J7MRr6S4qz7MrzKmgESHzW6OxbEPWq
rQYPttmptLuGfx774zLwCXDR2Ia3m1y1uiM15OSXxCHwPD7KA7hsLfL6sKnaZWFL
U2H/1MXLln8aQB/iNY0Gl5lv9fDaCPXIZaPfuOEheqTyRKvowLB+EYNWO9NvyFFc
5FQOiQLwfB89Ju/VbeUFqdIkXHc5mkhIudfU0I2tZVDEsy4R71GQzVPGVXmNuNgq
Rox2psE2SOOUPOdXg5dOa3WFjioGjbOmu/cZ1rkC4rYd4yyjqpTmpg1kMSK0Ix76
+6YvYkll08YdzONo81lnyWo2A16Qczv6NwHO+RYWMGwDeJ5dXSi92BFkGTn7ApUz
PJPe2/OtQrB0+uDcxtbt9CO34tK0sezi/NoAYXmBU5FU8vtCdVn+eIy1GUQ6m9cj
MmGOWoqSVbAeYD4D13M4AbhCKhuo641Ul0ToT4dNq3/3X4Ujz6DoUvOnBcsYDDtw
ijH5EC3HpMy29NZEB0XR4MTddKcr8qVcerWTWqnNf/2IIo6FPGtNdLXl+jVB43Uc
raRwZD62Ni6I37X/FSh03qpKdR4lC31NYdGCjnrUQJAnUW3xiWhpuAUlb7C8ZA93
YyAec0eMaY6ei0ordZ6r9H76yJMIkpudcX9Tu4ZemzelVoZ7Ioe/3Ln6iNKSQCAg
tUo3/UGK1U4lFR9REKT7EZWvmLaXg9k5vIatH6cN1WmGDtwWTjfZJ6GXQTnd2BDF
sFaTh9JsvTwmG6F0aN1DcM7l0qUJ+e/J/kKh3qrzAOXqvdMBU0nf7CcfbJx0XQFh
boYkqZck75MJK/hm8dFPkbinBGujDQlGDnl7UJUwjZoPUOO8djKCzOlY8xkzsaMl
OcE9A+eus262sLt3cF4+KqYYqvCTcWSdNmCyRRFYBnWIngIqcNN9nPTe20eoc4D7
5w1vJ6KxRlnkoBbIEuP/jAdfffCXyJ+PQbHkc4PZ5/q2PYmjKQMHZcsgBVREn+Go
/H9k2ATMNKsAurmuV5UqH5J1ZOjrYzbbIoIjt20y65sGySLlgE0seUnulUv6uoyA
teIH5n2hsthPBsuGIDhmwG9VAVGBwY1ySUmkJim+YUDzuhLyrwdLdhyVh+ON2UlP
2pq4vMFdbgUjBR5bXcI+HZk2arIj2rqOyF8/HGEB9c98G6hq1CTcgq+P31Y39H2y
44sP+laZhlZGhH+6Y/AxC9upDE8iPdpA3tTrYzMN5xkJKvIu4FqOggViWJRIpe/R
S976uBSFuiI8Td2yD66/b6og9D6mvKnsdWiT4Fpol2uNY6OwXZD7Xrp1C1v9Scg/
r0Q4xLiJiwxE85sQPiobGtOXim20oSQxT3WcHg4jOetE8WqOHfrC0twOQ/WNyEHH
sx6XYA/K7DbN8VCb/x3Kxajt7QIGm25gHE0pXp15RU0nrrr3Mjk2Tkjj/RfL/HxO
vERhz9rssNbTmG9CDXdZ4oQRUnEBc660R/TP7T85DMFvmq+Pd+Kk+9Ow4wGq6MtW
0oEYVkli+VvB4RuMFDu2KOkQ3L1lGVvwtSxraiKV/YBpr9p1pAqMzrv9qjGS6g3U
mDAGX+wZXaS7RfF4Hxo/SxubBhCZJD6O6LB8KfAxYPnfx5eiY1K/pM2W16mlIgRa
StDDCIcNOTx8EVGCD2dgJNga2y/tkN+yyjVzzqUgqnhVfbl7LZths6ROjWu7obNH
Y0rV+Gx9yvIfAQZD4g4u9RMtkNNVGrf8Yj0ZRNo2L6LAYwW2jou2Enjv2L771zD1
WIwMVY1XNlBEfugo08zOvw7RqDYngJM10vVeX8GK0y1RNvQBEW4PyzLGnJW6I5RI
/r2sFzIvTGG3Cku1qHEflA9tZtIlXq9gWmbSRoIMx8jEceNzs44n7IfF65kSLrEP
Rhb91CxrleurTSXSebbE6SALN6yab8Wy5uXzSwoVA3HDMk27wspp73TmmgVNCtcy
I6yffM/1aQRLdhy6bWW0k/5HaTiAJuZv4tVsfKhZ3sW+0OdlEXFPCSsFHEUztaSw
f7Xi1IOEzGhmwY5hy5qPOr8DJHKPmImLGJW/uY9Mqr9U1HFKmXEUIj/tPGN5tsAG
dBVqv2P4UmvJl83K3+xN0GBShc0iTaQLJlwbwftktYlt+ZSeShIHbIGQU2aFshnl
VM8K7ZuDSOjqQ3aB4JFbQLAfxO+1KZDYcoUeKaQ6H9fWbxm/hmRvmxkWawA8WokW
KEhXZYviPDlCrNZ933seWcW7fEGH3gKGDzqu9lG37kjKslkYYuWYOME6WU6dZdnb
oRuGi1YEOsQpiJwSZM5AAIphq0a67De/wwqPA91zXcPLf37SG7nqa+Y0IHxBH4ww
i5d4PBUiBy1Lga9urtW6zmid1dOZzuQVyXCR7YlRQrKJuvp8tKMr/O5gKtvZeCZj
jLzKp0422ptJO0tbEMaPhrYZkEpfIJB14WfI6bOHT+GaHiamTEKWjb2bSXlbyrtm
t+BUlTafYsiCZGI6srLJqvRUmaKSDe7JAgIgaAYy0CMNCbmn1c7WsQJx7s/FS4BC
f5c7zLoXxPfr/UhtrSpv/dsQXoUOxFi48TRL+7qtlsdVogXyhnAz4EA4QX/dh7OC
hhKDNupE892KocmzjyYefSao+NcqBlCsuq+/RH+urjVRDgN5vvsYwIXdYcu8w30f
5HhuHakIer8pNTA3PNoFD3cYfDo8Q0nwJD+g8f4vL4ygf0gWJ1soSeschm8XfXvA
f0XMbxJcKndb5VTqkX+10ejPnQ06ZiLvVJyfaXkGoI3xF6kIusBMIwD9/MX4l94C
K1mUUvqkQlHy2GU8hyDkyLo8xDrsW4HbBGAjWGlkTJ1jf1HHsrw6zck6isGB34B8
jFFPKDMiX+72rOJJ35j5h+zMMpiMV0yS141GqY4xaA7EsXr1o/i2wsBi/wgbaTgL
CF2EuSuG9IwSwPh8+oDfzVUTp/n7sHTiN8L+M/dgMzdYSc06w20ZWrJ1oyRTghXw
ij8vg5Gfa6wqeBFOfr8TUllYz6EnEovO9WAbjfw+LsOu/CWbXOZl0GBr1SHG+R/2
IAp5zHSBlLaTzukYW2VvNSeHdVoC0ZQIbdL5bVAbGOVsbcCWhumAB0vru50fXNG5
m0z8bZR66IDldoiXH/1NfTM8z0tNUW+NJA1UBco5pwwLaIDHqlU1cCTQwCk2DlJO
zqqU2scbU9YkD5T8qvzsSrHelNx2OwkeN4yEO2rXBsyozMbeDSXq39Q7g7P3DTlA
ai+DRPuaH1+d9AHOU3iQw+nbZ1m+c1//Es7wl54P8Y+t8SqSGq4w09xe/qXZMXV5
SjP3H2RnxcLC8gVeLJk8PY0nEMInUDqT7MMD1nOaFdFzFWIeNvyMAz3obPhaJN6q
sb45cpFDktyu6nMAbyDOOvcxNavM2ymjIvFTUWQhNmu2NxhlC7w6CoK7MNXYyg8/
xxvBbZGt9PdlhxIGHcCdjKroS4KsnpA1gD8xfdfooZ/oKsNtLCnHhvJtJke/4w2Y
U+doHFf1M1B3JnEfe+aAkQiU/0vsiZHRoJ0K39QXBhQ5hgfFI49weF5EeuPhqfcH
lUMNVCdN2e1KOsooLfY4sFdR3J07UUlGqsRxijkoqzc+tM9yJY565G78LHIa50GQ
BFizjU2zi42WlhKC5cCsQiW6VwGs+iLDspDKkP/UvivD5fAfhLZiW0rX4ATQ3DL2
ldi+F9i03CwsJNgGykHGR6zlcLkzAvf8E1hnEvDpzM+SEy4t6WqnVciShD5Iq/8A
6AWaxc+fuQ9z9jaSvuNDcoRzVJfKrhG3R5YT4JQCbtuUzMteYEKXN62YU2N7aWyw
K2eoOXNMmhxKa1qhvRMSQ+fO1N5/zmOS8Ejocv1F98lG9sHz4skvKEJdyxcO8xkR
u4r1YPWJrW9a+I+7ijzKm0ai4fA2w4O4zPkJy6p1Puh37V13BAXvjoIHsdPgoLFj
mVaswg8jup/Z4wigx0eAptKfATQJrSKy6KTeTet3RrugFD/9ijuBEw+cvtmw5iUq
LUON9MAED3dYvGmCQT1fvdClAjXah4TqHO0Oqkio06w4uCQTcMKIsaHL/fT0ivC9
Ydhz3ximM0QTozcg1faUFDkoaDn6dabYyyRSqym57aicy4awJWTWlzf4klFbfieS
YSEmfct72iyGeHPet+qvC1a1WBzuowirbV57Fzd0iXqw0bV2R0OkbOxGKNAsAD4I
g1GN56NEllZGLFlvbSXU4fyqmJBrmd8QWrJiBVBE99WNObZX4n4Km61ClxwFImWW
OOxDg4b/NFSiiOXKQHBmf8+MoLprK4gpPQcUa5Nl2AjGN1LY7/RprPXVsBM6LbXs
ieriqnVE352AoxC/ppamb0CKOckRvMPV1InrqfUm1YQRaCNFQLPKk9X5xQmNAtFa
D5/BWCiPQzfbX667EOzOCwKXH2pU5u4GAevwwbWzFMrDGb1Sa8nZlfuBQFhmQX44
8HUY4BIClTb5qb692ywk+/RBlPX8HerNUPUglXGNfQkz4zyIirYrQho/5pp6krmR
KF6zYW1a3P8Lbc45kIEZ0zNhBtHwsAFV6x5jFQGc0CNX/IBmArJxJr4a76HQl6kK
xC2lQD6B3EHSFYJQhfyLgdm8sgD3Bs8jLiODNjbDkGfvuYl0KwdDgsY1o62CPmyx
0kpjEPFk2WTBqoTMuhM8+sfDh8/cvF9Ve4XFJjWwaWKH5WET8e/p3t9Ce43iI90s
sm8uFUT+BVS0Fwl/Sb+56tMDNC9qh6wuqA2XWfzEnRmuPcpPzMqs8tFrZVSSNsuQ
MSUGgicDL9F2as3f3H3vWQMy9dCaOiYlRrl0abyOIkNKCumyko1UZ3xKhe3rOeN8
41VO/f0pBAhjd4Cn2+U3J93gnFesZsgeea/Sa0QTY1+8yWFqYrAdSymqWnC7zmbo
JaGX7pPwHquupHHc0MArbB70WDqfnvPLqjo3Y87rLEL9oxFZmywkjr5Tww/qj2pb
0RNn06+WhhUkKQhS+PY9KRwI020WaQItMC7z1Apy0dhgDrNqXNwBwRxrwTsWNUz4
guvFWVGoNIvLQmS/vEA/zBDnuHKrNA2L+v+w8WcY9tElpXbtdEw2GxwlObNftUBe
xL72gfx+XGWIW8bgES85206l59fz8QR+zrO/1udLbnttnanoDKW7gnsDHtPAkqoa
p21QIA5AEsYIV9KuT6lHn0INZEAiJLvuxDhFajhFjE3HF9zgRIJREcDyz1pz9P7j
IEFr0T+6fiO38xqoIjBs1lLYLzD/CcCD/UyQTPPIQYyRwAxTZMyGTT+Jd5zBFsUY
a4aVE+as8y2sbEwDEiFkQLHLyGvmqcDWwJuqFNLNwpPOStovCtkQZFoCpKCAM9/1
hk95T9xOPwP4s87mXE5KxpSRLL/2Njz4YzICEWZaG5PprSmYyGsvwxrIgv8ixgSC
bwIMC909xx6bHcSvfrordUcLi0zwyi3PFsYH79gGmjpAvexBvbR7gpc2diQ1otrK
EiOdrv0OWxdoLAtK47Ftc6xRQL1Av9p2e4v1rBLpBvPGQ2UAn0q8lcjR1ZoouenD
bh253o029X2bSV1rYHpPUM7f7i/3i8DKintwgU47ndw9hDB8bDJx5lOPGcxzheM5
HqsJvN+L4pw9Lz/5kPjzgg/iEFhYmlOCG6xb5NMIWLWC28opplLiEcESY4zqHGo/
JOK0Id9aRL+Tgn0NtUFQxqoKaH4y0w+DCykI4JrqgKYYk2Lz3M4HpFCIFSIoIbyX
AASg6bHV2PzcGjLbBFmt7lP3sbRZosh7l6S3xRdPzptKiBb7o31o2V9KCdZllxx/
46fziSssGBIlo4jRhWBycTeojfnOMR2W8nuhuObCnrcgBcoiwFhJ5AQR44awLdzn
4Ns9xJ7honMveiGZZFBWkcaiXlz2MAjqHjrGh2aTyusYF3rnyfmz8QHgABo6icIt
FAOU/T32TJdNFa8D71el+zQsj1BkSE0PXnD01CbxuFFvDhjNPm23fzwTyA6MPdk6
+yW0L1ARFoT5IbdsyUxTsTSAm+f0deX+QJUfTi4wpU8FvMBRw/c2Js07geQoPyvb
DS9uWSkS+OTn0rKZ1+rou/98aotCJ7abS+99uPnNvNvyGGYuFKZy9GUdw7KAOly/
/NTow31z18l15EhwoxUBocGnFQnKC4z6mVPyrDxZUhszI2GvWzezToG1N8V610zj
3U/atYevYauXD9nqtfLekNajhgfkCmZ6FPYD5X6S0W/ZDfiNwRf5v8ClDoPpe4uu
jJaCfFv7UtfZX2M/so1zS07Ih7DwzHpHSnbF4fJRdTmJbkmDxVPHNdSJtaJgLICi
Y+DbYfZ2rr1Jzc9gSAH4wFpz+0ImG4VOSFP4L3HZOMSoxPQuX+xX0wIihO/nlTJZ
XwKkpTcDLbahxXEKWUlgfKt79TLNOh25BddBPfKnZLcR/eLvrqGk5U45mrZE1N3c
i+6UisrLrPl0MysUE62t+CiJu9LhH10b9Vm9o6ara76v5wI2qnYTzWcmDC9GSZL1
VPrxsK1fqrL1MocD7zTqurgSe/9wyBcxPu8maz8m/H0bD6GwS7DE+phjlfgFI9QH
DyWQ6Amh+544xzF0VPNnO1o+xuiKHQ46X5K5t3UqoNLdGQT0cR15aikJ8xdVZLWn
pG1z3GdC2oSFdgsl5w8Am4B2uROTCc+fYpafsGfN4tWwXL97jh7R5qev5955E3E1
J85Zscm8oXACl3jHqrhFrD31PvPb6obzv72pDs54dRqkKyDwGd2QKD5SG6mLVf96
xVZxtuLVwKX0ZOMhNicBq1+9KWQUW+Xu8ASgBpGopy3PEoqrni0LIDXi0Vw7zkx3
tWprstVzxl+U2Tro9+GEddroJ3L0qH9cQpweHq+ciqA7ZRvsP9NTbB8Qlwh8sfsv
q53qHPtLt0eIntRTHfbpoXZYO0ZkMBDUK7PCl8rdFz/wvv5cdgkeYe9M81qWfImj
aSv4Mq8Ad+kYfNSV1vMbS5+2fhikuw+rPjs2bpNHuUoIIwrCY1fw67MzufDF+qKS
FoC0B+QVuMzyMg5qTv7YxO9sBDjRCLbt4P/GYHye0q1gvwB26RPuTigPEWFOdxgJ
NUm2e2C+t6guH4AYfEyCG9YSTu21WYpweIjd8tetk4lVD7K1Wq3CxlAmZrVnEE0k
JJulFcY4OQaQKs+WQa7/JjUY8zBvnnU6a66lgbfwvYT7TeNAVr824UUf+tvp1gyg
8wAOmUh1IRusM/YGqdiLd1kRjNchdsgdz/xoSGa5sW+kZxuC2MqrkYhXbkofO4Mr
HBXVT+Gw9WnLY+LgQ/oG/2n81a4WMtrFx79nX0Xow2XjXvuOdvQnYfWDsM7BAQGq
w8BKfNXTi6fOjrfDgp8/WfqiyqyZqKrc0VENvaBXzIOgz0slPCyxBZCyHNxMpU6r
1HgPg3t+NRhwLd92OPkLEybYq7P/MOvo39LHYnNxkX2YKEKyVMYZu7Iao6GNKxrO
Y3Mk5MYntBYbfA+bhZkMAnUsNp8v9fXsndz4z180nmtZyP52s/MObXdWRd1vkSpz
xOlNwXA4tpythVe895nRttoiKV6uEJGWaXvVS8UoBa845+xVaKsTqSbwMW1S5cUc
WfibBIEWBmRPdmG4VN04F/RfuQM2vTUfKpNNUw5WqraFjnRj5hfVo37wEZkT156C
8748thMBBqGZovAR8owBZ6ubmu2/yPblEgpunpJFOD/Xlc9QDiCgzaY3mUeCA9gU
tZbaqL60/ahe7fEs4biBxpqk+BeR5OUlhQYSArDrMrdqXQssLRn5nF2WZ6ZYXZ1n
BA5T2UgUq4EPpeVTscfnsKtNWQXiCX7ywYZGlaa6igdMEFSIr+Rt36bv06CpGwaq
1UqFZGnEDw/xx9RyV9wy1pxOgwspmzawyjku5FcBeR7No5jdrVKrprM6Wk/JQ1Pt
rhLRQbauN8wdydc4bOMDcDizzFA3Am2gqR3TCW5PK+h7NezgY+Mt7NijLoXeuz6E
PoojjQqlGVyypq/iv4xsH641rwu/W7TUj9HzbzLrGqrJOsMeHMbaCD9ebR7hlRXd
BkoJFA5pP5+0xDix3IkLFKPDWY1V1AODzy34ZPv88tW8HmzonPemf+JV7eSFGoyZ
blXGNlEiH5Vj9W5fvxqQwPcqPHRcV0IBs0JOCBLZwNO5jR+NhymnSqNA9iSrsIMt
+GMRvf7HIAA4H75vEub0od/bvgwmyTTYfDdpfkd82H2xU2v9G5vK/XkLQRVpMOSo
+11rc+uRkvyv/RYFtBdZAzkifulfn62mrrFhKuMZql1cn8ti29XSlTlhAutjKhLJ
ZUrbNJRc+QTVbbRxxJdL0X+23hzFh668+NlN8X4b58PiAVvJWVlZ1IrVgbg2mPzO
Fm7DQGkSM6r7yK6DWy4JZMzWO7SOPH6sWx6TsSsQ82rBg3W0/JvV4iKMf0rxAwGy
UUQ4Knu2YWv5ASzTrasTl8zyZkd8lE4CvTAK9z2twsfpGWpAsenhfiQHmUdPeLQF
7xECPRW9ndjBpxEOf1rgtNp28jw7MSPFoAPUr7RNdFoJYfkVZOpc/MzRf/QWPiyo
RZrJXOp3j+lzrUPgLDumYzAfEaOManYUYzkvX0zWqZw/ujtpM1QwOS5XT60z4rmh
FyE67eVuw6AdWI90lEDo6utxS5QNJIbePtD+McWZomFkMhIkJaSaiCWEKxdmIBr6
pNJeuEEn/ERMdRhbv7Llgsz42I8zwFTsw3gzhQ0TlkW4UvNv1iclgQApGdvED3IC
H7f8ueqftbUmloXTEPTyLARIFtkdZyzUtHCo17mM/Ei2b6FvMecx4Kb4GaG9uuC6
T+yCUSxp2ijOdpCM2ao88Q4me0v+wCc2GOCkQ1kjtUQ9o9RdxQxVp2ZiJdKHf//I
fgCzEy5whhivdL4Cz/9/q8qeKuJDLxNPnRGVXQhZrlm+cS8BhruXXa2WidJ0Kc/h
X2Sh/KN4d0/WLlmcM8l5DC3RNVzl7h06MTn9NtQlf3bwL5pVxlK97sWPlWRvoCwa
XWgxFjTf02BZuYNQF8fjeR/y54Kfd4Pd6sl4aae6bM5kWCCLqxuB2843vGWHEFu4
ehs4aStTpPBLz+NC6W2gPP8K91u7hEBnePme64MspcQbiYFixgdc63wurZ6RQbS9
Z9kxeggSw1oXcyNxqpq+1nObA8pvFSqYfUaY3aT2yG7JXx6hgksAHBNZIJo5PwLM
Wd8AyzcUIrGp8wsN/tUvuByYDZ+lKtbRQFwuQNAKZuWEphHIG6yjGjXZcyiNQv9V
DeOm7lfk6ylS9QXoDU4dxf2687ABZFbQ3cYKmWLQonxBWFpamfl5iUxFzKcsjIC3
ERsEEFraJobjzHJjNkRxlKVVwS8ARixo8yWCZ+O0C2QYg3Ijvq49UszJ1pzz+EVG
Kylj0QYMw+esogIlnME2JQi2s18sesUPkHAcZ+l1h4+PE3w01YIkM0pzUPwyyFPF
SDs23IcCNagItZDi+ZFJTmSzx/XDNqY8lEYnG4nhg+VDoIUwi+3EZCOgybM6bIVN
+UzQkbjGGVFssRA+oblbldm5kOro87uHdDJkfQgiD1D07+IncZ3ydF1XzavFUclk
/7/7wPWXlo8y2EtKCJNc227CSunYhuRW8lnJ1CVkEi88EYUNF9avEN4FwGpMOQ1j
Hq2E3LEcZEoO361QLRKY/CY17ifsZCrLd1Sz2PA5LgI7oGfDVNpSaicS+n1ZqgUI
Nf+o74+R9fNwCJF3tFK06sSIocwmY9w1ZDQQrry3xU1qXqm19T98RWdLbtQkpwKB
DSFZ2mlTMhpa85koVW88lppNKgHNGkTCgpyVAUVgmUWHYVZGROPMG+HguPuN64me
UYGb2LExxmsZ9Ta8t1vYXPCRgzaGXBbPMfchtNx58FB5qQ/8ALg1jZEG4aclIRn2
qIN833R8rTfN8hXEitgGZa0YVD2kXN5ccHPVIyDqanlAceDHCcyzvsNxjRXcPnTq
RIou6jxifEXPWaf8P1EgGB0SbK1qimexzcVY56JkE8auf2JRXI62pNTvIVJiSUWg
qt/n+5teHshFosL8Mst96wIFXEDTeuDzU0Zo1TtsUvMGdu18hoRtaShr5Ue1+8HD
x5icpbzt3JicxI96YIYB6FbwXTU4DMEK0FMMEMOVITOBmvSuu0HTfWs7auHtoTri
w8v1bUkqKbBZ1ewIoQ1SZLkR3s37c2CzTPRcEAF4GCG+tExxvx4dfXvYk9cZOGN3
32qTsX6Fn1OjRYnrCBJg+odyVGYh9D329nbjJ5jWFl5FFqz+vGUOVhV+02T8qdHg
iWU1ziHMzBvl1RbzRqdBhkkmGigTfFcwQ7FpokM+0U0kzesuw69j84AaK2/LUzo3
JMm1cPG1wGerRTx8ijnLq2QOiZ+tYcHRndFl2kIQMfvyhp4vR2m/Ynv2lKDHbQ1k
NgBaf7q9e7o3MdEjTRVJRCwAMPv5gKqEWDKo2EMMhtshn/yg9H4dceQCH5dLAhSc
qpQ6wJHLZ0khy5l7cT99r3unLdIRkfTLTNw5If18vEVLS0esvKrhWwcrNWXMaLfh
R2PhJWQspoXI9di1PDS1u8wVg/8APn/jmstHuCj39Y8TpMAZRYCRNsOHGXT7rHU+
iQ5LACBwIA0BMhFuy4ScbLVvFM/6T3YsKmzwDPYoPU2hFpPOSQ0QxlRN+d+e7CA0
3feMg0Vc0qSFXG9OabPgSLeGhqsH/Q9iRab+KMhXfI3nGAS1bJgkT8EvZtzl/rn+
CjiacfOgmzli58ykAza7+b21AXsgXOt2mY+9BjfrAC2xTE8pac42ZL0Sa3ng5/iq
l0gp8JUBRNDoh4uiB+eg4SHQIW7z5k4Sk0XowuoutwW2T+jRo7ewt2tig5pXkaRY
B+OAZ43EAzTXTbQAfFdBBtgg9zn+zp+yzWnMiuZP7wU32N7lcjRIbBRes0gAiBXt
w0UQUUyRbKnblNyv6Wawm/8MeEJpKUMj2uZvpUiNxW/uFSUQ9/6Ga0Z0T5/G5z8g
V/Sj9cp9NHxgHrx3sdW8vOSdtnjE3HVWZnhdexmTjk8xTIfLzsGQiKJ1M37SrzrC
5uFi3LpqHS8SKrz/c9gIkSW0q67Uo8q4z2aLZXhJrl7/9qr9cKORX8fZ1sBTWADK
Xi3/947MhrF19JcQFGhKkyAOB4/YeIcr5Cv+vOzVwTUg3K1gEjDm3Uksnw3U+yRL
LdGa6su908QdbqsELOA/WSKRx+DvLPrEcLnKyQOb5ZKy9sJxkpC8Gj8kCK04JkQG
oxBn6X4yPOScWegR2sEZzeR6j+L+rNTcz8I0BPgXhNZQTJ7pXDXFo1664r/pNYlv
iDbLLzVUnD2Q9LTsjk+bJ2UTbR5p6qan4VCvCQijB9V2mzWZoh0VI6VDI3is8PZC
HAp+1i2WRqsUXi5FuiUm0VAdXLLCo6klfNU4ONVpZRKvlOZFMmqMj0kJq15g1vM0
jJNwdKud5SpwObpZo0lV0JwBL3/fxlnjOlgzlBLoIY8sOpobUzrUFYSpCSwTxA49
tNnT0fP+D8XaWNIs0eHmnyHIMyBpVd/kqPk6hKjQDo4GvVAX9Qf7HCDhp1mtqYEk
WlEoULxMmOz3tEBGlf7kw19hrJHgKnzeuL8H6yHGpr7mz3NshHMnW6tlndMuysw3
KZskIwU8qnuloG9Fazjoi4OTMEOKNG8M8ijDNuzP9Q7MXkI8PxpQD8U3+w419AyW
qZYcJdIfBqolZFD2gS1rVyCYju3qDUq5u4ZVOIM39o549440Pjn/jtzd0AhEXVD0
ntmXN5aM7MLWCEumGoRILwm9bDwaPyjc1YlUeEg+SY3FLM/NI0gJvh8X4tQL1kBy
Hpy8OUvNXKkYmiXU1+tnSnLGqwFBXGOZcfQe8MtA4VK0zD1UOR8C1EDdMt2ywP5G
/bYfTGnmFziCGz8+klqTh7tPd5n5NCNIXpNQ7SAaQ8yu6L7/xF4W2bfDfH6YG8Q4
jLHAHiZ/kNoqR5GUvVgMfcfeClJccIagO8/7Ao4mIjM4mXLe1hT/j6NNoPGjE86R
fxrPIzT/+lUjPAQ2iOt8427lo334Bzvqlp+B6G2Vc1fg/gDzuDDQcqIRKho3Nhbd
rl7i4TzD+Hux79NOV+d4d9uOh0CwbsGp+kXb7uli0ZXOcRm8xErTvU4PSDk9uVho
PLIermSDSY5RYJBvnetEAPME+1+Vl263Lva1G2CDvwLFkggLPiotp8UlaBANfjMb
SWXHkiRRr9YPax0Vji2RI37n8FG5cH/BARcsmtcbKYq5ZDlYpFl4ZpkcR0xhVUn0
WjiqvtgD4Htn9+6JdbbM+akjRve13QN98rHcwEzArg5BYezn27RtNeJIxvtxWe7T
uXs2IyVTz9wtLjyjVwccLVFDtHdhgNnJTl43r5lu/CTd9YJY8KCsvvph/k+vye2I
bVk5CJ8j38TldBUO3iFbGJnROv6LWycsTwuRe56+w+/VmJ17sRsDdJhPvwl1uZuh
7J/Zmb5ufoD8VPWsD4YXvXZ3lehheSAaWBSfnOn9yUnKZQVapZOsl3xTGzMSm12Q
SznutimEfDtmANwau1e4bsJhWgYVfH1r7fdigEHp5jOvpCD8Q78R3P6OmgMeCW0y
JaK5VhyCpaXTvMCV+vlUUejWoopqhEDZ2f7IpcSs15MDce1m4cfqjNXVh98LLMws
aKjpivdYsrmKCFMuEKshC8dr5LeMo6ALNidyfTJKjhM+A3jhzC2zbTIvImaI2wzl
Y6uHb2Bb/WpSiaogP81KHSsSu8fwSoD6FglTypQqvC25sVzR68GorhYS/bOYUV1x
/ZJVwbo5lBqzMZOY2hA+E2Hk339fO+xUw6YIrj45MJq8bSivYUsaEhm9Fl7GG/aL
966Lr8lTY2ClwFzAZp5Cu4RbTszapc8gD1qYa3d0yDeqjsCtA/obEcYGzIXKfmt3
/n4NvVZ4AoSezfFkLtftSlyIuxNyC8ZYCUubu7vkJUhfmZ2G0wmCSkJfwaGd4ZRJ
MmM3P+OnKuokh2IJqFBXJbzOgbEe7lgerwf/IR1TT736N2EHdSlFtTLRjN2LeWRl
pIfWlLMLCBVTj0EZ4UeiWysGAJPWasaGumkkTB5TKgyLk/hrKyIFzwNewoEzcpcc
ziSaPV58HuoVndGX0A6hZk6wmhbNw3mOGp13iCt14LyKbi0D72ejy6CWtFevZme5
ydoSsZinmkwuOB0TMXKdmXr0NLO65vQUlO5zUVDALa366wKkuaYCBNI1hvLHHmG6
7gQjIlEyhURl8ax9SntxppUyprbx9gFCc9FH2gcHQdAhrKrKLbBhuNwQOEEHLX0M
dYa8b6JlIb9sedKeOuviJoJRb2PuWmS2BXRwZmDgxkL49cJkhgLZwrNyUseLgyyK
pBf7FRtAKyyPrZ1+xPgefUU3ZgzxySLocdxgZ7yhylwJWq4PamMoMikGVIYzK8Sg
NGrYmfs8hiekvVJtpHdbx0zAf4f0Pv72loroUtUo7huAoyGDlMu9O8CcPplIg80F
m+tP/2iMcF7sOsXK7U0tXV47myZvCmkegEFwCqMNzlea7cb4F/HpwjApSVEu7HQm
IfYWo8tBudm6fjnA/4CSxV3LzuWPzzkQnU/WCv5g05qSLxXR0K+oHPHoBl40lAmc
4592NxvxvGElJMMEC49iY/iGPsEpK49rxUtcXAPuD6AdoMr8PZ0UlU0kaQ8U3Gji
pmRhoVS3e3+Li8Feh4EmFuHKx7zvW7b+IHE4KIXXRYC7vynQQV1Kgje72EEOJvPJ
LkzZcHqV2cNiO/vPweQnPFGL8DDWwXVU6tPuFE7VFBYMv09w21JxuEK0BioVoGlD
UYGIg9gKVksO6zGuFHsXaY/5baNmdvEEfwmPpaQYRxDBTHT/5zjOCKSUcg+k2yXO
eBGjqvzghUstOMK/PtURpYQ1lioCZJynpWBZb4uBLOd4QKitIRS5K6ue76QxDin+
546r+C1fqwPX2T/ZVIelyC42Ifks+4vKMYj7zdOfE5YIG3lzygp5n9QBw7fXYEco
MQpEeaMR//v1HMnLqXvKOHAR5rp88kywWAKjDyV0Pc22Vfq960ph/h962n46uTY1
LFmYf14uTC/aiLhWcFmnA6mWI7udcjhs445l4ZnumwhjyZQSFOHp0HrMyFn07QD5
eKbOVEDBdER8HVxCS0IBJ86sEQmPtpUs2JcIAFFu10taUEoTTVOwL5bM+0vIFjYW
1mE/ITFcdXsShEQrUt2YKwwRFK9szZd0nCylgxJJLvnmoXZwl+aCoPFcd7ZYEAps
/BEsff0M1WOUvSdqOJkPetmiU8PbZooZZzIy2HuAMf34J2bOUPhxNHOG0cH/JZPO
+FPmPx+QyvoBt7KYw4kVAQqInq65sqIchqhYDsBHtZWxvtmJZOVkW2V2ez6ZAMMI
8U77vQ4N5cNrherQgf4KGp9zr5KdsZvyodGu5WvSplmvFuAjzh6Bmw+BwvtGZE7o
BWAUex/8uo3Pps4EJKwjp/ycPjLWoQntHBPLC297TLkrp/ET8rxepY8g3jStqT2m
Og8Zh/kWLNbHViBEw1TSH9Y7etd/PthWMygb7Y2WZorY2EDDs3Ybbm7xG7MOKH3H
djy/kCjL+sfDdGYQYbh8O6IYFgxXztf1wUfaBIU2/WbRlPBHoSnBYPjuwavRZPif
i7bt0oRUnshzPjQkyh0tEb82ONruSP9kkkZ9Gee1ugblLqsZ5EowxNHNghf53opn
43AgvcUOUr6Wal0TZBrMxxOU2/8+58KcVAjwIvGsmCi6eYk2QKjfRUVlDKMLgUn9
7Y/QFrHom6U/C9WE5N7CNeZQH6K5i2wE30zC1BFb5CSuhoTJKqng2A0jSifM+wt7
en/MMcWVS7JdS6Bl5gduOdkdBk9HVz9HiXJuyzxMBaCl5SSXJcoqTckYaCW/Ranf
sfN+tJ37QkmV+b+ESv3btqkwmv99idUnOk83eqiKF9isEuSGTn2WA8BrmhmOUjJB
aIHfsvYGq3WUkOhYEqccf9zgfXl1qMzTdu8/uTkgvOwtz0GL9KtLfLV4H5lqWWsx
oeVNykwvjPJYdPs5W9Ejlelxngmpjy3ejQn3Wf8QW8ediOAplLxmcq7JwBHy79p9
SW0WTUkMN6re+z64RTgcmjfoUrOFg22UG9IPo4Kv6mrONtEfm4fMmKwkW8RaQwnr
Zx+Jlv3iZ924hLQMyTzHZ8uNoBKqnZBTs0NuY2moOl+m7InJ2ocpXdKV8w9JfNMA
hAtWlnFum/QQZwtsU185H/bCCMa41vm7OA6YyYbGqKYVK+KpuCVa+KNJcMmpu2FA
ACc8ARt9bqKZ78WxLgP40zGEL7f9dqmxTpryKAgwR9DjNVmKKs5DYjV7Rn725qH3
k+7kwRjahEHiyQnTtHfZnc3LsqKy41s9Mb0q1sfBMjvSGxhVPVnfYaQ1zW5J8SaQ
b3Fku16PeskNvHQrhn7rUnCGITgrkwGtVSRmM3TSEaTaAzfk/bXHRPdI1DL5/gE9
JQB5GONh+S7BYZiulndNn/TPpRYIjRJZHTpQA4xYiRd92nD6JipxSHluFiWzbTkG
2uDSx/1XemE3B7IG2qJ1V1/UKfkxbMzouSvULCteTgkdoqd0/5XMi32kQqsUxoUR
trmzD8DmxpF4zHcAjJw8xbMppXxnyB/uqg6jV3k4XdKkJL7h05hendYNediXKzwI
Ifp9kkdGtVGhxCnUuWvdKX7oCVO64WR0zIaZ0pzqx9RWS2Q/xeDv3y26YQc44VLe
2gauU4KFvs1ctd3JSVMLtv5K8Ecl6oWjxmjOW3TbogQtjGqb1dGliz6t5uYaPqsc
rgERl164yxdWOfh3VEDcqQROq2TR2YaTZjLpI48aFvCZBDy+s3yFDo0x4uAOe7M9
uMOIlZYeQIIlcwFniFyHTZvfbMd7596cTpHLlSMlG/+6EE7DhRaR/ggEk6Z4VHu4
FzEUgkvpZjCHw/0cc31mmHjSRMiTj8+T30WwAse/LeVzwr0Hsz9DGvxTH0oP1cd/
SUhBkXAjBAH42kf7qthqEa8bAc2RqbFelEZmpbqIFTyLEfSqdYUEBZEf1YxGH5Wi
rHcEdfiP0oHPD34W7a0nBsF+gHbWcMwaP4J0uioc2PsPL8TbxpNzedFHKu/v66LI
lSU/DrDcSiqkLR6EvmmR4BrsvcPfLAVR2zSKIl4ywGIJyL8ISEVIF4U8/IV73Uis
6rZRtaq7II3nCZHaq5tdZyGGzZpyfzaJ+ArQh9PXs7eM12NCvkOO6eTCzk0AOEcQ
VvG7qZrPO5U1SLHp1NNmriEGHraDaPh2Ql67Ur0S5rLbZ2ku+ggTXUAJrRBz1WiG
WyhZQu/fo5nCibW9A2s8mtC9K7jue7vzuAGMnBsRJz7Y55ygEJ42L5Inci2CDQOC
nwpJHPKIyDJaWsGOoZD4OdfrheJ7Gyvf/1yc+nr+EtTdpTZiclYU+9oUsRbc2TjX
guX52kgOEzFpcxU4+RD5MHK3tYUELOx7gc078MoGLQcME71JZVshTR88zroeSwsA
zs/Vg8zkdk/5Cdm7l52uQmXwaP6wudRFRUP9dy8i5jcBrghRSibep1/fizxRTmiF
7GIpi6Id85E0G0zgAgNHfGB0nac+5knpz0aH53xtn2kjE8EtqH3kaLxq7BnGXYSJ
6WBzJosTCGdxAPJj/V661Ot2G3hzWQskBU4MAus52wMUR/J6PRhsRIpcMJe86Gtp
zUOkuZ9i9wWhxzEklOpsUZC3VNRlqVGhzl8AMAcLSRPZCtchFcYprLsrEJ8HNXI/
Rb4C2+szlHP/1WsC3swMSviyapr+SA4t5eTl5GVT5QIV3Qgcb9rG6WFMLqg5HsKg
k1HowafvpgIY6iaQd0FHFbo4SCl0+rdPx6+w/f6tvQEg4x9CiChwDisOfv0y0cOF
JMW+MgPo5G0LpqmfvQN9O85KfYkIKMNBBV744Q0FHzMr5Az1I64BuHV74W1Rfe57
uVGyWLPLIjaQ/507Di68CWr7bnYn8mYxO1zYw2HlF3nv17jgxGQjghymcIdiOhto
C+KTFR1yFi/MPn3xjBuGWrYIb0PPQ7nI1fJxUOnY7Y/IxjNaCDga5qgs1XQ8QfXo
KWFlwqaQe4sOasqV2Q8Ve1rMnNubWHhIdda9JTodDxuKtJ9+3XzWlgc+xWr6BmJv
CVxWCBYHOdtQ67OVUvTmuAHaCMXCtnK6M1U5JSJKHs/79csRhV0etrtgvfpB4M6g
u6apKj13TLMhQnkc58SDog8xRhLBwrFKpampshtaJUd1eWL1/rZAQe11HP+T7MhZ
Gymtz4yIKigJLnMbHbP30Rwcp5m9WohPagPaANy/Rj1fYNzLX3Y1omyt/EqXRM+9
dPKO8IJUh0kqDD5Y9+mZsZZalV0VH5EPSnq773gwYPbbPanF+STghZyOt1JbmS9m
13y5/T0QE4iIPMlJzQ1R8Go156MpidQHbCwVsoO4T3O/e7ttXDN2UiDUpyfd5vmZ
E6JoOSedCY9pnCOJPqGrog85+rS0i4C6SoUQzo+z12XNkB/ftDqPpWfZXT6GEFh9
vZ7Dq4HSULVV90mckpf6oTpA0p7dwBN0cKHnekdkHDjrtWICrNHn5tGSlDo1vhHq
fEH5U3k7LCj4rxi5DusGtzJO0M0RttFUFPa+8fSiAMWiAjGIe6wbERGQUlpgIRAc
qx18sHVjQH5agRP4jI1UvyhoSv+6r+ZUJvTsA9Ck2QOj9SaSCav2VQMfLU7jD+zX
rUtpXoqmzc8/tM8v2pXEn+HO9Krayr40HkGxeRhZQxUmk/YlH1SHbNaEH5evrhW3
lBuh0dcl+IM5P9jNbR1NwPGOb/Es9R6kZvkCTMOGo0EruylTBOmXGaK8lTYzpcxX
fFivzjvlzL+Ae8jXua2PNjnvTYQcX2L7V0yY8fIiup1uUWqmKW9JMg2mRbwK08mN
Kcj4mba9/MGBl/Kkw5pJEcwDjA+gRShWQuSTaAW4sbMPxc5D1RoS4ALQ1iyJtCFG
vtkRGcyXivXkwW1+J4VKgc0w2O7MHho5BcDa76SinIK/Thw1bGZrfqQWk08jhCH/
GJun2h8HgzJViSnHHzJl6V8nyLB+Cm6gCAfw2w+TSAwk+IBZ3OKr6FDr3esJBZxO
9ooaqmWbQj8Q4CVPgWd+pATXPFKmo+5BnBv/NknFtqK+xyUvkHFZETOyHDZ5FXMz
lNi5twocLFFdvPFKBbfiKFX4kXEtqv6axS5J0asfmnqaItHJ9vNi7tP+OHoSRFz9
1K/CJk+vnTWBQtPwNsFRJrObhmuIWP75O3cz39lFSCuZa3qro2OJXD8K7kdaQ/9I
N9l8aKRPsgThR1TZ8M280VxYDylPMCj4dfUedGokP95cHY3gAoMpF8BVBf2Zhdfc
7B4kIaxm+JyjnxzjL50WyydNDc2dgs11mxQrcdW/GwXh9gmNfx/1psv1rTZbJbYN
EJ0LdE2B7mRyP448v+tmj9Z42ieZdcysJUV3nVHYhxMsEYQWvBtwdkpDaoFdOIRk
rNE1M0oomru+1O2oYa0ny+H+1OxTbxVS+TPYokMau1UhcuOwVxZvNVtkW9RCzSMz
C9FUzo9hq6brAkrBcvZgO/ci7aUZxln3MQdAEg49C+xRdXLwUDyAG6I4qDwGGjvf
gGvqKm2H9tHD6tRv+v1b6/5wom/LtUzXtGhLB0yCx+vO+WMO2pn4hqWy/79W+yAW
hbQYbJdfX69MI0hX8jO3Kvth9mOyZ8v3oKw0wHjmnJXndPt2zyEkfavtzW+bzLmA
0NGHesi6dFO4tdayl19BL5ulwiqxis5nZ3+irz/JKuvkf/6wp61FvV3ysx1z+eCz
6NgQz50USYjbIw/UpaLwiNfQ8Y6lTWP4jTnwfHAtsLH3S+FB8zytsf7wNBII+Rbh
X8YpynGb7Mf1RIUd1wGScFTDGt/xbUWotOx2g1kxFXFNQPztIsnZAf/64/Eg4LEs
UmF+HEYlgVbnvFAmlBjUxvzJyNuCoE+WFV8HhZkFBn2+knpbJKfZDLWJV3k8GDyq
2iaTLxLYiXHP1snfWzNY0zPIv09ojPfEx5CrEOk9hnWec/ljvTjWhYZMiAEXsP70
paR0b2++uqnoAmNcBzZOGfEWMV2LYtcxOHNpmat6bP9yVuB2OvNcoBYBP0tDrYwX
KF6y8Dig9u8BKykFtXb/SIHklDUAtPuKk1qzUqKarH4VSS1hOfGXy5rzhFCD8J2e
+0wtREAd88UFhe8/dUTCgmh0onnY/XT7ia67HRb/6g7zCybifW5kHasDOxLfsc+N
onwzc/JsQ6W/4k4NOd4SB6LbV0RzforwWQMEI43gzjPlbC/9x35xb13dCXxpkG1o
12LnyQaVMSDoBVMJX+xV3CLz1kw2e16YB8Er6o4/6SE75ZbJ1unM4NdD1MSVcRqm
PA1n//9zNDQCVerM7pwAZ7m1yE4+/MK2hB0A1cjcAniysUTKKqNNxMLq98jbmxQz
UnJIvByK3uqYPWYGTHTwrImVIWrVnEktbV4ViSaXlmWrij2J9SojxiZC7hkdM4ax
02zVaB4OJC3T9nGpgKMR527HlOImIXScajeXc8bwi29dpSZefZVFls6eKTN0vgx6
ofmd4e6KgszyQ1OYqJZ2LLAzZ1Vf55sOR5QQChhlzbRcJ1OnoL8LR38MoQ9iWx6/
XyjktaDDWoXW0CwGQ3vxZ6nSv7YgKLfOvnbOCrnpz/kFZdTLCOYCfSaLg2BwLddd
ROLN0ASlkQoeP1dZFWtIkMEv0DC81A4AM+yWoq5Bb1OqVWrAGJpf+T8PJBvLYImZ
u4sEa7dhhRsUmG9sGFIdOntyq/BaOaC5dgDtPTWFbInzJekyRin75w/Y1EE7nF3y
Kta5ytqxZ9RJgn1nJDZQtRljtfviBYbfyDpf38PW+/fYzwOWc+PLNvnutd1byCyK
wKVbIQ17KTvW2sXm64qbCadRWjD2zfjArY5y7xiWYf2G5B/RQfC+vHIFUEr+qnuk
faqtfyn5tmfo39dhrFGPh+qtF7meDFRZYKPQgfH4u1Ylculo32/FF3KZEIKx3bNe
Ja37ZvhmePt3XYPpWO6iYJHKZHwuJRfHm+dz4Oq6iSK8R8Dd/iV4j5AZETDlBHEp
ZQqUx6b+9M66qTujQ7P6RU/lwjC3GkZ3+LjvbNAnX1p0/30C+++2uyNcpY2FLe3r
JM7kbpu0rQXAhSBzODiZAXYsoqusZKcmQwV4gqM0K9lIAjWNpje62rryaPJ8o57t
g/90IH2zZEN4tZSPIteKfteUZ9Nyh0JBWOQ4yx9JALLJxteVWSC0coyguNSf+/so
c9wAWy1i34BW/Rpgk51jBzR3Ic6eZ2qVew9j7HEvV3wwl0rYzTTOsM5IEByV0ht+
Qv+nnpRUpjWiylFSROyzxdMTTzRyMOuO3uB9CZZhEjhgaYiz2lCcev6tSo3lm9Cy
0VW4afbDUokSJe/eFNRR3+2+QeRndK+DNZBLATkyFZlaSBy+jwJ8atTZxZgo6C/f
OJeJlTFIvqUhBvg2RIjtc8FIKtk2s0V2bHo+hEPUAXklIFeWxATdbUz7THfTmdx4
wl81pZOcJO54Lc7DOMuQmwh6ZkEcAwFJOOM08by8HcQweg30WMrdPfg4R3vUlrVP
KtxaAfj+E2c2o86L2OhBdjS9a7HGsjJeDOofZnYxOTTuwSKYM0XDejNNv17IoRfE
J+qkQRWUebU5qSosAmUNqsjuIJDyWxywG8i6lyIHmks8QuKsA/OI0rl/oT2Ls26f
h55+xQ6Qn46b1uD9zpXyyGx/4gwBhpTrXqcgVaF62IK3y1CowekN8TIj8DnzxQHa
LsnX9xbGAiGQeVUGkVtgwoR5+CCClenpCRK8+8vIT+ahlWxBVIKLt4htJOehHQI+
Vp2aVOiWwgs/ZDeNbOtDdEui2wZKdyRMW+vT1twA8SR/2p7+b8urA3w3EVM/X00c
bvkyNey036cCakeXuVPCRsa9ckZBjDf1a3sQ4qLuJ7R6vXEZ5wyi8ctK7NylnJqg
ABm1aqdqqBTYez5bAA8TVj4d6aq7syrvf+uN5goBb3nE4I1cpXTmTtHtwJngsMjv
hQNkcdru9gig+GCUFtkdIuDhoNfIF7UPW6qyniV8E6DpRg8/61A2o5Wbk5mnK0xK
xhdc3Bx7Y08L87ffkUAgEhSJpjmCZx1OQZ/l7uP1pOAQPk0cDADEDwINW/PIWmWO
CCjobIa7Dap2qGvBwFcvNfHuE6AMGpdlYq9R+LGGXoSVIiqz6Yl6TDfyz9bcwwN9
uAHit/YN3HW6NlFXMbeWNbkhNZKAGACkguhwrg6/ArMeliSdVDBcFUUZdINRSkA+
uGVmZaCB47KpVgxhkVHzo34N+HpGssWdU8cChDDrMlgyWuxciYPH/YUKTJAGrJgR
nHfHtN0b8GYkQs7I6Wj7atQRGGJjyMsFEG3NsFVy2O7ypv2b4XoNQPAi5s9IaHof
67KRu+/p9npd/nFa7pcYwTpqZaJvJWDtZ1GC2MLZM8f96XILRzyTD7cw/gOg60gq
AiuHyCWB1GSloLfJSxmkm6QU/grNQnKgW8nJ0XyxUgKPQIOGB5soVg7cIBASvpL8
6zprdROUIvPLWDjeB2leW1UApS25GDyVSn/hlBnvKJbNtq80er95ZY8PKWJnGDh8
/JwQW2LfT7ZoHZSJ2uA/mFHPgUGRB5IsZVTDAXF+96HziGCepiyyYA6s55Wm/E38
M5STD13OLaW39snU+1PurObgF01lSzVCWlskK/EEIBdn+L7hovT1LWU7lYJU6gdJ
MjFbCX4/FBUi1hKweEsLS6HH2cvUxuXX0JCNle6wjWfH2EOiGQk3hgyzFxAKo/Z2
8uuW2TLxfKpf3PKbt2TV1y0aUUF7DsbVys4mdIwWRnuzTASn81bk7bUj9YKjMhsB
R3u+Zd4kNSb0XuZ+ZA+ickiki9jRpQ3r/oGt4kGCilVGAaY/pAcek35mFgeKTTl8
L1gEDo9nQ2T209elMAnXbxsT6ljQHFpjqb/3e4lJwrIiUlFEmIdoXWc0jP/PhlNn
erkPUv4C7fDAtDOs32lcY8NasFbAu9izZ3i1jWYdVhtpQyjhI5NHsewXIXaapFon
sNTvXuCwKwdkGnb1tHarmFteqcOQDXlUc9B6v4kOW1rQARaIhIKZwX9cNgdk4E8E
Bsn8DbgiPSJv4DUdfJKplfiCAGS/QH2b5WJtz6uZBychw7ePR2oscm+GrutrlRpZ
S0MS44ld1nnE8qCVwxjjOJ5DVkGr4vqgnTIPxYDSBoALgs33W3tMv3WsCd2TWr4G
uRPwxE2cufL24OYXLxmylBx7NjBuu8WSGLam5sbUcragD7rboXOSPmIMl5h+ckE7
BrpliSpjoXG1HX+6yRTtbLtNR/KfcJTzBpc+tjYcJAlqMcDDllNkzsxkiRVmxU+7
QaYQdwO/1lHRgAdv6bOgFWgNFKn9TEDRB0JlAR7BC6IXOE4he+YZ4LF30WBVr0Ls
uRhFhlA9xJuiXo6p/5q/MT5Qn5Qy21JQ8cxvfnHDWIeG2q2x9D2iuYSVGJbJVaTB
UYxjps1Ai/V68CYOmtQzoN5jIe6p9artI/vU8pbUMiyGufEYw5X8GdXWc6M+vAAa
4VI6UficTmI05y/q5DMrZYieHYu7UgIYAg38beJVN/M2EIvZ1G2EymBMAMzXTRLd
Ypm4j989r+1z5GkJnbzjauQtyGBpmEq1+GW6gTGn6cxAMdedcCS+O3nAGreUe8v8
VaS+di4GYrvvurRL0xBH8d8xVvdj81m95ki/445d4Okxq1xrlctb4HAzRojwIEZQ
hD8GrzSI3D164/BiVFU8w9H2uhcnGWeqKq92YxT7+iITVEyx2EG3IvOVZf5EezKr
Op8Ph9302seGv1mLtLN8gKeV15m2Y0+EWOGwaoiuAFRl85MoZVZ1w1Rh8EB4uVc1
xLBkBYPwmsWihtqvNHnAJ4mQqAN+k3I+Ws/0Ai3NIcVmhrLIMpTxOO/bBiQjXZOm
kj+m+Liy2EEGH2lCt1Rm7ASa3cbI23k/Je50sclywpTKDJ50Nd8Fc9NNdI5pU+Ta
68z9R9yEl+8MXXvKRWELmgaGiefoJZzFVEdnd4wE/sflNFGD1iekVGbWuUJZBq1o
ek9hLqUokoDraVmwiZ37naP+eUIrZuMT+mu6vXyzmjIfn+rI5Jy4GVQl3zhlux5C
b6nLnhdQXxz42SVVTLuSYkEogEqgVasyamAonux+Ijvon1e3ydlePefQd57pdBfC
As5/IYh1qslOo3S7QT64GL4xUnpAUrvKKEZQ2JehhxkD3luzsQ4YuN2swyRxXNYP
AO9ymjjZaQSk66WADufDAmzgnmDs+0Ol2SvJLX5wfDUN0xe//ZxIJXk8rcGH2V2T
6qkkTybqaVlmFVCV9w5VWDytlE1VUwn36M4QAnF9l6cDoDISIpS2On3lNm5U4y7q
s6DGVacRFkXfIu9s6GzxSfn+28Z4cnU/eYm4uUaHWuZ1CeL5l/0/8qa1yakggFAr
4YQOwOFeEVLa3mxnb4mlCjt51dvJAHuwo4UTp52xiTfc02sHdxrs7dG2FsfJ9obl
H/t7Gu7v8j2Tll5dk5xHsV13oHrD1UtIAK8x/1j3apT1+XEK42WROyg30aO3PMBt
dy/dJ+Fa/IltDsY1iJ65Xp93XrCDt/xWqQGc4jVUgURE6AytlJDpQqvh4yaL0i3J
qU0FrvIubt9fbPyb2+ggHLk+Yo7NCYzzRUlIwePnnpAC2htKqUKHXXVPfANZKaIF
K7AmaVdVgRaPuwllpm3rLPYZ8Rvd1Ykd7PK/vFSvyJ16uN3dqMaha6VKeOsjpW1h
4asdm5zM4NYdgO18Lyy80bjJpEgHz/Q1woZMOoT8wenqpo3EePB7u6UL2WMZMq51
EJEaL993vvK0W+qm50BVpVkgVs0V17sbrQ/h1bcmfuFlJWjwAmX+Qe02ZGGUTZGb
2PnRVucvmiQmnbfy1IKyXkm/htEb2GQWDt8K/uZbwppmwWB2mQL0ar0oGhNAx8Gm
ZsnasiofmjSeiu/n0b2TaXszLytbitL1wselfbNZ7nQGckuyFbxCe+SqPbBAJPXL
Hfop4um98yT+rb0e1wnTXPZJDSW9Or+EKUHx0mgdT9Yagl2ouB+Dui+u+U+7O4bO
9Y562hBR+1b6kF2XofB8E7ILedENacb/VCiW6SP/M/vj7oDa+nW9RStME1tARhas
qmulCX8Jxk1v7Ag7Ttq+45KB+2cnnsP3M4tbA5KgVl7zW+SrHUV0ic6AGb3/BVNP
auVs8UGQjCBsT17YVeKpyWstXht8I38tybAzUjWlPmrow13BSni1c5oY9sEQE4gn
JqVtfMvoxNGVzH9KR6ZTdjOv8latrPDuOfsyZJb1tBw5xtPm207n/fCt+pj6QSHn
BiwDoh0tDXIDorbAqoUoOsEj8T1FsX9Jd/WXjlbyz7wr4jAGcuvHDwZR1Y7Pywlj
L1BScTKCt1wdJJJTR1Hua2hJUbpMa+rpjE7WO2U/cJqxbUEBtQyJ5AoIfZtr5eJn
Capele9LH1rNFa7rW9rNjXYDWYh3nRci00gUudm94ZzgIN1LmnQYRI8I8KEmjKNu
uXgp1K5AgxrGfwD9w/hAhpyyR8LVwK/v6bRX0PbNWMEXNW5wlk09o2KYQnYKRRFK
/sXxdf94Uta/3DhAh0IXecWSZgEXpCtY52xMKuRIozpurfP9oXLi9POpnRqgqHv7
qbqYFvNipBRBGDrJAf+HRhcbVdb5E2n1ok7n6Wjs1AmxpQGk4TY7tq7u6gRhBn7o
Ok1QUAcrWyFWbjrCTaGm0b/Hi97cAwjYEhUt2MiNcfEJtBLCh1u0dsMqPISaDO6u
jHEvZ1biHkzCCF+Skhx9ma7YKvPMDCskQg/FdRywtnA1TQPYpNepLRZUbsGdWTmu
ywdMLi/lvl6cKyPp5FSX9wSK7n4PVMIT2BJhzLr/fc7/hegEYFx7bT1m80n1tgRv
UyQ80Iot8bAD65zgE/nLxL0RGvbu7o41cAKedrHEpfM1jmEHyexd2V7TAPg38uVt
xP2NgM+rEzfN5hZsHLM2xl5ceIonhPKGhXAKCUVqLjtbWzdy+L2gBVYXBMXZlmrU
TuE+jPWZZnSW6Zztuf7J+s8cdhqvMHimAUeQlv8gXXRnQcNA/G9oMuORmOhSd+rs
0rIT46FGRGPVkCL6IMv0KaBeNClOXO9rv1Z39UQ+OaG+05cE9/VNL5ooxZQhasZN
GmRAK70TWSY5htSxRLa2RlLEYYil+o4NJ6xrDXOFoLSI+MjHNceQLmLYTjokLDnD
XFgTS6CCd+Ijl3eKG1cZBjc/WA3mpla0FwaAlI8SXySGKVcyRGdTkS6uh9o/3AGw
7mMfwdNM+o1Ehs2gETIQvrkm5LMyFceLaLBxv7uloAEkQtOzqEiTYHX3ne7RbW98
K5wANjXGHZW0QogVxcCQvIO07nFHv6RCu5fU8Jx9Dyx8yx93yEr5hN2u6bjeV6Mg
UelA/jVAJHb8Te9eLhzC7bVtqp1ONHTYNNBeZxqCW9PEjfGzi5Z8nxXn7hcrn/de
Yv0gtgU3enEu65Ni4msNO+70/H3pahWfdeJ4Ns6Opl3NYvUlLEAHm5M+zJPpbxBF
zg1Mwz1PvwMWne4TzQadmZpJv06nf0UcU2zYaKEFhcmm8TGw9Ua1TO2ff+5VThT5
HFxU7p8Tmxa5N8qoEQGieDTmvaf1hHKYfdr37zhaOvAiUZeSxGq6G+HAioKAr/sO
bBXNUFCX5vzAkS8HU7kgr5jRGhAzDspXTtansIEL9VPYKeZDeveR/QGfsDmwcEYN
3Xb1YkR0Q9c4EUu/F/zFI/T1Y75yTa3cToti79Pwng2Ng2MkMvUD1qict+VqN/v2
m5Cz1JkI6p37evMdVsZ351yRWQCVjMp6Z2jnUL+FGZxPfU6d951Tgpwq1enSdSzO
DOFYHdyTIqAFl3p7MGUzYUKXtDDo+/tmBkrtjcLzDa5HB+2tNv5l71RwwB1/N1qo
WCcoVSFqI5nNqvLlExa5CumTU6tPK/QDRVggSphdLMTeFPXRCkFafyrMqHyWBxR3
xalfb3RpITuxHVE08fQIiDPhAqub+GzrqQ0fNUDAlEqMU1v7xkJZxtf0cw+IiHIA
RFLI5ng/EG7TUEByK0ePF9hjzaI/JkPjRppX0OZJ70QPNgRwk4cSUwvl0XLrTdXq
UTlYltIuzJtRYMGTeRKcfggrV8wGLLObIDRrjWsRLq2ydd0xgcK4HKROdrEQW4Qo
o+CSJxVl7iCgNO3BNtwZCPtJ8rDxe5pj+zo67bURMQ3BHkhBhLphO+2lRMdStVnK
x6t5LXBL8bw8YQjojWHgjXDxRbUISbIoK1X6iBYpi7KQp6sxFEAP9eBxB5WI3XNe
ZiejhuQjp03O5tFincnRBmJkDRdvDbW0y0JRSoadJvlLqOchiuddM8a8uM9ZjSmW
JmeqBoYjqaxMF/ZBwAkqqyBjdGv26dsYBRygT3k8GHMaFNq7+7SsatRFKxkw1QdU
fSSLS3feb8fMswdZUnaV1bMOM7uGMr5dQv+k9uuQ3SFqwxGFJJU4lYhp2SpWp2+f
WxcLRJvJxbDme9GPecEybad0VV/dzPOKCuXH0N4D449BM6V5fPiItJdESN7G1c0g
M3MdJOZlMYJjieZwCk+JNAG8T0YZR09ezMHJuupH1RuKojhFLAK7mbQBDcMSzPij
4qfvikFbMCq7EXMg7fNHhf0pX6cmb6UMOgrBgCVjmBF+eVkAgfa/XY/ZcCR5noWp
Z8jcaqOPONcCf2sLnsziIy0B0KruL/HKl99yz6nab3ZsH3uWA+XepaJxSK0FmBom
V5LeNsEUX+b077mbyJj00QTvQh4C3gDFcZETTUDscn+3w2wC7g8C70Or5WpdQ/ca
tRvJH5BtKC/NZbcdZY6t2O971P+I6Ipm06EWW9JrnTQ8Af6QuuxiVmS465sYQuSt
/ano/E37l6fIVqdky6TxcPUVwHryFFmfwHjYqu6zDDnXorOvs3hXAoBRN9o0ZegT
wOEqB45VGBhMD2C8wAKFSKXgu++fp87Ut1JRYyyE7SAcVev/0XQeFhto9c00oxAe
+bSVEsk/OJaUH7L85e0DV7TCe5dzpR9oGRz88d+E7GdaGxEdVda5J2wqHVVu+QmG
+P2WnwKlalr5XMw0zHMTzPP5hYhNPsEiL8MyOg2K/neCXgXp9dlS1YvNWYsHN1HA
xefENHgLks94hRCYkwwO2UIpIaNFALWpGVGF6S3V5C2u2iCxMScU4yyfZjF5qvuf
G8zSPMWZ9fmrEBo5QvP9CNyd/iLJ1OiR5iQ2IVdiqHRS+nnPGxLuEd3F2PD7RzRI
lZG7Jn3zLhv8eyQg1tn+1uDCa3LlmrlM5BeahmQH4Z46U7Rzm5+K8VdPLZx+UzVb
UMLg8Fi/hEFNIz2NUjTmTy4XVVXTkWesShxYtcYhIwWvx6CcmJnLHb9o9eHPeCoe
EoVFJ4PIR45SauDrTbpLF7uzTxIxMHHIOdhbwhkvTOiAKXYRLTplb+61/mL3YrsD
4zQhNElsOTfkZxprpllJDBwRveY1v5Exq1EIbkT5mug6vhS80ablWkHObTzGmbEU
JExHnXcQTOrRXM++HQ40arAmtr/nWrRV9F8laRLuD7EdYoZku3mLqXoXCHJraSYd
q1AbGv5Bxj2bKSSOnFYKL+rs9pn3vwkEGq5PO9fbHinsjoPk6gCf44+JImvRskzB
udemw4UJqCEEvbDsmNPeN1yXTGxJxwjnJyadDpTPAi000uAU4nszga07y0fZBLMH
tpIed0w/DsWTGWezq6X5TzxvmEDeLgIHj7l2tQhOhxlbxR20i6l8jx+wyh4bO1e7
heEie6ekaGt7khmOeU6QQZ0wAaPDika8ylAqGTdNqZgzq0nUGXQE25ZwYDi00VlG
zNrauG6UwyvX6rx1RylDm2rLJExRvBblf1W/AZZgEN2661YjKc3BkHrh9Fev3tVx
0Qvo/RN+uty4UmXQ1qlaE6uOExZx/4cTL/3M/qImisN9LvLd8tCqrq4rZPd/tjA6
A2HyBtW+5mt92bOlYGKMzGtFxM5Rb8DhoV8Q2kB+GZ0d+CgFZBOH+d1AWeb9UBr1
kKT5PyPzVtNl+DQoqBeaYBJXeL8XS8nNqUSw+R5Rg7iKv7GR8qvB5bGgTsQdPIHQ
70Ued5KebVSPAKRiL1r4lz9Z1u0aLL/1V2vBVMbzrXXZEFI0pGI6rcYUmJZ9N/xH
lvBKQ+83X6YAALEhLXc/opDpDNCpndE2gMaAXVk7AjUVNPggm2Qu+RQnANCkxwGw
w9GBu8tU8roHqzHj+GylO3tE8y9HvOfjhiV4As4xNKqhBVlkDAxU65jTA0eJGgGS
dYUQE9d1mlBQeFMTJvIbqgPGDIhSw6u+cZlqY4y1/6o+jjnOD+XckysWJeQnR/wh
mppCASIkc7N11U7n4R2GoATrLIoTu3bBZz5LO8azLsXmCwmArGTYqCFQ7omvCixR
W5jIzEujme00l6i34+/hoXtdDjp6wJc5Y+wFO6vsEWSdItlgKrgaG7Za6QsTkOnn
7VVJKZ648SP6V60sMgfonosBtD1maig3LUPbrEUuHo1jBUiftpY8hhPaXV+1tSRc
qdtRkT3bjtaTsG3UtWas+b60HgoM1DSq5xHOaI7W8AqBvPVl1D31WH/BNbUuFocv
wOYj0HCSlHgVpPCszcRUQeEvHiI+uxx9a+ryL+HzykhOX2C7hAnJg3s/L9JMqdnV
nBKwARYjyG2tbCjQytIf2G9vN4yekVLc88ALt9VKv7qcEnDct+WmQTsR7mhGgdwN
Ryfva9kG0oQAk9zMKwqZZ8i0qfu0aK0rvCkMa7xMs1JD5GonQv5i/k2k18nE/nR7
KU5wwq1B9qFc4Us/J46FutztO685NeGgWExDG+LXqE1gs/sAZxB+qEp3eccsvVgy
1SfHgOIpqb11meQCBBqtISHzxKCjGBVLXSSSdx3FgwzU9BHsao7tVkN4pJg1cx5r
eV9hA1CLp01oN5n+Y1WraFo0DYhYVsGCfvDa+/QqDe8pV7bEyBy9tkszsKVWuDik
YRNCsJ/lPtKgMVNq/HUUzYloM7k8Q0eAT6VbFlKBX2dZ85/VbDly/+LY3wC/WWeC
hx7Ue6vVYQKozdWyvVrq/+sg2DDVBpmlfs2P6EjAApci3PHRpBtV5E4FJCW49wm1
uo0dqsmRvVazsKK1LJK87/k53u50SXZIjqSxXYXCc322EbO54GF+qTlRcSb7GkLZ
vcGzCaEbSx/pcRjvrVGPR78hYoeu7Mq0TGmgm5372NL/O7/A3qv6BxvBzdrvl+l7
Q40Y8DIHcnTsICbEUEigg4zfXcGbnQBR5n7Ki+jezr24r/ecgYGQfyUFw8yvgXOX
/DwL8mV15lB7WVimOl1tRd8Ac4cxvkTCiO3vvsRNjFGQhVWgO7qgPkITxzeJ0SzX
85xdE8RYi2LEfIECj4clFiFSNGRo/A3twalfbS4S5SgeHwL2W9TCymLm6pcjg9+h
5FsVPelUObkuXtzvZ3HOpXt49Q4axhTRJjgdpfNRgQavGWbMw4AqvZq/LljhRPlU
Mn1lmLT6AsMUap+7apu+jfUfxEq0UlUYuAdqRboGKbdmhm5DVtTeleK3nGrQ8ux9
bT20ZsRbEZYSUoDpGR6NSRKy23xG720zJtyjT1paRGacQ8RL8AoxSRFN5fu+xrhY
MMmHouBsbF0x0YQjPkXMme42sewaK67xZnmI11wgTpci+KivWCxZ0pc77dngLS/k
d+Fu+4GmKLBpzjO0BNc4r6gkugN84mSoitxSzCB/NJ9DpmcgURb0pNB1RruwIom6
dnF/CbE74ODqzhRGSH7BJEN9hRaED0QiEtMzyx1eer1mZk1xhO+7PVEBPVw7wrZY
ag/N/BtahP6ogLVkJ+R9hyT2TTsmsW6Ebvdv3wJw0GSSuDQq0Yp81XpGiG+SOkzh
HxUQUABiAXU71lT5S8+47Lh+TMie6+XY7GOoxW4Gk7lPANADo3+iLe7h5UAoHizp
abT048UVuRc24LAyvfn0/dAq5ilLjJ+owgQqL+pbl/u+EbiJ/GGSE3d+anZ2qp/r
Fz1Qo9AHdmCtyd/qcdPFgQoRKPOHA9Qz1sgj62OjKg+5R4Cn8xRozmvcy4GB5G5h
nuiFBqJVTU4WCf4rahmbW2azkj597oVs4xlX1FwviirTASLVNsL19/Xce9tO53wf
laosW3E/b8BM+1MyTfmiZin0Euum6nJhE3Yots31sjH2SibUnLLWLIHn/n7HwtZp
T0USKrGSvWKIEcD+Ljm9ypwJH9RdEqXZkiQFTChjOaTpkVIwcbYKF08sYGrMZ+81
93nsENrhlXyfFrmvZ4oK1j7uJ1+2nDoB1Fb7LHs3zNl45DVKESkJrINN+WLRUCd9
Mzn3myGcK7TuVCYedF2Omd7iBdFZgDRK75HW85RTeNmFgFHdX6tvodNirskC73d1
uVFUIAJ1BaE1fbIp3xvSIqGefPum5Bq/FmE1qmz1FpUriMskMtfed1eCpSP69hGe
oTJZ58BSjZAC8QjAGCwPrYvshB2dLexFM/KoCdg8lgEpwySbzsXsxt+IuDWypiGL
cg5VGggznObmgeZoCH0RsuNpjgZ5s6ZBlsDzOQlHic9sAsSJ+gB9VRbpWk6zS6CY
VVYiYdO2bSvhdUZsCTOBZzWdg3dpwnpEx3T6JoDRmiT7H+XFUD1OPMqaN6kiuFeB
9UG6WJjCw+jfWvbTTYzp9lMp4nZo8pTQqErd2SWd1ijMgcN+nGEf+V7LVeZL677z
9dIXlwEK++uRRKwPkifBvxgt13OT09tiLyo36cpGzjwKs8tmQUtCJon6zFxpU52m
Ye4g6ckggVuMqoP8wNRU0wc48KfDcO4g3e0JjqP/eM2sEPDYw1xNrbYcRalauyc0
kp9h+KeEqdEgOlU8WYRkUBHdt9zy/m4Vk9JvoWFkEPGkWb2Q2/YhnlecSxDL4Enn
ZbF70agLJJSsw86kQWqsH+2Ksuo1RhLyBqxiYPWTZdyXQvIoGvHxPRch/QSlsXxv
RyL0wc3BmeB5pvx6XYNiPmeHgdzckaW/sCogvL0Y8ezJICM5DyObeZwHqFD5NqQk
J/wS59eD0/hNIvbXpDFkb4fP4JAbV0L9sG3F4lkiD1NE+751bFfAdEgAOGNB0lqY
5Yg506CF6BWdkdWcgdLsjD2opAwGS/I6So0iqzLiFVpVOwcEl8T2/mdH/gxPpwn3
6cAxR7Ndl3n+uQ0pHVO2XVVICYKr7id4slnE1WHjXkI+c/R8mtRH5jGKtJ576s2Z
ICRwn0GUmYM9SKeoOHQhkh09067pcBeOtpnAZnGSiO534kPob4RnGhTEtPwmlSKY
niERzYMOF0epGPAQCSxOLu/ZDMZUx7cotWkj9ii7M00zwbc5PpKp1WABq5K+KOp6
5jdQm9yl0B9S7uMjMp5LNJUMEa+6Ig7Dvf//SrjE7VNNiGYjltTKhdzGBuGleXzN
z8rYo88fiE4F9eTscx19JKF+5kprj1XEzaiFPioKXiiw4FKCPSFhjTe+E5RMp4yP
HPnmI2FvhpoSjddyOP5JneeBAUnfm0deCdA1cOCy8cAxtBgYe3OrofLZrsoxTbK4
+hOu1zaarX2a60w8ET9J/RzIFKtnfJmdka/R/jUQr63oaxHr0RnX615BOo/IwS5O
2BUYJgvOeAa/6Rw3+YYuBeU88abhnd3N9bYUddVhGbewXtIActfafYtvdhUtJSVx
UN45GmOB7zyQc2bQGDZ7VF9g49HoA/N3StBbGr+ZnsNWcmuQfrsbsFhcGwHps7te
eKMnSUDZpN44HwTC6lQLwUue729sHPdbw9yl2zkpIpc7/ZUunqHVttvfoXHRJ/Sh
gzNrbqWPgTitiyJazVb5Y67/p44ORTuzYHitPhdYiGxn0TWmsJjyLuYdyrFX7zCH
i5zaJU+oWEX+ptpTCVDE18xTOLzslsuY4b5ATShYCSqyDvlyVjD/LqzA6vNj9cBL
c+I+pJ34mIdENHNhJ6aa0fR/FR9WtqgaKgK6O8CBfiUjIluM6fAmn+lBa8Bjl6QS
uCOlo+Ff32FTe/wzRd7grySl3SmECDei4pkbLgLSFdSgXgWqpIMbwmA2Lpdqn2FK
zHisD5tfepvgkzhQYkePnac17fn7xPcylOBDD4swFVz13uLbdTaSJcDATU86FVAW
GIgze2NovmzuxKLKCcTJvQm6tdrD9Xgxagf3e0skQCoLmXjv6pxtw4Ybf47Vw3fl
34GjvU9xUARZhtzQhfFzERgbEU6cOkkCi4n/IyVUq4p2oPUJwAfPViOmkGyvVoel
iduCnB43C/GE7mkYA8QnfHL8yQGpJqUTDAhKJNbS7zgt98K3zbDd95qTGFK2Krm/
4UBjqZkcAWo9ZVsI83Ti4LYF6HT3lMi+Oann+TLK4a5lQ5UOw+Ie3SW7ShHsit2+
5phE91lvz0/KFY9bQrS2blfKTaim1BlNNpMYQYH8WVlbufpIQ+5OraS3pm6LhzzB
KyHfTOTsV3jM83REg8RhG3jd+rWFFj86N9FmRiFPwnBfGsAuNv/h1YhIrExencAJ
ls7yA2eolzwzCPuvgU6VpLlBHBQF79vtoC+GESnrnZ7wAvJ9X+dC3qkRtHdJz+nW
974HabhlXp+u6dEG62vbp+MNub/6x1Fk6BLea8qZo772n3QGZl49r5nBloXwyqRW
kFtGTIAAZ+Kz4dRgKmYMGtaho+g5QiEM6XDAApFyr4Q7arMfhj3HKrO0BqIH1a0r
Df2PmiMe97lZuP3NOHNA4dSgNTHPNBMEvPv6kq6gBnPPiEZs9fCWPW9YOxjWEsSJ
9g2wrsw69n/QLw0+9Ockr3ogMPaBnFW5MRaRGTBMuzGsVV2noaTHKDMT42kFoyWm
5ADYtBtiCAGzYjnDUhAAf67XRDMA1sitRzpfN1d4Z9CwOwtV9HNIjXPweEg8ZuVi
fabKdbsGmDrya4yZQH0P3IfFSiZwNP+eMGo/EMuigSC3qqpT7WDu8baJoIjMqrME
pS/STk7RyF+k5I5IypkhCuzN8bi1e7JJWEkw00c8YGqsiD63v16yv46yFst8LFpK
7OehHbm9l1xuV+1Eawv/KuqEI84UcI57oEiLlwjlpFhIt5e3396EoT3MLqsHzo54
DKOIBEu7j4sJxHgxKNLLhmGX1qcUam1F9/8ee3ehbQIQ9Njz6X5yNNvs5xqleUuN
wke49IMoxGxHTwL9/+0nD0encGTlPDGpGkLYbQxTqmU4HYYRnP8sv5fO0oKU6nyk
Q4qU+bQfDIhxKWLQEYJvB/aKO274BudfTE0RGA72YWjhE5htNkr1+2AGEUVcm+sA
P5iAbG2QXQezCuYcNQU1tgJEd6HUrkfrjKNQlsJ2S9LD3RMKYKWehCneKlYYgIMV
QZ5PeI4ZwY+el5sAIQbKp3S2YvD9jYuJr33U9YBHGZNFNJt721Ql449PWoaYnDi7
ntVN9J9qCpWXpPI+0yJ0eUoU4WUkL0goTZS5yvZwlXtRQUzX8trtwuutEHHYMbie
k8bEmhjOIU9m7iLJNdkiWL5NlOSAPLC7zT3H1+zhgoz9a4aNXN3n9bUiA6IXX9s8
LHoTH3ms4JH6fEeHn891sZvVz/9/DsEt4N1VET26yYCfZYGj7Db+1JDZEHIcoawA
Hl5v4wyXE8dX+V0EleR12t6EqWjLnEblQpBNZxIdxlhKYsxhLRG+Zk5UV+uQrWf8
QZ/0hXTzIrlPp4gUDfnh3qHR65hQ/pqn7AFo5IaNunWtXqyKIwDIww2KTCHAD/mB
CKRa7eXEIClgCkzZJmgUGzgYbPDJRbmkDeKQn+ep12pFBh3yBqYGTW7gtKvzr3kH
siznsJLzNU5Db9RLS7YGnb1Wai82i7iz2Bk8w9a5soKcFQxbFEZA8IXU/oMxb1hA
9LLkeZII03bxfljENt4UyiG1bmiWuiuxEnz5pkCH5hN/pXIM+Y5q6SiEgxjmZ6Xb
/HPwq1ns5HZbsXCXuGnMUasETqgOf5SXE2lMUX3Aq5nJB7nzyoyQ2tkchzw35a6a
BmohBsdSd7Mn8MKwuhe69UUa/JRLeQ7BojdzWdZ58i77GVK5qNqS4GdRDUC5r+36
IOUkXDeeq6+o2r26sXAjoBqPbNOpqBmmpilKelkFjAO2gcJgEnqKuotMNBVuBQav
yO5w2V1VVzHUsGYEL8u6AwSXX2rqaXMmfPm9UpStuHYZFdZYxLayggDbtJzgqebP
IIJqcXMbH0OWnDBQJtvhol3Ob+kMMN/33mHN58G5bwjplWo2RpLa1pXWpu4rvb8e
aMNcb39rP1pvnRX5lHz1HcaTo7lwilNLxGwL1eMRrpagLDY4H1NkCDBiOlQRI1BQ
P0ubzn9kfXUBmbfcEr/Ok99Y582GPR8BJ7WxsZzHrtYw/D6PexygJ9xOYCk03DFt
g2uvQw0/FIhWGrJ5qK0OakV+CfwEf0+JNVqFwxX+7vq8i/tr2GE/Ok8rrwDGdMB3
aBpE7/fMGAMYWkC80n1gWb6pmUfxP1VgmJZ3ySCYdpEskPe8/dda3KnQkI7l+LaT
7yZ9cse5e6/2wuX0QfDzvZtsTfLHxBMFJ0TXSgIT6RIVOBWEihvlaklos9Z/tb9J
R/2ZhzakszHoxxskd+zOM6LOGfjydYQzB8CSmb1fcqi1nBCzZ9Zx3erd5KjzGyke
Ihs21/QkiXNmBIkdMrbvlT+FKp3Hul1uSaJv29iZyLZn2M/heiQEXDYI18DA/AWQ
iai+9dXjMsjMYdxoEKZJWF3Jp854EMKb4Q2B3oL27qg+vZVOGUjzg5Eb+ODABsMe
3K1GHFC4XoHF+PYSlKqrmAcLQWixCNfJ/JTpDaMFtBoYb4E5Hl45h1TTON8olU52
QL6nLzEd1/OjXiQBWrCZJAjb9kTzFA+ROygHBtrL4V93oBMwBbgzboL4AIsepJgA
Kh9xNpU/SFi6BbV7wo961Qexv7aULkZ6Wv2AfFSHEaYaINfldLM/pWKPZ6cRVAlY
FgGlM7RQSkqmGkJIqz75sE+OTBMQzruTr60eoQQwbcR7LMZ6W6Qo1K02iZOJoOYV
QapJytNq7m8h5C4tG27ICvIASN1Ur6p4jKXFXwDy3BdqI0FZyIBxdZnfsibcUY9n
d3DAA8ucO0vEe4Vn+ZV7FfhU8LYo3E+EDz5+IQ9espY++kn8w2N64bFAeJHXLnRc
ncpiJIgZL+zyP3XIkAWRXOzmbffeK6iIfty/qewF7ewtwyPYv5zcwdbUuGbWbyrE
Ied2JWuNJVV7suG12+TlcdVUHzgYr3xkw+kgPwo066dzEWJnue+4kbqd5OpcW5Ao
tx19RlbfTzSH+a5f5/vF0O7qCcaV20O1jaFHTVHKKzzEifpYDWBzYW64sGeQHyCW
8nEc+NOpeAVKegSGa2T1ynN9blOHDfprQ/FZqQWwpyJxxibQi+FqjZox6dv1uANN
pFf1Yr74xAF5U4QHMxSrUfdCwcY6y/vbZx2xu8lCaGdWDjqpWg14UVF307+C1ALw
dnyTz7GyIiNwpET/a3fXw+9LpYD69R5y2gZfJUrCJrRmY2/G/ybsYolgrz+ym+Dp
sQrr2SlydRBkw4c3852u89ZraW4aEOcbWP+aFt+uKzQ91BMIOFUt00JtTPczkljT
I5DuVvV+l8pDsauSgPI0fZufjo80JGOyiHL9MVV89n5TOQ/OqhRLkafCJDo8WMjy
MRW7cUkyEUzZdlmWI5HdwPfT0qa251tuBBPOmS3eLDCZGYzXESLBQXS2VbcB1tfd
fk68Xub3faxRPdDEDvjZItEigHvryBDsDvuICAwDPoHeKCKjLtO+KRXqFUwFbjOg
/dZchOuHB+gngruhMPA3QyBM/A5hkPnMAraawX0j4cnwjF/qAfZMOFJSzZMEAv9Y
1ATFiusydm9+4P7hC4z5e8rbWGrvFUOiGuDoU86MQfIBwsb2U2G2f0FYu/PwWcSv
4xVZ4LjoNkoltjVC/lwnpBlfNPo5IJxqkGlVLoN5q54yTmP+D5rnbYibomI0h/0K
K6NU1+K3GC6m9XjrKWTsMHW9DSz8dplNzrgoArO5qpMH1IC8BopUB8g1sggx2x4e
KfI7xgpmJvXlbuexcVUjUnA4Ge+cpM3uHFIVjnlUXjcnQVyRAYOwnngBjh/ABkh6
zOZc6xho1sYq2FfckR4ffkVcfcNIoFQd7o3f5WnSIi53TuHi+Xzhnj8PUtz+6EeV
cjuUTD5Sxt/0WofvmNycUy1trPBKu1LN1sU+3z0LEiwj1tS9xeVq8LDrcEqTHS9q
1wacM/m145h/Q4ndLK/rvqws26oAUKrJsrRea3sljfB4jkzH+vJNJ4P8MAxZXQgz
JrRuTe9rlY7qzufcwmrTRxMSes2J8OBFRfi7821TKESfL5+L1ZjlydTvTNy4mAj2
GPPWXNUMJf6kdWTtyx9W935TATfzzE0qp04RYRI0us5ntQDuwQBiPEJWHXn0Bc55
ITrRsXV7X8Dyb8mc6p+fnvmmUdTK3qjhvWO7aN7wNMesqGTLjinVGRuau7/Utf8U
jLcLE1NKwRa25CHplB5myIX4Ns28hz3IuKLEm9KanH9XKLBZYxusde6RDfrUQ9G5
u4qP6ubFQuXsvF72OLDtKMynL6ItCuVf+ZrX8nO3Yzrt19OR5ofPHc+Ul7k+0AtY
93vFBifK6AZR06baPCy6Jx41zyRZMH3BYN+NUqBgt3+9YmVlaAXqOXNiwJYAkeVU
pZ3RJPmPsIYphePNzucnFtDP3joqKcl4bOz2S1m2FQvtlX45mldHBaf0ADNZxo0p
IXqFK6ph4fs7l+L+lo/qC0x8Lr1Y8FoYvotqnDc1PxTYDoyQAFLg48ZON5Ragzgs
aF2Z1M257KPDuSOXNF+EQJJIQcrpmpFT5DeLMJHdG02fed6a7NEsN9Mif4Zaw1JD
3M3WPW8P+K1Fu3qFMMXwHGhHcbFvpaypvKjbmJSTI5hbfQbn+ajrKzgNG8iM27xZ
pJfbD5yj00XNuq865zAjyra+VjURX0B/OO0fN3PyP2Np9JqMIm2oFmuVUaNgHHzj
bvEX5N6+zWqNO2MoFvCJyAJXXjeFA9q/PNtgOww+cwGSkndeDvgTAg9EfWn/Jzd8
2Jy9a5FPQmVavr+r9OdUGnVwsxdAP13ySuIpISkzTwt/5S6y1SoPosKwqfpPtbBK
wucmodE4p7vltJc0og21gMCjUS7pdF7aqcvSFfJtM9nV4bwAO3rKuyeB8W+gytyi
dBxSPMLSWe8kV9PvGBiGUVHjYe2UhEoLoS3JwLhrAUbkZ7oEzlON3Bn2C2vBVMwN
v3wCOb5XVo09L/KG7ud49fNyCaXwAC379PrXg3JI0WGAbl4Ub/KuKEit/6c4E8Au
j4W6PvLmZCLwVQ5YMiUXy0LdKuYS6AZ1YhpgYyT/8qmF/b7eekn4I/Bd8kVIEqxG
PZRpKN4GEmgzrOa2MLU+0dP12pPd1nG29Ud4qxOHaRQ5Og2FprRErHhSCw1ybeZA
7wpFrTzg4SiXyqpe7QP6R4X0eErJTMfYhWhBr16weAeEAOqcjFcJfPoudNNybQu6
n1VkwUeWXHnTbPE/Ft2tXDdLqO/qDPQgaRDDU3p8hHEvEGDEMrRFQIpwzY6f50j6
KWdnbQpEODg/p3JDzuYu3y8VeAaCSDfrgfioppRPI6tabI7AoPHoKfUktuiRJdz4
bbv29qV3JGf3r6qV/oMpfVE6FZeIrbcWeTBaYi1N89CRs775mknD7TTYX03z6gCL
YyFRJJ5OgWxnW3Bps1EJVC/bk+x6yXf8FE/LSm3ZQitc7WUF64Zzdk9KCNi+/CFb
w01Pn2hPjb5vEQVOKIoBsQn4kLNYHRfVHnsSUpFK84JckMAqK6jkm5YPDov3/TiB
T3t4K/yj0pepCb15B+Luq1pYmbH8adwpzk0RHGtaJXrzi54RSY7dHx/vRTjhUqQq
GZZRhzk4WOCDhUzpQyEbccwU0Z8rNE6xN6J4hGaTKqrad2wT8fy4k1ZSYOPEQdXA
knFB5w0IiDC0lPpbsmFchtXJaeJ4QZayegSLoZ+d62pfLi4vmvlIElQYIbX54Rzi
2p9IohNOgUPRCvHLDZXsLfe25Qfc4LPa3j2viDUZpvCSYz9oNnxGWdg9pDVbf/Fo
r3VE5xI2r9EolGv01jgAOWLPary8zLGlLyU12SBYmmiA+kcagmvw8yhX9/wwKOh0
6erOKplTstOpZ/UD1ihkpyQrmSjsj93yxS4EV65xGb8hVpVKLWNsPoH2I6DJtdpu
T4fnNXjYWxtK9Aan3yMUW4W27//TZVaDDFQTMiVxKNjOE5v6Fd8YGjb60K/KYne4
2fQJ4yKEGROfuI8kvNMb/TpIxitXvEj3MciHfJuqeZBYWHmtUGJJqGAnRkvhQOi+
I51N1q8yLl2N9571eisdup2obUzJywIkfQifv/Y5OHVlIDvYj8Y4s/4diXi0xyo/
dRwGxA31f/JY/VAeNw0zj1O/ePbLedWue6SGu8Ek8DBGZbDfnWWAdnWFRHh6ielg
8Ik0HStmI3cGRIU7A1RnysNDxtoZrqQHL4kKf1JDBxA43E6EEDEmMx2JgjU6X/Gu
sw7QfKp1HJXA96xJq2QFB3u5pQHqG2K697Nut00DbaONl2wsLUMFftIlweXWntDW
t3WoJSl5tsvGALgU430U7fpbVcDaQtqcg6UllgymU70RrSMrj4+AToUOO2I/bxPS
7GGxaZft0uw2FxVPCOopdRCK2trjepR4M1My2f2QTUqXaRPKQ5r8eOpm4q3LyqGA
bn8gDIdr2uRqfF/DEDj5rHYQP712VoUq3YRcB4fshYWAu62eXIEnFPMhom2Y5Oqa
XJmuozTvZ9twSpyKijpKFCXwmbnRNIFbEZ93mnMcs388l8cLqjdyGGbu21bWVik1
ARh8NEA1VsBTrqXpvFDTb7lvOxdN5xYKu2gVX7nn9hybLiFrEXFn4gP2/whMvr70
+65AgJG4jD4ZOiLdrVxw4Z204Bnm+RFWlNZHGAHO805yNjRSCh28vmLLmuweZH+K
abKUY9PA24lakfrYnU26Og1VdnWt3FyGb+/yFbijG1vZYoEXcT9LCZbABBERfmIq
lDt68BvI+795gF9SydIkTE+PBxGTsfIC5kUYyYh2xVFH/+qgRL7ZXOs3IksxdJyi
nBT9N+/oLWwGv0hXgHjOiQtjNaaaECvVJQyqRTtQ/wt0+l0+Hn/ikC1Dkb1lfVxv
t+9z/KwCWu5XZKPpe1dnBptsTpP2kmXFLL5oHNTZGnz/5JKHbv4o31e6AijL0Fuj
yZroYMNDsHzsjy5H7gI1gFFcPrYNoWJXHgzvjtEJF3CISisp8y4hI0V1EHFv5MYC
kn55f1Qr5XvDdZkLw5pdMqueABSfQRvYzUgi4/3IrDw/DjJgiQcwXsdAQXvUouLF
OQui9FLWMTE13WTPU1JarBJ2h55yFS9+l9yImR7AU+Ct0Q7HMCgz1PRLnC2kkFND
4ss8rirNUoLiMChTmkzF4tbaKziuhnmXsduQQOIhaZ2xVEm7qRRVShysweQSH/it
iF6pp7semOonJ98HEmFykftEea4XNhmIRNYgLK4iE/72FlQTVEM+2hTz9fiwXeQ2
R3U14Sbyi79/5CIw7Uz7KuVECTssAwAxI1jR26Zn+9aWIwte2kDqGLlAZ3udD21Z
TH40S1N+rJjcTuX2Q7JaZl48L0rzr7AADx7XB+fT6QQdFQ8N+vF5XxMV0YzCrX2o
3v86Zc+f0iDc8ZFfe3AZsvwOjc7xMsvOG80DcEJszoUgL+1UjaHOpLeG0jbQoMGR
IL01l/pXvGzzbr8l3ORRy+KrG4f4lJoaQzp3/o9gJu9F5JujEA1qye2Nmgjj4kCa
BIX2wjABJNftGpumc+N6QaPeufYXS5KjnZseCjRZzGmU5kFbPdQ/J74FNk5z7TaQ
OwRp1+D63iYrXCOKSJeRClwaDshd3PgSW+ES9uDaSs1ww4rcwht5/oPX8wTgiKqg
pkfzYMKFdi/TtSpBS2dHJkCAAFfCdrqIWnyzH6RTovCRtILvLEsl8jE7djElz5LZ
zsB1dod8mdtT0bJSeDr3hMsWmJ9GIU6l5SoMqR7U/LVE/T2wWVqCMXx2EqcovHlW
XPxb2in/EmCyoReX7IULwfTcEGm/pEs2S6qbzYfkMIV4Oj1ZVoLg6O7i/xCAvD4a
6v7qpduft6RKODRNQrXMNaCXn1WklOHCTKaZ/p+ap70regTbhr123roTiNHQ5ELX
3g/ukpFbVSLMBSoB7+Jk1scmhP7VeInrY1ZFaWsIFLbltti+0FkFHH7tJ9/VwzZl
2Dgc4nWpSDOBNfyMGZAnpS3xCUYnMZvnmcGEVOPNP3nS/3VVaMvLhgpqkQcbjNay
7QRml+ptIJ9Xk5oNTogO9AVF0P0D9eJqfF4qX+YejWr4D9KdEwIA2cHjfNMMhQzj
rGscSMA//P73omJp61VI6n3cXNVh2FxQDxEyBrt1O5HmYl+su6Syamq/kYAmerWC
lGZDHKkprCcjJB4XQfyi7yPLfyhyR0xiZ6RDGMZfDFnqiY1c6bhejr6+xlfe0Tlr
5puiGQs6Cnbp+PbX6Wv14qODDHHhQPqmuZqT2XMwVlGkmdWvgVWqTu8VnmWk9t+/
LmT6skRIqgZRKeOTC7R/WvicxQxzH3Shyay0MuEBN/LKdPdq+mfjETzQMopq0F0/
Rkb+aJF2W89A6eP4m/PIrmvyVacu2KVoUTHD1q2PGAR0yi6n4PmPTCl9ccsUuOOe
9m8uZkCnpsKDwvGBW5vlaXA+4lmqfDdhQO6pBIbz3d7m+Gv8yuH+8EZU215YxduN
Z63tOOfAUhSaxVocHGV0uBtz2f6LQvcTwPcMx0A91jK2z1rhZDZa4dbiSLD68x8C
sQuzA+nU2Z2klbY8+biTPlND73R9RK99IDD08bG+lhvhxgpp5IZZKFckYR5CMiqu
+eClDTF9z/EDvjy2obOIC4Iex1AvIGdcMyWTxjC6XghcnlHHEL/N7Au8HkZlXRVi
aeOtPjSuJlecSlHOlzVerRD1srjADbkitR9J80pDu9WKH0pQKWX0Ed7sRp7fQVOe
fnyBnK8VyzIpoWiO7UIjN230VO+JaxAVrDlLDwGA1jje3Fcm9lP+LeSrr155AdDC
9nOD+xkbf1A0LsOscVopVYiDgdTq1av/QxjdChVvG0PyJswCnT+Uq8uhJfhnodiW
bVRpfnOJILTu+pSuriqIib6R9frWiVWnRURMmRv0oyTsoO4sJ4gtFGcqQEFP7b3Y
yRjkFctDdC1HYsxlFoGt/K7OqolzsqX0AkvxKb+5VXmwpjP/qtSEStBGXSda6xqS
nJxz791ZoO0IWgpT/F69HOIKVQN026gTWMEXIXjJmLy2ARjQIB32qmletC3yx21F
KAm7/4G1GxDIYPnLAqLX82SfI2yXqPw23QYren1aKG0ONj/fctW0n0aAdEEU1YKv
CHNheDu7IjUGW3w3SAauPKXhnVBzDhdmqEQZGTJYqjr0dSZhl4zlTJh91k2cs6/q
uYrNO1r2BexRhXOjVnDuGI6lDH2BNzg6BcOHbyMsFYusrw4gkmIemUTKR0yfVneT
YMgko7MPwL6vV3/Hrxf7N3DrSV1RmQsConmtUnuO5TAay2xdx51eqb4taeZ98LRu
Hc8jlZeNZthm+DEFwZI57XZjm/JX9WLZCVXeinc2u/n/AO8KKZM6vH6KxyO91/md
sKfu7g70WEY6rwLNw7qJkZij1LjMfx7THBzP3DRbsvfr6rRE9UCv7Zy9Es9MGK6h
hUEntoR1JRj11IcLQtOEqThgBEvN9omxw1HBg9FXWMJXTHVILem2kIBIo8xr65mk
F7ZYlaMAL03/Y9wrAC7nsKwbT8thy1WM5UT10M46/D2JTCCp2wlmjtk6VfIOrHYj
CTpjidifWWA7q84pa+ICEI1Adi3pz79+t0TdY6L9OOhOfFWMB/Z3DN8iB5KA6u7w
odn7A4Q05p6GwEcdjX7mXHhRo50kZRXc+JpzJlbS1j39PY01v2XMnyh7N0dyTUqy
3cTmuXkH+3x9NHNK2eZUfDxPb5ZzIJzuniveZlk/7PDbXjew9hNcsTIvs5lgoKuP
SfpmZbX/4Ft5aQFeUuGX0VC25aPNbOJJd9IBmGVADONbT6v61G59u0zajo2Bi8NB
BV+6sjAKKB7C3w+vn9vomG5n4CY6Lk+9u9EZfHVfR07vpNqmRR7ZUrQ3wRp8L2wa
ip0uZoXvjfs2ze/3QFRUxEp9uf13S3ZBaLMnIqdzp5guIovwEQAZgTS2wVLCebMz
cM5k9Td+WojVOMeJ6SHM03nvyAR7cZdgm5XvJC5KGaxZf/kkkDfqQkLN7FkdKfxD
E9fks639NrqMrTX8vIond/G8z1I5+r2uHTW2FLICKjr3zEqTB2muGnWgpW6HU9SN
snhpJrFNCRPAmhzZy1baCZeX4rIOGpJ3vH7938/GhcXwUlZi2VMlp5rHveCVVfY6
iJvWdrl/Qy/5Z9wYtLqE+gyCBbBan4+qrf8OoaRdAD150UnhVP51E9q1dMbdmxWf
+FUwLchHhgDg43Z8BX+ywxoKYIQZaL5V8nZF4662CREvKLQp7Ch78E7hrH3LwgIy
a/lX6sYBdJIWldHnMjoQ6xPrgHjitFTkg960HJIsx+xvJPeGuTIRSl/LD9bsFGko
9BMqf4BVIzd3le61ZeAkbxgvPIebStU10et/8IrY5WZz0zry3NLhGTD8r4QqU3MX
/xCNiyGKAn8pct63YsEzLJrAfY9mrDq0KgSLOeWfeQ65d4NvTfJv92D8L+JC8RMX
r1MAHdn9K17Rcng0ICsgPrxvs5pcjNcp+bbYgflH8UOMVqllcEN1veYutaiUqLBi
ZattK9oExepCP+CjGXvPh20rNo365vJhYqEpDWHDf6wfi8nBg4d/UFfftw+GBz2W
rd+mzE87TCQQlYvKF55HZQu0aReOSSUIZxjLN0iDTAefmHxNoeY24GMEkfH2Z0Jh
YhJOG6wrR3TkoAoVq7Ttfc+rfSW8/3Q0FPmfOyCNTndz2ccVJpwybJefXm08tvdS
NkqA4Hz0h5PiklWwxnRk04adOdIshcYqosYQUS32N9nNsPYkRFUIpyP1ZhIxDljm
LYmr8TzmSQV4l6A5YSZANzTUfmAWxKmTqxWTGxuvEQSEksFTqcGrU7PfkoPn53E/
LaP39X//Wcenyxv8eqjWu3BVhSJjW8aK+gnlRnb5AIiGtnLS0UuskRQtysqOz8EU
pC8tY0MuaXMT5cG18RNeyU65DkjK1bia16AXjIk0hHOcOEk0gOuB2f0uJqOYaQwC
n6XpLKEqa9/mUoOR3idzwt2QMv7tAVlEF4In3ca/hBitBxwAlhiXgHvBXGvOC9o1
9tGpuk/8hOPhO0yRxDOCGsiBJzmFy7j+erkyApVfcj5DU43Y/Kb8RjAshYTvjtqo
cOdKUTdGYLe6yvWSf2k9dZm2xzcv/cm2ZgFcR2Hn+trKPLB2EvZqDyzvIAQleCC3
n2pvNdYJj0Rb+EUs+Et4eI9d1hDbahBA3sgPkgufA5Y/rmGRUwBLf43iX5c+0yro
Gr3MqXRmrrNL1ns1KPRVMVmURAyUofXA6QHvblveTVfdMZACBGQcBHa+W1t1AqlZ
/JQrKwAcDl1ToZB+CEcaHoiT5MSEys0leDVG1kPd73u/8mCIZX0Ki4/Ruo12MyxB
IQvDN8mkb1iEXxq4R1ZGtPBr3kNxgoD2JU6qhBmaT1Q8k1kS1tJMNOeFTiX+p3jD
YOZUqDd/Nst09GZGBBL2AogWq1qVeepTRHCaXjesBy9a441UaCiBpRe0qkQR/e5K
pyGnSLwlSJ8m8gtEcFw7PZ/yJWd8PYJLjYU86b9Ds2U/wKXjEeGDsWfMtv74VCyI
HGZds4Bq47QZ81mpNBDOnk/+J41EGtBavDZERd02dFwoyBsR/ByMnVwaTQ4Bigiy
DpE/iig/Kei8dYlx4b9VFiGIE4wCItuPiUrhK0Vx4dUPZO84AUjFN86vhuitnd7p
g3U59gB31BMm2NJ33BoMkVOVuvtosCwdGHFLRd83kpPg0zxVz3u08N7auj3QIAiS
C/WYQr3tqQCqLomJfhX1wbdRnwybfyO11hrtN9GcPaXvDfdwvTIOnu7a2M/rHq8w
+r85zy6HVnvxW06sHruSuHbPKJkGtUEN7qsTBtLfHZIS3Lit+PV2m7/QtX2xY3r2
C9pZmJtynR5LzruG4rtfZ/9BL/DQp6flRxw3XcE+Ppel20Aqdbq7RGeYP5FFPQGw
Bew0pEbNIDgpuGNdNwahRNcBwA+LMLYsd/ifLomVr3pVj8QPWM5UqexbuyGHoZPf
K6R3fA5BwtXBhje4NdoTPwURrWK2vIyrKRWEfxBEIFco/Oiv6fq7wiFhliZftWgQ
7AreQQMx0s8GdsT+2ds+nsZPg+2DVtkpjXFbxGSwEGBoGj7J4hUZRdeGCeliffCv
6mlSnND/MymfSIUy0AfDOqOoq1XkB5Rkevw5xCt/PG4SdqOR3TD5MJdn+z0/DrJf
V2dRRkymBc992TGtCLi/Li0zRknqoOyI6F1+aJAVYSXS/Tosl/C8SPSzHlVTClqC
ZwZloHngMCiJpKQu5d0SRJEweVhSbhGF+rtCoESM/GKOIX9VlNhlMWUDE8om7Z1Z
J3BFZA22modtNflI/ZXag4FLIy/Khpq9X+dkGEXkZIAhNxFzhdvroxYf2O/nJzBg
XYFJazkHYLyG4rImsj2XyfLYR1s1t5rkd/3mNRM5fqI8d2WoKdsHN/Wq6yIhF5C3
UNKhWHMbzDy0WR0ioNs1qOd5ENlqMhzTki9+/1QY+xofJjxl/FLeQaxj55EVvwCQ
LVWc9hzhH+kn66nHPhdbEbTzCXZRf6l3D4D7MsBATQB3CZ9kuWFHn7wwsoFSKDIZ
8Q0qVC+WgLmVa54G8p4eQzIxaDa8K/+f+aLZl/D30oUmj32IfTwIXFts2ed6/1q6
/Jo5G7mj3YzFrn3TsL/O/CyM3/KVFc4clEc58yqJg/EFB474GDugptie8baxHLGQ
WXbyjRCnJfDulDZkBTsr1aK48k2e0Q7KVpXH6aoJbDm9VBLeWNhCqwKd4LtguuZx
Tb1c1U2o9Mzfnjn3ncbDWxjj7EhBheGUkihZJAPzZHGaw2ZmaTkiJRlae9LyNqiw
vxSq/k8UmSazYG/RBndTw0ouMKVmvf3gPfba5M0a3jTnZ1q/2e9jJi0mpTgCHPqR
VkFnPHAEXNgKFgsqJ7ebLfNL2tXPvZkbw9FNKlnxgNDOAvbyn9MJMUxJlGUh3Yco
D4RmAkfu4lXpmS7DRRBuWzzQNIQcw5y/0gz6s/aOElPlrGKBxdTEk3GIa2orahNM
ES6L7TjLqKC5erzLT1j3Dy0LafQJOqK3gM7xFtG4sqbSIbY1hMtdzzB1vGojhgbi
dL4cYxQWOod432I9ZWx9deQCi1KkdOQuLUTAj3ugeqc8EiVIUjTWPsb0tywG1v2S
oQlBGffpQJM5LB+Dq/I2mHM1yt/C6GlT541/WTLiAlhctDTvmim0kT7DuYOeN5uL
ePeRjvdHpLtJ1SKL/B9Hl+U8fWUJ57kH8uYt/uSn+DIYDPmb0M8KwBjFuv49kAOj
DmTuOsi3dP/pi9+AYHYrKVSNhFyhYf49zr+TogN2enh/bC+cG58EQkgH2/91GCmF
E63Nm4CkX8UIod2dWXrwRls6uA3pLIEdNBYEAJVyGCR6v1br7MpAAnu2xo73vNlX
wRq7rUuRTiiKv9B8z4RxyszwRRbujqzM9ESJpACHznPQ+ll97X4XWWPpj7l1GHpI
g/dBk5J0Z3j74D8Ss+z/+hkidyesJ4Vz86LO8IfE3fB8IQP/Uv8tJq7UialyQxit
XEAsjYjdTOUZXRKn1OhbeX5hrToJUaFDqCIGXN04EJQ+oDgA6RHQaRjz6q85GdVk
39erUVdOkvibcxFVrs2WGt7uXwpNwfHg8hZjPM1QiPF58cOzgkiix0lAwsZGigxc
sczHiJrNoPRVBEFeMAJ7u0Xp7HXqmH0+c/IhdLECih+6Dpz0vKUQELMOW3oYtdYs
1csPwQMB0M3jFd7Ierul5gbrIYeU9Xq/4zF/GdJxNdV00w58LffexWzXE6RWnnZ3
kxWx4oX3cdNyduDBACjG6nKWnV0D3zQDeO+o84TKd1CIJQwpe9iaEVb/Jx125Qim
ZoO9lbU5Niqg7/9Kk8hQ+1SLmrLd5DGx76k97V7lLH+m4UVaSSyxyXQ49XB5pN5O
y4KkDAqmwOUbMkmF7txnoOD4qih/wVDWBEpgXO+Xyzja9Lazw4vviSoK/ycA+EHT
J1pcBVNi7CXT9gpqNwagxdNw8BNhb0ywkvEm74ouVKgtT3GGJIr8w4ir3VQthmZr
fpJZM5aUWscmDR/ALCv6ZqDCKRtvMlw/i+bCyJieCoxe2Ltt5HRCcYN4yaYxMeGp
zXCEu+nEHBphWIfWPPAKFgC2UNWtdC0SUpwnCBQrx85ezjmVUsWRaHNL7zozmKHC
deVG+agFBN+fYPw6BUv241877n3xJE2fYSShmrs1661Vy4P9HjhPkO/bAfot4QB5
wJ+PtMoogEJw0DaguRCUwG9CDBooO3Hjads9ITjRZoSPphJdS8BKZ4cGiGNRtUhm
5EAV/NCfe/wTcl3b29taqWFdJrHl1/jYqerOZptuSbG1kwrDcv/QzZdd+EWRY59+
GSnNMDXe3eKPs3p7+6zTtBXWroLAo3ufE4Jmq4m6JwS2r0l7xK3N8juDwQQbAJ2t
IqzqIZTeGH+wPuhLX0j+Qi5bAbfwaQejXSsuP3YdBvu8Akj1LTYrkPogdfFWq+uE
mo//MDHkJGblep8bZ2z/27cRGQmq+SklL8UaA1EhY7nc13YRyKHrhx++TO2s8Zjb
6eViw4CmdFdLOudxSa3YFOOuxzUDFRQ9Cj5UbiSc21X1g9WdwQOjTYGzrwHo2p4A
47ld2M1n4h5wEdIwtRnQp5Tt31ycIegukU9bCQGGtek9O5nnpg3Io5EKoce33ZLZ
/97XDIEMYvhi+5JOrV5Eg8PIti6KawjpxGi+hq9Zib/CVtsghaeumzYINoOfHcHp
pJP6CjXkTBLNBvrm8V+lBmilYQyJI8qLyD1nkLp7EtB0rA4ZxNuYeCCLRWMrLVwH
9oZhNxZSI71O83XTYARI1yp2L1Dxsz0mAToqIEk48Scoki3V+usF8bCB3mkZjIEM
NDQUlfgHrUiV+R67NpdvYiwGwU93zp5IkbZMqz42Pxhumie39g4KoMbiR3E/Ggc9
28N2MepIZRQ0sICq+4/ptQbYiS5qEIsgZjdNd0L28wWY+jN9w/cmWkrV68TjVvPP
/PCVerVOIp3inRvJSgPJWJsdinDqjZcLA5r5UmsEJgrouCAARk8oTB2w79rG5ArE
BlBCX+PQ8NTKAXoTC3G3xYz7OMdtjb/CUUvjt9vZkIltQ05fVA9k2QFnO3u2jGqz
+LCjtY7zAs26JCLHaQVlvNnqI3KkcgP73C7jCIAb2TNNXnNI58ndRuJ5upSPbvCr
eK/FfvB+x16SCEudCgK9qTydwk3BtBiSl662i61H9e6FziLW5Q2LLRPTOwYqR9ZC
qdQTfN7Me6ItXS3g6UP25tFaY5A4PBhF4b4GbmRQ5fAyyiTfDqGGWjCqxwp7NVA/
Bt+sU+lPBc/wYNXhp9seRjt6kbxsOaL9rVTCc7crHIdMjMUeOc2im2hJZuWMuOA+
iS++O1cepwRHrOWSRw9Mdp0MozFJj9LlI1U0vMaNvLv6HiBOuTlmsgBU/iZAYyBR
EAYNgCQUMHbix0adlyS/IQ7323m8zGOksLk97xqzaulumuJNeNECgOYBLrXSjJmS
FNwCtocOcS3AxRzwpmpsh+QWTwwhl+bSLUatzwAsMUmAQcWEhw4/oPMHxMgMpc2o
U0PQK7+1Rz+cBaQV63a8if0mbr0TApi3gWThjS9JnZO5sARwwfttXJXPJFxxlPki
sFdEN6Vzj6qw919F1hzsXtKTuJXYOt886yFGLbeecKglJmigo4gGOCvrx0FV2PF0
tQfeiCDJExnOLVY3lSlQShbQuDQx0w7NXxYqWWC+8v5QnqhwzNWrSyleZm688yya
zXbsVweMf6nrrJhduXYkC9FIkEL8tO2j1kqgZYN7xw0jwT55EIk2yndJiOH6Pyoj
cNQHUaOWDmlibGcKqgs28csi68ryB3eHYBwf3w+Mgj0nBtD5KmCQo+47q2YNSTLj
RscMZEMfWvpxhc/IQg9QP/SVOrq8wOg+jfEPC4/gsG9TmTYxxcqIDZyarPFh91dn
wEXVAA0nrrG7Vkozcs1HdzSSsAfjj27PF0tph0nRPwJdqR4+1TH6ImkVJ0sUugdg
Okt4A/w/w6W6gr3hSqeVjDnwXHvCEFIeu/8wnUYMWxoMNH7mGec+FLz6AuzHc5Dh
S6THm8h5pSv4o3NTZ11uMHNKPGQ2UpcjnBzgkQo3go0ElItnxDIKc9LffEEXpTOB
PTNXa26R5dGEd6XQMTN6gOCRlH/RBmKunBP5+gy/hJfULVAxa2KyTttAlo9hAIBB
+R8dZ8IFVipV+0U+8j82j3E0HMpOwPQssyDSbC0Tz9zsoZLNRszmeqZFf4RTp74Q
CcfG9Tn8mRNoy48YVR65FwE454+RdepafDNb96GanntWFGmirVPppD/9bMqjwhtK
3DjQWMdEV6yyvzjrAbCgoV0xeNLSbn7WnU/hxpNPgBef8hiQSh2SZrM9NLGxvMkz
FXdOGF1I6N2WUSlfG4YeXiMm3IfGDOMX858oyaOt+P1desxHweIpfNpNsAqRdzTl
vqE8ey6c6GjpNCwl1SDDmj+WBlIxhotHkXMzBs2eDisNLjmp3Ovtvz4KJZXGwsER
+cJEeQlopbhh35qngTcCQmZmkm7CZQmVgGeIQtgyvd9tR6M+n+dhoe+KYKTd9cX1
3/CFmkJz4VPtCCT5FNjqSFujPXpkUeSJSJVDsKleEZuPfy3mVLlHERtv97xNCxLC
jnk8fQcsKb9BysO9zSckBbP1pabEuJUxKVFd7GzZYQGOIFjavsQOFc76ZO47HZgg
rpHxlCJ1NYjBpSU1UdE3yo3oTTYrF49Ct+uLiSLZbZXiHck8OVt7fQaPC3tR/wFY
jsXyim7laa+BcrXhdKKM2us2rf9c34TYEXuV0qrHD+SKTskzEmQJOgKLI7qgXDw2
80mVSyTMpGRnfwtEqjmNIdABeHO02TEIFfkUJn5glm3BayHaYDuCn2C9JcvfrWbL
p6QiEmwE3AqWcz5hmZ+mvmzyt7jwa/ocC/Lus6xXfI16UlFPEb2XciG4yhfXeK7J
lXjy6PnACO8J8h3KB8D9d+2n40aKvLgh9OC/p4VAn1C6GzlKq92UHOXIoXlM0/yg
zZZE7k9NlAz8DHObpa8QjHrks4Bli6r6r/K49SqKDoCoIs+QdPu0yDTr4cd9mC4r
4FDZrNMXOYK7FAq1fAphsrcC4Ea6fneoHHMK3QLfrxJjkmPXlw/JR9Hvps1h3bc4
N1yn8OwL20NwD8/qlom9ids9ZZGL4sx658BSfdTWgHnUec0iI69tPPe9pfXFA1KT
wSbFgsQ5eYxIT5FBViDXptfxW/l/0NFRZtBseetBClWmCtcV/fdK2QoSuL7lk0XA
JiDwbzmxf3spuNRbcQcWC16q2Q9oj3k4sJeK7aVYkiqd5yK7XihYe67nYAnCDRcS
O3UFVRM+yZdalx+HIZ+bUbh2bN2e5KXY46sDr1STCqRQUwpN6u/pDHWTOJj8Sd+x
q8/Nckp6izK5+GbMtAB5QTBy13Jhhk538RTiSUvQdkoC585OmBXA+O9kmrrNM/Ul
FQQ5qMP143t4Go/mOcRa9Uzg4+JA/bz9vWqnmhTG4AECiYBrnQcnl4HwkrRBGNPq
f2SfExNGuahQ2Iy+61IXX1apCMMyvzE110tSqwRtfE9zol2JaR+SBG42cqDLdsWk
Q+pxzrlNEPiglGDznex4jZZ9LTaq5xr1bTdHtvejvZtDW09goAIEHPnK6xhalich
oEV7/I/y5bfdRKRsYvNKqAaBBRstiisFCZnZt/mzg5asicxCoY0VI5L3EWDzIbUk
GaR0vtw4q6OMm1evog69tHSLtt/NXJLRYW+YItOxuraZpi/E5jDa6HgvHDUQVBoG
csJm/fOnN97m/iugZvdF7xS6vVGLoBSKSaef+Zib3vC66qkldTechhbJ+Tne9o+a
AYI9+7IN22WnpTdIVtDGdOG8jBWlYzRKLopKAeHiQVX+7HqlaLWmCnpmd7Cf2TJO
APeeDLG/PEgJrZf6zcQcmWxiOiBwQRGbiubRMbm/Mt14KVxyot3oaca+1WySNqIJ
jWSZ4JlK+g2YiiKZp3L/epRU9dpBnoPk8o31459hUBb//OEmugBWAfxs7TKFxbA8
jlkyPWFKbu5O7Fw168F5eGwToa+btlIgTLmnICtvKxpQFEElBW5Ht0O5jOCc6DPu
JDfQ17p5kkkaCG5jeHyonKmR3OwO09VRswqxn9sUvT+OUB2cokx7n0wNbEV7LBIj
YgmZaf/wKUVuz/gjQaae61qbOK6Ho5+FMhSHTQhbIMeR6t2d9SIx40nNowc1wW9z
FgxZR7YhX6sBlXWYAlqfYd3B8Psi97ZIui8LJxBc/UeESVAO8WPZbMHqB1y/fAZo
DO2ZB96rgw/TFxc7+MjNgLqQtXxpH1LFW32h4a83QDODV1vZfp8JBac0t2wQJd41
fHtYH1DzViHQkMr4K+BNVBLJ5LSha7O1PwrCv/HypFJrV9dgbOdaujU9OqOD0iyj
tujCx8Gbv/fQ/aAwMyDWTIUCt9TvcYLZQGU27lx25+hRV87bW7mgnEZD1v7JFXtI
xt2TrX1rPImdf1+dPnWO6MTPFnZkHdJvpKBn5iMcq6+YX73pxvHF6k8C5vEM47Pr
TrKcM1xbCPh1I9eGRZdqcKjgMxajqwBfA0QtLMcI97gBdNoNPg5ieh1NrBM3S0xi
hhfDAeCPtCKS2vgc+y9STcoiyCRF6Jo1QtKnXE/MzvYgmpf+rO+KlzFAtMIViB5q
uuf0yrqzNaLWrL95Z6vqhqJyQ4kyn9c4KEErEliFydHz/1+Szkj/E4KHwBoaEzXa
wgcfoBufanC5GKl85iq4zkxOGALMD8j9AV1GzwKxls2mD+8fTnCQkmgm4w3ruw/M
Wx27gxcgwlu5/cTGBYn7hFwmsHSamJfnUwmW5dQaEY/dw6m1fuDsQMYQKlebEg98
mDcKjr0fq87C6bfi9Tr7JdWFJ94jv/JolwDbPmjhedJwmrTJ8fHkSXp5wps+VpS5
1jUXm4y5j6KZvah/i3Fys06I0OyHjk5X7JkyOxbQDBH0ccRp7MS4XAARfUWwgfpl
WsoxTotFdWyuuBB4h3DPPgv4K0mI8kj5PZAGLB4cxK8PV4GHSISl2xduCpWF6Pqp
h3seGrdk+XMhb3HRH8S+VGOKlAuorX+X1oORAR08oE+wc7jzyFyLTI4s3pRcnvDG
HeQFWSaVCkU1btImPTXys0LLoPCGZNNtqTTOvw+jOBW3u1WyyyPFibpK1+Tlvi2l
vbXAi4Rou8wMJg+XoMtN+HI+8+vQGovFdk7U75vPvOHNgW1iDM0FG6zmfgKix7Sk
jIppZeyHs0LnuX1KwpS0G4aoboAAXNxjs9VO5XrRbJTRfhGUo8sTsv2hfzY9U1MB
RdNFK9+AmqLB4l3gaSfYivV9fwzl2/GZJlYGPMA2fcUhDLdPRdGQVk6xyg1C0D0c
VwuXFe7gCtu8o7dFdIfZDUsTjraXg2jUA2gWQKt0CUyRjf8op6GkN9BzOcl4/dmX
LUCaiS1O0wr4vAzabqlIRKVhFV44GNQz5jJ4mCmdO5UkBgj19tYBjHobS44RloBd
dTQCIEGN3OWCmWDsbROKlC4QNoWp31mDADWMtD10/2fahhnoCauMVG68oQGXRTGJ
liZuMm4dddM+hBfhsOGv7xFQqGN1nks9LNCFpoxdfMbeupNRj1ALSKYdoJZG1Q9b
F0yZPuRR8/ddzldXtj7qCOT+nSM+gd3va8KbTZewb92+68YO2jzWpWnYsSeLbhd2
u+nFXJqtu3PzO1rUYwYIihhfgHW5fElZXyci1EfoxUOkC0jOafqIfWFUGmehWTYx
fzMH3aWwXxUQdgp352dnoVD/VcrxzpME0cDUrJrbkdbRmNDNQzm5rVewdZzp8yAi
xA/uAl5ZsQkx73kS4pJppgZ//i1H/kNP/TgGy4iAZsstI42MktY/vZvEZEYABHm/
IHwF6faBA6gOIz0Yq5VFfciGb5zMkjdNq40zGF9NzKRvSko5jvluN7NPS+Bs/Rt0
zi0+WCzWx4eC8M8cuR9EBBjVbGW2Auau4Mcd4H4KjxQ3Vu29AxiPejHUMcoRo6dy
wa9Qsxp9jVxyv+FjGtDWZSleZi7gATzbzG68576GdRAF7pyBUsL4mBv7hi4p6BLh
IIxoEth1jla73YVegoVrLMsLtQX+HvOj4yDy574hIZ+5Z7oFkCy4LtVLTNLK4XHg
khaLQOxm2iE2HifUYsxzckqFSHjQEFQU7gvGjq0B1rWoD2ZQ2PSRGrlnHiQQPTb7
Fd3Pmkz1NbOh2Cxvz2UDscpAL0EuvOOxG7rIM8qVEgUQVJXejWTzimqz8rxl9VU5
EHIPVBL6OKlGA1FKgU0xgSV6rar8CiYXd9UNuLlHKANhyW2jzjJ8TvC0QlEw2bBL
8tHyN71WPPF9nQqkyEG7JYzSKPVQA7zig0CkMHpWFCoBea+GVpMepGa/I0fHpzBi
ZBMMlfACllNPq4krMPnrKwJfpJZxzI5EY4WZUaIODami+WfdhSe61stjAFPxkHNL
brG6xioyzzdOjLUBeIN0U6peEI5Dy+e/E5Xqb21LPV+XAMTL9AQ2guZ3w50xpMyf
62VFQUtuG89xxQtVgJWl9wrfh7R/R2LZKu8ukVeZWYRwFl8hmSnwUTxg6zokrTuR
u/QViL4ibLr/TCvVdc4JMlWWoEW9FovaF/bGvycylB7Pp94/cuwPFR6OQDO2Mk4R
8zN5heBoxl0m01YLy92X9rvoWPp6DBSNozqnvghlsxgS/vU6n6y59NIVOACl0uHi
zqu7BvjgKS+O+VhXUgVPopTrMyjUv5wnr6GGNyxItUOlELg4vN1KNpRWhOcZhmfe
aTUUTfaOdcsceazxSg7XWCWHM7TsaYqttK/kPlyPGOHgysLZqL9bt18KlyQ3cLr/
NdGxT6mwSxyy4kemb6JMyBfwC8TsqnoHSTyUfmor4Ki8CiuSMhQ8dHXHNu7fqlTe
wfteZhdn6cV51EFzIvZ1JpzWWKvWtgar4GCaf7Z/fzYT3YZm2XGwhjQbCTou3CRA
lKIGrfIB912LF2Vnff+BBRu9qcSsPMQ6gf0GSKU0nOZKmazNGN67spqetg6j6skD
9+MHHxBIsPRe1Jl0CKW5kzIoKTCQom+thFL01eQQj5j3yMZJl3x0MrIW6zww7DrD
+RUajZgUxrbvFJm2NstrjiiQWBjzJ7pM2jxqmKtEF3xsLjbs6PxEC7Fhz8AbTjkO
NyTqp+PJ66wzbxfPN01ywwSqwNNkJKA5bHqkilpVsnb2R+1qDiDYIJD1van4jGdl
4Qqod+llUNGEQklfdRoCNmhgX5x9VF1oiNoSuOFMFI4GSFz+05nim2QSSB+pwDsD
/YUXCQyQCBBgP5RfaLkQx7SyVFtV+x/6Q0k0jxHDUL902DguygNA+mbb214KVenP
kg5L2wiS19zcAsJr89ofRfOxc+k5ScC5yRavaYA0zBWkX4WVJ4YMIypf/4ASl4jo
SGeueaFlrOGy0UEPd4xgwA7I/Pyu+DwG/UMEYPiKkmhTCJT8osBwV9K54EWqSxLs
/CqGwxKwf153RghpCIk40pR9567qGcbwJCm0PaLAlh+7jyAQlaZ/63pPbW0pKlW+
RQnM4or7zyPUjQ6C66fpO6uFNtW1h1+2YK+pOcBfVChLCQg+X4Yz8OtochNogvDP
9khnHVz9PISSb2nxO8paXvZ3KFlDkHHkxFxa9Xnuv1qNnOdYBvY1PVIy/kZpYTMN
Gk5k5zscXem5Wfc1AUIW0skvvZjt/wj9wqB1P/2WMayv0zRS7msbtrTQIY/lbjsN
Z5aQddA+ERwQMS2XNYdxkztV3Xzs5yniD6wrwKhOUqG7Q4O6JzGS0OEf0sKH8cCo
qb1CHNS8pogYf/HsCy74IxRyIbQK0DcZ5u1LdubnQiP9mdkrZgcgOfIJ7Prn5o+Q
/Bh8ZDsAW7VnQ5ZKoHDA/SRt4LfxmBvjHcRutGzcgFQNR3UTbMsy3CYmPH1nmWHt
mkzcXCnVLhvUWxkK4Xm+cvGKexUqZekWfWL+PY9grai4o30eg0NulEVrWfbA5ot+
xpUAw3C4YLWbEhw/76wBS4RPmDmvMmA49REZg12rcViPQM59qjnYNH4MeIX0sLck
1b90jYUp624EAUxamyVlPkF22f6sSVhdIXuJwMN6kT/fLBKuzoHpj+ics151MVnR
aRIIGccEouYHoK9EmYVuDV1WaqBC5oODEG9lomQJCPynR4atRVe9XNI2kN2Uv1Wz
aKxG+mesTHFBDGN1CtXnLPaEW4RpauQ1OhgDP/W1zOY4Eh2AnffPjgYsN02CBzd3
LqAmSzLqzZHXjPwc2d4p5A5tPe9zjvafJkC5ntwX9L3ojKNNPk2R0kZvliQ26DOk
f3l816/Kn6zD8jtK2CFq0b4+jDzlJeTrN1+dmFm1FSOzic1wYIbyifzIZQs7aIWG
vEklSGbKPacwH4o2UptdTyDGivyiXGKnSDf1efi43jGu3muvOB2iNh699Hbga8hF
zV6EgfnphD4LNVZhZg6VGL+4MMFhxetcOqk2kjdrN7MzFA9eNXtmAfQ7CQj2zTa3
Z2GcLSqCXmGuQP1JLUxn0Jc4pn2Cvt59kL/WwAzsyvYWWDAoBBT93QC80ZWNM2rD
lmGvK9Yn1UscbQUcgopwfiaEWo3XRFEKH8pUqnI+dwzfG+X9ZMy0IaaycXnUcXRD
tSGZvcqcm0z299WkyvHJ6J/LElz3uWh6oFb/blUO8ZEN/+t/pf6dKH9MDnGJT98v
ktwmdgLp3hISHWRdpmwOhZVxIncOVjZmUSKkcRarUK0INcdS1BjM32QfdQUtGe9u
LRanMvUGhq5sNn9HP2KYYxPkWkb+/CqvMnN6MAv/exvIPDfY6euOSGakpatx9bgD
TQfJZanYtPF98IStwZ2NAJs/1Rw+cGFN8+iRn1mAlCvdWML49yM8HXc3cVzXvSOH
nP/RSHkdzH59GAC7e0yVcXvSiynoQg3SX/MH8vZR6EJtQH1hlhjNoV2R5BnJw4P1
z80GpNWEfumr64Au0pz4hMlwx14/naK5ine1UxiHd75KkYnd8Q1LTZIvEWUp+A2q
qJVas4xswrRGTWfnHhp4yjtDfSkTz+lZpt92ZzcxDCTm3lZoDPKFs9AZxUd3QgRc
CIkxRiAFKN/nShMORwGL+qk3pO/HRxTjPhwCSLw0uPDZ8dUbVVO0TUVfHEFvPAD2
Tq/ifme754i1pN7jnWI2dAJ+E78Rw9/5eSH/hLdLb0HV4vnPQbA3KV7E1Ob65rbC
6kERZu5E/YRbWRBxiuH6iQvn7q9W4CfiRGL+BOMf6DZqHQ7ycNWi0QAI6A41Go4u
YZTSdzQjteZWvSjx5lpM7iq6Wvuudfr3twga6rIVpbOqhus100FvDtz72mYgaoS3
R3E+fCScEXveIaooQtkpc7ZV0v7lzNVbR2+/xGUBH1NImV9zS1nDZlRU54YPGrWY
W47bnnYPmycRjfJIak1KgJQfiKzLuthgB/YrxFHpdd2PyvlE2M46Fl3FIkpwcjZN
2kitNL+WMJtK3vQ8tGrvM6ixrwLUcYLYRaZoQmRp1Xupp+K0shsJ5yBfzXbkQ54K
ALghos+SM7oI3vhEQpDsavYZ4N5fi7P6nPlvwZE4TLh2nCCjEVZaujZ3cb7RZOtu
gK6qp2GUPBAO5ueGRR4803ZKU7XsJSHol6KXPxWDxgG+pOYRXcbBpVR4HnNLO5U2
H9SAtIEMcyVqV8jAJgEPozG6mi4VpypAWWyBlH2rHxoqkCpKQ4Od5JWHhmZ2ZlD/
Tph87RcUfpbJxQ9viKPIycsNPOxXpgfpB7wmD47z0OvM46yThuv7nhL1aAbexSEr
+n7OhfMxYc/Cm3yt1Dv/VlQzOVX22QNoxqQuapAAimDMucORg3xBGhpyfsue6LnU
K8yareR6qaGLE7IpLd4FbViNh+KLXm3tZLOaRO5dMQR0lpc84TBJnGC2SBgeORJ4
fRQSM+1DA0zKw6SYdB4J+7r9LHS/nT9unK2VL7Hr3AJgZ1JwjiWiOzBq7sclhbur
tWwQ4GjcHDaOIIFcN9uhDzPyafMwb85VaiO8jVXNcsW/ec49MxD/sPjQyZ22EAdF
5wmjxCBYR21nFKTYI7oyAlj30/66ypMyTV6/6FK4c2u15YVR7g7Io59axUYl3295
38ktU2/KMxjAJPnzDwth2FSwdd7Z/xT2U88eOUUBuvJ66s9QgC11oTX/ZCFv7k4r
bFml3EaeQRTWSwCVM29AgbVB39S6mMRp3kTe78qpg4+ojO8ZxulNJfK37US11iTl
GFw9p6cYlW5n1F7Ly3qLLbm2jqQlfrHidX8DW/gkCKbaKvuhhWTCPouURhvLMzmy
JMcC1R22bYY2V7jBEbofEflDPbow+Sv2iMory7zJXLPYx3iaPa5r+h84qSI8pJ0h
6zdB1Tl2/qJ1O5tmD4zzS/4M5c9zZsH4aoDKi7N2GG9b5/INVvm4YioE7eKxgjis
fPZLxrePxUwQByUnsed0HYI7I5QNVjosdi6ZjtuVYRUObDyIRsM2LweEwpY0xaxx
BFHQqDAtdgNQAcYqMWyCfiHGyHkLIQgVggAa7VwnspmQkyINHgARyo+Li/kmg7Mo
hz66xb7KxLUjOCcVsso+6QJprbxd5GJQvHGr0i2BcuTq+chiKkuufsii5aVwsm74
BP5Zi55NATS3FCqyaopSMOwYz6AfOs7kJrABm/F7fI4DFo5e1reWNap9Kamn9njA
0O8rc6USaGJGiXjrX5PJbotPMHEsQ4izVMAPg/3KxGaYlSTEfSfiAfgmD7cl8QgH
LC2GtxIREBBHR8+gqW7XtNva7XXp7VO74BMm1tzo5FBywmFQVc3EwNEFg/0f7Ovk
9f1Lm8uAyJlvXYFt9xFC9mVISTY+j7/3YisR09a6HWjvFtt51B+79byiaW2kHoG2
+UQCDR2XMSlS12atOPjoDja7sHTN8L8YEixqJCSYpHGBe5d/gnduv596J/MH8wiP
5v9jSxG8qZsnTr/kbTwpEZfwAuhrt2UsVnSqmcYrGlrgR8WCE9hlED9+ra0ELR95
KZyr4LoMwMwEqMdMPxVMEkhGe4bbjNEYS2a/kVAj5/Ig2IkitVGpxbPrTYnqm4lb
4eXhABpwXydqsdw2J9sMCxzPryVRFBUdw3dWRPYKE/MiQkrgJAy5RjqFa0rmjCAJ
loKfou5mJU+m/tqdOklBcoU//UQi1cddQjvASA95srDRVrr8a7l6k8znEsZCGxy4
K04Gr03050cBKE9zSmsSn3nPUWsg7hcixZf+LwO5BQowarIjlz6BA0nX+IKlNzeE
hTcsQHjFkYSIVtd4aum0T9AuksYsCG6Trn9EdHjYrsaccBEPUcc6AaIGR/I/gEmz
hb4pnAsOxPepPpJyWALj1OnfY1uvHZM3syohVpMq7FgyEadD1XQW/CbPImvhlJ+z
EX0fLcDv3sgjR4KL746u1R8D4vu70TYyvu+1vn69pout04udOv9GmvE5RRQAxhl6
XpQFwnwtCJgb2HoNe9yEbKKj8cexAinGGy8iN8wMr197N4LmepPXztYr/VhQZyc2
+Af1A6AUx6hGUJV6v8y2PGFwqpUe8kHNpH8u6+MbqB4NtQj7BLd4IaOw5dLAj0Xl
cDHVog5DqTQ1de+a0jVERp0BoS12rfEf+YMyIYc9By0AmaovhBVPFNrIiaBNUmhP
bPr3llFTiKP78+xaeGtMYmxUZKCo5RVnsrXr8UDig7i28QwqKJLQvO/LdoP8LmVY
dTKAY8GBGM2yaidO9kjxAD8GFlcXoCHwyR1Ogz3iPTDRFyN7w9OAp7FV6ciT+zHa
8fApIeC4H6Vh5Ao9WxM2zl4HKuiPDkLmGRVCIUhpqJ+spnU/lqAouJs6W9DJA3AD
gVvi5J/RVjI8kC63T9Ns+bPFO3jqeKGigkKIvLO+Kuxl/uIr6svQd4wGXnb7qt/3
nJEWDDhdgyRU1SgfvsTDVzWM8airLS6wOvWnRCUydxmtuhbfUW9jw4XItRFFioiU
VHCVJ2LNRByodDfPNGOUyCOI7EVo6jsZEBVkEKXNAYC1VjdLHTU+8l0S2bpH1EtJ
MZ18c9JHT8nfWNBBGDy+u10KeqcjjIIHHujshK+9TQ3GZE8QGH7eLCcTs129Z11U
b1vbjGRKEB/HiwvhluT2UeLxv6ngcAEHXPbpbeaUFdg/wK4659mauFg/1vuMwgJl
EsTxQ/Ikx3mzoPcOT4/3/p7v1fQBIQb1mc95rd2BDCu4P7osuHo1UEs8S7LefU8y
Rn6Wy7MSXVB52YoN9sK9SiAQ82oP55vREfUn9HnoFupG1u2klC7oJXjvkFgS6ETF
cTr0ukwBbc5T6SJYjnaazNYLBzGNkZIX5uoVyMhddK/VDS5/BiUrZ4jvHis/BP4P
PV/BS54tWwT+D7hKcWLzQEBPTGysgoBlkyKG0smf6wofegrzj+rdnMTB9TZ8I1B5
j22GkyjP78tf+O9lYEtWMoagsd3p3lmBMtz8Nq5j3L8AyWVjvjRjfHNzt7w5EhMl
cVgUYOGC3YZZsnk8Hp+JZXL6XDGsBObzFcWK88aG9rE/OZ8kuEqdhjKF9ugAO53/
clwT0+XidEgIMDBkUEPCGBSKBPYaZrRGH9a3E/aWnXFQjMpAfJBITd+FiBD7Kl2x
OJQJK0FapqarHi900snhWcTToGU6K47pB9q23yCSS7g9io09awaP5QcUBCZipZZL
ozi5x6nIskBzzqWTi8ddMg0KRj0tq5DnIqGr9c8fLOLC9b+kSwryjQZZbSkNaBHe
TV86yOlvI6V0nESPV1lUZU9s11miAzKCHvsxwl10vM2U9u5rMqlPKbfBzjkRHobg
ND0lobPSDbeQe//FfoSuN1k5FETsZPUAQiHj8Le9dqFW/LiVFXdu1xNshepurR2M
8a+91PN81wT4x/0tGZwfVK3/Ud5arU32UW92YwvHhj5BFklnx5Wa/gvzfI+vrlFc
5VjC4siipRz86DZOuaXfGP5uvI35v4eMELRuYpV/ax3lag2Iwkka+8myPVAhdKHj
XjVkmI89y462iqQD6ruXDtbSjy5PIUAsVSVWShKIjCMyOq44bU+eawSArgwlxGTm
XFw/3//N8Y1UQQwLqgIut8wHccc2EPGT33gU2ZsYQo4E7RDoO2BAcVUvOvsQIfg9
LvGBDGZeYnWubvacJ/qCLTdFJnIEaV/kfdlQfKcZWXB7s9hls/2YLJBBWcWjAKaT
PNaii5YCYBwTk+hhsP3PP7zwSyG3bRkrmY2Q7P/4PAmO7yllDf0NasFW+HxUW5xE
7znEPU6N4odmVOAzH7wOsg+bWaCWoh8eLHLigztT3qfypROTh4IHiuZmHhnW4j9q
VWA7Qzo7ZXX6FCkf8LahdMtV9mvJgVYPqV9F4YfH3kMIdN9EH/kih9/wgbhPHrNf
DBm5lgMXsLw7dJnj402lfMnLkYju/xNY3frlb83mR8mJEEex577fkxhCqJi1aQk1
1BpM9NjzWQCCKp0cQ4Hh5gzV6+ujJkN0kDtgeH2tCZJEj0xuvkBY54tHvYuP2t9J
0vNRFWArhzUhbiTg3NsFQe6Xbr5RPL1WiqmbiFqNUfna9sOcivaUvJKKH5tvW6Mo
4TRo4LmsuvfS5k/iJ6wQhKDvRJg3xrezb64HSDftf2VUfHQ+XJNLfMzPvCbRh3Wh
3bOu9QEoGobJlbL5+xTgau5HiJVJkc9xTtGUbHk43eJ95k5w86hSoAEhYZj2Wv4g
TKVbRYsQuMgRWwAW+w1OCTTk8Cx1hm/L7SwtK/AJKDnpia88/Ghou3fqOPrbeICP
Qb2nUYsjoayGvMBNEeu/zeW5PqIfekRPKpp9VtnpoewDTNWyNJEa5J1vwedFV6/S
X/oOMqYD+16sotQMXs/3SMsnafYIUfuAOPuYG3zf8reBezrkLIk+PFMHdS+y5KrX
loXH+rod4H8uhzoiCs/5H0OUYiJQBWL/D/gSenS+y8gkrd5Mq4oof0mdhuJhggEY
wxDRtsiYS0aKfb1WPdNTA5p+BnDTj6t9alv2Dim/Ycvwk/JIQTbqu0/Bo41A4UYY
MOBvNpKVPesLSDll7/HMRe6njerUnrLKzf2u5wUJ/pp+y4R+1lFT6P1lInXu4OLk
bKesn1GtJ/YWYNH02TlMF3RL5IG3NGhDLGEUIq8GM1uOlXV5pnW3NuyGrbLn99zs
xSWsFaG6O7z1hJ5UfDz48xlWUc84yKEXOYVUgj3wUjMokEwV8IXCDsSkwjdMhXb2
iD7K6OalVrf7FEI6CCzg2ylY33G54QKobsDXRqtaMz8aWOAByI0eM9aD/6qAhpO/
/Vr0qVFTGWAjRjspRK6OeD9ltKDGAMNiys7eznASJcfY6NGCr5ooIW/xjWIzGJGA
WRiR/R1s7nN0Yvw3nlRniQaNYuA6EyGGXtG1o9iP96qYt0SkATekrtPjgtoLQYIi
z3KzlE+aN0usKTkhZ8IBB814Io7BD2lY+EIQw5k8HaG5yc1iUdMvWGxi5Uw5r5RO
A/qQtocct7nLjA7VbtQxgBAD3F5YrAuit2eIm8UuZqkdU+9VFTf5s+DXPyJfa+3R
ggPOSbpJBZTu+PYWgyUfLbzXrHFIgTYWLKcRi44Zfb5QPMcuwTvuK2R1PNAY264S
kUY3Jlj5FKqH8LswFj7Q/yps7+Ck6WlBQ8UZjusyWZSvGA6RC0gsRvU4TiDmTK9f
4oWfnXM1t5ivQrIzygiPEw8CAuOQp6Kf25sdJJ3Ey9fKFiQacMymfM5USwIEqY8f
Gl8nyu8KR6rQpsQtMuVgL6yaYU9ckn1ioAgXLROqwz0mQkDPlfh0ZOigxKJ5OZJt
1JHwGXZh0/Aj1uOMHVXgmMWHu/APfMIyVjNVBNe+0p5fORHw/FzcjUSH29g+Xv3i
6NyjuG92n1z+DuV8IrX23Gn6CTIXvaGcih9HoQ/S+d1RzkSGXVpjGGA+7eImQscR
PR2Wedi251EGQmTGfcmpVmXf7lYbT00T5EHIEkudj7j5UHXQfD2QFv1w5A89TMXu
M3zi1lFsqZEXb0g9THtwi1tEbGSg+Y8+xH5EbWDP9LGk4ZyOgSOESkY3kF7HCtIW
etq7rdfxil4diOgbpXF2z0zb80PQlPCnhk2kMyy5NW+J82uptzm/DBHSXKOD1D/L
j/K8gQ2ln38Qt9Y9YqDVnpUNcEmZmg/cXG1fp1d0amA80pePYztVl7C/1dLf3u0j
nfwy1qZN4YfeYZtqkbtOPlidcbsMpKzVybLynobM+dCzq9TGgrWLcZ3+w1o9tU6Q
41g84Mx35RLU45vDqnwUFQNUEKPKUvIQ2DEzABlDDJUQOVjvOUFcaCcRfyecBMoM
bh93bJT2G7PTFTVRgZJPq7CWADVt2Ikh+I+YfhDRHo1Bygus7Mc/AlBoi7buj7Ie
OcIJ+mG/LmwGTsRwNgyR73mgrQPJQlRYqxlzZ9/ZCCiWBM/nQx5Q/m/orlDPkjpw
WBAuGapZfuaSDi2OVV7fxPRMk1LYJ9U0yR/OvH7HXSGoobnwEYOb68EEnMo4Tb6l
akj2uwkqJjJ30lgtNYMgR7Kxxu5SpQDkMrsQBTtZlACs7hH4X8Trq8+TKRIsTW97
4VqlIOEXztjzK26735RI6d1O3EPcAfeQBKIvC4ayD5DGiXj54R1WQUvfJIV15tI0
DLQhsYmtSm95AQp1g+RfODyAYpQ66DksYTPWFdSYePHSevpXbVqn+ulMzuxU9n90
8m1YZrONxsk3edcX/g59Hx4keIKXOBg4FzeBOXD7Xm22TNNUT7WEO+dSnC+nVSg+
5/ztwDYY/CudwfPECnjKBNTpjjP82Ev+XXSJRpgla5x4sCzf49Y+oz1hU0oGUC69
4U08SCdM7QbSKR9tMhZHpEIbPaVCGOAOQLvHGVY/a0jS7Ea0F40w8pBtOWfbebii
Z5FVAW15ERq7VaqXG1Tw6U52ZMqkx9aq2Oa4jfkogM77yjdYz9QGIIMx3jdcukDH
P8R1BMBwAOJ9eyUi2iRGZjzChDd8CMgxw+Ur0y5an6js5hP601qp02/9Kuxglo60
o5Pu6C1Enzoi+XSn/jmij8zVmVuBenYNXs3bc6aoWsJ/h2W0tLDvPTrQ+Ct1pChA
td1W+QE6ofhwQORxrAt6M4CHUSzkLXGxrKfwSTHL7LQEohAQkA9pGpcOaeadLcpY
bsmOdxPKo3cT75bfCQ0LnSyVZ5eKQCkBmipnFMcnunXis+38xxGMakHpJxjn5tEE
xZHjZ9x14zb+q8jgZsYR+4C1GqgyeYCs5b/9B9Jpbb6uK6UGNxNwsVkW9q9S4jbW
G7e4SbQg0A6LrrLXzm1IWdz6TIneiFo09P2LIYHPXnEZ7FVWw//GmIcsLLJgx2/b
fF0lJydiQqBSKE4qU73fefeEaWQ6ReAfDg+5UCOnR69wwKfhDNsGyEwswgkev3hD
iLaI6QWBNgWwhj1kBQP9iW7dDZpW9o9/tMMqF/YX4LZjaRnjg/HzZNFGoCGIPova
kGlX3mYObWOZImPb+FyIfotJIbr2324FQ5imNGgJtzxQIQwP2U7hbNQPZutvjFgE
ai4199bKUZcasSri7LDTXEVQOjLKtFy89r6ri4mDpYv38/c6XS45M96gUstd9Cem
vrHg2rJaoylX7VFHjT68ot3okzKNoYKgMvmtiUP8t4FI7PEphxSkoQxypnW7CRdX
r0zIuXFH+9oC5zwmEIfg+z0dD94UvIcDiIKP5N/gcKjLlT9ipXDVjReHZIB0fySv
sHq1pMclU/NXvAAnBYaMyrs//RFROeGve3BrOWz04sBx+UN19r8bDGe6VI4O58I8
/kfsv3vbKNVdfafIfe5+o+QBzQAKsUgujFeeX9XD8R2y1W7s2z0dLx1149Pf6GSk
wuYSdfO0OXoUeaGzna1B/FLNqv59+XIV4UutApu9j2P7O18gC+M1LViz5K2ItR9u
RyYlgGSb22Y3l6W+wh6Od+lMJF5WxiNId5m1QZd/p3IjMqxqwQFFCQOmuSdRpckR
tANGLq5KDkiACTa2qID2a2snYeOMEMVlEA2GcXEhNogxXLv5XU7KWn4gjieevd/5
/oQ3eUjjuI6SWZyyt+KToYxjH1hRIQjwVmk89v9LQ6TJVicq3KpvIm4Dbhy/PV05
8MYVgqvPb3ujU6s7LWud83KS1egs/k46x0FtxuI9++4Mo3NdQc7wsjJqOxqMH0kD
2ap3fwZkwhR0SmMUb23P+OD1JyIqCW8NGcXCEKdU6339ysB5A7ImlPAGWUG6mtp9
PaqI/4uMIvXPUmt3p+8X928uvxdzQtzN/FL7Eew40viroAZr4Y3U7jWbRw0qx88T
qrRGbuqxNC2EUGnZrTMRggWn6F8cU5dSe9hKJ+sU0sOvDktO/qB5pPWluLe3qTL4
G+zi2DJXX02KRzRvFWKyzQL6OmTMybc524SK4PsqqARnPIjvSCvf1f3syqM4iHOz
fhy0rb22IQIrG9usZyiDTfVf/QTUu9tOdJiNNUY7EBbgC42z0m7TEBHx9neacAJq
sc/ZDdAtlpJCB6m9MoN03YQajkV4rF+ssz7OUFn8S8kKyWDHZvd/QP8wFnMo30xg
yDne5Oatij1C4d3KuDjU5ct9IayBuQwDsJHgG+oXEhmzaVmtFNu3kAdN3ddMJ2m8
hur1QgylHnZSRUBBgdrFmcUOBc8uJnOzdM63LNzi6yIm+DUg4rphtxxf4gp1bQQ8
ckjaGXsSQY8k2c8tcJWbbu9zHUXRZUhGWWjdpAbxZy6czgCMiWg4G5sm/ivOKZXi
UNC1yuBKcwYCuB5Oz43l8U4rctNMlBovr+H/Nzy3LJl30rfh6wv2MYLhgNSauGce
ZHesKGEe/xvjhxbp6dE2N8JYQMHhe9jvPAC/LaeunA1W9muQ7CNQEuJNnvTV9WLn
WfcWck7J6NiQbVvV8VzrUPgsHI5QJ5T1bsuxk0zdXZuLc893LyNcM3iywuW5gZoS
F5/ExTMOfSTE+Xg+93Bx4YHlxfIBUr1kJq7zp6Ns56tfoTbI7orxgl1M656v29aH
+RR4i7ZXMXRg+gALpSA8Nyawt3wrrqxwScMM4h++hmox1vR3bCyKmwtKMoN+MwME
kKpSBhJBfNi8ylVskmhQMnwo+eyVl75aL3PPkLrWv72xfSkFx0hUZ/B9Y5ifHQPB
WzyFsY9aQiQ3RNLZmeFvp2i+U7kYsiXd0sDHNy4CcbywTkgPVWZCKWSEmF3jNXph
nZ7ajUV1mo52PmDSUVl2Us1tuIoooDY+jHtOEhsIy/WtYT4skFx1TfYj3vVg9zRR
msr7O8DxR6rAo7dV7JJ0dJ+sKoUuhge0cjH8Rqg5pyCN6gM9MVt/zKkfLUdwaJHh
CUkGmToSx2YTqrIBlfmxSLWBn6GJe8erV81BnSpO2AozMSn6D0EJ4vRfcGIekTvR
H7y04TfktxULUrZidndfyFcFHsGD6gDEKCyacfDOcAVlixkiYSyusXrWb0Bj+BQN
kZ2PxqYXhM0l7f8jsZ/FytKmce/YfuiyLFa9AkCDlChDKU02MpnJFxqEvMV+DHzX
ZRJGM8M8x9VDwTkfcqPaNNUps7npn3fea6me9run0aoysJR6zFu1XavYj+PbdAXE
a0+1MuIXuzsAq83Y3j+yxSV/y2iu8ST6sDDZ5sFtQFzmBSNJJB/gKkZnLkp4Twxw
JBG5WSBsrRVYTyQH6Uqem0X23oUk9TGIiJtxDKA7ut29mjJAeOtlvLzYfsmdYyzV
N0QAbKz5OfsIxaJR7wH5wjva/T+V3xz2FXJzyT4xmIsdU9k5mw8+kX/MJYAtAOgp
QgenhXeGAs417Fid6cbMCs73hBcdTvBYFMtuFSZSArJwoBSPXRQyab0Ksg7n3iYJ
TrgyCAynkXtahxvaLSwje2ZM89jFvga9/lz7IY5Mytm0DHsw/9yRc0jU0JGEbp8z
uA+EqeqTMLMZxP9kZ4gjAVHgp6TqFuSdtX7ognJyaEv4D3Nba9nsN9wawfVPswoY
4N5kv20ttiyP3DpdFpHv1WasBKeS5IoLHA975tdIHuVV838SQjwN3q2FnMP2ZTj4
XA8Tbo+C/F3ly/5G0TZ7HZYP2XOi5KsVS8fZtyvtNZh0HRdQowZ341h3CSYgvi4h
1HcoGdC7ETv7X4tI1Fr8yFfQ1f6JR5g6JRaxB/MwfBbPKFFaRYrJ6TGroVYpctEM
juO4y5KfzMTDSCrnXsKO9OWuv5YwZ5qF4W25YAQe6+ILx9XeLxUGIRHSgqYAVTcG
2/kNNi95XCW8DM+WRMajnP0eD5ZEuF3Bo83s2Sx48OAbl7BP8uYJCy28KuX99u49
VS6WUe4/iUy9jsgzcLAezUpXt5TBp5C1oBvklk0QBAHCAW1v1uf8U9R3KPgSI87o
ukzup4KBK9rS45uEGSJa0n87D8LHhhWMl/4Tv4h9n88I5lOfKOj3PT0QenFXEtVN
oygL4ziyBzT4jEbhdOy11hA09q5kUgMHrhU9WR7tbyFsKl0NbaIe87HVZOn+A1CG
ID35SofPSnd7rMwruQZOy5gXK+crzPAoooGmkn2jMlnWppg0ogdA7UnJhv2gPzjw
Gd1/i6aYRY+SjH7TLgjsbNZgnFCtWveeaQQ8E1YQSHqmcMAKWHdDtaST5SSpGXH5
7jPLaLKL4mBrAx2s1NIEq+qsBZQX9tSekf/gi07X9pG7elRge8IUnNxMMEKwf3fd
wIYeTR7uOTxpXXt3KV0UQeb8GfzvlOJ5s+4ZmZx3aIBK/DLsinBX0APi7laIk6gD
z+kGHVqlzwniP+CDE2vdZRCbw6Ycz6qXlI+nefA/0apQH9bHrvvpYwKXTuJirqlT
k2/QnhendadLVLnvokG3s3Y3lQkZxXoQvcYJRo7mQcxZvXFfnK6KtPe8j4/HMSle
okh7OpvtgNudwVO7cnpTaDL+PxbBmcmznpYUqzRNUSxqXAOAZjYe6wRLTbCmTlOU
jXc6NGcZzpRycvH+1qp1MqgY+qq2I9zglws9y22yJoqPunuhZZI2Xtkcx5bt0EGO
hTvoeA/Shz5PXQ4cxHN7Tltjx0vDjU9w3jU6mZR+GwKbCRYw9pIk4fda4YvHKXpf
LKIkygf32jJF2dEpoz3rXqKW82HjD+344ksWZayE6JyzBQBhTlUntG6IH8k6PAdV
NBA7K3jipvRPXLEdwCwHvj0/xs8wAmNHrhXKqCwiTCunQ2EAQWY6gfo+1AP/+dji
D0xL8mkHWliHO92CeUed0bjnAfM9E6pcmycym5QZMRLz8DCxErp5tIMVfJmtB7of
4MTDBw2U3XzOpOIrhTtak4MTbxIuXVzjkx1IcCrJk7yTym6z6UsAbgbiRes2kdVk
rUwRNg9fQ86RlxCprINOMcTKbSFCEHMWKzz3O8x4lCweabDTx1YJWM4deZkmXKpM
J64sIf6yZFgSaSGwtjCznQ6XpKkR68499SQtCseAVuZzRk0a15eT27HlpWhH/E3H
jDrG9+WqR32nH+ZTVuA06uz0dBrcbJ+5mQ85VJMgbWCA0UbZxfbNzqWcYijawzbP
Z7rZ8ivC0m4TY3aSPO6DHFUBr7d1iYsgt4KExTGgiKEmVTFNsKEZy03cuh7hXyrs
Ros5WDkzIOqS6ROHA/0uXF341RCeAWQDYxK0ddDkfmdS4/qsGIMYtLV3PGfKRZbN
oTL3CaC7/RRGEQCorwyB2ek+1KaaYi2crhIuqlliOPjC4Ev0cQXUcZY+IDcczOs2
rUZSQpXvVp8HinHOeA9ZvaHaeopf7aOiUkkWygODQ/NC4W96bJ5sNk8nQcJfMPMo
4eH6DL9CH6jVYpAB3DcmcvB7MjJQE6niyEjWSbz4SYCoLqAcCTpjFE/VV8LrNiJq
kr13z4+0Q3vdRBkUN1kKtVCtCaMzLruVdxdvfQ+0oB/ommoQBe9dA4MmT3KZOV4u
WevVhcxtYDQgWyHXGiuOdBzZ1Kv8doSVeOXJin4E/OBeIhmuYSOuB80ZDzYyZae2
Q2uBgh3ZO5SuzFaK4/A6jfjwFOpyM59noO7/X3vmPQjawe7ysdgRhxD1PeCanvr5
JqJ6oRQxV5OHXMCn7GdYkeFwZjMwffKYOwJYkkcqU/h5+tiGdhPfhM/bKIi448Ch
RmwJVqXeDciV8iNITkpcwyaoxEn+IqlXuujONfPqqxIfK9bJo/ykxXfj4u5SaUC7
k1ZuYEiHyQO0XO8T9jK6PhCyREU7yPyA8KA5d65P6MaWMYdfvrzDGNUGDQfW459b
qLHgBobnpDSEdktFImGqA/6yA8lDvG/avfajn1q8z4lWiZ2FfAoZ4OrJR+kT/5G9
cdBfMWGIFyva/lNTvtAsy6IZTYfwNcseeZU2u3rDaPs11j6sU0bNMjXGtUzwagsx
03I/dcsV+tozomTek6qSkP+O0OtEfCnpG5sAbaVa7X0baJjN3Ds9U1f3CbQMGYoC
tERb2MrPrTGc56KhqVRd95NG8BgGrjD1QLiruhpA9WHPatGn7EeAPNF81tHt3Ulw
Gd2VYH/T5kpFpgarEh1rhswjZnkFTQCkXTAGqAfVzZgOziJrprWrW7lLjJLKTv/4
60JQu9S2jNaCRKsZqx10gm/GKuMXgFPrp8xQFSppW0n4KqhkTOd4AQDfO0uJE0r2
hAP61nyqNkVPO/jt+saULG3lJMD7nvUu+CQaV0WmT1eYYDpmIGg9UKYLgkqitRiZ
f37Fi7EDxhs2JwfidGlVCArZYj7JbDa2SNj/rygbxGt6tbxNg/mig6xJXHEllxFY
MdW/KqOIEnUFykXQP48xsyvWYOtuhiPNovZ9rY9WwgV1InQ6DaoxBGNEzEvDVsV8
FjJvNdvC1h/hPnebx714J0IxJXZ5eKYI2xW9aNLMfDqPz0BLUTsYdYmFbEUKPRLA
ffBl3bhssKND2Xjp9tcAnRFzPqFJCHPVmcl1QdQ6COLzxSwJWaiRHrpqxBErLKY5
yTEVKSW6JU6VY1zOYPuFY6uu6hDJlKUdMS81DO96Enb5EKCS1rJpGAifZ1V0yG08
+Wi2sAmebN0r7XcuQffn2rl7ecBDwjDYKxkJiW96qCZBS3d+i9Dj/KOL6ovQbX7d
6BhDbD/cRL6osEBPdzv39Mf2edbFKBK1j3ZhKCxj0yAUWRgTJgnJ2FApuGEgtxUg
IkP7rS/JKZYpp8+xwXwcCSJUSGpWxRWL+PNejqllZzlgkJChm0NxKOZnRHa9WaPH
NFL2CrDC+ywqzO+1ZlQDEJaCII4BOxpTwyRDOGr/kR2/T+bcuV9/OXF5E7Czbvsg
SJBg6dCGpiHiOKOLkr1CteR/5Y0Qn53IMR0v8m9GoKhEu+n5GfCHFPOrzKBi4+6i
ULpyampFl0kd+UbYXWr6epc3pKDX7nWqmPmvwrwoJeQ3lqg1awQsuQAJz3yi4UkR
b+DCZXEsm8W2odhuAILPSxAlbmYIYHrLTJvAnNA/zrHG4/3yxIiEtY9Eh5aK1gkY
g0joe2zOOQsVzh8oU9DwMz0tSlls+kRNKUoSL2McIl8ZwdBMmU6kJcu7H0SmIHCq
YOBsb7ShGTTGHxqJJMarxPvlfg63NJd60MPEOk8y3g52KTDsvxIRzlcyQoOpU2NT
1Vn6UKRUrWTlC5M2S2NCD33mQTuxJ6jTp4QZqSaq1HYUbbnYQORyCllHhkHYnzcQ
9Kp/hes2VHJ2qdxuHlbyYLuzp6XSVfk6e63qnRAMRtVcuemvV4R1Vvzq4Y2nF5/i
SA8LJacUwqzLNKfeGi7tmbRgzfZbss5vWR1enU2qZgFy3XXc4TciSHX9N4qgG7Po
s6xEEsBKR56ZFw/pmRm9qsAVhdGLtIs4t8Dq7Z7ZS5lMrDaHkzYnXi3Esl0CmpTD
mkEBssBjcVgK01UM55xUbez1RoDSlqznfj4CG4PERcj7m7G2q5Wu8iTB9MzGKGbv
Cwe86Ab4N4nzozvb4L0lcSgOJG4c6hPX8SQhYtJRBVdvSk0QA4g5i+ydDGjKhqXF
egw+pp48nab/7e1fpEmatmSHN/v78nBfrCXBeobzc+mJF79JWbGgIBQzQaStwYtH
qe0mobOuIPc7gu771MvCMUlwSVZiubuAmh+JiljUSrGR0UIgtpXAKn/w5/9vXcL5
eUimdBvTYnSwrW4zIkHhyaze3qwxyfmeW4IgQWhndhFxivv7UgDdaiINTGF/eLXs
W07BFzsV/l23nqRRAh9f+SZuT7DKknW5wew8cPV6huYnnmrutGAMeXWLzwzY4lNr
yuFJGIAz+C5n6hYj94fdaC7u8cldbRpEWEGtf3B8wmwxj0ctxw3BicWDYXzhZR72
EgeazXsP7TsfNc4f1kXR984CPtAc5fYwznyixEwUCQKtIHBHMhSkGKAXgbJF8tY+
KDWq9tWDYvlprwadEkq7anC+MESUjB2s5Q5s/Je9sTmZC11AGM3zw1oRaQDMGjOQ
w/181wDy/mI1LGS6nuVx5Te3BRfANQz+7UVpug3Ta74kv56Tj0vnWScxKCSstSMf
f/+7Pnc0PaAnxA9Wl1ecjMmmsvlwNXhR1np5f/HI8iDlxUBnZI+zCrvUq98IO4q7
gEI9PwRlaeKy5FXVrMQoQynNfOXtwn3hmSmjS3pF8+fR0m5dtV1/8Hw1tjKUvENS
y/QUJN7kGPjOYg3uQm8RmhC4XReG0ofx4PkAOgRG8a1jOLYxnm791stoE1YOttEC
Weyek21B7pUt20+/Cs5iOOsVXKyYbtSDg0J8Bu1hcwNp1ypy3Yu1b/GgV3Xu4y4Y
QHb1EzUUu+tjvIwCTJDl8OoMqJybC+8D4upifSm+8pnI2zliFB8TFQss4weImeDF
kC3XTWajwv8Wms7pBv1NTBt5CJeZJ0JnaraeZmZc8pQIRloxVvh+hy5NGtYlr2Dl
WP0EfksJe8TKesKcsPllhWMSM+kehpOuzft/pePKiEqSC3FIRlMU1f7K05+EMK5l
ym959nyof0Nqdgr8qxZLnYZw/lkV96+qA3yjHeFQKkwEPyrfWIhiBbe1Gj5a2V/C
FRSQE6A5tP/A88ZPIiqQFG2LbV+C3wPI8/jT7omkkYrQitkKxUyu3fSIWLtWGD6T
w8l34ODUmFMlEiOhr5nUgw2s4MezZCNs7brg8Fyn3o9RFWNY8i8f8UKa9SRfyR9P
fuGpjeyhRjJ0eK8Ct/OHumdZuq2mMaXRkyMPBN+Ezfa02KJhZLG3QpAgqLWyWLAw
p+Mc4sbDjcgg5kT1cPlphwUr5gbqsdNkLHesU1NUlHoFH3lolW5t+/6tlI737BOk
Vi+fPFibrLD3SLZ65oyQVi5zvDAlT81RAuu3+xkKjtFvlStGIBp1uSoO/Zl9yg7f
J45iw3/YsPDQ7AEvmWpVfAaihL1UHbIVnOrg/LPGGY9DDLiqjnuzW15lCEtyzMPQ
wWjr344vSYUy4UBgoV9J8FvhzhiZRTgqM6cxrcQ/YbWB+DxkN7xSlszR69Y12yfa
cL1eS0lym5BXxDBiN88Id6qcGJmEeWPQSN64uqt1AjGauO0W7O+MB7rkNJMzoVbu
eB8jV2ROpElJHWO0hXsKoa6s2QM7TTtVO+JMZQrdLB14hABNenZXwNI3kV2H+48r
VfQK4wA2RrWXttgR17+k3jatq1No9a7jeQIUFf1yddwuQnvchi7TdQXf0gH41M/e
+VRkYwd2JNoxPVmB4yaHwJjmDOBKFCEo/MNb+p1wsAeJ/eDdDDQ2KwlGy7c+B0u/
xGEdtxPtNTztTCOR1mu0JDywWPEzj0IEh8SAdCMB82iVaB0AWB+L0pJ3yYPrJ0RN
VVwETGZljDST5l4UOt5ks6qkSUlpO63tfcUyJtIFIvgaeOCQsYLtfwJx6SpAtC4C
r3d6GU5qwhYIkZ1YjOyGSD3g76bM92iMQ06UYqDG2/NwblGgSDKGwlMU8bhW2XLJ
lPpCnWeS6Fc7TkMzF9RamCPisAk3W9J6zcLNUbv1PKMkYHry/q4N5QoZU+NAiY6x
/tabe2fYdAiY12ms/2HLydSB22HTETtrJ9zAG5mMbz3bMHuR1sxIu8Vc3LDPAsRO
Be+kamhBcDAV16+5VQeauhh3S6Ndso3S5UkzmXxtk/JuhWTvL0AwjLMsF8HsZAHM
aGdwKLsmlqDckfz2yP6IOxw7kry84M0WrmxbtOPk9MACVgUp/97CWVnBb3MlM/er
I4iFCOL0xFT/A9yKJeKnlp9RbudBhJXDvqDyTSDPBL7m+KnIJtxw+93r2h8DM/sm
rkJ2hCu5uggPBm1BHwCd63/Sj5uyfTXDoBcT8GaIQSekOETS8cH0/jKNodCSAMF3
OcdtvCuPKKuxfoM7IUVgmeASHKvzPn77cUf0T0qRTX99FLWXRWRp3MXdsc5fFKM1
JV7OTGE9Whi2AxPVYn7juW8KSp06XeU8J4NjLuM6rtnPINih+y0q16uUxTe1nt+u
o3nAlG8os2FpNYihyYe3uNjPfbXo2Qb7w9vD0LviGQj9F8Juu9mBr9tVYnUkEBT4
DEweL4Svoc5rOH64SQ6Bf4PElJwUbwb+Fbx/AqnzulURzSInOdkF/7ceGF0GF8Ed
l8Squzk8vhJJuu1SAizFYFL2m/ueINlHCNZDtAA9Q31ZloOgCqlGiUUGl1WTIqOP
cBLZHc5eRrh1WsLC31Yh9qnpELnHoCnomNqfYcLN2r0ue/lIZT8eM831UNNsCzLx
VVwLE3GA1FQeo3r2KRYEWb8fUa/KBQE4zWTOdnsjvBy/IRxe1DqZdAMUJKQvyZrc
7km/xaQR/XQp9ZhHVG0RdrmgpfcjkmWzUGAafMzTR3WisyMFb7zm0KOv5UwIs066
jQJ59uapDCHTIH4XEVtpS0Xs1thupXAALZ9AnmoSsgsRY8wFV8nPqwoGrgl9C7lV
tUaTA6ZA8lh5/QR5rG7SdsnCy536sw+dqGInKMoyKFBxHikAf7eQnvB4vvsEw7eO
7raZp2hrqc7ZrifrrpWSVoOq0G3Aw0PujEWH+98KZt+WYXJIBQQcQsSfhUdqZ4xP
SOhC/jF3u0+hEuZNQ67OfLTp7Ht2p60tyKCGfQdpWMMLWOPe4bLYRV5T0ii8CgKk
8/ZVk4lqUt37Gf5Iltp0vA1KZZAMV3+UigoOjD60is3ttDCUi3QsRluYHyDBaKq6
hOn84ZFHgnPTuFRny8B26PTjGzrjAU1HHQXtnbZVM723mtiwnbp+2Jzlf0VSgJcg
mpB2SEoKD4I+IGldHRjUjg3oAsuftv2Z5ODTtPhLj8gGX1SG7dLf+eJ2yzD4j1ge
Q5xWuyWvlolsuuAEyFQePgAMk1uUnEII9oVq3DJ8WxvZbyHvrF+iq5C3X8+khFeM
4O+AXXceMo8pLPLVqYS/0cfkgG9fmwO/+s1rIHeeTXtOrnykDEAM5dP1ECmB099z
DzoOU7zjxw6ak5N5QdVpr7xZ0G16rt9orH4pLfAF03Dsv/vdNajbw0a+xXposYGP
nyVL+IvPKCVmrq/cqQcMGEWG9UJzT54d+DjITz6HFtDg2f8YvqLLnDN4fgAoqqxH
yqPSCyQbyOdEfMy568Hx2nMq96bY2qkg+K3UqPozqkQOkTLsGmMsouEjvhNbqcBb
vTVcataW14RG5QdsePn5v/6esRgBE068pitBLJrQmCtZ8zX8ZvPjsafFeAZt5zqP
0VsNqSZ55wf1rbdZzwC4nljYnFhE/e1KVC/GnwzX5Bh9/FezgFCkQ11ZGsY60P63
e4B+3b5xg2L+o9yh/YE6S/+hdl+sV9f3WtaJA80zbNXB7JVs6d5EdthemsBFK8c4
BXa66aEWSbPD1ud3gOixYFsClaSzXOov5zDKmpWPf6BjPj+4vjW25VsThOlIcA/r
RBKgTp8mL6OyY0R2d8XxPgCMZXi6vl7pU5oMVE5RADnqpiAj2Dcf0FXaXfwqdXJv
qZs/ITiaQUiaw9c7aEeyH1rWRFR9oZmQdENfaTq5vrHVTqSAEYfk6gImJ6QmMBMd
en4A+cVlJcJBi761em7YgDZkkvvIbP8bHzHjKGRZaUAj+73Sw/qvuoWMjPPOGLfb
jC7p86uxY0Ua4c90dDYTUe4CK4pLa4PS0SIejjLYOmHRxz3POBzFNzhPfcrONz5S
te2oo9mrFldQI4zFchix32O8a1ndqlQ9A1SnTZUXrJYADYgzjPuqJvCP5ajaEzun
FXuEzDUmU71kN0KnaPug/dqqqdiGI+1ZXqkwbEqGSwO1h0+CjPw4LSHQBQB3STqV
yaGcLBOBCgRrPucM5kUk2oP/rIo8ot/2rCzD0jbzGNfVt/dHN+vHgRyw+dc0dsHQ
PdmRMWaFKxiXmb03QC6CdesmbeewYqyle3Wi0m1eNglMHwzN5aadRtpitu5V1LEU
KZI7OSrOp54R0Vz7FoCRDvD/1XJd8ZE/nKQO081X1PtF45tG9x+9sVjm4/Aix1Lp
2D4kEl1lufmGHgsKwRNAepP+EK8FWpoqVY/esz3vZRSMwk2O32J1t+sinE4DzFid
tQCwV8TrI2Xm0wuELhRKF3ixGJzlcOGrqsZKWGIi4oOi1vZBaMP7Km3qdvUmHqp7
uZrapA3RqUmjRbJqDPVMBUk46LZOXWYBID7nng8LflKOI3mx9JE1e/4i89qVS9xS
wOUtsl9sQzrS/uKURDcmwLzZDlLalDhoTAIS7BMJBJdFalAEC213u6oJtrB+LYKL
8s4cZj3HvNS4dw7nWGlumbSpGHUFTAfI4FyjpBra6l1qZk0Oduh6VJ8vlXNN8QKK
eeY1hQIx3Lpwz6xvRSVjCD5ZNGQjayLNAGTMYJWROJEKAZREfb6GgQAPy8/inmpD
XpbvlOyqOk/g2BlUENXgfcG8Vjqbm8sWqcqc/WGkCgHEiDeV5eUZu5xglqCL8+vE
5x3waJv2lnnW/dHDnQKs1kQKT4LBMh6zHAJYAz2BQmNul7ozZOqSc19hyTioN+lM
BwIYKgQCx2DtGkvwgu/oTw7hLCicLthgpdRCaXlg7E3XFvl4mj8NLAzpSdLve/T3
07rvXzOeuh6cESDhXSipOpyhtNkow1r6sf6d9Wwcsp7YgfJemRspy8sYYq8uN9xC
XBA0cEP3XlXJhZtLxHtXPT1Oq25BzDzIskCgustgkC0dnYd+wvNshWTLRul2Ib0o
YgZ8nRMTUR7LawC9S1WaOcopydMUykMHMualdN9vwl+5jF+lQ0SODpawVRK8/5ey
xkdYpUqgB23O7Pap0eSYbK8OSyaPJ9zqsCBh5APJW/vrqDVNv4DdJKxZfg1hegd8
3ACI/OVEnO3bjt36vVYuIjfcN1V3RG4uQqR/LJwKopEa1OJZxaFDyiuxI9l/K2K3
FHnkRThtsxv/75guAxFUySlU5a/4z8hjd3J71cL82vKILhJLBHr9viqnWNfjm2a0
tg+O92jthiNZn++F576u0MA4sWIZLBLry90jgG/x2cA3iZ1i3mDEqym2+wG4fA+S
NitDXI7C8vsA7ZSQSoFvfQgPfFR2zO83oRA4CvOz5HRSCX5gea0VrbYSTRFtSibY
lA24g8P+7PIJ/S+taXNBpKGDIZN/sAURBs2oWMrGvTMxC5bQiP7X6ERs9Vh3tWPw
71Fd0a6r9WSgHfJZ1w+yard9vH/jEBJy2oDNxQwGKPwdXDm2Ie3d0Iw+zT8FDDne
tPhLDDSp393gjkEHXkrK8HoQjWEZQSmczn/zEEs8zd8rQHjWaP9KQ+BizN4MQveN
6lHqIQHuFEpPKkDZ2L/0TrjnR9deP7XWiqoLMzvsWCXzqJt8ETeLtt5O0eal0cfx
FA6IDnH9glzPKJDkTnHQmsRHyij6BuMyLCSxvgqgdz2q2rwRr3Uqml3eRP2Xauog
KT7HKfklH7V/Y7s77hbcfZaIA10EqYZs7PmtbCZsWfwFhUXO67tb+jAlblTyFjma
DEGMQUj95WpMrVjtgcgUiSxMsVYALv74GVDwxdZcMfoxp8zI7K22NazlG31DzZ/i
EVKbbjffRZF14apGFbL3Rrs6fGcrbIXBT6HmzvBkxDoMC27eZnZPHgQveg0rdrMH
hzNd4Dnv8D5s12r4KQdbVjllw+wBzvDnAmZuRaseEtLPxyo98Ou/17jbmHivsX4c
4DUumOozbSy2u8Dd53nrpEPoJtTp7E9QYb2Ic4rFc4En4ZZud0XNBoWeDyZ/gEPY
Q33ZZQlxzNxOihl/71AIBjXbvDEltI6539ovropZ5HC5jsqRMcEsT5TlnPwNnff8
Pb/RrCGuYw/RDf9DKx7plozr7L9ZAtlJQ9BIEcZCpMxlwLQRaeiRYQSyhPaU0Kmx
mRF2dWER+p+Qp8hJLSsYwbEL6KKlY+1dVrOV+g99W+9f6tGfYv/9uVasd2qFKz6F
+7i4t2Y14VQMR8wswctGOp8aJHJxvohxX+ndxCzusMnFs27jxqySbmoPfwkAv/hc
pvB7QECsYpoJ1FGZE6P4NgK8iI+VcS1EVPhRgm8SPwZcj3k2caKRNjq7G4gemSmI
pi841p08NxIM7TBztiLBaQ0Lq7T8yzpb/0DaL9+Ftaa9kA9v69SK3zKum9aq8L0E
fmCmWrYnBcEC2hAMcR4GRW1Qorsp7Si5Io/vijHGR6HoDTFeFeRHRDbN5Dp19p6R
FsGCFDROEXLIVWlxtz45qeREpgbxk99eO/3UAq2JGrSa+/Z+pMpXJRvzfA1c0y6J
kpISp7gnFb0qV/ULLU/u0nP2skJJWBlAZXMnNFUT2LjSWYluc6XAuZajsKJRopMP
7oOuZbqqhB7/5q140D5mWoJLevR3+k04nbVqS7Zhd3CgIhcJD5UinQg0Oi080sgv
9OKJ1gPLKLtPjjmyeM/5EQIpYl5OeQifzoy+NgQ9CRf9fxsTw0naUnIFmsWggjoy
Nhyb5bFbMeEwHB6YmZW8A7njPJfZKjtm9NuCuVTkhPO9EWEjiaosdtsjwRuse9KX
+AKG5SwZ2KmEUe4dEDn5W+9iO4zn+dS7OUlKJEbqQunZqfR2NCyveVuJsyV0m0w0
ujA3SgF1HCYyf44ncuVZF4dDKWJ+XgwAdDQ/zlPGE6vIO7D61tQcU0vLF9vPDL+t
lTEXMWCptzZyQBkbSy3MtsCmbvGMTE1q9KGfPJLWthoPJ70Aoa6fPeWk2BoLl+Cy
6Z0W98e1KFB63dPoK+D1zs6p2lbzEr4hTpN4CnpBjzdMckRFi4T+BP5SZw036K+m
nSnZ/gytCaDeNTp4HOQsnDa+k9Tje5Ysxa4ogJp0AV8/lPewL+EhUdfsBQPf2xZf
Yms1OWXdd6EW+ClS+e3pKWyDUvj3CBH3SSCUQ4jpB8mqHS7Q/UFxcrDvVhNjl+ur
M7+98P/3XbMAV2NvJ5X6cv6OVLWmiGPWgGoAV1eVz5e24ZHMjMs2w4GBDMKY/+MA
nxl20YEy2utSnPSQGWTOjgModYv88w9/nD46E5voyebYKzXV2VpV2PzSPPoUlRcb
6hM0v7a4UqN74sEBYCRthfwVpNAUrpWtDM5NlusRFxeteAWrQj/8pi2e1jvxVbim
5HIgThNWX9OwjmPVaWOEgo2RTIh4rzhGrnEE17oGGIK16qWnilpER9GIWTQCD0nn
u1wSbTIZmP8ZCEJOWsWVcYRvQ/duDzuWIiNx3j12SYMJVzZt/WDZshYu0yd0ho4y
/xzpA9dPsWVUrF+qXAo4z8hGl0l7OM587Is1fcALvyeO5dd75YawZNsqEJiPwloc
ITaJxHCuSLsJ7kjTnGmPUMum5uJlGr91/VjRVR9A9wN9zr0aWkOEZEW70dBKsdhq
FI4TDpvqXH/NOZ+L5OF9LyX/zOvIw8mGOJIjxpognWfima0+bYa1p4BboNrEbauE
GKHH+Av3YVVjafJni4Ck8pL6PBT35wlR2Zn6Tulr350Fg6uRvcTXwUPQtWaE4mjQ
oUU+On0bGUEXbbWNLplgW+Q0yiKZFxQokfi7D6iOlns2/PKm9xXpdFnZ0Rz8QHSg
b3DCTxsMm3Mvcs8wMFe0WIDcj86gmWPnoHdqH/c3JY3GVJUJU2i1JnmKMGUuncA8
GbpYhArCv38cM5uRwkmJ0vmi8wtuO7RVk5BnXsHZIV5ygj13D7MhvfX4UlONFZjR
HgmaWqnFg0I6tETe/5g6bZH2KPUoiSuyInjtxKjhdoNIabSJpYtnAYh6ok7e10a4
tQ2sxuVhqfgjLeYMJtA9X1iTt0GbEgk78iMCa2CH0wNrq4iZ8ACORQa5IsY+d/q0
/csIorRYJ/ncjgAdAloAkNzZBfq7SOgHMOQUbSrcxBZ+j8Yljh2PZ3GsJihLgtdg
xKmvLG9kcFeBUjuLMgcKZxcmLf1uQU1UBFIjyiK3sbhwlxxtdCpeDkBI5MyWfoKU
/QkGn2y/BUwiadciwXQPnpruV40XQw7/ql9v/TwFlXndyiqvEKSqDOndnLNEQpQ4
ozVKsuO/f0I3gZm3Oayd92RMhqrIbk0Ewok11j+aAZYUJM6nBmYl7Bs75e3y6M52
vTPYNYefmsv0DHA4XZRyxAVDiDkQyuKUtONTaISx9Er6vz7sJ2VS6NlhixodnkMb
K1MpmruTEyobfbR0UGlB2rkRhOrq9O2o1KQEONPDY3EhVlHNubq0A8tJSuGkCRlc
LyjChIMNvrYag11FI17V8FtAikaxQ6ABkoEaVOMX6lJQSIovdy2Xl/mhhyx8XXnI
YUGllgGo3v8AzqalUp2YBuEa6gIGU5MIlwqcJ3woAvRc57yQ2CCYOk6Rfx1IwEt/
izaEMOIWfk2UzyqZm3hA//KneT2nxBVRKwYAta1Q2FqeDq4my7hzJrgMVVM7GqTz
Ez2m12D/jMSeZsjebliY7F1NBcqwe3wafZrPwOMPfN8/L6FAQJJ2xF9XbiCkL11C
ZoQqlC8x7d3sCUrsHWpYwtKoqkV0H67ojOahHU5ZmI3YxdkOeOVKBuMJurSg5uEU
c30k7xtukFxNEywZm2KYOL9m/FMOMzcAuSpGlJGgP1SPT0VcRmuDNoes4HPHyf30
nZPQXft/133XfKnEcWfFnw720tjIhFLGOQ0XwNAj68X/N2VDJV9aLPlB8T5o0538
zb0GFrbN9M85RpdN/daJaJZP07dvu6+Atnrhco5H5G0ZoZpEHWLaJfHDQfG780y3
QW5kYXh3c1QkKumv1MiqIOn5hIKcexCW6luMPH3gLpj3wGeEHRV0asNFG/ue7A5o
1zpmgCkw+zeWvQfPFWcDk9fpwny2N7XFjeYTS9mKTh16wODejjV2NrF57GNjB/D6
+0vIFcg6uv2lfsHfjV+JK9QIE6N3tHS56a6/CbBQXAaSsxdX6ttuz5zV6Qbk/k7K
QFZ/n3BMHBzF8/xf2OXtNmQrO7L6PVjr+G/P942lgC5KByN6XAatyiFUG2wn7EPD
eomf9SVmt8HCBr+ecixXzen/lxyuZYMfY7urO9++Fmsc+gV4C26iytG0i+yF5pRS
EnyvX6k7RU9HY6/w3wJ0xAQuUnIzOyDNuT5fGypMLDcP7uFTqsO0x/fKzlNMdd5i
v1NKxu2wxiiYPI/bz4NwVFckqQ5g6B/6esQuUJuIrMjNFwrl6I8EARyVz59oELar
BeY6O/hjLMVIS9r6Jn+Lz+1C2HCd0YHTr/m5ZF1y7J5dqJ/4/vCr2ZAr92DE8bXB
X+k9DknpVuRL/mOhbUnfRcVL7afXrxyE+qIROm2Gaxf9cbhtfkBVyPulFR2zpoSf
nwHFR+H9ClnqQDNv9kYxh1FqZqMysDXmCLCHSVXWH2EB6VhB/nf2JLyAMvhVslHa
hb8m62FNRxf8i+6wOh8zPTl4dap9KKmNDmDOP0G3W8fJAXpr95L4OZ/sajz8Z6dx
mxQ0BJRIziDys2b5P4dsSwrciGL5wCf7ARI7nBCjBD1F1hqNqJi+YcGysbXfCCns
msdUa06qllZGSDbjlGOfXE3MwD1PnTExBPF9R0Sv4BzoTJC6TbrKoKxR3RQhk3FM
0JVZGCBclX5n7edtvS36VrmasbCeWleg6qgci/trM9PHkWHCl6lSzerugTnyQXpm
Ff4Rx2ey+Niz97G2l3k+Qv4C7PNb2/ao5kT0D08KpsD+XjpQnuvmawUEvGxE9Ilw
pH33vkc4ndDHu+DJED0YkPlh5zea0x9XrlB5Pt/uS1cLnMgEkmMenWSXvCHmvYvU
CK04KF90eyNIFsIUDQzdsom3bbvTCal8hFmqWVMPN+/gICrmMVs9mvmPgbgmErcj
wWZig/NalWzCcbXgLIqtAKiyl8iYrDE5MEMySdhO/W5TwqWd0kqTF1NAs2Wr5JcX
KF2VosREn260Ml39BkxcIZvW49PQOxsrb0efcDGMH6OOQjYdsMXwxaTMT12Dy1cV
ZUo/16eKmUj+sRCVugwPbTrf+EaQQ5gguqMXEAr1ro3MkdU8wpLgLM9GosEETsd6
mMLHS8I0OrpkQwtEsDH4rSg16E+q2NrPtDLLwOV+d2UKgD8z4qVxBA976lqZCfHT
ZsHwBse3122RMPHqDH31SWAArPhCzv83z+4TNRetCNMokg96HHOcGdw2ADYyCb1J
AuXsj4aSiRmMMPERctp8vrO5UQ+PG02r8tbQjhVCkA7k1kd9tNQV5RZpdcDNS42L
eeqFcyC3LCR/J3Z5eacTJxPQ/8atDwyTpj2Q8lL5qrxEQvL5qTzbHEUEVSaVA5eM
TnZrLrfeQF3BxvDHyRrnIeTorSuOW0mPHaX8atjVS2Vsd4MwM1pkeYxV0JzPFslD
teyROyN3FtxnbW0bxhHQWD6nONlkw/DaNUlA6lvXs99TNRHb/9kwajpLvyQOf/Oy
SeTzgCq+2de7qVtoIaZY2s49SwqLc59irw6H1H66CKOjsTrNMM9iaEL8+SBgXrFH
KEfzf6cNndYyISodl5VbtvxlP8seb36AOCoBCktynafFxa8iSp33TjuS7a3mG6sO
ddvDMGoPcdz80BIWChbzQEn7apIRcQWITv0PAqMPZuWFujOsn3UodhfKJitrV74R
1Dt/lOyNMd+8O01MUcnhqpJlFfAr52ev21fIipCBkp9sIa5UiSFYi9vilP+FFp3y
swZDRTxQKbBFDmo3Y7xhwS3zKERMSm2lFmXJ67MQOiTlXKWMlExkwfH3h9e+opeN
5sSclJ9ZmTAtoRc9+znKCt88Bx3pDMwpEkIRGKb2Cb0HQjS2YumgT06LcNIVLvfc
wXJ7Pt8LAmTtGEdH5d2CarrAjfop81APnTilyTv4fTiw4Zmp65QnPrBIN+dwQSvY
7IiquS0jg65wQW5AXsSG6+tCVsW9ogI4M+EV++JpZjQe5MPKlIE7+RM6df3IoilQ
MjFAfYx66GE4WfwFqsYmHQpaMTRqlo2bBAg4a9pcW4i0owohuak3L0m7bm+kGAMR
M9DmlYyPRCZ2BW9Bq5DRmqb6kW4vaCIQaAY+fgvPfcc5AALeRG0r/mArUROkzD9f
P11hK75z7CCzv3IiuiSusFw8mZ75S0QZHvxUFq30ivy2zfQ1WNCsg4bWfmhLxeV7
Zwf4zWiiX4aUY9stZJROpWTDDhgjBD8wa9ZUbdZ5a3d+7Ua+31/7wFkHipexoeqI
XGTET6kWVhb+/16XzpX5Kfol+0uMwGk2F/BpVZJPEtwFYRtmdaAg2omecAxxKJFQ
5sa0Lgw6nNP/IFpQIYFbQlpYhi/uDfWwBfVwPcCU7s7BLlF4PaM7xUJmf7LwlhMg
SvVKtHj+l96rd7Hj3OkdDoUvDdtHENJy0sh+Pjjo2XiIZ53fEQ74iZTX7d2bfVBr
SgB6bx/YqjGaruq4FXSaoq8zEuDVcpnm6ocUonT3nAHuU2c/o1udNi0F2+Lm1gzf
kVXf5iOo4g5I1VJspb4Wh+1MbwkqlWHn/p3KksptT7bIPlXhCwygTKlpjIuYLzF7
yml1mSoSMOS6RCWuHDT3kK/yHKrnNS905rekVQUl6ogxSEjxET1rhC3yS5MiKqYq
1RpPRX/ElJ+U+s+6BQqL1oYrGmQr5VAjCnzWfk1RDvAWcsLMGx+/4tAzbS7yGFIL
DeI4RMDeCiu2odbIF5E/OcH3PSosQxdmqnQUXtjVQOltuCkOzQdtSJAsZxeJNOFG
Y5sSiUqEJIMFg+iyMzpq7f/ETQrzsYOA5UKyYPOUIT/FeXNNXXTfDRLDi64vPz3e
eDRds/4fqobopyorOo0grkA7ZYNx3F9dRrMbGk1x1BnXx8v5ByHjAYzK5tJRPxGe
0EuqFcsCjlqQ9sTKEZwzSVIQWZtC7rqZ3UZ2BP788Ch5SfcC3NsjKjBRHk06Y7fc
mJVeQZgGcCIirSkq3tDUTW89L4OpNAgAYaBSXP1EyVI3MZJrTJ+nRwUSSaSEG308
REo9Bm4oJ9G8vpILTj6wzaAvo+uqJQ55uErE7C0ab5JSssCI9QfSHF0OC4KDwzHv
fnF0RAcAGvNZVzI7/pcYbZ1XnqtQOLsW9VzaF4Bm+88Ep6CsoGJSugO0NmJjvTHX
V7TUcmasI0l3OcKgaZ5lviH7JeTyL5Uw7Oqp1FHGkh4vKhBe4c/hDucvz22sgmBf
ENpmJ+BrIl7WTyTl0ENucD2McAPR7MIRFrsuHFQcYe/vHspuMYKCX8mmXicwlAMa
JqofpkX2Iex3DcBSBayQYUyHUCuD0I5FNaT/hg9cZQiFAGkt7RKByuyQaDkh9iCJ
6klsgjtUSKe3gt7kCXjbG7RWID5kQRz6IvqAH1xmO5N4pMyU7TILsehQoi17jWZj
5OzPLxhKCQ/DXXWTU3QtvWYIdNgIWIiHOKvvWmcK0BdzeqoPDl9L97j+IDQkc2EB
Sv20AiehRNs/zBR3grgj6CMWhWqYZ7RTXzy3SxoOOT38V3eTXsqNGwfPvPak7n8J
h7yAhK3xv+In2Dvnv3nBWxCn+5q9Oo5exnpVrvcq9m4bHVceV0iouD9leCDFoRLE
MsrRQohL2hs3vfqt0+KXhfNVGpJOfY9KFmGiukL41pq1tT+sCl1y7i39AzDyaeK+
LNiXJyEd19hc0uOGVPuBc2d1S31qcjLRUwsLQPBF0gC2fY5a2PfPryXw4/iLG/aM
CWyFHLPCYO2WL0OOwigFWeB10oxamBOOP/TdYqOUfLyiUGkdMGvSQ5Bhf7NT4xbo
pofKHCpJAhdaImYHSKsjPgp+lLttY705P7IGXf3kdtFU0arSIjvhgLvKJcOY2+zc
A8othult69j+Ktu8LJXok4d3Wpm/5uv2ROnbHmuYgQRmEV5BAlhM50R1KZjsuNX1
dIAgDtOILPWO2SImGJsbhOliU/j37PFyhYAawx+5fK2kLUJjSM6i7y6k5o3vtGOF
tc06eS2MwBH6DvcoZyvxuyNJzl/pkeT6upgEYZbR//Ro2aFmd7z1RwEQ4BycD7Gk
fZ3DJhdbOtqtN60JJ8rkc1UISYSCiSBUZB+uOW+10CPjoqdt/+8mpC1TKJC9kmmZ
F9bPfVAiOGDFShsi+Rpq/CB55NXR3mdejrR/6ZeHEpGhcBnSJ40cgkCFCnKJg7ii
oZ0Q8xxd5fjXso/ufUSgxdMn0MIs/iZcO76zxR5o1AefrkgXnDk1vQBwiXxRRY9G
1GclV5ia2rPr/yV2lEr0zjSvY4PUalTxS7mtPFISJ05gPAzFBzuX3Mxha/FXpnk0
SQuZcTxtBhxvZdMgSDX/sZMpX+kiSaPKLxJi33piH9/pVQ4vcudnXNqaXqAi623q
9EqI1onOVprrMqpuAPVi2TyL0cWxF1DM5TyCFLa+7xbEFRzGvZYPOc2fW85W579G
o2SmtVtqCwVXoZD80m2FSfcFGm/oBYela6iTsam2ELxJldiO8w/Dp2JGGKAzyvaR
bcR2izjcbvOJs9Pz7BKn6msSrP1PsR2nan/Eb/6lB4lVEbJHOII/M2UJTXwE14ck
9Mhnq81uJaBz4EQ8fdiCwIWVEHRXGXl7HpAcmIdTqAlZ8JQbh1YExrYS4QOF6Wx0
lhRiMGOnGiTaq3GfFbogOD2N7HimgYFCW/woaqcc0XdRJpUWITuBUJpGpOQEfA5N
uOasyA/9nnRLYPd7q4GpBGLOg0t2qmR7rGqou2jaa/GWs41THX8BJeLokUmgcXMa
QAzHpsKeypNgq2LAg7PJn7Y85xubTQGvsYxGdDt0miTBYcMkw1HBKewes1EnLJlg
1FqF3Idt2czQr/jCpz6Kb+Wq7xVzGqmZy1alkjrww0/ya102BKBHLX8y65GJGjM9
2yi5GtvUoqaUx5XwbVFBP1a49/fVGTzPsUWcdaDKa01m4MBlD//dn7QjdA8QVS1j
S3Abft83s9JBFibPONDIf0chc8SC4YeOdu3jOqTVlvD7U/at0pQzrNLM6pQVrc5F
VmsAA0dYIZulvdg/fLMkrqTz8pBWsx8k9KGqwQEyz6T+FMsTcmE2mep6L/zW2p1q
VR6X3yqfRCIHr9x/Si6vw8IYgbZDacsHHGORueYRYas7foA3Gp6RTybDiAQreBg5
SWTbk+VPMCoBx2NMelpTex+vsItVMIBypRIAfEevmq5lXwBuGW8FCpX7fYJQtYy6
S8LTed+kJvuI/Fnw+05ws4HDX0uYHFFxK6eMLMYrbBD5btoL8e5w1VzT3W0jd0gP
EkPzWjno2NLVV3+mC1oDMkMv/ggCJ0IXJRkEpXb/ciHo0ajY/x2IBhylYKetY4Bq
nBnJKKJmcyrnLsu44P+tCenL8p6ufIUv3VfR1pTKdoQTef/GKU2xFD+rwFDJD0Rm
NNY6PbaKgt+8qp+Bn9EnmmfEh/zxpS//QZoHnZx0fl2XAiTwnp0oEGM51O2iVU0v
WWPoRt9IjmVD3GKYGo49Hm1hmtuvCfb/L1iyWPsUO4HX1yvUGhvFwMvVBRz7EscQ
1nPeCwT0JeVUXEDaCpnOh+rdEFbmbZEGGQJbjK9Wc1kqT3BRcZM8zCva6tTTA2IG
RFaouMCsorshL9Oa775jvgOvEgcc8VTrmshaw+8zc9dT2dbAALG1cmU63XWjQNtD
ZSPhkT8ioqg7DAJKG13ThKDVBdDcBBiR3YPVo37kJmjygmZRRUVLSW4wz4x2ngqe
xZIQXCeHf1V7KQwe68wOjE92AqsAPRkk9wT3QFrBSiN5sIHpIJGMkTfAH59MAct+
cnurvjmOaIu2RnQFZFxWfuVxwNjejgzXWpDrQ/hHSlTqABbTILt8MVuonqNFHB8K
XARWbOs/GvCECyF7nujzqvusiSwPt/ywIijdC7R3Rjm3RoWIE75ELLpuDt0Jq1fk
zglWcrfiQbleCQcPzgOi2y3J65GjC1AiMhCScvHE4XdPl6bJuU3SP1t/5ozAK/E5
4mHSmocUa+RBaZI7hJzkvHi2U6b4bqi57m7RiFuvI2MMoZxOEldvomN7tvmJG6ju
lFCY2tvYeV41djrYz7wR290n4tsEtKXk34RYrVK4IZCyxeg7eVekz00PUBwtUoH1
+/CfKrHzGQE/T2Y07WjphRMODoUGcZj8d3/fV+Xp4p1VHOKCfnvuoH+F69Nt/y7Q
bcrquxV7S5ixsgFx0v77SDZXKB/h41OhPxt0MYQinuBTM6zzjBqdoXEbOJfQROPT
fkhyxVzSIL9bbvjjbMTgO4b/bMQgH1eYWoivs/2PaRemwXctwEILevwfpeSTJnRm
fpzE1c3SEOhi5nkuewlyCoeS/ghUZ5lC5iOx8yX4hzqSJFnAea8Rx8hvvxVCeeX3
oEXp0Ov2uoqEProgQrbimmAApKYWny0k9jjsb7kW+pta6wYOgFhfoMp1nu5Uvsx8
GT+3SdmbHgXJoEyxJoD4fMkQU9a10/T33uyTz3bcWIWyJDarkEGbYBczIbOpIsXF
aB3dtlaNYHt+stuoHNLtScLt5CXtpAgnN1qdmsw2g/5h5PZY10wZADKjFFNNSSlL
7VwIrARvNasQ07mT1KVPPnzyy4CWPpl+VS33a2I8FGFmtAyOr61a8cM46+SlQuVP
2pZut34llWLraozXXCgpX9c1baOpZ7uW0E/J5HnBmUx/xZwthNIIAIqlh+widLs5
DlU2FrN7kigkZxvrn3kfIF2NIW5H0qXxKgQfrh0VCN/OEFa0j5NX+Di98clJa2SR
yEyNZ90qHpcRg1P+UVdaLe087kJ7v+yAjwFvTOR67R81/4r05tkFsqVtczLRTFyc
GGVT88emO7Hs99rJwjYryAN40TawF1AtGS2adVcK2cXMDTeX3ULdOOTyjx5P3AsG
St9odUG7rn8PyWwQmAf7BXNPurlqkg6dlHjjPBQfk0V4N9gbQDY0fwZDlQemN/ap
gi0gsjAjN000F+Z2txnfJHftJhaeiv9j6rikG1aXGqFmxp1Y03KEXCAxJ11zShvP
xmT5OXOcRJj+/jQ2Rbx8nTVDVuThIKlJGw8xXqinOsMMTzUUV0685IXshEFgKfGH
KHM71qRm1c7XqpksoptQdI4L3ZUIgEKW3QKjkrQvWqtF++i7lbZMZkNVRxdDSTSy
7Jbs7uByfYA1B0MDlcWbMjyV2fbgs+PjH0QQPNGlZyTZwaOe2jCrKNLwQ1NzBJFW
oDcyObJn1U8SqeqYjmHABLUyKgiIZTGwP6D0i6kF/Yovkjc20ohc2/e3bIecebgA
Sa4BiZ6/MVKKMyle21WH+JgKdMFuLsBnEvS3/PB6XjEW6k8K9UAU1l+e62iEKQkk
nF6LpexNHUUz03Abr7X7srdRs6bOtgLrkslkWUxjY1qhCwSFnVSuxtUtsAxzxWsh
HdiiSeJoFm321Ua80/YZ1qK/r7VsUrADvn/4ha9tnPGm4nOBE4DsFfDQt+NkVw4f
2MZPsn82G/9gU1FkH643XoQigqZBFkUKCCiNMTPE6gR7WUxbXeY+KCDUMlsZfTqS
xMV5YbGXKo/yzgBzzBID9GHx1ADZVRFziziLXV5O6mw0eOZ2dTLESBNhyvqSn5p4
ONEBPWlLBEDxkpOPp7d1pTdPNJ40t9dKZIIzWYJvfuckWP9oqXoURFOu0OT5bhOS
l7CL11Dp6jsCk3LrQ7btF1k1PjGivJAI+pv0C8SQVA9Lmaxc5ZSf8CgzoPleFbCc
6WHzv69e0XhM3dMAO96Bn0yDAuSSrCq48yPt04uFB7CwbawqITCfimg+Y3pYAN5+
6U+AT5OOSlhDnKnEP/Qm8H21xWGaKVVTHPdrtYfUQorqfbWS3HXr5fBdr3sSPpSO
srnVaV4gEx7JaMIXmmLTQ9ozGcA9YcPQ7YTWMypkLtHFWU3Krx2t5ICSi6rr+sPG
PJMxvFw5HoFldsW+nqRZeXI7sgakPQrYUcc+TPuSTcgYFC8+DVDrTYUKq9psGaDa
EOfXJn3N1Ad6baBIZjCF9t5msjSQzvtRaiC7e178JdU+5YO4MqIsC2KLNFfTDmqM
4cuS3Z9AiTH3MHt0cvgM2XadLv4/1Pe35ibVdEvzrSedWjvtm46ZcQ/9nH59vwXp
RvomiqPXwdTIqD/kqD42wc74Ed6pRiFr0kRAhRBAMV/JFkhDs4EW/y0y1QPYymjf
pRMemeXAxVZKNYunybQuSNwvSt3tBSCa+o8A4xHnGhEehd6j+vnaUm0o+n1kFArH
o/GNBCNo1FbDJtyQO2p4lDJ5KWonLb+X98FXzeDCdZJkXQft6HL4g1zwhUeLE/Km
FH3Q/3c2PO6sWJv7Qr3StCObaJ4SzOC++Vujz0UxQrEYH85f2Vb58DNO88b5XT7E
AcdRog+bxZCC+fLt/XCM+72Ao9hP+NItlq+jrWfKtY5lO1F0qm6d4jgckVC4mDv0
el4U9iVmB1yXRTQHQA7qgjYTbNzyAC4Q6h4sOxS155LqkwPCc0E/U+LX2BNeE4D3
9L2PRQyYJY5lbXA0PgghlANr1GvEKe4yvmS8hoEl0RIYbqkmL6S/LPs/4iKsPGf+
QlnAwO9Wlfw/ra8FxqBOrZPVPfhL5O1Y7j2YO2JlbrTB03Lwd5NiCY7U4R5pUxyt
i4YY3sWdp4dB0+ZHHU5YZY9oISCOli+9CYgTVz+cHD0ErmTQt4yCVf0eS5veoKOQ
IO7s8FS8DKvQlbOu5MFtgsX7uJWeJLlfAYS2IwIm9aceRCa3AJ+L4Jte2QqU8vje
7I9du9ltwLcTAzE9NtFaZotGOsILLs6990v91wukf6d9BhT978sJ5tYhtKvzRw6H
8Vdhf28M0GvLvAx+lFugfoNSa3TB//pf8mUBCggQXU+OpdXwCV7finnrBhdPMDpn
PrJdRGwbIj0a+78Vs8tKhvJ3Rea64A8eptj7NXjwhvGzG/hG12KkdY31GykrPXW7
IO65Z/tC18F4Y2BznNkaoOW122rxFrZ49DmSikQxKX9shl0Iz/XaDCX4mvr9FVRD
GsZ8db9j/V8FFxEB6EmdB3p+TeOtCa9/gBNm6nEX7Ubbv2jO6NzyIKKgs3//pnlS
jX1Z4X9wvym6Eu7788+NlIxQpGQ2pDfygxafbhq8xu6duqRVYxFJbJVI7236qCy7
rq7LrEYNNyCLAWH6TiA0p5ZTIcFPsEp1GyFR5TM9Jmqz7umBoV5Ucj8hWcMaGF/H
xK9MMNPZRHN8CvEODapBTzMjpgrpasl9/5vH9eHXCmbwBu4ahjOyXmEOhZic8z1c
gtUSwxlrVYZXh7YLvDGpj+i/Ehis/wqg0qZseN4UglCg6AAPdTZD/+RdglK3Gef7
K5sSRTUvhCy/LqGljdTr8yzz9Qg3CbPdWv/HJP3Q32UNxovX9cTfh2hmVqNZqIme
yUX3+YeDEcv9ppEBbqbU449FHHKhRBXrSrxT/wcYUcQLEVmsnBwgD5BNXyvFYIIf
lk4gjEzBtDpHWA3dprgYgfFlyrqNQRnjt8fdrFtxSS+xSc1EoEE05aYDTvkRfEeZ
mYyneVriSfANORlrR0RZWNcaKQNpaaU4DwkrIhhXQBroy54TZHapr+YJv/il68JG
d902IDJTCcsvkCNM03K9tdeoV2WVgZuO8HuGXzMyJXbKVg24w2ivO34A28K2UGSs
vBdI3wRLv1ocmWe4PQLMnn5EV/iKQazIbKtcxg+do9DPBJyL/y91DWFFv9J3x+Im
9VMGLgpX/KTZBEeZD+z9J4dbDPus5Nz5rj5tMeeS/3egFq2hCO9EUkI2XuRhjfCU
phNuuK2NGM2RJAHUvMwWJM/rKbBbY91BYqw8Zu2809FtiNUOtwZtjCJGuFz7NPti
E5CJnfE7CH9/yQQ7TsBGQK7rLoxziRTXDJPyLl81/CNopa8tK2q8DIZJnT9DZR/E
uVX4cEhg9wli2YkIUjomAeF1poMoht2syla5xnQSF8DrpgRLDgxxzy4BJt4xjZ3l
R9EgSEDrMLPkIlXqI6+D/qoc0fPb/uZ+xm/3wCgqUb3Uyat+kzCESCbbm+V5k3IO
oyjPnW6gWIB1jXygRzBpWF7Er0JxM9L/jq2bZm1++XKXQhSESXJnzS+dwOE1os40
InjYosXzLwGXGBhS7Rnzr0nAwQ/SUjaYm6QuzXYDr/XULABc4BeC5sPUUUNNYEPl
G57QfH2MiqZ6Asj8lwCv5TJqeviqsa8EcUk/sNMuALxqLwNmkBkKAcWpTrA3BdOv
v/XKcdV17qBlqMdzST78dhllG8VcwFqV6g0DREj4ThqEunwFq7qJmx/e0ZC2kMvD
+qAME1BLTNUSsFsBb0QgY0EoRbwtk2w9qz5fbwkN+wxN5W31KwI/jiYQgEPdRdkJ
KU6A5vHPOc0LuHTpXi7zTtv58/QnIR1xfTnrR0LakCHk/+AwkMD2XQ9ZrjbQSwHR
WB/kYo48XYztdmYltUL+sqyyDg8wUbSFj1T747kxxivwtQoW8upski57ZnD7yrzb
iw1OSOBbEF9OVRxtu44u9Jv1ri+j/BHdwW31CeoxdfamxIPiQ53YgPx6McZl0rsH
o+hJO5SrQzG1rq4cid6F+lC0ukql4KMO5AK6RDkaDAxaTxzJKaB3eiCwkdBjkff3
amPYpqD1Vzt1QNTKE6v47xXP8qqf45gbOlS82ncXVXJW0XMeMRGEWciKAOewikoT
vE34kKEooywBdv1KGnZEDqxZIk2J3k+ZF8fkkaByAUPFdjAcmEEvljNAz/7zJtXl
CHzAchBytskGSCKraBGWVsHBKRQeCSZusPvTeQBObL7m+pON5dR/HQod21mawoo5
wxW6K3ftUV8KRVPvI7/tczOcbb6xURWHAk0JtewQemW2/rI1TaHt9SBwRjt22BeN
gC+9oXIC5CHKDNPt1Xs0e7Y7aEevJbcWE03MPtRYodldDZMAuXr19RF7V9nj4G5m
BByUcA1AzlOYQOkWaOQXlX/ewcIj3LtcB6ekwERzKw3YTtFOgOk1AlnR1Y3jbdle
q2kY8y4C3luFUKJZB0FhkWOXup3vwcN9W3pG4pimr3ngxB8D3kmtQkLdVTC8fu7n
g6KyPVWsgeDH1SjcyP7aKndQAyKw9S6QmWb54QG8lCTpuEV86gD0B7UTXykkQvJU
RRai+9WLdO9ZxOaO5b8Bhhq2ikiToKTuF7C+1e8y+JXFWn8WiaR/C1ZQBvXhnTHr
gRJyqT0cGake8uPf0pi1GPGlmNsP1cUbxPf7gZvpb8T0GNgfqvWqjnErmDkK5UbX
kP+DVjtjBioj62f6rGUHKLMqnkjobmkMo1foLLabFMMNyvm+dF3qud8OY4Xr1qF3
Va3TnGD1oPLgOHvYnHbThk8+UQkCCWrTpZNe2Gfl1pncIPTYIUjedj+ZWmYkotk9
oQI1LqRuEV0cIJjafGpYvvDtUDpmA6n8kdLRFNPg5bC6YI+oINztCaVYAUmEHx1l
C8V0oKx/kbNgldWN/pPVThK/sromo0SotpRtEOn6X+XFJmNBOOOxGuuzakMFFYzX
rfXyP+iox4mJ9KI4au5Q23CFyjqZZnfyizTnk3uNeulIkcV7ZtQnVnDjqKnHI9eK
DVko369wh4gB60sCopJ5JzPCOhIw1AbTd+9GhiqyGItNizF9LWtA0krJA0IFvOcV
MzwEzPsYc/el+Yd2DLsQ7eA+l29PGWGB50x+Qk/o+QAHfXT3Rs4Pk9BWbIS4K1Tl
ohesDWN6P64H63jeDmZIDscKGWhb4TjkAfW4wylI7q8pjqx4RZaQa/kQRTG2dHEs
H4va41IrlmR803gUiPys7/y2z8+Ym5BX4zwmRn7MAjp+X7MeJlnis/GrVaL/EPWn
jECDrl4g0AvIFSaYuZPLVmtaVpC6AZ0sPGSsHbgnl3/UWg1A3Ck3atVe9pT/1ZS+
gOuVVHmlya05PQPQfl+qQO82g0cQqb5bNU7N5JKaZcFwmLQgOW7N/m6m+cvrG4D8
cMYZJODyKj4w31EkFCaSaMmGMja4SeQ8F3ORe+dH97rWtWKiqUnAiYgGtphhgeWr
VzD4vMKZpxe90ila+EVepQhhuvo1JM8YgxFBaEHG9j4LlnBVBKem76vm72K1MIrB
vcv1qG6q6hxdUNav6j73acZ+CuUiuNxlDKl834Qdf+9U94idxmjJTODW7ffP1b3d
anoQ6/3BKdF+mPXUmn2K/blCqnNHF/zF9tX0QpVJ06s7z7D1PRI3JKAXHsxCzKol
cj4Y17rrxLQEQEm7Kjl23c2/f+jCAAmwgO3/CWMpFBN1QTFy3u9DRi1vniTwubWa
FUll0VG6eCxmQrKyHu2+5vRp1nbQwVuD49rDg1aXOtuUljyXy+1KVYQLGEeDpZ1Q
/1xnUN0sXx4jR6HC6bmX31+2xmpL/WSAUK3qCtIDKeJaHrSSNR//NJikcuwG5dGz
ayCown3GhcB88nlQag8rqNIFNShMBakYomlW6xfLZdHAEV61NDrLqkWGukTOZrf3
tdBOQW02+lC3VjmM0xUhsgPrhkHYipDYRqrGYCOm/If0tlQM8lNaUeNoC/vmX/FE
HcMJ4Yy6Uo7KTLUY+6CtueQg3mJmK/5XrrkeEmuK6yHMRD6n2GtqufA/M6TGtKXm
SrgFryeqBBPQ5PwGqOPltboaRaTHVZ8jC2TYFEdock+Q6zd/9nw9GxyiOCxVCb6i
PQXfidSZu9OYkaPXk9XmRxLT7w2gNsxLHQNDT0LZYCMlXqPxkWgMX4wgeRRQc9hy
tCD8+CH7YIi26COOHSY8QCVa+Yuj2y+NrkAF6ZjmTnFCQty5ly3bKs2kdlf6eCfL
Sb5kKINuV1mHpsAwsGtandLFY1hgOfr99zUqga/wUbNH2s3pIAynR24speDGSrZT
0nyMiTzaHxbNGpVgraHJPw27Bl8b0tGleRXJdl3ps96vTVH8K9p6JaoXvIaswJG6
r6C5K1kJ+aI04X/uwUaVpywrfoDgnhboA39/cDmV6oxQuWKIqt9DD19zXy/yjt2T
aEPdPHaujeXRU5qFxwJCOO8rq0JPAwh3MOQQWAhymRjGc5ng1/ZopfGyo9Em1Pqv
HekrXDM/OO9NqI1+ZNGFYNGZgj//PrHyWrWDdyOEEf5GWYf2EsYqqCH0FAVhLuZ1
Uq4YGjFAf4n0G+ndeNjEPdG3We+TsI+bdAmnJ7FhQPaX9oDc7KuGe1onEX1zwDHy
slHOo4zzVpRxsHRIG/b6wvn4GR4DPgl+SbFLke3zf/tCK46FXVFKM71TxVz14EmF
7rX8mAbqDBIBn1B+CDsTso7iL8/j0SeH7ZQIBoN9tmQVJP4jboy8wTLC1C6XgBcu
5m2+dmVs5NsB9WX5C3wH+FZALApumKplyBEzU2OQdK9fR5ANsqIUQ5p7C3pAXRxL
ikwHpt9LL49vtzJCIhC63hHfqyedAKPMISIrEAnYWGjhB7AL85fnE3ocWNQdFVLZ
Uco9b8r9Ys6ju05ofx4o/YS2PGSo4zyO8VwhPE+SE9q5lKwF2m2zRy8/FTv4WX/i
x0V5y+CLil4DrPHDl/K2wjeZQZvJqtUIne9qhcBT1lhn/hd4fn5e0Gjtr9f/kRlL
iXw8MOMAeL3iSalXFJZUJkwyU+XIydpv9YFfD3zLU83ImVcoOqc7MNe8SsZziKzP
hRGeSemHuscsogm6P/jYyltOeV46Zd3f35bKtJpi56yEb25WGok333sMuJ+LrdYB
OdGdTZOlAf8P4E/HpftahWgcAjyDl9ieJPpJgKLVMRdzdIEomp7Hod6KjMW3JNex
nfCEjqIqd+iqQAl89bFnZDRTtfYCojGdUXgqu+wfLTprPPQ1a8dWfelNZ9DgWu4m
OOdT323t92sRs3DhJo4idKlRKLh0aCHv8dVX7jvtDXvYiIrUMU0rewMHZCJXj1LW
C6Hv9tvb+p7YPaCEoNIK6HjGmgxY8ZKPzxN0HYwKQCk82TG4vk+B9H3gYczPvJrA
d/BRQ/sMMrezqBZkeeCLNDAukuKu8sgTGwdWR26kGzGmmmhhAt74eT1l7LgzJXxt
Jh8u1EMdK8HEH2obBLZxJQrc7c0V5pwx4STrlCHRefM0xdemc2FObpoPiZjf0cnv
zo8ru81ZFHi9KR9xPhIpSD4Fm2iiwN06KETv+A8KZFcyVdkZxxOyVSU7dlpbEdiW
lJg89QdqVIYx/pu39UEhiTfkttRExj1sPvQtbYT23HACM4wrOZmbgv7iTYF/RTGj
1iARbCnlv7lwa1562sbbwhIKNMIZZgKjXLjRIXTQHYQQYxFRNK+fo61M2ljn6mEh
panIaxQl+jPrC0LpDw9LsF181X2DBkgjDdPRffDbLYCxU6DiLtwgLogiObZhVH5z
TyIskdq/w3p2POeK+FTAaXSydHNAVYXvLoGBIgg76s64Yso3hgbElrn7JP2EOe5I
GqHqFtyKivAx7/YV2rUtl99ZXJdJ75Y+/NtEPFxT8riKpF7X3/1/HunvtXUvLLkM
v1NU+Nk6dvh7kNA3MBOPRwRQLnOCJqA8ja0HX+zzJ4TVk38tLXQ5fKoZhh8F6Pnz
4spGRnCJI29H6z1RKQhpix9KJ+zjU0Ehns3UNKuKOSqhXHFTj8O8ZOnKsmaLNsv+
JEFepaiV8YY2YrBjNGq4WIY9C0HFEBmhadOeVMc39yauUx1Z26W+1Tr+ov5swEIt
MjCxYK+OjqqkUJrL7thkrhFceiwwfvIzdXUcC4QDMWOrJrRTmq58vuaIE2MdMHK8
/16qq7W9wlsVx4boW3t4o1IsYWVijsBa9mafmyWrF53yAuPvsQ/12abp2zXGzTBR
iPpAPY1YCjqUmXpYI5nmCV0VeeT7GRAQampIiNNNubfB8VDkzOPqXmj0FE+Ft19T
3WHItLpC2p+ox5346rOe0ySOVGu1sBNeZVaDuFiwROk/+ba3pYwwDQQi3NUKCgvM
Gp4L3LK/ENOJG4qZoo7Tj6rTpqBl6/r1KAJjKtoadR6pYP3k6HEbiMCysOSFqmrV
wpRyBxZxkHlab5cnWk+pa3wbKTErYDGMr0XxbN0XWDsGuMV2+GxwfDqXbnJIUGyQ
l7/+WpAyCa9OLyDcTjPkwg/soEnfBPA2i8hMiEnhAvh+36KDWqTM5EXqQc39KN7K
sAc6/b6oG4QU13P+fcJ4MRH8C6EWzvY0eQOeCC22Q3aweDQiJoCJ+oPKObdYRayz
yx6N5fTZW0VZmZHLu6CuX3r92SxqUCwz7VORm6Cl657P4HtuZe4kFsPf0am0OT8H
1CLh2ucIaA0uWRDSgI01Ingf3Z8RxW4lGPI52jTiHJA0HKZg6X4WfKEdMGEA2bOY
yWLm4Fg5oreehEboSS8K/IR6lcp3xrbM+o2qdG71MIugnWUmdm5pmOGgvHRqwKhl
yVNjypvMtJjfUjsAsdqlJD6hPGn+BVs2V3G/LGezAKoDfuiF0IE0bwjL2l9mCEyA
BzxpJOPImJ+hxvp5klVIXMi1f7xuLfK3HnVfZgOMscOoSzu/S0IbLTO3bSAKoK+p
4ogwe96jkLOzACKDsfw+mmDkgNcuvH7gsfa3nMXonx7uB3gRlCu8h8rmKtfXe4xy
rixnhfDQ45z7qrb+RguxUceTaSSTIyPq6E0asvK/0qhQ4WltTWLlDMXV48y31Fnq
bru9SkX09sNUOPxi121yotUofLq2mfIGar7rwz7cD4gnV/BpqFStd8JU/eYPAt8l
EKMCCy0Z3vz7jkUBweyiGn5xFYMPJ+OqkqVVVP2OQ3xx1zUoVPMB4W5qMxgyTve6
FZPbzLzmriaWJXPUB0fJ2ffUupw0oBd6+Pnj4W0XYe6Q7PKMaaTJ6Ht6SAf2yD+3
bmz1rKzeOeHaSX+/3R+OAnOvnGdSrJLMeGdCiIBMrIMLtOFPf8gER1SZBAWuOK4R
Kdx9pLMX/da78k4kg9Pmc8xD9GcLeYLpWKNfj7Ub37eIlpanYGYg3CmDLVyRVdV+
EpNTtFBuitMrXQmTEc+Ypi0LvULquYoe7WpN78bwuvP8/pEW7vHIi7uJIKE28nJ3
MtFAMIjBAvCBovUwzLLZ41XSZtVZtKmuA9xbztE6qx65jfwn/WoQMqHo/SrEzE7b
/SQZtsaEDislzMzwcQP1CLeB/rsyb3ZFb1+mOPKV0X/vLoWjrl8cySal9yNhvkUP
EUuK0sOHgow71lpXCNeOapHI16xhEojsJk7wAceArVFOnk15qp8iZwKYSkqJ8H6l
l6Tu/hWcMxopbnuQTpzuZ3o2lZErIvYql6xXC+LUgPoGUdpGVpSdtngPJUK1Aaj3
7A5x8ulUBZMi/tc46R2cYi8NKoumVKZFanTo+YJoI9Yddlb5eqDCM5xioXWxa4WS
RX+1vG/TvmeWUO8LlRyD5Ps0BWraZtjrkccpU3Sf/V/YmG2W8dqxr6YmuTUXRIwb
AMAo5zUmhN1VSA6cbq5i4erKlWaLoFzOxDl9xvm06Lg8SHzsMsmg0A/+NA1MBquN
BSdk21uc4EjV1XiOiKaqtCWas5PosZoMMBqaaT00+H8fq5vZWKO/Qv88VsDNEYq1
0vzw4wRJPdJSFn/wOdnVUZExZLghuSbXutRO4766lZbL977T4aGv/wJDbSpLbjXS
mntKm3U1IUOsxygrGo4lRwY67ipukvDMU41bgNcGwVrtx+vo7uozv5z0MBpn8En8
oTS1N3TB2AzGedb/o30VAXKIYlH1F7h1DIT12wA2PDiWGf7jGVL8xvkGGKa7jvzN
7pE0eD8vuyM02YyD64pgCSg68D7QIcVbbzW3lKbRXZBtw3FxA9k1TGpZxIzxubzN
llj4a1H92HULCe+NCo8ocxks9qWN925tfU0QFwLuXOJI9agxKNfgFKZbDjFLGjTk
VGrpswO2Y4uTLCZ2FgAs8HcPhcBRguz5s5Qejpw8Yh4jcrtkmxhajtTMrjXCKIhA
XAqs20L0jl15P51ggW7/1lob6bwsBqNxiR3qlIkIetXJsFF5dsaSsK3mfBVmkEd4
RGgatrFbneWqLDWuy7HVqKenVxd/ey579te8YZB1CnkOdkG9rTRlcOiEwfzwaQKJ
FUETWpN7n24JZwLAB2PCECJpHYIK/5X23f765J8m++ztfT/fOYGHvXwdn3luqYk8
F3JmHhWctFI9g79osIBOQlQL8T52e5l9srbiyWbG3UgS1TfsKCfYiWXJKX/ZgAvq
p8TIol34UQz12rzDfJfCaTW0UH5+fEBSnVCpglf+KJxnL+CHnLvLUPbZvVC1gyVG
sU45yXoR1PyL+OAr2Qe72jg5hy4Dcno/x2540yZL3oBkLb/fLhkvK9YvN1zzpuIW
f9D3pL8HjxNfVcneLTKRgUezOlo+p+xbawG00gvUe6uQMULs/lt4424NaHNdMf42
ZC/dYqvDQivqt3CC8t7MtOWS30EJCvhxjr0pxzNA0rMKMaHmADjLZOGRmtO/prBl
EWFJqkHDVzM9Ha1MBnhXSx4uxhLQ5zpp/xrh69cBK1A6/K3UJhII4FHIarMJGVO/
WImV+kwHIS8voLy8IY4QQZpUDJwVlmeWjgtNoXW85b/2ARWPjWLEtW6iTjknl5Tp
vvtCTSsddoSaJTBvAaqeQGhD//rHG0XyIG0vYoj9rPqqF54tz4ld6wvHkq93i1tt
b9IipXiFNEbLFsDAM2sflwT6eh+qL/lAU8/DvXzn8pE5B57b+M6/QwhVfVcuFzDC
mwrdSgvc9FGpyu2TmpDXck+HAel5Ty5uHipbkEFPPOzNQWI8JFpWKg8GBK9llw5L
joIi5M6KGCwXwIdtjkXH3DvAfU7TTsFq9mHHhOQXeWwfCysqj3bGqKBvLTcZyHH8
2/3nmCNRf6xAKEvGXa6M7s1kjnWVd3eISAjXb+Y3m124++42wGiJghaIcRggQPAs
YqccryF4BxwdrWdeb1Os85TOHyFk+SUqQsebcwKHzCs2sSN1C/bbQtvipUl1NB8d
XQhtDwTCeIeUsK5I6alneaSMM4XT+zk9Vsf3K2Nd+VQvrUxJiy4zDgX1w+omjeWv
hkmUjBuq1u5Mo8W42HoHj4M7XQgGaIFGj52Eu8sZJD9InADhBPV+MpzjUkyzrtOZ
/85T3zIWpj9xKz3tVgHq+b5NKVrCIv4bH9Yz0dJEW+zRYaxRFnhtliP5JvvrJROy
qkkAL+Oh8CLnw7wiDm0043rdib5u60640dSwLlFY3zjR5uIe9L5H2YrvxpXmvOtg
6OspOul9sX+1Qzr+9GIuf4qKUamtxpawvJNBPEwYwWvy1ZUBWzKl4w5OyV2if+i4
dumpe35KrfskI704ej9tZgRRWPQ5GlMYFMIu7jbvsR+YiIwb0iwEZEnJByBdPMEA
XQhd3fcu6AomzomQaRD0IXf9wbxdsQDwl9zvrXRr0QhMfioz1wBw0OppgtClzz5i
F1Fxq0nouRkBqaj9wEVi7IajVE1q6QkrQpszRWsX8EfPeULEILDhc++Yneehb24t
THLviTxiV2apCwOVrKTOBbbFOi4/pp7h79J/aN/786uqbP6RM/eDMSiplC9OrN1C
OESrJrVi8dr/nffuXtirLMy+z3xOz6gA9g+Iff0i88jFoRUGDYu51I8i0Dm+DXPX
WMAhmNx/ImzuAzz8QhHiEnCmyQRcbYc676RsFiosaGTNvcU34R5QzMc4SN+tm9A7
PhdD4qCQBWl7m37r9K30L3+QJSTbrqZRSmbdZUq0i7amz3gLKSppMA7T1kK1S8wd
rAwWFp4j1eESo1YKYyIgkyQUd2H9ByM+fbYSiBmqV64RqBniQKfBTx5TklANmmif
Lsdkq/VWA+PfykGoJWaH5khWHgM3uJZD4MvHIlcgF3VYgoyfLksakNy2mrqrPekj
CXt/k7uQVNUhVrT+EPLgrt97KmxzlKm6f8WiYPNF13Y1vAs68F8xmek72c7ajtkw
oY4L5BLBBw6jXP8/rgUng7LasKVIyisWShkC/hlS7fqjAN7WVa0B/iC6M+KopYE9
Lyur4RzIppYQzJmDNuKdvRA9q8+aBVmy5bd5MhdN8TrlkweXzdMlew4G8jPRtEgH
SdvXN9PuXC67BAKUYt1JFqyenLxNlYHRTfp12eEv9hgiAuCSZpwse9Q5ZLwAqrtD
NuV+4DxTaNmzp4S871C/Rc9HOm77XfODv6M1u0V8KHCm8q5dd/c99yf69O6B3Bhq
qY091hMi7MG9oAVUHyOSEk40g72GffzM8Ib5iEcvslIl4/so+S2VLPLgblONbzFL
Tmpy0af5pcxol+cvBS1rz1t2sdyc+EBkcYhItHr0k/OZT6sRjQ80cijigCc6jF9r
lyt1CEt0Ea0rev11IwX2AkljwsCdq5LARN+qC3eADET/A+E5itxf79Vp5dsmpKB5
xo5WacIxU901Sjf6bL7z05mn/BTN1Trc0VvBdFO7EIZ4/qKhjMfZFD8DwqTe2IQ8
GZf7AboFcLFRxvFQF50vGQPijai5yEc4JQ7zUvnVH+6HWLKgsCIjLuc+qeshs/Ug
HKQWz6IvKngUlNYGD15Nu10DcZFsc7ak2Heo0VQgg4OjDr2UOrD4fxTfzo2RyTNm
04Ir9HT4kvTkHkP9bczlARjJJZ1c0bSumqQ5mAHkDVyubvTY7JxDbSUc6IN3Jx5Q
jBHcwCk4OB8oSSYg2GzZLe6hRzH6wP4LFFkjCFdBLa1wEEvdu42R86doygM2mCqt
dUTfwkdnG06wf8WbMaTWtMZ8oWXqCLvdM97N6DXysHx7szlF8hnQP0RtbvJfmRnp
z32NGJce7u6jTXsnIwRv5HnEHNCs1Vb0DIWDPgprgf7SOC7O95ShF958OrRxaQX7
A4h6e2TUBHVUGAFdx9dNtoyZeAOQ7ORZBnrw4L4xVAIcE+kTxoSDGdQQS2A78V8k
P6IuEzwUfjvXrPQt4QQAZRWVkCp8rC86f8kWlTt4ObrRGV8uNl5dau7bc+f5Mh8J
LvGiXZDBkxSFBEVsPMagNbpGzJnIntUbT5Bjr+o9sXeKH9/13wqeXELa2ow7ivW0
zY6Dd5eADWpfx515ngXBJ7TZ/Yh+KwGH4EL/MsnZJSmZKGie+C+Gksuxbjd//IHB
MaVfu+e0E+gCJScE4Ogybbj75D4E6SMFtvNerzD64/sXzBvpuTi7k5iVe9JOsl6r
0d6WKi6MC9cZiUuJlvVHLb3stuKwvI6WkmeP60noSEE3y3ddC7tHX5Ya+d7cZrYs
8606dLLAmOO2B2HrMGwS65FD3s2nn9eDbCXleulmKS7Ry5NoU6BCBpdrHZxKxp/N
/vnHV+lD91m5ek3Ml5pA1esrF1CKqce1njtUltYXmKj0jlMXOsaJAKjVFeOQ6KeU
u4t8mrMsV+ROZ43b13CthTdDVw2Y9/P6H0yp28WyJ//EO7z3d8uhcw0MMpl3QW2g
9+e2Q2+RPkhoB0K3YKQAjHyCqUoIZzLc6WN1ESwnOAqDZDQo3F6bdOHzJcVTcgWJ
57JGO6+GICwcY+EMb1sG7xlt1hbws+yX13A6Ly8Fqs6F6OCV+iM8mewtdsYTKMzO
3KqxwqRDHSeboCL/NqI95DsdWR8b59DrtCqGoGM7mt+jZPbyvoflmVfdlbuvD6Pd
awPJeA4O4fbofvBN1NZURef3UuI0uOMZ/NqN2qmsXUbOBCAgT1LSqdrQwgBh9yex
VH8/jzwb/8x9c/woQjPb4DGjZCOYchjFS//mpbKMlmYb7BSwbTzCjfqe3czOH3I8
N9tfoznxB+XBBxROBndYPNtnhYVJAnCb8iMixMGWKCyxaJB8t+udzPgmaoZk3puI
BYy0voR6wbmuS4CxN83zcafrSiCX1SAF3WPPmYjDdfMR++FZiX0yRXbM6FtU+gvb
wpX6N7b5zSuH68ofUi/nTDgcDLRVyZ+xcWXRKWEKXnrenA+tCKnHsHIHPmlncvx/
M0VT4chelk/wjzWG5JLtqESzLDZM/9ERSw0xhbWAyacxLauA60C0WWiUrVBOpGe7
MmaaI2YmdN64SV0KBZynXY+ooYtkpw3mpE18CokD3JhmgKBvl0cMUY/XOkA2FaC4
2NcsE2hdV3UZ60UuKLa/OZiSFNxX5O7EPOSdAyAWR3qUHmgVhdOrhX6UkipnAVXI
xm3kmGGcjC+Xl+qm9jfYoxXu9A2SKEhRr9hlPXcecK4iUpH7AuxP22MZZOnd3TeQ
S7NPjicMAHKks5h76Up4NwViqlEyqeyqS0OwvL2WdYwTmpp/HVQg8epiKq6gmUPE
R/Diz+mdUnsoUsL5iKz8oIxafiyjrxXGyqLHNzRQoTnf8pVJH05u1UF+H3wTNOKr
pYewl3ZMTcFtipiyIKh6TTh2vk1W1eKjtON+JCXIxTU1z8A3gYb8UBY5IIt0u9GL
LwO28sHISTdcAer1GTOt7/abBKrqOefztT2cqPeTp53eU1kqnbVQydnRWDmt4KQk
a/xrgSrvxXAqH9IbdrV7Mv/Wi3sdJX0LqPlTqOqFEv6jC++r4Dw2VRirlqEiPVoc
t+wuugc5Q9xe6ClDNI0GWZCEceXhFd2Yd+a6XEutazg0q1PiSejUHVajwek40PsW
yhVKj5Gw5BP9GJTq9d3OqA6t8d1+n0mZ+ipPeV6vlp5lVRxPtXRSI9Jfo/fvsR1G
AGsop3TFPwMWJ22nD9eO1hNdOukHwOMespM0dym3vcPB97aoxpm636EHlr4sycZz
x1AU/Ol+jHWDSoazHEcpcKSmeqVKaKEyLHCGkNTzN8ixaxeSRBx6lQUAPfh3EqHQ
Q3Y3NM9xTjG+GM9Cf0pOCbfMyPm3GdQiuIgwPtaMNsao6EhnLPpro9o1ayDq3FAE
rOoMH1hew/pyOfNhSTMZwWOrCZwKC0FT3b0+NvKp92lkjJ6hbhLSw0TIimSFO7Md
Z8l8cPehKlysAqciXD100+FicbUwxoQDv7Gtt05pfeQ/7G8DgxWzmhhkUp6JFQrF
RaJSBSVOl90oo/kGypHc3cdw0DZPkRstEHO6VnRr8Ntp0Su7/ZvBZLDy48bLylUZ
sDoFA5q4pwKJYcpVvnkC/0d6p1ZGh8FtpBkpBqwHAx9ASnWXOxDvbWOuSlY1jzJE
FCbgVnZpfVHcwN4De6Cgr9cb/lzNqeUiqPNyIxWZZI9iemh5sNtTexHGpIUI1b3t
bpXWSB+o2bKsH5pGtxOI+Oh8PndEE9rSzaMUmCc5TlOrXeeTo9eSg3nQvZ7tPsFk
yXN8PRGzY5TxsnZO51RExntmqahZqZWnBznm4yidi0n82nxGfz7E3ZB10w9he9wu
EWwgtwRFzwGpZgIfLLyzrNZSiJ0zLxv2M3ttipVo135e5PuU/yaxdpyffaYuZi5I
l+EAnOk/GiN1ShV1cn3FZTJc0YA+PZNVnpM1UyGcJ4e+zviI/fTZ30m1eIui4YiQ
RkDhQX+HwEDTEhYN4X6Gy/ahqjOUcTX/S7zTxyjtdQOKX2ZhIckbCY9NwOz81iLd
BcstwRV9nvevJ9wdNG16jdi+qBztPTPcdVnKbvsPhHxYnzE6TjWjesMid27WdB6i
57+deseQLdgwziWfE8EtVYy/iSGQBfShgWKQh2UdrLOTnmc9rc+Kw3+NqIL25SZT
gdQDrR0fHH9PCMArFIa4Vu+WVI349cgPJbo71/Pc3gM04RVOCX0BUx0j8MBOxIgT
ZY3Xftb2jcEHVujKFUnnNKkI/mdz6uJ4ZoQSN9Zrt9sehcFYhz/aq50te1E5VFGN
jrXERwMkn7ApEc1ETKmc/NYgrnXYATNwmCRoI4zzM3J3YoSAca2flzPPGIqdHc/X
uFt/e0FsNUZRHiezgJ19IQ3N9J6U2oS+a1S/+fy1QiHfrMKTrheiXbfPWltrz4wh
L9nTzNIET15MP9ml2MjoimGetb5/PKmPLMFDMfKHy5P/nqnL1E0V385P0n7LVkFU
Imtkpp3rJkS/QrAidq9AHGdZKyPlh9XiGsAYrHiAhAGsu6xHQhtmTvSJOWfKoY0p
LcoMcA6qCb2uNuyF2MasC51Dgp1sXcPvZ6OlCm+XcdkeugmQBzCYHqQDf1QlczDU
1iJ/RGaAkNYoMWSGLXpZ4biegH3VJHcouXzPodFXhy7u/t7/fl3DVmV8UlOAaSCJ
JM50p3SrSI7y9bk8xE01kOarJdKy7sE2MfFzjUFHGJ8dC7kJfLnUx+DRBXd0RSoW
88jIp6mRybzNCfHmvBgfxgbXakCqgzcWJRfDJWGS0NrXD5wUOFyvgCqrLnO8PNfi
/Ps2JISkOsdNMkn6+BlhwtRBrUezMZRnniyh86gEuBLm/JPsmExoAK/JQ2Ly472N
ehCTV/GrXWbuKLj7MMYXOj5FCcoymDLZZrx7H7hUW66KZxCv6zfJ54UcGZv6HbKY
mMzAINA18QogbN29GPcWBC/eY7AgKqSbpHkn/dh/aUREZiLduyOkILnrEy0WgPiI
VFjqbz2YI5myPL8NTj+9AdB985bFeuFKBB+t2FPoBxdZwGwLc01KTnxSNbA5RqWC
8DPwLuQrq6yEJMGGvwShfJf5QHbizNqH5nBoCdjEXi0WLk5lx2FOffNO23HXNEjN
Chgfka8cdGdHth40u7k+efqtyV1viUzID1EkVH6rkoaQJ8k2shUA4myLsIA02A1/
zOqg4wUE0Vcg1NQStKJ171YgKO9pfwlJqoiYVxYHNUdAXwle9VsI1qryySTBm0nZ
0aGBhivwWpWqF2F3F/cLgGGVUYfynS0PQ0ekaNqeIaaJMPOtW7ul5yVfluin6js1
kKEGkBzhHxaTbEqRlQ+IApLtMysmfK1FAeXCcnvx+e9fjQrhvVym6pny7MjwBwk7
u/7jFrhf/P47eMhWLKh+Wt7NUsEEhyfzDQdaQnAhWMDhN41P12q37uz3N8kmeoU0
Qsl5HuE3F6pyWg1LSkKFuVmvCrfASqCQcgTeIr3k4pAvElJFRX+7sIv2ODNZTGoN
ESzxgq1cEKARF/mDv8YTWcPYeI7rpIe6oU+s0Ktk1D5wmHQ/wDV+pjxGALdiqzBn
2fUEg2ck6pgnyafXW+AmJnzxNUzh7bxD0xIkPtbuKnYDpsmdEMvWvYWO7HBf1Qzp
aAaU0ygG7RALY0/2V5OPC9RQurmXHK5rLIntaSR6bFU10ccczHEt5OpIbLCvw1gR
BW7swomD8k2qu76KBi863X65zsNqRKrLoHKxzhslxUPB7tvYO7Zz5mi2ea5usP1s
CxeUPS63xEXOT9TKLPTLDMmIuwFQeRUdP0NdqO2EYoE0JgXbh09CF/CfgCwz8xUG
fpLabVE0P8ZJfcXXuPhBq0iG4/C4HpwMe5BzcfDCSRbifdaE/SdX9Eg9za/ufGpk
JyXSBeeIxAIFazFQZwgbGu0yQBy+xZ9dtAKKZwlx3TN5U/o1ozcyDc5VaRtdXp6P
UL6+F8xEarxlqAq8K0WYfNMzov4sGi42/aRk3UibY4Pdq+idgJCcWXFUpm1Nfk5y
OPmV8sY780FR6sFI0SSQ0JvE4npl4X0q7jic2OZm6TAq91biBfV0UQFUVLeucVA0
e+c0SIGSvL7orpfjVWujCCu6ViQ4rh4jW7D3uIGOwWBCljxUCqwzgiqBIdWL9pc4
J9xCpu7WXRVQirz924mFs5/XZmeF4wms2SWIhEseXYro8mAYLaN0fN6na9AQIH+3
8apqoJ+NKk0CbJzo9CcSArf8C3Q7fm+1g8Bt1RPRccqSihAXW3ZhCrxoVKJymHqz
xy3N7RkropOuCAXGHFiJq6FjlCuwvV1L2gqNWcnGVAJ2xW9R8nFPhsAG04wZadX0
RNWdKOTW2H+QrSZ13M6PvPr5Fu3qWhjh4jvBPTC7gwYsQgUd5kwfzPEl346bpyHL
kAyUaK6OHJW18/cwd+vFpaBBUfhCs8ZWi1+C2p9fU05xjYGb7mE/jYWglPElap/U
vrmOd2SXjyL8BpbL6qg29VDBJ+aX23rqfVKSz7uOVG+AdXx/6us/EZj2aC+lGzz1
E8tJbD5IByeSpgxaad1RE+IGi6CbtlZSsNkj2R84xOGZuTtJ+NyzGEJOeA1EzQ95
jU2uSnvkLqW1oUcGo840DLeBpanmeZTnhKh+DWURal/2wSZ/75EJz50SqEnmKMxY
vjNa639i57E4LeyF7tOMFDy2hIeU/Lv5Jn+F7bsEcArvfQg49OOdmT0Ew7R9+kCS
faBKoHjh8iD0W82P32fujk+IxzvEx5svmiosqInODLcYL5rMtqeGExnIbJNPbIsW
tumNI/09lq5QodVEnax0VQsmA0OY7UkKCo/rLpffO89QQ4a0jbokvJTUtdn72F14
YPVDz7cfRXgBnOUeU8YgqSBZTZducXfqS91qDSSdALbs/ZI2KPRrHyb6EL846hQX
9Nmuze1T3Ss2a3rr96znh+2traNDm13Lj1JQiUeDDysgnr9xjpPQya7bUaRATuC+
OG+zh2qzkK4yzZJf6hGUAp05ysrl29Ny3dLPXYaEVyhKbwZI5rWJVVoSwKStCPPM
9SavdVweOr2C1OeCUDsmfbXSHKIVcf+UxbeEEN8HRHLFmmPXkkS3gQgBS8jPSnTD
nxz2lUKvb12m1gR8ThbHslo9vpYlavojJfWnDItmX3HYJ2NSrBylPgZhKY8FqXQt
xuXw3Kbqibe/T4w42gTICcFNBgQ625XGQ09/LSC0ZzoqybibxbKNVOhKV2AbyNOH
hijXlwOzgCsVMKDhi2ghrXJIyaJbqKFVZQOZzb+x2rJRyEPDoxk/axlmw/y1OfmH
hLgj1cvciAWx6KKZZjBNDE/oYMFMdYLFkff6659G/sxSoGqeTrDgAadl066pMFoW
wCXiBoWxq/N+m0TStQdvf0i4g+dDvtaUSxYltLzUkE+SjjbOnOFEk1i/lF1xxGqH
W4Iju6V5M132tPz2IUCLC6VAtOda6lY1vF9FSb0nfaxBf9FMpROR0u1OcR5AZ302
f19erMhwmn3WuwoppsvvmLk8NJcEWVyAZUkS/rCYkJYz1/pf1/4QlAHhWGW+WSWf
kJzPuJyKZ61NOZma6QRs3z4fPLqfyMOPNf5Wj2uGlQkqq6C01HEdbgBl0fD9ssYl
6cW8BxEXeJC50l54up7CvC8/8za7p7OtHYa/uwqwsdHJj8M6thTMf/N5EgKd6ZxE
1Qfotcdr8PAnc7zMn1dZpIRX04OG1Cxzyf98puiKfYYrlMQSk407B/OcQKa/ukiQ
lmYAlwJWYDm6IFYn++0zf6Gfx/f9Y0orBkkq+yWbHcFZAIv4h36PjCsDN56XhyHR
sZ1Xs+ST5UJfx7eBLtMX+R2ow0q8l0ukzwo4YBu8bjJeVf8vHJvygxJvR6TtQN0J
UX/HeKZSmOWs8te5/ZHgO4wxTro5A8Zbd/YsXUK1YjB0hE8s+st47UlmMgmUD5vj
bLEpz6r1hdK5TL+gBinti7tREqGJAtmTr5123gGoIzrBJwdiHEdkVn55y+TF1jYr
q+oFv31QXUMXWAEYF+EBGS+Jnf9SN9aWBu7qdU40q2wD+8WQvrFspebl8pmN0X43
B6FcCTNbTWkvz8zEVpWrlXeZ5k4tTIpKfPL9H9FQyo35wGhLQmCXMhntONo/uXUw
sV71z+nnYbpO/sSDoy3aXxQp26MRUzTo9P1jXKGCYw9zOSlwW6WEUY0DydjaPWC5
afela8lDyA939nbJQ2vzlG3wnbjstgkDJ7lnfC66eDAYwjAhYzMjfJkB5rVs8lMP
iJlCRQoKqmnhzcsG2scRoz/zQ+/OMyuUL+QlZ7lu6HpTv4CfAGLxIW1wNgYJ+ND/
TNPFTxgm/GTfxu6MFBXFYaL1FvCfGeFgWyB/p96F81BDu/MdLyTGLM4UK0Fng34T
Km4iNf2QECSBfV+ZyIGU4Z5+VNIKtQbsxE7FWI68fto100xPZkI589yWEtw7T93N
eRKD+lEvgSmCZHuAw1aj8oTcwOVXBBQDz86YOQsYNyK+QVujT4uQMRf4y2ag1K1w
WNId2VkkuyGbpaWMuvWqwXkA1RZ6DvNriA1N0HYekyUfZHgIPJ8QbYLZ5VEz6EMI
tHSXKHOIPnYHsF86PG0osEgd2CMBJAV1OGjTxfmqzsvJzjbALV7RbpS2TqrqHYUv
/NGkCVQgKjUd06HVV0DxRAlZp8eJH3i9Sv0+P2Um9rxmBnl0YKwl4mhy2gfvng5M
33CLVDE1NkdeXyRuRXV/PYE860zeh5BMrXFIXILOcfumLFRESQgaAC1s6y67T1xF
xIZbOcFomsQzEkYcJh6bkZQqmQyIMMga7Vu2zJdFEAC6yrZ6esGtjyNMlaq6v89k
lRcRAj683pgV+2jUrb5NY21Rg/80EIbCmhvAhxX3gHkon864oTNDUoENldwk8piB
jLQwMUgYNEeK/4mBOGl/rM0N4Lv75fDLejkg2AG6jMP01FEz6Ro3xIwaHS0qhaOK
b0e+c6SQsdGBOM+XALRMuu1JKCNZsGv/YUzE6uOOIrkdPGZgemTuSDe5yHBrxuKU
p0Rltnr+1WJw3YzrWJKOtDcfMRrzNN6Gyo7RwRigcKg7yXNjqGa8E5gWN7kIc0fB
dUMYlCTI5wd0vym9HvvJk+ua5BfE4tUbQcYJ39u7g6oyooGW/C+oMChM4lQfHLVM
ihhsRJ2AC/iLsq7hIN10XIWGPRWBebiwNBr/P4byJp1EN6JHQ6f/mAUqNtequcuD
oVjWR6Dt7Y3U+VBINENihFs9awTtkWn/Ww4wzASas6nRauAk+fL7t07GqSXtTcC1
GzS8vWDK5GbwqifUFIOstMCR2rJDmJMIgi97M4agEUo4v8e9imS+zJR7G86qHdMT
CpBlGvK+vkAyxDhXysI9a28REuToqIfc4TLlwmD68B1/LQKDqRrFEPuU+fmalBgX
Y4dmSXtXec/vy5uFaBCvDwdXwA77yjz9By20PL/lGUnzeo2NPHpXK9RaCfPAkzDn
kpq8ZPttH7sUVRLL9+ohvAkLrSAFOg98cUtdouVqwP3GXTmOVyCrNJ/0R9bKSF3r
Nd8oPVpWNyakkXXv6Q07fLYiyL7vqRBPnp+sgR8IZ88QZRJPDaFue/Dwexhvwg/R
GruwO5d+92Dk4qDyaHcyC2IkYVz+jSTITotoBEVkSiAfORA6CovSxvZuPzZDasmt
p0e3rCBPFdtZ6ClD82ZfTq7SnxEFNjd4KPDlNkR35l8S0dJ0OaFdo3x0jVcFDnL0
AEl0nJfkl/fCDNRhQF/alUewsByGuEV0rN/5UmWDlT93vix62fzyzkbziId6ereZ
NGiOkKwhGjtXhvGBdzb9YjKNXxM8ax8fKZrZKPBm1S8njJ9o5fPWGb3P6wDJIviA
GI6zU6csy7u8/VLe6Y7VntzEMsZ5fVTOraylomoomQNxaTcYvAfX1zTgLnE2mSuh
Zyi3M+9L3IYcoLsktn9UkQwB3rp+SQoravT8QtsunQVN+HMxuQ2vYw8/dH/Qyltl
R3qNAIrPyVYQg8B97vnguzZHvMZXYBPg8iqK170zHG2flgHZj7iP3rYFwCFUSRO/
ajX6t95ctV4/JcKNKAnOA9VQkU5CpABZB+uqo49uQoyVDv1s84BC5YhESrfe4Rty
4EKbXH6eY5mQDdrSyb+GXssOEzXj8sSI+/44LdC7zOLYTrH6BvQyfI8OPSXXqeD8
OwTDQ9mpShT1UJ9c2p5+F/nDnHxS7kWK1+RzPf1tveCzDQ1ZtrOPdXT0TLw1O9zf
G68LmYQPb140gUBlJBAxCkW0fyazc+7UR6X0RTjvzbMfi3Lh4YLez8GiOzxIxKIz
MN/S73mttd3Txz3oGo9+zs6yxiZtA8woSehwooZxYL5njDkekjeBY8H30ALnDhVg
qDzy452qRG5Gq7KF7m1D0AxMWYONoK1mc0Gi09RGYlrVaEuEBsfsZpWCmGA05ic5
x54WcJNQvOazOZUiXaaDJVyKfqAq5MPYiRVY0hVAA0FxPIEebscCqQhnlxbjturf
oCo7l/ZHBun6RRTtRpOOdvKK7GicYv9vhwGgEGEA75qUMZfrEdo1mCHPBMBti0qP
7XduoFXyk5I0xlkgUms/ojN/JgugX2OYU5upw0aj0hC2DFj8sAy5cS/1y+qFJXjZ
XXReRnjgSXiP+ir2RIV53Gyq2QFp74MDNfc7RjoTPo19GGhnWloicAmc7tyDArG2
8vUFXKMyylPT1o9d2HquEwM7t8JPaTobKI9sc02WcxrLMWwYc+2p9lJ6WMvW8/CD
7gtmIoreXC267I6Oyq6oZeb8unxjYnbaUVesPhGizX0Dx6+DBlnD7LD87xr++Chd
pQ+y2CrW3OgCDlbqapZhJ2aM/l0kpxzOmIHGUY7iQxA++y9QUhSvMF9lwoLwP99g
uPID1WMsAjO/0ixSyxoqEp7AGGOihSahmdVKBVij3hM+F+NRbABFRHn+5FhyOLoL
ethagQGmQxdEm+s4vtwjTZasjwEoHoJDpWprZbDtDyQdH+pNjgNd0TabhhEe01Ln
JzntMSxkJo4B945L2XQT148jOlyk/RzCJTv/jRwE0ZTqICYUv9oiP0//tnzOdHvq
0ZgbYgvZR5g95GanX74+uEUvUjBizpQKMDaeTkMuBuQjRy+ME9ewuQhflL4i1eqw
T0PghnqsmDZT2cXl3eZQsfe4DZDyoz8HrCXA+qUyZh4UFoO1F/yNzf8g0DqZok4b
W5ByYOGW8WSXWdxeamS0+5WsjzLJllmHAthKvll4Ul3ooBW5IcMphQjQiNemmLzr
8REOR5bqrnPF7vgL8WVGFau/v/lcm98ZV1aCw+160N4J1FpVuyeelm9aFqwMXhZQ
mqVyBv44ojt6TPaQkkrzb/F+Ujgeq8ToUjtKDoHCT2IxTWhUF8TZQCHtr538hp6m
c+Ixv8yREWa8SfKfZ6t0gyrt9P1zLbcAuP1IIzJrC/kOM2bCfYuysPduFlAHzm3P
9JeyJZVcKciKDK8yRndJLJmYgAFZaHDznyhLH+WZTu+Ha8QAr79eO/WHro3RwLNh
3EUQ/0QZ1Y1Mbh3MkdhAw0hq5VdrveQ9Mjk1l5ynlQq1nJH8MnUTElo3oHyZjsiy
ecBsPNru01BU/NnuJyeEfsn4xzjWKlCD1tOYbeUU65tq41iC3Y8qH8P9bzTau96+
mBl3rZKsqD8LosX537XLthbfhkFERn8BXxSxRbCnfqEvLXtGnGZqCB7SNEhxmhyy
Fgu4bMtUUrk2EU+sPgMM5aHMbVlFQEn71SKGtcGOorASB1/5elj548RAIqVrWyOw
d5QYVRYnUZXNsrm2e5cwnrRTwbVbV1GN23TL4U2KyPQI+GZ1bTdngmGAH6wvUJBM
0UBqUqPVyxk0vkAfUeHbeOrd0jffjIUqxHbuJCDo0+L6frOZD2wwYV6eGgQ8mWXN
V8AmdjXrr79630bbV4dRCWqxslwC7a4v4jJEZuvlgh8BVSUZ0V+mNjXdAg0B6LJT
0K7mGgU5yQEI0nxF1mRe4YZWWnMzYNETdvvpPSoPbixJtepd4DYVvT6YJ4qVB4Rw
BNzMjO2yI1qMz0O5iF6jX9w+KyBi7QkYR182AMbni1IPV+W7t2kjnhngEdThSw/J
EhWortkOPLrh9AaS4NU5cINrYWNYaW8oVak0vMcB8w59MAg65TaD99GXXZW4A3mT
SQQ+1UzG7pA0z9uzwzyjHmpxqEwGw7u+Ompar5Zc3PGo9MdRQKpL/tuprzqlNtqN
gCiYRp7m5eDmLHfY5x95Ds64BfsKfB1PJA8WTXVUCkiXjC6XeGjCTvKgjwZo5K/z
F0bXX4kWlFW5LMCuHkYLHCO3tHx6UvN2JV0+4UGpXhCBd3PTOtZUvBSfiQFu2i7K
WTfmyG4ElPbNFZCKrCoME8ai2GwRBRaXgOp7xsHIgSoeebgvEtj9d1yjFInqhbfj
3WWK493QvskCbEUyphTkocVylJIB08M3QkxGim8HStO5BJ4pE7jSUwPBtNvzalH4
yD6G3Bwrxub7nhS/WW68rKFIzh7IE08rLaBcyFu3r4Xqpy645rdk41ZMMT3Ccky6
RsuFnZ33DVSeVECAzgGQUNJBGI2EYoBu49F3Z2ki0eXHUX77luQ3hUI/GQH52Wm+
I8YUu3dFRKEGeYzaauHJd2WCLNMIqdpMzJ6haqUkhqvTRIfxkoWFV5I09tvVFTwS
WgfMN8w9vw+5qm0IlbaKXYrHP7N+/DIk2pVPEHkWQ40/rvVZcSL9I+C2pkOugvPb
xpA1JBnmiU0cEBQCUWzQgUvBDFbaBdWK28/Vx2jb8rCBn+OEP3nnk7V83F4fFpM9
8sZdC9ECMTXFCCovvW3pfIcpt6MXP5BBGR8pIpNnmD/xz5vGuKp8uAx779HOlAkO
YNyblXrGnWCzFTMW5aiYDmjhafJfAM+uZ0LtldAkfQM5GqpXoTA3Xp6GgVy3LuEj
QZjNUIHw/vWoJJH6/ZPfl+cll068QsYjPbgx3X34XA6Y3tfROcCv+t8oV+pJL04D
KnpafNypri9dZ2Ykeb5Fu40oLFJFvELkKA+J4rg9BfoO22MLte5opqdgGQNdITSf
0ZIZXSHPukOe8J6W5WueKoWD09KwhrJkgjRzhOZ4tIEmB3cAYPkv+Ysb60GAZ9Ut
OVImyPW2yYKAcpgsgEafD6zb46l776RYnXVFfvs1/msZB4eQCplBd0wpK8ccK85c
zqP0RRPKLO3RDyiFvFALY7ZFqy8Azhn9K5Nc3gdEr9L/npSnU4ocvG4CpXoc4QYv
carMmaZsjm/uqte6cjdMIeXCnHwWZw58aqx33UeqAyjwayHAwI0506sP9mRK3IKW
1GkECZ5FzCY+sO26Jxz24Pin/j59K30Rf1RUNV8k7ylvbggcGrM/YY4bFSoNNqPb
viJUuyobYdZzzkk4dZR0GJvL78fM+F/9AOO6NS2zNpe5wzT6xCY5pZLrpTFu/W33
0WagTtreRKEJQxgW7SW268Shl3z0nT2uuTpyVy3vqReGEHmKxau72+eB644aAWHT
+xLmAfy2n4HCMeeZmv0cKZROIgYjDaAi4GScKtvpxaa6AFb40uH9fEBF02bFtr9f
8DrwPZquaXsKLb3UeH5QL2klbWkjbZG6LySgjxWugpixIcPzKSAmG9gazjTACDiZ
VBidCDI1outcLcIugPEJUBTT9zsNbudamHq/IOFi7Q/O+B7Dr42FCngu7c0wnNrX
6EcSeImQv320SPLidRxBCtnnwXixmMqQ0F7V/Z6B1jRXyBo0TLHiDgONkCF5YnyY
DKESdcbL8qrZsg6skeAudv+RBLgYmzeL8OmZL+/JWX0rxaUzMu+o1TkyTZ3EfThi
xvHVlPf7BwtsvvqQic6Lcf6QqJauLwP8h4oQyJ5v2a0KdfF7poeaaUIzo+nUoOgu
70FTUviPwzffVFSjk9G77acAHGqQK9bCb62K+EPKaS3wpL+EBTu62mV1rQmc2n/s
tkxIClFbY8q3W1zD10PaHXSQGLVB9+hhs7TPLn4VAmE7XkUYWam3w1pYdMsSSGoX
mMLRnfjxGDUDbKLrISNrEH7yg8PqhAf+v53yqFG1ySdBenJwhVdfsvh7RVZ9X9nR
Avi/BMytmHNg0wMJjDq07/aPJ//cRG1pW0nKG/CHcEVeENtSjusXeEsqkAtKJOWV
3Nt35r+fM68Q8KNkE/ileWQBAnSSWMirtlrvBNvI7uKjNrDAgisL+Etq85crdYDB
eGkI00ABUywKALvTm7z0h3BdC9W0dtHa1Fv/MareQ4ABqdEXj5I/WQ0rXv/dzCjn
+AaakzUFhb5GZge3gFDc6GNPpAiqdABteXcvK/iuwoWnk/9McxCBgyF4jUmh8scc
zUwM0vSPQiBFJmcjib9jhnuLQu0QL4AyF8wn+AdOMDyoHFh4dbRFM9LsCTmbORQI
nC/E4ZS8DazzvZ9ygMLiPAJSEwUHhinRbgwCNuvsuyEChP8I4lrI/EmqnnSfqHGC
KfYKLYyGrY2pjh32EU3syOYQWekYaBO1kTP4Qmd1Ir3QHwSmynWKNuLfKdrqQ+mb
M5Y8bqnMXOajaBO5aOJgKBQ+TjWu88l8qY82b2P9dnAcF8SRya55aAmbQDRB9Elr
IuGOfdgZZZXp9IqW82AY1cPgBc48+wrGtBO0Ea9sYzcugGq60BIW1+mERn+W0bLu
3uBWWWgRIKMqOoWuSmQR0PU3TYZolz4XVg6hgoC3UQih0EmsGWnbKqxi1marx7F+
xBiJ0RQsNgu65kzu81EvUpP3bsqZvViFBjTwsxGMQDPXQxqilClXtuCMJXtnCH+K
LomEqhZH83Y1EuPu/ieiltf6jSYVMUtF9SiD4KZA3xoeUP5EJcTshtqs3R3xGp6U
RRtdVzvKMnwQ/D1XCjsduN3LXtVTY1rsPgmsXSEvwKuLjdNW54jY5APTdRxapg9Q
RydNKiB8b2R6Ns3ztoLEQx506WwpiJbap3oxW6su6f7/0+iuElIVMws3wY3x/cxj
dC3jx4o8t256WVIXrSETQQCHIU+QwzHvS+wVgnbxq2LQS3gzzLVXruC9xcQxIoiu
rkoBO68STozoCr5f57u59TrspJ3etEqyGcVCoU8+Y+HbNlsTnU4SUQL7RST6DhoR
0cFc1tUrFT4AzaP087ulUrG8qSb7NKT8trFKe9O6FDLCy89UP3RSSgKtWUUsHluF
EuwGApFqJ6oKQlyJ6vj81qqRXNhumkTjDeQ7RlAxweJBWXV8a26jqFYncsoHR116
7AORTtEsNEffWhZdF2vD5LX4ttmV0SgDLKikr/I1da+gyvDB5emxCjeCeFMVylWC
pIV0jZAopEJMvQVQ8rCJuXnZR6G8YHGSkVXrX/yByZVmjkkX87hSfuoFWKOPRg8c
dj75auDBiBsyAYyss09BBBk7HSU9wGeSyfBBkRTrpeFoD93x6fOsrU0EWnTG07i3
QJ416Lb09MxXP1VThfSxukRfJasJFeadgSfu2wZ0oFH2LmZAGvFHTdLoHyMNrVPw
d4eldmW5dZkBjU2seDNs54npm1i8xvcWM5ia5HhQTSwSn68rFkSjAUT2MzD80/qx
TqUTPD3bil0rG0zf22I0FHC/R88Hl3rh6/esx7g7hxZk5IdsdI+NdtjtoGWesbxD
rYs60OQkTFF2o/dZ4cNP2buUD/I96HRB5FKEfeP5az5bXYhLGyEtYhXZlkl0OjDE
PAO6S1K7rCvnzSAvgJbO1HszIseyDgDcAoKBGINlWVL5M9xNO2ydcDSqZ8N4JAMJ
X1hF8j1kZAG+AH9cVXAwWZ34JVPxPb9abotFsznJzMM1uPkSF6fQDZOmjhv8KBU3
VJboECRKx2KLlyebO2Gw82sXujpRLuU/xmKhRE1QYDIX24yvvUY7f5dtRkZUlN1X
3tdjuKIAANs3coc8Qh2yAta9VMjKB1EQBqm52YHaaAgGBh7qFhbyNvL8pCahUEvy
ONSfyH33obGTSp1jbJvgWMgeBuDJIXp5NKnP0FXcKbl33ZnZGsOUBB7gDGiNcmGr
GaL3ynkdE6oflklddrXVx4fsFCrfJXCxH4wO7FZDiQXYwS7Nz3bslL15T27D2DBI
FRcf5NbYP+K2tyPsTJqQh6zrudSit3hoxcvIh4Y8ddttNzKJpYPimknwDN9Ho7pU
ozd6JlHX+9stjA7Evxz7+gRYalbsSGQ8SMzEbd2YriT49Q7uEXBdnn3Z6yR8Rewq
+lppRNbQPwP/7kqKbKPM28wRNNkfgWoANeWz5/aP1tv8xPA/SgnOZNdbZjNbH3Zo
gEvabVmyKyXvrOChA67tq+sYgG7V95hl/8NmxukvXwlWItdwHDQVg3m1la0982is
Fn4EuR9HRltxnAv0iHsRZFIWVXMZ7wNnjiYnHx/fqOabmaCxECnGR0pvB3LyGEiD
3J5Qwbg+tZTQriuroldeQPd1//HIylKB5NfvyNKtoK40iPNpMkcXmnNB3nmuaqjW
YakGgDrl+/VMYcgR1Gx+pjd1CVZM9tNUcJ/HxDhANWMgKoEUsmBnDWPdG8ntciwO
b3bDe+r4/QR622mlljgIOMLlkZlyGjfV/j3EPaKUWFtiOxnrZ2qEygj0r5TedjFe
zaVv+pWxjFLYFtyPU+fqcmC/eqgaKM49l3RDS5dCH8vG4SMW6WBsyddvenCN2dMf
gWGmPvQG+rAIqLj3LApVGuA4CZYQF/xwU/r3RY71an7nNvL3nCdJlnG2CkP6Z3K9
g5K/gCTneBR+tCgpZ/3cjwIi9HF1la9RoOPBe1bE43BfFGlo54RwLJCcl5u0hK4j
NMKnxGOL4KoRC+Zx9sDoXq9D8BpABur2E2XUl8vz+HtXO+26eqNitrIU4srjLzid
0M5XCbTJshSzQCAXkO7Di/U8bVFdg9h8yAd9QoQ5r7ygD4DIkHnnJZyi7vkiwFgB
E/DZypPsUxIV767NRssPrvCy3T6um7Z3Zb4aBMWcl8pAFi0RjxhtTQArKgQuCopa
rlFleyf+4XdRUW7ijhGZo3qtCRLkuLS6kqSrdGN4bao/aarnboIF5BheNZxl1xuf
/ALYqGL6y8ge6qAPOPgVMuOP1Z7cavWoST+ACJ7dwoK7jJpqkz0Ro+rQjb+WiWyA
seQgFd+FV2QlGRB9PqNZx+YX8C1dixu1vf+cqKd0VwG/7f/hsdaoV28VySfDiaGZ
H+GXmpkxtNs8aHgUC1440qx61Lq+8ZbNMU7ejcIwHqgC8q8m/FyX5PryJD/uaVJ8
f7E/k6TvXxnqHi6gbwQgnea89mDZALSoGTzhMASmIQBURE4+1y8MszvYOhX3nFF8
2eWl+YV5KZPUu5NIzGLOlBuWPoknsS41U9h8+gBdWDBOD9Em+XCXpZerZ0RCsQm4
ZaeMwH8ZDotX9IJX3mCQDuyWqJyITrbCGSlsQcH9G8BU5QiO0+Q9diy86b79fdUB
gOZf13EKEHEj9aVstjB0K3bX7lmei1LwDYqlbTJi9jiuIQfxw7cXwHMwWlpiK5ep
j0oRtZ+6N/aLPYc2LYFMxYm+8vqRU7GNV/CofJICmMst/STnA5RX46o0ewFA52TX
ovC6hp/lOUXHMeBydWRD++9wsn+JZh5Q19EJr0Z5q3tS+OSqgFOivTeCeNqSWDPz
+PXXU8LLKf0Dhv616vtzV+j+cvNPUgJ2sa2Tmg8t1T+UBi17e5Vau/Kb+ngwE2/f
gKNlFufCwM/wmVJpbrD/UzjzvSrGXv7W54gx6T6c+lnJoQHjjpMt2Hj0ObdBTktb
uhJK4Z582csqhAdBjQdcMP3nsj7/NCCByhpFUqTb+NVA75yAznXallvmK8siUK3j
9JKz5ot9J9b57LZgcMcKSFb9cdWGvnHNnx9Yn6hvFBvbybXGFdtAHm1PoLXInnBu
5HtMS9LC+gzqeuOb6fVUtyO1KJwyRfdXgSv+09cnETMjid6rgkktdvnV1jpOBvXh
4djjBP6/QNGLKc0/LUchmtJ50PA3zj7DcIzbD3TTeH6LbR9HZE7DecAh0Wd87ujt
XfwpP0THi6jj9qDXB+5DHgiZyAJ9xZcDQSk5bpcbxj+5S1P7ig8IiCclSUgFa7NO
M3ij2wuc4tIREIZt17cmocQAEcjORMlEjo/kPuZWPP4ocK00mauyra+bbRjq4tUy
IiA4T4ME0h6Q/jnpzR98JGrkGOTSuWRySsaOrt4wN8Z9ggHUbddmRt1aFw7AVziM
96l8fm82gGjnGR107AC2HjeBptQx6DRCSESN/HDTvwdIPV9Bv3geBHdQCSCMttuX
1RHcOXiIrM+eVwz0WqWly/5cv9Cew7GshI6AhJLQT5JNjCBJtslnrgBXxaJg/igL
mb4uKYFU6rkAhcJXAKKqBCYoV+U8AINwC35MSe1xkadPodOsAapEcwlXIJEvuXw7
b+Qou823BrR21tew9n3tyOLI9I7QzUecsS6ylrQtH6joGlW/DdaenMoV7Uqf/tLC
DGVGxSFpJ55dyJatFCuVvcwWJaNAVh+qL8zI3H70eGT7sfF2gEX7T6JB4UgQ2NHV
D/zSgcWu8fKb2xH2V9ptT+wQQkn1jszbjrQFXQbKJoI4DsvN+QEsmiDaRa/iiRND
wXgVtJWc/uISrcabvmWAO4AxGB8rpzu/YIxoGwyu5QACmEFxNmFrJZeLSn8FxCg2
Vi3ohjlXyUnIlw+5Qu2aVE94OEWctJXGClr4is11oHDq3S0zGSP5VGM7rOg8snrq
Kk+s1syOoxa+jjhY+N/KAg1khnH+0krWrmcofTOW8F03N9/zak/mpGkO+ddTojV4
G2X9Lw+7kRgt4DNNhFbjPH8M5kkTPlpehO5XLbYQvI2uryzTswdNadG3MYqaOSOB
jaqXnjzhf9Aq9ycObvH6Fabn9UnRKLxzuXBW7CAmPTr9NmAbyxEZHbyyTX8KKUBy
xGTVHAGdEjqL6BiMlr5CMtnHGQ4T4jbsrUPl9qz58LYk3XxDNTz+sufPnw1oNIAy
zwDJwxiVaQR01cIPrxfeWrkQ+qrk99teOLoq/Foe3LmBgqj1UE4VSxa8RLoAVSyJ
WavkdEobAKTDiPQHDKuiEC+Me+jgZhds7/zI0PFR3ZLIXMmy0SdqVomR/BfwC+yb
wWgV+K7BoNfNz+SzL3qbRpgrmxplXdzT87QOdqAATXiQbzOpEUEdzvM7TQ/sQ0Fr
J1TNho0iYu4sSKOAaJubrnxPf2Rz0VYcXMhS2//AMtgv5RMpyqceWJpLgffeP0il
PAysZVEIoZFCdxPYg1Hsrm2t0YhTDzT2EwGNPmyR0huY7QhUYj2omtJ19eVvAHnu
GznuUXbJ51NK+X7Z74sWCZYdJji2bvzEzhuElERSmV69+vVFf3GN7UdIeKi7Kx1Q
7z9GVjuJn/VFbTQsuaT1orITNEhGEJmuMEX9RcNuA1BKzqIvBnC3oxf58yEjlBP9
WM6XF8395PR+dP9xCMmUDEyiboO3bwEA8XklCRgH4ST25OAtOWQWdegpckiYuC3L
wnIcGaop9o23uSdc7L0RJDfmxD1PXwlheTpkFWpaYgk3y5ejpLiLRhmaCjSy5ths
bajww5SmTeJqHbGSc8mzMQ+OtjBiQiOcPuvfbw5qwxLPbbkhH2ov29D+QSMogSt3
gMz1UkjprPOIoQ/gL8bScXn+AKUkGnIxBuWR4Z/4W2V83IHyQsB2jqzoubGLYyGl
v6hBeykqdhnGMCJ+NFVVqAj5Ck+VmvAJqGSNKLjVuzVArn6sUgOPdsLLZZ+Nt8sH
FMh15jYdhtkIEAFZvdl8bcc5vQsPQxYALsyNyikZgzs6GNPZJbNnUdDc6Gvwy/QQ
btXH7lQ18pb5EyHFIids73sToHV5z8MCwn0OzrkzTE0xHcNk2T6WOGF57cM52KBM
YMK5DUUrUU0vHTzw8sOMp3S7fRIYhkxC6YRMifzkjYf5TnYosL5Lb8RR4wGf0gHP
2cQsoW+Ky/t9hvmz4bd4q/OCYn7zsyZFBLJJumLHqbUDz3hBORG7kzCz1VYC+Y7j
7WEANykcb+28qc6nIaD/11V5o43j3hQ6TUx0iTLiLV63ixlRaRbcaF4juTGDjzVf
Bb+NcaVrq2GOysTzEvSNhMJvFlzsbLmgr7evsF1Zlnlm8IaFqWby8ns174fzuP7x
ceSyAmsu5SFJTpofQRx6QrDAABFtEpR/udfU2mitlxQIwdGzoPjL84Q3nJd4Xvq1
YOXcNUktFAs0W6wxNVqiOwcgHBEOLBd/gXmj2wXT3OCotAojZbTPXv0UU89QWh2o
oH/pkpcJDXp/RdIMNgH4ua2btGLw3ciz+4JyrIuvTxbPwc1yF5aCtIhO0u/Ikkxz
weLPGIkZnw5d7jyc8zbHsLD14eMwV/cKDv4MR2vaXjY7eyXy9ugUytV51gCz79jn
xUVlgyXRTZnHMnhijll+AoX09M5OPYPBQDCrkHAIkU75w2p1PtDV5oieYhIAUhZL
jlxcbSWX51hPSmYiJ+zHiTHXoouCC8jjYuvF3dpqTv4EuwuHqoz3q41SKDi0CK73
e732Q+XOSyrAhH+SdtpvLvCZfMmINwIo3vAtsexOAklI+X4xiqvTv9eEg6kvQdha
TDtEY8jChRgFs3ER1uSFyVbScYf+Yk8iJRPQUrwyB6FM5B1bupnzI1hocIgLvMiK
xbDt+gTWzFAP7a7FD8qTEZCo6lwbuRMari7k6Ix8VdGu1juoJ0I7GCYEfBTN1AlI
ewzmerW8XtTfC1dcCHlB0T879ZwOjIODgYJMH38EPWL8H1ZdhSedFjfSPN4ljgML
WLxlshLcOQ5UOMo4kcH1sp0oEKkrOx9rTqtgkpUnjj9/PxD/kFNZI1XPJftT84hg
61WHRBF/sRetrAM5DPWIhY+rUS88mIXzSbLgscuWn8P7YXlBfzljs/UXkx4cQuwK
EuRyLvCG8xpSUi57PBaAKuOUqt8TV5NvBF8wAE70w4wW7jngGk8i+0qI9ROTFPOK
nw+Rc7nMRsQBa44cagkotlj0Cw44v/NnXWzztUJSIIX/sKthTDmJ7LAvEFGQ/iFv
BWh45DJzNyoEa8aqs+hiVJJXQRR7GZXJBgC3WwgB8DntZK9wmLa7NT79hI4djtVs
tWXEiV3sDaYzVwIJX7xI867fo7SC6mYvM7SeooJGV8D23UqEBXAW/fXY0yK00OVs
cams+xiLHI20qa0ZP607Z1+AbJQTK8DqDXdlLz1MAD5flbHjlmcdIV0UF7Zju1WZ
p7vTk4Eb1sPm45M9FsH2vt+unqhSgigt9qSUZ6F9swEk0kIJng7batWOiNN3su9/
m58efleIqwbqUCHjznRyAi+hEEf8omdCebgEug451ViNyQrwDtPGU3JQQ7bg5oxa
mJ7xf0YTJRDQLHeeWRYVqJ4sXHiGnI9x/bPx673AJzDTFD5Q3jmFzoWYJsRpcZz0
wBHzHOjeo1RByjJ0Ev5PZ2hlDhhU6c4wrIk/NEpIGOKSfTmtIXknok100gr31zkF
FzFvJ9Pt6vfNqQ8+KrBvsFSmeMJwjgf6wWh73SXa8M7pvlARiJ+widnBThFjZ6S0
5H+4/oRNxsaPe6j8dO9BFN7J+BD1e7bt6K0+ya+YFhWObns1foXvuMycCMnSSVyk
MOfbaJ3QUrFiu/FWBB/L0rhEJGyalBIwGB2spECdfiG65r5tJlRYLnenBOrLYvLw
GwAbcf+NaQpxQCdjoVpQ5O+ZUSrYs5LG0iMHhpjQ87JyHBG0Xpf9WQ+rsvpW+HcN
DwqcMoesBTbpIY9Jt8bWN4jk07+PvSlezN8NqjFoeeG3vwUudW+nJvzWERPm+2Py
aU9Eq9Kf2OTwxXzGBxSI5I7CRs4Jujz/mUl54eWHgS+n8aHm6/e2D1DM6ErnlmVP
Jg2qwRP8YgXcpl6i2KFYfenDAFuLEWqyKfyo3j2OjBPMQF1rfxftEzEHwBp0J7sk
zg0yihitmJCdD0PFG9EiR82ynsQ41Z4Iu7OwDl3isoH2HETPBGSO3xMbO7B2y5Go
KSlWp+LqKODFIpGflnWl8HQ3uQY5gkqLJlRGHT4IYQz3RdGdsD3NkW3/sYJfUxom
ZoGBU3P01tBjwH4gxSOLTEqtMTsnO4Wq92b+1V7mRRf4xOWPxOyHGaMhxp0+IkuC
of9E18FcbGy4SqKFBM4eWG8pI2p2rI6MMVv2mBIfTnNJu7o15m4rrH/Z7WwWkvno
GS0xOvVrCV4VPcnyRvoLAItox36i5z9+IFBjG8yIROWz19CnAN0GnFe/el16c0oE
UPXFiwRr8Ft6B2K7xKqxtAI4PBp8d8tPOcpy7vqZrsBu1+MxJ2mMfPGLc0P8w/gB
asUaM+OFvGysLGJZMOumpKeFKJRks0eKXWlN+Q/4YLmYStGod1na/5OtAbtDx2if
1X67tubjjllJk0QjrszrB3KjEMqwD6dJ03+NcthrBgAbCmF+SW/DQfHr/tg8aDAy
nNpEFyhSDWoAQZKAM0N2NwVIu1g2NQtteiyHG/fqnosuPIdweMXvQsTMdYSPs4KY
w2p54bzmIYOjVvGov5ImCHReiAGWEuVoQ/eGc25J/e3Af52sa81+T7P50QO6B9TQ
iV6lLnvLz2yQMmiF4LiV+Ag5ndSw6rRwHFzEiQi9Is7UkYFrAjLrqMgN5AU0chh4
jRWVAw46EJkKWwdI4DWTXDy+gyuHpQKZTvTbbFhdmtbSCytBzvPo869gyPQIKp+y
X6t8Qc05bOdza9siKfCK0Rj0KTCRUbRaSAWV3NQJu0bmc7LNxIWxUvPuPuj/Tfpy
gYEY7EUMnawJOh63pToPAAFQib85kpeqLfi0fuWUjWXS1mBdw69A96l1xDAS+g2X
OWSc9DNrIdyqZvVubcEE2CLeHjfLuA8X1yl3YmDGz2a6ZepDdpJ8FRhY+ZLrNHMo
XCYfA8u38M1dKyGmTI8NY2lD+4txkIGdFp1RNuDcNLbj3N+a/yn+TyBIiJwRDvNw
87ttPBUWQ4LyvDW/vpeWX3W8mwa7tLsqrsyCAbyfCntXE3/txdYcguBjLFR4umNs
hpv+vCnaA+FjO1DY7man49yyGuPU3ikoGuFRn7zfwvr3K/8nJkUg6KyyJ8bhKkP2
4y8cR8+Zuw1RSfyw5FuD0UzOe4HSHDmZmL+wcQrn7mQ287xoAT2VrL6rQuZIwduC
wNHwDo4HhHREul7ZDf4jdVjlbq9cJ799EuvzXqf1ULiBYT9MFiU5fu4te/osLWv2
nfK5r0w5LRLU1Q6/GtOyeJftJbOg+1Q3RYaqtoIWVCWURj0NHJHg6/5kB65Cu/RM
9Tcex3WPFRJlg+B4iSCd3LMo8AxWevFmRHMQ4rjAZDUbILqxLphx2ZBngeKiszip
r9fYu8mYFPlIeg7C0Zcsjcd/yD0tj4o/I94IsjJ423Ofi4mrzQaKyUAQpJ6WH87j
PT8fpOW8k2TUUVza3JGAfuoKL91uk6dsF90hP6Hxtx3ZmdZoUwIj6eU4LHzZdGp0
q76A+wiZ5Xx/13WxuSnlD82UsW4Gupxz2hJrAqvCBSPq1xFzLJOsqt544U1phr8L
3UvD2UQA1sMBPATHHDXt+JZn3UGI8HElS2eP3ESUK+e4DO3SY3OWqroQIhiOamz/
Z8u/unwEhPMBExma6GuKdQuppafe33R7FtzY7YtC8dMeUHPE0vlZXFQlX/Bp1w+m
jvktKMIJclCe/6/Ok+CoZAq0YzfHnoSr5MaFF7zSxRFHTLIkg0vUCo4PT0t610Df
H7LmIr0JVRUgBe2MH/fP28+bWd2ElQN46B3x8+jxiT4RvuMSLzshUYQNCaxN7Gi7
UOqOZL2Djl9U4wYlc1yRuRUw6h1s1wqzucHe0nBNGLBbUMF9iNrvdf5RDIfOrn3C
hEaj7jizwa8xcfdpd/YocJQJnGVRYLPmfTRzBBA/3bjeGUe78Jd5y72QIl+pkil6
kpQ0gdP/LCxncFFc0cjZ9mJFGoTteCigXcdb9YXf0Xm4f6vhCGT0mgiDlsMQVIch
3ROT0Yk5ISzooY1iwdzPMCpotxfpkKE+detPnXRKD9IqT7YQRZODBtlTt7nVy/nK
oZYBV+1FHrWyKG06pr9o/izPFQhYmmQbA3ms5Lw/FNWDnhi2hES1bnPQGgANaRuk
IhvIuwe8xKpvtVXSAXZsH7SfpRTqV3BVK0sN3bA2VxDwWJwqK+pOdJJNLAFrArZ5
kTHao0P7yPKE9eZ0ovHLFrXMJ0yMkTSdyXX856PdTYWFjchkItBH4zyIz2W2abJE
+0fC63KMvP3PAIeDbP7TBbhmWZ4qrcOImkeAzjmjAO6oH5K/HZP62e+LJ9V5cj7y
+6Lwk7VqHmMmJ8fQ5RZkpnD0stbHAwbeJC/ldt4CVT2TfqjtFfjtZRk9m8a3VjqG
al1EN/YkDiNFXTsxRC7EFhJxhVe9eZMOqMnfnvasqHD8QoDsBfaGnOZ/uNXxtAlk
mlugBJ34CbMtHOAIyqDQ918HzPlLb1SdPsIp469Rx+3CrKamBkGdmoKVZtEo78bs
a4azi70IxFi+FeRx+7Ti1YV4zTo2cVvdAVDpZ9GQdk/YMv+1Rm53HrKntTzEDJiE
s4iORi1mqUETVCrKQgdefLx+I+kORXOtQBkqq7SRT25h+5ohmOFY14tZpRwOV/Jr
cB2x7zWMFgyAaDWcfbDZJXjgDbBx3Q+WAgOQS0Pi1ZGEnfPw7syJp6RpUbRgifC9
RUYioctgTW8ROXvFoVnrynGkK9lt4v/55ZIXLytjwcmqUaFCqNR+CmyY2GlEnq7J
ZqGaXxWdweBW7+O10+hgg0OeiZMpd0/XIfbHjynJE2rSXPcPEb/DnWM9fEFDH6IZ
cqlg5+iHUjzhqrBSPX6reM3Z/PpqwGLxyTmGV/oqf9aLhAaR2KNSi/7GqAOfbVSp
UC360yE6swc41fuRL5GFPajvmaX+KD5j18XfDYLp+Y9iIYbSj6w3NUzpMatc9nrv
CR2dcpaF7m0sn3CvkekDtUlhC1+zQnaYmawlVw+AuI6s96/Cki72MOuQSHSjpSQF
P+E6xAlZIaMeXUThPdFcxoayym7QKZ7mBff7QN6VLi79vdtoWEpJCBNKOjtCqeLD
dKmJI7AK5DS2fXuD+h/zdFN5/BPWjOeap4CmD0HI3yHZIwpG3DxaWCSbH5au/Ltv
kI3BlFdzBsPo8bZI6rI9VyRACemt+DTL7jzgkFeJQK7eFnyHx2YTmsiQ+NAxoRlZ
jXwort4yPLggLxQXzn9GdERtiAuqWFgM3bbhffhEp+gjx/YhrrOLKcGMToM2bgdL
KRc2mypTxthK1sifPYKdKoSpajcI3M2z/Hi9x990leFG6DHBr3Q4MS/UhbXY1NNo
ISqibPcrJx2Ga3ZWOHLgXPD1F2dsy9LqVAUI1hUt45MOClCupxJ+YtcyLQhVDej8
pUyRVqm+7/08NYSV/ynR+k2ZVtLjKFmP02hP+HlbXPiwABO2VP3euXEt8VHZ4c9V
cA+fuevEeva7kXyTgMo6VFXZiPcBs/vjiZaxiQZxkyhzE145Cb7nRkIE4bzl5szW
qNMbG00ieVHUAosurIizSrZZH+Oww3NuQvvPTkXrTqAkhnSYCzden3zKIhOunqQM
SigJ9poz53J42VvXOAWvakKCW649QT2sweAuwzayGllZ6nTtt+OZGs/QAbYdA2WM
NNkSEojMg1Nt5RaERF9H4YD77JyVP/mhT8MZuHiuouZBRzCfxI9SD1HKQI/GxHPF
X3T5ivuDT19I4wgPks1tC7E+eWCccPU3VoS6lwtNdB44ayPjNVcEMpsHbXJqxSt+
yr2dL3Nv7DYGT5UdqY58XBp1alhAA6zoysrQ8CUAnjMpFJNjIDzRgzn40ardIrRh
WYuH2dqgygNoqV5DlnI4aJuETkGsWv9EB+Fb82FxTsuzFBCAD0va0Z3vkpZ/UaBX
H464U4LvWEmD8jQJtF8DauyK47wkLkjPdskPgBr5Dbz/9SwvRz8u+uCr1fi25xDy
y42VjcAWQD246zDhi8xzTY68tHliWoPkisrdCRdwRFeZgfqg7xBTwbnDjPmOcDx4
xM6rr/dhO/2gLU5r+M3m9kgKliIZRT8VSdqWEQ8PWmuO/6x+m9W06tzrUEYGTSE8
TdFNIUWOrYvwlfCpv9EIgplmY2jc9SsAVlJfPpDSj9MBzUHdztc36XcVCAccXi5I
EisOafbxGN2Tl1y1jAp9GiDrtiM7OcGB4++3E26vwsXZv/CUgyxDuck0WM3/lFCM
xhhVLi8xo86x8dhrLDQkXMjh9QDXakTUb0UXY1Bk/Sw1+/+vKTKlDryjwP0fnuGg
qlaaD9KEOAXQ2L85AGs6pXQfy0MZAR2g82BmeYXe3zVK+0cI+YmYbBJ7+HKgynzN
SJa3XTt19CzLnrHLErMuU+rOvqevxKD0sZ+6SBE2njOhTWaewU+SCLVGypxcqq1o
GHWkTk+lnJDy9yuSkNZP/1yywCJ6xdlMtHx6lgb4eAKcPCuQAnxCmwQ4N+PaJ6HU
AbOspElNqxC8f2ljP2wkjqvIULt3mj+llm+5vNvfupsaXbG7K+2+sgmgUad0ovEZ
pPASEFf1jwCUNmqHSE0XQTvI0uIIc3VOZFL3WaIIvclD2DOnAXwzMC75nehtpBqQ
A8Gy8xZRMNCEdQ480Sj+QBAR/VGKOGJPlppdvLb3PESufbNLv1JCcmacZdGEUUkN
IYtNuK3X3tYL/COGsDqcN2sabHQ3VuutqbodLK/qUnwMDeQJ560QkFfm7eCdvhJo
i/4+Y0PqewidG4Ir2llzt6MbsuUxVGEOeBZJi3IH30H/mC90TO/vSy81fXVofHmi
OiYvqurXqA0zOLovdrOhczGC0pc79epZ+KfmqwmnIlTzw6+ooKytZweQ5+D50XJ5
b4OVRhxYG5OqZvEzKvRM2buToOTO1CDCVXk38pkj4uCZxDTmjf863lI5Fw4iCOFo
k12TFc/m3kk6Z9zSUAENcQetSWZU6+MlmoMAGxGDmlpP8XD41CckT5NOpF6EyVrg
MLYl3F75l5EQ8TXsGr+L4x9R8vVmSwxa+3PhPkcSGGjaK5saxAOPCEOQ1yYH77xk
+4MZmRbbjLsYcyhMCAmCul1Ht6e52jslN8uO3lglIQMIeGsPozaJpn1AeBtGzouI
xpEaa02XYSF6vcKW9LWGDuj2hRDwf8SH6cS2ISco2OUPA9tutS5s+RRMZfh9wQkN
5Yz7TB1J/rR56AMXJc5XDMQV9UTYOMXF9JrN8Gc8wW9GyRJnlCAwNYWb7ypG1s/v
8J3ljcQJbJOOqBKYtIphxGZMRWbatf1795Aa388jqUJ6w1HNxkKrYQ6XZHDIW4mW
XpXUf8ImzZEX747mwQl0tFNvNOr/wJnNLUXGpMKvdLUjYl3+l/Y+YffNsSfrx7AZ
DQkxjXpHhB77/tdviN2GXa5q/8p0SkB1cXt3CvPO/uXaWs2ay+08liTXBChfAneG
KHsOyvaYg3+trbh4yiSajIpkaEZCV96jTmlRoNvU24wUcFy4JVK/zvnYvnT8h2xM
H6nvYSKOyxu1vQDbypjx0LFJazP8+VhQXhcYX8SrRSBNiEwfNNzeIo95O4a9d4ha
mgGJetgI+oiZlA3WEGRYgGTWwiKEOrKDAffv12L+6D3Kr2trzZ7MaQIBuRYPfjPc
5AsuuVWF5HRYkd5PGhuqxUR5aOfLN95nInHuK3wJ/BtW6lnns2q4XEOeWeM8erBp
CnVmcYmWSqOHvkYwy9t9VWORBsrOn0svno/Z9iML5rDDMFaeS9f/irK8ahtsaN2j
yigjtZP91Gy0aF9URKBvm7AabXYnWn+2S9eNlQIkCaowFj42wna+IMinYzpyy5yK
UjE4eZesTuQL4/MgB2hxIPJnkiyHvbBOm5eeUs9MJQHwFhnunvoJJ8uzgUmj3/h2
E7HRxydnjfo0gZ/ZYdI4MHqp5E0GoRkkgGwfEEjtjEnmTgHnwdzWBadJ0M9ZL7FF
du0BpfMsZayjfx4gKLUaitY8b1XciLy26uCmTy4aNsZPJALeOPsOKw9GqOXqS8cI
PioOEYLTu7T5lfvZ390g2a2gS25/nuwVbcJ7JpYQa/3NLEbD2J8nCSAxyct89gqK
bQX57Hr9yfEFwCvGu0PRNnl5M139sq14oR6l+33tWVTFm81UzeAj6IrfOwWBSjVK
YThx1r95/NuPn8JpZih/hmfsuxlREZyp6ots8DXuIUVGbIwSSw4wNmxHTjC3P11L
8UvFIkskYqH948pu2Wl+sCaFPDZMOhbjM82ffdr/no+kP7Io0vzIN9sdQ9WfNY97
fuoeyq52u9p9QuDurkT6ID0ThfaP8CfDcA0yzP99oWd2/rz5z+B8ODAcc8kJWvnZ
T9TSe7xg/oJavdFgJd4PvPa/iTnDCrzii46L6HTe9lzgi6uWKe3lEyIJqDSSVOE+
KexoIzdUaznlnmIg0S5wrz94cC4gcS4Tgnqc6KU0c6zup20CTd2nPUzgjauM0uLm
7mXUm6wL2+6mVlyjXd6K2MUzs8wa78ykJ+Kbnp9RL9yAfC5gPbbf33poy5PqjAa+
4EQJJihRkByDnOEgUuEo5O+A4KtHMn759+TkaKf6tF5kzEUpBEpgrOMOhLs6OgRo
QsIb2drJ4X3tseXtRHxFayxmUfdzUbgbwxFLF+DhU5Jx/aqFcD3GasDoaIsXiI1g
VYobzFah9WAtBuNNs2Dg1AKLhuQ4kIW8byjkhUqaA+5o/IVWnJuiSt6DUBE+7EsD
rH8RxfZeLdSp9nEk2EUpzEUA9AWSmNcyplityfZ/O33WqZqTNuCrT+LbGfb7K9S7
jRocRLHA0E7o252/AUz83emkSpLQRDUcOXxiHNwymtwOgw285S3Ec38tKhg9vl9B
uDQ/ROZHLSrpj+9+hlOPDx8Znaa0PObHW8nrqs0GO9J11PKQdytK8pDS2I46wlgY
m9HsGQEe4dhANu0DOpOOUMUgG/QhLjj6cSy2sR4jk5F6H7MmmXfbH3XEGrcZZ6Zw
uB12upKuvyPWMj/N3nH4+fQhuYlDjKWpNEP41qtW0jSqXFiVtYUAArvCr1JupVcF
JXIAI7RiZTWioSg9II6/OGC/TwVcSncJGt9TFDkt5NFbPPr2MytRcxp4npIQpjGO
HlH4KjpdIssF5t3yc++HsxFEIiCgIKqotnte7gm1K6O3A49T7ApGzZJeQZZ3/NDI
Exg8+Jemaz7/B3japZd7E/JVFWEw23uaNgLRMca0xfh28YrWmN3pVOXXAzHAVDNI
VLRbrQK+wODaHN2HxqhZhSRKqjizpFUsTLbSb8r2LuN9VJptrgO2LY/NEUhD7fxZ
EckZMtqyl3j1Q3Zze5OIp4lSPFiiJuGOHsVbuBBFG5LTwWVWWonbZUunAYe4V1W8
Zv/fME7KD9U+AAA0wk5bB8e0ADO6RILj8Ag+5LfJzpGJh03txiY4yvMNCahDffhZ
6nXQ9MbPazkYgezzxikwBAj9rt/pGYNiVpUsA7Qp7B4RstE18ljfHsIDEa+2+qIJ
bJn4ZzZNAplTjnxuUd74jDdXhyNH4oNGiubIND8WHIKLq4/Qb8xS0JnBQut9Yphb
FKFBhffPT40j4w7R48gAGT84K4vgEg8hdPm1bcaSWStz+7lng7Vhbm+c0a1PDMwo
HDkITYr6lmYMSyigoYqe2bGyWBP5QO634CkR1P7VhDPy2j8fCpUX87+3w+zAOleE
S37g5tiRD3xsHt1HacMas+E2stgQKjEfWWl45Qxb3LvyOZB2LV9xfCZUDHmD0vvB
6Y5AZ0kpFUwl/rSewx0hZ8v2URq3UF42TpnGR6CG9PJyKPRJOqMybpVgQpuajfY9
W411GY13g4NmfunsG2AGyMeLV+PlEK6nDKgIc+FRoDcAiwpp3nNEcD8Am2Mx4B2C
JjGjFfacr0zVXHBC+iPXmQ34r0duyEv1qbzMBRc2OoZZKnfCFXXT1W0IgIZ1dBsq
D1hl8W1AiElx1dsHnlXUs0PutC0Y6QNgW+H/35Qu+fYjGhgHMhjTc3Bm0EDZwslV
jdgzF1alSKac7vb9m17N/k1uBgVUlKHgxxGwOWQU0LlnNS3l2APCCzZn9dOlbGU6
VC1nRmlxHNZDBkdrFF8+DN7yaknMvYyRPxQcKCz8g0GUf0cyt7d/y9+bGXp2nx/Y
MCPTLeW4W3w9EH98+N9mnRtclEsbCydlkW0TobVXaUugyT+DqROXoDmTC85avGlG
EurrKG1j0PczWQccAjkTxgYQikDroZhsyG/H4iVzlFakAwFfl51P6I4HLaebtT2D
gTVC8YLCHC8aDy2oPm7TDRztsF9ElbkhG4FR257waXgXkahqL+evVJXjNJYrA5Gj
ZuRbL0IrV77BDYRxwMP7D63RWeXdAtS/jfack++en6THYk/Rj/MkGXGFBntl0tlR
7YbAwB3cZAIiWDaL+O9Fm6AYcd1fEGLwjeSWS+WaBbJzp/aZTV2kvHACL5i62C4h
du2MloDLX6JxqmXczzt3HhF1HRBbFLtPjlwlnL/2rEBkc6rriosKpz1N1cetUF73
zF2qi8qQvRNS7iLz3yMXWxBo3QHb7aZzFn+KM1w4DuuLKcGghFyD80A+k52Hv6dF
xnSeHyMIWsOhiztMF28WqD0wHGIBfMt7koM/ZwaEreKKLlZfTJ8l4QzugGWItNEw
/4ckecQDWEdwYpZ5A9Tf+0jQYOTWPZAUuaJp+K3/wj3+ZRZRjvf/9fsaR36enIyx
ZdzyLX4FcOa+VN+aITgThX19zmOMmiUVkas/6EOmrTu1DfiAiqmSuG6pOeSonkRz
4c9g8lc0s6fgIE4++EO42QjdT+6lgOimZ43xgoezTgH29tWlg/SQxblp8/YGTTks
K8fKiYcjNz2rte6pb5MgTrWDMvWzWs4ycZWWBbuGUShokirWyBDf3Uu4ba9PFAwI
Eq47JM1GMSvvjTPqfgHLmviQfendPT1L4VMj42OhTa9o5UIw4RmfJXQNJAgFvQDi
YXbi0MN6y1icgkPgTuRlnCnZi5b+y1ep+J5Fb+Dmr6iLiJeyRDWoGFsZ3a4GDIh5
tdqX3O4s3REEgVZnb1KiVCWjlJWZ28xtBaFp7R4ddjNRDt+2Csab/QTUCWD/rAWm
i1JpPGGAPKngs4RnP8LcJoT7I1cXxtNw4uoZQXG1zQ9c3Y+UZElKOnGyOwxwYg8l
YsaMpdopZyltfvUH7RR+8ViZLwUUOak9ALFdGovw72WlJf2Q5iai1eiryuNhmWdY
acNXJZLse9H4b28AKSD8uautStbs6Ktb56kCNlLx+MGyvClExa+RpTLOFike3Iz0
/8qBncb4f8fpBCZeB/KeDn5rVcFyy5l2LURUz9x5989XKdqEVcuxkktdXgN1EVN7
gh51+tmXVVDhkFo+QXJv2iKcLLyEeE8J+S87a80xfAsFi04GsFBVUFQB8HhDgKbW
Qnvpdnmi889MfV5TnyFgLEBgnIKquEz8lqjMiwrOOjhrNA6SLzVdo5AEK0cLqg7+
HOQgVUGdX9teL74DlkB+jdqdsf400n25ftEmB4Pkp9fzx8ax0J8zbfKOFqDyx8EV
irP3tlHSOAdjrB8BG242/u9m/F4hgcqt3Of/rb8U+7NKa/XQheZ15KUiMkoUG1pN
husnILFivzCvzBkO4Y2uEsInuxD2IDo3Pzx06kGaVhZNaXAcC4Mytx33lM8Q77H9
ZUBQ7Z/K9dnEjX8fR8+NwQ4rAJqOyCZ5jI07TgIk1l5u0HAI+hswqkWcfO7fK1wf
nVFNBFS1Enz2KsQU0623ymtxSgdbW/MDstzDPwGf06E1iah0oh2QTnfxdjJoZTrz
HZhJkW9NZH2ypjwfWJrmFU5BmknXXE2DxADYZpqtOU0HjYx2xwpQHPiV6+YjnMh5
N4XDs6RBdB3HyzLKq1cOl9g68uiy/QWhLK8HySVeO/oubBeyXaDMz6CA4WrdeUXR
eegfoEEEd/e2lE3xYfVhMabkcH/5dvfAACAT6hfy3X3T+Fgoyi4akvYBU0rUI16r
BhovdJuWd2Qw5UZ7d6SEM7peSjc9vxVzs04ZnZgLdEuQzVw8e2fGwuEH74LoiZ1p
RA8snEo9axhbDHtJEjcanBBDHDCu1ZHXoVb/lP8D7jlLkhNTlor19FNWn76HN+bL
18PqIRhv2L8oW7DfNIR2acidkA+e/3QpBnHe/0Pt0e2Jb1xPc8MnVlYrtThfcCxT
KaDtcOCnWtQdg3P3Y2/DVGrNxBsgfy4L/OJWoXF4+XZ3nVE2Bqa2yHC8ecXnb4oW
yhTxUfV1DIMdtucxY2O/+IKFYcqobKWS7IGSUmo6fJHw8Oubtvg4qDYUiILdOHgV
HTFc2VVHczMJqWnnaeXM29mmMRaYJn+ado7WuuyFnpkRI8OckA8u5adpTR/W1aNn
EfTgGJgxHnWlNNy8meClMe6ogAn9KaMbag6Fa+J/XQ0+pQ3axZgeXWrE9NmAXtdo
F9QB5pqEz9PxYD3oPy49PsdoUDBcnaWCX4QBeZFFepxeDo0ziTAbsqPiErmKvHV5
jCxWzFXu5N/9m2hfGgzdhXG4HYQJyE05k1NLug4U1WNWlcQ6uAG5xX9xT+G7w6N+
zwJh1YwlBiqrQBcW50pTsj/Hb51z0GQDjjXcvkAcPp4wSJYFo4QSLOkCZiM5YS26
H0uFrNb+DULoLK4BcyqWsJS7PAYHA1/MDq2PiSaa8VPrbjX63OIMT3elnRmSKZfK
b37CV4vC9gHIpZS08uUGaEJAJVr3Shw1bO56AzEz/myhTbszr0ez4L8e5qu/Ac6t
uTna22ZJHDoA2a6mtxRdPw+e4jMHzSHjtNNtl0ZJ8UAgZaTif9F9oJfgMyJIXM3z
Wr7waY8LNqPEpJP4NW5VyWwsT0dXBZ7+R6PY/k36ymMMSJoPbvwQ0ag0dcyFrJe9
Lx4EqGPY3saRXzfc/6G284XgURylKBdehCZ6f/aNZC8s4Z+oMGg1cL6DIVTGal9N
dmtn0yti+tWsATGWemCBAavh72A2LYyIiwbobqP3qG/aunVdsk1WoWlMgl9WpiOs
89fBMrr9Dm+kyTGmMDMQkRnsNiww70nLRbS9Pu5YrgmOp4mxCTxgGoV0Bt9WtbxQ
2TzVzjW9kkYam4Y31LugqKrYHjRbdstHILohGoXieBR9DoJK5VZRqdFavxv8Afwt
wj0vhLRDXJyxcM9/CsYVI+hZtLHcd/1bWKdaOFj9TCLQM/wx6MPGpmD0VOgFTeMD
Lk+kqNDMovzGYcjE9bOAEsg3GHbgHbKr6Gh9FjiVKWwO8Oovogt7nQx0AwKugYM3
VBhn02qL6GvNYvtUObU1klE3lIvHtxyTnzHPNnzhTgmqnFPK9kM8932piLKzXA4I
cvm5GN3bGKAEAESk4S+2U8O/AvEeFlx1eSUBPWBCWw5PfPZpzAztrGRv64SW1Ugg
XMYS3xBxK1ZNmLgG/5spN32LOOA2vs/zpk8FId1FnfMnKxEyZHt4RzjDCC7SjzTg
kVdbFYqi2iU0XxxWG5sy02oG+D9uVmFR1yhRQzKBCH4EcOpEfYmDAph/w5B2n+4s
jFoHyfzOPEn5umzeQQ/w/qnMKG1LOPFQVx4ZUtYKiT3x6rsmYUbI/2OitUSEcNaP
QzuaGr0xvT7FqY1iih3JZXsQ5ti63iIsOO61edmiuuptJyPvLIkpmoptmrDCQ1MG
9pxht2rqUz0fvFn/1JOoSL+ZTDJkMmOcWptWmYIKuRGfXXnDfJPWiNkS0JorV8FG
h/6WkQUo2BZ599JofD1Z7b0cRcEkfwBoWhEixnoCMUSPxsrxqpOHhQPllXj4uggq
JgjFlWsj+B45T+4G5WrDYYNT9WJRAZKTTdJSWIB5FSpF6+V7rZi/81t/nLbJlt8/
FdwJ3WogFBpMZITmlQyfGHFvMV20DlpKpGB3HL63IZLQsrlAcQarlxs5H3Y1ZDnm
qYTk7VOVODMDhD6xoNoRy1anJbM1syyy3m1xbJDTWg/Cdg/ueRljMNlo6LLUwDgh
mfh961vu4YSh5HEfNeGnLYIGhMPzuPlUhdNlc9/gnqc8krnwJdBKTcLdnh4bIaCW
fChv8o+et1kM3ekkQ5mf/i6vGW2Vbmif2+QiKY9yVikMO+XRfNarUi+G1nNCTWp3
yKbQFg+bFYmfQQsFkUGBMcpvJlCRE6hYguJAZRsToJ+Ded1Zyvtbc7UvX2Nq4IWJ
6Ten9ox1cPEB+y0ZP5avW1YmaIP8vpnAE+Ksp0ZZTZlRizUj3aTlzYU7W6JSEpeI
d4UcfIj13DJTsR2mwL1ENFSMpxjsM4aW/6XRsnOrGdeZsS22ukig44o6gEFEl7Fg
7CJDsof/a/E76NhTBBkTYFVKkJf9cwpUVcybdzi8X8vZRKbDXxVIcgPGhYI/qavc
erj7kkPMbt7DOm0tuImPEzRi62ErAY7Nj+ZblV12b9bpzZCp0EXgNmNRtGAfXzuh
BU61CaokXwHelQxOipbtxTU0ebM7NrwPlmoupoVPAcojyc2ZfkYyRSmqtrv77kkQ
qDxsktc/Vu9xkBUHJbqQj7QXyw6JnVKZLzIHWjOsOhw+RLMrk3R/t6r2AH85HOx/
BjuG9EYDtH4ZoW0MC0m3VOugt+CQ9SK46xuLettz4BVNLkSpATXLMPs1PaHjerOI
C9g/ww2+Ula/0z2nlMFxW/06LYKZnZ+XmdI7SALLOFabOS4lXvo7HCBjQXKYdnxF
1UyuvPqclW+muLNdd/57b4yHpScbkE9idBc7BaaaeJrE6RpdW9L01d4y/fKzfZBu
KzMF7dsQmjNvqt5T7gLgZpxEcH4e93EEpZvL5VMvEEFqw2L5pFXAw1KNFJwKIrsV
a/XsVBCB0pBUcWsPtXzXYNQ/DxFsgthOaTRBgf5HBNvhBzzgc6T2HlpviU4Uds0I
Euf3epnbS9mFCaaqp76QC54SwCC+eVFTcImhdRmY6TCQvs9Hfpjwyxgfv5n3ZgQI
cCQj6DEt1EDA2HyfKf0oMfqEKMANEzPbqjMo3HBbzNZyGDWqExodCrT1C8y+BX7l
gFrTnM1eW9XKB/KAxCHwhw0eOOAzTZIL2ZIJwQRz9HV2vSACpBjzvpm1CoJN/4Cd
uZhCsYObg3s2+mPxrWOfOgATNtLHVNqqLQgActhwZk7MgkSMs2x1DEk6B219I6b1
6iCCJSLRas35MdqRM5qwCyOwrPD+PhOoAC0GEHqZn93fZ319s649I1vUpCWndyTL
6lWi346pNdUUdr42K564iorSR5Q0d0/u6nMtuUT3rS5vFzSXcFNhfieIntcfuM8/
5Zb2IFBpAnue1IbCQ+pb3/BhlpyFkrpmAH73zDzxDupqR8I/uEtaBKWx9g/3J+sq
f9gmwojCHiUU7iLasoGS8kQS/p+5VYyPZLfNJ3jYCs89kMszO+SkCWWFo5uIHy+T
5nfl/ot87W7ucArhYudWvu7EPZ/1AM0biLZX83c+svUbVodQ+clR2LMOLut1Kk5j
z3jV2du+9oY4NeRcTaxn0ID8BhrCdJZIRF8L27nYlp6HEWMmV+IJneopEaFJiFDS
aOteFz/UN0jXyUXg0no27Jwm33IcYZqwMVZa8b9kkyPXijYx2Lp2TO/PAJC41UN5
odofoa2L5TVN0AdqLGk94H1sWVfy9m41Y8o3QjD6xMis28HX04I5gZ5mKb1y+O5c
lPtAXNpgyItPGnIArHCF5W3quzhEy/jHYbZ3QkUObFdzNYVO+tojVhqP11lZ89MB
zdVaF3JWHVjTw8tNgR30qDa7lHjKVXWd4bu4MxbnbBQoikKNQwLSXgCxRKF6ehfF
IWgIiZDxyfD2iV7TQ6pj0FpFhFkiBApsPfPfQZXSCdadICElybknoBGqkLcjMx/E
7Gi+VQKIMgOL9XPwOZ1vEJGf/xZXCtci1wOm8TYwNi2Xxp9vfsQIpUHDASbcxA7i
GJUFnnnwa0siMqbzDJycCGMJYOoqTVsdrFG/Z+Vvo3Ds57ua+jPcg+dH7WnKZo73
5NgDH5a/K/JncON7NZRanh3X9S8ukW26TtL4eZpLKn10CYvJqoHahx0ShNsCcgzh
pAgNA3IKxj8WRSOOGTjefOiGNA6s9BnLgumNqyHUvYa6f7ESYi4G/B3R9o/XtTHO
2c2bomDgY5Zmkjt0Gn1dwJFoEEGbmoGPRxI+dwUYiWhT5N+FDg7knBzkGKCEjbdD
IZhN4EnCVNSouB8z4s1kNhVED1GI9qg/mQoRdiOC4GiP/SX2McQ0++E5iZ3lA/hZ
Cj45a7AL+/Fs2E6xNbFWwJq5LqhBm2dvbRjwTq5O8MnO7tlWeMOq941Zu1J4xbSV
wPlEyvOCI7XM8APjHO6zLUXjFNoP9E7GesP1O6CUxumOQp5t0bJmKkp9/HwdJ3F5
+6cyRldeI8xiQ8DsurPaTTA4QJQMzmsJJzqkWVzE8Q9oDNY90YaAjVEI9RcD8xoL
Jq3UGohmhMEMp8sZU5vjAMv83Oz5jPJgjpNeEEjgumdXYk0uRuD85X8RR/kdfgJi
CGNYe5lJIcV0b8FOuJ0RmNnqAWbiNXBtBABlp7x9dO6bHdDeab6g67jVEVXGVsVe
UZyJF67LnlQQV3ezkXhFsyLA9SZ+oBT3EYpzBn/0OcEHeDmgysb2OtXx+TT9iG+C
8+eUj/q3YiDX4bbKsVMX8RzTc5LsoxLSgPOjfK9xPccGojm9L4R83SxJdydkBimd
LM+5sQ2gc6N9kDaOYNQz2NG+DEeyiUrZeXxDPDybpexzdRz8+uIKonxnzML13/vS
1Hj+7FvqFHhlvC/9WisvM4csKfa0cPC5vvOTpEmsf82F+oY1ghY967BEUndmS0DG
nei6AEzZiN+pvDlHeJFSN0onukvuV43le3JXaLbYPO6E2sbkDfiYdi97HQlueyr3
fc7t0ScYb21aoWrzKkqpW9PGQTJSTdKjOZj03S7EsY/P2dwBuHfNQGBRmcxHUQdH
HX8ZwhXbxm8GsF17WSybmfc51VWRowyaINwkXvU2I5nkWrSEj3mdd4mREERXNWxK
1obs/5MOxRULYiRxncsHqJdbzYIq9VzaBqGMKOAdhdpNV0wnbP0IOkJ8w3UrUDHW
f0rhKwAcqTLR1ohfYa/XJzmQDjoofCVo3jQC45x20B2qaQdVfCHajnZsBmW51Yfk
ZtbHnlL2P2EspRiw1BxzCqFidPGZ9CFjwzItNUwXQuH+XrYocIs84DvoqxtfXlpe
hpmt10PwLpwPJ6GkgjBO8w/DcTQq/FZ9UuNydWItu2zyzNnZF4O4l0gk/3xpFbee
Uwd3mpXtku+zebJD9eQIHhsqOVRpVB6bhKMbI3uL1nbLwI9oW/j6obKNbZc9oKPR
awqol4OCNOyweSXOErin2CE9Wp9P5FanXvPjk/p7HgBIL8gsddtBw1Iz0NWs/Vq/
nDLKTdLuFDNdjA4mDP1oqqZYkcuGO6GgOSjP1QTZyuNmgLeaf8ufqocxSsIHcwT8
fQbM8UMHqPOq433h0GP6AmqDY2DFyXmDf22QoIMWssRJrt7y2A8sWsnKUx3GZfUU
f69ZgOoixxRNqikyYo6LxEIy+efpg8HI2nJNZgfMckrB101dep6dJ9kAeCzUN1kP
2y6cLBkTCu5GbwfCuEokI8DWlT4hQqN36gHLWZJlc3RcwOBqQ/nXNU3tXzO2qtn8
BIjO+YbLQFDUXiYwJ/FChA+y7G8TAjOXgkLfRi21y81HTOPqCdIBy886tpBOcVt7
q6svDioqRdIa2YMX0XsjJUkcogoCR2WfjhoffodYN675I8UwijCX6+qKfz3LLXET
3pdgsl9HG4bQSBHeSqoM4ED26tZqAYGI6aVupsDEPgjOOIZly35wjfI1uW6us8pm
UD685xVsctEaTQBFbJTtN8SgvGefeGBp+sFSrXaOVTNZU7TnTSpYU0NYTijNhode
/5n8IIyaixoZGkN+k5+4O6TpGd9o5uT2OYkPUJBIvXBe0WTMbP0U4W/117eUHDUN
A2WkgZV07vuHAgl8SCxGPo6lCHwLPFqEpRxhS/9P77SiqIDUdmMpZshAaH3GKcq2
LbjSwff1C8uf/pH2bn8tRaXYAXMrDXa4ipcGUZoYq0tEDT/2zRJsKYXDUOxOecUa
USY75BxZnKusOZM09E+TAGwKl47vy1YnspHgLuHcDvKSxMVVaxQ/aTsfT/yISz2Z
7FJ2AcpjDKfOTKPWmhY/EXQEMUHfNtevHqq80SpHb+ne/ta6AqWgz+QA7DrZIPIa
zd7wHewsJafVRlP/rMqvg1vh+Y07Q++pW3cK1hly/4NxunBmTgPiZlAHuE0M4+Yb
CXSxQpIDK2YBzf0bHFxTXNesQV9gRgXXHxXM/vCDbCTnVdZOhYWfeCHKzRGRbpu3
7eU0QMMUzPOyrVwVgdkvl45z+MmWtzIUS1wvwWHU1d73XddLMf4w16VLE/UNiyyb
4uIEILmPmeyUbxRu0X4JEWF30IptPSOFezrT1TSV2RO/MlfbtygUjPadeQiQ85m5
L1gkunhwCaUSOgiIq9JJa9oNGrs7DzHhQDZhH9cVlMU4e3XJbB00WNmgibzhB5Vj
xUiDRY0g00D8LGO5/bBGVNvdf0FFk2y1TfgnRn9qA04d327k6z2C1r0LgTFZV8/T
gkohWMe/O2XSeF+3fPzyE+bDL4bWoyCjvsfBdWswPJaulJo5GgtM19zc8F1+UY0R
ctXKbjbCO1/gK+q1xBfSZQsej4Xt6MEY3BU0fDiuWPevov5nP9/pyva1xZkPiCDA
oo3v4ZHGkYxrQiJk7N/e3yvOwAVx5vvmjy1KSHWBLPucz2F5KgJ39Qhqbeo81H0I
V7KM08jvWpkLiolWbnsYFe4/2a16nsqJtLXWrJFZggy0ghyvek/7j/6ULjpTW3Hu
Zvap1K9Z1R8iWK44D5bQIHjK3gDKqgfCd9dA1QyCbfsVuIU4xBsviNJYOZTkBDc9
rZcHLxXhRHuCwvOIDFIjk+Yo3d63Co0aURX9ApwOxL4z/qk14eAwGIy269krqS/8
WGuGkmaDLtgqoZ2uToSU1BsfOWGsTT1vot/62PbWC4qoPtcnFYLUD/oP9iVkH2gj
MUbdvQDwCFKn0tI8xB4Zy+DALiM/kVg35DIE5YMj15j9slP/RG4zCu7JVwTcInyA
u6BYccICAAPM4r+4nYQRkxfqA0whArMQbtBBK6p3JSZ06n6JK8Qc7GAREmtUvtU+
qutENKXnOKJHGefthSB0fN7VrdTKjsXp+GJhotFs3JlIJAYIid4OzWHwTvlegcCg
lEgpNuVyNpB+wfRPtQfngst/VdW7Fj11qgNCvYUeCpVkbTpDWDdAoAv0WGFgkGA/
UCc2Wi3bS+weZ57VoUv3ivbJq1l6TlTL1eODoj5IiOhYR3yDGXUh2RAY9c5mM4xV
OuhBEiwwKSgCFnql9zVgPuF1HPdi1ayD2ac1NrLN9QuWUVkv5vBz2QOtMSvbYTWd
iGdfTevgOKEnVGx20G4bX+NW7qMwqoPOkyJ2Bz8sqSpIW/mALn98cirm4GLoYj8C
V0ewtD5OFx01/Rz0OuKQXmGXZCR72WPaWbZigpPdzGcQNehO7FrBUDMfEt64l01d
3wwVkbwnD5GyyXPKvLNArZFvh58qPE2gsW4gboQDyl/7aqI8FzQbCtx1ipfJ0IQX
eNpuwhfBLW1qlNmkImLEIzFmXUIC/w69RhdkDljxFteg6yX0vHGCMwCUcxxOMM+D
Xr7hJeyM1IvMEee2okyacUbtES5enZRD2ODfMsBy9q4g2OjhLN+ZjnXwLO0sKyIB
d/C7tCrdgRDYirxDkOv3sz0FWQv97o3ZBJOvgpBh5Ud/5yBU6BVF8CMET9JKKCEu
9e0YrxEktoMcPIscyLAQtGHXvN6s7og9Kk1jS/Gvkc86HFDcnxvFt3KpVU20BFzh
+IU6k0XKeXF3IV2skhOqe9bW6VWhp9jZtWAjFnmMEnqg/Za+VjSW063FE/010TGF
thAxJED70uF/CdUSgvsxS0n1HJM+kIt3rKltNVAzfoIStz9/IVwZiy0sxDoJXHSo
eQYC039JDD8t+745Ye8n8BbN7mcOwzt78YNSQVVrzP/G7zbgHAjEHZbK4BguYGSk
P0z324h9Wpv5N9kjsKFe/Nx74pUR77ktho5aaFQni3za+RutuQYItR24BOMHuQHH
Ha5jwGO8ZGI76ATljvaJOdncXzf2zJE8wYPCNEB03sITBmofnNSD0abX8oOZHVVA
M2JdGfWgoiKhm8gHlmpSjFm5AkOTT/M3nQBDXHa0qvt8RaYvfT5WHT99KYMTPGZp
N9DoIRnD1S6wVxCSEjQqXDHrKosPGvleWLrSvL5ETAS1VWOM3I2U7+0E8r2yGpla
0rlFuCYN2feJpA4tAPo+4bKJJ/+FiRg46FVv/G1NbTibnM1CB3XP0HSFNu5wJCvl
kJiqhCY5sNQE/zU8D8kJZyLJ/T3FbTsDKieQbbFZ/FCPRTAy3gWlhgFq8rhm5UME
LAYIdO+Q7wjfLI0xmHvWT/uKmJAV4LVl98+XaOIGyIe8dj8g0BTQd7VtW5soheL/
oolWqLCYrlTvNLis+njN6f6XDK9y5gQ06B1bPZIjlddtKTl3B+Ao723PkFwOa8ct
0pDU3+44aB3gSSlec3sZObnV4q0f0REMPAEKS+N297Z5SjnD879ZiAR19SXjH0gS
qYPZbDoD89l3DrbfzcAdz75HT0UEWuABLNtlM6grO67xWyoOOv4e02l7zb77TTQy
Sja65kje9+BGwz9zzkdYPYQg7gsLYPOVPxqXg7oYi+4FdFworTJth4DHqkSw7F+K
gQ9ZBMMcNR2gpsFGLzSqVIASGfqWUIx6BG6dpfqNw90C14DadlfSHWxHPp4I1AM5
Zu290fXP4r/BI1FnzADR2UhMwfoXLJIxd4cHoUff5c1FwtxCoTDPi7lOvAtxGl9b
hEjhhYBb530HmYVuSf+qORiQRP32vt13IQ88/n+bHGdv+MlzRjbc79rgTaCw27Gs
ZryE+2a0QR+52qkG4cJCZBnY9fCwcukrnWLSjL75MfFYq9mvXZcbZmBEpe/LAwgE
OQNdkwP2uwl6OMetKU3d5IZrX6U8/wV/qstu5QYq/tOSKfuJZvzXkbjfI8JsbRFE
gjEWTmRPAJswPbTrBHWP8Yh1st3cVcnp291keMOhSAydOeaftyJbTAV/4GOwsArx
ZisWyQKV/0jaPOttZ3uRIJzNYOalqBX2p3T0U/kW2fpTfxuOIWXnvvnG6dy4G7gk
G3Pg6R4IpHJvIFOcr6oUVA5XU86fltVUY4uCqPA6G6iU5eo5hx894bzLaFg0BeIq
hc/DF/19x/OiSSFCHF6MpPLBJwoRJHP/EleEtCvrxRePm7IBbtgNB3HCVH5OX20y
AMwro4srI41nDjewbhJmtNKmftF37K6e+YM6LjjmKAPshpj0fQVkS32xGapgoJkO
KtZFgFIkDDDtkNOrVO0e8bJyD3bCmTUwIN8YvF6GmCvzh3M7G4vb/yi+Tn3omEv1
6/012ieCeiXcYU3gPy6iqKcnVsD0Q2SKwIUkMz5j1Ww8GFn0enAQlULEjti4aKbg
gQBTYyN2Q6vhR3fPg6DCKx5ckUGkrdBJtmZufH9vomhfxCF2yyUDQPTur/KA6lS+
TFqd+CWFJmj7cM3ZujjC+tm2KhBn2+mtSJiFd8xORImvg9RMemG+7SCPfWCz9coE
kRCatQB/0Zqky9zAcqw/oeiIaBc0n5Uwcau19D95gJN1oyn/FypD/pRqlIPaxsYa
R9hyQSCajgrnYiXWosKzI/ZchEW1ARel9eTsnbtpkHrJOwJdCxe+DdhJWC5f9fBt
ztmqE/1ggTXslaaR73vs06ekdYMO5oIS/03js5BFaBTilkNvuqQDAlzSKhQ2r757
H5pK85TZifLHQDOkIiADubkbkdcXWWMHv28iQBA7aZaCzc4MEOli+aH8r2iOr+0a
IqPHQEFspdh0ps347BIYEDnuBTYA0qE1lyJAie9mLxEEOCaPD2+Fb7YC6veayiJJ
5cbPC8hgT76XoHi+3Ap+12047yeb5SSTSiswZZ1N3cz+EmvtcjGeVUShjn6oI5jI
y5S0MFy2+u2bntc+tnQ5t0crqyIzXG7Ks0hSYGaUMqbabFnjGU4E13DZsjcpo3uA
5kRkw881pl5ldIjjKQPnCtg0a2fA2DRtC4qY9sbwhG5VNzZmht43TF+c/o5bo6O6
ggYmP6SF7T8Jmf0k3LtRWH0dY9tyKbMqiJ4HU8VGtVE17O6zRyDvEDRX7xJSOq4c
11RvDErxrkk3K7Mm3mrkyUEYmzdqFGhrbtDXbNw4AEkWEPDVjKqR1/3IxQmTjaZj
9N49/98hzeanU2GNRx4PAXnSEjzZMxrY/mm5Er14RHvkGwlyFGGqydCVbJx0h8ai
VA8HgsiEtbabgwksGbEavhfkPNzuYCasAU/HFzaM5Fa8HUIQpBduzF6F9myZyDDH
zp2TkJ1ekp7eEhO7dYNZAZUWfs2ywcECQvjJPDSHqT41nSZisoRHX2+PKmClxLvJ
7vRU86mgv5YsMhaJljpkpl20pHMbJKuJGVv3ZGqqhUJosNMuNEHtfLWh333uJ8vN
QXmdPcHKkevZXPPHWmH4EVFwLMY0Aua9GOI21USQ7q0wqrYy3ckaSFDuK9dmCI9e
hDtS7gQxk0bdBAMXiktoyS+JbTAC8yMeLca/NkeQgLvlrrkVVG4Ii/GAbDGv/8jA
v6vB3YHquVCFpf5ufPKe1D46UsnE/A0bVcW28wI22NbwD5gjBnwFSUaiieIu+hy2
3gnEcuMkQRhHfAphtzS51iJrx6YU7NoWxoV5UKd6hzaR4T0hn/421dMk8CsCLKaA
epJEfKRRmoD1E1dUZ2vJrXCXKhtokLpYMDKmPZGmvw8bO6tkVJJgZgpWzrGBqBTK
JewZvMUDfm6uB8Or22yrrb/3JyG0xSf5zLgEZoN8PX4/UtdM9mqgNinN/sBzZddE
sYXJkwZywSyGpy7bCJTDpfSXLfxC2lJdXMHF5OD8I31tEteDv16KGvq6U/30SBpS
U6yOoNXkt++WuZEyJ/Fm40T5e9mOgMEPt8A2KzicmY7P18FeBkEUyxGHBgB/rjRK
vBi42h1jIu+kuk3BCfWSKXFQwnXAl4F8clPiCtJSakPv15DHaDV3Jvf7dC9poz7s
+ASHca5h4+dKKCWSaKSAZLkgDUzqgNsk/B982Y+s6Z+5WtEtISA+UZ5zoStMKfzn
uOoHS7/tfLyELlAoJHPqe+vcwtgeMu2ZM3L8eZLWqYRdUF21zmlWQMGPPEDGUiB9
0qLu3GRP7e1b5oeNtR/ycekx7JPIMnIR0YNnMijvcIXWPMju6zg+kY3DK5Amc4od
8osPi96Jw6lrASbe5pfvNVX1tbdQ49Cqzc0Jbub1L9QZVaGfbgfSJdxWOIcqez/M
VhBS4q5Ys2gMkSTpvv5XlXa58N1VEWZY64Oa1IZAt3in0xiktaT+9cb6QmhlZMjq
/geaDd/HryG2cP20qjF67Wc8/sFMDoKSjcI6eMBTKrJEtN8lcmSmsgJ038eRSAxE
N3N8wSmEVVWjCn/PGfm6xLAtvNkbN6M/biGEj4zi7AtVC4YYrN6q2ZuCWY4v+dIj
SA4a1cr6yiH3qjL8ZPz6Z/rI3l7XFnUpZTaieXg1Dl+rGMBzPI1YC5bGvSVx67GC
+auccCwxpY0W8mUUwOuf7RApGnFQvWwCGKmpDZhMWPDdCyV9iCkAaNZ+PJudmGyV
iT8KlmF6D6aY5aj3sR47IuPEHENBoGjtbEh03LOxOuRortiJOlDTsjtpibI0xrbZ
NfPjH3pDo+sjC3T7KwfmM8mI5Vw5+6YIYrzCRR1dpGsDB2VpH8kP+ovifMyYVfYm
fQToE0KSULDAiK98d3j3qAgjlof3u2zdJTMv4VKB1dLxCnxx2xHvUxOJUg0WO58y
b1ZOZF+ZCCrwvyNyzMy6hm4XPSF2yxRP7XfsKo1MaCVIRpLb+O4Qov476UhYMFoZ
2WWkS1JNqHFIS1bP6OtkcNG6LWYyAtXgtXoRu5/0DkYnkUodUX3J5xnxGFy7x6pb
NgRn5L6wj22VInG/Bp5zoH9n46hOYFlo/01a/6wLEN6JIEZwIZUFsqgcTHPuOZnL
NBJ5loNR+FAOnQV3dcXwMcdk3+5oILRBzhvzjzb6wzjK+L+re/s8RL2O2s3m7+YZ
NHrrf/EhMFNILb6BjH91CNsCa5sRiGCm2ybi9ElACODkSXpqHlTI277WdeNGfCKZ
8X1aQJE2zUji4ow2GgmplQuIuLW7P/z0W/Pl9u3R4EUVDYpRYNMat10Kl6exqlUT
xL9bXNLKa1zmeuqVXJvLFSxWfQ5B73Np/sSFni6XIl4dIeQhwQJEEvxqQoqARF+2
Eevd19O+lD7B+snqtFpQUZSVi4gKFBDS1/EEz+JrNWbbPG6EdeiPt1GchYlttXf5
ziIsZhaJUr5IqWsQq8+76gQTGh5wFNaT4wtmfQkhZ5Q7oM89XO+aZ9SRfMJiaAD/
tpqKKOzHQnEIrUfEeD2yPdqEL+7y/6pHUsa/dpTncwYYUuvanWjPCL9htMpXl77L
9Ae3RQkNMeSRNNw0WFapx1+2YKs3CWew0ITxr1Av+xM4tyU14C7R25Yfdev3NeGN
eu1rX/OIoCkYQQXyE2MTNKUM+3LtPKfd6zfO7RN236orTPKHwRiZiS63gDaLwboG
0aSySQwTGudqNRtrfDKu1KffTY/e3XnPgr8vBnY1PlZqhRjUlbY3In8saccBv79Y
YwksyRXXSDfEZn0EpGkvsvzlRyoGBh5lUhhyivqBUbF2WPgz7IcRRSzlQx+Y9+iG
/Pbc6uODUszwyUjtTXivyAApWD43vDvxWq5fQYdGeojWGE0fwaiNFhcq8BEQeZKh
Xtp0akc4X9TeSA0xSFiMLqD19X/3ZFt32EVAkoV4u8cZmPOkP6tCui/vsD0ySgjl
jdfTcUihpqXx7ADEr31fyAxMJDi0umAGK8fZOydCDSkOogK/RPicgJM1W+WUGKIW
pDr4WwvzNluOpvx4bBQwXavF38FYtJiJjPry9YRcPeq/PQRyyWI15raVANoETYnN
29pSu001qnWrwcpW/fx4Fkj5y4Txnuo3HTuiK3d5/iweRtokSTqf7DI0l0KEYxSn
M2aE+TJ73oGYuuPZ6BIFZ459xpLsiGE7OWZ3kX+XTXvlFAa/vpdZjWGEGrdx1txj
SyVJpgwDDYVRWoZ6v7+IuYQju+muLkY0dJmxT71jLxSXEhuF1mwe7IGb4mkQBW6f
blT+Nlr6UwkBfa/l9hZxpaRspRgcvfDv4Od+C4AkWoFtEv+e1gdpRXLMoqhV8qvS
aofVyF82aDKlCR2PdJfabeyWMSDDVLo7pYxtaPirCGN13gevoLPnkA9M6037O+ev
Grku1RcAxGAlf9uj5K7yJkwF2Jc26OX3P23aazLIK5hCz3ixb3HHqbGxZeqMPuDD
vkCDX0xvRR70bk2GQHYgpboXjY4Xhoedum9SmKDdG8LIU4ESboXnlJAvX/wX0f3d
02DbVR7deqbxMViZUn4Uzn/E9pYvkhN+OxJtGVJnr0/IUAF1aaOKbfgilkBTeLHM
pkmrqDfOlhndLQAO/cXkOgDDDkHkARACwStpplXSzro3ZjeJMJ+7s5Uo8paEOhmt
chwIW9/vkf8jOTHpOc3GPRspz5wPLHA917Oo7g8LGqH1chMSJDlN5vxUYGEQAPBK
Nu0mG3C45YL1Sg0Tc5TRcAFUU2v/0qmS/ZYKbKH39h53ftBHpqO44gmmFUJXf6FL
Aj02fkjpSBx/jIT7pmWTNFDQ5L391SvBohYiXOYreejD8N58DsdrWg7f9DQFqAu0
lDewdWikQ3VNofQz3hS0tk05TzezABilIMiqSRM/4MWODbcGPH6xbvXkTX0CblX0
cszAYJTbe0p6iuO5HTjDoU8PsNCn/VsQeBvPm8vOt7e6KajyROKjqTu/1DaBArZ6
gLh/d9V/I6pBxCOHAG5xdrUPQDx81DRvOAX4QRJ6z2UB0Kf0yxl7mVlz3MI2fEdk
dXhxpvQzAbcwDN5jO4OGHi0Bvef3W130Rn98ZaosKTze1rNnbpCrqzAP3etXej17
1xHHEVz8LDMxJP6o7Wk4pSzdRnbdeZMUjdRJgGS7Ttoc9oejydWBvdislPLKXP3j
LNX3qwFESBMp2fIeM/7cjWQfo09XoU2EbfUe1l4PMr3AFBnYdXqoXA3Vmu4XTPgR
9RwtmBfyDv95RhES1GyVN0a/l6s/ORc6Gol2bI0msruJS9xHb50xAX8sgd/NzFXm
eKvTxR8bPz8D3WD00ISJnbVCK1Qh/2a7Zqd7QaoiFrF/9fhBuY7NwIBSBmXkXeby
glp3coONpE2ZgFDv8eE3on4CPrxJr1+OER4y7o8HF3gihxP3EH3Ug8CHXhFD3mZ5
dIb+EDUA9FIMccNsNHRZpwPgVDoFnijMFwGNdqa3LPWd8Pp6k+pURKbFvy8666Os
6U5//2XFChf7+57y0ngbey0nLU94bXgeLd3PDPEk5793r21J7NaCcw4vKAHWdEfB
SI0y8iIBNRgJiD3L0T6GTXkc+IALZghNvt5Ns1ehVYuK/aZLqrl89w1knqVhy0+l
4fNIAc3+RqKLUPf6zucJSb3io70WTbkWcO5dkfvt5m0n0Pie2JgwxBh22r5vBc6j
9uBaoFLZw3rN9WqM/eoCBYTiXB1EHmGWoZLsd7LmGtXyTRuSglnbZhHjTN4RLDkW
ibf5MAKbyrcdMUOZHM5M+DtfAfwMQOsHKwgCMULdE5X8a8k+t4qxRYY4jwzi+ciC
LwGzYs5CQ3JSN+am7Oy6mfctspETdccDxVG8DvrP5sXfgqTzj/XYuYqJjWpN1les
F+e1Ttz2+nI+o3qe2mNSjwo9JOFeNvZ5HBZ797Hph8v//myqK4X4Tssq1DKywubW
c4SF+Ol13yJ9LV09Dg/ou6udOYaL4dSGDeCytKFbnbIeqTyXAmcSUj7pjLCtauyn
47jGqSG1OlKJOYHQKdrAqHqMe1C+tNyphVse9bV4aNKQae3fDjFbf9YNvV3eDFcV
+N2M5N9dHiynf3QL+KN3+Jlwb8cX19WP8t5MwC9B7WNwFBr1nAz7yr8sbn3VNCOV
37A1yHsEsjNm0WzimjQg/o05nAdyjmEpNRnzNTQPN1A65a2sSUOLqJfEY9jwr530
9pkFSVrwhOpJf0vbXXR7VUVtUStGl1j1DFMw5TTo546EqJ3R7lkixUlF9npVvcpu
EFFEQekBWBPagTmr5cG7txr/5+h/IYEJQJLxINZVjWHUL7nfRkng6pbsNvAt5HbI
9vA0uuWzBhW8IERu0WeWMB0hpNGe1DpGriK9ArYpWUBNlfroPNY7fGdiEjlYaHuK
NA9r/V8pyfaLmju7bQTiek4PRpAvEiiPUu+4anyNQ0MBRAmaOfCrr+iQewBODmvN
fm3/bznZ4hdgjEUTEu6Vw22Xnug8vTHC6PL2u3U1tfww1+XMVADa4n84wV6v2dDX
wX4R0Uh8SEfujgDsbeD+r5kOkGJgTCosYRYXHvnaUEfmT6J+Y0dks4xmuA6/njk6
rX5aqXODZ3fuKbAGjNXoP+h6RnlW2OQrmKgNSogS07HVgaZ/fMnKzWI63orlkB3h
4TnuPYaQT40NFba5jGS51DWJxQi5VU60LurJkRSuCTCSGzTzFGGhZa4IckAq62V+
SeWLZpGaGKYzbSM0LDqqLtTIpHbiemy4Qz1W7WWR/6mUK9Qs3OawZCrAQYWs8H3r
UsiAzTUnFGH06ph4d5nmzHM0L8IGS3LJShGZdLS1SCsbxxuJOVVU6mvPkc2L/nge
VwTxVdsy+86J4XM2FvyNcjouEQWXzerTQt+Zrw+6xmEcu2j9f8ZF0LjKtE8x91Yh
1dXPZ9zE3S4yRX7LHGMQvd6hGa1XxKrwQBJjldeb9BPoqlRfXwp1MEAt0ZBYeCjs
urMw3boUTlJwtpqbE4//AhXvmQPSTqkb4nOrUz4i4xECZM9JAV9eogmoh2H5OT7k
jRMfEujv3U5HPqgJv40PWNwsOtMjPT2eEFNcPupXT6Fk1DRV3HNqb9WhIZSTcvoK
w4upKiUJm8BrR2Zs2VTsKyqer2iApHhr3lHddYGK4YvagG09BSowWFVDcUUCbCPF
cRXtwO6gwZyTYsHWEkn5oF6MEi2xTBHSk4OuSpAicsq+r0CRkThZP9dxEmSXxazQ
aCgOjPNrEg1pyWOn86zUNuODTSwQaJ48LkH3kwPjsl6xzZjNBVNFxzxXEXEoJIEm
wLQHnMy1TTvYJE96WdOlW87ysQkUCnd0g9mkYHiOd6xl+ri5W8G65SIpN4KmvgMl
Ffq36qMdmpoh0A60zb/JzKyp3vsPaY1WqltEMwF+NOqtAt4pkX6bGBZSY8udGQIr
JLRvQUMxwd5c8IxmgnrVQvCXAe/qnuz22SzDq1yv9F5qP46hivaK9IbOzwgWJZI8
Pl+Dbx+BL2EU6a+EE8r7NnSHPj394MgmQycOM9yPd0NQhOex1x3CLUemilhfRMX1
GIsXCHTiSV1UHq1i0RyRts/OQQjqYOCiH8JbM9zlv2w0u6Gb+4Z2jPpR3MUyhp73
9HlLuO2vwAnKxATDmFL50cl9A5X217XzlnETmnkJ+KiRzr2T45EOJrEvvvDyf0u7
5VDoi5Tn2tY/2qtYRVFAnVkIsHM3pehyKLtk+OLy7K25FaxexMM8VhABsemjtp8S
4k02wpfuNGK+gfUGvvtsu4wgQL3e6KDG5c5cqK6jmp3fMVqvbfc1ZlYucN0oejPl
UKicLXLPB/ZBPYmTt8WX+lBkE1LKUgWADqmuPER7/BNr6dcnnwnLMD50S+PMDJKD
2i/plgMjKWuJRAxCmEDAPINgv/dXKaDOWIhlhfR77JCYqttC0adtjKZ+Mq08C+ZQ
PRL6hD6OjpPUKXD7bc4O4pY5oVFI6C/RUGVJUwFDmxH6u7dr5ILrSeIF5aGTbkMu
+Pe+dikTaR4ZjpLqKSnJO/ef5GfU+PxsQV3Yqq38Xuray8i+ybaxDz2NpQySzehF
DB+YwY45clVItFSZOLBTNHij7sKiP1i2IPHB5h7ehcmPS5RFPn2zj+s4Ne0HWWO+
TLLje36IvgBh1js3RFKErzdOCXzZZ04gElqCthhwHYxskPQsRTl7i0xFRVx5hd1k
q9wCQICvhzd7QHe4WwNJsNP2YsceALijRdSEG0p/ULY0AqCVusPW+qcR1HCaz0HA
BIm2YKXEJXivB7jy2dI/eYFDUXI5hvO8o4IETYZizuEHM2X9Sz7VRk4RJa9cz9LH
fDaUErZ648EGPKpJeoCogLx3Qx+pNaWV+wFSsOd0/bo+ybi5bebwPaoT7G0hKjm1
OlAHOhUoOrR1SeA2MHFgbsZsEfdVdjbWvfhML1qRgvqDmuwwQT9Rs9WNev3EEueX
yW7uKsdQFLH0GaaywX3W5eJQQRWcWCPqSXMZVc1gVbuMGBUpjOYvFfY6JOHy/mZO
Bq3UsIVy12yS4Miqi8qEwHZ7MLkp2j7UBQUx0MLBRyf4zrYCxm3liMkXY6dL/nEj
aokjHWBcURclCct82ECBMb+BENGq7KqcRZ/zZfccbzRShM0UhtKNWX97YhUxmFTm
wbVUCD+SBuBiPpbrMkfobI515Xz6C0LPex5MFwKMRRkXi1ftGs5tpaZQvtGTAyp2
GrMMsCcSCHSbDWr93s9rrEmy8qPhkRbmPYVZM2DaHyIal9W0z9kLC2/qLCCGVRJ7
jZ4XIT6dE3Ai40xt/xdfB21TCJdPzHO+xLZGo5ilCYIIGOwHgPRcpC34ND4Yc22P
5ND1zF1ADZTfzksfANbkqHuVSAGXYMAx2A5XN5gOWi54ZEG6RWOipRnKe9q0PMiJ
8fD1CbbPgZKUaZn1om3Y6TrBcbSScxZETQnLtapSvl8kxmkKPgkhlLG5JUlixFhs
aMPJyHztY9aZRC2M9+6DVk59iD/DpYc3rqRno+tacra6/fvTWSxUY4n535p3N2v2
wFyUugn2g7+L7CgBZ6ZX2AsJGzkHh0TqvIl3KryECXQB0F/kB6ge98KrH8/EHhWF
oqCtG3n2yxz+WA0rj5dJY1i6lb2ADEAOHxqTarSKG1lfBKYnN50SU3mByowraQUk
fZCWGgM9Mysz9VR9KquIh7ND7bY6ct2RJ1h8CDywR9OZgcYkXDfxoC/4nZsv5yox
0OjG9ewmiCHQuRnNyeodbAQJrVzfovgf9bf+bPuyUOSN0wdtwOLRkbNTxrW+lKqM
Vgevz3eT3uulA/82B+waAFWya2OYPWIUWmwlnviv434nen6V5Xsf4LmzMrmaqw4d
ukqF4q47BwAEAwhy5RfbRt6+c3fgmysOqZRUP7KC0/KtauomALknK3v942novDHb
G3YdkhVpOukHGwFTbfnsyk05zR5RtaT9lPG3B2kQ1AF872wskkdZLT0G+JIPzxvI
x8zPCkHyD9R1ZacwO4nhEqmbz1w1reLjBWr8e8YGQgh90Ym+qQdTauyP3pLf5fbw
ekzOZpRPQFO8c/blL8wIfETzL/T/KESbrPlQRsPVLYZyRQ+W1jvBgn7umryjr77j
CYAzJuoe3TCo6QNpJwftC3mcIVSHgFdzCwF3p2YENZSNhZLOFCPadssHGpEi+43h
Zk9H2tE1olhfQ43BxsBSGAjAImZWeDgDifpLpjhDfVkh5tJmq64V49BmpIlVYGwd
pMWfBhNkYqulYs8boD3PKQUQBN0mbSFo6Me9xfkAAZG0dBiG4ywq2L6eDYNo+YyW
Zix3d8PLWCIv0aZY5SK1/gL5meXkVXerw+blxziUaKuBA+HxCpvgdFM2p1B7go0s
7ucGNFbvvpNgmY0J2HmCunk4kwdsJ7jLqSkUxoEhpyuh4OCRZDOHxGyHbYEWIskA
1/cT4m6tYREFc0YUK9hEoINIW74hD7tyO/LOZ2ngmEAjJqW8tmlDfQiCf42vwJtb
zDQAr51P+aVVewajFNM7/nnpXnOnsx10fVAo/lBscDox4I9MOrYrKxpOaM5wYqnS
QyfYtiApeXuVjOOgdRKYgKMhZ/Bk46zqx/1W4dMHYvwqWzBAr2H4R2wz52e5dKqf
Uka30YZzo16RulM9D4Z+1Fon/SSXeRaff4lu9rkt2x6eXXmLPxiAAJv5ylkIlyLg
y+NhQIZ1yUSL1raV2KtBmwXt8j5gpTasL7uzN7fLAKvzNzbfQM562hxfxW67RkTi
1qEhH9WwdV3G4twpatNLIVt8dDsqoWPxZeDhWaOHlH75Pj8c7bty8AZI/po3XWVn
mZQ3CPUgAv6frhJYjhsTQPryOo7LZML8geP207QRlBHqCfkRugT9LO7bgLK3xS7d
+/0Nsy9+9o9YoQZ7lo5A+jSXNlx/KEVHSHywrFmwSosPTRUPx4LJD0rrvVPwG3jE
pMqW4mAhSbxxaV4Mqo/0NMtOCTZusKpenOgQofJ3EJxf9aSdqWJaMZYUSgyZCZ7F
sfq5vKv8GsBEwUt6p4jWukuWtJSKM3twvVqisHodj9bo6TzbR1yKBSScs11+9Jvd
gdJFA4VLtnKVspFExj9TXlxBOd9KMM7jvlc4VSxvi6PTGFBtENrsIVaegWaGX3RW
KBiFLNZW9OQDjkEA/JLinfIr0qaTGH49G0xf0Zwwhs6JbUB/WmlMe84Hm8M2kAPD
l4jOO6FcAlTYkWtQy2qLC1qXAmlhCp86UB7dA4rGfTxrQ176QzQabCDaA983f1e6
27QltP2GjVkveJOsov1K9ophIxiTx3MU8b/kdN8eahminMSNAUEcpDZGvAV65qMQ
+475vaeR/JUToGCm0g9+dvhI8rzSxg2hNzBvEbtFnBgwhKFGKxCndyMc+khfYAKu
Zaj1vTUWqrSdFupMYciwxnkG3oGvclR0omxJoUJSp7V+6/dQTFcZpa3QwB3SJIe2
koZf5jDNfxwDqYWhTBFjm6QJ0Z3ENHedykaiW8jpxzNku6fTRfvsRSqaPDTgHBr0
7PmDFjcL1SZKVEUXsy+OlOKSCXHq7Owyar0rqctDzPdAEY2LiUcuPONn3N4M6rID
hZ7aq29bomozdfZnqcdBp1Jcpsa70GW0rIf1tRmmsLv/qP28w9ufiyZiwHk/o5FQ
mgyb4br/BLmK961GMjA1/jk8fcElMp2iLbvrBAqBjlLcOHIzSWW/2SVuJ3hI+2Vu
nzl/lm9N2lsJL/G++11zCpGgfhKFxFIWQKFO6TsDAayxLD3orc4oNbwO/djLrcTs
5pSeBSu8m3dxSP9HMlpG3rffZuMrkVaETiBx4rnAYSIR0fx5TKPvNK28iEJQHJ5z
KTq9pPbMAMjKxKcbmLzh3MAVJlfgqqWN6bU0gBt7sHVAsa43NEZZhgmJChUGRVfW
cnSe9pg/96WR3udah1Q0oTROgNPMsumU+J4ZOZ4ivt7Nqi+1vfrxcEwIvjUYtztt
XMFOlVg2n0NJGk6m2RG4mmMSZighJTcwbAwH3tSSPTsBZNAir7rymxf4cIu8/sFA
qbjBD/UNA8KT2pkOGLaAVxnKkqJMREd76XXzQI7qYHKV5HfkWv4Jo+D5QG/o6uAJ
7Yt9UwXSgWTGbvNMWMAwyy0P5YmPNGssSAS/4JPMd37rIWXjdUBj+AJDXdojypWx
AlbJIQRgyRRc1WpSIfa706ufUBhhSWe1hTXz7iMYrCSLh2GD8JLsXVCmzkp7Ljxz
zT8ep6We+TP0uLWPHfwbYSl+88ih3cNp8wMM2lGSEGcXwZR5D01oaYnbspaKACJN
ho7M4Fr3xyqrek3o9Mmgiy3abHyPswTXLH28q2zHrgNRsxMNqzpD2kx3fVy4hlQX
4Ff+SCkoVg5O8EAdXlJJ3+sMXbL1qT2TLinv/oeHZoY9Go0JVHXLT9LrFLAHCoF8
VdQwse/KHsglYGepywmELK5q/wIGZnuvEwQ0Oyba3I4XtFFhDTH0rWed8cY3oxqp
hr07XW1J5touxXS+lOHeFBJC83/Wl/Ny8lkvvHevsfWMlyydDEHRpnV1suO+IEr6
j1To2Ig6LlBtA7cx6Y+VtdG5vaWy7axtqLHSbrPmKE0wsWNPUlVvsa41DVypbYUK
7E/c9SfOq79DUtbiFb733BQCkHpcJlKN8QuNNwL6nnziRIrSBknYoT+IFEeo4kNN
lzlK5HZd94D73Cy4uqa84XOqz3bm7goiu4p0z/srBd1clWitFPdJqsWL+JkCuKyR
/lW7BPTUikWjdHuCfpfM+5n/76aoxX2FXpkWtvJv/TD5MxkSMaseo5FJIDAONG57
PjV3DNQ8kdAz7JETtqLhuk8UwoCBQwGvSSJ4GUdCjMOlUaDiib+K3fHrAJUvtbc7
VMdAzLuHRAvU/nHOHWW7wLrtShH6c8KuTGj8oPRe7+H4eAvHj5kFWTM+rwg4+BAM
S0ihiHS9JtGjzG1cmn3ljQIlbm/r3EKRHCO/w6adQGg8VmYj9KzU5ehmsBbCU/ZI
tNKkBrAXAPWmdi4DxXcmRRfMhRQV8SxrcABBbzmvWIiHmZtt3sk8tpOG+Ud5gqEr
e/TIjuWICedcRIlhrLhh+mXAyXw/Ldiw7m5uYlzi5W4WYxKAfV9dSTeX4LOyC4+q
/cZNlOVLBYRw7cCO9nPSxhWxaYBOMNHnrUTczjbo54N2E6s5MvQJNp0nCVcUe7NK
UaORCkzKFc7VGB1/57HW4lxYNUxY/yLidlyB41F9rIGatC0Y5pIL/Fi9QNJC0s6f
fZJg22DFtOvPVsxbD+0T5LVXRbGEjvdngGbba6r7z5tBvE6JW55OJaSxqNSGfXXC
GpXDfth2+7UTLaTfbaGOL1LHRbgzUydyTdL8l6TgzY0jHWlO8kziZqh5xIaI52Vi
oh05qLIBQBp/SHI9huVk4M+K50sEWUbT6H+LvkJg13/gIEoaXELV7NgnIWCce8LO
dkhMQR3XgA2uoQI1xwYdoCiT+q4834NQrCrW6mRkpB/dWcx22ehArP1l691FcA/p
zKsEWq2DFuoyEuUtqEGT/rrzY9vzn2Q4ue61K4CR/pjkfw5AqvxtsT11igyK2meD
Q+cAZoXkSg7K5qFAkP2eP3mwNJGOT22mKkRzEDkdHa2CJ5B/oSQaXpWbpNz0H8bu
bTXH48hd5r/zmJqSMWjdcQ2A2QQV/zBbB+fpwwHK3FHQH8mr6rrJWiKM+jXZIWS7
A6x0neprGzRLIrG29yJbHM7YvNWPJAvHKOjdAz8DSgxao0ybNGk0ilBcaEaiEEeO
xrA/nz5/zBlYW6XVCWj+M9hNlALlAq8RE0hJY0R2QcRkUwncIipm80c3unuuSIIJ
Ziv8Hv+ObQoBnAdGQLatijs9/LQuEF8XUVRyeDwNVdOLAoP8utTsxIoaQNgYR2uo
fvl8jqSqt7z1OlR5t1Olxq6M+dLbI+p/MxzI48Ey4QPuFN5S9By6nhgNBnHwK1ZP
zFlzFYn6hAIFMsZJJOc9d4ZHR6pCkahwN6K/gu6WhaWik/K6qVkhNU4aXH/rAYZV
ZR3PGEgqQRpAAurvWyfSEP3+zq2zN2yDOYGgeT+qQwPAoaAn+g6BY/GAuyTsQNSN
v/ZDm4cefN4TdpV6IusCTLLCGEOwfmHGSNDbbv3ZVOFr17YDyFiUdi9bs7fylPQQ
ZhpolVDkpfEUzUSFejkTKHhtAf/wHkvTzCSQnUHDD34/v1N6AcSM5Z1bGxfotrD3
mAj4x/SLcPbLRefE7NnffkvyqOHSMM5l+QxOYFHoHtoQAqYhmvJlGtXAJrJvGpg3
hf2IGDcarkg2TFd8ClxHI6pXH7CphdnLlcMWzdyiOFplUebKQt+Na1g/szTQ0vtQ
3NS7xAXXUh7cyEKXxEJmKP+gjPBhdYP7ujdrJulSHB+Y8kaZ6TLD2NZfEVfI5jlm
qiGfDllv6XNwJujXeKvTG7wwpWf47vwS4lDaERb19e5pF5S2SXTI0c+274YKR3Ip
D4cR7fJV5Ko61wgofn0YO3iSGQG62rBuU+9GRKBRP85HG2vuBA+Ih+E+/Ibfp2qz
3Fs3NzRBLPV+cjMoQjdr6vs35yKzbVqrPsJo+SU8aZhkS3tkVBEUOW85ePllxhAv
10n/+7pJssMCYQLX7VjXoNk+656CBIaly5CVYvARG6DBnp9UQylZf9b8ej7z9ID3
R9caK26u0+TQoGSgdXVJtQ0egKMmXEfkLL9yZqxbv9lE4lebV7EgxpYXFmexqDLj
gKvUJIhyaOg/VqHN3RYY0nzGj4mqF5wUoErZbL3pXGkK7K/FIMDNUuby548gaO1I
WOTSA530WUBwPfku2MUua4mHCFugdlHP/l0hLUw49vZDm+lIkcFunBqj5WUHt+z8
wuZX/i5HoDjbYexTFZ5h6d5OJigw0/DrqhgGCIUxA82mHuVQ07M59AG7IU1fwBwu
qZiHrxyeU4l227HPXWt8Fzm1uoVsFnWeyGnk5k+tQ/LXuCkZosYfqAouZ/sP3Z0/
255VWnayPKK0Y2g3yLjg59tpFxRWWSrZWv4ug9aniDebu92lKxbuiXLvAAFJq5EA
Qx9N+sFaDYUSDa5c15aG7Fr3MyBP/r8fm2o07qTBaN2H8ML5BdNmlS3f/Cz+OYrN
8qiEx/kbek5vTGHNv5SyaR0wyldzTUpS6cQxTKgbz5fYVdgweqjEWMU1/AS9eYoI
/g/y4HEJKMeHt8fGRex05mB61Cz7DmJpaRmAQhIUj7PhCnRBTK+SCk6qCR1Fp4Ha
rSE9NbbEx9ygXWjLHmQfCECWkZvig1A7QlMaurd8y5nq5nj+RY9aaSL2QU7I7ClF
caI3KBR1hcD2i84kJow0lxKyq9bal6b5RYupX/1tSyapwMDQwMEQOpHbKwx+WPWj
DkDpmKq6oHo2Gyf2Aw+RVRMKL0LhS5hTMxw4rOmFU4cLxvAtgWhCyGipQXRA1yrB
h4EagQlbfBfVC49kX3/TFshemGAkd6a8xart5ruPk7K5QcPr+/kdGef0nw1Sl5sO
nTxrQIrI+fIxNI0Il9pH6TZpUDMHbVbN9dH58hK1wu67x2XuUuopC8pItvHGAdTz
DG2L2ULEeJ+33Xv/rFMhmdi2Mx17uQ6c2JGleFKWT/8DrGEO5yGZtlaUd++a30BX
7g8o+8agt8++1qOodMnRRIpEDyINKIzvPXXtgfn9VcDJZSJ0bXLeV2ifJmeiC4N3
ga055hcGW+eClMy64WFlmoDK6OzBSc6Hcv11mE1HLGSHIU1HQMe5oycllAqXYdMe
On5QuhZbFgY+OYBoGRm2v2vg3zpZfdP18PmagXN/ZXD33xRvnnbG6+c6i3LK/nVf
6txd1oKw+yTz734yWrSfFVTFDxc8Ft5ylcaLKFWAMQ+zdaFwJ5/+DoNgVbg5YdD6
X8Q79o43KtCoUOOBq1UwOb+I4wOSizIk2n64X6bbtMgCUWn1jOk5otVlafJyx0W7
ObUon1diCiSYecfBr0Dpxqi7aRcLOXPCJGUa5JUZ/4d4Tnd0vsGrxiChV3tEEgUU
SkIyestsrAHpQVuEL1uvULbJmogsnfsmAQ2/NiwRXh3sEwmBbduVxWjGW9+Y7fQr
TG6tNi0vtq9AiIyfxvgRpHiomQHXIn+AQum2JRSyLvo/Zg8J8J7K6eYVIkIyNzYW
6woA8zohmTTwRCUILh6O94Af9SadqtGiOVQXseATnWKJw7VQnVseV1uPP9WtrjWR
GwtTcOxECDfujX0TRtY3h7bi9AkFw/D6aI9NiT5y8Jh0aq3rlj3u1aein17dY4mj
tCMod0zFtZeArIpmN0c3/wX0H2Yj3Z16j2v88kmM8SEgHaLyQfL9eXBEyRl1i5iU
NtaOO1wRPvzMb1YI+nJ5pNMignWF4IWv16MjvT2NJTRCMwnWXY57LFXkf+URnX74
7ErAjLEdyAVobKRxe8aJErsrK9xAj+RVrfVZ5cydFUl4aG8H6waVoljpO0mvq5Qe
HxTstU5qsYCSpqZvISMdbjf/Pjp48GJzvtHgBTMe6seGVkbZv1uwYqKGwB15aiWb
br3/23o44IbSmcHpkVoZpUe5B98mkHyzx3UaIxVUpUxwXozJSPPjvxODs7grFJEM
LRnwhNQdMTXKVlbucwULcyJbxsDr3GFhxj3QYEHXdOxIvKpXChRjncscmJtlUxSI
VAUXSzP2mH4gdPrTCbziL6so9haES6YIPuLoQKei0jGCBfj4vCyzOeDiMcR4FPRM
bFlBY91eVbdIKsAEN4RKe8Ja/lxtdcdDmcZ9jabSn3GHlyzOojntRH8YJMAaXYxA
WWcB4GNfQ3xETxqqgkesa/bxtFne5RHnkj5i5POqn9TAYdHUXdo6QfaRss1OAbs4
paEnxrr91701ZhMSFEOecJu+39h5gsuwtxwj+2tZU0hDCCV1R4dHZ3RiiomFGpSO
p1TSbn7NfEXy0wmSqmLm4nVvPFEL2aBJPTAXN3wFF96QbzKwLQdso7bveGRTqn2r
R3pw9SSIeRoesrQQ4/z0nGRDA5xfpZoadmnVJwTXXBeh9QLbObFuVK9e6AoJZ6h8
pTkB8jlx3AqONphXu1N/3c3xFxt76he/YMomuYSIzuwVgFLnAdWHo3hQwfoIOSAt
1Iz5cKQbwgs0myHCH10Tslit6bMPdy5B0D5HlgBXsAg6TwKPRA4+gcrg5wkHS5fz
5Jl2dw6JRvul6Aspr/Td5DcAFLUPUwW8gxCzQBMmnH0LCR33Li3NYom8kY0/VuCX
hzinRmDhgxNBngNc0HDrK+TrQP6j6yFbkcrBRPxGsafBN4wC5X+D/JN8FwzE3L+N
PfhK9hItou8sUOyNsKL9iYy+Y8zNCN84ks1ldNxesMLDwyMIL1M8QH0wI/1vx9cy
h1YijOpJjpKlD39snVpchMIWjZp1x/ipf09mqYCJgYcFr+rrCD9LfPnJegdr6PFz
ByfADe/O3OXtYVKR1OQGmRiaba3phlNbyeTEp2gLQrAh+NfcDdJn/gxb4riThTm2
1k/1b0kUgEz4osariSO+e/4XQjVFsO6KPyM081d+HzjhEVV680h3EwovaW8/a0gc
3RX/4WjsyER8wNqgFgY/Pfq/FrJQ9ZR/NpI6tnhgKfL+GOOky9NAWeltzQMp0ELN
EpJCK9BZ3y00lXC7gBTNuYluM3tTm4Z6QvZxhgoCDR6WndieMZeKFcMl/y6lJTrp
jxo9t+Cck1V86vWZtl6WMbCeaJT7QxexnXTj99MxTauHIx5ELOwo0G1P1gDNnjFk
QPF27ysB3GCYROfCNxYeHKArfcea9Y1HVNmbgOYX7xUMBtTuVNaIKkolESELhj5+
8iMjiCmHF4I0gmOtvi5uY9CT40gLkF6CezK6uAvqQanjKyN4YiX+IdED1xhcr5ZN
InDi3q1UQK4TQ02vjLzz0/NxnRoufwedvDwl/zxQR+gNK6vz5vYxyJoHvcsoFP7P
5qWeOTYTeRCE89Ds4w8SMhKyRsNZwmp+iBp7BOLXuKIOHdz8FQUUC+8bHpefr3Xx
Z6ozq9AoVghYCaLG+uHPEobtgDp0QTbq0qjYMl0LgKMIf4aMzc4J2wdVYbyuj1g3
qJYDt/VgTMuI1zMuBM1fSg8+HPfrn40q36PHnYpSRgT9nWP7N8pOzqEolDL2OhhS
/V69kZkt4zwdwxXTupBcOqUUCg93vJWJxLTQi7wb5ZoOLLB2rbDLG2IWyVW7g19S
mXnky8XVq9lmJtY2/SX0rosoMIwyFeN2eI7iCMHOWXjDYySkAa3xqccM9/OikUSb
2hMCGN5fYt9e6TljV+K4zcBTj55m35C+tCkaLFNTjGP209YiEOwt1f/jVbG5ENK0
Me+ieNHUsFiZntldAXboB6W9yuxqTbbJB5dVOIxGgiDbhqj1g6sKPaLZcwPb7O+P
WtltoONJ3llsKp8z7LibRJj010Cwc/n7mhSlb3ZDNWKpVMT8hiqFxoP0kv5OIRUf
LpSoH/o+NpwKugC6JssY3vDBMv9/XQeaXbPt4389tBcyoiLrR54KDXq7/nf+7yif
QaA/od95hRwdlqUEGCatUkgNe+usBNvWZ4qz8kZrEjnAmB5y9JyPxCuwFya1wEc0
brzMDRe8iDO4aM2MAy7vGXHN7ozWkSr8eho+UlsslQGicrtoAAtYVgKa/q8rOqwt
7m3eutLHpMutXESylkZxvmdqBbAQ9nXx1tJYjpJi7paLBKafuKGNNAtvwJWDoLp7
ZgE33hS/ybS0IKoROrnKCH1rT2xMkjFNujylFDxSov2EO+zIFaB3uwq0i5qRAh5w
jrRWFTOuSTTG0edu4+yN7ZNN7wYKzlMah2mj723622FLH1gn1Cn1/YVxpDXu8SCT
CwxPNyj/ABNkiEFDhty9I23/GZJk/Gotrbt7H8GD1xWFo1pMcnmjpiwl5vZynoem
LhNNEhyqGoKP9lo0n59boff5FdM4cttazPkPhxlmwpKSyEojXrTmYQqWeWbfZ3aD
JXGlKN6SnGoN5sXLzIAUC8NSapX6STjcwFzn41FEymAVm87EoaRi6Emb77R5zQGG
XnfAuzcAF4hg3IHAKy2Uwd2jEEn9yIKdA6BMgM/gsd47qqtABGQDmH3267NhyAla
C/+gxvLzviWZDpKjM4tOrrMiLfwC8y/1L/rf1Mb50yZ1MiL/dbXaP4SI8PGkRMgQ
UWQISJzqu8u9ex8kDahVQtwuvMwMvAPDIHM+3q/cGkLmJpetbVCStiSt8RO1gmrK
2Rj+K1MZt8y2jngT1fHryVijvrfjXaVD30CjDFNLurQo1hSUGdyfHstwQrmDaaTv
ahnukcvgQGTEUpnsZCPbrHQi1KyT+E2F8JXks9DIM+6YRInZ7QMitzLsbBNcQiQ9
1wzKQ0IfHsf2lwtWxPZmWZ59riFNXSoePgpUHZXSt1h3yR8TZ89T0pc36HxtG9BS
QF8ZPSPmizP25l4yAyzyJ4T8toWegr0/v9I8bo41PzwUZsgpWLZ+qjj0Efq8r+mW
WTHwtoJhxSlI69yciHfKSWnRRP4/7j9yByJuqLpusPy8BYp7+k1VD+lrEDC8aZyU
U8cOnBqVRvATVqI5Fb2yhFNWG+GJbCryrR3YtXWst6rK/WZV9Qi2MJCh84bwsiDQ
3rdonSnFUXr1pkjui+oo806iyukBsc7DBtXlfcGaV1Frgkwh7RclALb/w45osaYU
f+1gx/V3cVh/eYjy7qd72I3FR2td2dLx7XomntC/qEAVcgsnUJniKymHl7JwJkE7
EbHFzOlHuflJIH0XeOgUeASeibRRBBexbHtZfNnQ7kkCl6vTaNxG46qLnOQgOYhg
ZLtmUIj7CSKpg2HFKn0uYHCvL09/2NtAClBKLgKetpskQilhIjqx48vIo8kiIT+U
1tqMN6c4UOVfGU4byUhLw7K5Vdt0iZVvr1unStZTSmr9o+6WauJJkYEx0qYva5o1
nPf/MzckXm/DAedO62Sl+AAVqz0Bj5wrjgxTlGEDBBqsmkHeOL+vS1TSJTDdASC0
giQ/875TdFpaLp3EryJFLr1iA3GMh8tYrz+OVOYni05nkJg9iTtPpvWnUDpbcvoD
WQlede8DXHzaGNWU+3UC3nPyw9cdm1YbXw7GrmLdjGC70XhjjsDkYhemzybu77sH
B9AVd9P884KhF8JJsmi8i7gN7hR6m8MPSQgPqLyhmElaYSBieNJpQcRCih+Pq2Yc
sCEEU2wTDII47NYr3xGGl/rsYuHRvXlAKv9RjqNfGZMeofUZDmvRyD7F3w3XEwuv
uMZHVmngVz69S81FMA4M5SCL/cyuy564+t/N0wTJdYK5Tggw35ZX7QrAj8s9c7N5
ZSzuv7WNFVzxfNwWR71yPkMtPY5ihb6hTTlvf7QETk5IQbgQrzDZ1bi8ZSdbU910
Ah/b3Qg0jlAunbX/rk74tol7sMFUo1xXbxTF1IT9BuZpGaPDTe/Hb+A0BjN/94BO
4/JIq3ZFdDcA6tjcl0IfwRFs47Sxk1pMcy2WKHnj9tn+CFcgz3jo0r7vqTLkLDVU
Uhu1CN7xpJ4gtE9lXKAS2DThvHOV+GOM0T41D4jWgkzSW4zOw9XNCZxKQkRcRkmE
DGAfSyzqQDiUPnk5Ivbimx3FsaXWmg4bmhv4ktMEFdA5uUmilZK5nIeXKcHYWiOX
llpnJVs/Zc80Z/2b5b0hGV8PX+nstMtQ0oqdq2LS/yv6LHcmO/og/nfVMKaavPJC
7+KjDaGHIu2D6eXh355e/MNBULi11LrSSt5Hn+eNXgjGcsIsogmbTPj8VhJJh7Hh
21NXef6ifI7ng3S+yPNBHx+lVcjsWB2FYflpdXRWxYdVIfEbmwH6QI1JehzVNOHO
aOzjGM2XQqFT8HmrKh0bRfzYrc2W+D8PGDwUX9PUJef8zO+WVAd6JahcviAmfcr1
rpbZdHxyQMQk+hPG49I5uJ2wKpSn89gg2YP5ELJGIdUEbG+OHmFW+wHOJifRv8K5
KPIZwcqwMmlwlbRWp6O/QFjKj+eyZEPk4gliId/20cNwzzBhLysIpfZYcFG7YNSL
5MT3EE31vDcWNXMm79ovwrjOrBkagcGt6pwu/7FVXozVeht6cZvc7ExE3AdmMfLA
blLM2DpWXwsEWpLk7CoIo3liTtOCEYzJg1fn4rh8SaB0k7hmXNR8XlZAeK9nC4gu
tRV3D0T/eBIwLq9Gv/Mz8oE/VKtNBm5hXaR0CGiz1wdTqfyI9yOkvrvQnuatHrw6
lXiww3xeXREK4MRqQfXPoB5o30QuY33JO+grMhUhKnlX1UMZI1CdAITbZbwjeyoN
1tzFaFjPV+F0+zfGflFZe+eoc5HH3tcCo8qoE8/42J5FcnNKJtokWXvKH/puA2Z8
y25BJzJggYbLCLj/mwh8ICft2pTkcxh0tWtWDjV9vH2Lyg9rt5KBuHXh581g3ucm
rOWbMmi3Bdt6IegveKUjMMe+q0d3IkGzeqJ6MiZUDHWgJKDDf6mLe5K8anRnVlqc
sDFkvp1T5wUaEGlnfwhdyk81wpFc4TR9eh7VxGvl/ilATcnSNm0KohhFP2OOTOUh
T/B75oZ+xw5Ae3lOjLzOM3nIejBsrmvNjqFIEY0dVbcYlrZ9bLNwGcRAERgMGNv+
12+OHFCUFowFkDxxDBEHQOBlEF+1pBDPtjvvc58K2b45Pldo97eMQjfxkY5F+sFd
F84xrKcG+/oPyREJTkOeePNQlXWLX3Bz5OGXZduuLmiFqyEn6svgOnG2S0LCNbo3
pPhTJEsu7VuV8pfvoY7btq5isqz4IaMON6Kkf3JE/VdYo/4FWJ4Wy0q73njGORnO
70O6d3GGhNX461vM6CG2HjZhCvMUp9j1bBaTk0TeGBL3w/UaFCLnR9ogMVPV31h9
CyAO9PHMK8usMjdqCiO3wX4qUFLdTVpVrqaf7Wgjjiq2TYM0ny327DSXPZND2Hz8
pE5oi1elNU4kuaf8Dzaki7p/RI999dRzp3pLTr2iLRMCqadLsoSfcLJ3p/YeOwjS
aRdUVqFgMXQmU/136nGrAfPY0FKOdlk4XMgECJG5H/pQlnqLCNlQC4S1bfYh1rG7
7Y3PhtH7ue1i5RIIlpApN1tH/1Jwmf4xR+VuJmyzcgmOyyzfsBiaShUz05e0lnzR
uh31nOuKp193sP0DLLcbig1ME8UBxXFudQfAw4MYCRIWZFMJF7iQ6FYst6XVjlWc
6SwBi6kVJ5NEgVCnq00BjCIxGZNH2BoNczt8jBmpX388eB2DjnBXcwg/B/o+eci2
4BXK13nQQlEpdX5YaP+/XLA2nT+By6fU+TadfdJ33/UqcPvdlatze3Bf2O/+PKUr
1uJeQFNucdKFP36rnzUP1h3XNsttypc3CuosxaKE69bs+uoZbTMq2/sjYildQmCn
O4kFoshFMriAmHWjuhhUuXu5a7OMVhgpQomqQ/Xzs00qAk2DbP/4FReUWwce/sb7
v5vitOWtthLpy8/lqOenVZ4dpkxxxSWGiHcJPjBT3z/lNX92UNa7kSGH4mL83kZg
eutMOswPtn45SKH+hd7EyP451j02rwZd2uMu+Ii2lh15eq9gO30YHdht85y36SZ2
qu5uVnqtjB2aJVHyCzvIh3P1cPTv3d51kfks6niiPha3nZFxFOxouCFQkS4sk1fP
o1RGioPGePJOnJZYeQtfahvp8kuAvC0GB1bQPVPaZ3lsIgVj/TBGgjcf9XLp4O3k
PiYr62D8YWT4V7YKqEQjDfZPKM+WDvUfTDPnVvj/SPHDLEcB8FyDTOLZdaRPkRlp
h6LVthIJbipr7yFL+YdzcPIl2otd+QkZhr5E2YjtNQRnGSNtWkPdqYyt8ZqVLfGR
/KiGmm5Zu4xtxmePlTUyl67BuabyXbblzhFoRImVODzVCzVGs6tPfVTcJa6AqUbV
tSYU1fQp1Il3pM/ccOjHHHj7DtF4ki68K2ugxUMHzLidSbqCV7IivtwHRc3xdxtl
ambSCPubm/NTb2y2SeR/vkVwFsaiZMUWp+rCFLyqpuxePVsQCSGrG6IoLOlmAStz
Q22jbRByTbta+f/5ZcqeeIrc/EGckkcVLw6p3NKzP8Q4D9MxCtFBdYw4oguwxpyC
yV0cvvADcJSRqwVQt7mV5SrwMD99Czt7bC+u2cWsS2WSytcoueTXY6svGDL9gIyi
BN43tLjtjxEsMcYlSTff3lZcyL6Kg6057cQZfvSOqF4g555yRLVwyau66MGSOXd3
fTOoBy9b13xxEI7yPRESlYmI8iq2B1ITyr3UfGg+OhVnoS2hZhD/E4uAKFjIhnNs
FuyJll7lAfTTq7LHi+gz9k8Uz696PmdoKwEB+Xniu28e4N3HO9C42gYb1n66I2P6
Tv7LfAzE7vPVWPW8MHqaVS48d5t6U/S6ang4ONaINh4DIps9UFWVajRQS+6ZMj5a
2nweplhgmy+sSuzmbdpFV7amIP/ktSIIHbhPWBrnI1N56GFcXKfIXcueXK55UuWy
NUKdHQt6IxR7dDAvnX/oBWQOwQjadrHNeq3UP4uYtdLyN3OghRbrp46AG8BE50O0
m3Esv+YUUeQUWQxg8gnVAi2v6eDEl3gVR0qhdAwYryElr8AnzXWp+lgL/urQGg7E
YydOEN97IJtZ+CN2Th453+C0G8sS6e6I5r+3E7NBagTgKlv4Rk3pETBtOWp1aG/V
Lci5KR6r66SOat4IoJg7S+jJsXHfO0YIfew47jZOOi26YN3VARPSK/oCJr2qS0lw
cE0J6VBk/RplWyFo9k9WVnymJZrno0qFdv4KuE2awZGpA5OwvvJ00JG/0jVxjMWi
HdjndOqrtbbZY3mMivwIj8wwXInt/upjWTPXZ6YUfR3OXdvnQzXaj3i6K3CXho8L
EyVfJpV0q9UwsvVxRyFPfFoaEbZEPATFfs8bMSH7cBXcRBgaHk+nuCN3Ut8GGMft
pNo2PRuwyJogxC/6HNYGqC/YIRhsFK8zlcCmGxvfIN+EWSYVSCkNomPzh+y2nE+f
hF7xHL/UjE3Y/e/PLbq2JM3p1x+QQNh/kAp/5/yNuAC8TvprXsHC0DtGiszX2qzG
wSw2aWyV/q0wa2znfZSEia/TknFVYz6DqI+HuXLf29vPIN4mGUeLZEbnO0lJa38h
v3UTNdEq9FOirB+P4DAsTzjMHjRUqoAx4BRCTtbUFMGNmie/Nih+BOLej37T5/mc
aCQOqL86lTAANWoS4FK176Dk8630b9l96YGiLGEiappE3f1JgLdIsPEDodqky0ZR
ODXyWrsGMIQCRfNRJD1tSNCLI9ZhJ/kvSvx2Sh/AUl/MPrdhUue6+/qhfXF1h5oF
jt6WCchVhDyK2g0lMrSW5PZH5VN5LE8k24kP8i7vDZ9Cu5fQZswZREi3ZIMoqiOE
uoSZUi6Y0h2nGlbjvnQUk76ZBGliF0jr9o1NaA+AqPurmYBbLJX7TSgDmv7TWbML
gSlUt3rMif97s9oHUF6Vn3b0qM1sjvJ9WHSONHbvYA8a7bu8LvIaTjYt8vNFdCMI
uoIlYEtCfxlh42tR8ohZ0u2fa7YVGRy2Hzftghb1gFTvztkADog6nVSlM2d7Wk0K
v28JLM1NMRRWQ50RR2pQBNvvZ/zykaHeNVxrKs74bn1KMNhcVKy9LlAge1SQJeqF
m0UF2C3oy+WoxIVCUncl32huI4faQUKsSDKbb2wwZRnziahWmAnqjYwEU1zZlNnm
xZjKGckL2loaNlR/sA/ia/ev9hu7AISRpG5Pv3vOwo39VlBc47amkPP6KOV6X7VR
vS+W49Ak+eTxqxskcKMp6Ejp8avkbKPS+BhCy0akG241pOoo7g3hvdlREF2Oieqe
S8eurlwrdinYWRSCXAkMBltG34dms319YvA87eYSPOH9Gq0vs6YECXzmVa91sjVm
uF7KonPl+p1m/1DEZhHmi53z9UV8lrDXfbZW9H3xT5xswq80WIwBwzyCuapw7aBX
g16riwEyob7Ax3iOuthbrtpRYqVscXSy9SjjGwvcfabRP99PlNm3oa1urGkb/HZM
/HNf7MGQw2UrkKZYjiJY2OrcmQwn0i8g3FMznHDlupbHjgff7DHig1AAgbtKpOzV
TBU0E66l4XhjQT7GwgKYQxd3xP4mhcYT6CXeVTSw/n1kocs7AZayWzyMr44ZADn8
VkneOPvx1cBAc6jJG392SI73fJxtVaUz0en7x6UtEy0NXU9pvMKsMjbnL6Sp/fh8
E4kEATZ7J90LcAAhTffaCaXB9uCvC8IttiCxmEn3FPDoTu+YiXyBDf/ZaHBkGhA+
bAR88z8LrwneisjL/s56U7soL8mvC1YeH/BnFJbWu4G3TRIsLA0SX5H3fw+izHkf
zd4UgEenybgod8SniCZzdL+oELPmLjWXBNXxwHWnA3MMHKbvgUHOseXUepp7P9tB
t4YvHKPkmRSqsE6N4eQUzxvqbdHL17BS/wn12MD8Mb7+XisiSV0t8ViOhB5VjNPQ
dwwMPkmhw0kB78PZxQ5KBpN9whZS0UJ1M1ODxIlBp1gw8zW6H21CzbVcMLdEz6eh
YtrqcDC+3wSNa2OCTcQEV2Xes1t5euQFv2DqrmxwX2f0OYMIVjPALQvNqWph4ILV
wQ92D+yk1HX7kMJavgftGfRpu54GW4ZKLRh3ly+2SoyVTD4S6ZH7ceIjXLQNyEYN
vZZeNFAHKJXJ//hSEmuw8pgelWnP+dbyqQEOEfbA0MT90VCVzmVo5PIqDKWNEpd+
8Q5OYRtIyiURBoPwn5v5dSpgOe73h+U88KLZpxqYw8oS0W2ZUYbMbTwEz9NZmuvv
lJKBIcvjgohdUG50gmH1/Sy6ou2OuF5oc8111fVpwsydU+x6fDUfMhM2IU7WsqzK
SjXqC/u9eA/mSv8MytiFFMPAq3fQa86ETL7ghZ2rBGwGC2HcPP6LmZaIizbZlqu2
H2sJ2yWYYqBh2epO+iRyteESxLZU9vYoY4ZoPBSDnbXjQTht8AcUxIlVZihbWw3x
d1TqYL3AI5fzDT7RoAZUbZzPaTLYyqngFq8ZTnZzZ++hCgz7FDN2ct7bdlAvPLOm
C/hnlBM/0WM0mciU7RIIZepIy9Mkxyp3ima8BWp3cv3bfc/c+Pj4LysPtGsroigL
/ZjZtfV2K46bpfm/Xv+hTGmQydFfauRIX+W++P6QXAhKaeJ4Iz84Yk1Fz3+mxUGC
gpuhTvYqxZtAMzyFI36yWYSYoZfB2xCvIT+doYCN9HK6blfz00CShC39iQLGRfor
flXhl0H2B4SqN6hWV2uh0mfxiLyG4fVTXBWPgxBZTxZrCa9vDIcECmQrv3Zg1xyU
YvMZsF+SLy5zgQc3q0nYtXOAvXBR90JOIFHe39sWmTOLaMDNFXrxTczdv7faJ2+J
AqFJ4NAj2y4vLf8ZihVNIHEoe2kD3WpKAARkpMOG2fJFuJzPBRgAMf0ig+kdOzqR
rOh1/duk9fcR0vyua53qkBHMQ/4gkVyL8BIOut6jR1SX6txXU3aEIqzDu9t/g6H2
uVjvnhEzY7XKCKOZjTtxy44doN3dLLTHqNN0baq+weeQO3V2vlUjN93hLnJCEN4v
Jv+HUtzM4pzR3nwSzBLP0K52ZJKF0qKFz8kdomHDFi9Xff4ncCnvdWeBcf5CAmnu
XOjsI6ZvLbXDSEnKb8nppMmks7ECPpWU9r0RHw0oV4Egh/+M4sEmqT5s2Z8szByr
HUf2u4YwFRNvY71cG23aibAI0/LjvfypcP0xM87K1VwsprXMsSukhIRssTVLofFG
N6Y4yFEbXqL80k+8blczXcXRFsmqIWQRmbQ9V6b1IKNR3RiVNUIfF4GHvltEs9Kc
sya9DIMPSByNQiXVteChCmvhniSd0nBRxH5nfCs5o3+Yult3EyOzNjRkBdkOecR3
MENnnfTYXWzsqSJk38G+3Z9qeGYcPN8mhQxr/BwcrfmY+WqJjDL4V0Mp9sSM8Qiz
BeOoh4GXtCbj7TDyQnbDLlK+8hhU+FkGtyQOn2/4+pL84jsVX1geiXnccD3Y28h5
SBMVmd9Z5SLxG3oqSh4jZJnAg+0md6w4wZeF8AT23x/3AS9GVPBvspMWXt+mHgpU
59ln6gKKufWJlMXjlTvAxAkfVNL0XZDkhWjiToWgQRi7+qN1Y0OtPVF9jJiQvpnl
xXam/npkLT8c6NwgRLOLUMrJmEEMMQnc8NA6G/phiAougmZgiG0LLEM8JXN79Dmu
fDiEOIALuid5LVs1hUBisW19U2F6jYQa0JDHSqOWd1EPR29ezj4hWuv6hCZM6I2X
wtoI/Di/i9OIVr60Kl3UIcgMfcGdwyHTS9zGIsaddmNIBbVxrXhsD6wTVEFseHZf
K9RvNfoVlR2f4JV/awng3CjNWt4Sjb81xEJWXNZcwrwLY5cAj/sckwZGvBMJrtMp
aUiIRdlNLeK0/CgTSaaN8ERgDZpHKCpW880LjP7zid+ud9crB7+8yIQCsw4EI4t8
tSS1v4wVg0BjFlX6rHdFFGzVjO6/KtbaLtsq+QZ1T+ksQvOP95FtbpT2IHe5StAL
rGcG3849cDHMuzrN1PvNJVvyjNwekfIXgTWjWIZ5KzEBZxzJnnBmiouxHu/ycNRJ
2ljeqKj6N1PQQzJq3vlUrwdWyQSW4OxeEZP1TYXzH/L2k4GFbbOCgCiWaOnTWYcj
JUgu+jyamacJvLiSUfyki2OscyKlhvxXC4oLX4aQp3D9azlAQ9nt77Aadpz+jZYa
RUZAwIJ34NA+QEKe6yJOw0Z4XKpG02PGQRGX3rBwsS98y+rFmZKC/2P9dTVwW7GY
vojyz4qil6L377jEkp7FK77+TPw2GB6ZTr9tbBHt3UhQQzAy88snp0QnTPvzAFuc
u9B+2OXkBCsjfGPaR6JSplbY5I+9pGs1MeASMn87T7ETv2cDg0bhkclFrtFMi3Oo
KxFsurijSMsNtQVFAID6xQQOpRoO2ZjCPjMlMVdxsHvViStwvNTe9i726ffBsC3c
WsDv95MV1/o68CvbZ35inu4zp0qdOhgbs9btA3iXE7NQzYZXp/uX2On8FLJv9EY7
J6L7aqYfZVz3dQZguO7WopGcL95f4yeoDsV02zu51rFB8Y8xDyQascuaLFA8TrF9
CDVgQOq1jIzDss+kpm+K75d3Me75Ko1esM7A8MId+nVAhuKM4KxAUE70CMtC/Gnq
XSH58eUl8OvQjV/BARrkKeJtYNuKmjwXnrks+16X1asFrEhggGKyVzMedZwlrNHe
BNoWdS7e2h3ZvrWoqYvIlljP6MCTyeTktdSg9zvpw/vGO5h8eFb5qWQiyQhpmx/C
cx+XriqTOrqNyss4i6m7pSkYALCddAi+r25lTWX6/WPSg021T5MXcOUnI7Qh/mRk
su+/mtPeDEUpCL6uApb/QFCcE1ypw5D75N6Y3ejWlVKofk05DLuXNnvrgnjlydAQ
fjKHVokXNmwkdOqmMFlI36LpH4VuhdSTeAH7whOIy3jj5GBy3VxGQ3XjAZcAnoVG
pMuvS39tgSEKbnQW5kKbWFDQnif3NIAQ9w86DpOXnf+733ya4nEKLVVyn8LfmNHy
2hETTIACpp7VeNX6XHl3BKIXD/OLg50LBmjWtVy+iYuQ2+YIeLngLyhSClYt09FY
5NB7gb+UdOwUeKTyXuzJinYd3xGud2MOSGbtAzLwKuDYTUkNPelrMXO0zTR1uPka
6N2JYJyW9fQ5iCSZxrW6GzGfbwBsHq8P9knwuUVl3sbwf4T34VhhVa03fx8RjOZg
7hnDBTZR7HF2PvgR43A7bGRaTrbHPWdzD70/ZOUoiz/kqglS/iBmdUtKNdWYQZ/Z
D9g9hvh4FoOX2B4FI1AWtlUWHS/ZYK+3hlfbegFZubclwlQ2qJpJQMT6HdAzthV/
ZHzZATJbOknXJ0q0rUJRIspVQ5EyPjgFfj9EJ+HQatina9/TEU8kU4LOD2atJRAj
Ae98tDhctvX+Nbl3pXhLgtz2MCUsBR96is991uX8iMydhL3f9qxkkQOaJGFf2XM6
RfkP2HzCEBCeN05YJpQ/wqNWAetd5Ed0GUtUudLsSoDUHTJ+NeqFf4OVzwLENQuT
59KNc8UkK+XJai7VpScudTI7la+gVBa1cWasBu+6+EjnNnEwKEyObU13k0V8tHIU
B1OX7gf2ty7EoqyGHd7CUVFlQ6w70rIxeW/Rxl9AWoJLIamXFlA/esfkWVrq5TLE
zTbS+2pN6XB34tmxBG+zJkfQNwLaoejpCxXkideGb1uFykhFW/tET1aBWf0PuD0H
mF77WaxWeChAyCIdW+nstR8HLriM0pkhXhUvgunokA6v0vqJypIXudTk8wY7Z5UT
S8r8m65t+OgZCqMvfRWxTbQjq3hxg533rUmozN7uCJn+jUGKsihX9hi7aKjw8yss
UkMxOsgB4gfHbCfN55F1PwaAGAG3iOjf0lhLETyVJKXTj8S/LGjhltJImJdrL9zu
Ws4/G3iQzatFlvvJa9mdoXnPmqOhFzbOZoJFCJyXE0JJYAksnQLQ/VIcuNAf7YEe
wWrJmQGtt5WC/Y0EqbHLyturHfWcKLGDyQqRaCn8bqJaUE292TthpUT7j93zq4JM
zYSQxzfcIt4+/1XsZZ7yhhvKY2hc6kEr2CtpkBV2PPhdWYoSFyAJgrtEI6VR2xYs
c25ruXIq42ttkVKdOG7rVSXQMCuZZULasMF9tL+5xsDPd/l/BlMklmJ6PMptbPKB
FTlH1QajUBRRmMJLk1UH0mks3nFMZ4tnZkldHM1q+1YoUen73UyrGKrthJ9hFRzE
uUq6ZXgDZtD3sxwVA+BRFhP2aGR7q+XeeepOeR4jMSn1Zs+5s7mr8qtxAt+RnmBb
cvYoFvuGaRrHgu0S7DR+imGOwInndKP5Y0YfTpjrtdxA196+vLrHkLeJBmEUnFsi
nJ0Iq+XWLw2m6hWnMDsiMOmqtx35CHOGOg9pKjJE24ZQiYRdnUwB6CyRQKGG2KYs
cFwiGfHv0GbqD2A4uwly3aHjYsZ4BOkj69KcZ5S63e9bVArDN9sS9IzaYI2dTWpB
iOFxY8ovCbi788LPyLU1cM9gacQW6gLoaA4cvjnhzAE5P0n4NX2deWWk+PvXN4SS
+cZPAsSewAA8YGnzLUInN4UlKgsPDfPCJFBu1qp6jVDevWGURVtPM1Sdr9KQyy+E
nLd72kFAbdhkixX/zFlKGOrr1Jo87TTACcVzQgoDKJfn6r9I+l1HJ0DSN+MU2yni
CevnUi8fa1S8hvHojyHFdvSgwT3Q67x+raoX+EXf+mNvPbLBhWr6UKkO28s9aVts
j6DDeH7gU3ywnOhu05NL847yfljEVZtt47uufnmypz1nIKQAF+lzydHKjVQsEURx
vg0B35lc86wDyu5aDSwWoPi7HzJViiVU4M9woMQqoOOcZp0uXt4yiibBvGEeO5sJ
1hT614ntji1mnstM65ImXEQlsKzJwTHI/HinTkSOoVns/NKnjnLiMrvSaHKcPG3V
s2m+DUzYxwFcf8LD9JY/N8PfpWwxz8Tf5MgOqKiMwKKnM7R5IACVSRhwiTg6KSAx
tK1D87xUy1ttWHFqAFEOzVYhJSdD0wloQnVU/7X2Omf+gp5Z8Ox/BTm0R67znazS
46IC/wFqI6OSkdf805LB/ZD9xv9qDHgDnR/PdRE6Nh+G1qnmvlmuAeZB2kt81Dsv
+q8JCQgnAtf8WyUa1bV95YoBciiGLHp2CDZnR8A5JTA7oacpa3te6gBj6O+0JOkM
2VSMMKrycf16Nl/FbKQvlMtkQrdu6TciITynQzs5gPPD7DiSV347CLMxtTsSRPXw
8pE/B2i8YIes/DVWccTZUc2W6IZB2UnCue6EBLTYCheFz9FnpKdiyg7/zxGJH7X3
MZkjz9Qu6R5zYiS2f4JFx+NTCk+Kp93Gv4b81TJ4bFsP50P1SYCGaMNvbBzW+lSL
E+oZoIDwdNrwzmV1ppz5PJsWkRQMBXk5m1oNkuDZNQMGcNWSKnn4156jS/M/unf8
u/lxYSBM6w2YnV25y3f1QMh6sxKpEsWc8LzTpAAran1Qx6ORrGLCf/2m9xdKdvZC
jsUPgIHiRy5T6ovivoij85qAaek/77a7aGBOFRgXdfEELk90I4GucBRoZQ0eaZ4h
pv4Q2bFfLOpFRVmF7HkoiFifGD8xyawMR2i+fBuRBNG13JQrhYm6bGqmtjp/03Fn
qOxX4Ku7AkyYKQSDuLJ9UTeolKw/1nFYryOLOljbLYPifjmQPv2HwnNlUZj3nRyF
8OBK3HeDhfOjBju2noh7KOwxuIoZaax+H3HHCuNYTY0kjDL7gx20YTcjha+cPtun
oTxma70PdDZ/Rb0uxB+E4mhJ/y9SI/j+dHHBXAEqen9iBvdfZLYNqr5wg8ztaAM/
tH8FQLVxq4MJKMpjBfM0iYqtvxkXSmtwQ/dX64Ccs+C0gBmnG/wB/H5nkS5rKS+F
g05OYmU4iYpuQtN0c3ikp6yx2QxzY4e3MxC18uBKXoEJGiRvDfWwMOMiEKck5/YZ
c3A7QDUBgc93Yz3dlLbFVB5aJdLAN8zhNrzHd7321BVQaIwxD1rJ+jhkII0O6n5u
emujw7ESYjIA0MirmlLH4gsdI9uky1WKLJTvFYPbtFYiuhc4VZXvHY4ZhvqV8x+y
EcLLQ6Khlug8/Dj/51C/fSUHjRZNayoy0Th1wrP1UGaabPUY7fX357D7BM0udPIM
+K50AyRS28Uu+0gqFJlsffp2mto2Jyrahif6g3OTW3dHnIt0bYLCZOVbPaS5oukN
Q4/yUUuXKo76qHQSY5co1vZRzEtJ129r399kIQl7BZTUhBV/PCBUtRhZEUdwgbkU
R9IhBuSJW9xMC4bZeR7Hy1u2y30A1tI7hbisOARPe3ExN9Ur5fAGfxT+2wxEGWH2
ipJ9603NlAs7zIY+BLvu7Ubqq+2rMKPw8CJOW8c26daQABIeZrWeRKZdbxnNhRE7
T8+ctTx8eavr5980MktCa7HpBDALTIwsbn9t/PF/0vSWiEBJcbz0jYDZfkA2vigb
E3NQ2toTwChwqanf6Jn/lLZNw+NWNz2evfbZRJ8Q+ZAFUBjCGMzy6wNc9QfVoY28
YqiZdKsgi/+Nbg20VSBac76iLRPHp4dSzR+Ulyn+yw44hW3B7CGX8Vzlbv2FvbxL
WEJw9cgyo5FPnxfLjJkFzugdhGrZLfC+oO8nI9D9/fIliCDw7CNJLrXxpoO0Q73C
eHCCS7TOS2qyxwyTm9QFlu7q3J9za5vspafGYZc3C+Sgc01Wb2uBWxIJ2tfqRDHf
aKtZwOsMwaNYreg8clJpA+++Dt0m9brNjfIeQfWWSYmxnUyK9EaIfqkblUl6adYb
BNsj4M4pUlFU6sLYoyadn4axCI2W35LJNqnxPS8GjtbMtWc4L7MXQ9/o284GoBwC
W2RLMHiYaRd19SqidA24EkQai59QaTzoY6Q6fsBmFYiMdLZnhdXXHh7Z/5DSvd3Q
D+e9o920O3JBANaS/xbqxl95Raz12eRWGQqdNiiDPgqtLcRf9FWVQzgK6A3jRLcq
YnHMxkFXd8sLlzTj17HW/TVUCk4wtTBnOXpVgcwgxQ8n7BlVIIEfslZUt/1kaxqU
e3KtvrXdEixWWBHoZaP5qmPDuoychOfcSzYcTT6bGl721UtEwNmtPAyZb6golwfU
NhixmEHQa4nSP67Gh+CdXGmdLgnD0+TpnIOCeVkeg0gLv9HpfPZbkGh/1fSzXtcc
S8qrBhzWFJSNvQbn+qHGJfYem5RQoVnwax4SVMjVLAVLT2vATPyhO0Xo+LH7OQ9T
Mbf7TOUGgqg+2Y/2yMs4EGIdsh0jeAzQTDEsJ9j+F7XYK/Z8bvMAJ+hHUjxgTFxf
MVj/nYAiW6Y0CS0YEAWrRGUxql7i3vG5DuBiKylR8K0RF11aYw7d4DZ/YvWg35xh
KWIOtEIZVGZPGZ8FezeGsu4NZjjxrF5jazK4LbTHB5ngzKDhx+Zulx0zD8rWA+OP
ZDTfLYtpCOyANAAx71n4PqD4S5RnRX58KL4Vo9m7SCkqXVe7DiHhmEO2dYoEmj2R
2DYlKcq7lNdZ6KNAhvH/JYQekM7Qt+LAjua+oaQi2UicMoBp1hUsOa7fxuNI1BHR
Qh0HZenOMnw1/zE5xvbVv3ZieqA2joZXtyVwTQM6Og/Kox6MBWp6kcEUwdpq4Mjq
NeaQe2kLpa9ZZaPx6FzEhTUZlTZ8mKdAIv9oekGcSivhJ+oD5yZc8/BwwYEAZ1DH
pGLPk+tNgZHJZDJ5X9Rx/wHcXysILcu4qQZ/rjvdWLC6L9cAaSDPvEKYI4m7/OT4
gzzgl5TR4+hEZR33YT8Na7+Oj8IbgJVLdetzTCagEfMiOKR+W4l/O2WjJ7EZagp7
b9/Xzto1nZcyhX4h+en/uOUU+1qlDNlKqJN//UlapE1ibD+zgs0RjtH4WWtdf/9V
OANSmSAa6hgf5Rs5+mAgbDO5Anv0RVI/UigTRcF/HNPYD52JIf1HLj8GGw8nrPXE
WWUAmeuRdvrXjYP4fS4L+rLX2s9vLaGaNyO7CB0HNyejoaUBq45bUkbe6I2V3vRj
7fdAasn0RbphrHnFlAqtgqo6pWTX7nTRKdAyOGP6Ul4xk0CxFBCJxA8Suh9+4xF7
0BihDQKyMceaRCYjNeL8rDkKlrOdUBeR5oBNuTn+8dXzhIBgjpOqAgNjlXumJ0UW
e7XDBG8Pobl0ZLmqzFS3pAZVCD30lLuZCC0nxHHGkRqGJxRv7eY44dxlC9Ws1r3I
FLXMPY9NHtmsO/rHsIvTxy/Xtjegd2vru4ABMA7No+Cd7ZfbQurZtnwz6QF9IMbf
Z1LyL/TypETI38hjgnTX8+93+ZrJzHPTz1d0lmp+RHhRAMoB1nGcy/5jDUNFG1Ds
2jitNRWjdT73NFjtf8IczKVBVdYlrUH+grojQuQkUiplGJ7oJcqnsv/dAwNfV9d7
9r/fFKJMHX9txYUrDLQB/oewTWNOW+YAzATx+mWE/E9RGl95L/VjmFgxLHab3e5O
CFrkiVdDKS7Y0dkpNO8gVBYH5FNaqz6z2FwbjLXbGeXFkDZOiWMaBlJcpkb9cK/p
G3m+U2+Gzu6P7NPeqhh5569RcUU5YYV46CIWPsoaihh26pPIc6bok0KfvC7bWc7c
KABNNxygf3RVgPbRuZc+oG32b0PnLGoKIti2cXWDS1Q2fTf5eSaX90hep/i5kteX
vI61q60mmSL/zRUzz4+ZX3v4wPiWBf4zg3bQ4O7zx+HqNLbbuZgIb02M4ZQujkwD
E3ulhjicj1uwWrzo1BF7X++M5nmTDlQ9sDWSCfWFEXpcLQGru0M2y9uZbT+dyVUJ
w0fIORUEaBbZfOqOQ0V8/c7/MI+vgtFt0wdq0Iqh4Kds3Ng+TARK2+x+xFjkLXoF
/mF74corTpFUq51RNip74T//VrKNcvYnfsCaHY8/bJNLB+DjnFv4YhTvvbIobtUD
SQ0gk875G6e9e8Mhp2sRpIJOfE0o/5F7CFjOGbgM92SErSrgEno1GTSoNgdV00x7
L9+OVnHhqGXySM2+kFTnw2n55rXwujHlRggi2CjrWoKbp5FyN8pdg46BaMkpgt5e
e6weKWM9skD8ocYH109xIYwngCKHtg33SD4lyRoHRLiQs2e6lL99jpNlUNNDiXnj
HdUCGZDUSnyywdZqMBdsUAmg24kTBZzvH8MWlyVbJMxRhEofUM6QyntWMC70w3mx
EHNR+k6RQ/JpoaKSuDp969h/PujQKINQ0PPWfwDwJ3BW0FKL3OL6SCasiUDkMQQW
VaLFl+f8S2/VG2CfSTuwnYES9/BAv4e9fyHKkaOGWlta9xpuBnmIND3RPFTt/XjM
2UZXHDkwg2oY8l+wzgO6rCu5zFgcRyyn9NUUYyGx6Dmlv15jI6S1SNyeNAe2Pthu
J4qkk5qIPbWmQI+WbzWdI1woSBIJ/FahAJpHDV+WEbeGAT2waLPQm18itPCudESC
RJ3thutkPaCvRb9/Nwa0gr4bb0zC8RaX0bHJoUMvTgTCG/2EgCGc3WpnU3zhacGx
StACyAxguZ5Y1hWXfeTsZ0hcv5jnaATUaEkX+mEYVUCF+uZVG999CjbLMCekeJKR
MmcA/w4/IP4oQXOc1mIKNz1aHh1dZOOAHN0B9/PF6KFRGWaF9fXtv8/DgVfMIpka
Hryut/Kq1u77Kw1jJQ3flctHMkliARD6CsYKAKQG+U3V4P0nsnmrbbDhoFFzJ2Hj
ieltzMKhWJwEfhBzsndCAR+R0h9u7bZ+3+cLDgprC3tzrcCv+a2x8nLV/x4s7nPX
qMhzLAQ7xFTRzejoAhrNAsw2kqCrpDDmVcfzION3QxbIPbq3sRYv4E6FxxpABZM1
+mbcQrJay+6McwUgpXLEKL+lzVMIHH0sxHfruynJ9Mm63KaJq0iwut63An0tXr3h
rIZwoaiL1SyAaDTU0cvKTiCPE3L9i/pZ2D41ktV3ie31bEJXzG6/2laigF1aAkZh
n/m95x7u4vgdCGHSYOReLFpEv5R7dDDPR19FirM0eoiRRkvHD7MlAJ8rPu3fcit2
hEeCaYGa+HKf/T2rzAeTfj85pfGVO7gx3pFszDp7r2Vx3sIHuGvw6/0pZ+Sy8J24
elMLWhPTIH7zSR5VjDnCZ15uar0x7090l1t+zS7C32fgs90p0beIcb+C3fx1s6rL
0ZVQ+GU9I2ybPoEnXkU7Ntg69V/5HzwhldrXHKE+xTxJT6WbmgI7evG3iPj6Ql5G
7n4c4A2DsxklLEq6DQ09qWkTcqC7ovMM4/DR8NsMwZJ86Mhom9viXvgortu/IZV0
ldiQC50mOT6NuyvLQFe3ZIEISCWDhJWlV+0I7GIeY9lYOdt3YTdClsIyvIV7pIFy
lpfh1R3qpO2EEY9BzypBQRm+wpjed9J7Jo5WY10YDL+KtNOrw3HfROnLzh3qtKTh
xRuWA1azcQ4ioaTaQXyMpcxeBX3mq7Tj9IBVKvv5xDEUVIQ8wxdn572CYWYphm5T
ojcNUwQPZwmPg5Hf6DmcvoUrTcI9L6lPRSmVbAO2NZ10gb/T+oOzKhVzNCVlkpDV
lrFAd8dNMI7bTp8N2VJoi2fNR4iLmJu1NHmIf+f2PUPuCFT4uA7KGogj5yQM7bK4
vnOrniF3059/KNQNpVgd7+KS/at2fltVI03lmez1hg7l6iKPs12N/jrP8OnqRr+V
qVPjlvLWDLJQvobmMIPPdALadARD3bdDRkXUpJ/Nb0RDAPwiKVQyWZ4lsD+epKsH
OWgqT7hezuiaHoY6HPRRhFGaQFd9ET388MDiwNWLAZ45jrj9qM+0tk2j5BQIxJch
J4g89Kd6Jlc2FBiUvxP3oGaIM900MhWlMIY6z4SYRqwPhokOu91IvuigjfeyMZHF
rJ0unlTrAzri6cQYcIsBeFPCRFIA8ZJDYSncRL8S2qgIQU2JNlcqin4c+kX0VyvC
LTkCJy5DJZCwu582lKJYD7P5Fqph+fWVMHSrR1QgICnAoTBho4SdD/H0flA/Tt/y
W4GqTtGMI331mmhFG2NR5EqyvVSfzGQu7E1Js8LXp+stGE6eZhuYBsBQ0wUsaP4Q
KFwIpW5CoxjaDHZBpyhcNSKTSpxU0uLH61P/jPEWAcIrmxsv0Zs414EzhOsm+9/O
DqOth/1cYt1YeWUoCVLeN2khWQ9Vv3MKLDDftzpUdrJtil/QpIhNmXWDzWji/hoT
IKrRI6z2rh6R6v7yoxdrkLwAl7Dzd58OGrzw7HVz+o1VIo7iHW1KgmGUNcb1+5MR
M0Jk0GDpQ3yWZxUwtm7MqPuLwBAbr28wjqplP75fLGNFgTO37HhZu0ipOvN2SlBP
4D9UoHYmT4kOhNngaBGoeZ8uZmGYS/VshhkZsuqXjL5MiERhaup6y4L5vj+387zC
bTqgj4saghgE3iN3T2XZU2hhM3n7xutEHHL7waK0Df+MX1yRwXifM5HygOtl1/N5
zYqDdK71P6I5U1ljOqYtK0NPUlK+v/oscpg9aw4Z+vrGeKGiNshN3efuV594tMKM
J2Wfs3eeYBP66dn5YkJcVoHlHMAj8mXx6DI6VnqKJrWa8KdGUmHEJ7HHq86tZCrc
VDFUKym05+nClqP6prrCKtv0q4p92qQAJotJfqKMwml2kJVBm8MEA05WGlhTy1pF
IfWW148VRKKE4CeuqQmdli2q7zYSU7gV0SST0+6cq8B6mGOIMXjh0jUo8tG2SeOW
rmLSy9rKmygj4LcJKn3q1LMXiM98McXlUb3WyKykDbiu4OzQWazQrAsVzAUmJWu0
vFknVrk4RICXABFxaErh6cc0I9pGYt/4GAXtLkq6naEgtJb6HmENl0gmNpCmV4+r
oc3GDefkYU1OQLeMlWdx/MqGl+LZzPqpg5Tt2MCj1K0pE91PXqpn5Ig+eNwVIxLv
O6H3MipjdmkQRWRM02ZLtezjkadbKzuY5LP92FH3Pf4q+Fm6GPkhPtb2jst44rvZ
5UoAV5BlqlbEaG8CjxzdmPOaNDjmQFJfiDlAV0xnj79NFAAGaP5tv+ASSQEf8Sl5
ljjg6KXVvwKiWyM/1Yl246PwdBxSmeMV++G/kuk5uEt87GSBVoTHxHUz1lMXgfZV
MoinpF3/XHvu7zg0zUiLWR/4xsQ/PLCGsvQe5PKxg5FWbENnbKY97co4W2p5lo93
E7ktgdlTOTBiRtSmmvzxzU7aV7LaHVa9cspzicMiz+I/y+bJ/f1eLbhXjDjzbdKT
c5epCmpGc6f3yuNhuUydLhKtxKm4scrsisvSugWLwqxXc1pTIwjGImlrUnnTiFQk
IU0xbUl82CtxShyR3PENcntxLgkQN26JOsMZzlwZhIytl1jz4N80Fyg/s7JNLyEM
DXKOVe+E4t+Jo43J5LX26b47h15vDkZ5762SUYDzlwjI7qj9ZKrLW4U8rc81X4sk
O4vwB3M2d34St01Zzo5YLedD+Tiis3OpmI1VyEp3bGDugPwdP3s9VnFNYY//OYBz
OyA688Bfo3IjfYKY8ga3Z4Dac2PoGhlSH9+0uHtz/H0z3l4ZOIMVYaIIoLrWAE+I
Age6EksVbBT7DKNNC8rzHQNQBoMH0VL7vX9S67Q5ZZmHvUcGBFxXJ/rPSPR/vGVo
+k/KqKaVOq11k4s2qZEngzvn7+9roANNNg+U296u1WK9Kk4523zx4BIXm2kbX5mH
BGLbCJT78xzZO7AoOTpSeZ4QNWs4Gcv34sKLQ4qXHgAgtp9Wwl0YXpS7PSmpWZzb
zTU5Xt2xlIeZw0t8dGoUboFQcU1gRDNz3TdsCxPvzGR3OiAjtMWLAfb2KxDk1T7w
I3QSeYO/93TSzjRLc/fsklHm7KkabRfvagUvyiYmU8Q4xQIRQDkEt7Dcs9qsrYmn
xrGoyPqRSHhJaYpnVguR2PlDOr0Gawjq796eDRtWByZT6ESqwWd3RTF64BPvPgV+
Y1eZVntLLpg9pR5vZq/FehK0Tv4jwT66Ys7mOgXoNi6y6IYHyPaGnVWJzqvzOEON
/b4ylXX486mrxBnDyaOFeAd12Ic4hNq6TbFAoQAmRn/HgIXcPc8c6PcZIeWC4Q6n
tCkzOZyXpMfJfB+hPfKRIHRZkBKXQSg1ZnhfJzT5wunh66foEx1Q9zHPDsgklftT
BpFJm4M9WB2lDfvBt6AhNjsiRc9/CU0BTAQ4XxPcMi2Fp9NG1FzP1aRJLjAHWuQE
iE1d4h+O8a9kj7RJ0gwZ5AdlnjUIqv8PN20X9xToCyqSdLtaCVIwDEbO8GW2gdUX
oYz3m4S/lDt36iKcSkzcjl2b0pVkr3HxxphwWowzuqardCX8ijTbOExSpBlNR4uV
xAknXEeiZQbjqVo6Fni6Z1DgtuUSoSXxylYUSKWD1xUlW3B8LIa6ZL+VKRLVpA32
kMXgCczpxoNRYpHp6VUzycE4+gR6PFsiYZtJ46t1l3VU9zXjUST2oQQtNOVEYd+C
RuToS82Tv5YgWqmYLhqphIbJY1wpbHahSEm3vfM042l3Cz1CmdQ39T8/+qxrxRJM
NG3dIvfuPzlV/aiy4XtidWfQ517PQhJtP2OKfeG/M8L2tzv6d/GEaajCiWHQQxUs
ahX9gGv+pqD7FUnlaOymmUrgyw7V/a6cUtMBP6WTEILk3sdkm/iTrJyzToHgl0Wz
7hvG1Mrvl2JAF7V23Vct84U9FXjSyNz3HaWuChfhGlqs6/lqWOP5UrO7FhFRqa1J
PYb5NQCCcK+wF6brHXHyl5PqC3QcYf28WInA5B5CX5e8/2McEBlUDMFmRk9Ni3rR
QuMDg5/aB9QyNScQxvllOAUGy4OCsjPUsDdeX0Cy4L9VHjRqVeMU/vt5wJMGOF3Y
Oo3pQaluoLTHDYmJyHYkFqEvCJOeSiCbT49+aiMM1dmy68NWwlcOFvfZAs2u5oYh
qTfQ0DLZhOe/d/kqMGtAPTvKa3xeXeudtkE7L+RgV0bAX8hA2CiR4mj/cSKDAwUq
80RBEuzEmmzUQZAhJodFNIP33ncwRKjZB4O4uMYtoUXjbJoQJwbwRwmXndIYBz78
BtTb4viweczi9fVQGpnF/P/ZUUU3/zzw1yjaQv87h+NX7vv06DTC4furHtqYUJCb
Lv5OTOb77AiQWrio+jmn5G85z+aFk4GFWCOad0ziXN1XNYJSPUH+9bA9EqfNlu/p
NRWnj/pMmaQoz/V4PLO+ZgNUd7UWEHyOIPnvaAGA/6WEbxaaW7TEFUh4eC2jQSOM
ZO+b9CD+2YWyRj4LRNzKVmDMFTJMT/gMy+VpqyYXQOvR+Q9eW3EIXMjSJbH5yxGs
T3iNYg7w6J0rjhRTJc3vCA8JhaDuYhR503BkvatZ1Y0bm9Gq2g4oJqHumkWMPhVp
lBh+Mf3f1ibCuVacn5R6ic/+rARBVZIXUm4TC37e1y8CtCYqVNyD5pTPziq/27CE
AD28HEab7Irq3WsFPCp82T4Cm4hsD8z6xcTVBItNPNNPXzI39CFKsOhB3ygcW6yo
BzmK807deMTYLem2dxHW5psQTlbvPmbUOakagnFkblPtih2cvFDr/bfnI87YkPZa
gnvYxc/e4U8YLwXIHPd26kzSOaePe1Vmrc4pmLm1lK2bRbduo0/TpQY+MNY5NrJb
6C9ZvXTcEjYOKyBjE641hPSZj3Ym7WLR6T6sXksjDcPk4jyvmp7XXwo/B1x5hsF6
a7KgaqpnVmp3JEr54XmKafxvg/ldfLT+2FIS7ae1LWGmXt98DffjQzhkzsjsUttV
OBZWreqzroETNO6gig2+8mgx68Iu70nvfnIOWTW60RAOrU+T4GO0OUUIKAZ06/4Z
YWMkzAz3UlVxmBajHiMs8w+6XysiJJi47jVsbA5xW9B1QHMQtywitZ2FNM5Xox1z
5yssjwb6jcpUb4C1yNRYggjI2P3W8sX45GUY+tT0OSCNNxNqWvNcF0K/N3UXyKUH
4nC6EyGJ7il/uyZcTVOCC7PEwVpghI2w1BjU1+R5HnltZ0stFbNY2LpfRA8ooJLB
neYv4LzkaDVlw/bdr0OFk4MM7expuMU/0x/IbeMvi0VgxNRBDjAtXFNNRt5EV8IN
7nGkWx6vwfuS37ZPb5RJ0GMz3XejTwrt6sbbwKd70ONVKFyaNkmyw+feQYStOioy
yf8DLz7DrN89CawAyh+VSVJKBP4uTaH9j3PNSI0LIcL/Nw48DKyvgWLK19LBF/pQ
Vj/wOIjGe6izhEfs551+lRt2Iys1KD7rHUymDgPJQ5opnTj6sCVVfxdqFngxHOBq
CVgIEH0rzFUkjJWS9wl0mmTkvDtCI4KLvtS4TPTKFv/ju3qJVrx4xiQVaeGtFsN2
8oLV/LLO8KInqe0Ace3fN0wLulKVNX/5M/MHzXqiv3yW0q4ePdxdgSSaxAu6wmU4
GWRjAZh3vMdgUV7JtM1swGU68dkWCnohTdt3iYpolr4NRhPWpRUfohKOIr125lIR
NOAlU2qQ3JFgIZb3EEw1hNRA75kzwQxALUFEfcmWNT/mn1l8PQUTPSLmGfMMuirc
QFyS8p56D/+0HwB/xyYG2lJ6T7bf57/ZU1YD2u+XugrzQYiNGd7jb710AHI87p+8
eBu1/go/ci/yxlD/tzfcy3Vbn2xMQoSVsSyZl5amU59hXKW1w+sOLrCzNgoNIFp2
84GBxd1Isw0gRb82P/byhg8aEzzgDRhBynXnq/Z9L6RgFymwOcCYwQ4buVYnNrx1
dv/dZQgTar2E3ts0ym89frsfVo4fjJiauixWN670GTK4Ref12hxbQfN3gm2l0lTC
XfL0OLCxMfLvKihLT0yN79w0/SGVc2nDpZFhPTKrMZEabxD1AtX7t2J3c2W7lK3c
EBMkTGhvzsUvgDjPc1NeTAQvFe6aESQXe6HwRnPu2YZ41mOrNNIn/3STuI9cT/84
El0zM8fBJP6kA3vliKXAdrnDLVKR3r6W7Gntf62QcISjHWEz869Cr6TxFSR6BJvG
zBlihcFooVlTlV4PZYMt6R6NS3f+N4F2vCTUg9RzKElNVMI7w/lej5l4aHdkbzoN
zTyDxhCSoCOtId7iJ7mkIOGPG1vWtwcoHCtgIZVbA+FZNVQtfohn+9S1/I1PRM2S
GNzi4B2Pfqy/4IKtJGIIppK3FfkYdD6NMgbp8OlUnePunGZZ7a+/w1nynBGmSUhf
Xo8rLXFNuTAamzwJSfYdqX8M95QjyGaXIMvXvLJSYCKM4pxnmf5Zi/k14AhOE6Hw
UX4oREYtmP9WvbawYvZm0NiMcUxl8bLnXVUMF+G3wQDnT340XLg9SBUExYiNzVtM
c4kZRVeqBduTtvGYJX0D/1uAiqScXbuvPdMcWq98MzRIfFjIEtRbzs+VP+wNglnw
6ql1oQ5aXVG6Rk7lmG3AX2vhsyajTvwsRtJcd6pdokpgJ8AHczL7+Jz0re8wo8Yk
appNoE2BcLPLmKzDHfrjlaKyP+qEX7ns8KicGa6aQ0pjm+T3BhWPf05SRlQ1J2E7
rQyR8VnbEXiz4lOltbtgs8sk7oISzjBwCjkw9sWCfJ9nv8jxc1kgkkqbrkB7QvGj
a7zVhPI4/rc0JJBsanBe7noKC+dw/COZjN6hjTDsqaZpxWwTK3jnVKOqntP/cOvd
BkXapvgkbcMEMwtxrD3chF/w0ogR2S18eTcUeGuZwYaMkAs38NwTpXOAq8XjYBJe
4cBd+Nubyv3FAK8w+QtpGWH/3oTYWZvYW47a0jM8JBWauchkg9z1OsM5cuJpxBz3
leQBc1Onp51nlAHPZAhWZxlUH+idZrz+zXXBOPlVIkjYBv9dL0aOQl78h1GX+tVy
wWee/h/HfepUWTQRfRdxNOXYupEN46vlBuPobTbKfu3iwGFs+iL49V5NStt/1WG3
ae6ANjIenDoD5TwUmXC4IvxgAKPQcG7unveV8ixdmuJ3zvhmMxTHGMB2UQScmr+v
g2Qh6LjAGVTFNiDPXljcVL6odxHb43UJ1UqhMmLRSrEHrzaKQ/hrOTWEedNyB/KY
HsNKSpHzDXB0T+jnRYTKmoQ0HjTFqBw1Wa4sDubeFEv2tEWYkckYMuA4cjoi+1Lt
6llJQeAI6FHygK8z/g/uLirVLbLc58K+OfhbqlY9//ygZXC09kq3fLsEstF9UZOH
cThlNMtm081Wd+twbLMJM5EylUI+lCkqSxKu0DJwAlASZKSSbg1Ei2Yo4E9bOGPv
WN4OQTtjd78ZeCyJFHz+dS0DZzUpJtv6u3B3F951zrRugulCP3OKPPoVKJfDCZLR
Hkjduo7PXQeRh83WH+ifEMitIqvm/+yZtc2UtTV9gDwQlcn6Wu+iQS6rzDWaYy4s
gjNkZhwSYWgDa0UxuTQOis//iPulKiY01zWj215zZ3gqk1zLU+yewN6aLv/yIJrI
4CcPehNhRk6e1IyZQ5ZMOp9w051TRByHLnG3YGo/3Cl+atP0Xm2BdPHhPCH4L0M8
iqgGrDK+e+LRxf1PDcH5oyevcKq8KjV9yO8d83FDefIYR0e87hj8SRUjQXq+Kusq
FuqM/FKMfa3GHMSVoD8jNur0ZFQ0INWzS8+AftTRQzD8KrXoHKFMtBPTT6nIh1ms
yzyLssNnKkKTfbqDQ3PFZdYcTvxInNlk+u//G0J0igZ1wKVNzfFra/+3mbAOdsww
/tqkTFeXAlgGFEbtm1W2pw0+RAqfCOCqbWbRld4TjDKbYeaI6m8kGx1qkrvFawGT
RYGeVxbJqSHzCjH9A1/6SsNqyMnzw6eXbufWqEVVSCguhIIurR8oemmKSsxj4hN2
2iYf5EbBarFRhRjmqZF9sRXkxoE5V29xQUHnWKC9JpPejgHsDlEazf6tmzqkkSeY
MVfSdN5NsukxtO6t85hCRiKwvY6GerNOSNqnT+A/UUXZHR1rjB4CDwi1pr7hLMWN
aCSnQ20nm1pUm6LcsjX149mvKNTivuVcfUot0DtvfjX7JfEoLqBu2tWVrBwlijJy
OMYIPvAEL+7j0TMjcSmva0PRK5T863kLAafJ1DzbNAWc3NvVC99YO2DSaH++71Lv
rrxVxjeAcv9iM9TCufDZZmCibbkIaEm/6RnKmjAMdltHa8b/bBB+Y1gzzxI3Nvux
lIZEngJaQ4GPUDdSgTaQtxlgPxK2+bQta9v9AaeYKwoaxxEvWA9kqVAoVXgfH9SM
ryfU8IY9IWHovo5zU/adilviRjEv8wXNbcCvEqsVXColKHhEizhNqCsFmVo/PhV3
WOuXsopkkttpwZrleIVVSpkhqob3Jj/xLKQwdFRXg74yMtHARRjLkNudIZGcesGw
1v6H14TFNSQwHo2optbsOz31lT9qzgSY87ylaz84w3iQTg4Bo2sTZSX8A3SJHyn8
92wmmBgZA3M1nBhaBWBMPtE/W7+VvOC6MJjazCjDP8jTkXhVYwW/Cmps8SIoIaDK
XyW6qbJUCt0sRIRmWp22YYLIAA1RQA05BzdI40VHhQt5ql0znq3pY/siXHcGz7YR
cpjdTVyYVWvnuiH+NES3S/U3RI2t0S66KRp3WnYniHdeCjALAiVMaDx/ES8jjStd
rbwrIBCzD104IPQYU+f1Wui6k0f3CbwSQ00AyQ677BxN6fU3wpDZwQo8b9B4GEvs
MY+gLZVHiAhxpvuFgDZ+JSDG4zF2lUcPvXOKkUdlJLiM2EVAkXdR1+2i9uoymPUW
PgHl5yQUePLRbDql85wqjAuVgu/0nB/l7Os9zMpnegHS+JBmbPDZNpG6JB2qijhQ
hn9fUbEFc1uXizBZBAWokbDTCNAn/T6KIL281JtAtdWynxAKSMdj4EQeDU25Fq7d
tj0ZginYXwgbDbkrbkzx3RkBZX7KSyEVmb2ZwtVD7zFiFnAk5G/zG7ol4eb3keEC
TfF+s2EgmfVqz+j9MFxFUv9BLuUYocb8YoGwSX0ay5E4ZDw/ySXeRHDI5g0cgsEI
ZJ/mjiL3MMKfs6BmifAAiZT80cr38JjS7ZGDEdX151Hvap+zuFjn4AmSVMUXjmy1
CUhdxL2rbi70qEjts45zKQL/4Cj8ESJkm4a89/Ee/WTacbUqtFwi+s2vPnj6nEyz
hMgukG9akdNv4LR3bK8ve2O0eSX2Va4oTYKGyTIn/cV4F8ZGI+823quB2aUDFDKO
8Y6RJBhxXxJOAlzvXKuumQxpfn6EIbBcE+uLgh1xFMR3Bg/45Ff353VbnqAOLfnV
2UwT7pALvDVqpVE8jp/drhZtkwR8sCPEl83Y4Zm7YyQYrDySqhI7ovjju7crQ9ZV
pU6Pm2lfQMDPYvX4a5QJHpmOpHOlk8eDIxQWGZ6BYQhmA8uvOqX/5QnGQ9MT1NWt
1Ds/midIVjHOVCaNJzD772f8wDJfAHO6yNKdWDhzPuQk3ZN0Raf/DMghfzzIIBWd
9dx/Yvx2FTE4I9s4AodNbRT4+2HhH5b2y8X3RaAYN2kMeoedZNWo6zJdvGmFjpCj
S5QaR9fQOt40o2dzXogLn67vtIdlfdzuGbPtwV0Ev14nHONxMPydNdlXV/y9ROJg
/17gBWIvzmGtXBrw9Qjqr0JrnBMtPcA+2Vyb2YaXsoaf1LFQaFmSb+p3RmKwZYEa
rvwUcPZFCOUEYbmhqemUDh3niVb6suZmP659IDDAEFqQSQXtGeduwvuNhGs62b1q
9gFzTfnm0Vn11eY8IcW9t0V16eNfnR6I90F7mA/ipWCMVAO9LSzrapsDqtLSr7FM
VpPVr2s9Du2KGnMs9eZNRKwB1gql66+NuavieJ/a2TIGyaMkYsW1FEH3fQT7enia
sh3C3sZ48VDDU3L/7aQDkId1lxym/9t1RjoIOINQG8rD1R51+h10yTj1x4ktK1HX
stkIJ+neULjmKI3+vhVhVQcGPEE41sz+h1xDNMvVjbxQsNUuO1KvU0W/LuTxtJFm
81zJYInKnG1wRBj1+FsbXDFyBhasSNY8ox3+MKkrXSxfXUp9LV6mZaebSDECLZlw
qGqveWpPjwRf+imtnLDqtHhFomqaGiv+mJuVss2yd+1C3ADwW27LV6tMROAxHrQW
RDl8rFg5UXbPfLA6PKXiJJPKZxLci7ESfG13SEeJo3pF9g45hXNZhMNcJm4JVlxO
Rr1PvhK+rkgob3ETCzgTlAImIWlGPuuUzZYwOPyr0f/4G8DDstsBvedw03S3sfwT
1pdR7cMjLv57jo4TVF6djHM2S7jOVONyd1pMqjtcbixBc2eiCEr0KcTr/ZqRBrHJ
JdZDxwCQgNzlR2sjnGq4tZ6HzUiz3EbtXzY6fp4crUWG0y+nRcM5VJdGyDW48QBV
mEIilDFbUPdbwl787eNZmOl4WXcVyot5/b7MkWzDGzhxtXlaq8W18P1C0tIanmKM
HWQWg34olRdT7qA7jvn1pV9Do5HZem1L9r6l8guL5IB1pj1PDHu1sBZuxf/wmEJt
iFmrmlzCy6qBo/RaJa8ObrD9Vory8ND+LdMUWcGgEIpo3iIVgp6ZIARBfGyyGzrG
mgVosUjkPJU4F8JuB5Di/KMzpccZhE2NutnoYkZ3Vqez68naxqxMpKfpjwftiUie
krszwENbS5hRH4lH8G+VPPBbPkIqYkBlxHXXKX2GurEx0mQ9lJCj5687OiH9qXm0
aFnANdj9xZaofq09C+urtIoAK8HCgEDqVlASolzNYqHkwH5Sh0AICYFso58UPbLA
DmHaMSS8UbfO4LT075g45EtqC7BeTREn9SA2gWN6KFNeswMMql7y+KdKZc8XnwVr
B8VddD9iMlIML2YB47xFNgeLWMhGBdx+5tIMRHFG0b/E9WYiPt00dMwXfGubCSid
Ukw2SP9N5daYI0BrPWHwlNOhVdEZXAwyTuIW71ulsiWH1UQ8QGPQuq4yoZV7fgzy
/qZXQwTbYu4w954SHWOdfvqBs/zOWLXw/FfDZj7xSNyZLy9EpipjesTVXo78/jmT
aPrLCq3ic0XDJE0Jz0VgcoppkifnJkPgXS1KIlWLjEZTh7I1YngmCmq6bGhocjk8
hrgfgmDfXApSon86b2NqWUIqlLdbp3Y7sbiPN7WD3e9BPZ+Djupc4QXytKwqN6YK
LsXZjoH1RpsFUwoxyM4nd1ySFEWZfAqKYfac9Qj03kgY2fZ6+usLoVyQ0aKqqjpy
4Woa5vwZ69MMEHXHNMHoSDbz+rv1XfsBICf0aPCl0O51hgycGKl2eEGPyKxCPfZ1
u/wlHo1s3y8uOkXFJZweS2z/lbED3D4bCW9ARh1548z3TZ3fjmTRVrtrTxOl8l/7
0tcodVx0ib6y/TOuLgCeIJOdFAEMK6o0/zUdhOheEzgpUAzAAuw+N81BaVmskFUX
AzSR8OV021Si2rJU3E1XSnWk+VjMTXcanNekca1x9SNQAiHLA6whTRtQnJwwM9xg
22wH+DSDBHEODghXyLcS0fCNK87UZq2qVKGG3/lbkhaTaHzPMeDrrCq66Wy5cy4c
njCb1MB5Owllf+IY6mMv4CjX4DlSZQtVp4bTAVV2+LpTmxNP8MzdtllIonl2AowR
wEysPFUR+DhGhPXEjHpeXYCPV2Or91/CC1E/XZ+YbdBeULe5tjr9wkTkQZWK7L/d
k5rX9D//NtM/ixMj16mc9JtNYZcYNOe/XJ8M0VCiDdv3p6D6flcSkAXhmEhInz/U
zxytvGk1sq9PLeOkDwaQ8IkMJp0lHX53fH3RCJ4Dd5dcvxUXT+Q8JkD9N436kXtH
M0uKMohx2D4a6gk0cxbu1QOIpDJ3kNCGNzcdHQrzKNOfKKIMU1T++W8N8jXBsQhW
6tTsb6t62WPQ18hsg8zTr8WhcfJ1Ql4a9Y6OK8ow2Tuy6tZ3KPPcsywh6WsugLmK
astJyTf+q/tu/NuTcAQ5wy1m3agDLSAkTIZIn5eljyQtdvQcKqP+NVaSS5cx1zqx
cCvUAnCQDxKzcdkC7cwjkQro+Fu//nNCiiKpd6PCNObvHX8Vg1biddGhNuFOFjRo
8s5SbDpuJC5Cz5dmfQ7d9f/EsKP9e6WidOW6UdxfTTTcV9t+dPrXdhle8a3uOHnG
PIcC1Ik8yxqkiCThfFZiW74fqc6gHJehU9colhORIk8GK04aSfIp//NyUjEdBjF7
4tLPe8i5f7BStBHzKY4yIDPqJJLi1MRIQ9+7YAb2oD8liVDzGM1lEr50z601WkUD
C76IG4obzuChnZyjsPRqs/BNOF70zh3Lyw049RkDqWcKIHvzbDLZVcZYZv/NY1xw
LgTNub7dAb9xXGpSm1R45c8coXODJir3zwwHZyTY792fqNFaMS13eyMBPvHO74DL
N/NUnjf1FDqZR8qc1iVx6mjwCMB56eLgy54MQTelD7yCQSQha8RMliOVgcDi6tac
vsswclm41vhtvgDq+QU41t00itsf9iuMPGocOOBmbJAtIl4WvAGrsdqu52L6wcBc
VR8qMP3EZRjHyU6o+fzS3L08uok4Ry0eKVdzKtTMffEqyv2e5xXOG3F7Gy3wMhr1
oaVajKyP1n1dbsCz9As493z/1Olgl+aw6z7Ui69QZRoNdkPrtjoQ7hmdASLo2Dst
4/GOLcd4GZxmmQ2U3kIbpa1XUi/hkgXqyzQ92FPhT3J1a8g7GYGvbMZlElc4yU3f
ldX3QbyUSLhsnT0O/l/0Of44gK6pohASpBb0//DX0WR3GW8SucYlYrdHDWDqinur
lJ8HoUs1/VixHPklRvlMdMRiF0Rm1gV0BBBTytBysd3zgjLl9EDcBss8vHdWxOGG
dxsH2CoCFm1WicdYAQ7SGH3MiacSbN2Und4EWbL/G2b9Ji11RbdR72mTaZ4hpkmH
O/EW2VANge1C5wkajTMtg6ng9xt3aR/BmDrBwfsvOGxo8ZrA6CDOml+jwYLmr0WF
5TTdcvUVM4tnQDr/d6uxiPcYO6jpNwj//SLr8ul7UZLshx7ok6uTfBxAPKOzU8pi
8vCeL7SfBf7hXYWGXpFxTw0R8VeymKtYzcqOHPAR3n8/R9rqYV7eqAJhupp1+bTG
sMeHNMsdeGqDjAo21neTnDWqiKy2161+xV/1QtS7amDYa0ctVsw2ZNYG8efriphK
MJCsRAkQIx9XA4pZdv5oBYW73J6sMgXR2Znbnf7uwHFbf2lzWikfnPdw+QK3N4KN
uevIEpvh2pATtbTfe1XOlzFgu3PGXkCsQKnM7ZG78hYwpZj22Q3QGrdycYGIpM0z
fbGAHkNT9RbIK9DkGre1PO4Dast/JMQS70ZfS/l/GHPLOh5CtRaFIzVI98lQHV1m
8UxB81oMFDXf8tcFXCHSWc7HqxTqX4AakxQ+3bNO14422eZBHae6rrTSYAxmtUyE
TM0ATHeQS0wVD1TQQhFsSY6uJznpC+IpKbc+uF0cSRq1DJS3Y5Ql1wRO1prHsAf7
Ntcug7g9REOpl1Cc8XyWNJuq7r7T/EyoHEVbi/uwiV/uJFYjwiDQmlozCGSCIH8b
KamOW0adchQf4YJb2aHjWHp22M4DDnvf5qqUI0DNAZL7gnMehFCPxWvoR6LH7+0S
I6PqqQwZ+MUHA4DWw2pYJ80w8E6/itKoWQIw6gJ1bscEZ5TON0UtAey9DKGnDwt3
1q3Yu4E5Of6vS1zFoLaB1dWFQf/nbo5SrchGTDA5OpwvQhPxEE3bfbkFbjgclOzD
m9loFVxf1yneV4KpJB1E4QJD45S3fYFGLdl0C4r4XBbZpiwII2bojj+NIFi7TqLR
FtwT5ReLiTho1rYBBMNZwrIoVTM/PVPznn0xixrAVaOnfxS3DGM73ysdxpA+LSt/
MaT5mo5sB4hzC/NLUNzs5TFl/nuXcqPNxEULRmuM7k/+r6+ifzeFeugFjEfWqXTK
FfvXtYbc+OQD/9yuiBibV20GTG2Cs/U9YrO7KSxgIwzjulq6HdlZLtR8vvVEr5hT
Np3Vi5WYk7qHGyiZ3ReOUCOU0Nk6JLJQ55fec0U2RBW/szNYBiom6ZoFGXnloEjt
AOZfLxIUQZ+b7TqL8him6SnzovovNjLtH5NNvciXOF1apW71s9QBedsQYIeng1iN
R28Umk8i3ChyJYcUhIcxCErhrOs2q9KBBSqYvalUAAV+1BcVCEXQ+LHYWNHb12zD
FDfcTHvQTZ/13WiVEGjyxqxSMJALawDiDpeG+jyz0TwLLdLfXSv+qsb0R6+Jn/kN
tjS7Z9NW44OK48NJlP7YstOrQjPjy5rGh3JMbxJGAf0yXL/x+5hY73RHiTqq6g3P
ZMmNm56/RnMcx3OyGnCg/oJqvsK9LgQEYS3dXCZ1OXjK3LjKMadxKwFesee7PAVR
7gq/GeX1HbJ5AszRXLenHCury5grutDeGQZKs+X7HAk08iOjrsjlIJh1MGrIrWHE
uZkdN5BTKlpIurEDIrdfURDcHPkCZDgmRKmg5sxHhT7XZOUVHK4a5wjXkJeCva9e
J96TtLgy/+JICGbGOvVVZRxZA+PRortJp1vyhO1Wn2N2MQPJugEb9EAcOL0KJsyT
/n276vkkIc51CoaN9l16ygTEMOhlBLokG4bYFB/bwIkPun58R7kRxCIfh75A605G
i0fTYQ5Wiz+DM+KSQiLOVEfLpjomrE2ZVSnyc4evaC2OVbOa3w0euMjTrY8KvmJe
SN0lzk8ib+ed1uSQfGRmq4ZQPs99dcJJw6MOryIUQl0cD5aRiCyPm7r3I0NnlJQk
egdFEc7CAUzwoyYVowl2oa58KtBt68gRCkhqSfhDQnH3Dt1n+QxKluzoGQfLSk7d
XHZdcK4hiU1YeE/mPSUs87qyOMvamTTFfPBXAMs9eL3ZCnnh+9oMiM2vgDD5Ri47
+IVIrnyU56PcmKmuGqZePKi8cDM0ly/wFpFKbAbbhfKdmwJqnWKq2cSGrbzvEC4R
7TRxfD6HTrFvXgSxhJULRYh8ZS5jeJyCWMS3N9O0TiZxVvFY/8un7Eqe2ikbt94g
cxe0ZpdkUYm912hnEdnxIG2hPFmxiGjH8LYfoDnLvFwnKxMs9YdHcMgpmlfah+Yy
J6kF7yQSvDEnz4QDIezqEl/ZfxWoR0OGTs3b1BX9ZzJxnJ1tGI9Jxkn/wFmWOyHi
moZkV33q5nxvgP4fXd3VIK1l9p4kWvyWX/f8Kdt+F8B/wrYUSZmf2GRIEa9mGUj1
WfKiZRjhtMuLoREVSXbWkcq0R6CdqnSu7SfURmqy9D2msIGeVuAo6A7uuOUszhk2
Ywp3hBCg5Je/ny0sqKFo1SigQHoLdyxHF/mvDqYN/Xt9GYPacEJYjYd1WikPtK8t
fP+q3I+OGlbGWoyNQexQ9zMdfnVX36Qgb7POYQJbsKohYBtC/Mv0L6ZFmrbpe18L
9kinVTQu//rKGbV+ndqLnkMDm9Gumxv+2AyjYaXY8QWQ3/YHspanNBD2ueDgRAHN
/f85yWrh1rtxT99RfIxYYRazc01Gs749wCR23mC9AxSJ3vRvFKgekSG/wIiLAcaA
3Bz8FfxSgI+Bj5dovTR7uTK1ONNwHyQRA0sIykNmZl2xobprtjjEnARJkolXbhFm
UYAUjQfslvAyDhuFUdrmDLSgpR0h6Yp8Mhn6ODiTNM9LWjWoO9clQ4mJsLZoRbsp
cj06jGdU6GbCdCw4q7rBLrdmzq80yBX/sDWzMO03rdhjHamHLkgwuqKOFNbiocpe
crxqmuAd7NKvnl2RrSEkyYEI+79bN21QvJ9QpYvg9962XEINEuE+Rhcz1DAPt2YR
+XYHszMrrW3yaNKR9U39CvOyhCPkysSg/u5wnZBWHIkC2K9YL42efyJkGfGV3Pps
ng2J6sO00vHUG3w7ZebZkgCK9pMT0hMVAdWJAywx/htl2lxtUWY8PT3M1eUrRjOs
4SntG5pLcnv3KUt3+OdYhguYf+o/vd+4V1ZKuq6D5MnDtk3TzWGMQqsttbD8bouW
n0jWLpFBUYVtkJHMYgy8FnrAGasPHDALuep0ivQCC5Wh8QX9QqfUbMPZHCYCRFyo
/2UQc+n6S4lLdER8cEFDDRojydiH7wuwJJyXUtlKJsQMFq9aDXO8SATxoqH63I9m
K5cgLkvq9qSifrKk6NYMTSGvf4UpzZeTnZ9ifk5HCEmyXvYXa6cIkheNNzQ6Uvg9
Zerz7V9ayWnohBm9yqXxziv0xGUxDNjgo9g0zaezy9eB+Y/xiYxMljlrx60j4dMp
U6iU7w7Sh1+VQNgq4VInJ0lTZxH2IJY1JzR66axQIHp3wkfkXiNlGyhsTHTB0CKR
iDpBSBwj/rOoxxe+Lr7cgGxsn9rjZema+gQCRLw7etNbW6dye6SLMIdJ79uMu3ua
nTbKmKIFWn0UY7VrkVTnX3tONsQ8cqQCkfqn6N6pzQioHBtM1PYIFMknQSp6/xKu
aojDB5KwMkEJw5Q9GFCUMwW4lIp3dOET+wfNYtASZSjdPoVkE7gdMh4fJgo59zJ5
A2uNkMWUgKkhTCiy0lgzsMr/rof+4RFJQSY1FwiqDKnd4ESNDk3426MiaJgVE/BI
yhRUJjacOox0nx3KEgt9NMnAZT4vjbsISGPnQGyI+FFgQOgwEkkpXoaC/IY92AD6
fm+DXRh16UG/InbAPSaXs3vqVCC0HgT5e78P412F2xYMp3bX47BGv/K6Sr0ojgnT
517VDDu2IOYAmvj8SK/6ICJmXpxukxCaViu1Vc96VCX015RV3ZvudOjyDFSXhon0
WAxGwuHcynRtQvv6DYfVHGQ7Mu1uYRkQdxB6vcEEYCb3kaWdqogR6Dn3HlQCdV0s
QEt7xXpt00YXfaUq+SeUp0auk/YU2+Nj/bMURU3qLIlxs3jBQU8DSqLmEIIe+BI/
pZHW5b0ZequxiZL/kdoWXowQMXt018d/SMkQ66NKbHKLQNUcePi1M5kwnYU6Pdc1
2WwVwFbg8kZQzWbDVxB+m23PSA7hnTtuM8A6wV4KBFZRrIsIftU6RUHQNkQ5h1MU
B/Hu8qOCMkJ+z4B3LnoJiGNaglomhYaqA+RrOKWqzYIN0f4wQ8qk9+006jHAHrkU
TBTmsXaqIzbe8M763G5uZi6AQSVvZFcFTmCPpAzqHdoEkt/GVcTfLBG5aT4egyzm
+ZxYNkzgHqb4uArs8PKwGN6SCDVwHUiE5O5jut9CTYA3IhgXuChE0+wOoX8blGCb
FbxMmxXXCPGUlrJq4FxASqA6o5kHiQjTBy/qOneScHF6wHjTkBOROL6jILiveUMW
PKt3BJ2MysNCcpyfqyjDy3h4Z7WBxzCTvTqLnLEepM/xApSKq6eZVqarVsoakwhc
ic3XxWJsrT+OwhqMb0PB+xiWtK98cbbX3qWH/K9JqSAiLzta+pRiLJ9fq9sD9yjg
t4VQmF4a9fp1BgInSAzAyQvgtH6A/BLvcyGbO3M+j4PTmCrV17fVyzI6F8YJvvRL
69oIZKvjgaZ9QiXwBwrAP8kRJz6Fk3cuqKHHtExfrxQ9jvMDrkW8BlGQabnz9qcT
NrnGQq3YMfY7yPsVazeiWfsemdV55EUCp9Zl3iYXqnGzjFg8Evuw2tMDlx6uQ+so
76GAdBq8BaMjckxXzIJEJZXbcT9P8gpcsuyybVutm3Bl7Rs1bEZAQWVkI2vXY5V8
2LEMHjzU8ozECxeBtjFbwmPK4hD7NvqKMapHAdWFbVhfetVxDSurWM83Jy/S2yjj
niEiqoe/aqK/nxoTNaJAAr5K9cOOrCoG+HrQP0aWs/lFeSEFAZutPK+o2pw948IW
o6WuBmM+xJozhDTm4qlvalj/LDy7UxWLKLRquX2qvw3RFvY3IqwnCHuwBsNltvPV
TCW07d7UrfMAFWT1UVXd/qmWsKvn33y4lJDM9ExrZmQZrMebgAzoE4M/5o8KYFns
9lJzfl/AA56v2agXq8p7YZ9QagUiEnrOWRMGOPa0wolaKMC77pIGRllRqLSG9lCW
usysT6qzCDt1p7Atm5N8Ql+s6oUDsD+9C+5Praoonla1JgPX7J0ei1OWC5w/enMS
06QuoJu4uXwi3FocrnBWiEHuB7cmRIsmEZfGjW4PKSm0D1Kd5FtKSYllyiFks1AE
U9jIhoEzIzUJ40S99Jae9Ke3+25E9aSGBJuuoaUaxZGsnIU6h7TgIk/NdFGwfYvF
jAGaiNPO0TbxRxI1gD1z0ldQhQeRp4+Y7hglWXV0YdOpQ0o87FspKxYkYEIMMq5/
WRYrFwp3rOVO3/IVeqlywk3vfJZ6ZbTt32FcVMY6L5BZ+Hvziw0yJdgnCT+/ayc/
qtnaiBpWRfTosRq9rXJ5lNSlJ7kRzAUkTRZp0Cz9fBgO8NwvxYVQHtH+rVaRD7tp
MN+o2V0sn3UHP0tHyaOqeJ2cVaDqRSVM50k68bpjm6TPujpbT9oeGW2TZGVRP1gs
YUBAmWMEzWsKWRqYn/4Mrb7WJEYXejDuiAEMWzOudTdyOY3k+0u6XjKGTFf2TPkN
bMOTKFxDY5cNtduRfzs9emg62EeJsqrxfSDIV91E069xxOMDJzCguLqvi0Hz2ERy
mQv73YPLK0/jCyhx0oexJ37YpJQj7BOZgpq9Aqfq68JCiYkueJ4tR7fE598JgDlV
qQTqaVYLjl8z0rmAl7WL+8F5Y4mImZOuEN6EEdXvQ64rQ5er+LgQJO6fTr3MnH5p
wigsPId/tQWVh8haO4SnrSUuv7ENOBbhztf6wT3Ue3luyR3G2RZ0zMYdPH45XqyE
WLXH8DnwTEpGpLJZTYaXg/9zBpFGtGBxqVabmKZHGbLlEsgk+iBKXChS2Toru0CA
KbVYPEfTntXn0RBjBibHksEQ2HfHbCxLi7QI5krpv0lElZ0h/aSbCGeiV4/lG9vM
mW8ufSkCQ9BSSfT5z2oEL6XrNs8xeiGnRhptwUZqdxwtCbolR9PpfCE6NM/l0rfx
OeZ1V6T98PqhbqV076JT8f7V36tXUUAIO2e0F7dYh1HPcYNBfdXjzFLrze6E6bz9
Hb1ajTHapVGxQeAlskTkMbzNBdtK7QVO43VRpnVwPlKtKpGOTJm1Ucfl5toGzX6t
QK/HjFPt88u47SbO1c0gRDJz7i4bqEF3hgsm/LY4vTNZ6xaGbFx7KDMLJYFPgaJ0
3UijES+GplgDJDg6bSYDV8P/GKwhDgGCDOtZIy7F3YLFVszx9cpnBqpZ672J3e22
vO44NmmjFu/nhwF4qkNU3UxRKzA62/YHESaJFgnV4Luzu2dSb/MS+PmyI13S2Yeb
mujDT3KEWcd8Mxb54jXOQxAHJCt9KcJhb3jdHX8z4knfm2flv5fjwo0kh+suHOw2
u3q5l0jQErgwj/FlkEfFW8go8MBiCfFeL6CXnWiU2DRPB8nMXyHc7I8cFFHFrwRj
AVZ2bYYBip038qVTtK0uxGuGfmX+x2N9dCv4zT/DdLDcksov/bNCshCjqUSpKZEY
8vZxor7K1tl27cEqb8hILnWyrSi2oK47heKxKgMj3hejKsqrIOMIUGBzyxkVNLiC
MlpaPxuL9r5jXmf4UW3rp5kdYOsL4Qu4qM2AtIK60jGodfeO6xL/jbUVRV/KPfli
Sg4hgkajt+x54FKMbd1yFcE6EoLXgwIhjqbL4Mm7uRS9JLL6cgpRh+V9i60oDIXo
S8tbIdMlWTYVpbSd+uW2ttXw/31IPQ4u7cXjj63F4/6CRVVqMzkki68UVtAbovrg
b/RUbJU+bXs0tYf15w9UdsSeyNS3rBl2/s1qHU6IKjDzimZPtOWkwwNd099HUDgs
28IstF5BVEHJDE0akHGaD048wNUYTDzm9BfmPWKuGIRYwAhFaEEKDDTFiuBIbphb
gE0aINo/GV5kIkrIQFLL95NtaK5N5b+PHR+yw2Mag6CP8wwrlnqsS9vm3fXDKtap
dC7hy5A41olVbKacSxUfyignEofBQdciZ2y6SMhyhuHuo0brx12LEp7dQfw13X/L
4xBdmE0114Qd8X/cXUd/kWlWK539XM0ovySMIDTmxCpbsbL7DXIBol4nj1T50Huv
OiYVSVjogXuO8iX2BStnO0hjhvDMVangi5t/3MFYPdHHKHKziERz83qpBTh6gSma
95En0PuNgYE3Gy+idloEq5n7ykiB790Gx/zW4wtr23pQz7EdAUiOvhg6u9WfCogr
77l/1KmmER6Ng4mfkI1k587nf74X69tDWTC6RwHYRFQwM5rGQHxZdllyRu41Spu1
71M8YuAwBU4bSSt1Be1/9xkrzCc7lChyboxSqFRKQ5iFx1/yAGukY9dn1Ttfgwrt
2XJ5hq5dlEGyhJ+O/rMkkggzWRY9IKNdQwM2Ib11spuPB7Fkk8z+c/hNUXPSNGyY
LRn8J+ai99rxysKWgUQMOPnNAWNnC6fQU/dnmG3sAdRGSz6DsXcMv14y5cFcHCEc
AtHc3F6V3GZ15XzOEaM4paoJu+XfNimfP2nYWDgu13RkNzdAhrMmoskYdgsb34HL
orSyxzY/jP/GZLhdMdrcHyICoOTV3OXcBG6lZAif1H97gPS6+8CfRJToFI+0DQDy
NdwkKWaTqBWWF3YAz7nwBMKJCF7/Dq0RtOahmEPgLEIUCU/DZ4kOi6UD383znpiG
AhyrwJTM706M1gXWGqolfOtFzqt53tJLRagHZ0qzNEAXVNo5s+zK7dABcsO7TTf3
eE5viKw2CALifPQNlRNuHAFQ8Y+VFcYplaTFHH9iC7WL9u/A3t/MvKHnXoHi+vPJ
qcjf+VtqHwgrDkamffzL/345h5lJX2mc749uO9z2kO3JIPpp2WBM7SPXFnbFvQh9
fA9BG2HcR9kCevaCvkOb3HtjnWX29L1fyPW42RJB3fRfySEUBOulpNRB0fxVg2JM
b1RKg2HFMpDiHgpHOl+tzG/xqv86Umid8smDPtDo6OiivHcmXTZAK/bRAlpE5CtP
t3sSPOlvLxPB0M1C/2ax4siOWN6NrbdUNR38ugrqoq2JgVU5qXC0jZgiumxro64n
XfPyDcFASHKCqr611InficFCqruigB2pfFUoJUBG658vIdTQ4cCbAK4GaulCj8bm
SpWyy924W0gZ6B519KYAhQzCKnqU8mcXlyBNWqR9Y0jNODDqYyG2SdjrW9RRnxjf
lYex72dzjcwN9vKaLLpA1eNLwE/u01wi3lrOu9jB4mWqBNAqbDYTK4Sb4eAPu3eF
UIunch4RKlr5ECJo5JFE+36TUje245t34/XkVEaBnqtg7iNb0292kvzPgVfbgbPG
8bde568KiQaZgTQKF+FfkTX+KLrsV274zWzAxzvrxnsBCRFOyvcya+bEiBnR2LkG
A5Z2iEy+3TzPYiP1DWelSmzVtYlaILKvvBwrr59LooXMvYzfLmBIId6+eWRs///I
TDfFDaX7/E1e/O2092AlXcfCNI4Injza3n28nrR26IbIF+DhKt92s9V7ylO3ljvp
zzoz9KkUFnz2NjtGtUE2J7jO1iSho7eeA4W2AOUyxGWyTjo3N0oC3Dg55T+T1ikt
+EjK6mRAXCt1ur33PiFl1aLU8M2VT2Q5+ZVJWMKPj+zYTfFhVyqGsVZP9omuaIhN
o2dV+NYrVoe5mDDhHkfDDR0VZ3B4j08iiQM/FkFlI6RxgLzQ/flJvlb8jOgbTbO0
HB4IZTr/YX4zn23z2ex04N4OouACbUrL83NenscOiXX8wdCNOmcce5DR9FbDdlc2
e9y0Ckf4d2bAiZ2lscd0m+TYnuxbOQalhPwvaXRs9nn7jA9yzghOf6oV5Wy43S37
MeYw9kpP9DpHOFZjiBKA+KrJihl4sXqYDvzdRxko5daYpyfLBvaYOnOD/Y3muW2w
oTOd+6oTL6Ynct9sI0D5xIIKlUqMP36hPhPcxV355WThCsgp7iLbXA/DXJUbVgaU
Rm4q5t52yLS1A5aB+VXMv+XCJWv8SmoSGfFnpwKev2Ij9/dJs5ukNJn2xAZfWBuo
YnTCRbl0zKu2RaBnpzrbB3oL+GX4Dtn2e6ZpqroWbuTdo/cwzOezjeYNKF+je3Bt
Gb8sq3v8ZcfudOoyZwQofBacC1CQ29SRqNqwGB9eRgjLdxI4N8YVz4MvrL0pMlnn
EpG6RMS6+u45gP3/B2NpUVD/IqwjG+Z2WILOYbZTaJbIT6NNghqcR+e7IkOA/jb3
n+500Bdu48dP8aIexjqljffK1TvDU6vQI8YJnf71uWjlF5w4+VCJATxlUevFo0Vg
LxVqkM9ieaqgI/wgnR/0t0M26qgsKnpzx9GtS5xxS3cye79HCdFqMtstw8ti0KY3
RYQJLJlwYOvI722MzcD1p3GVcNmCaKhLSbvMwU9TR4XXKEYFKcFl7YKRFSbTwzXY
kh2XnS8u50oxGE/iiaiAiOkOQpRLul0Qckvr5bwAwfzMulIhox8tFhHc7IdrqzwE
KxxFSrn38MwFZyFOsQP/r0/GokbEx+u6G/O6cXkGBWJmcqfqYgK+jNzHub4008pI
qnidTC5tNEhAEentFGIokICrQPzHDfoRAliMHMSvl5Mc45m8eBu0ygBmhhtISWM5
azZ5EbFWnnltnkNNBwPSjOkdzWUNI/g78AYnMcnDimE0d2FYQSe8WCmnTmC68CxY
cTbuwnwUL4OMROp3xWce0DVI81HHVKUxNdxkM6rneS9e5F+IAB1E0xxlWEDp/cEH
cwpaTdTcNwLa0JKkxOW8oXgl5jjzuWS331Hiu0UfDM0GcqXurGTTVCxh/04gM34Y
YE1qytAE7oMVWuvgv0fiCX7/u+8OSnw37tDTLPqqkz0WwAodcaGMRxhGYvi6Wse7
LaxAlrHO5w1Alham5j1S8s7hYiDsLXd4yS1R5W3FGoYMV6z4BepBUyRQ7+ezjtoc
qWrj/RMt1rUA+HyMhjlOtxOAG09o4lVJEJHEsbzZg92f1ZUqOnkUBZ1iB7R8/Ium
EGpPAsBh7KLPDRXkRKuVBm1IhJOgy1MWAyGEVA+C9b4IkDA5jQ3+qn6PgXkc1f4h
9Lnoho6EDPNwx7bJ1j0qoxuR8Lmy5jNfKkmc3LY3MFfdMZGSfKc6xaHcQh9ZdpPK
g6UyP9UkdpGzcrl6o1uEV7MrGj8umlItWUn3CcBSnhQSD/hsy6gslKWlZmVXdiI5
0sovegxYk0bfk3keY0/AIn7LMFgfIxbARkdd79RJ29IB8rosOcfRULC+4zPQM3nA
meqp63OnjMpMHM0GljCDo9Xgy1op1CtZfNFFvFZg33IsfEy7Sr0vbfM+3+lGJDYZ
0+QMh+/wsbCVyhz1Xe6/Uv3XVS4kuxvjfKR06AI09EMa3xI1FPmIaqSLvm2IRMr1
+fi1j4nZnpnowGjiTY2ltvlxrcqrPhVimwjCrPispHAiwvVLCtzwHhtJCTJ60BsV
p0ce96hESVqtM7u4JW0sbTdhHNTdSNr3RmUSQFHu+pBohPQbNziGRYAiczflUJxA
cs2Q0IKkJ8YHWXUqo9cNzYKtwBkdY2yUvg3/sxv0VfRXrCwnPm2B8s3h9zkIMqY3
4OI1C2I5xY5YXvxQJJS0dheSEZ13dwR2t2PENHI8V1q8fs0lNh57gIXSZhaitYsR
rnWqhnrqy+njDyeMl+vio+GkodAwKVhB5ulTnQOR13wCGWxOBVmWIk75fmcKDN8v
lpYkUo21J338tUNIgrV9rfQyyaMV7TNY1mSjeLHQr0y5beemlKF6qQd/puBT2dQ+
v5i38Mr1cUpV/NKKMJKqsUNjBrxUJQueqccgbk4n4qKVNtmECSulxjlsF7O4vkrE
swnjDReg5NQLX9Dcup16sr7TzQOC4FR0eF8Ey+7vCAmRXzbbsdRyQlG3T7+wSlfd
QaXktj/FIVt/K8F8eS5M8j6Mc+JZm1YD1ed8VI48i9bI8/ZrBWHU+/apk0wXu5OR
rGJBzmGGamgYbmRc/kPAzye8QzEf8NN4L/Hd6DGD0lka3oc3E+UXOMdbm37tSlRI
n06SCs2CdXAXkjXXKjuSdpoaxlBcJZaH8BJRK8IU0untyMG4YwXHDTEh/qN+UlcR
Ft1V8yBqGfLbOgcf0U5y5eUYFsQuD1QlICIX6iQmgZlIY0h4YIeB0SAAMCu0AeMd
uWaGAmBvlB+ZznkbHDXlQfnm0OXzMhVvxvm3GX39vHNQIaPwUBjlbDPrnbbF3OJ9
0YXJhxcEY5A1vncSA7fwrGZ/e5tc7UF8etsB3xQ0CX+dvZvFpM335s+PtBwE0I4D
7wEknwB3a/LFSohC246RTCaLC5yLRy61P8T/OwHzkc6T0Of/4xbxY517H8Wi3oid
uaEzoutTq8YujWV1vREC/1kJjoPGU4d2CzyjSQGFMsINhy9P6+tvVOeW/gqngAz8
ZGTdH8ZXeOQ9dyoE3uZmxQaoH2oZNj/9jWHcCpTcS4Gyg4E9nlVvn5CZCL5EfHBX
DbDNi/StlXJxmx+pEpieoTtcWVwqb3CeiGl/CvqrxZqw228Spo/Vw2jw6XC/MdKl
5awt0HhEMGbpxyAtoWLC125wt9A6KpEu49e/lvSTiA7ngF2vAnzM9vTcewW8IiQJ
ocJ50qXY8ZF7WrG/lTGqMRTgDpYLrpO8Efu7hcNGV8bQn3r8kAepX/4muSNVv8ht
xTlTNDQCTES5qMvUPVoji9TmBwgQBYricpHb5zaqDXd69e2Tg38qn0MvT8uT5A+b
iAFkLpT2/v9vlvbF7SlTNUfwtaBcsrzi3fYYo9BxEBSMAig6zw1Romh31svbzeOF
j4yEKUrCHFg8P2VHHxFAn6iIcFgQn0hNV1ZEoz4T2K2zoZgsNevWj7wSp14/aR6i
DavNo24chsoXefOWKLSpLekvHZpuMAYxNuUViHUgJ0NPx3UjsiNei92rL07DO0qP
1DeHEJFCgz/0wAxDPwtdIuKxBItOU53uZ08c40JDowLLzEqpe83zXEHJp5/RQf6U
rtH47EEgPLGHo78z3rL/Mwe3lx2gzHvnK5MLZK8rXChQfEVIj0I9xHA191D5nx6p
G0kn8JMO9oUhxd572fJ5jIQwckztL8OPdcO7fiZ97OBM2yFQc1PWQoEIZr4vUMZy
+1FNY1eDtF4YWx+4q4PFEUoIrD/zxujjAvbHEGXgfvyEt8LSh6OXrlbZpC4b6V8a
4+w7fYFsknti3ija4uta02FsN7hKJ/QDfhYVICXmGXFLgZtI63DJCj79LR/AMo+d
2i3jj8U8yQl2XQ3xUjV3ky0xHo/vtdgSDgk5HCEP8LveljkeeoH5WfyNtKyh8JgQ
vA4HihmhIyui1CtnOVjX9Y70j9shLLSFst3pI4PbG+TrCj4aOscTBfaY8n3uQy9C
HEz0owxN39YcSu9fM0Aud3LQ4dioIjaBsuzvJ+dyeo1dQrkdrsHJLhwBEUaYrlkw
lMdLk+Yvikz2hEN1lc6V9LNMJEXi6qDiosIc/00ibYWiSGcRqG+n+vDuon02NKmn
LPqHk98dp9MiRcVMn95vMv66Bl4Cz4QepseqGNsC5CTf65ICdO59hO9laQXbX23j
224Fmt2ITl4HCSjJ1kLW7RmsTEx25H9lAF1Tic3qCqwFx4AaAlT4NKfbeEwqg0OM
2/MwXGqlDvLET73GuM8VaW2eiWhbSLr+vnWZhBv57Bs3j5GsnsbFZ65HCjAnQrDy
ZEoMjy/C9572H2SBA7VraJihOPBvFIVuTrtEzjigWsdP5lCxpG4P03hr8EZwRwWn
OVALYeMy4v7AO7Z1ANG4XVRMiQ1FVoVtwjKxbhcKxOPVsPyXyVo0dhWHtykbH8o4
DY3nxHu3mwujKEOjsN2/RZ1p2/45KH9ar+mr8raOH09rLgc4yFk+L4I+jwKdurfh
8jFCmH4sqZf8EDx5qHI8rsxf8t+wFnLIxqEmiTKGtCkL6oLFY25+Pl6GrUp6B7hU
8Izg3DXw2T8OdXbwMFWddFqqGl3iJSdbmzB9uw1iNJrlrkcM5Z3ChzM7Y2JJPh4+
OOrQWXlsqyiqD9GVejUoFdwVk2k5mdW1BZEc7IpyD3VPfkdOiBzxQvE8sgHYAeLn
GgFsTHuIvLwzTgGve4+0lcTTRARVVEf5lXee1tFnqk055DBEco9lElPXzmrDiY0u
st2bF44br+vgsgZ1I3bhM/28KL+RMf4plvUDaaLMLAanWoTvN2L6+gIliC40DhJs
75+yzIFUoaTjNXvLzvgf/SPvE6ft5LP0Uzoz4trZodLLn1JKLz4002LOF+wCt9g8
V/glnZwG49Sy5tcv7XdZoCBZH6UFSsXXv72caBYzpQLTIy4akiWHMMqroubz4nwx
HqBBAzhjXHNEEugwXNZxmsAaFTWgrQSbXYv0RdwRRxArQQac5kgH3J+g0lkmf37h
ZipcKKnVJJlWMsYr/wnD8/NXxns3Ss50Scit/Sm39WC4XtgfeOIsAuZrbl+GafG0
+9kmkGbskFqERm4NJpwaqfPqSLZY0QR5t2hiYynX7yWGUQMRim332giGe4mV24h/
GyR6AudwcirouA0GPNiRB3UfV8OI6WvohkJDOTCP8gnsVMXgpl8pmzfdgXwqVf0R
fHsOfikslVbTBbTu2aUQuraafabcVrvidxI1QrmUgvALzcj0Cb5jEODctrp6Rvtk
u1rXd4hBT8ubyr0SRNIG7I10Z+JWIYnp2UKWcmgcrZDvWqmwF6349ymfJveOGdeB
LGsSeGLDQtpKMH8mnPhkxwFcPNpVoC3c7L2I8FWiErREdnqhpN61+fyytkFxsiqK
ygctahafNVexGk8777+8aiA2ZbwizOw2cezE129UAjKRePxJIBPF41QwGQBkol0t
9OHy6sGXCcUQOrq8igSxagW0rUPaNkWGtGSGWmm7mRHtN4BkLGm0A/eDtfliyCm9
IVE4I/gf9dqF7L/pottuZYYyS9b7elbJefju7Y5mWHA4jlpSpMVZAOPNjxfL8N90
6Sq3hcqM1knzSIAI/WqNdNREokOarm/Rgk9uBc3+oXW2jAme4SZCaHhHVpSW+88Y
xV7qNYVBmpQq8bx3ww/Nk/CKyn5V1VhkRa2SF3eOblRVtodhM0xT6uS9YtTdFK/S
wdHShi15RMSxu8jfp/MzcEQgMV7g/6vZKaiuuvjmAGl5Cz2qo7SevdTbTwEXqFGX
hsVoVKQp7Ml6MBYmZkYOCmKXjeaIFyc5hW4EzGrbbyML+ArCN30YDfIfIrCyMmEt
FF5sxMbHKfM+5fMH5VnqBl+rGzjqu0otDplWTDxdQwQQKk7H/rLYaAhw1MRYpo3L
Xe6viEzWFmFBFGmD3A1HIgXIl5Vn0QrICzb6VbVSL8cZFAokYHbUpQ2xDqo2EaMA
g376JZtkmJGaXXaW8seqne+SvFiOvhIMWyiTP6TXBWEsiK3j22w/NVAfZCBP+zpB
N+2cCZSbOfL2DUQbkU/Nu0iG0lg44T5pTDufwyMYAv7rDEJZyU3v9U8BjiL9c4E+
DphWg9yvjdxaKZmLHN2pN12IoeK8VZ54nNZNU17Cbz6v86br3xy1It+aDTG9HSDn
SbibmHjSxbrUn9z64M2oL353vULiz9RhJhGQcqcy+hryEtWd0lWekQnD94Qd+KDT
EET8b/JHwD8WA+fwOqg2hptqFFkRb9WxmMl3LjIR281sfegUrE2lCUZ5J6t+NO4n
Jak9ZeVaYug9oGN3XxKzCSrSbK0KXwgDO/fYrPPPd/0Xfk2U++OPSDNyy0dLRv47
S7gNBsx9gR61b7SVA8RXWyQnBN5GlprTHut7B2GuOzstUAcuB8AgLiCvmTKQTgMV
/akXa7Uqv9de4ZdiBh+TobSU3BBpkHGFoPlI3fX0k4MWSxmb8VdCw3BeTNm7dmZA
lQpPmo8eWwEtq6N49odWAX0krw6mPLbU5/JsC/lhOq04pZ/QfSj/A3u3lievhm04
VC6/ZOxBuGLD6oQNu2Bs9DYp8nN/ZI/QyVXdm2lS79xJbPTYSgv7PTj0d9tl63JG
7ZNTBkAOXrELzL9YqusZl9VT91iCXZbCBxBek9bCUW7CodKVyh2P6M0PCCxmoSTn
27HnStqrlF/x9sliHcea5syZB1qkBCMf2+U7RynenC9olRTsXq0+dF7y425pCGhp
3Zj/raaug84u1HG5brvtYs41FEQk8QfGy9UZ5bYFtMUt6oscxd4eOX+nUZTX5zlM
TMkJHhhF0nqqzZbWObFUg+i+ARzZxD525N360RWhp8Iwxefw0iBjOaEDbP9vjtvP
tB9Zl/uDUjfv+RVfv3RTla9wo39O/ghr9OKfLA+F9sjrkEBaklpo/MiEzINUhtMB
+avv/jMqiF4OQ0TnYmBvibDDwNhZvT0ku4u61vvGWtaQF7oSXEUgEiqtWT9YOhbm
x12yv/ORh/TSkyc5fTUUIeP2pl9cvKmVi0Bjoq3KGgSzkvP4AHv485G2WxTppKzl
0yQOzglfIhcTeWjDM6SiQILPTEJTKXgFeyLQNoqItG25gC9pnmnjXH39UKcX1ZgO
q04jqs/g4Oa6UyNj9z0luj7sV4jPCqtNoqRcCYTBJ9t013GavsTtHYwpSkQi54SK
JF9iVWY5UESljeGTbMmBbA5R7cz6KQgg0SaOPnINwvWpaXD49pdW5lX5jBc9dKvS
umxaSiUpeiYpMu3yb3Pn4eIZ1/VevtHuxkSwQsxvYKIvN/+ysML8JS5MZJGE+1ag
h5qRqJi17mRprGVjrBZup8XXESY2dAbKNetWETnmU0lnGaZwiKZDbfYWNJqGDALo
jMPDH2KdOnw4Z14Ldv9VGLkYM/8L0+xOa0dekVW9tcSBD2F5By8N3fLBVuua0c74
Xcn4yMeKHSEWn2zNfQdRVVj2kxG0HZSejaWSX1Wh37xKBKt58CL0JbLmSJdGk+ny
I54xFj8V+VI+2DQh23s+SEtemZbEM4+R+wZURpLPZGzhItrXKrBqUZqhc0oNvmrz
YdTBQ1Pi1L4UfVHfsjlinSSGtv9cqDx84avq7EYFzhSWLST4dWuU2leAUQSv0uYu
hp30FhZIY0SXSTTaT86PFZ3dDCYqWa9Ae7BS9VCEu5EWD45ma2UC/ZPbKYw86NV2
kxFHXBOR6HspWRqd8RBBopfzYaceCJjIoJTwzC17zP3VhiSY8X3+6qftfnecHYMS
pNti62iKpb7Kz81SfLaajTdRR/mno6+YqkKfTRZiraZuVHyrtgRyKSd/+DYQiP8E
fzBS9/5tJapPRfmwCrSdPObT1Mwba2BzDSxX71GaxOY5Cu4ns8G1js1nbHYURKoK
a5kQ7lGVHrw6bMRL/Tfz8m1dF1WrwBur6cJPKG+O+5qXaPuj1qstIwec66ibvpkp
iulANxCgsaRT1tTeYRaZuRKe2nIhB4HxGE+3dM9A2d0LmHMwMAwBs/DuzyaCuEov
ajOM2MvXBSEwikLOuy9TTm5mRgd9tG4se83YLAl9O48jt6SBNLOnparxwy6pfriK
zrCU/tehgDOpDOnHHG6p7BXqE8J0FeYzbtXdhBp47snhII3Xf6NYKSAIqY8dXw6l
TcejBvLbyl6M7PQB4uJmb9PWGeQu8nxwSzNsJ2i16h37PNuFBz5GsBroy6bEv+Em
2fb4AH4euoc1rLCChzCJ3juld9Ssr61bTaZVCfoKpzjcLpjDBVY/WLqgbEzcreF3
+khtVHZ3qexYN9qv1D0mmFmRKFari4RT9PKLIB5cIOKBq5b2/2yWM8lZnkqVvgjE
eJegW1Yv3bxNz3cO1IeObuMLyTWQDD2u90QxY1Bjlb8oCxBArTjgDGHJniVnhH2Y
nzqa5Sedr5N9S4A1BhJvcVmCxbpOJd0HxNG0OfMNX9hsvA0c673v34eD9hIF0J+X
GxHEmopBAtnVuaQyrPk6wPNa2qYkPxezudBq+SPbUQCB/Ni+2IjAXj5T9tBYC7uw
XYfAOX2XcZNin9lXLOPls/hRf07AtcZwWeI3thhicx7Yy3fXyL7P/OP+6P+pKd10
Ih9X5ldbrdp0Lc52O54L+esbKeXuQEPvYfAbPJW7P1LiSBBYbBdBirUbkL+lJXtG
iKNueKQARujDy0k9goGA7AnlXLIBiBQDq/H6kC6LVc1S9Dat6G/ppZfZupOXRBhQ
+i59/MVI/Py9H/PLXjjceoLRAXtGJFcsOwqmhfE9YqZbETPIoaqDoqwlM7bnzVUe
G4Sz6AOj/em6e4rujh8AjkdSiRw/1a5GUkd3ETb6BNJBScWWv8bW38tgZzH80rJw
irhFKAk6kkQxGjy1DgBLm24c8Y0h3WRg6xMcqsDUCm2nQj3Y6yzPL9+AjpN7Judl
OybujV5f645iEbQlDVUcrVGYpQx2psGLGJwfqavPEGrNf8wA+1T4MDTtNRtx2Xvi
JPjqzxqf6doKKreqWdzd5jKW0731IRLmmRC1IPEBJXLAq2QPTSt2jM/Gw6599UHv
KE8oSG1+NFPvvwE2r6Wb5ny/J5BFDyz4lis2ekOw6xhao0NHyNGO/GbRnAl9LM87
Yyl9SZA/FtC8nfzG6XsO+ylxdfmGmcE64a8hQnbz1Gb8/yDWBqeDIRZgwJ+N2axj
OOYmB3UwRyQ8QDcoaTexnVjnEnXTFsO5Zgek8g5Cf6r1pPn/+2Xwm3hC68SBFD/a
0oSpUaSn0Nxu6WoMHOoL8pLOpSAHR53CST0WdaoalU2248mLPxzoQhLhgiyDxgYS
7YtjYEhZgkQz56RujnnOvKTHSqBRc1DIQRTAc/Vls+iI2SXnasCusjNoRrS5RwaF
S7TSuK2JScHWrku/aNDUhXTC5zyiygUOp1A0TtD41ucM1VwPEkhVesn5dPw4Gdvw
1BbzjCO6fRt5/uSSTkTcKDQKf/oS2qUpnGAW38RcW2Vu9tukpUn0F9off8rJXsUW
qUkMVe1rvBwLv85Ih43iAfHJHWSyEudW9qm2tXBUZ0EicRl5hlfehN4W/B6HTpn7
e/hFPBlWEhElRu+oDJAHp3h4wV87bZNQK28kvlJdVBZeI4Leb/vp4n12dRqr48rH
AYmO5umsYeoKtG/V0Z/GMyF788C74N0AHLw3mLe9R+lbdE6gCzHaZDEClKVwP+5d
qJZBjdEUck1e8XNEyIMaMTO4iS6tB6dn7OKKF+ypDAEZx+qJvGxQImlniEVB2rhy
fRI0vTELQN4PNQLSlxp8K5LHBQKlQlVwmgzo06ETk78oMpSIwwe6xKdYJJMYzfem
j38UsYW2GskP2KGFPzOl+WFiVChla3wPIfY9cfYPu19LLeoGezHb8U7iJ6eHyQuA
AowkGxPebdK3FNBa3S9ABp3wiNkUfxogTvfe1KXSj/rYHXQJqHUsKLp9dHYXkVfO
aJlZ5OsXn2vYOogiPRaz/oKLG5As4lyVzbV3dqG8h+rzOTY/zemte3QC16QDdZqw
nQx/A/sUXwjAcYnClZqBgf4pd6FrK/Z2Afj6s6+PAZK7/PaAhCft+G4jWaCtU9j0
b0Swh9QKIm4Vd1rlytde952PfK/1KcaGyimp5HLniTOUOLvbm6gp8ufpiTmOMAQd
04IOzgR6R7gxAg4N75QeF/x26/13HYF2deMsCpBDugZDHt0pQuCSKTUsoclYJGyh
FbpT/bwH+nt/MR/Lcaw7dNuRIgaiG9Ou8QPA6ZkX8dVCp5Bjwu5sE0YFfrIUoqw4
/Ev2OiLF84D4pwOpkRAST5Kne2XhH2YjZkmZ60wYXHLibzSpH9HxzSFgGoQTQiAi
Z2F3Cg/eut7wvQ2MHH3LQfyytTaL06/ELyAeun3dsb8pJMREK4GTIOV2AKLwAmwH
/LU/0CaNkVCVUEmKKKx5vdMkwrzizqVZ0SkZBq2gB0EOz8ZNuYyXfYoHH71jDWm7
OnbhZX5Z+hrJch7WlsMc4Px1m/lY+TJjoBT5BTc4U+TUZKl+Fue4xmhY/2fWAhiu
JSI0PryUpFg3dJ/SVn2bPDls0z3x2yVDnUY+f1s4Isc7hE6w5am69BCppJjwK99r
sxGswCGGDcmHOoX2tWjGqXf89IL4Z4MRoE+HCIUUJTZ3fbi1u8o11UQ5MZ33Xht7
3FvQBSuKP0NuSjjlK6riEQ+apSRfto5+ue061LFZYvTxMObGazqaqD0Sbu/ixTb+
1nYerDIgCqGpEaSFqsT/O0DtDCSmZT8FDz6Mh4eAM71QREs+qiszNJosQu0zbpQp
tpiraNxKXZymen66MpYZJ9vltyWrERtNqhp7CnVUPEaBeILQzjvXVWwn/QDzDrEH
aT8m3PpXjr55s4bTxlo2r2YSPNkSVtD398e4KMVh4+MQvhvNotOCZhpzVbO/vEMX
3GqzJAja7WRMUznhw3apMYTCoDN6fNIWFO0Hgxvd1LSdx2s/5+TP6DanC8ZSe1xD
UJcWoKRsKkabZQsf5xbiIykXpu5DMvyWaV2wyzcA7fCUjBXkFqm1usunD9ngehh9
L+EuBiBGTPEuL1ZKXOpSHxb/5a1oIpjNrCIMxrai/d497N2CdzNR+ZMfCYuKFcgL
953mP3gV+spt9uPZPIySfWKOLOpOyK1OuNSrfVVhRbjuDx143Axn+HwNQ8IGOja7
c0sB0Ej3WUPYAi4Zif3aNIQrTFX/Gtda0ffhcacokgMMPaNHG4a16oOVDiW6ITZO
stSy3GEePk54OvGJyMGzkdjOvwmdGcGRA1ImadArLjzsiXIZD+vuN7AO+NoVL3BB
TywUxrW3vgC4UHfrP/kLq/35p6wR+k3JKuo6DAuBFJdRfNZnoYn5AjZeMYFb1Ra/
HfMFngRY8/IidfWCS9uAVvUgYuyGX1ZjHUWqrv4pCqJT5AgJmz0pnkt1dTy8Q9jr
6QPaAPJKZtGh/cWdB3FKlSx1GI9zzKRP1BdpkHs4EduE0gIXhBuE0lPi+4qvzbLp
QJd+8TxOkhI8otkXGh7a9sMu6kY+uTQQq5dz09By+oKpM20NfwLLYCow4o5v+ic9
L93P5kCJ7Vadnlp/KGoMdZZQI37Or9i8T/442/wchAL89WA0wfAEtGP0YaTwTwOb
+ybSXUXsrUr7+0haoVb/tO7og4y7YQBwPyGZeM793OORQJqBaeAlhMOqUS/iFAl/
qRMt4fypmBK9urU8ei9TrOerDnHjq92AgKlqdvvHJxTUJCt+YsAzOq68UJpQTm6+
5L95OzV9Ur4GAPm5wFJ7CsNFsBEWEixCMFNhc7jiXEkM59opvEX09dcKkR+ZqiFj
J6oBZ+6bdCpf8klq9FZ51yytuALYXQlsinpBE3xhp/+Q1DuG8c6BdAD0quuid/hQ
r78IBl94egzn/ZM+3MKm4+wgYE4R0PrFSsMNmEFbkkVuK0tu85bDjLMPZRSQ8RbB
R8GzD/b0An8538zyHW3g4QxsXrW0WGDPA2jRcyjfLE8wQ7MfVkCX8bNq/8yBlcN8
Yjkj4ycHxhhG4h7jbr0qXjXyrUcaJ4ZXZyINq+kR6qetWSPoRyH+58LbslJHTKpP
IprKFdpT5pafYLzIvuXEJa4Fd0frgEwQOMPjUoBh3xVUJ4e8sKvzUTFGreY0+v1D
0eHWSMQ4/xsP9OySWwujgaOL4suXyhGzS+nzbQuCeTUoEQE68aKJYfBRLeFUNeIm
5AcUVq4xN1DTH6f9YQQMWeCUZB+k2FgVnBGFEwbgAddJ63cf6r9fzdWYMeAwbUzp
M5LkWJS0VuGdy0fBjHX3a5WU+EIwePizii/olXFOQ0wgGQ9/CrpnAgQ1B/+X/WzT
R+NTpU6AABvwKxYi2p1n4eIcerXGrQga6+Rb+mQ6EnQp+IRJ4rrD1uF+8f0BuMkT
Evd9xrbg/VXqIFukzT02N72sj64r0jApdO4MlYErQOS3ovh4cXspigdrWIThl6u8
9a/uyPGD0YBmYQsP+tb/X2FZ8pjPd7IXAVzHTgCNPfL/P+jejrr6Qn3TkVbl/O+n
2MnEOgfB3YPAjyYLDsk3/OWVf4l/Zdglx+sE9trHnwpmgu5WsibnoF3IiCNko6xF
qA1gFWYIr2VaG7WRlwxfXCuk6soROzBECzDCdeuMh3pZ99IgD8SSVJE4SrQilsn2
ObXAX0dWACCJP0K2U+MLQVlJQw9lQofvbB0zFcebawd/MTMe0syyRbKnxx8njrfn
U5srrXsEe2SVpx1c8ZPlKGW5CFqOhdFmW6uRX1Y5nZXQ8WcIRDZeAoxZttYnfd0I
hfUpEaT35qnY9gtaqAXx32TFvwgzz0PfxGywfFCiCcOgT0YtT8XeGNr7o8VbFImO
YaIvyOa/GpMeKASNRbVEV9vl2kEQIZWSZ8aoV9P8zM/uYq8XGwOoUMPnuPfNZC0e
57whatsFEx7SDmzEBMvA/Jao+7CUtkGAnBVrQSGWzdWTTBwc8I9Kai1Cp7ltdCGI
+V//mctQgoiXzkP79r7HNYKg1iXl+Wh6GPpq0NTrh46SMWSolhGXvAlbi2WTMVTg
VdBu3iG269om9zNI+sp1JSokxh66gBLnNb3IMnMwTJfbCY+bOffYFbJyKW1Jqgo9
O+xXQufUwcLz5vX6zB2dpqXh/DJP5NcF59hIPU7C3gI0BeGBlKAToZsTX00u+KXn
ACOrXQzpzIQ6n/FCxMlL6Mb83r4KT0sgM2CCizsnRc6t9mqwXyoR9AFEumG6qj0f
BYXKJfvtDXzIeeQP0bHInx82SUh7A3nuv4S6Khw+FlIhECTqjRDwgwdG7/65chVI
xyrEEPeJ0OeNdlstj4axIW7AdaZJazv0NpAsYA6QNDEes71EgJp7yUswTuDWfesL
m6Fcwp8EpQU/iQvE8xDfxxgVBZoANAkO75N8JYMksi2mbKwSgbtHxa1gUgSc6OtG
iUgzhWoL38bTC4tH45hHudWIO+t5VVUQGNV2RFGatx+07hDbW+jQW5U/8CSo5k3E
Jn350pk6Jf0edzFdTyQ4NbFzJEPq22oj33r0DNjsxSVHz6CrWSaRX+HESGC1DWQa
GtgL0upVEOSkTPjGjus8R7rrVDjbRpDjZ0tVgsVUCqv5jfkZjB0FLiIEnlmreyWM
4a/f58Rygpab4WL7r+xir4ZVedq1p+m4V3ObSvmzoNPiooaLjFo0e5lBiIYKdJVS
ZBkef3GU0jI/6MRlUC++YhE0ewvWPd09/Sw4aEoeZ5UzfxRicpjyXj6veEVVzgtN
jDqH4vN8P5r+U/NJivyRr6JfszeyvwiUBB+P6pg+exN8VLzAAGxCcN84uqsTlU/K
fRwEN7hQaXD01CSpT8g11LI+MGknXlI1zveo9FP0iGPViAjtUsOsjUFIS/q/iOfP
jLtIAxpFk8M33LBYKcOmMy7tGcjTnKt13FJIQoyJ5+WDoIIBPdGrgbRGnTvBKVbX
l9/nqG8txBa4+zJLjSYC5fu41Tgsm1Rgb2psuscbWVTF94j1AZu4pSrqfhXhhCxK
cMELvN0iKwk6Xen0hqEt+d/q6ct8ZRc0rhtBiYPhTuP315tXarDJqFFllatrDBqH
gW0r8YMNo0zVkfhCFFuu+ID54Ad4NwDJ6R6rx7BaXWpnT7tKsk1lLOfotyp5hPYC
UjIHf0osMtkktvxlt9iuj5ddfW8baIZeC20b5ex4kzjPy/6tlXfeWL96XN+b/auT
6osDhks1f4ddGrnhJY7nW+oRhXqbxzJf6PRxFN0xVkUlSEe9IbrEaOEHEvRYn666
I+VE5e0nmL+rjrNTDGljBQHJgtiPZ28ewVoj+je6HBQRAQgkK/U0Hxrs4zwSterc
L5lrPPyq58zX8xRbwytirx45ek7Xwf5Tj4M0MDFBZ5NaPv/9qJW8YTUwbts5YlRR
CXZyZTWalADk0ToDT3jlYW5+U6tcai6mHHkxoOFAGGz1TIjB82yimFPLs5pwzKj9
qU+xqU4piY7PC2FehWWK9zBmzjz0kp/ZiG5f2S73mjtl6jqoUvbzvv4Ld+5OF6Qr
Sh6aek7Jqtub0KMsj07Ne2iofMFJAopve84kcawnJwbZ99O6qH+gdMLq/PkWuETF
Ea7dJ/JSVnuKMUDbnjNfha5v+gdKmfZOsgofLJ0Sm0fYIDvi55dHyOoR+YJMVgEy
ASDOnXWqV+MutQnQZByichHLCx0JlNu9Fn1sGezalU02jL70Bdu59floTlRywjpU
kp5kLLfzSnvTwL84fyhzq6MXGU/Z9nDL3SUZj97+raPjFZP9NGWisBRqdPG7uhAE
MdkjOZG/NGycNJDakcPiUdtPccsFwVawRI+27n9FeY2myNPJwQtNjNmW6BV2kcI7
2a9WQzA9KZq3AQEDr5l6W6m6ewD0c+V4OWwF2HBY0fJM8t0L6YbbKBwBP9D6LkWP
BhswLsY4JJSmsW6haUMmhBwa/WlwfSrZ1hLgKryMxwpQ5WioDJvzciOJ/dsh3lrr
2uBfs7EOx0SWA8NUf1JVicCjo7XOo36xO1XCjuMl7MH+fZTKwn58JwWfCE9XomCi
Oc1g8djC/WcRWX0Xx3/44bkypwlcTwml0GCQ+1V0BdxXm6epdYid/rlM1RpeVbgQ
V9mnXDp3hR19AGGifROBHtc6pgRvgaubptAIDfP81GmsQLWcL5gXfyLrJn/bXn/8
vojUmKNvF81DHM2UWX2RXRLTo/7TIuondiRjJFMivv/zibWljM6v/k5H/VrwSCGZ
vuPTSV/5AFpG9bw+MiACqUX0v7wbW7O1l2grJPEV37inb2/+4X7WeE2PgSKmqGL8
8fd5TY111mjPBYA6CmcYoSMutC29nOL9Pmphiv5XUz9T2Mij0pFM5W32+2q4uckJ
jt15GnMG9Nls8xs5Omkdecq18brBe+QoW7kxkPlCC9Kg/XMTVfDMmlfDRamwmJAu
g09Usqky9hiVXluMsWha3C36NF/9NoHdQUKZNK7P6KVxUiX+Yd0zJqY9gLU9jSBe
oIzlqzBeBVykmazx75mK0HjwNWRLNE5IU3lqex6mrQN996/91MS7AWkuKU6M+KvU
Zcdl+gQIeevvs3Iw+Re5bmrF3TZxNRa8xyQCgNtyB7qP84S5lcBXsmt4dosncuMC
+S5QzaXbpfh98QL3oqPf4i+qZo7mULrVwgBgMRTYK1s/0mlT0+LMeSAlCvezJMIq
kFm37YVSHLm4LfNfQYpw2sSdItQGdG93d8crZyZCmzhdvuG8Pej0VqThLxtUT40C
7xuqEOy8iYP6jGxkTZ63g0reVHrwhkvkUNMQ8ZD0Oh3lelXxv/xakhsdp7RI9Znf
8MG+b8PgBWE/TboA9yjCoLXQ87aV1+WRqy1/IIvP+5XYXmyoMDlBcOUUUoOD61fA
w30430aKRxI/WrVFY3VMImbxb4DzYUcdc7GXZxezVTz2K2eaV5jvRcp8VUBdGtYc
JkwMRW67MFrkEyuj6vB/OVycd46vi0ioEZqk/ajZUAoQTplHLQDG1uK8SnDRMOuU
KJ8gsuMTjGJArQN0XUEvrD78ZFXYzTgf2IpXR+3xpZVG2vAQKMg13XIk11WPhmbW
0dXaOC9x3vGSgiGlr/o135sB5QGNnIfkVr5WyLQAPEKgcdl8/XqZ6UtgtEZg55cf
mx3V8Q1LkpeH6uuNCnn6FhTH2DeIhnlL9SK8lY8qHIlmpF7/KxMYD8UZbgdU2EtU
V0nVxBo9BdwtXbsQQD3MFnbZucOimI+gHftMkfMtgrOQGuGSsDafe7tiQTrLiySG
QQWOh5PTut8b6n8VmuC4hm7c4HZg36OGVNS81uA2xeEdTjQlkv0P9k1CuMUdgKi2
n3q+DTAbwgTqV4PvzYSZ9v9bLIWA8cJl+evI61KdBzOT2AsnqyrahrKnQBsecu3p
yI3jjfbGHRAC7aEeheL82kWv5fLUaGX1Q4ENJ6RClsxOBqLptCNujPxH6kEDaHRu
LUA6mlGy/XIByME3a8i7t3zYHkH13svpZlIhRX7fMiJlwg5C/3qnEOhANpiE1PtJ
/PyWz7gO0vcxCGhoATvPjqL6aLsaIqMnsulj//iFEy+F3IZoL/Wl64HtlsgggyKJ
eupsOZEixWl39tW6+9VFwiCZKByr9m4/bRpNOAz4RQ8fwqw0ijI2xU+LGlZlTkOE
Fnocra20HN78UhUBFl56nru7lPg6VT9R4fhJkPIw16XA37lKkDT4VdOGd/ZDimxw
20kW6m83Tm1Ifpmgi84hCpBs+WSnUlTjrrgzhBvfmiI7jCnW3/P+kWb8xSOubAUY
TsrMYwYNlCeE8w8McRK7p1xCH6LcMyU9gBYSrwYG0zt5ei0kIfNBECWKQmGGmERT
7DYOm/MGT0+9d7tnj2bIf3dTSn78wU22qOO7BwZcQOSskRoWCe368pJiFMx601rg
/qkUb7IL/Z21qy52kDm6jL+JdLHPfh3G+rsahtEmSBOmzOG1L/vfWWT6FDhc5Hz/
oObuSC2kkPik2dS+6O1NfEIKmQIyHCxjKdMWakasYBM/w9PXkZgleFu5C4Kt2NAD
aOnF0bgzRUKe3EdeAlEqBOT+d6D7u3zKMcjWxS99/VPVGn0ygBvbyTl7WnqmBgNO
Vqs9laNKAgg5Ucy/AYmsiEQ3gARogvCdVkKx6W24NbEfM9IU1r8Svqc85P/h90To
ZmbzIGHLif0cvzMsbXi8XOYEumdhAGLx50/yawqpiv/XbnH55BxvXbyGfYUN+DjQ
Aq1ZAV1wXGnIa88k7wsX7C3S1z/HOF3kEdHt7hWL27BKRzqjfwlWrOB6mGrWtXww
jeK8+L9MqVLA049xdHZIPgRELg7gqbVMUyIQyXihqL49Sztwi7bB674X+RKnIMqb
Zo+gxefIbVzWt3XrXCBIopaz0Era3ElXS7x0OhzmIE2m/JAfczxtY/dkz/LD/TvT
iDYHBta7+c+EgJzwExoYp9o8KTqYwUxVS+gF6ERtQAq1bfspQjrNxyOT6RbzSfyR
NTXQBFTtq70s3tdXdCaXqGvLKQC2WLoHrreyNKankaIZpq7hRwXDS5A1wP/7W/uW
rXR1niPbUP1GZJxcrd/bMYxxcJvAaA28GZbJmbGWcfu0LJTT8igS3PO+dMjdSl4v
kiX4kU/UgY3b69+UWZ187cZOACqBfHUva6koTGmDYwjno94BoRZCQloAT7b5vjoS
9QrUaKFFYsjuoPmtfBryJXl6DHXC5+zhP9cDoRXWSW4LY18ykXi8ucypvDmF21EC
d/BZBfrsPmhq9iPERvUB0EVJ+lqjcs//sYLI0YO/FTSLBL/oUsoiQfbmqpOJEJoO
tg5M6r8JN59ByvugjdzK61akzDTo/su6w/P5POXwbnQEkybYl9ZTYLjk1lZT6x1Q
y5ye8CGsqtObM9niDovzTwfv8eUpgmu5euPXQu6mMdJ6in2ySEClikix0z7CW7Sq
9MepNiX+//j7l1ERlYS2IeR3RsWIwkQwk7Fru5o6CbGR+uklfnkOjKhTggKmB7uC
tTYcq068zpp19njBAhlzaKTuw3M56rewXq8pwCK2rbtbgeVRCWx+9jRNsHQIUZa5
wfzOAHPGJ1tJkLLOcw9gMeZ0ZsMcY9JlNaYAfRe8f1QAI9MtA+ueVVkH5HMbEKVa
Z+7QKXz0A5Ed3u42B1PmaOMRpTKml+xtaNyeehRcgaz6gZ+WwIgmo1HDt+wecOJE
zyJ/c2N4kqT2Bzvl/3pARwECOED9tTwHsdVNnR+PkAFjB4RdFoZ5s0ztpc+Zyeun
HZMpp3obYKE0DIIBDqbo1TjtvHg7GYK/Rb4KhmuABD5lwCmKF3xdovf4rEDh+25Q
c4JpPrXVjt0lYkie13VjAzlcws3nHZwdnJRG/ovNcJIXovlxV8hBrL60nWIJ/28X
ucXVhSTAFqotKpvi7ECyj3EnHK5QFJDRQMKgzbwjoNIGNQYUF3QsclHc5o9i7v4W
63MIdsH9a7ddVQg4XaS0YeX1CZf6mpZOkzPqi106Kf3lYBWdIojHWdJ1TtotF/Gp
QvrTk+LaD8TBGdbN3vNcc3z5uHoJbH+KDX9UqAW/gkHqhwPonq4Va6RJQVHukzWK
fCkNi94AppqKq9ZCQHzTV+hyvcx4XpColJANS7IiPlYTpinzNkAZHwBUKU7lN2Ah
mU+RO6lxaZQIijzFx452DKardSAkwsZOr5Avaouq8u+AdJPEKnC7TDGTkravtjft
yx/Ue6QiDt+AXikLKGdBKRc3DWhbJ8uXZw0Lfbtt8swGFnKqbvcmrSCiNqPJwgW6
vrkPWVWNqVcBEPvPx+K6JeEzMTfEGNpcJ8GW+epXbgkK7X5TgUemgtqKOzA3lPLe
x9yxwiSxvEpqYybYFHdgOX1mgObyU5lS11tG2EsTnD5635FMKdz1Th0mEkSZcohZ
Pd4hOgYus3EAu7r3YWLZM2heL5o4TgodHX8BfMd5h1u+Wl0CMtD44NM1VWws5/J9
gLWfBqpqFOvSKVznY3EcOPXvNJwiQWkz69Kb/z3JRzIcW0f/yhY9kCXNeY18SeN6
HCNxRvl+nz7jO7LQCGI25a20vooFW9Hsyvy7ErM1rPwWVFd0/XsEqKXBcrKUaetl
PxRjbBN98j18R/j6i12/CKXCGJlbfKQtqCU/4rN1MBwf1qURiUXg1w8cnlSA6isc
z7JsOB1t3i4yg82434zVDLqtxNC6GnbiiniemaPP/N0tcHeyfr1IoBiJiEvfQYfG
OhYApAq8+FNNJrvc0LQrj2DRTeDTqt3FvfvFQrXOzw2Gw4e4o/1b4XZzFdPtIzUc
mtYdEOqpr5gR5bN/KaXwPzwYDknpp860M94lHcNg73yPBg5B9Cfg1CiN8Dmkdsr6
38wN1xvz7QVKTtmgr52oOj4Rnl9n0dUJuEn6JgeDi5+l6RMaEXChR/iMcfRmcLDU
V/cHb0MluY7tk/iTRIVIYbPve05gmVZCJ4LOkGCcsCkKyL1vefK+CPZpfyUqFEg1
4sz48flxO+rSCa27VlIqQRmdnOm0PQmnEGTkStMkqMOi77ZHQ0H+SAd15ZTU4beQ
Yv8icXbMNwpkghr9ADYuVSEVMwFDZN0E5Euk0nVOqzgEYwNVa5mJ55L+4DDxaW3C
BOlSu5ex+wJyC835uy3VdHAvAPAGWSKomqHS6c5a/koJti6dZr4wzoHlmEuAUVYt
SA4/E2i9vsKB2Fy/tlPrPk8sp84D6FrWTg2bBarBao2wNpkT18oGssnNvST25XQN
yymFfIENNFERLqnNX4QSCoTsgtJmSURYb+Hw6QsIpLBxpqrXuE/Fx3PAu7Heuz2/
remX50JBMSPQnBQE1DNkrt8fe/yKYtoqz1asZ1A+1mDkZufcaMie5d76XCM02mwt
lai+tzYIRl+V3ymzVzzUCn2w8P8UP7QNyje2bW4fY0jq7w4H/a/ZEPfCOpATWYEc
Fz/Wv9/cCSH7yJT7X9vo4LKuybVA0zbyBKv0VS6QeVHyKr2tpiQOrWcsM9gPQPRb
hcR+3MtW/4tzwsU6/jCKBlryb5n+nXwScJAyE+il9yMOn0w5xiendYpvB2AMF79h
PVWeTkWCLEwt6yDzfo/Q9o3m29jUbfx5wOB8ov8Yz6dIXF4u2ChZCk26V4+2f8PQ
+DYaszSpWaq69ZAsH+LWJZILSocCqIAa9+tVNuJOjx/cCHDYOIcO0ieJcg0o94I9
hmdUM3OsTQMDX/a1+4jZnaC43l2JzsFjWPAw3UAEFDBTDUdJebNf7JU4qnb8n3B0
rAZeeSEKN1WPK6DiNZEt0H+1NCuIL4cGNLTHc0x6VzhV4EAZ9PqtQ8M1/8VlnHyM
wrcVrAbVOhW3eFL53qb0SR7Ik2Q6tpXtxASri9+STm78itFA02mgoUyw1EOE+4+H
icZ9VwT+U0An7ailrpdH/9/1gUV704YhkblZDfRIdcHEIDH0B2QwfrFajoVjnek7
npoVPedjI0BEtBLeYjt6yUAzpDvWVaFDyAeYcnBkf6VAtYLOVzdlgjluKxyzFjdw
zPo1MbhyqUyp9O4NmZPJovGP6gsxyD+xTJ3e31yl+0ivpsL0dhb/dz37mAqy0em1
ZFoPz/VN1MzescO2ULOcUvCIdazCBw6ZNN+NG/Is1uimvWehS+A2t0Ty4f2oLYKn
We8rrjzUJP4N2YPi9d4pY/6jAzv42Q/L31OT/3efGl/ctr2+l9FdLCZRhJEv01w5
zd1naNLXucGv2x2ISzuQ6oB5jm0RCBS4LrnCDAuokCRvOmogCdgco0xHvHXKGwhg
gcJeNOW3tlhIWhva7ncWVU2QucN39xP/Sa7LDMlZAwz2VGkNohqok448+ysve+Gy
y5KIMDQT82WzmM2ix6hGDPu1MGYTPWGWHM+nf3F/x5XpPTKopdTLeonkxlaVeChl
C5psieutGmqev5lycH9ldWnSXp6TxXd4MQrF0YP3UlRx0uaLs2R2pPd3QDo9+B2y
+fHsboShbTa/yq2/92zyHor+dmb0aLtAfzidxT29mByo814Hx6AtusAFId0VxUgH
XQOFWEVn7G7u2V+Be9j/Mhuoq4jOH6Pw52e7KMso7HHWD4+ETzXC1nYZeyPQ3nU+
zGk5244Z2h2CLUY/eKOwNLKMU62P77ACL0ElWKZmdhTysFidAr09DnbAUhQpPAMM
/3MXifsRAiompNtfcGMo4vy5XLelN2CJ5tek2jsovymOh5Ux0m/kZGE/qtEnNvua
WWECyPnmIE69vuJUtsp0vK1y1fs+WDWNc/lMMR8UtTVgRmGVMtATxZbiVFUIjWgN
J3PSw+6osVRGbH4vmqWqVuCC9UdaNpYg7eJ/XgDij0fiNNGiuNb2feg5te+IUC+Q
2zO6quKbCRNmStILe7KESGfmNAHPsyIduRPz+DrAXLEAxPRnWEJW4BRoCYeJ3Eg+
biH2aq65aMwP4Hmyb9XGtNyfiKea/2XO/67YCNHvq/uMrJnBg29g1L8dYMnEOU24
jmzoRHxwcjOyB5p7n2TX9YfOnMV1yzadaZnuxKgPQ0yrJpj5C4eiRyelHlt8NJkA
I32SeM9WTAapkggBAYiHeKNz347aUIQnTCQACXgHcAUb7waBa04ViyYfzK/Rf5Dd
3GImCaIe6ok3tNxo273omksUg9WDOUe19WjS3EwfbPQElpJrLMjXpiiPsfU3ZqO/
s9kWiHhiunJA+yqTJ+jQ7bpOJZ0mUoPOYmQ551AwLJEgMV915ZX5k64VCY/dd//Q
tqzHMn4sb/6pGjsrdWVkKWlF5imJv9Cq3pdZTJPzZgXrede4TNZdMY+u9vuX8lLw
D9lPrWri2Mphfb0AYU8aLLu5Vs27vBFyxgQYl6K03Us48XuI68w9NqQ5kof2st17
wpvUNUbZOWGbQIvvnWIGLI8pLu589P9v4aYl22T/94JvscDb31CqI0KJiL0hqnf/
pqWc+DnMzkg6ww4obIwru47lBI7yFNFhT7BW8sCUgarzwNoTjcvGoUaOetf5aCa0
z9SfTPoL8M5SgvI4hSPZTZxFZYAC8W8u30tXYgvsHgLFHxjAx4WGxuijWPrao+fG
IWG40B2rxTGK/tZftSD7fGTH5P5qOh8WdPyUwjkdC6eqfC1Cq9JOyfgP+hxlGSYi
9J1P6ELJdex7TzId5+k30TBV/0hs6cvTM0C7fDCN0lyZPkNkMDdRE/ZDAYXKyhHo
rEBdJcBc2S6RHpDuXMH+whKNq2zQKj/S7UA6BNLn8uqtU2xx93HZ+q+dfW1hfwnj
MLCUp1+4T9gXnLRnJCyMIPev2l2h/Db6HhBt0yPZOBw3yNwS90Rc9Y/+G+DM+423
QnA9mLmkzKZ7z6GNJ7d45sWIyzTJSXUcEXu1uoomfuY3xj2WwmnqjNemaMZlRoir
+5yUTVzMr56iqv38AK1FM+tIbGfGwK3PTyBsqsfwkaxd8IVnnvz0gTrEkNTsGIs9
wWbQr+UCnBb1Nb4ToikTrPlzRxOLoKAf9KHyxglJZ0TRvJASl4gsV1aRLEwIptPz
vB36J+V1pgWO08rkhr7uc9og8fAl6wSaUzLoQhyyRHLOH3WzG2VrKwtLXW54pGva
vQmDFKe7smaAO5T3RcnizKwf3N2p/CmWGyrLgiEkH60YH+U7C7wEoVHk5/DHFoaC
ehW8hB2H0LiNNgvTCYbZeIGIQH8ok87RonQ5A/YSkh4UUZnvh9aMqtjLwZUYQMa7
VEi0gKQVKEetj/aVh6CFJQg2zPuoaHROb7htzJGzHvT6Ev1r9orB4xjRCu/iwGbj
yAY2iAazheQqQxwRTykKOlgRc+aN8A9YDmzy53rDane0b2kX/EKeg3z5QCpn55n4
rgLNrztm9u5/b4Ex42jEMOgbigLu1ujEY3kD/x6GuW5hq0hnCche9fGdepZ3H0ZS
YmiQkLOpcq/6dQyZjw/uBAOSNeMDvkiOItBVJT8s11RJELgZ/52/LjdQstgKVJ1U
BAUrRGzKdR/x+R+qbco4AWRqHVnpVMz4G0pqqvbqWhdSwPYfYukx0e2RizKZfTxQ
kiK969QolG05Urd1hVMuMFCkHZJvRmUB2NK3XtmNTBtjYS2wwjeq5IDz4E2l0sZX
eGUA50vtvVaifcFZn1zUv78UULkBJULv1EHfkQUlkLgRxVW9bywViR15HYT9KlYf
yFI8ytoT2jqvHwjfq/KwGWmgXaZoU0MYyEteg1bcPaHbTM0Fv2zcQi6Rpq4LAI+t
qLaz7VST60LVsTgPta2qVDA1l3OSLmQEU3aOmkfM1xN0mPl0qETUtbYwrzuL85UC
HlN/fc4/hx+br/d6iwOrttLGvvvRd6tYonlYZYTmx8TIoOP/kyF2xG448njTsIwD
xTIEPpRFwYNnR9WqBNRgrfwaZBW4AxH3Aejmi7xjvoj1DAbHGFQMhVeImR27hMSD
Wxpih6PwU7GAFKnL4x/D4mMz0OKSQZKayG14izhxq2G9CuGbxjhqxLYVaP45FAjn
ceuMoYYJSjUNBXOXJWIYxEVOZd4z/eTgMvCovMFeh1RkZBaP3pOhYerer9/Rc2u2
Ce7a1Pf74IoWRnyn8dhC2J+/x090kL42I+VbvUbe0DvpylDBI2spZMxeGfQ7WZxW
P1bpQIi96VDirbIhABBGbQhVqowld80W3HrVkodp+6HoKn5pMzFvuZfAdTQ/hRx1
S/aKT/vtf1+zEFQgUiLQzCeO8KyO5QLs6eE6iAY+FbLU0jSac5oLCfhqdhpGBqp2
3KIao7arcrDs6uL0Ke6RVKz8ZSnvH+N3+cG6ExYb5ElHExTw2GfRPHuXqY4pxgXm
E18a4KcpyjQnkrN3WN4Mc5hoPhW6kBe+zIUG1LjTmsVxiEhJkGCN2teaTMFVqM69
YsYGjxnB/16UEv4RHpA/gd6P5DobEM0B8vHScLg0WJITyQlHQsZhHIKl0yZ5gxIZ
BEAUm8QQRkYpB5H1zoArYzQAJaZVgMMo8VAiA2Fii9OdPAvViR+q2IUVwTATcsUt
KjhAI1sYKMjiCzF7W1zUPIJJXeJ8FzAOX6MXHtmlhYoM0qplhkuKhg/GhcWLx8fi
uVKGm7VDSjBvrcp1WyI6weMzDJ0cflE0CHj9v5Ve6MGYMrDZT3A9nDXuXj3Jhpkk
Tov5NulteAKRGJmf+si/PRZQwIqj/8PyRc6R43u/R2tCQR8mLe/hAvLNw7IaQKBn
Jz8eAz8Crgm7IEy78z6XDQzecGdTyUrtoqsXjTkbut5+9WplucdWWWI8NoUI24Os
deLrYmEU/6ID4QPkYFdrO+eBco08UWOFWBqNpxvyrjpcEtUS0A23j1OjFSDEi5Dw
bUc4CLM65/rXuzX/7KeSk+8KwmWrYd1D+oOvPBz7CQmbowX9rJige5IgR73FV/iq
KxMLbiygGw8KCg3F5DoyajUUm94a4ze+/PEkX4Dkt1fPX7JUwUsGzgCvACCOBFKn
Hjez3U5sHQ/glfixfiOj/NaKvSYMgUa5zVUifJFsdp0YN7dPy56N5549lGXsJFdb
WhwtR3+HVRupCtAJ0CFVwfXGqmNAx4InkUmfHXRPdi/QxC4Dp96Dzc7ZmNgLN3K+
Uj2YK0ftUZgw1ELc2LYBdj4CrMwBdIRcM3AyK/YtO//ENREeqYNFJu56n8amPYqJ
YcOj3CVOkMl0eqFcCcE0GbOIIq3D4joXsecWRWm3st4hmBGqEKtmzxqd+zfpB41I
iV1yaVhj+Wvuyk1zbKjF0dpk9yYTG+N/Mul7btcCGilwVHyjyMhpNXeRUsTgZY4T
nbmUzcXZ5Bp8bWHdwcQz4f4EPebJUsZWHGeeutKCpFZxPnOP4n01RBIpObIHjgtL
WJiGshrZypQZrMH5Bj6gSHQdoaZ7CYrHgEDS1q9XaIF8F/JQNup02JoGRgAQUm6C
cwek11i8KnNL4JHfY4hy9lN6xs8bVqD2bAAzsMQwD8GfQbFx7KyO1nSSh+FSiOHc
1i/5jvARpH5nd3Xs3sIsHhfJ9+ENlju/1HPbrmv9tKLQVkePZ4dF+3nYQDY1zEl9
Y8nVTwGnH/LQ/YImGnxEtDHMNh0ewWGrHjna4+mMDIOMkKnumQFFtqIoSlvx4vEf
Xec4lVqd60krVDikcTAEy0pT/MSr9e8fz/3JQQULk8p/iqLCZpUi7O7Bfzjvsj2D
zEmMMqyQDRhe6vMTFmBJgF4iiVki58/7JPKkSMfmDwmMMrCZ1m5xsuzSxbgGVEzS
J5sj4TYUmZToUZARa3BFq1cHIyRuhd0ANzswLVasKe46izfyBSr8SZGOmScfr+dl
CpAMudg61iDgpgOtRlaMXh62KtSe5o6wG775WPvyT69E7r1Q4CckbVKT3tsur+z5
AJ4WX7ubIZhLCTJuNPt8BWKuMRV1Qnr6g1nnkW1SIiqQdxTz2J7JPFlrGNWoDHtz
2/qy693GwMu5phglkRrpO3P4ZslkKngo5VTkfKZaPg920B7XVGP5qPcFt/sFlok/
R3VgzDwdxBqxuEKc2KlB5B0p465B3es0kCSvd0ukb4BVZLPDkThIu0ECBAXt6tFX
ogVVOwl/EPYBUBMnY+F5mMOfYzhOw2ywpucKupxpYATVzNwILiD9oEINuMRm9v/4
5P55z4Wa9VnYJjvcxCba9tFXlsqfjcW8OhaXF3c1txG+yrw5oSrO/rI9HeDqIhE7
mfo/cxc+UtPh7RSaUXgIHUHbmDhTqqIuFil6RY+7A1O3Tb5EA5/I1OcbmIBPeFoT
hdQV/tRUKensqH1X+v0MztT1k/UDQoqUeAXnnVa+AaDfnxLHLqWtc5UX2sa2mdRG
mCEltG+/Y3nYAkaTlmym4Hb28RhEKx6wEjVFilloCPJfpC1q2kL5hC9qe63pAX6U
Lk1n+JOljSf4UdENWhbeOoiIA73Oh6qdCA8CutEFH8w0jacSFt56/epXSYRXaBGL
i92oNHk2AOjQ+Za8bRAdGFowSa//NMEvU1y0rdoFU25C9K9E2CZ76WR992qmA7P6
0U3uxeOH5L/D6s04B3oXrkOGOLUHWvEiGniTGWC/G+mRiYgIpLYtsbH5lCzLbwrq
Hpl49rMWJxqzjlTD8oh8JycuLkhqQ5iVr+lIGiEZnyUcdFxgs4SGjspluL3biIRT
nUrSoIJ0ZmRcnx1ip2cw81zo+hKcT0DgygQxfBa8BDU07SrpNKGanTw35pbjP20f
f19PAKGzv9rAZwdyPhLezCmo6T2KbOvFdyEqRifm2iv1TYrOe0p8kaK6LS4eon7I
/bUMxUJgd6PUGih2St0PyPtIsvbYMYVfl45mEdItmWFaAdLSG/u09i7B5PF509tK
QGxTRlyZopl91fcx3FT+V0QkwlzqgZnUAhR/sPlVdZ9agSu8l3/MbmzQ1PuAGc1q
zfmCCiDTifO/VcLC7kcY/WbrPzfKE299FkbCr9DBEvPaHE2d5Y5adYDiAVn/cy44
muPASXT+z8l6+acVsmXtmTG+75IlvJ3YGUxSeWkDnJP53dUyCVoPnirrsQmdQA5n
H+dkzlMbIlm/XX2JjgB7UrmcxDFqASPvuMm7pgWr7k15p2UnGgdTSWFmAjlWcIJb
HZhxkXok6kN2r0tu5n+cqmMF4VTflyeo8hitubnO1XP20Bk4kjF+TTgXHhou3Dks
ThjQUQeqkQnsdsjI6dLnkMxct0d3n6BqoE6d+K7sqRvMX8Rf5lnWpBLk4KfU29tp
wUdK04OrAx05CP/8oRh6CLhRjMBfMI3A0JIYub1OypEFRq7Kxh0QpPf2eSj1Q5rP
3rSuos7HSB5MSbmQIyEOuBew7c59SCdhSZL3ghoecAZ4CG7/kdHwFKHjlqA0PGQv
LSryB5IqJGSvGOkTJls8NQs/xIoLhRFCLCxffHJwQ9RAiR2OZ7KmhjV9S+f/j3IF
QfTg7gH/cW6C+RvAV9gKhB3wavSpdRGJCvg9yk06xYS88+wXnpFI5AI/t7gdp4ro
mWDI764fXRZ/X6sSyWQFqlmcOVbgbvfCoiRr49+dK3uOgUKdPL9De4+7avnYoKTs
T0BY2/XRXZA8l7daNncJQz8aBvYVrRZbXpLNRJOEFI/7XfYx3vXqvHlkF1s2zyvk
bYhFD10XmoaPPg9JVd9kbeSgbdSi/TtXRLSko3Gw4xK7JJvRMFDWFGZ4YA85G+0t
lZm6mepVdUEyT2IeyPbB913f4D1YP/j8tEWJw7qCkI5eVP3+idKAW7Ygm5UHYkpL
salBtAjxf81lszW7icojLRiHg1WWnXWB0hY0bKB0vQ5cYgdxic//rgUQQcNPoh67
nOvf0JBYo8QTecj1w48UR+dR/9OaiqbVG9+ejCSQDOtNE898z+n+08RY5jODBpr0
FC2OhVmbFyXDuk7xNjgoMRIqyXc3SUHIvbFXXoL0ss5cG68ToQ7j467oq35Y3ZKq
IW7XP5P1EkPrgBxHO9Mu4G1kITRLBeiHumiX06vcMPDhSmqQlTSxTpf01VSSYs4c
eQJESDN0QvWEhad25OHIIdJ/qSzv9U+ngE2NncnJJ6kAvfHfhEnRP8QBOWw89IEn
dIWV6RZz8chIWD2WA2qO0Rs7nVRUbHpw9ZpFwajHqAq2+sh2u1hqPRzsCoYfOx0j
xEwdFKMYN1fsEPvHOnp/nJedx+P/ota12FT07td6FUuEkZav3BtTglm1XPTNcT8n
mU1ZN9RMlyQQjkEcZHhZfVTiK6Apj4HU1ZAuO10LY9SW4DhjaiuL7iGlkaBk5OUH
w4nESAzk2zx68qdz/XOAqSCmUj+MwyaEYmndBRDLAZN85LHi0AN0IIqjPEcQZuvC
tDyllBT1BSijM6Jl7sCKVeK0NAihFvXwxQsg4aAFN8M+XHtz4PphhnFE1pzLhRO9
eQVipTykoymf0T0F52Ejcxz6VpB3z8A8dotd7z66XBcCgGWnJldTD1XG5Jc7kmY0
mY2EsLQsHcxSLt4K1rpfXjA6hvjryMSV1g+H93Ac34mHNNX50R5D6+oOz5u5TgBH
eHpk/BxjFrWJ/C2uECyjCxBGERIBJEmNX5lzULIR4F5zxgkt890pNfcBTwSxNlz1
6wYY6ZsP6NmlCIhuwWBjZRkqtl/uu/8X7BcLyjOW0v+GouSz/sWF0mcRYQuEoMZI
P1uVEbyN6lEYw2vgPEWEnjiHfahfx3eKAuVKyxFOTX+mMltyp7bNZ6lx6UbW7Fdc
sA8mGTn0KO/b4w1zssYJDAnw+RPu5V884QnMdqsmq5OzvIGlo9YIX6Hb2Vkt2XhS
syFleKk7upCvSkSMtSjHrivQdczLWO7pE+R3m36/M7qTRCfHE2WVxGAXjz7+Dl9c
+7a/xK/riX/31LfDK9UAF1B3+g6hQaJVwyTdCFwShZg5tXkId/igx62H9FooFdo4
uE59b+KWdUM3slaV7PVyR7yM9WGRYP6emnuMOApF2ZySrfIlGoJLuqNQ8et40NCQ
As1BborPRNjpFqpVe1lxBbJEZR+jjZOKKNv2aSisTA/hfBWP88Kt0cnjnHDnQAsr
K4reJDW8z/XbCop7NWFAS1J3prFRETsfKe3F+4WLy5C4HgEwS14Ge0hCMx3wSPtB
DTNgX1aAPxBJ0EGId3AM3q+rB9+xoBqQGEO0iUwxfsc1wXXCMFDojs4Bx6aU4dSg
AdmmgCJ+B7EE2tdBdgjLeIPd1PoVtfC5mgYvI6GuEG+w72NwK3SEH2JKoi/JKzuh
yGNywBNM8j+XynKt8+EcAGLlwf6advFBmCGHlNSBjjTx+VRp3Y+irp9/zQ0qThJy
s1m35Bj8Wth47h7CuQczjwx95exrfWp+5e3783l6qdgHJCmgnRYiSTlHBu+OFuvX
J94X6XUQOozFO1YoU4Rhce9Pwv/XGdJs9TalV0mUnUUi4IUVtBe0M7c0I5MoH2qg
cnZUfpHLtT0gJWcYUDudFFRF0z+gk31LVYeETCN44CqmPFIPvk+63JN8E02vK66z
9aAOAKT1kpA9UcqTlLE6exEeaxn0lTIxtVJMjrkiTVjoYau+61xpqf1HQVDF0PXE
6aAdYSHdAskm7vWAQIxSajT2xRCc9yXedYdUJuPaWk6G57R0A1mVySgBcpL9EdsA
o1BwZZUQMIXSh443VmjHKOT9FiiK2S6r4UmNRjawFqFcjNzdfjB0Nc/nIa+6vT5H
D4ZkCTm8HsDEvzBRp/sKZDrVan3x75DWaJHjAU2Xprj6c2pCgwZ64+lMJs6wDRJL
CAAfk9MtOtOhI7DoYnBsxUN6OWbXp2IJ9nA7OxXA7oNIi+QHYaUYCZnqF1qAvBdN
ZPPqQF4beU9Q9VR0VEmRGREiDXzjKvqqbMznl/hUiSARbLxS6cby48g3ZZTjo8Z/
wnDWdY633tnxLRz1ikiTOwyew3b2tdTu4aeHTCMgEJyk5mrvwP639bbPVBOnOO0D
I9GCcmVPT7BwMI7nTxtBAS6OJzkpnEj27SeoP1WQMHWqDSI/AXb7OxwSoGajs80s
3rT/z8WUUmFywaBV/R+vq3TxEJd/WbNH9YNSeRd3+osbzhZ7ivBUp2Im+0t7Fkyq
6x3hULnmqsQ8ahawXj7QeCYBnncpXqCxfdCZfGFsu9kZWlUPPqh5+DzDEuU3Jgs5
GfBavJbadoHz75upNJGWmcrMm0PGPhBCTQfMPJD/jGGGMQPdly843xJSYE5vnWNB
hxswTKCX7cdEZjBunbHtgKVijHAbLcqnsHuA8ES5/fi0UTgVsLN+okNajgJ/620I
0kzyB2k4V3JWP1BmqyZppxZxeZpN5v2bOsGwCS+BLOPIflOYrRejCj27DAsYqJ/E
UMo6cT2SjtqZ+YhAp1PGyDqBRfwtJPanFK/cdhS8mHB13Gc553G8UvgbUb58B+Er
nOkWXepzv6CT9sCR+34DiCtsRvCVkaypZHixCWZ9ErjyRxKK7ZqkKee9DiTmzVfR
zXvz9RNe7LVJtDIotkq+pGMIZV9PCa4etdL1moVU+Ztm2tifKsXhYq3SvOBvNJuv
pQttm1TcAXl0FxRJpaQH0eyO6cXdGY+0gR4iatFNuqjnHBcfxhE8NzKgAe8ob/50
9U46Ik8XsA4ttMdvT0VG9fT96ilbSYua4WUirpHMck85snNTGkRZaRWyC4ftATqb
gUaQJPgTV6V8OJ6TNZlb7iK20v3bWSTtjkfVOsnrVW4Rq1Dteq0XD2F1tvDZRXxG
JVcD4thGd3X3Fo6Xy52KhO7TN36kE6HfXLVlVU6wHzuXGsBAGdc9t2Ov9bDQ5Gpr
CPpTuGT/V4a4sg3UTnLK+uOFNZqwbFSDZV+JnYtrnjIYBCdmbmTKCo9ExDckHEsl
yUW7TtMgyKcUcFe0Ri9vuA/xz1P2iTxdEIvIy7jWbujX5N0A/6Pi9qws3aoQDvX/
vo7xBraIrEexkGfEDbnXItofgs7dE9l5KEl63AUEibL4DKJbAc7BLlLGRQY8tVPG
NDAxLeE2eqE2JgU926BszAoLqQO1muAxmZ9NAGf1S2GMHM1qaOVmik6Paw1hOiMP
3Tm+UkZMsSuoEbdAyeShaBFy7X664cngDWUDeordamh9PSg1Q0p0TrCLecLS0PrU
6bQLzTxRX/F9fTbGgf0LWAcqWUzrzKn8rcfY1zW9pBK2+2A3qNc06crEmhwNAooN
IJFjRKwwASkNlqqodWQeXvgJyXyVP9Mj9nRr41GMVXLzIkJO9yt4ncNm55UYCUOm
AiO70eMkXKVoPWzIpXysQTFmUJ1X2UowMLTmKXBBYx//iPWpkgzpooFgxOiFuC6s
xvVuJMPHRM1KaYieCmhW0lgeLL02O6KrECV1/kc2e0u6N0IcJ9/PtrLbmzpGx6RJ
w0nYlGFiV5gP3MBrmBi0agXrCWpG/2irDPaVFqa0Bkg6pQTdgRiiGlYnKUGPJWvV
e+Z3w/Pg7GQGeknzLtBS5sTAQJsMLg2Au0yqmPE+PP1UuipQK9ujhExj6p2vKHbb
9HSJGzmnOpyMkd3dH/9k7mJS+EQEYifCWDIQjGh03CcUkIWG7bHJXF4ECSMsY20h
/NG5hhCr913CtwwOMicD/QgxiaXFMvHl3LZRZZQbS0BZ1bKXLghbinvxFWQjq1Yw
fRWgQ1odzlCE3C38wNSGcHsr6DpMAwnf1eyXE71DckRlkOR78V8+tThMaAX7HCF0
QWCjpqHoBYOcn2BTgnjYVg8dWGqM9Br0pKefrLT/9PxpiWbOCr4jL/BoKkRzBg/Q
Bf/vtwDX4yb3imtyqMLsXbgZ1fpImJzPBChBGZCk76OlqviVkRyhelmhSoRE7saW
kM/sZ3+jCc54pjmChElYgJzjU6ZavevILRlfrNHT8K7mngmgdnCK9/rKe8shcdP8
T0qBZBtEOtTXPT+p4Vue3nfOSYlqpBlejdjAhZ6Nly/Xi7iSTWVG0fcISdIP9YzM
4UBa9nzwO2J3otelCLs+pvMMMXC38QhoerFSGfHGoGAxSDCcDWymfilrB23i6xM6
q+JsTH+9PIA0VVUkUsaiJfNirE4RxjPOCrhdh3x6D9xNkCBFfW+x+nXgsVVJE9RU
5Dr77exniGWSvMBzpWUXcUnFkRDqDLa60ZwUNbyVksNlCOd91saZe5l8pJmqdvPP
asCiefJ8G0tsjrvfjy2uu0pyqV9XQ44ux5HVI+SOwgVBJGBUd3PzCeCV6gwvYZvN
ixIIN+TE861f6hElFn4l0skl0HCMVoJXedNb0VLBixDaRMJ3vIKY4nLFGOY1rgrH
9b2npXz8mFwXl4V4UtI82CZ1Kyk9bFRX7BRAjWF6zVzhV/o2vMvMgxWB+zJKvJHm
kFmQ4zhkua6hCSjn1GzJdZUebT4OH/oFEcLNw7oY4Sfmj+jh9JdVP787CPAMMuV9
lnN+n5VNjnqJEzs6zShikymheZ7+YeLT4Cf1f0EYeJqDR99GZFJauRMjC93QrUmh
lJtcuZ7kV9FGSY1Cx/dKt4v5F2H1qIw2owNht0BpZwzDWgpB53mgNmT/zgyQQ/L5
3nh9Re4vphjMHtL602fVwNj2twagmgnHtjfwQSiDRyefG+dPpAHV6MfxK3NwM5yB
xUqPLni2TNmGLeMNd8t8ZOwLGkClHQ7s5VPhcKmwBNCpRoCNmPedu9370Gd8ukF8
CAgi7Egdf1ZgX1rX1GM2jJELf16P+dpUCsSbazEYOsXf2cKDJTuGg0MlyMHM9urn
PeLhwDQdfia7O4ltSO8kvp891WsmKQ1JFTkahZBWwW//oaoDCL30X9CSBInRPyCa
xWj6knYReUTqj4cuZ5RqtWWZ5L8uOov1tzELMFkP+eJg8KE5DLBePvR1hiGgxU2s
H45I+OlZKYsgG4Pe1nELU9Wb97zacWnzTAVxMc8lSs8TgLqLJvQ8WzFEv9/LrCzu
kcK76wnIBCs3J0ZOYoXDgOJYQp+8GluD/wkBkVjXo2fmIr/PDxgElqmO5Or6IwRu
1+/S5X2HlsMviJZuO5tJiXMZIJFhtW4dBwS4nlRjp1N0/GmhqXZYwmtJw+DgHlk/
wYyR+a7DfoQ56To6cvqf0HCt8X669U6u869LaX4aYqWq8jsspmOb8ZJ54K+qG189
tDSedU0iW6PIHktwIb3GJJ2kDeBDDvZT2jbqycN6Gz5H2tV3q1va2YVozPHWXgDj
zfD6ypEZM2bCUNFo94k2v/9mY0hIIK7wIdaXPNAGWOL+0MQlLmIhAeMNsyOKtcei
ff01E0RaL9EqSbw8kSd9vFCAU/y9tQY0BJxR+rsExCwHDkfNwB6u2L4n47EwcB3K
SnZVPRcS61ynO+IefBZiXe+irJdal5E98u6cPygUyTjrMycbWQLf0iSVSf9ZogfT
kZCIw/+n473yv8sSaVbFQxxEEippjAwlOusHmO3EPpw1ULNUGQ22tSMzJa5EVqBs
124scRmAMZh/RZf/yMBM1dHbOVUH+l5os+ileTjV8Ul6FLw+RPFpRnxv80PRwR1x
C1BQsqMtMwxBNnQ46412WfLKsHWJPZS8CJ74BQ6SzpgrSCn3nXSrfndmFKXS0+pK
bEXj8+84g1Rt4nurqXjeyHDAT9fDfAI320vm78ltwVIUwb4ou3ug27i0R/q6ZMgU
XfAl78LRNuTzwAcFpG0vk1a5P7tBCTTwDYQ//R2/RrQy120J47bwDZ7SKxJgTqhZ
WN4YNL4KMJM7Wv5iRJ16DqbrixgdUx9suADLHGRyM7SJ0E+zJwHSCFmi9h80yLt4
SmMxvb1dR/kqAEi6lk2Mt7AivizbxRMvE49UH8gzQODEFIcKHL2DYdOJSXEGOjlu
lu6cAJzR/uZJ2e8zvAozAm0XudPspnrYnfwjhBTr9RV4/RWZzUt4UxdIs8F+ZPwA
m+zgIi6dpY8vQOH1Nhx/TYsu305/Q9RDp54CveWj9VpYZxhdV2w1FGZ5ftXj9sCl
Qne7Z4XbRBVUu4f9P0LyjicX55CwFiVTcK7+my8vDzv1MuN6GtsPxcHOpdp+pjbB
X0yxzN3F9P7EUoIc9rrfQ1uxTfcr17GGM//gGLhldlFmeSVa6fkPzeWCeMm0mB+0
goR2zhI2SveLd5jNmSqm91zb606qZyxvBPdqalZ8HFJ2f3jo1/d4eWAQFPVwLgoe
dvyYXUiFsNFGKewAC9f5JRouID4RZTNOkQGgT5usoIIA0C9o9hwpQXv29UAHx5Cp
ohMx/qAgo2ZOEpZXzciuD3ka6fsyk4u+AtmGFhtB6RTwdWsydUU+zBR/iLtpy1jH
bNTOZk952ReB8NJyeGmgOfVrpitNfULBkS5KCNnjPImZfXLoftQHjwN3l0v8TuqR
890X3yavpZFjVc8Hjv3I4u++ZLDqJjBkNrKqGqTynA6SLiItnRpnXN6+kpzXXsvk
GtHd0YZ8+kQPSYADwglkoYdd1trAk7Ex8IOL7Bx2Ayr9QvrI4lXDUtE3z14s9gH9
UJEByXn/1Vc+fNaJaXA2YmLmwPRa8GrYhSM+xVhWqpB9s+OCqJU+p+NpkBmuypAN
1tf0PdPRXUoNvaEzEt7l2QYu827Zmxj69RLx46nnKfUgJshq8BMDAcI0DiU9xUwA
j57jGcza6mVxgcC/ayaat99p6XbtdTypSH2ki1egDpnH+WxRsyr8Kp5QUr2/ldv3
6CBtQebPlSb4bivq3MtkN4zVAVnreS0pWAyP1OlfdfOwXiKUU5W7SxKPohYXyeON
MUOa0DWMTjaHcs1n7CyEUSyc89HM12da+s9oclFDvLuOHytXVfE5HpNieJ22Ub7u
a8SRDtI21r3U1N2NhdURGM62SvBwtjUKguXxY07EvA5bGLnP4lvFrE0j1dYLKt4M
nDukEOvlkA2BVfHcsLgMA390PWQ6sv4H86tQ0fsZk7fk9GlDRp+ddVBK021PkoFz
DHksBxSxaX2haQTK3vKHmFVlv6dghIBoa9Fhn2YadfKSkeYm3IFIngG//gJhz4Lz
lt7z/5u7BtjuxGugZGBxJH7a9cLyYCIhnh85gshvCx2FYZ0ICJk7oTRh/J0dILZM
QPEMT9AlRs7bm8DbVA5Ah0BHhdVs+niT99fuk/c9+FA2Zb6D4fV8DCt0aqj2FGFr
IpFKZs8EpH5dpHUGenZSJ/HJKijva/skUuo/pu0Y9JblOXJO0cQZA4mTxkQKF1+E
QeymLGLKW7X/Ofybokw2/QY10C1dWje8QpjahG3/uC6HY9kAHp5AaX2/sH4/eIPw
qae0O9MxHSKTAzcc3z5h9U1XkV7UcPHfxd7aB4NCQj40UYz569zGWfCaQ+C55myK
t1VY663lQwMctkfYIoMoL0AMHAmt6fZqOdM6bikqal3Zd4GByxuPhQpAeG/7kJDg
H3PsVMRXQgGgPg/HMhq6Tn5hxM2m7nlDn8VxuX5FU2OyROq/+0XQCyL8P/edmiLs
aDQndUFZIHICjJs51CY9ayaff92k1kryKeQvK3K61pGKyYNO4Ljw41w5DlSrYk4P
wPhJFSOknKqaTt+UwVoXdubLMYxY6D9olNYxLNhwyUpiVDL4WS25thQeNhnT+mlH
Kh4wMp0ppLxjOJyNGz1y3oIgImN8b5a88lwcYy82HCqDqaOhduoKM6SQQiausdyJ
PE6LS8jfqPpzXXxrqPs+hvAVl/llChYWS42eLN4j6shkhnK0+3H27FUkoonbhuL8
gxPBk9pfLeXC31DAptGuUkX79pVbq0pOIAQ/FxJcD3tQtXRETUNfIgqKquB649KV
HdaC4XmILR/Tkas4n9IGclplAtnN1k6Zy8xZ6FaZaDxn4GKRlvuHP+q6mchK55Hh
f0/N5R9v4jN/4erOR02CkUBMO366FYBNxswTYGbpKgNmbOWjcEF+EPdwLEGBklkz
tauy0PFWQEG762gI4b/TmkRz+MYve8H5x4sk5Yk2jC4oHeAYutg8lSNfMndwlsb9
BpPiD2kC92XnyOysc9xTmPVieNQQXn7rWrbhclUvW1jHZwj833k+NElvEwOBn6YJ
4kqpduXIH4Q/mkR9nwkD0C8Enf0muyhvXZPXdAMcn/lnI5R7kFVYotOMw7kRHgIs
71XKNaBm6JDij6FD5rvKTfH2YiTw+97fkgIbwr69+j1JOt022MXSMPB8n22QrbJv
L9ReorYOFdxA7HH8xpNnSgdOnL2tX+4zymbEKdcEyyjYUgJI5TE6XOhZWFXHsBNe
1PYPRPjwIrpoBF8aT9qT/3gWz8PnBbsURfus4d2WQnKcBxBfcEfbBCikREQvKIvm
uFygnxWpmR0ZHELQ33rf4qGJ8tHIeXa42OwEq97hBRNFrkuhriuJ5lTjrLqskRxt
4lpNqzu6pA8qW/S07yai9DXVplKC+XppZ49u6IKBxhxQC4KZcDJySUWP3g8nD3B4
nHiuTXaPd0Cx7kFvrRDTX2WbqPCnjkdU5ln+sEMPwuIJvzYunewIEI/NcV5wsIhH
FfdvwUiCjWKvonobaXz1inRSXHluQkCeM/Obh4qqNoo2vrK0DK6dJoDkN+CAE4C/
dX4UrK+RpqASO5+SJAqx4vWpQ32mHmlNTaJRuMZSoXv09Q+TcVe0rx4r952nONJN
PqPZ9VHsltKDKx2qzeekLJtqj38fTWlZYLcGS/55Z2SMicI9v9Zq+dZ65fPb4p1I
Mx4DLBaEs/tmh1gZvxU83lHpoghwhvL84ITFRsu81wpx98sfCtiDuf5YieTHkvLh
q6Rc8/jgPY1mGDP/9Uz0XZGC4aY/ne77YrtBj3fntbWKdg/MbSVGTeDX+5lb4i4m
/A/wb4wi6rJJz2gxhg2UkxPZvQMXTf4/fNc4slaU66JuD8T2G42LZ/120Tau+8Sm
7gMsPlnmBhi+U87YnmaP4FZcy+hjgDbOpvPOCWx5FsQ7ifHdqQheSfmEX8fcJfCt
j9LMFD1bkpY53zdrWk0ZrXM0goOxCKeyXBY4A7tMHiLtPBgZVJhGsY/YhGfSnyyU
Xq5MYamnrhThBTnEis5tHuVCEuHz8MJptvPh4LP4xoqLz+YWqxRQdEi7G7BGhZWr
AluAqElD/AvnIb+j73cnFOHGZhnJncPFuhC43YcHc8bVvsFhdonQXyhvC7kIqjdS
5DzB74+bA6nZ/Y+47AHSjFadUKgx5xUYnZF4sENNsc95bo7q1rkq9iT2XUn81ly+
I0CdC3tsgbtHj96vqD+M+PL6h6d5s5pyc9JsMU28I2Yef7qrI9pdWTYAW+VOIyZW
i24YauVLIOGM49h7t84M6Zeyp6lji1/HZFBuZgT95dQFX1sTSgBH2JzcFNF2WCku
06gNbjkc9IyGvGM/EmB1og8PbO+TWFUXTZvFGC6+rgulV4nigcfTi8y/WGTB9fKF
n52uT3pbeI5s7P1NIwO5mEPPQh4+lPM12QwB1cAAXIT20+l4vJYJ0Qn4iAxVMT6B
ZfWVcBEHenUIkzQNgaaBErrLXRF/NE/CoIorqNRbXtPypPVgkjQFsuxyGxpGKF+C
GVO0IB1gErGapJU8SJdJEY7GQjFu1YxTNuO/Ehpi/UM4AJudkEjjwj7J/yoHgqvd
FH4mhsCujJcjlari29/ZYmIQv+OzVddz5+WlJQJtxhHnx9pJHhUAjSFa85Ng92Mq
j0Gs9tmimK5P0n6MH/qW/1MfwHF5Fpm8j6QvTvk1Zt0ORVgf7V6DuN/ofxaTMkiR
P3ucqfYe51fCiq436Rz8VWCVyGElEgiOdp2ZzfxMArw57SPU9A5gINBzU0sjlbbe
Z09sCq8a+nxXBfOBTEVV3MaxlSxJwI53UfKD0uCZsXCRERpvprGYQv9QlMqJePuf
AZCfJRDRMmAORCaLBbIHHaJpfthT+cOQWVmtiPm1UKZcZqb7ZP8CiSxxYUsDH9W6
TD4egY1eDCjbrFimV1F9GG6o/9Tp3Q0lwiSDxj3h05gWwATXZfIxkzUJ4d/AjgD8
t3jPv3OE6mLNn0LR90V7YFmbqsHeTuyWv4j1TSB8yN3WXnFTUC7+Jtl2S6XHVgOF
R1+14T6oTKm9RMYUHHAW5pVzpzNxmVn1MYGYFE6J9T4jbdx5rufKlfPH3LRmmEPb
G81RfiwV9ji++/s85QKG5UjtWJh7eFjg8sJSA6oaT0cw5cMBkBBsfJsnsV3Ei2T4
p4EaKIDgy9lI9Mu/Gan5UgI1T/iAK1/usse4pLaIM7TyGO76D676QmkG7PLgVJf9
K6W7aomovLrJg/p8kHTtdzUuxeTSzd/upOvgFlFR9OoDyJIYIBZsRNL5zB+aOxf8
fLC7W5yCzqETkduNg0IRNrkVGXKM++9KbtknkSAbETg+Sbdr0C5ENp4M8wIczUL5
0OTIk2cbECJLifQjirIKtCXlb9Pfrm8ify6NgRPnpmewC4mdIk/3ZNhHBfXLKsEg
z8bZpSbOxrCGTFR4ZSbJFcQrvw13T2e9rMOJvO6GAQos9GebcAl+CRK7nSmj6T36
oV5sPtBu2rhw7m+eRLPeu4ENmfBq47ozX+29fGNfztzBkrjdq0fihrraHDNXiJE0
ynuhKQeGGY6MEpvYDZlS1vcXuqLUoVh3t26U66m1PMQ9+/Y+8dZNxMB1DHEu7Hb+
mycRF9wLJzUtQOYfzo/ZJKX6/AMWIQbMvL+Rs4azYpxQd2IdDJGi42BErGkPoeg/
LUunNrhdL4PcAX1SSy1a8vwAhiALOIwL1WWTpSGyYR6VbEiS6ZBfdSa+Rrm24H0D
9ITo2oIAB59QNk2nUrwW4MxlzAoK1eCVahih6TQmMegUZ7yVeXVlWF49rXpTBJNq
Z23s4PweUzbF692OUfo7Wd0gOy4Wb9c+k3AvEH496N0T6xHmIArDdC57lZtWHhMw
5F5H+fZQ6Ql+bgctPLS1nnyfZqabm+X4D0mtp86Hk1dd+Vh9Lo6RzD3pCaOi+rm0
hx6Ix9Pb2YYU0xSVN7d4sujbNs+J447UzTdFBCfF1EqndxYkZX7UlivjPWow3qzL
HXK2ZaWXAVnfBuPlWNheTtXTucEbNUqJ2yODri56UHUHyeIvNGJYl86ODH/CjJmF
lv26uPpYRrrTdv2w2xD3ct67is3lJ/VV6bx4jpnDEFnFPn3RXevhy8iazebIK5Lj
5M5rRAbFKkqsOEDsMH8JRySajzYklvdw2ZjZQPTm8BbNk5/PAsPct/7su4KFZGZl
Ur9/gOWy0Q9dYZaTfC1mMHcptxcfDrFc9vQlxfel1J/8h0NPQgb8EwRtlbPfwm8g
wX/UHnN0OyiVKVltjugSeyHAhZg+15Y2lh+1KxKklZkh2bI+t22U6hABXDwRpvpz
dTBJxKijMCNiQFwdVMLeVQn38unUSeBIsVPRqwDKZxxE1Nu6jEbKPq4vCzcuy458
rmbZJfj2KHIMbgLH/wfOmBrayBZLfgbJBz3/yJjMPuK4zBv+YZ2UsgnQ6RKKum7Z
Y9RzBC1nb+vUG0NSiECQiOqIRq7/gm6bD8I60W6HM6b8Ho046+6A2i8EqbokMAKk
CPBQ28XNKhmWVcf0P8+zqzCeL8PVHcHKb4VKoaH9NDw9qNiYK/tB73xyDjKRvgNN
TSYiECScZe7jdAzSvealPxx2Pn4O3sYrhCqNapN57URQ1QgtbwFY3fzSZ2pT/B6j
51V3QBWP0/FGeHZMPGp7tzBp82lvJ7Dz3PbCTxhBX9Odm/1aqJBwvUYTti3CB3Ra
bUoQmyZ+OZMTb21NG7ojAJHlhFeL69P37oSrsyWPwhfGhzlZ280tZ8vEDpvomPcf
SR96CPQl4iqkpFUZOn9feFF0sIyhxOEUmijbueePh0m49mN4bejSELuEGBANXQhm
gpGW6/c0XRmcGc735Or50//ZLZgKa9zskZV3qJ5FVHgahKW4ZQRYCa4ZwssihipP
/6zyprkTscNYCYmi599YSjtdeqVDUKhJunXLLyjePQFg/xySQD3CUlntAIBXZixR
Shm8mFxlA7x/ElisRrsYWKyIaIIttIlb3/GCKDmfWRpGGv7I0YXabxnYR6sHKtJB
kD7f6XEE3n8levHYu8gIQlUA3K0NYmSSbzw/mcdAR99SIhNax2L/5yy9bPjrzwLb
SygVJPWMzrOvqJaehVGrccBQxG7Tdde9kQeE7p4zu/ay2ll7gZNA4H8tAD9g+gmM
S37NdXSjsJYMEVUQReuj5B3UZGZacenYLiJ0GrzzJT/2GO5lrql+0yLXQcAD2sMr
qZ5gW1TBQzA+fGpdSCdqbU15OzCoKb4kESV5IeFgacwbqBwHeBdk0tA4Fz/OhF9n
T8FJAMj8NMOjOq9TbnwnTSXdqEFqhlbzw7YoS2jMymkvVKpThzQxOmxbZhAzehtr
PLgxeSbzshJk+S1VTS6250vXr0HShBpVI9Kp9uXML6Nr2t3sUGtZgxDTYM8JgXii
hAf7zo3JmYgKpEQ3xmQP386nMk0XQiHMUsrF9BCMBQmJ+ImI9V7NB7y5NPmPQiii
9ujwLj/Ffie3fOcT4PP81xVsxz2zLqayHRwyiiNorRXVAJx3Y6otNWwmEDlsoTup
Sk5im+S93rZ3xpswv0OBxj3vU4r8LTpEKm7Gbd5XoGgsRaXSvkNp7Ef8ty106qhF
Hh9hft3ikHUibmKWIVKAuNArHOGtJ2XQFuzhva0x07Oeez7lEMEXeApGfkgM7r6q
5GYQgRH4zaZd9nb6sbu653xokj3ZlC6mieLWOpwmhRA3SsiADPGCDzh4o6c0ON29
zKfgY/lGuL08c6+GwfVhZGInfN3YaXMOCNJMDZwWgILL4sg7p42RtuUoleUShU9g
9D3vy0k/knxWuJoEcckV/nBpXnvR6fqAuX120DAlCNGxwsFh8vULKLegQ8dVUStD
Yt2rllyibcl0sD+bY95jMgeCnCFVSSwFQQ9VWV90LDvYMKIEj5XisJg5y4BKA7dY
bkbSDeVjH3jO/72h+SdV55q5PXravIY70O3ppRZrPbeVQBYepTamtIQkxOcf1PaZ
5mTliVshpzuk+0pJ/dmjmxU3f8keIgEeGMf7/86e7Dtkw6wkw/S+/Tn6YJ/s3BpQ
97bd6QZIBoRvgEkj8V8KI3RvddBXmi//T12oGfBMZOy6urhgDuf5oT4UqKUWT3RS
ngaeAWq2zAaOyfXNTkwJml433aKqJRUUVy95kWiPftYD7sK8QJSSUh2X5ixAGAm9
OU0/EeXqBaEspcMbS+ZN4YJRGfsDwI9vx7VuxOz0Xhc9uAsqmJ0NlNx8GwDxJahz
NHy5xw6jycTHCFlX2RnGySXJGgXO4Q0xsiDcSX3Oy3Q4yf7yOC0N6nmr0GZEarVR
8Lgb/wRjcJEQ4DdjB0YYNye3SPITad1iliHJAg1Lo8YdtFO/ooaQ1y2F6Fvj0yXg
RJvzCjm/bQS+V7IJ1UR1ldC6dy0sd2TEAWD9ufhC6mzL/urghnuMHfh8sZCr0ghx
pYpP4Pn0pkcVO8mtokEpAWFXRs0MtatM1nYINqiHGgtMfeWaW6h0+2SGYRFC3Qyg
dBku5FI1gVbb2ZP+x8K6PTcIXhgablPUfcmt1ZUTga76+sMyazwibHKbHjtCLp4C
kZ2T2Rs/glLt6RNp3LSyqodYmUYmI28vw1qc7I25PIbgwE0dm8U0ln/laps6uMua
gbr/qzGyAafN+J7CwYLJCK9N+DjMksaMVpbw5Oms1QVu9qadKBTUHduTSJmoHZkR
C6y7VXDHkCly8QrNJ1w6WVMItuzMKEjsl2nrJzJkcxVXjBg5l76QwO8Pte2kiZue
YgMELxMqAJI6gC1P/HKheTWPdEuBquwaumU5L01yI2oYB1ejVBdhU+Z/fdd+x3qn
BP1Z+ncMsTp/JN7XcnJP3ZRHRi5kMJ4nVMwhphHCabygdZk3QQdE+91hjiBykPaX
47+cgAKH8XUi8xs0wzVRUUuU0ZM8+Nw7xXIZCUWGeyB6AnWiT6TMkCh1pGkKBRSl
gS8ycgbKWfaHXkVAHyi0AdAU3u35ZgpfcnfLxSuxY7pqCOzwMWkwruQPkCf67vLv
g2iY0t22mQtmsI0ZH66Ooto1c5m66rgXk233O4uOPvcz8+vST2ggr61yy50qgg0u
dc4Otv8q4P/fIETlp28MkBwEjGGD5k+8SPTrZKHK0XuqjOvSANeyKvAGuPNyfJdo
Mdo0Pm1rJCuOuIWEL8q3jW2as40ryOZ1nPHT1KauSaGXONuprmhHIYqdDtPGf21K
jMwAg3zG6Slgc1sDCTE/sCJCWmnAAIFQ3lkYZvh4nLMWqJ4XOv7vndrYkIRGCaWt
SrNlJHmW64jWeESItbYyruO6WdRl4Cz4OH6nmbAfeZ3PuV69IFpguqeK3lRxXpLk
mTBW52cMRkuiCx1xeKKEB/eL1926TdXBCs8g2FUGhPLBRww9H9L0rVuEVCQsRpep
G7l/D1gUJz8yPFPuU0nIbASSGBEJWyguNFHjuz6bqJn0TxAfz+8FAFrthSPYfOQG
n1P/7UoQky79x5Hap5XxQTZIfnx+UCqOavYDS/UQ8khac75jzK22Mdqmbp0QXO50
tf46XCYrh53nXtpYalTyC56R4ZVMWYtGjK2nTINqUqRHJtpoa1LWt6gtxhJGNzXy
GfWc1V3hN0Y5o2vWYAIOAC2dN7BDz1MOlAtuDrH96P0jxMtLQASucLPoR+8MV4uf
t8V/inTQ27VRtByDRXJrOiYY2VvdMwdeVLI8SwVoSDcVeAa4t9OOCUVJdF1IC1zL
pO/lZ4F1kMFHQ/2HkhEwPHYUxWqo9+IPQPW+tEAgVTn8fZR+RNikA5CBZkLGjcAC
0xImWtUa9WMEi45cnKR9OW9KScfp/zq/+uL/tTVwowaM8pFr0A1LlViw5gIx0Rb7
AA8wRzYdfI+3T5s4K5+7KTGMqMV6ArpI2vzy5yVU5dWIExDv4lJ/JvlXiW+oMtlD
agnIjZUhGVX737iZtpaEyCd2yr2MkXto9FJF1n8dPtETVqLvQGmxmA55dtmrLmev
BeIVZOkemQHrA56ltqaRRTslzZJ0qe3jNmYKf2Po0JtsZOi4RiYPSanvQfb7r40H
23z59RrqLkDfEhT/GamB2EHowujTj7HvapwC02QCOc9bP5WeRwZ7X2OzAWm+h9GX
xViKyirmCuZB/ruvY+/3kEeSHrVuKWyM5idAYWAfTDVV0lYOxuEswA0CdLrJ1y+P
s3K7V4Wf2IayLjytM3pQTZQ+6YCAId8dZqLyk56tidgaJ9UyWzl4vpEG2+kUsoN9
jWtB6N+9iHE+0gL1B6I3PLeqmKmZPIFb+KwYqFLRXI5hAqvlqAPb3oH3EzmnGfwd
kAMCl/+jtHbtFwff3+UuBfTuZLIkSccSdFw3V70HQxoxhpfpTJ3fPtcTlno4PN/0
ftnAbKKRCrPMaDaK2YYmz+TbeKcmC5UuuE/ys4A0qdUr2sfzk+4J6wgMnciM3VX2
m+Jy7cA/01ZSL4+lhmxnpoxYBzeH8nqFbdqvqAQ2lrmpgZZ9Sv84jwTB09H818K6
LOsz1Be/x+Ic+W/HfQ1CDfl+UpKgsAph5rZCHblQXwIPt872qjkUYOATRqE+THIY
wlvhlidWPkGCI3bp+ENT1OvJ4KV7a0SX41HnPAOOtceNHqC+oDRWvAFfBGID4Kc/
JoM91lfk4TiBqne7fFnRmyuOUsmTxSUFkxs3c6UdC51mMkPiy7oK6PdFMEe0qJBb
bQYsID6ONawS/EbIZ1ANM01nqMJwgJDZVUzu8Y22OfDBqcKfRIffG3WrURgwuKQr
bpxJiXgKFpyTw/DS4ruSqlf/zAyyUh9WyPSos5msaIGRtjpoVD+wxM49aTKyRhxM
QdNYU0DbHnk+SaDqonDEN5LvJu2DsQE+C9JgjXLs0XqNR6Vt8knfoQoAmLvTtNgB
qCQht360uhzdVVpoOqP4Vi1FRfFo5bunqksrlrDF95o7Fl80g2IT/G7EIGds40BM
90b6m1LldLV60ihpTH/qFIjGhyzOAI0ZCKH8aTRIvBpz6IdsxhlkPcMMj0O0GFbX
tTlsysaVHnkb6yCk1ujzEMln66QD2aDxDrPtSQfiBVFQz2MDyy8aJBQJCfMrfSNU
y9vxw31hU+oE/jxMTouJuyJVy4n6rQ7BLprRU/Hqavw1AgY4C0QNSoZRx85NKm1J
nqDRqXBBLSRmBqvr59a9+BJcVIn4qtwWPOamFf3lg5FWULKMb8NID47ueRohoc+q
z/1ne4AjAbGR9MPzeRg4p1pbTDh1D2WxkmhELa4iZEbyInaZbuxcxl3vZ5Mm4cSl
eqzR17FGGSXPpzWkM8idtQF5ShNmiL1QPt0XSxwEB6x9enfbi4wdUmzAlhlnusfI
nE5/1bkope82zj4UhVECiLFRAT2Bur6Vbery60Ey8nKMaW1LPiSQ/UvJZjd3LNrD
k9lsYGffn0OlayenhzgcmLcYd8nXo1DkBkCmSy8kiB2AmtUVCmPXQVgXx37w8a+j
6l7ccWfQkouz+RHi5TwHKflLdnJkwm14vjvy/JEjIOE1a1Xx+/PyLVf3RNlsecfQ
oj6iIMXGL05mpH+H7w4ocbXzI0XWPoj7lZDT2qIUD7C/Aj/J2JqqUNCQzrt0slFU
7Ezq3L2fJ7yetE6vdI6uSS51kBNANwFPdrVtt5Ps2Sg8njLJLRLwTFPdOjuwtMWs
AxRyjT5NjNGkFCHsI6PmNlg03/T1kuxjv/YnGIo3/lfdlVKdlaQ+6gFBjgffxK1x
4resuHasJ3i/z0hsEO1fmb5rj+ylaNzsryfnenVr2gtydYn/X8dJSxkiRC6lXZSL
9XTWNkv2FLiz2HTpX6Nmhb3JTBzxgeCGptMVhN65x6zbU6YHvU8XlBHXwdTBV9Ui
VxwhZshJwiHNwAyF7LBhkDeYEVLX1lqm/76JXa4VwKfgbYJtJdDDVpB51EMP8Dr6
3iHUIxFR/iAxYxqlBcVDYxRoBC/6VitqVzQ5+mtRHr4QYDOW12U2+d/z/+7hMcAL
zCa2FvvUDKs+FDXM8JKGKqusd4PopKb0AdfxgyTs/k6bjqgSSvaJlqjcCtL5U/iu
6DccFE1vM1a3ibL6s7aWqv9gua64u7jOFt7gjTucZjiQNhADI+BS5cZBUjdoRwJA
JV0jbqn4sW0ji3dLfDaM09hqkSLkWklhNjhsi4p0nhyLc+HVFPPY+FbQi7AIxaT4
oSq1/nTFA1im0CcnClXpGlpUbJAOUr6AD2oKlkXSOlSwb7mTXV+8KDPsIVD5IW2x
2JrCXPjMD8baOvjQ5MsxsWFR86MQfh+TBhM6/QqgxcM7m0Ll1Xhzxzdahd9kxtlb
E3BFaBoz4HuwFVRktqFck7ZGmTqO2A8k+n88/phD3kfcMgx4jTY0QVPNinAdRWUm
sa1nhmFjsHF9QDK0TYgKXgU+rznBMXuGQUbnEP7eOR5R2DMkjgGn8VKhYfPT7eJw
fLw0R5URzN+aehSAN2C4hftHAgZuBiq1t0i3R1NIrO06VGwQ5KFNRMkNtjYzaSE6
jqXSsc+4N7QM6YfqCz+PVrJJ4QNWp2LsaTn/1TzsePDoZMB7CrWiiehvBntyYee/
hvldWv48otUx2QDNuvOJsTTs3VrT0Jav2ommC52W0TELvfAlBK0qD8aICeaoogAQ
aJdh18zfDid1+ChT4yXgDBS0ST2LBx4ne2tpS2+J19++xei3wGy1yy/VVbDWB41L
JsOQ9fhbGCbpMhET8UWg9+SyEpHADfksyZPw16ZXZcguizOxjSrDlmhpRg9L2xC0
NU77sM7HOTQ4kz2TASzWIa3GfikFj+zihMOyYgSMuVHh/6lQFbfNzU3wva90bmqa
mp5jOrUEbtobccMDg/+SpU1dKki+FRgd7tPyuVwSM4prXCmMH0D8w1/CIxBP5nrb
GnOauXy2MDF3FOQl/w8bIclQU4GOCsquBey1B44C3epJinIdXUnuW+rE0yVmKHKC
+RKoUcim9hZkjbbIm2OhsKPeLJWv28hOhWjQp5iH0X/215MJunXRobonJwYcypQe
Rc99wg7ZRz/qzHfzcNbpVsONsvmAp597UyNh90xLtp9HXLYlC+cPuTZYawNtgy3+
8qJNt0z1aFCp5kJcmrWU/wUiQ/qNZkZrDPcBgYruA/ZAJkb8TequXyYLz2jitawr
q0NaA5VwPbf4n5ifto+GZsKS4IRtsn0VFFK03IJmBIebgnZ9O4dp8Uyj2RmmvAMf
3XEgFNeCg5LxVojDjSJOgFM6ERUiPpNTip0e0R+iNl4vmgR35v12JRcQLn3IDZhy
L9OB25gI3zrXOejCb4k9ojcRl6CudCdKaPusyfuuCXswUOv0Npm11aSI+Tb3urfv
mIN6B1QoN51QNtCDxj//slQFJuaXocI4+mr1WsmSd2bVgAuLyocR3F/eFk+Ii9+2
XfXeHFmBMmKGbHAiLkGobYe5nZui1L30Jg7wCortkjkdP1WOjSeAo/VVhH3aQ/1m
9/G5rIm9II6DqzzIfMS0xZX/MJdG4K+qStT026HdnLVBpEiEoRDfZJwMrGWgRsvK
yVTSVj1aO86zGsVdUaxQMhzFEROxahYMplRzBZ1cEzRFN18hx0NS9k7kh6hj+/n2
xqcOgDKClelXPaSf89ucRafbIkF71hpsui5xPrObYU5s/GFBh7u2L1e82JFJnWjc
M56U6rcwRBLi0A5kwasS6lOFmFhywWeJ//aP7eSi7NdGvGcKnA+kcBRs4dtM0IcG
GO3jUGzdLY+E7m4cZJ5vTs7GJ2XHxRj144RUlycsbL5npFPEGmnQCkKRP78aSDIr
j2aEzDa0CGqr6zdAUqZoRSNibv3BXTofvI2s+KZwzwtTJ0wTjoN7RPqbP+CTfeQx
AYvVYSK66Pu/jnkwESavmKJYUIP27ROkh9TYeZ2IbHKCWgGqCMR5RSmCs8VN38X9
MO2z/2lBoCDGWQxCLbewlor+KwGFJr+7T3Q6BY/86DucH/R4Q1+hSdejQXyFQRPN
TJnaFIzkFT8QsglzRj3Nab4lMtBh5vSrF6cLQDS4VhrRHA1zVM5wYppIGsN3Sa9x
JtIt0yDKy6oEa39EfLgvVknZaPMXGZb7Eh5DBNMjvrsF2kmV5rfnUBfs4JtiDS/W
nP+i+oJ1C16+Oaa3BvQ/rrnStWa7GTs+jK8515d4pvQfx/8O6itU2kJYafKbQ9CG
X3heCvMuiyllL2VH5f178TrY1DDLbmbcAIEmaXSeNeAEVFREwpfNIq93CRVDh0fW
QXkndCA2OeItywp/VyTIM6EuwzGFz7i8cXCieoXkgZcpc+cJDtzAcQ7Mf8ecBLjH
xjMn+vp4mF6t7wlnCjAGA2bse4YEz9dhs7RVhz+EkysHi9eR/xrnb38XR4pGLycO
dUGs54yRbT/OTsuRDYjOUPrAU12ujz4L55audnheHBifY2mcscgtwaRi5TRiMxio
6EMTGf5Q6AZ7GxTWqNyXLpcYCWt3XVqSLutTdNzBnkBOcOZgcftyeqUxBZYaLWNd
jebAGEGDCGJwBniYNS+tWNR+QftYaopcRceuIu4SZKGRjylx7Z4sKeepstdxFuJK
KsqxRezXe1uZ2Minu0UJPTXAGfcZCS9dJ4Caq6SUJogk6Wr7vI77cOa8FYha6b8x
uLbZ3CpCWZ3NIsJvgYO2/ZDhXGfQNBSr8Yzt+ED4Zz/uUgvegr8hAgra9PSwl9j8
YUfcooOICaV0UKG4GF+sxnxAgFzm/oYll89uS08XTWyUcSjb6uEMuk0kNsr9xsHg
3HEAY24iHAl336Al72W0DkpQGaF925J4/obsYhpettcFWVZD95j2W6vTpe3w86hb
kk2b9WcEbZexMvcIztTkZXnC8qYtP4InSANBkKvnn98b0u1Pq93gR5geSoCNiIEI
874PlZ2OnGwzaTr2uk4Uxtm4r7Lxlp6dH9g7txl1cSkZno3K3qFkWJbPGdqHFFM3
odlIi9KqLMUNvJmm9hFfk+B7d5OVXI+KTyJGPswBx2IzG5eqaF/a/gPEp3nnMyxp
a2l4LI6Hix9rFFOMW1aiJ4NjS6Topb2lAzt1tAbNx2Ezn8kNt+04nu4l+UNiHJad
RRCpp2bZX64yKMT3QQ/vjuiEU9/oLhUMf7bFxZwnMVFSy1LGuCeSN73PgUFEF694
/1ZFSqzb3gdWnb9BqZzruFEJaol96o9jmtBEWX5QEVJSR1v9A9tX8JWUrF565OUY
0nXRP6/S8IAmj/r74hPduFO6H5bL7sfJPixVQtCcVB0M4DmMqrSJBTowroLsn1en
k5BZtpEBC4HRhVirh6ZYh3V89LBtw2+R7OJhPmr+5uVkWDMMP7EKVvP6ygAFfzXY
bJT6cuPHiF+4crbCi2I9N+IrkB5Yo7wLY7YgecbnSa4wPygYikfm8G+CMMgMAQMv
wjLwJyo8Muk+Tsr9E5+vKskVv8IsEwcqXnIE9n/taaUnEsUedQIEIbIQyc6Cbrho
Kyayd0jyblnnj4Ww1YmnSbWg+Kq8vVYIwU9yBz0TNvnOnb0sOANhJL7C3/bYxeP8
fqqGVr1m8MDJQzd7IhLHd5iZW2vHWa3yHSvdCdXtcS+GO+aLZ5hN7aM2fhMG6yoa
w5S1ylBamR1E4aT+GTD3Ytx6g0b+oP5lieXAuYyKThNxFNV0ora2nCJEAAD6NS2n
+WSBKBxChFtt/IUfSqFgCnqRktsYDQXS40teqe0pgKijvca/tt1YRHHaZdPzKzKG
UeIBl3CUI7Zeob0vni/budcT8uE9XGwREk8jXibJeZwkQIBrQ512VDjmcIPE8rx4
/IZ5wN0xrkMexugjvZzHLc4Cw+HWl6ZiTkJOVq3zEYpxoHYq3DJWOS5lklanf/X2
zEWCIHaEPpsQMAxe79GpYem1vZixtRUV590cctpHOngMIsjL3OwVomtOhfHW2QwJ
SR4++IsNvhdaGuYShPorkiNf1wguscfuNw0EeNdyqkXT/vpuwJIJW9/Mis06OOcg
nkt98mvS7teWr0/a7qrwdynZLD7hLtfSsv6Qn0+CdM3NiNfMPrjJdboyT1fTZEjD
U94huq+niX45qIWFYl4IH5empQJ/GOMSgTNuJcEUaTP2gJzgm63h73Zu2CStpPXB
WHaeQoYCvGdQUSXeOxL6XOYsvfCh5c7recKi9lBBnMNjeYO/HkHZf8PnffmSZ1/p
3A2X7FCtOvhf+6D85pTTqPU1qCdnSVwO1FJprPAH+J3BmBDlut7T13RkGN/Msn53
709/4lyLl+I6ER4ileDnFH6VMhrzkgPORVRm8qIZs2rPNfkVS+a8iL5ODXMYGOs3
oNTUvxVvorZpNzGo9o8xSiGyAdgMaDti3np67u2nBERVYdOrgB2cVltaxvQKcRL6
efjCFYyrl23zpui+vfnNwAFqxpz26rXK3NzQFowr2mt6xr8W9xHauIfQjgr8J8Nj
uudC4KhejSvIp2LJUvNOwbvo+M3JNBVDbA2DJCHG+E210YBzD9NN1lab/fJTNpz1
pxAIM9Tso4+uidW45dH9TRaxEvmBgWyXqkvijgTEPFtVWQh1WwJa1f2RTlhfxxE6
mhqLCwqQuEMHgkuVSlgYSjSfELCtfOlLhybE50vdyh1ua1QJYDTqdKBn2b0R3/+B
oiYj0vacWRuAknloHrr25GwQFF7QgNYQQ4aCMMSEMtGPNKhxivFi79k0IYHMnacd
hp9LjFjVyO1aUY1BVn1R0jFTnLjuNXRxEuh35UGPYgMzzYbWm00RsztyLrMdqMWK
9DTzGdjNdP4YI6eeWuN/8RRIDylJGnWMM6fp4pdE3GAevAnLMz1yGOrYV8AHM+al
5CnfXWsCmFk0Os/OJ/tRw8MmhNIHBucFV0h6dNbbfA1cbHy+xmmRC8FZqerE0Oz9
wCL1NRMgPmoKQbogKVdM3/DaaPH1Si8s/lPQKmttA3hjPT5EoUJ1DmDImLD3K7w5
Xpu74KSY9bkig+4dj5rtIsrdiBTOB1c4AR0jsIR//PgHQ/cZvZ5LMGvMfATD/ses
f0DyK+FLnF1tUO+OmFyjFHtbGfBIvoGI1NBbVCw9+AtJOr21BBASbFpJu+D0+ofX
AmALqlTknekGX6zyRFGV7cVzON0vuXmSobM2wrCyEfY1mU/uTwJGgtrRJm4FiPBf
C7BIc8wQuWyLd1zjzYughqN6xTotEtXlClhVLGJl7ABFG6vzmGrNzhfHt5nsMVkW
boxm80L9J91Azp65m4H6RvZBNv3DpLCqny7DIo9Sf9XxG6pCEPl3tcx285FO+Uxo
41UPh2urkFnWIMK8GCkpmrKZqTJLM0cGhcTaSptrLAuSQ9wcVd5NYU9kRpDZpgW3
J1Ww2dAEFtmmpTIuOV3qoU3w4Sw4CPl+Ns1T54hAn37dVLHp6Z4ySZKe5U+wcjtJ
lXOCuu26jVvFnL9udcEAJd5QeqLrLvLncNqJjdQh3HyP1QMUIqGuuVlGtrZ7FLGw
5Hro/PYJOa3dgg4Vo6vxRvqIigdIm4Iva5u+MnWU0t2q7utkjy/OqNYpy4DIOAMY
YRgJAnHV/V/D7HYBUaKg2G7jFwYqecDMByA0B3fG0PLgavvUoQgBDsHtI88OsTfr
f97yMcFHqW+fgkMoO1JGXaY7ldu6uNQ9zUfaFdue5uBM7KI6QQBHJRCP2cLtpkiy
jqMXpCvjH9GMq+RIJW0im7ubCJ3sQyhLh8999+MTPP6lZHgNYA/fOaiCbkFPAnca
shNgh08YoqBfxWFPb+cPjkafYiHSSmS8nGyleZ+9jj3BOoH6cF/e/M/42vxwTj43
JmHcuzfpfTViTYNO7X+tJBjeZUv5tlPDX/TInD7ihGMtWAINzS1NYRENrekTEraJ
4QoBHqGjYlQMbxfBI6MSdFkn5Q5Zb2QFUYwEwC17KthIXqoAdQdJFVNjNlkZMZpg
Rjulw/vOayN60dIdzEvn96G/XN/wW2lxGGXmSykpE1RnQ+9GvNWqyk+aSO9Db/WS
KgygKxYoUPG3MQMlCHhkDj7g1ArFp4rRwbiRHaoc6lhn/A+jExgF/OYNKALegcqM
6LdF71LDqiOYocxqMSHnHXkxLTcZK89evMY2jXyM5M9RIHE28+zQFPoD2lSwBu7g
BrlJ5dvrKdTJjkHl+YacHdLcUERI0JbH52BF7DeF+QSn2Q9lj92hz5faifpQAtex
jiECor5B12UsfvWL+ngBWiJXN0RRyly/vya7sg5dVRB9wg4WhT/E/V2zpKORg5F7
pnEKbhB4Cmy45KylH7O0EIQVgsY9g1DmYWd+IKDgvoVOpDdtBY4M56XNKqx/Ua8R
vXStv6VyzRy9gTD//fsQkrzvRvUDT50BTyKahQDB2aveSfGunDt2IIZPO5yv7Qbj
m6PNtnJUQiV80IODK5uwXlc1euVoTmSHUzZME/8q4SglTq3BUY7X6RvXD2HaTZfN
bnwlMAk3I7o0tG+MlMIHdSwJFoBRR30CP/5TYxtYUcy/HO87j74sxz/X6tpdUPFq
eUQzJkuxNYxk2hEZZ1yPmKxEd7TociRc7Omp0ZEMxg4uOB7nLWaR0llrWNSchhQ+
MfJy22BpPxgRW7tulLp+dVWZvEqSSLt5LLDZ4Y+M4otQ5Eeys2Drwhlc58W4ZOok
A50SemuG0uz7pFaTTFZsYO1gZnOjab//zD5iEkNCqpCkxQhBxbaadcLQpj5/I3VE
gxFXI6du3RmGzkN91jLCu+vZGoaw4YgS/4fIhTHimc5uL+CerR2imktHevwX0QL2
aRlMipOUEBMTXITRrfCIkgQMzc+fgZXNjPa7GN4mJNNzXgm3oAfrqfal6Tdv8Kd7
eyf21lQk1TplGgkgvaU6WJOjQGFArUXAt1UZa9+H+p0Yp0iSp0oQd8/lGM+HcXot
VMm0hRN77AQacQKL9QlX77ewGrekXzsxf9RSymf3sjUz51hvGlOlC51CHPkxA+1J
jA2UAffDTW2/+mX210ZqENrjnoMmtlLMq/pfGlP+KP2MVEuElqv7g34AqeG5aVfs
6PtZnrtVr0AtqmglxFNEQDcGx/iDkKFomVaC01u1x9L8D6IQN6UNACA8SISX4+LI
krtWTmna2YWaNBYZaIUnrkktWYHoh3NopuVtTHMnKXiq1jMNms7PvK6N9uByRJZE
ukWr2G/lOZWlp9bhJFSwAG4VoW2BUiAJLSy2HQKg8PYG8mawaj/eIhnTGygT23JG
Fi35IBHy78zui3IVjyO9PJ3P/2QqZBM13tEUbse8sVJz+eXcseveKogWb4pkXA+p
8tiuRh/AM8+YAmX69zLobMqZEqXWkIII0FtBtxPcxWNfFumJTiQlxK87Br6FJ1vQ
LJFAPtr5ifC03N3aHeQNvb1KW+zUTkqQyU/phDFfQpeYRsPj64CNY9Pv3dvZk/MA
oOzMyvKo3/eFoYhgDka1n6/Fh7Humc1OLyuRhJcxynB6PEC7hDqOppeIzD6SoqVr
l7CsisbCslmAuQyQp9axQDC7FfLKSomHHqhGhljlSl9LChM2HcNkD5OykzdIIuY1
GrJGqrebN+9r3oJXznNmCFyfB8AqBVbPsNB0xea4A/bh0qR6kHiH0ZpxgF1v7zeJ
26W6eS+NcPZIKc2ew8Pc3jbzBoFLnAhkC65BbyUme1gxE9SiOBPEXroRmm56bnqg
hY8jDQQi2ZNSiUfxUk1GofA8BSNThY3g93f0ghFcql6Kc5V1q1/tXTr5aTqmMLIj
/gZdhpZ+tWxK63h1616oAmRfzgtC7T0RQjLFw9zhVOK08spAYnxNvh2gTqdmzut4
YIUtPIkBxfcl7VUoBQ8xKnP6hkclYeYTdHvWFpiSmcIGzoVrfIIaeV46pQ8bkrH3
iTTQ0jV8Dc0H2aJhlA0pWY33LJHlHSb+k9MTICPBMBneV/AslrPBXWAhVgirhBZG
C9UuaPGJvgRZCmRPryMB4Udke/HT6vqmeRpsy1DeI7dp48CFck3dhjIHn4myuSas
To68bM0Gi5pOfOHB9p4Q5usUb4/64tfUiIbObm6syeUJ4IKqXlG09C0mQlKDN2CH
aARVINiUrPpoEWJOF3YHAGsAX8oL0HxtcXxbY+VFy2x+4Ai5ELliNuZLLUddfmw3
SIVE6L6PStTiNP8eYsnof3WBnzJik4mHhpKBVswKhLUVQTalrsmRFkojV9WfeNKU
kWSXeUcEM17hA++aHcrGkJ1px+wlG2soL+oeQptgyi7m+q5eUOCMnBHPAdCleyYL
z01akx8odrPAQ/LQjQoiINx+t/3jJxKMYaG1Ok8vJmhDroRD1diWYchScuwvDIZy
NMwqlNSQAkmP+ll+eC9QfY3Ow7WCmW+4SN824e3FTNrTJyfrP6IB3C34RwNWTwpa
D1X5WHM3lGPLlFIxKlvikzLR7eX0SAjCR5A31KCSacwsGFLn+YIDhmWZoKy1kxEt
SazhB9M/4700yvshj027xbEko8Rr744Omdf6RUJ5x8Wg7NsBuZlfOmEpS96P24Gg
2PlrJuOcrpTqytZ+1WRBy/OnvQeSdthv6mQ4nkPp86FYjj8afGT5Is9FE/+7iPiX
nVMdq6Nl30hsTxU4ZHXixlpIfiQ4iAvFKiTgGsD1u1bPWIZr7nqIT8g/NLZfQ6Ct
XiY1S6NzUe6xCkjxXpiGuNXhWjuHkLk8zvpPDxW19oxuKnDQnE7PV2qCEmnKvzpf
qW/JQZrnPrp+/VbgTBXvjGsH+RaxjopCXh/I1rFfRH8UWT/AVKfJUGPd+9zMbQC3
2V6pYqV0Ud4x66YS5dHByOlcC+Y5kyGezWwDwFlvwisuo9JkWlXgswFWEUG8pxP2
wCe3U7gwshcQQPxO8iFnlt5bv0OoV2HDjW7DHuR9WcI4JkN6WeujGwCpnBwn0+Bu
xMTPKMn1AnTkZcjj7eAiz5JLf4vdggm76TQatvbRWTnM6CAR7eT1hzaRAFzGnBJD
uvgi8oKhhnObWqHjvwKNoGDGZgAeMS7mgz9XyqfpBnRO8y5qfXuqf/Qd2J/WvIDi
GgK0qdgvfUaC+JAftfkZYqdN91otKND67DiKb2puEuJq4VmxvTjE2rnVM2ETNaIT
EKP9NS4GurL0oofWUolrPzCWtofxeKY+UVz6n/6/p01umKwTyd1PoX6QgoNKzpip
7/CW5ZrzYVSPYLd8tM6h6F/peTfxAXZ+zHep++d2iZR1wYDPkN5I+iCc3tjTfG54
dJ4do7sflgu/Cm64R3nOV0MjfvDkNG2lNLIAqMBuKy0IggmA1qD5M3r1vgklQqZf
/h4zjjnk7MFjtS/hUamU3q8rwZrquvBeQ7BtNxkXiYYfvlxD+s2Mkao2gbuprVmO
yjM24si7W1GnOGhJ39UvfSBhF/1X1eMnzlfHxRiGa6fXXMWfES5RQ9JdetLd5fmn
DVa+MiWy1J0GDSSpVvvgLxsE63qUXHBnMwVuD24uOKffZ9fwJC+C6G3Dvo8AN9FE
hTH8KKcAkxt+jSofPJbUzwCSoJEkK7Hp20PB2L5DcKkmBV3w+vc88eTRD02iUQDN
IQDacbifL5bqBp3rVGivi3EITLnQpcDr8qW5YjkyIpjePzCNQTRy2CbeDYFyWuyv
DgRF8/KGHAcHC/scGvzyq40ZglMcMWc3x9jYRVXbC3fUMA6llZLloCnCSHAn3dtb
9uMOmVH/WFR70eAX+N4OEbnIJpArOQiFFYnF2O/QAAIoXI9AUVkvhtsS4h4s6z6q
mrCLzRjdqbpjQjVIo+ZBj0SUIi7seO1oOykryzJoARHZ6wiIyV+I5/7RWj22Jw2S
/EseZ2IkQN8MRCENRx9Vn1KAPEtJMoywIcCX5aaA8eFr8IgvguKIodFcwBO7v0jj
yvag7g5Voo5g3m9k17DXl8ppNUGeDx7HGlDVNj4POkT0YtyhNhB1IeTBLgrIcnsb
5F/Ftsm2H3mCwZZh+Nq9sgcAtkZN35ZEJja9ODnU+SRJ0vKEp2WZMSahOu6Nqsys
3X+G27DVkEnQwTx8pv1i0L7L7kAzbkkcfcFKrZz9HCJQYzytea70mAsYyFg2dLBZ
g3EPhADltLlpxWcoQDL9D98DOG4HqkDDIV07vTgdTqA92S58h6Vm8nuwyLwykrnP
NTVWzgq3ZIasm96I5iqYjfMgEfpfDo0AmRVnbQu0EYYYEHLnnmXxA0AkBTuyxBxd
7D07zfJFXciy4p6Fb8FlDjJZumr+5zH6ES9u3dEDMR+IbiCdFLnDvThqgBNWu94t
/Uy0JwO13Eda1w85gPpltamTUxeiaLmMQdqwxxsCrqMUe+h5ZqOnUfaXNmH4ONE+
3N+1PBo5FwYXiAo8aAnpMWI1DNCXunb5nErvhxFgKDa65ao+/9DBUpvGPOqcillZ
iBjsCL4l3aILr3saYivk9UO3ifKxvES7t59HSDWfG8a4dkRnApHker7xy08R0tu+
VhWNKZN7V044/pIOUXuvbwGi+nIMYTE/5QH+910FHw0I5VbA6gHQxSB/sv3lELu7
lltAGvHfRwEzLeKYQRtAZ26TRSnEs3XDeKwn1NOePWUjwPSHP2vOXvLT86TBKReJ
m5L2om9/hAylUlW3tYt6Kde87bYOTilVo7M23bIMahTFUN6XRC6iuUeX8DDNHu3k
/8g8xzaqytzultyoAt/4mYg35/CwR1dNS9SJuOJgX9+fkQibZzozVtCvk0mMi13N
/LuWFl+ABzOwH2tt7PemuhFJXXn8ocWAEzN9F8epg9fbRLpdM/7WN/BTrcJ14n9d
DNOMjt0SXhpU7S2uf9Ndir5Q3DNUKQUPNeG0voM/8JTabDHDR+TOt8c0+sw6nrNj
5UZvXzjJ7GCq9AzKmRuPZfFCbCSEMonuzj/Ynq/XReo8Tk8i3m4X4SZN26sbromE
tLT2XxUUlcHWni+c4KqwHF+kTiGkwKT+StCAAzKWxZtqHMmFMk2vmRIh6q4ei43d
6e7THzNCi/P/T9iiKyuTvBghuDMw7Ig69fJKrn2+RDWJ97vSkp58nqp41EDo8MCP
KEBsdttVP43WaC6Al9XMG3xozGFf7z56Z50y7EYutQH+WUuMQkuesjdwZM/pYFho
nniBBdwN4hE+i5YNf5KN1FMlCPmLrOUhsZyTFx6Y4KwjazWWINjLfUrLm7Zl1jyy
IeBswoCkQ9Q4kQtbGcgq/ScphHDgX1uG1f5aK72mMwJW6xzb7x88XxJyMIAO1iqs
sZsjvoX7rDfqyGGC/jDh74AjbPaOWC0xygHNTt/3glCHA5vHrOjmXvNqjqJl4wP6
2nyfDofE1rSZvFu4rCjKBrFOmF6uyZltsi1JXwdMZUKFsj/xg4+X+QQQy6cawaDt
JhaPWmn6QUmeyV8R0BBc9x6vTtDN/WhXxl0iO71N4ZgT+/RLsWLzvPrBsQ8zbOjK
eaW+pY37eJJ3jHXP49lChw8/npfCF+W9a1+tJb4piWztUFyzLZxFn81HS1hTqojV
3bEJ9HIcWfy5XzyYoj216BlBHcqe8oz/o4m5M1kphU/zLc4BiXuw64nNVdEkHFi1
uj4y7F/1jE0Mb8XQ7/T5mIsG1kKj/HDBnhluff0pZXlP5fYqpBpqqrQGuJCQ/vMA
RidDzEIg3bvgvV+vJ7Xz5G+EmzITRHiEm6kZbK6o/muiiUh0zUWM7ze8iY6FTaYR
0Koih6jhMlXqpV0ICkt0+le44P7AgZqM57QvSMWAZx2NnzpzjHdoDOqB2E85BFMv
WQz7q3NNM23PMlnQXPm/YptDiemxVVbHbrst3lxI22V3Vsjy68RIZZYE8jzM5fap
LFvQDVj4VWqqHb+lFpAAk/09OV0oQDJ+nxoMMIQeHxBz5fLCz3eklVJRzP7fPR10
9Hu61u1wb3tATUb/hA++oVMp85teegNFRMrVZaaIMKQVi2Ml3ZMU9NYCUM5RPgwn
cp6vfPm9z8hU9w2fLA/pt7m5tBQ+CVCeXNG3GPzNGul2g6UclilcSQ1I8OffV4gw
BXMwYN8jELE9s9DQPsUNjmhwhz2O9NeG9TmY1WpoLj0q6aF7y1/nm26pJFzipzUN
yGFeV/MWF8dRlb8BaSK/4+0uk8cOGPruDBDuU00vMr/T/ZJ9ndeDwPg6O0P9cWOp
yALZjOupT59CY0H/mwsmD69InERTnk04kU62dmaRLvVXnUy9LoTIr/y3BvtJJnuM
1hFre1h6/NXK2dTrJNNA5XSKx6qV+xBgKTlgNdw42HitRRMnjyRx2EqEGFtMK642
Pex2SH5ZRQ4YI1caGoqyFD5r/83DhrD136dswD1VAbYoAkFi3YS1XUdJflptRTpF
x+dZXvOspK2jGEpu+ioZ9tBQbgcQTn6j2yfzj4dc+Vrjb8hJsDuxNfdna2Gs9sNS
ZZpuOi6AobDA7EURKPIAlCjav74iDirSRgYzvlyx12kxTVSZP06SeG4Gbe34DKaP
fNMn2o+BgPjo0amVk+fF+jGChRznPsxtFcoKrrJ1f3q6zZGLsk5JBwoLtl+k2ewq
AHX0f7mW2yoadj+DX1FgAZMYbaHA2ZEhXEJATLvoGfMeOcXiNP4yyNjA2hmGAHvL
K13wBu8s0yt0q8Xpb7NGspGLgO25tYiDaUouLrLFD2g7BlEdEiitUBcPD1agESw6
FWGMeNE0O6iE/Tyr3whLqUOFWZx5q6WNzFa4+QDvm1cttOri6GRH57u06WIKTJd2
mA7fUEZLfAkeRBTSG+AInoqRHBTNpXaOoSkdi5Jbrjc7Ro/Sha8wm5K8I6WrLN4F
BXE+RJvzMVzZuniFbvHjmMVnf9QWCZq4d8uiPizW8UAItrJ2FkmjzitO26tPvfwC
iKBGEbYIxqkRJvHtz97WCw2bBJovG8RTbEbCf5aFXKtKHSGCNkfxroFhoEZPkTvc
pwXBIVPy7co9dOjC9MAyNYDmAlFd5QDMoY0BYb41E6GGu6WhUyvq3Eo/04eMxRu2
g8hROVxmE1AukxyaSEhR3H9yawu6mrWaFYapNkCsMkSELV2HZm2W+UKf6X+qhlSR
/EVwtfa2o7NKXc4mO9JM1XtEMSa0143K9Jo1iC7t5imjx4KTqH/Ejvwd8TpaUAyV
FtGeuq8GD6sKfDJhspMmWsTsjB9zESY1k2yLuExgGl//0Tdg2kHcvaMaMSR4CvdF
0fXvyWIVdNPxEnWNNOpY+9o69iCnBMIAQNZXHcXbYsaLPOeGZOdsRwIGR8ZZqEmC
4U0SwtcI3CGWdYhJBhkMm78IvZrIpPEA7dFvCmTxl+/y5WqbIi0t4AI7t77B3jl0
kvjNPZhzwf38Lm+Zkv0bLq/LxHrZfPqKfDnSWTg0/u4AMMioJegpCsi4WRZfPGTP
MpjhCdPATE0twna9wnAIDOuDbyMAWAmk6qApovprL/D+YSSnRnYy08i4BWzyR7Se
AW8pcrKVs3I2vlRsGLL/JhE9j+fVZOc/zRWNi0CCmbyQUL9GsMaBPw++Z1DLu7+9
tGIVN4oUszRmT86hK4r5gwpXTdRjsvND/Q53ZqzUq3X5tvVBtqJX8bWWFTpkyU3A
BcceA5CQXrJYiD38cvG5OgHkJdJLRZCIZMvA1Su2KfFWGVwtUTDuCEpZyx2pTkSP
6qdA7YZtPxmttCvz5810J1PQwYxtW7CYk9HlY/d23GT79NO6xoHpxSEZ+2j7i2uu
H7X+EvQbdFF17TCCwqQpY/pE/VyjFyv9iIMd3nHSSTcnQci38YicG1qs3aCwFRZp
kbjZ2RFTf39R6UzhD2LvF3jU4cX7RGfVylo1BD8Vw6vNUbBynnVItkdEaO1x+mhQ
SMwKM/+Xn3+9Xx3zD2WQExyhF8dOiz+pNP+OSUF/QBnLf7xTnNlebYrpi2HwlU7c
rXqCSudXQWOA+dJ3zyzJvN1Igi7XDb4iS37kyE9SkX3Xjyh+wN/pOmpS5rPC1bPf
0zqFwxgw2xQOFZBX5DL2MzABUE8a7+36XN8L8WD8+Dk03hSPC0F9y4Jd8OpLTZDv
MxZb+VYvw0aJXbPmEVuTSeVWlEtcz8MyQoDJusMJFSqFNDTw20ZjYG1CaH7hFxBC
Iml66R5binINYD77aOocsNDkV5CmJHx4rbQiX6CgbsxGP5v6fmfIKEtSePCSg1bH
VvH5LLH5toEXCngcnGKXkz8CXiGNeFuK66JNnndkOVPQhO1e9hQlhcjHGZ/j2CV6
aBWI58IBo/XAzSiLSNAWKvArmmQcHOVTUQmtpfXbaY4I0/ud14IIQfXY0eNA8QNE
YmEL1+mLPLa3tlVZHUUBs2gH2zCa/4296CE8MqL4eeh++fckEeazBCxzOcRoxBmk
qVFkV4U1wThIu8BABZ7xc9y+oHR1CIOjZneDmiycCTdCioIecKZshXEYwxz+bf1P
Dc7DEGi5cMZ23xKwfi37H0GYyw9frKDFJCZVYnwsDJQbl/oDz1BffjLTj+QMuUPS
9UYZJLiqkK1LhSPszBupgD7gWtZzNQvD+VQMETORFRV0EjspGwUyX+IG0xrEKpnD
zhlIGxnYp+vfYgaMffTACY52TLRaU7cze3T0QntICCm+TL7sPLXtIYRU0zzkbKq5
wBqlwaubPY7RbAb6NLG4n+KTd0JIferOmM/uLzxxZ9tm2QraNtOOurj4OD1n4Oqi
DZhpXWDhHPYcu7x+QDOPITG3sWZkYqf0HyJyXWHkp7iLQaWJWwlgwi9UZN9571ZA
INob4/EEVNntn5M8SP9BOPQfE4qyULfXmugE6+jUPWgTNfImBSTxY3InYTtdCJn8
NM1YTh5BCa9SdvK+HK6bMLpL+UKaDiR8GuapnsYbProe/vqhmdwAGPxYU1ZxyGEs
ewBU5+f1mu+oxeDa+SCOOAd7oBes4PCbKSmPMfhzgFv3ELrb+zU226Vsv3nM0TcA
9P5Q/n37MZrTSk2h8leA+mWcwTENNZ1x83V+TmJeXiz/mhLVQTm86xLVB9ktcyrM
y0aGJF75aQ6IRsYkuh61qTa06LeLp/IhNQGtNCb7zP9BB0bMFYgY0+pa2qni+GpI
hjirVsWSUkTez9M+jGWNrqWbvXH+rX1XsMco3l2HyzqfU7bAn/5PVfQbrTyjD4MF
+a+Mt2JTHphWkAmcM/6kUzFiXOuQ/YBw5ZX27AxByfSrJ1CqlBN4H0Imsy9ExOvp
cDTYydiZE9NLYeUYHQsCoM6E954ox691oaHf8Zp19BUVfdCDteG0IDJOiOFFEAu2
ybb5M1K7zDuPpUpNNHN/pFiz/488/wDU32XvKPVdssEf3g/5JrF+aYoVOnDDGF73
wqsIkRy54J8oFr4E1xnbawiFhd7eNq0JIrD2cSL/DhO97BEe+VAjyXjAaU2LIQ1V
Nfcpc6vHuSVGU0r0wACwvgBxtT+LO006yGqdgE7i6QqhHSqBIEUvO7YaK+FyiCPb
mRc8ng2WaCXeOShHDtxEAzGFLV81AQ0bYcHEAr0wzMMhD5JOu9wnoQdMOhSQdIux
TNCv0JbWl7WxBZqmLBCqOiu9X9B0KkXCFz18DpspJrfLuN6yBNac+vOw/5n86X3S
Rxo9Q2mGG96bxKRISA3qqKS+SW/p8QgBJLmdPtfBAjHWSatKPR32abQQVDnSP3+p
rOR3v5vq4q1RAeEw9ZwxDpF0vLmYnKApGB8UXjsJ+EUxgtGlvFXuEDFSDdcTL/+T
xpttroFSTAJ+eChBcY6i4uUPrHeLqm40f7ZpwHgb5q3N52V/5DgIYQVb6ey/ESiC
PtTPDrjE3v1UaqVmHaa+aMX8Z06zJe38m8zNWJvebkwBpHM2c/09RVsybVX5wNbB
PpOnRWnEwDuXOlAhotXZMBCjVkQKNVuzJTY6cAydu+dl5RLLhLfrI1m5mO9Dwbx1
jANKQw5Q9kO3Q86NHhN4Gk5+k+BUG2+n64xWxfATnP5J4Oqb9ysSgaaavGWvsNmQ
AVutHQHFBtySW2X08Gw9Ezyov6gFA00Nt1N1wJrCjExn4Ln9iDr+R0EKe1dEtvAi
fd0HmuO6XZOYj0AAl+n+vuavyvbMDEPA2S/kgcWufUQJmd9BxT0juJDUGzXGkD4S
JY2Nwfv1ksPCgWtEZNAzDxqsLDvWOudalMKNkGWbBdqupyjoyfoJjlPIb+zrPXlq
g2jmOtD0rJ2FxcrpQv6FxjK11noJY18K1hRm0eup1lS20I4gFlyvjx6kMbRgavl0
5A7YFJNXdbM9ogwuWCRKoTm3q5ESFrqEOcHX0sVE+SBWGpFgM5Ama21XlhB3VreR
FEszdBAoPy7jFQi+eLxkvfN8Te35dsXDIOcoQTQNV1UjrggDbEuG9HeQwzrzAidp
BCfTSFuHBYeYr6ZvoQw56aDWa/wvfmDLeQvbfSyiqdYbCSgPWcxd43DkpsPx7NKo
FZ2bDlCzK2OgFZbWxnBEz4o/NQjR4d/YgzPHrBcelmecBPN2CqgSgYvknikIXFa7
U0i7ACraX3XFBT7Sp6v0f2wd7ZD+G6myD/T25xiP2LBZ7d9Uqs2W5BgPA0mAehgl
NRM/yCKjQJZDn9KQToLU7OOmbkZSdoVjIpM/Cc7IHbmnFngglARz0AsSUfo7jlbO
8j6CRFKyzgiKqAtRVNQcFN8cs2LoH5pPGGpJ8hoUYmCbBouxiSSdNEs+goUbHRo7
yVJuExgmi6tJvc98Wu1ibSa3/EuH6XKQfZpI02zRkdYIGEmcZ7uRUb1sVkYLSMi2
APwunnc3RlibpqDI32tNDBTMegMdNicABQgpGv5tioVVFoOOKkXlmwieE0hcm9vw
FrpVD658qu2nmK7zc8+zDzvl47EXDzvk67M8M2ynuAKHzOkA18qxcJA8fS/hFy1A
vxwOABykVkTbFx66z/luFXpNpz+c9P+d2SCdwKfKM3aSUOj+LsNRSchtphZKviys
53xMUaS4hvegPWbilqMuvJLc6AgZ2AlZc9nGCq4MwThVXPptQqYBApW++RrrguIP
5xrQjSvuovc8LXpRjVR+Ev4MqvmL9AODYq0hTFUHG6hqCVjUWb5rImHvOXgXKNCK
c2FDWmwXYzEH1w/gB7cuW0aoXWwNsk31UDb52fmHeaO/Zw9BQLdVwdPJK5y89l42
3J7b67oCclNvkOBWkLr9eSLxL5Xl3WGaPT+K8tDAzrk2oKB17P4+WWSDeqOEQtp3
oJcrOicqGMPRapa7CngKVBYzAeINrEHVlHZI6ShiDJPJ+ek+XxqOutoi65a8yPsD
hwrLg1JokR3Z8+38Ta8ym0KuNZkjGXm4gUzk8qPzTV5ge9khMsGPrOzyc3kPTruK
ucHrjacJE2PsRyNE6OLi9Iov0OC/h5Ot4RUsvjRRWdp09Qe/775Iv/fteJXOVESQ
JquubonkT3tRcMeHJgjTIbTaYeZBtQtj0WKBOY9gzflTbTmz7EVhRx1HHJ0svSSU
cK02j6MwuB4nNsmWlmmDFNiqaH95MBmgYVbx7Tvr1kd3aGxpeYDwzJm4rCJYyZgl
Y/6y1SwMKMNKTICVFScwOmkYAlnlkbmpX1m7c674Qeh1+3WZLaYYHwQ9VtWEyCF4
KXqJ2HxvrbYmDBt9kKpPcq2wZLJPGukXWZSJO7mPCsZx0oDh0C6Su0A9UvZz4FsP
n7OHA1v/ZoMZL4bRZ+E5vAN/+8npZ16UXFOoRWHE2eUEGhoK1EtAbYbk5VDXG2pU
hDNW7F8xYd7ZsUHLyN1TQ3XnRhBfWNuCTedBxhxzmK0POJxrtFtv3uXjc5zGSuGb
q3QSyNoIxSiMBNKLXoshwXcG5HgD3GUue/yvHWBoFtbZLwMnaAvGV5xEdMSuJZqB
gqtOLkyDW3vmM24jq3OLMPnDfKCVxpzMXPKdnlXAQIaSwB9hhijfdaHUCX7FIv4j
uZeixMY1fxem+9wFh5pggAlXEvnZohr6BCSiYyWuzpWzaqgEaDa9F8dCP/v5Crlo
NH/pD0jw9ItmoIW69PB/S/ba0PN9UhLwnpufJM+oXTU3u8TFHltWnmIfsN7EUbTB
fOhDd6oifHrzU07B276DWeVthN7lmvKUCue8l8ltGAZc84mRexJwjQg6mna13lrZ
8slK3ium32Cq/MgIRs0wEiIPflEBjXkiZ6ot6hCq3ioH+bZelWuybG+GIhArW7oW
EiwseFjA/kOoOofMDNRQKZTjrt1624jwoUgzezpHCd1bY0KMKnsskm2eoI1KPDcD
tGPv+CL2foZne7/U2vzA9FX3WtCQNaNvjnYUkV/bpjqSYn2VbqqlzcrlemkujCz5
MxZEsIjxfrBasY+/EDJ5er/q+plVNcrpMELAXqpTFpQIygs0dFXX+lOl+3hpSFMu
8nllK8kymb1m2m5xXDrUlv6C6FOjTIPFMwgAu+Wvl0SPoEZlF0GcSIisWrPyjDxb
XDoRPxOq6zH/kdW+i7GMq3hSzQTxHkCxB9kTJEOH9VKDX6e7VslHy8fHkvJpf2Qy
BK0tXH3b0Ga8Hf/xk1R6mquNZyiFXodhR0vlb6dH9XIyKKQlfe80HjiPzuuJ/Pqi
S8Kbef2fkj1E8SmrcI8d6Lw2stun4waMBTsQYyF2GLkXgcuPAhRasqx0vQ6f4Mpr
vfmNoyB3kP9xSzLht0x7FviYkvAhPbZUxYWKmmrF2G9goVoxadKqonel5haVpX7+
o/bKk6szm4OHW7oz6ywEwZzkR3AF78BAg3eEaPfmQ0CDnGC4U8Pv1hAWGyCXrIl1
/ToQFHIgydhcKX6asXMz7xrw7NOTa46RSjz812+Ogyam1dmArWXrB8yP7zhj7ddh
/nb6xfRTLX0+JsAHcAJ3988hK3iWXAZDqJYKDpESQGc3vT9e0mVDQjpHqNFk8tRo
nMIP33FftllO+yz5WXFMT3RhpQmCPxTD37cgWvf+dEYTvRqc5TzxBBTH4pzbg3ec
zPKjnpxoIFFNGIYuyHIB768cKi19Ag8D5SQgTR+GUMrcG0siyAbojhcwAvFMv6az
BymjDPdQ4Za3LIoB6njJy7rlTfBK4HonUFu00zho0JaRYVoQ+2Z0lqq9qqdMUGGZ
KMcHYTHO9L60iEhXWMGiwhmIeg0yqsNIhzuM4Q/NnoB9qWo5eJbCntM1UyHNPqpf
7gjBc+PyLXmzAXGXe+ANnDRjokuDSfa01JQyDEucAFnzw+/IR/SHhBTApAx9HQau
lOykiqENZdWYgt4t83NG26CUHbf/GBCh3A+ehcAJ+Acty2etwYQtek/dn3tSAB8Q
S6ZBPX/totTMPifJr1ZHD90GWGPyGv0467GnH7H1Ok/NbaqUKYARSiIfREBG3TNZ
2TAu3QB42S89IqgVOX6+HMd+w2iO1tuzp8FFztTfm7sYLOiv6lAy4oz/8RgO4fcG
ZbuHsNawpzE2rE+BvBQPm8hhKFZAG4kf+y/mljM0D3AqU/3oj+RyArdgNqB6kZuf
l73QSitGC+x/Hljnld/sNPvym72RP8M4zHVNjSSn7iS7yvfdEv9/aV/wUqf3KU2b
MK5rjyBadXyJovzw3yGTZgp92L0Rmms087gQHHJbd+hJKxK9PiuRMb7lbBDOKzZp
DKKJwlSVnemJDvImVJepFKIILNnQjw+4R0SSOa+BDQVSGVRSshcE7N+W6HwhLjVx
EmtzFtEzbn071Akbpd6Q1C77ThCVg51gSTS50cHSLIHI4z2SvTnEp+oBnqDm+igf
KZS55ryBz7g0avJVy4DiYKZm6kmu+b5G/3k0jj+heqC27gjZKEaN75008q1+MTOq
a9O4fGLouqeV6uyJJYg48xz98D7veBOHs/cGH9E+CB3EU4zwvLLapRVkle7Q4jVG
ZBd3Rl29pzr+n/YdfzGE0MfG1b3pR+rHv0FEg5CR1Qq0guAE25TUQ9ytPJ848jLX
InNDFN2QmhEV5nF+73jdxqWwSvBQLzStS9p3FCzjdB6h7mc9rsDQk3vnhlliWeM+
p12Aa/oCDCprixBM2t5/MYju5OtiL9bLUIj2NQ6qTeDLDskS4PmU2i4dAQok4+Wf
P/YcQkM8CHwTudtLhXQnCH6BDUT07MKc5gYIaW1zU7u2VweBFozH3N4+S5vL+MnK
J+Fn0E3fdNn+8lC0cNtN06dEC2bamiqUoXx35fROkBE6C90ghQKPVZ5awVTgfcIw
XT6Latrc771vCv5Yzz9/hITUHFccjgsLlTamK4yFWpzWt91tLm0jUc9TOsHjyW8u
SJkx6qVr2gTE71D05b0g6wf9fHuLt9SYwXF9u+QZQcQtpm/olLOJ93fQkMaT8GWS
e+t1otQGdPzq+I/ITQkvVrjwVCFFHIoEbMKZuRuzaOdhkzvXaSIFjtG3uOak+NDW
796/0X4biJWexU4UsH6cG4wjrWRoaa7XODnN4VoBylQqhvd9xo8F5gUTK6z6TCjL
2EN9MgTf/nG7Qr8nWE5JNmkI6FtxTrWL3QnbfaMagjgWOFf0qoX64Ve4c0WpUcMa
ooNG9KDR+a7LQlTs++VIm8HnrRJomB+fBeGAa92L6eLbzhiAfmrnJV3N5fVlacxz
3sGjxfE6lynkbqnndZbx812+LOsI647l7EM8qVTvrwzkzROBF/mj33QaearRZbQT
6g+bfGC0V9ilDMxznLq0MZtbBZXjIwgvzUTiCdzNA5afDdoYxaiOuQgDoYB8f9Ml
JNR2EIuNuyo8RZl4GNOvjfHYczlep5/HiE3F0Y6xmgkHqh1k5vPAmaGY9z+rJmSI
7mxWn3364HEm/oeADD/UE6gb59N7paJJxl/uFAbtrlL8xD11MDogBiE/Q0WsNkgP
nJGrWMGCQCDV3r7JupaD0Eg7UqaBSyTv1fVkFlClqA4Rn/VWskeyd5yiEUtK4URO
6sgbvOeowyrhtR3B/2C0YyS4L8PR9jZoyaDaKOIFIUL7rocrU5vfWQBMrJQuUCYH
rBcUYO33ImqmEZVNaFyVxLzI0jlX2gkKbQWE75ifOYEAiARYKtPZkcQKIkrm3Xjl
91x75na2R8dQx1SI4xyowi83K0cqzHgpBOieldPirk5Pwf0oFP54g3l7fRnCjiuT
NxmgK2MPDo3lUFL9ryDeDGisMVUe9+RbWSCtsb5pqtD6n9PzCi8uDblgabGtxmfW
Y4R4H0qMX+CqagZGkpcI7t6UC7hVEVTHxOsphOCuk1hX07k8JzQ8wT7s+ZiHEimo
RxBIowGGjg0Wo0B9o4K+mUE463gYLSuaKg+/XCK1PcHCTgTaf2BUM3BZPvX7U3oJ
YnHx+m0j66ZYx80IddtZNem3AaLB/lw+fZGsmCdZc840pdKScPRfUeS6fBMqwXpp
INhso0PWKP9KA6/VeFl35zibRGY+vmHglbBuF2RxJMElBYpjFgQ68OSxfd2q59hh
MVmzrj+b/Kty0ik8dT7ilH7vxtlifTAM3CyXRvPWPehncXSkOcS1GnC5bq0F2eDw
f9LU369g46lkcR/BOAy/gGbO1kDfaaaywFXyP9CBK6kO2ijYxIeo0DcPyBgDYJ58
tYuj2z+Qwc5YErN+a0O8LU0zWULMiMtQFaVeuBZmbQAhCp3XPGB3Pbv2k71WU5hi
aalwFuihh5m7Fnko4IRv9Ifn6kEUq/CCz2Om2s5hKyfIVpJV7UYtBvM1CQ39DGjC
mlZvgKOSisT/29PCNRGHdgdXMzSzWoYHMCJKLKZwAxQMiobUzDyv054fFVQo1eG7
9Jlt5zzyA2330po6TAltuuiuCw5QsZsA9zp0oujQURuKl7EKKZd4pNQNVUIpRPgu
prsAcu0WGgab4m6jxPRfhpMESoEBXax/Ka6+EtAkvNtQHCDdNf6zz5sCLcgdaxL6
tKkj6cKw4HJou5VP+3vYVErUE3LacRKX0jkkye0Lc23kvIkqnSCVGdjhPympdJl5
WQJ5g21Mau9dbFX/66dHwG9p1Pk/zdLEFx1NHhcJ3YDyUabIHr6fIBdmhhXEt8Xo
SDwJAwGPgLvmu7W3RCy34JgqnQl0I/QTz/0kmn3QV1Bk8ZQxWkSKKHFW6Xb0E+BZ
hGs2lXIdDjqYh8+HLD6mP5KF9O8A/QvOGhh5yxseF2bJd0z3Q+vGGtwFO5TsRqoF
ls4DT3X4F4TtA67FEcmhT3lDYL5uieh/vCdNkpY9FMZKjrMqbkLyk6veC9KY+lce
rEk86QtAhOSNOKYkzUpvsb+PoULJOTIcvmlPOAVU40B8fL46iDTNUM6ENMfkarV0
awowP/KpjFFUX6plY7PfmZzMYV7mXKW8AEOWsUrHiwIw7OTuDYdC/8D7QdG50uvD
8lsP0B11MV7iwu+XZmGIeAQB6mTs4vY3qwhHgmEsZ4xm1VBs02+SuosqU+EpTmhP
9y3csfTOqIO03gXaR60B03vOqANe4cGHHLg4RMth/W8rEwp5UTKVuHhcf7TKG6KA
5WolQt/16OoHjq6UbApsDQ2/YHKmdcZCdR6+FXrL8aAtn5HuJvcuj71DQph4QbOF
aNqu5O+c3w0IJgwkovrW4SIYM7iXrcoRr0DPsvD3Aua82Em1HftKDGucQz4c8WX6
LvvlEBkH6gttvBnukBS6GW6FuKytpECBE4NfVQ7OpiEUxeihPEEu/mZFl0h7/LXx
Om01UMDGGfzCT3y3zlGedgB3tbKCX3YskTGG0Ec2jM4SxFtDPhwf894Lk0/eHJVU
fIF7XEyU+AHnCvphlRuNsLsyizqk3suMC+gRVVC6O8AAkOuLEhRYK6WPgFwqN8SJ
/0kZZZdQQVdRl9jmEOXt4kwL4aJhFg/LxQwa9mX4lJuT5t058T566H3/SED/8bY3
bOlpVlcO1ovFTyu2MdFNNVm2M2lqflUB6x6OYA6PqEriKJKQEZA+ihb/6AUKytzL
++1kUJuZyj/gM82ZEkRBk7Mz58/idlxA+n/Jjf7OrX5npGrw5YLFacmYfu6PI21o
uOmx6KVmuClaVIeIm23GI7lTm+hDJNT/AM5F0oA1dbpZiSbRhMRQNdzrmjt1Ad5e
vZ9ZE99CeRFZ/aw35YHSziK3hQ4ssxSEl4mhftjcvoJ47axjGyQKWkWaruS2zCkS
WzOdcmtma+u3kFXOeY+gVtWZv/xWAcbMexrL/zEmnebxBptCn09vRySQEVnmqX++
kOmQVEODILmX4ozoehPXH65umHIZ/6MbW2++dKwp9hy69nrXiHzADpqHP3ZsK7ET
o6tTtY8t0cm/K0ULC4TS+ABZnzwToH9EAedCuM3F/R/I0U0S3CqNFBjoibl4qeB6
XypeGQF3Lt0TZC8xtsu1P+EmjpmX73iCCwld/tLwRG8R+8vIPdcYEul19zqLMd9k
oPXO9uq7fC/7oFlkmdP2v/p7Ttj7ofA+8XKqn1FKpLfF4ydMgWs10aZ08Z5mQqmx
a8vaheHKpas0lrjDyal81FBBYX8129zx6COPqOkmr2sgS3okiaBiQusJ3RbkQnOF
C4TFZ/D0kRy/BH84WpTI0kYpo19rZ6yzW45YuPCPjDTJnSzgPIbSZg4/99Bxlf5M
VlDF5wXgk09xWMkvEy9KxUxa0sdwjLuZwnNdrBU+XoUClV2cdAUygbRYjGEW3b6q
Z8xUG9nLKJNyMfkDlHN1w6A3IYEyXx2+J5j3ZtBVvoPO6zck1IiXU3m+StXEanVu
AfZRItmpXZY3pBFSMZBcYoCmWm29FwHqyM83Jvk6FA/8nfOZ+xPI0jKoAWqePt7G
Ja/8QBp3OM7ZBUnjmzho9lEqwcpeVLuPFgvqnkdP1i6tnbpDkXxjbjTmdh351WqC
iLjq5iAkiSA2SoH5ax/TBW61jQcUGHR99EbLNquTUtI/VbdHEHUGH7qwRh6vhBUg
vwh8APJlDZboPwJZbBOErt8tm8aDqi29HR8rzQNhn/ciOHV/txdF7OyY7sA1LU3t
cbsEGwvSGwL4J7VMcDXW91lrPYJT2XbF4d7O+jz1NcAsLAi+cfu60/bHPsDv5dp7
fBy0RaE8wvHwAJmDrqJ4aefxWdWuRp2R6kZtiB266SSJy8oBas7JFnvTM2aVZeDG
jK+Km9gB8pgVK43itWWubsF77oM2v3dS5AECrCxp/kZQ5R0EjAOvhzKqrr5QZAwc
I8eJy5QIVyLyFB9vY9C9KDCGd8LXullOBBfhghbAOJzWZl2GJZSs2yoV6dX+QElz
92oeiRFy+b7RCv9w06CVIfroYea3FdpCiRqDyBxs00BiE0NOsp85tvQZyyz9+vCu
4Ew3Yk0bzxvTLrESnEM5U/X/LWTMgyA6qpC1NRFLW0gx6UYkhzt7D6HAxlCCgRcy
oVzyCA5XlxuXdHCWeveIsc8K+l4WfK7GyKhg8q1Qons2AStXU8GBOMT/A+JVPydY
44f9WG/g10r92MxKSP8OQ8hEmOMuDSjrLopCnSuhZv2S81rzP4gU2bEB9oLZvfC3
QWm3IlXATlRDq+i2GlJlrhcZ27n9UTXdnjO5JCneZNCPhOt1d/Gcc36IXhpsg65T
H/sjFecRKTzWiOlcfFoISVUjb9aiCLkTPXJYDaljwaR0S17ilcdsjsZGs3Fcs4Li
C7wm8HyR07SyMnS2DVPETNsCXiPvfmmZuqFP5To9d2VZmMmhBe+2XojapxxQccOs
5bDbYcFaMCYzZCkVCmPlgPnOCp281iyxXDXcePolTum5UM+d2wfQL6vtU98yQtrE
I0AEmlgELkD+L5LoSMI9t+gX/z/8/UyvbLfOhKgJaO3jMxU38+B50sc7KBmnAz+C
zeQGElkDCKpiIWe1ts5Ogt494tCUuVDgCoNv1Sp+B52yxxXSrVIzUps8lFYwowzA
t9zlgmQCIv8bh408DME4xETOEL0zXw1ZCXx23LLdZKspAZBqHXOgJmQSl9JkfYqN
fw0tN1xdQj2VlOEm+L7oq+HKcaKXzU3qTRvbYPmunnySgqlHc7kW+8X6mxIdcxAa
TeoofLPI5v8avZAz5gXrHQUD3BFdmHhagmQ8GCyEmU1Lh2lfPlKA5x+B9I0WNhYO
c9knJg1c5mL/x73FYbqtyLJ73OKBW1EptoG6+kFYdf0a1vy/2kAGUCAeaFERzITU
KxlPvAUeWNsqgwEyxdhLaA3FEKPIJOrhm0oeKkLsHDNKxWppN8/rcw+50kdYPnB/
+QVbxQbZeYurqcBguRBqtRbtXxoWGxVMT3Tz+EmlYsP9wsy7QAt8kKbMJR5AY5lr
8pnqktbeShOWITsnYzbEtgmmhXo5XNuZ5WivYxpt63KlNqOWM4+w7JjZm4GRr0wN
WIljvNKJOh6v+05DwZSwelKemfWedLNymOj0UdQ5pFxyMdaqSNVQSIR+bXgL4EIC
Ol3dSvey7JCua13aDqw4rqMzfUxYGQSLEvohxJ1QAsVygc6ePHdLpU8KR96QQi1z
qDIqbc5yhXpgvOgm9mAcCdzxQk/uBcdCoPqh05PwaXkY2VXdkGIxTxM+DLOUkBZZ
s3uSzDVDlij+FfZEDeye5OmDl3BwbwIg6U5H2X5OdT/Sin88Td5r7vUbdtaorcrr
ukApi/80E0ABvz3KTMIkAOaeWlJvsaG4p31ymK/kmVkLArecX11itx3CrOdyirPd
CO54DYD5t7kfVrQo5nRglRlYd8KlqxT+dm/Qhy8YCOC8ECM4VcVehf36kNU7ncyj
Ntytd2af6blFcwOKLUSoXPDtga2rSJcULGP+50EThNUVDOrsilUD4+GTAH/y4Vby
P5yoHXZ2l2vQHc4g4BPWOl7CTpBC3KsCUknopIRCAOoV1/b8FGaUBEHdRydCQFQ7
QZ6pzHOMLFcr6H3UziDwHWj+CPy37jwbE6OZ9kkSvFBmeSnFmPmqqBX8p9cANUpF
+UN1MEiBvIEgPOHk5uBMfit5M+dxO3P10ilv35ZYMwACJh8F7iyf7WVY4iMYnY2G
bXkqhTeZQDRG6KK4fbjVfJhijnQBorlq1fgsNpm60+lS8f6Z+oEwdzQ5MnAfbYX6
Be452e7IS7GSM0phk59TgBO4tGIc41rnkllJgj3IpAeM3E8XcjG1MjgROvYOZEVS
7l7uAgHLE9xpW+P8T77cPbys5fZwYj0OBn+E1UpaqzaUmmThhE/I+Zj6woR0nQE2
mMeDeyhZ8LgMnQ2Xznv1Fx4Q9UnCEZldnJYBMghHJFa7HlrBSjgxu4BpErDY9BEN
qDAlnnHmEeH+BCNieTPNJYlkhRpg/VKa3QzP6mf/DrMQcpilBflFOO7O9sWPkcVI
Eeriykpq3SggUipotlotm3CA7LdxJT3mI7h1F6Z7iN4eLGr+Znk1OWK89UFx5vXi
Ov0TyhmqbrS2D8LfYhJlhsoJArre/QpROMkJSx0/8FPXfzEGBi0F/zHT1qvPmNjj
LGJbHPqGUDKVTT/9OPjVFQu8oIDY9CQXYFZC6YNSmJuuUazu9jgK82QlScIo0Jaa
8z4TNUOK831BN/11ahdEoQlcLZHDZScPhXXBvh/WPMNHECYEVMoYO7P0QKfgkHhR
Vpi9tZFVG1Al+Dv4sZiRZJJmhh9K5/x0eHw7xkboJXMsVugMX8/1hMfRHs9EAWUE
tFo1g6asc9Ozo0a1uFSg39ti8JtCPm+lOOLZn61ZGvpjF71uJDXQ0/OJ8XlyLhGA
pzW9aj5kqDGgzjVdNF6vD4f09zmaFDsRm0whSeFFeSBfzfOhC1DpVyu7pqGF1lPm
FHXzYEJco5gPhbGM7pcLQ1vphnGkFCRHxdAskyhMz1XRBc3o+Ay0azMqkIufMAOc
/bNlBaYgxzoIm07+DnoBR0F5PiAXw1p6hVE3RQ3kjMfC/QY4REOBUpGM5KKRtMpw
qcfZjHbFh/oEVo/Kg8OVZ7G8DZ7+VysPoo/BldYlXd7ovXBGfTaj5J6TlOVFkkvd
v9KZVzUT3WO38+g0+5Mj0sv7p9usx1cKhnyoIzkT9aNsnSOrFyTwMkQEQejlUPHL
1VZCIHI5fBEBHyP+EWoIzTxp6KQ4KAPDaksvhrb1QA08eeoeVm1jysRvHczo7L8Q
jN8RQuQQ8DL2vofs4aoUbCVhL4nM8jFbgCczARhNSAGBpi2goAR8besjPCLdnUZ9
t8IL8K7xFq85gNHXU1YwFRr/bsiZYerVZwjsduxrc30lMvBJ+o5JA+yOBESYbaW3
/VC6yLehc98EiuJ0AIQB9H5waANbTgjZRJ5uaGzjY3sk2kklSuxvRf/0zSsrGeOw
bLrU7cSX3xEgKRc1wwSCHQPpW9Sd6X1ytR2iVM0Ph3IqsW3Qld715kT59d3UpfsF
p2Ul4gqFT2oqRKc9hqfO8HBPVz3sF3RL9xS6I014iwHwUzmohLs+gz4Ak9n5yy8B
MuCh9h9AXUKFad9RfjTvf7ovZb7uxg4Yct3rhdIN5PhHYxnPpdB6S4xW90Y26BTi
NVm4J+inDBTgjN3AlROYbiDJGQbUOAvRyrMslP8C+9NWo00UjwNXC5VSAU5P2i5S
Vj0gVwb7iJEMoAO88XCYijHK4tv9RBjrOg0Go7qNFk7ZAwKz89GO0RZMRGK16+3X
NAMECCmAf0TveiUI0A+RwH9b3O+FTwN1Br9zKwM3+NCYsx2iw0A4km2gyu7K955O
tlmw3KFEr2P6lH6G/nY08rxxschMo3QMFPwM7bTQBcm2l3jGVFW79Z3u3HxG6/fq
cZmnLSknhdD9cCokPw3QHoJ1kmrxBJqmCaMuqk2abu1z0TKLytW13Q3V5RZzMbTK
TIFQ7EMLFDy3Ymc8YS4DmhjaXcsM1Ie8QdpRkhTek79ZUkp4qpizLGsyX0DoOSR2
N6EySfJzxNOnVEcIBc/IWIEiHaM4jsSjMT6d6rELI8n5VwkKNWNh890dhZmA7jFV
iByDO6TyAoBUKd0Fvw/EPCR7TR6DPlz/RfPp07+LtgVBk4AGkgZd8J/fq7K3KkWo
SlnQIiO2eDh08og6dW+SjW7ISiAysdNsUVeioYLTfnIFzyVt5nEx6qLuoSeOZ1Zf
vNGQezMTxKcQqPuNWl6j+pTkF+dj/Idl1Cu4XuWqiK9Ur2zSJGD9lLa6s2fqwDDy
h9Rq0gnZvhUiWBfQLBzaU6uS05fajPPG35rUctbY5WvsQPl5+Wdu8ajCsTqkv8cp
Q8bS4d8D6Yb+Cwk2mm8qtMrGnU6/pCSdSKytpCmwjPXR1z3ixmlwl1p+10ITs2Ic
v8TEaFwQz1YElgIoZ7URbLNKFcXVX9dOQG8yWgbDqrfxgS3An9w5Iztm2VQaBLQA
spGTAcReoNpTJc9kL7BoMAy0BjHMA4u7KXb5BcQi776+uQy2LY/IlF1sfDrZpkBn
FM7vc9B50GD5jTuEmNbF3nENQSno4as5SUSk2J007vWMHxCW0jHUWcDv8Gk6wkwU
ZTAW2o/espF4aKxZTtpoI5kQiQK0de8CldWFdRa5HNZuYS4O2oVaUHoaj9TGNFBf
fAQv+H1Ajoqg7uoEv3aV/kVw0DVOPZmP2AvzbK+GjlVddFYcs/lb+aPsNAB6Ffc4
oKJ91AmbhAotVR2CQFFhGMPEeOlgxq1cO+mIEOQHNSnOl9DNQeluRDBp71NcGH4G
mC+SR9Rl/v6Zq61JQlTKT/evR4Uw8QcVR8gJS7rjGgOTUcVu1Aqeal3Rpfm/qcob
r6t40C0W5fADaMOwfmu6z4Kx1TMceNYJ5y9dLVkTE04za6OHY5aE8LakPuPJtSpj
LO/dGQjKGUYommTre4X+n6dI3QYSFMlXvO6apD9d2FRkT7KjGvRHFCDOrSDMBqGW
QVsa0PdhDdt8SMCsnsRJwb2fIUdNdo42P62VaAKi1LveArnyCuKmHYuJqUfQKk5s
jkcCCE5eJci2fY1aagGqsB/Z/LuCprADJvmzeJwNVMYiX0TGAZHJlhUdt+2lGbyo
KTA7a6pUxG5bNbS2W1cFizp6XGg2xrhPMdiNZHD7J4PdFGkZnf1w9EQCJEAcpzYZ
CH8NBU6nTJCWAJDL1BV9J5IwDQ5zu8mU5CTH0rZmFb4DxxXz780OgonCOFcbxRc0
hrDfi7Sa3IHGkwrTQ8rsLEFqPtxDVklYrdSXLmL4vEAdibpXqkEgIkXBPiEhn0Jm
8fRYjUf8s9yweEe0fLn64EQlIiW4cAEPLTW7d9lCVhTPn5UejpKRJahR5QBAHmVq
h4c+X3Y7COLV5/J/ZYUyX6eQAn8TReAy2LolJEheN2jdG66GREmZDRA2RRKSCkMf
YNNzOpLL3GQsFKn3Y+Opu4WSXEgaDXxkqs0/V81YLvgdRtddn5Xwyf72T5wauUT0
PC/G6rOj95d0w7NpbNnFmzWA2jnF6ozbEWziq+sqYk3QVLnkoqsJXv03/I+TeVi5
EXAfR9DcbiyzeUYwqmzsTWWU2Jn3ZlBmmBzpLTelfY/E3HRFsigc3GEqYbpIDRaO
akujQu65ni3iaDv23IF6O9+LeLtWGbJvcnWy+WupxVaC0pgCx1shXU8dp+xetOWg
7PJXLFxqLLx18U3IUVI6JSPQvf6AweaUgLfunSCA3CBhaZgO94ygq4UXwSzYwn7i
zhPGjADM5FbAD7YYouCCEeX8aB3i3VrKnQlsM7WkwdpRbh3Cg85+YbGIQvQzQ/fV
P5KX1aRGnjyLZfbwqLArZmF1BR1xAD8zGt2/ZHo/z7LzvfbDitHwC7Ahxe7V8eK2
NmoHepFc3iaZD4mJiDG9lsPvHmW+IZyIVDYOaHIG8MO92xf2HrPIl7Y3S2EzgRTr
g6YeaFN1P2JnVAcXVpOSHPTOVSz7vzNT7/f7yvgVbO3Qw3hpSk8lg1C2QLuVoiGP
7fIJfL1WbQTb4ZMBYx3tmfj6oMcgGFbGQL9XEW0GYRJdZbT7JPq5Ruk3kTIHkGSW
HpszzNsEzv/dyuHBCktQTdhggZRFd9J4iPrEoNZsm3GKQNe4pNykKEnbc4Ie6dVb
LKFX3p+frGNxk705F6VBDPKmCxfzT9bwdmuvnesLhQIlcPl6X7rwhPbQKCoiuL5b
l89nzU1v1RQUbOmdE3u2Ju0RVx2qKLr9yZPmppQ3mcL3OXJJk7RlutGy6LT/8Sc0
XFV1iRcA26yyX7Ze4PtP2oUfbiai1jkdpATyi094Y1yukg0TirfdBgerLwFFrA4w
Zpn+mRjY2qHFUY1h40zJ567jzLwTSAtnzECCx1Z1MMcfq9UThelvY4fjizNcW3oc
OeHgtBbyQXZJGGbN+ApBbnvsjq5EO1qB29VtRQ/rIKkXkMAkiexbPlSC+UjSs+yz
CUucQuS1n3o4DzcFBUaS4RZ1A82Wnk3E/pWLvPggsMcZ3HpkwXOqwqN5zAUkNyE3
Fm7fwsqVyUzeeoE+jzqJhodgsSlPHY+PQGdjVNtuVnWrvEfageS7wls/w94sfY88
02H2/As7QTYenvGX6tZXgGkE1fAwwmbKNmDZuG2adQdKLW/HlC0Nlz0U6iEIHrzz
4R3e/ZVQMM5efnFpNFa+wrsBdThLshP/iJfOnKbORFm5BqqX+x4i0rCL0sbCGh6/
61YSmKyUXdHdb6HuZ0AiZd8NLIoZZ4cNYFZTRN5ZkzRW09FegOi1dRWRZSknWIci
vse8f5scQCTdQwxA9YciKNBwdRL92YyjQzhju8fi0e7RTlfli+DyoNGXdqpBH1+A
dkYddxt8f7T2bdsh81SDNwdvfu6Z6ajdrAzj6SzuL+rrxkBsf0/Q4Wx2MZph6RLn
9C945y3Oj0wJxwsV9t5GRFU4al+g6MgKeutokfsQFNEinqIkQsnCciuwBLJUyio4
NbBHRFDV95TtQjJvvZZSSkowWvcykzlUdHLM6VNc3BLNa5u4fu19KHyIYlxvuRND
jNb/nGgFeAEcazIsbdpQ2XixEg7OPAlh/nhaKSz9LGoaLNb4nV+23lZYvVzYaCxH
HhqqKOWUGEgzlY5/xFYLj/lFW0pOGxJR5QSjt2912vXDhAM+b5RXR+dcQY97kSo9
3dWG+USsERQHAi/m/nuXw2QE/wxD1vBWTZJuKO62rCsRyyQIIIPHZyfdgGyXWcnW
XlYYRMDUgEURRUldiUA2SnYEKsvlZiRH0Avkh9OlP6wJlpzpPY77FNkOhQJ0rIPB
vyUhGvlu/07/RxDMBROhJvenVHdXHOPNsfuuB856bE00kKEVUF/MbLiLzKLmlf1V
FDm7Y8qn7bYh4/AIC5GyddH+HpxKdP28asPTDclY7f5Szk9BjzrrG1H0AD7nKqmR
wmm3gj3+GXBntCFQPfGCV97f36W/O8AkQA62pHgcqP/UcU73YVJnKYM7mNEXs3bs
iTTNpzIQTa07LXbEItThPLBn6/jQGQX5HQGvhr/L1nHJDwLOHanO0xkoIN2WfTRq
GW+TILTwoEUNcc8u/k37+Na+NJumV4pxVwOnASQ4AVJj5C1Nv3KUIfPW0E8+SvyV
F+HOFcqwHTTSgSRyZKig8Gcepn13y+ccD9wDhpwa+t3eej80pqljB/9/QZ1lR1sy
imHkuqxvigPO2/zgRDe348m3GXMqPEjmWEEFohUAT3jdpirDUA8NOaW+VbyIeyz1
GQMe3EFyQIxP7AYggfTrXSraNA+JRtYfRBvgjQwEGkgskoxZ91hT1S4koHLwYTQx
ftQq9ccxZznT+LYb9IHT/emdeeHNFa2KRssRPBnUT/MqJmVdxOQvtRy0eHPstDwd
HZGRifleAaNvOWlLAJ+oScZbCQltGpCmmhLqBT91s5KplxuG8Vlnisyo6Bz30B4W
Qy7BeLSwKRN4YZ14aFJkmsFWl1noIGoQaNhr1aJe/Mb09H5dRFLKlD+5i7g8zn/L
7OUiEGQaFCOCnLLLRkAgGrK03LRa6gbnD4VjNALV5j13GbpbTN12FwurzD0RpNuP
w9WlVWkJm88Tl5w0j4Snxf/e1+F/rhokLqUg55kiRZ9xing4+6jbpWzu8zv3YYu+
tnUBD5l0gqHZ+si2OXxG7zOQd4q31wRWmVIVqatRGq62+3n11zUAKdkfUj0oGG3s
ZG/3eG18YoxwCAdBDS4X0i/TF/xLgsParxvz+sO5B8s0Ja5Bs873Jnnh0tFmmx4O
DIRuWusv15fwrZZtVnKi/6z7YDlrOVH9Z9vEytSlkSQuLlfQqdOUFWx5m9qeZC8R
KqBM/WSdCWS77SqXHn88eAd0qreQVGRXBtSn4NzHgBKgFo6h9EBsmUivUP7LX1Ps
J2Mn+Gezh8M9gSgZmPjfEfxD1KycGynHZ1GVBiqTXZcAQ1EhvS7dDD+jCkQUqUFB
kF061BY8lX+Dh8f0U8NKDuWIAi6igSuNPiaDy2vqTs0NuNCfGG/MHtZ2Ma6cP1rw
5wVpo2JkfqbWQiezLEoN9Cnq6et7Ob3WlEdsvhNK3QKMGswxAoEutV5puElheGQM
l3uVnM0V1bZuIhGs3ffJaYUXxHTZa5YFeQcwvByl/Z97MGve5yzztWMOx+BJm4Ma
vGP4/xVCQ72YtW5WDTz5va6LIsu43jM4A9zU2+pC16sdStQeSgO2P1MhFKSEbZKt
iFF4PbOB2FAxYN0ZqlNoO1ljw4QDmgCv8/eV2KZtKLDng27/PuTuzBh9gmLFXnO0
KNC55qjBjnYyzF8r5zbhN49ZzmJGndS2choa2IXQnR8LCRTQNckx3GJJ5wWNEQIp
Oo194+Kn34xSLbl8F+Zjxg+QExHn34HDUPtdSw91miYiyF//RPNxHnAdtCHun4bl
obVmz0jwMNapjj6vVhYXFFNrC0HzblXGUCDCOO83uMGeRbsLlnxleSBoUillSI27
psMzd4ndpTSrcasBD4YJsf6PULZN0yO4wEqRpHdFkOsfZDdZz01VfE5TJkOdGRVk
97PLfFNbe9whDyiIC8OkS7w2XTM8pEt1LKJXjiCN/Et3iduPenkCpeNMU8P4Frwy
6QmY0AOK7Q6FlRh6v2XEawCJLL6oTS3RB+CPLDH41emW79dcPHhHngMxjBmC1XYb
efv2maqGU/lShQ1KobtZ9TucuPiYW0bEuhOfI2Y5SFuK6V0grM4NWdhDnY7zJu3u
wGw0zcvK3lyYwoa9Mra9ut3uy3Ioyh++F8nw4XNt4GFCO2Lsu1Lf+e/sPtMyME2t
IZ8xO/Xg2rCpV7wOR1ItIgOrf2NsojpJiowv0Cg/o/LFQaDj4BJEeAqK0CohWIh7
Z24yCcterap4kHrQcLeVSZT99oFoAtaNF9QeP6TS9fcyCqD1szIk0KTSMHO+Qbh9
uiKiqkyzV2q+LqwRKcJa2SillXxYi8Nr1taBWd1gP2SxtdEe4B9PrP5WEEMFhJhL
SXL/lJN86Cin+/GsK+vyHlBRP0FcbfytxomqjHH/tZhDlmMY17RDS7QBSZMjuzqJ
yZ5wdalvR/5ULWQN+Lx61xo4Y+Fj1qCXOYgGwheONRIpz0QyVMzbc/P8eXom+Hrv
mMuWUzfBRT8Auv+RTFxW+ss4Dffc7SdlrFEPSa22vrZF3LMWwI4hSYqCd+HddcSk
eDQbg7FWDJEk0ZK6NdIKsim+km6rWitkE6uLKqC9WCa1MFHxD64fF947oSa+8USS
qFBYdNLsDyjZ7CiKPTTmkk/mBVLoyhQ4Oj3iDWD998PaeuAIZl6gWfCGvM64cUow
sQ7q4OqQdzlrCPZZUnDuUdSnJAiGhUMfyTC2MWqbrL7SINvttw2u/P2gRN3c4ybt
X/nlaGiSOzu0zTt2jqp3AetI5iW7UXChYJeubqbjnEvQU7cUXnqRhIXzN7eaKG+I
0Wk4RBBD+QhjRzUqUVizrjr6NXYAeIzr9fWzyPa0gszYjH8cNm2DBtr3FtygoNc/
uZDEjdaHajhXr3rEfrhbbN0YMc/fwf1TR4m2KlPLzOWnmNeR0EIn6/sTgghdtECZ
BWBbWnMpq7sQLCHHH1q8XrcaiHyGkLRgaFkqtJrRgxaZRh8JMdMTyP+MvxlLzOO2
hJcuTm00NaBOJOCLny4JlEAc5vF3Fman40Gfqgiw49E0+PsyPBJ8oKbKcW8XEyU/
1JbGpEev+vuPw1UbFnYUgC+faudNGFfH1IUGlyWsG860059KAJmuN8+zdwYDAkpQ
19++YlhASZc6JGRywtd+QX32JWy7pI8PVQF6m2siLG2ddXRg2OILXNyE0loW8TyL
YUgibGFubboLUXDoW3Fs8tuOETVyTAwtOSU10ISaY/IdsS2q659p3uJwgZ9ZabAi
1r7BPxeePLsRY2hpTZjyYpbRZVU0OS5xrJGLgDKHOvV+D1V8S+YFImXhPGyremlf
zAlCl8JTF1XYTL3Ow48wlyrscCYGcCZ+XUbuINISgYKAKC39fMREsp0Ab1ARz6Mf
tHzBOocfyQv9B+dzwApnQPpDuxlNl6DAK0i5D378fxUTcIuKxUfjdpHo8/yuF1xl
kBZDQJ/9lM2TSRh+FXPdxF+8zy+CPFQHojS6VLfAQ7K8Q9G5+zalYVY+1ntdo9D3
HlqAeB+2JX0beXziFMFoq63SKzD1tuVl9r3KxU7wqdvc9FzhuEk3G3HXG0BfRDOV
k9O7Yl9c7GFSuC/r0xr98P+VtcmeDHpudKDN9Jtlc8aZDlryPPrqZZvdh/AyG/9a
p+jmFL62UHEkVnezMEYybmX94Wf75onIh3FG7nnmRml5pmfI3/Fhqsaf0zBHIU/D
JO3hJKfMT75RDtLIAfMVjf407JQYzbiaF/1ydN2LC2ueck+jemY2yQH/NjwETZX+
yr+5XiGe2b5GgjKxomAI0KpOwTdwSTNxVCuDtPOIucGgyNRuh8OWCEF3zA5gdZWF
phhqcuNkJSPQdM2Fb6FtIBBlmvRm0mrRuQEFzH3I0rkNgVab8g5qI72m5BWdPpCE
wxJq28HBlsd61WedN4S/HZ76hbRUg2PuV0C2HnH7lJysWiI5QxH64VdUZsIEAd/C
9REQhBi3Be5KlkAqEaqTA2JuYAXoHkI8IYqK8Hn5weAnqxbbLpKKjwAuzPnAgBk+
npy8qyN6u4kK3i9wjuDCbZS8AgIIMIWxfDDyg/Q2KkS4IM8UwcuFvmPEIu3L/LBA
d1n/e5PERg4Fx6gkkDWdLj19PehQuZ9siJnUZQjiI/ujMK9Jm/XFBnDB8uEublH7
m+xe+huJ2ZQQtH6nP43HPb+K44ObfcPbS0MAWWZIhM25EZNQuuHS4LY9aUvb3/Mu
JUBJfKsSbXOehIlnsgptNwCC0eDVzO8oBv3bJkvupnU2F36eip9BBB3T+gcDsPEg
6MqPdqYM0wQxZx1uBg/74wapAkrxBLG0T7ILnSti1cTXyUIJpgQ4oFJFDstv0cC4
gdMRbzS/8ggxQH0gIxfUzZvzfeuTP4wRypQuxIJCL0SkiE6ZYn+ehrx36lXwkseg
dAZ1LBkhgdjizNWIiyQi0QEqrgIU3ekkb2MoSFlrRIsp6rWtWGuWAiblhYXpkgcv
1amoPMe5PL5hrxf7aVhKnddF6KAILox5M8ZW4jsSXkRBxI1rvR/sYCWpftSjKSov
2BBRD7q0koJwYrBMIiWHq6Rab7WJxb2e8VM3+NMQ86/6Nzbrc6Vjpdc1Ho1W337c
JHq7m1EOsyMWh0brNGU/vLS7IHsF9CPT14shIb5fUjFuEztVmWkw8uFjNKWn411d
lFt15KbZmNcWBWMNFkrSrJy8/uJU2hSh65LRDsw6lf5DCT0oZadwr/ybvPw/13pq
BWYWaZemv8H35aRECjBGI/3H95YHK6NM7R9GKsuxZOMeDl/f+jgka9/ytL0cWk+p
7qLy5Sr7yK6gEH+hsrDIV+O4RccC0bvqDQYctq58OK5lQH1jvnFbWGb1Va7+Mki/
2x3/W94oxoHldz09EreDZCyKtVj80p5M7K1A2Uv10xfo8UrRBHdJUHXYkx+dqkFp
g9QXl/GTtz21ahlD9zqg+aIQR6yDlQGi0YiL7Gc/bV0KowTB0GGgW2JCiIhZEzrm
WXxCu13jBM0FJdoVXLnVO8tGikcJs2nK1esLd0DBliyfPDf/XNto/42kL8jwtlS/
nbwC5cHO2vldiJ4Sp4sbSZnmksmpY0atyu7Uy6FIz/rtwKdlKcXOWpOB2Q8mK6rP
JZpsOQPrvKv739BMSKqIL5PDK3vlblVpxtZ3Dpxla7hfvKUODlvmryd83ZienB6u
jTxS/JZnM9o2xXeIUk+YdDFkH+hOQFV5EPZfam3bUDcdoNaz3vTmBuwKRg3/4pvW
qqegLdzSnMi8ZdDnMZfzlY3y2/aClYKbWuVqnfUt8uW7QdMndMs3g5yTzj4t/7EA
74ypBkf45AMQI10GuYk2ZvLt9UgXqgNosC1lpbWr8gpCGk09IXzRsRD+m28A58gh
fuKCdDwjQHU+bF8wIL3TXf/PSMz04tNorlo4Boj8onkvOzOr/uL7RNnoNmW5BPvw
Qai6drZ3IQHdD2BfTIMRTu75sWsxwK7CBK5cB2VWfUcWwlhi+mlWx4sMdkZIJM7r
jvLRdeHIV85s3U8COUfTV39I+n7ok24rvsjRw0RCMK6ZzZzFbXa9SPXiiKhNDOZD
9Oetq9yxvpoFZpfWkqoSi8ccPi8dyZ3HBf67Zpo2A5y9TEfmeaGh3fF0qAcgZi9V
1Dnt5i6enMvvCWX05ECCiShErinGE4CFxHLYBrpc/F5W5nlzCeGFB1Nk+2PUq+A5
LokxTUDd1xbP46uEgPkgrGXNOjbjU45MUzlAV+tRSU/e5pPczCQ9tjF0pan1h2v6
Axm3WwmGM77JI4voBhKD2BeTGSyYrOuPmmntwTjk0O5jyQuVQesDVRo4tnPNQCOs
eZstGzBEBIK4Lofe/nn/CLrBiVcFjsD/hzzgZLwzTW849d4iZrkTO3YBMSb0GZyD
fDVDJBdzw8l0zaXM5mJVpuk5ehfUbrHBixUZqHguoetg3107kkiyRzZs+nfkTCP2
PTU2JoJjJr+ZRQCioo/fRgLVIl0i25H6r355UiTl2zwAMKVjCkk1TGe706+buFCP
0MpEB1dvGz6Z4TE2uPrm5gEMpGleXbxE/qO9q7DJhvw3XHUZlKY2Z+lEooQ2gNos
rZe7iNrh/HX7oQunSl40gz9Yhoy7P2Wov0vOGn7iNB9MqOiaTqLk/660Z5/WUbVn
Eb2Lj6RtAgcp72BCfge26IEVsSvu058Xo7pGwNU5JEDIp0oojFstLeyagnDEbbuT
Xf+k4/m0RexsSqWhstXmr2Mer7N591U10V9jVMJSRGvWnSLAoM8EOdoe08Ggg+9V
nPLbppdd0wy8mxy0Iw90677rjEtRKH7Veuny0v7cr/HFfplIXqCAsYNaY7RhZhUH
SmRD6TTIqptp92wmSYmwPAIN+EtF2IK72PGpbHFTF7hc6WTblcyiEM/oEuC7wtBw
b2K8Hllgm3C5zkqkIBUZHxuJoHdpkRewDYQp6U9Y25GAKfa6A3jLF1zQeH0lJiqi
fHngRExZRs/PTAgjkAKdR/zPUf/hb374aZ35x56ekkIkpM6xn4OSfp8/LogqKo41
eDR//Qyhe+XDbntpiauuZoTFcJI2bd4CISOJeKY2CBpvJnhiazBp3Lc+rS5x88SA
aBdcNPT0YTGomfdutNUU7P86RdXNoS59rNIOknk3qg8VhIbjwmePovFJe+WQ4Api
kKG9HXvzDcU+bNIIo0cT9YQMQqyPE+2mPqlbFNpq1jvGU4Rc59DZPnONjWM/kf2h
JKsKJs+7N8xgJ+GVuzHVdUWC1dp0Z3y1GQqJiBKaP+gXLLGvLSGvNRlLeMoNRqOq
2/DHffEox/SYntUICVU/jnZTUPcSwyqPQi9N/feFD3tOcs46NvTpyux/Oi2cM4KX
rsnA1axmxTNWUY6/8h7U+hALQqhwcnctyaV8bhhpnHwbLCMJu0Tp8/1J/h14q00y
qfOV9F1QBG1PIev+Teriu71YPlHSKGlI/yk0ME6JQXC7R815NwgX424TYiKTrISc
mUTi1vHQzu7blUTCU2eOo4yj9+cgk4ZnwIVOF4RgkUkOAzsdMyscaycVAYCljVPN
NoHdw0Xgf/LJylG0atk6O05rlJV4LoJd0TM9naXl23N5RFge7XjGuORwFbWt8rr+
Qzc7MpHJ6rTfWK3SXd/YIapFT4aFFV2P2bRu/y2bvSHGfBEQqZvEpNaT6ImoRbe9
XSaanLe19eiBLaHYB0vkRfgWN36sUtqxd+jRBoOaimmk/qesGyFEPrkbihAX/TYT
1iiNhRaI4Im5AvNgcMTHGk76PYppHJHOB3bjF7F3yQcXiaLFm5oeENjC0taaJZm9
8a09qMfG/9ldy9tUQTUCMa8uGWiABzVXXyvq41aPAE1Hm1FWYAd6z8dzhI6oMa0f
CIRglenlbGivZBLRoDUglvNX6h4IIjORoNgw1dLogXWFAs03Qhs9TiLxzrhLHYg4
IUlqMrN1oOe7nCZ0K8KqUmX4pLE/lyr6KPb18M/9Ohd7qqhJmT9OmSnDWDSkbd7f
xWkAE/wAxBEdwFa7ZnQrhi7+Qwf7Hyn5sa97PMKNSlCkkhv9XexkHJuQKFPgCWMX
c4VPR252QFijfba0wkC1ffjjX3LmTcIUqEhwfOnAyjCmtZUUefsktYE8Xl1eJQyg
XGE0JRImYfCwkr0IvISyThCH4QQ8l8MKde5MbbsB0eqTcsIQTLha8LzzQAic6WvE
RiEiRAlXjjlxTehe9LXqEBA3AdEjubY0Cu514md/HU7y6BIL/JD+l5Kkp4QQLbzj
RBl3qt8gtbXzGQ5/RU6wY65sZXglAeMIFOzrbmU3cLqYdc/EVlI+zgc/uWA9kkO1
Nfe0tnqB4LuR7Pcp7LCuYZX1ytRBDMohx4KJroRF5C4PSSr5X3FICfYiwLm3FpCO
DuT7kit1JxPv+QS6RYowbREoAQbMpVfjLoMbGyUCqFkPj5tQzSThZ4kvi/O13fgl
Mx+ROfMnKxhmJ7pv85BYHjxtq2SQsOHmgcoXb/d8jFBxDyf49rCzKsrEPoi9VCPq
pgELjrVhqqrk9d+LzVIlqYqTAEAty9l6g3PyjAvwD592Vwl19GKdpAtk4CjaxTiH
1RCeMEvgIqzMNh9fuYGaOguDYGjzOgKKcjVLvCNxQsGFGYsasY+HMq2IutWtCuDa
c+jaR8rLq9fSCKxQXZBkOZv5JaMEzNZx32TL3KyuDVZ57RG/ZF/EKIhumkzRNPVl
na4Nw4mFqxygYkrMZbHxfhryuZvFoIy3S3p9xVtUpLTcU8W0dPQNkD3nMBNt/UDC
HWBC5BqMdaxyrR+W1nf7ByEq09yPQCSHiX55LX9i0KAjB2eRYsKa5RfyAjB8W6lO
PJIEadhKdyYAYfijEeQYdZK7XngRhBclzupfTOMkhIbGlOKxd5vMoECt/5Wskiu3
ltqWrw0kTcYj+0W7gYEaLpnNbNdVLhtCNb5caCCNfQC4/Duw/XqvtbD5ijTSJyRb
SRzzXeb2NfCwvSOSdegAECyoX4dvCodhAL5rSoXZjfLjDucv7c6DftojJocHYOK+
ahImAzRR5KJzVeWgA+ySO3iptsd30KNUMr8E77w0NoTtMM3ZSIKMtjmcuOBrlVuq
UIBCk14Svm5CH/uMK5N4xgalaFPPOR61o2Q/C3PrDmO3OfG1ijMsuO97zJLwJ+Np
DfhauNoHw9SfxmxmUYHJZdCtVuT2lEwJm5d7uQT6PwXoxfo93MQyYjJkZVhzXfSh
0sc8Gp4R0epPUU7pzDiTr6H5Y1rlAwEk8f5eyGnASpatOv8RT3BMli3EZzUrwNN0
vNvLRop1ULU3zfHux/tcuH2mky7koPBmeFRR16SAzVang2c1G/8hkhQy0KW86YGR
1IfgViRcF1zmqi098vnxOjtmNHLoXf3H57tnppKKLddYSCUkRSjIYqsilI4N6ONP
prH1JBpuA5wwf27zr5a/2IikHtBx8ZQ3KoMlvd0VGQfn5zpZcycTF0wdKL6BmdZh
gKiLJCuALMXPR2ek3IE0j7LwEYKLk1EzV8ZEey8LIebYNQDjHFXZjBJhyuoPJcyp
FPbt3sifVgjH7vrw9es3Ciqhs9/5sNgjbHvzh02yIhwA4B30nTBgPjrBiknScNZu
T9VxpYVVLqoB1QSReeiE2md7eilGS6ZEBVgBHC9/Fy9wcjvzAgdCrWItb79RhlQ7
KIqLgG5s0P/uWEBtEvHQrPZYbCAGDOuXQaXfPL/TbR+d+qE/YmmwivdyO7KNJ8oz
zOLzGCxtsz8LCud9V9w/a18pa50nbQV89DXC2mVfi+7s+/WAEMalRwq0QNp+Ytii
cXLUq4KlheSbbXKfqH7di898fgv8X5VRka9n/3dqXzhqCVH04CRbbpfFLmFgtxTS
g16k+qffQXj+SXS+MIbjV+haQ4wcrwnvTuDKgzI40h2maai4VyVvIAnGoHB75Tsr
4/XudFZ7CzfZJWhx+3jHmvStTHIIX0OaeC13WN1IvyH9bsGlyI1t2Zx/KdbO431H
NjABlkjK/8j2ms+PmNhM5OmvzT9YXLDX/Q9Nd7c3W42GRYrW+7CxeJ5Zlxmmbx8J
qy3ZXx5XuPkcea2vK9YDoc/VqW/3K0ODX4l5nZpj7UbROtmgwkBgtw/Q1jmbj4iv
gZUXMD1VKpYsrGCDkDBrZgwvah9t2Q8PwQx+ml+3H3f3nunND0WrHij8XRnPP/zD
pUUzYNZ73NUtEMY9eEaA7XT+qepYYHKBc/lB9xXauC/s1TYHeR2Jb9w3GkLEMrWE
NMbTga1KDt8q9SEejf4k+buwgjJZQdBsTNbMqGOrDP4APvbzYHWAEwikaOFF75dx
Tbg7w8LOPtJUpUtq5FtrM4CiSwJ+MCTQU0tO+WJK9Q2MpKCzgf9tf/00Q/cRDZWy
LNa/uxxgyvyt6lQoCnx2ifNMqcsZKuRjdZTsykST+bfD1hwje+BQfbruMDggrpWC
Vb7guwYXBqsUQdg+AW1oaR4rV3GFoQXrxBnOrCD3jSWJNt3TR1xJzDZNvYBURiSa
u2D4qpnf2sAiZxKVqTnEYVPDNilwZheBYvTPXgkNJkbcmiAiohVJk1KpYbYzRsFi
8iQtxBD2h8a8Zak5Z0V0g2yX6o859d4Tfcsz+j7DM/j4QUmcBtqWx5F8t0wot8oy
1qblD7vrIcS/NxWKPHzHDpuOxS42WD8GgWiX1K2Hi3XPDAdoJeMgNghuV+tUYAvN
6cTsxFSD4yiCdyZSVQGg5aM759AHI3BPt1ohgxMSflp/uMh/kAm8uirDyjZIN1mO
g+I+capntYhWm+ESzVN2eDsLHKOomnWa+neHqweJVNrQzV1C1dLgCuP+a6m7ZClC
cqCCB3m9jgSHSj9PZOYgO45ZBh/n0O0BZEFIAXZkma1q8yMyHuZNX3NJM0Ol3EP1
EAkIelYRN0TGKNYAUwHpDrqAvbpFw2wJelZyVPy6F5VBTVex1yPU9kbV5zArbaax
zbuq/sNd510IBvx+rgXMxjginYBGeVET3TbEVwSB+6lkzw1riB6xYrijBnMbEZ0V
8FDMejT3HC7uRLR0awsK6f52b7NWFHZUA6PgBE7fNi/s5a4d/nqXxlPzTaOk72yX
siguoe6a/WNHuJ9M5r3HAAGk7zc9ZXYnCE6iwDJCcxqv7gN+FbaivYr2JYn4Yw4M
XV+Tga7LZ2q6RdgIVrhsGACacGZ4uaaY/rkMQRhME+NffN2WrFlhyidAFwBDOdtB
7seQn9AAzqy1HvDmJ2SCcDNq3mXMVHNKJ68Ir3gefkHsTphT9l3Nde2lTLNrECge
QmtI3VNZdoFeGoIfqyWNBDzAEdO3xv41AVMFcRa8vhUIW6iKx4RywaGSEqJgzZxA
nto4pn9g8n7ZmQGItRIQB0nQGb/N3n+v69Jt7tK9SXnJHhn0YeAQTylX5hSUDyBI
0oNXYtm0ZfypV+ghYdLO4gPWPl3Qatwfrxj/829Emn33UU5lRivKHrAxC6JN74it
KDoCQgVtoEbJT7LWt4Jn2oyxNZV7RmAt5OrDuVBGGQC3l7U5avZDbQegH3v1DwN0
hdvKY26XUIB0sLYi64CVPIufJRhaS+sKa2gRjW4oKs3vBhgb2XJLWsHbBDzBZYAX
XyJMrTWPHJJ/jZxYRjHqbwTw16fX/gq9bYYpjdsf2oAgn+9bBG1zEmB3r+yGBmR0
1QVRnAsMIF+ugUZGl8yAPhVbThjpMnBn4LuMIxrDF+GIXRMgdGVMTD6SzRlb7MF1
rz3xRLrWStC/YUcADDfxcXIVVs8cFWNeoXy1MrgiuQI+QUE0a4WtmZt+ccda2EJ/
lHPGeJIkoWi0Q6COvDkgvULAuHZ47rbBWDEF6clsjHFmu8CDB+nZjNSh1BzYNqIx
fMoiZiTnuiSY/vzmv9WNbjtmarCivCZ+pG+P7gypYH8T0pXvoxy+AXE84k283fZO
sWpHoNCRxFz4yU2c5JH6NgkEeglpRtnkjQLVqtSWQja55FKblJWAlEBZV6JFQXBe
C8Lj5kL1UR3cbnWTH6jIKplMOQIqkCPkSZBysFxv9hFK/z8AviU/NOgf2L20Ev2Q
xawNpNuYKC7vqHrNSaJz7gleJuTyeeR/hssIsJ/CbawTggznQyqnkHPvFGCL8rwj
7KmeresKGblyVl1DAhOcfl490wTICwG4CZi6IceBqNvRvXkogoHCC3kc774fJ/d/
X06LI4MZMxVLunVOXQX1EWyysj6UWpiM1ghBMUIJzuYKRoi0Of+KbJrfkrwD0mrI
bmSskCr3W+FJ84VNK/RDeqkS7rbczKViRkKPynG3uD5XMQdbCjhhDommAblMIJCU
QEvoof6o8PM96YQxP/J2G5HFiAcEPnwDhi6UsvK9q5lD+B1lZX69VCKch04nWaEy
PrJjk2Szqz41cAY8hcVnjMvyz/jGxUF20qBZcseDj1tmDhw4ZHEPXnNaQW406p05
vuqY6GdjwB/uKKW+NBUW3gK06g7L80rwgGYuj8oEBKcDmvSC1OwsoxFbH/iJLS9K
FY54+rCeCcJWVujG7IoQhK3D4Abip5RsDT7CNv+Ob0GVW/hxwOwG2Vc3BxuCQdDq
wZMbjq/bzEyXqgih8vZ03qiDpm0oSAdn5tnyRhDCnDPJidpv99wcIK8gVYWpdA42
wZosKIONrndOYeQWRxv2pI8oow0zVpF/JlEqvNBY7+V479LawwxGA9WnUOzkOWTD
DnX0CI8NOMG5E4Z6jAmvXD2oWfO6Pp0hAxzQtCjUCiu+853jlt/R4QORSxPu3lMr
resc1D4uJG55vVyzl86Wbn/NuBolTLPvXmZFM/dn2S/FHR50VzLfUG6PEPx6YLd4
ZpnqRl1pKYTB9tWYDFxH52M9fDc5VEs5rwn00HXr4HIs+eqdwYJq7vslg6r3E8dS
xywFzAtdSnrfGJqRYfp80Wr38PmBaGitrFEhjMzlx0r6jrm38M+gZpWB/hhwk/IM
3R9Kz9t9Rwz5n06sEAEA9fu+P1wqHs9HcViHAYWusAb5Ne5+ytolvQD8ne93WnMl
IaBVjzKn02DIePbtBTdOZWwiwxAQnQ+1ZtuCY5Qqe1gUS4Ef0BtINHGpLD9WDzaK
Js3MIJ/EmBqRXs18vgad7C+Mm2ZM95F06aLPMsrXfNu4VRC1hYysQwOnZS3qVIjR
bpNMCmH+2dlHV1yI3PMBaPgh28JgkeCGgfQKzGwPBx6uk6W0ly8xJXxuBwXomvJT
/th/O/5LhYsNq50KHxAIit0ZFzMwUDShlpeZfp3xq/1w5bWsZusku3oD+qPn/mSp
nGt98ut78hi94m5QUrbsFWxydI0luOcr2CzGpJXQQT0mHM6dQDRNjy90UBvNfwqg
XcFQXiBcmj4q1NWiCySTx94IoCcsT1OprY6OQ78AGzkqzQX8NNfFRziclhyrxTvd
yOasFoCRJGAXBBevvaC5d9cdsG6H76/tpVrYcHlamnG4B/5D/MzYm3NBmZV+o6rm
ckG1zAe9GUIbiyTK6jWR76UfyHFKizcwPuK30m+dL7ZQ1jfb+SPZ32m57xlm8ArC
lPAqSx9wHwCmkN0VYZQm7FA+iY+uyew/dNFdv8gl7IIENh9TCdnlD8YNeviSVFcp
GJKk+RvwHy+NNFVMmYlV4MP7mdDP0HUEcfPddajbQE/VSxjVQY+thL9C5+nXedCe
nclJjFIDddK8xHvgqIOT8bro2q63sDMsGEEHgktjyNZ/uKvoIJgYnJbt6qNm2IVR
x60Cuv5HI8Rvw5Pk/Fl7GhjHPQ1m/4AFwtBH24JMiEjzO1V6uTXJ38oHEjTzS1rY
+E1EuQrm0C+ocqUhj6CLUiTS3GHM830PrCh7PUvCP5HAnDSY+EM1FZsqshU8yPtr
YvYGMb2+3jn4xhTd+H4nAVG3OoLijJIPvMMrAIyftJau4myVUe1yZrGmO7aOy5fe
m5kDAMQ7Jk8REfplLBtlXknBkxAF+yfC+CjR1ZRL07pFsfkDb/LVsyrrMT7vWyY3
/KZjkQlLqxlvmHOEkW5QbVQZHm+RAKoEKMuaPGC8ijx2GQU4qP81CcI7fZh+zsPc
ENThrLpkkg5MzRlnapSIEiR+RFfthFBIgeZQtCoxeX5GHDw2G5JCy+N7HAl/10B2
8omvIiYAOH7h2/EPgzrW+00OakUMZysw7RUJWmCMLMHW5tSFt24vaxaUbN9XHKmg
q7spgAxA7t3t2mg/uwSTbIKCtH3HpAO+SuISOjsolcpH2LAqtdmxXzC2GAbRWDYa
/u05gOIM6w2B5f7v/OAcJK3zlIWd30xAUWENQBHWDUF4aZkN26minnuEr2vTbnqm
rpMOiPGiz+NUPu8pVMey4GJphMjHoWbSyHVkLYLuxxB81o2VnBMHd8H4HOSq2e91
bWvbVbZCyU/GfehAKyDHlJDI12FAAB5aqkcYr1eTM43xCoJQcWEZKbLQYlnkUYXq
U+BnjN6O2HpffhzfpkXsjHBMVhG9Kp2OLFRoRlm4jp2s+HmFtvRlgOoYVT0LyO4o
qCf5jEDzSUwPR1f/HQHBm9FyxmX7Dsb5OCwZN1+NQh2wQqIUOiC5wEd5tMWXrqFI
ZDOqaiBj15sGasPl7VzLGBwlbCpLPGvPVCwwbwJM1oRQ7An1HEkGXvbh3eZ6BYZO
Oeprnoig+0pId6XRrynUvOQRKwHEE/WlwJfYtl9VnHAZNrFHFfHWwjWK6YMPzoSo
qinvhf9qoPUo0XEX/YqjT/0PYu7p8icOPMNh/sRbJKa+ECCrUmbsUMJslDybZ49d
LLawDSLiGifAUzUdG97aBY+1maswQOez8FYt+wQj428EkC9lFjHpIng2u08z6tYf
LzyafCKaq1IjaSO7eYHdrbguGCmCrZM7I5/yexFuduI7QL6027iiw7A2ikVMcIkJ
soHiY8oaOZUPsYLhqTQHjrlNkBegk+YR+LxDAyVr/K4tk5MMFI3K+FYU0hFAinDE
uC+jxxEbe9sOhgoBjd9vHTQyWa7XaIEvgkonKTISJRN7zZoRIPzZs/d0CCvds+yJ
020+hya4bHY1WGB8TSiL9dFII3sYEQWBMCOx+ei1LRSHO47ynEPTWmEWBIeRVcFC
+Ej5qBLgCOnRjITFBOYm2e+wQj8HLKQGH0u0HJfB+GaYcQlspU92wTCqMKYoVa9E
2nhuaNurXhjjvr5qfsH16NdBf9BDj3Jva3oCDXX4yLgjmJx08WYIN2/5wcJV756c
giVSLoIs2OrrdgdMwzqFil9l6TCRpflFQbUTpvC8USdMGPnSJofmlcM4KG1lqBsb
MwCjxZQxIeEW/a/WdU8R1qmrVkYcs0gtCLbUO06XF92e1kI0q4EZ9A9BebzguZXm
0dPA4TJp+1P8bqBIgQORU3VP50PszqPL56q4xJvd7RX1D5JkgATAQo+pdrjx1d32
qi7u+kbHt04d2vtE2e9DOaEM4Ix16pToOPnfkXTfhBQZbsfunQo3TOVYvyR8tT54
SFHNsxOMxpu2O02wpWlHj+XtebUWFDlMpiBtUT9FMQM4wN/6Dcgc47KK0+JwIn1D
kItOnuAOH1EUL6f78hw7BiTrKmpTdh2upPFu9VFDn7u6PeL/jEo6UAN64FROUJRl
j0by6Xb2Z4ssxus8A1P434eiXNVoiIaVVKwYdiLICAaZNSoUweuYSn5AqDhkaB4W
JJX0rDPPmPwgrHnI8AJVFFvFwASc5OT/ZhTS6ndINIZNB5ICRq/LnvK8YnjzAMQI
25139WJkup+qyDr3xukJ+aF/9qtLUYtGLL53upPUjApA/Ud9u31/LWtsF7V5gRmx
ZD5AuuGWaGzohzOITGL0VDtJmWI0ikpRmPsusrvppmJy7pYMgvgTFA4KWSJoKfPl
ZEAx2XrPMpt/i9klYzJV+wZpziwb0bFt8KI0pe/YkzEJaNOV2EmjGMIMnvcI65zB
GY5drEjVhRfu1v0zx6HrOi+Ml9eemdPIOEyEG7vTHhRzag3arUOThthSHs2EdtWw
Rki4VKJdbf8nY9ofLQvKHdR4piTQUXAHqOUlcrNLY0xT5D0eyiVN+amDjCtKz5Wy
nfiqqV/r5Bm9mHoG47OZddShT5uMON1uwWix492n+6HedADZlsHcvR5Rl41fAXG6
i7vxM3cnjtVxsDe5wL1s0ZG1/BQe49f6e6qf15SK0ULjR6tgz2/BWYkPeRFVxb76
UYUWfS/vvTxbZWGDidbsZXPNBZH1l4O7oVqasacQo4//2QKU2oF74oufkj0MzJc7
t3ftE2ITVNg3ZUuXhWz42KGu2BTC/X3MQ4Ip3IhAMIwmz6nlBtxKEM8inWXVjimV
QO4CEsQDFopzD8mgEZMV6K/OQ5Wb0dqbZjn4y9JHsFURIT+GctjX/KHAEwMJHY7z
3oGCoBv68HJhuANWGpJY2DydD2gEHyes4MBjsnG72ENi1SGh6YdumibEDb+cftTj
U3w1Byqxk3cxFVrE0SDIwR9M1XqoVVOyBLPPxiVeOmIskHB55gCXqtZd2YXl6VrV
kuGf7i9Au+IkCAIfRcBocq4yuwtVEBviTXp8tH/fkHhFEgyM+gdlveeEdJJrECx0
YlqgkIW+P2dy0bF0fC1aemdw7cJg4RrzS1fFWRQReg0/n1ES4DYMrVGSiqZN7z8j
q8DobCMLujsiZSdEw72xUBqD442TaWMqiiwnXMfeQMvmNuPaXngE1P8EXoInRrV7
99Jc9DDc6ORfguXi8qtiI267us+e/gvhahqYfCd4TKjhaZs01MdwJmfwRRTRAGKT
T+83u7t7rHlKbAL7lXf0rQPyYQV8+J90S9XAu756BhR3JZmKRC9e+gV+5FKIMKeR
UE5mLvGX9cUlWaICMuCLU+Gwl57l2RFYYsxGzWtQPScn0sJFK4P+TIxteT5khZqa
7gb7cfJ369WoCfkYyv9pMXR/3JAyzgnRjhT65+Bb25dpSDeXdqOnlhYmjaeqMI01
H9Y1/QIPcCdUzv3NHaOcHvuu3Kecf0Ou81blxnixXgr7XOz9y8w+7+1plk1j2L8y
tLqKfIuIWQhHrkk+0VKdgfkqwf5Kk9vS4B39sfljSZxqH38TkYTK18voJTeCZtjF
BlPXrMdgdf1M4ws2WVJMLru5t3iKWkT4PrNyZOk/d+2WeNN0UEQjq74txMviinN1
n29jfTn/s+vjfHKwjDCHM9INZDZJW5rALfyG0GIrxE5j4Xtw/qO1I9T/BtzZPqEY
WARrZ3leJEZIVYks7aThF2eLZ6zmgsYGuFtir5CsuBgs1IuN+oSITuXE5pCnyhyW
5GAK4XbJ0nys7D8St31155bci/z7hbaunGCCbpEAldvkIoOt1h9OpTQOrrw1PneZ
959Aaph+rnETuljRMU6ftEcOUdD2SpB4S3EmXrlyC5i73D7Btl1wg4viVUmeB85q
Y/6Rj/UXrOT4Vt8UUfruP25wa+cs9q7j+8Co89EyuhHKBThTwxNz0QA89Rltg1uj
udG6jku3Zmt9MMwYHegZoQhoFv3cPJD7aIRv5qyrBkakvSWZmXOG2dpFlgq+aNK8
nOCIVHemKl8G35sy4B5ezEUHq2HJnR/J7wvQ8fMmzID6Y3tDZtsgAmE2+PRR8A5T
5I6mPL0EM3+yPNez6FHlBZtLi4MTOMZmxR0y7r6sP5A8NoOrquP9HTwUfO8i6czI
cwKM493PWivzAtEgNDkRtDNhzvkp+tJGLf8zsEKxVGKRoaZwbC2uY5mhhE642KtR
vf9ycwFEXPczWHU0ZXev2Ew5mLcCIlPoOu7IXUNIFYBWhT4KaWGjCFzGtrvTlJiT
KZjprs6/FFZ5iboqZeiKkUfZksfQxVtwR2iergZ2hraBwB5v9qQkCkQSCPppx3VQ
2eVGtVrErCwapkEXtW0xBiSITNV3B85BJHA2g5q2AzPO6Jz6QdEtsxFPEnNjSnag
bIKToMBDzneA7GtfOKXJWOzKMKV9IWbT+M2toTiv/SCW9v5CZHA6WdTAxM07vKlp
MDs4oIPHBn5d0u+kcf9tVhmLzzhRTyXmywdXaA6OFpq1mM0/EJiK+4THkk23x1b3
098OqkuhOMedu1ko0pu801aoLS425hOrUfaM3p3G4/V9S41EZkrES2wU6rw0xavZ
TEDAXapyP+Zqbd99fTRo4Xa/yv+gAzChla+ns/7aXlPKw0ogOtpcXBjc93zJT9hz
u4y5t+26uyFHo0lrS8oM7xkwx7+ci58V3Uq21+hi42SFLHBwA33sC+q+NjkqdC8g
x5zyRjASorJmqLCMciayGU5d8TPCHwlpK4iD4Pn4zShWDngpW4LoG67XWDtDpm/g
zfipC5HlP564OEq7Bw0x3dfmiIIWESauS8Wskep/DEAchDCiAA/IGpcH3s3Xzhwh
xFgvPc09msiI/Qrjl1vPb2/RdMnaTVPhT5rB6+E4aIBT4ncyF5bjY9FZkU6gbnLN
9MVwXbFs6lh1aOo3QsEAp0qy+1Ib09gyK6BsCZOTsFNO+b38B11lxcnjmIYY4O1z
Y4grlQHaPJ/k9esZ7KNvXVgQjtcTw7Ka0E63zLqg3Z2uupK4ZjFUFWQwiWzyGJZs
i1L9Xy9d0DEFSq+mOImrj82L698iBgMCG9WYR7HMCQT4wS1Sb8xnqxEiuf6FozhG
RvXVdPiYq0N40nMxZ/jv+nmutUE729TyT3NVtRkjW3+xBUObzIh4RcRQEdIxLxbz
Zh/kAPO+EkkpRUyfbEuURe6FtimhdUagHSM4xhn6Iex1Oe2YB1Drm8P/bz1oiDno
AglBWWT/AWONo8w14Ah3qQLdzXWgp1boMYBHormiLe+aKGOSdjyI62y/Q1zZH6g6
J7X6aUOASZvaAlvD6R+Cn0PzLxkpgEIJ/xO40bsPFSql6g4cCHN8OBLo4828Rjrj
v5YnyyWYqU0BY9Uv29Cz30xbDg5O9L6EaOrYwcVZv7aa9cYHqBikTd2VSWsYpWiM
fRW2AhCbhyTh71D4fLD7f0iRMyjin4bicoH0LLPxvT8GGGy1dQJQZ8VCO5z+FEnM
BktkjY2ImilEbw/jdHq0aVCfZSG9czns9xSm2O6qUc7uI5w6mr/j+rPtFXsmiFhT
34g3H6OM7lIC1MX9U0/rYneuo4EgdSsiojXfcPvZ5PDG37efAed3+q6Tao6Eccsi
pTkFBUTu5TAx4bHk9pl40TqzdBAT01koFm2sfg1S+ZuAurXsb4o9mTAu8wBwAjau
gV8EJCW7CtV9hTdUh2MS3lOdNOTZwjXmiBIkp47vGtKTZvjE4/1JLXK3PCTOtV7T
njtSAvQQJnLuzD74ZCpAoDNlUgMdKlIOBHAL9oLNq8rF3rJ0UB/4GPcT9HdF7oe3
wivM7/G6PzMim1F1t6mtCVJNghhCEMUJa64Qw7hClqSAvMV6GUNd/WALTuwBdOpn
TvD5MDKuh1moz0obw/b/8gQRKrGyyWI8L5rFwcvg6W6oRzwZLYySJbAGfRF1uQNz
efxjlfgH5xrEefaq3jvdkpvbdiUDV3x1f2Jn4A/lVUS2XmwpZZZuyGjHqr1YvDnl
uaVvIS73NGCnTt6yGLiwfXu6/UfM2YvpXdBUIjUpsDS+nXZIF6ylIPXt1jD8Rvwe
mNIC2DJLa9JD1VOilrD1YxDvdlrwzUIGNSMf3IEfxNdURCtwUv1Dph3obGk8PN5J
ycr5MI6e2Q1Xo7AKNuPkS1sHa9OLpGBf/jYZAFm7bwZwQNmx4ptNSFiVnm7pqrie
VW5xpsYcUOpfeFTGr5HQcm0OILGEtLvnIIe8V8j6IEOiIo/GAyPFTTLw/G4NOBsm
jgNmRa+QYjhOGRdmH4rfMN3bDWH43DeQa94VfsElKR9nySiRjH3U/UolIQpKeDVC
8C9YO+YdKbeKDSS4vY620Wk42hIZb2rwOxumLYVQNA8QmMfRK0zbkAWmCxsj6x+7
J/RrYco5yTmRR05gIuBAbG20KrWLV57cF+Yn2qcll812XJTDKQGxeikWdb/lZ7dI
qQi/auklg2M8/fYSctn1ATAwU+gJ30/TS7xdgfNMrb+ayhIIdSTmLURHeG1BntyN
EEAca7KaNOZI54EcaDF6+nJ6ieOAekn+uD9etbN+tqbuD4UX9ulaGDv+j6SZ92Ep
9gzGekR3bljhEkOm54Mdow3AtAOvwGH5EGCJkCLVch7G/WiO7jp41Sf69Khk/az2
m5eT0iMkMY1dTS0FZzyS4TKtZ7/ScNHNmla9vsuH7EOgqFqsVYD37hv0h4LXR6Vi
s14ATfQQYb8hGRKkU2VV/LAvyn7nihjkLooKSemhRs4akkXmH9O4z8wf4iNoP6EK
/Vhah8MKc3ZekVwK2RikDos/bofpF6Lpw9fcxpE9E/TKVljUDNd0ig1PyOYr3AIu
55i6DbO5E1tIqUuVMHs2w32K4hul99GIy16FexGP3EDa/k8aB7MbNLf6v1nzE74O
dVs/4CgonZ12ROaf6YgZDXvHVsmW4jGxothwg7YU0FcTwlYll/2FrWGmWYLUMG/G
EaToSSOBG8lLZeEawqJvYR+rLEqTxdcLsV/KRlpgNlwCVUgJkNPAz9o8T2bmGcdY
8jSndrI0nYFw5CJJTS9pS0s4ncsrlXY6VtQM7N1D7DUOFm8B89ht4Tb9VmaTxpcF
oi/um0cpQud9EPWV8DB1MdeEQ5Wx7xWbs1uoAAQK9yDRkGrJxwCmdCMQqhDiLZUW
fDzqfYx4c3O6idQOWOKJxPqXm13RXeHXy8pAT5iOKygtrwXnv8ojrijkpck2sube
1inyVpOj8P8dkrJbHc5Wlpqk7K0SkQjyhsCooVSlbZlw6t0gQkzaGoOalH3+KLrZ
aryc1YssRTa7tJW7xW065XbZOCuMbT2694AqBtN9+BZaClvgaWjQCiBWe1rW591W
utRaBn8LuVoQDHAFZlRzFEg77UCUJcSq7+vXA9w5h8h16onNjNC5QVqfuDeSE8ET
pWbZeS3Hq8ZL+J/ksk8ntypoadOhcpbBIGpgyp2LkIouReqZm2nbbar6mKWZg/PR
cyYqEOCtM9zgI9PyVIbtdODT3D0BGpR647MpTh+uL259xBP8XryBusMqHrRBSAny
rvn+XtpnuZej6i836NIkWSvzyXLCJAoLhxHZWKXK/CqgNcH3Bzo7+5pr43uVLp5H
o7iar+BT4AGtt8jbOy5A8Bw6x8ie9zohMDtYWKC/aXGGm/bKhRjeBPZhahvFDahO
0MebuAZsUkTlMRqjMxmC/i+HbDpLbduxG9Zq0mCbqR0WI8sDlyXy39JQ7/Yb5x12
vIPdRmqnIWg+E2k9C6TPL3b2w9cBsVYjf01iV9xW9MY2maIvBioTcbR0sNeDf0xZ
ljoHVZPINCjPmlsE2GIM7hOpz9gGv48d6AS3e8ZZ++9XL6O7/YThVpaek9eUVpKp
s3S/DkRYP0Tfb8RRhFwYQE+EuKrVHHf71KSX/Han335TKf5Mf493YP5LvKXSBbBo
Tn5bxWYMiVTJTu6OCgksmio0YEDf2bVD3CuH6XLIYescHn2zjX0mOxZrNEhR2IeF
McGJIMMv4FFMp5Z+vWIzgm8gc/W7X7YUTqfadTMIxVBGZTwFN0uGtepZYgLx32jB
In4FJaxiJvvEq/eXzftmR4V3EPDnZyTBd2Fb1R34qkPHI1lMsIqu0oDP7WtUrQnM
y0S1SrgUjOSX3xxAzwIUo6urZPvFWbDnA2SKvl4uQ8JBXT110TDkwtJ1eJR6pu5+
KsG6N1rCXvtiuVRa80jHexWRE50XHRFbpw4h9sSb+vzUbXjzRozmW3N0F3/VOKek
1QW8ElvO7YDiOn3gOamUSJlzo+TYFAri2n7LSwgahbI6Br3crRdwaA3MDyFAMc3c
Mb1cNfdEll12rzK/xdg6wB7V9/94oc6eowT14L908ilXWAHpBbHxBcid9RNG2fho
dKlCj8ILGaNYr7b4LEcHqWCSo64s28JJcAQA2TiT65cYGq9gFhWTwSnSjtpUdDsf
VawP1XXw9cVNf5pi/ztnaVTcw6qxpSVIejqObnLnFc3fdGsKYYjH6cyH++ywVUS8
9X89w00Sfen9693wMkVq3RoqoTXc0ymriIOHWIEZG+NGOTar6hmSPeY2tDNGPU8k
cR4izcaWKO/EUhfNCP19d8eTgzW5C29g6LZgw+hRUCZIt3LsbU+4rJbeNTSsPMN4
l7AmUZZ4YutGqKXPCzZZk1sKKj6Xy++wjwHQ4BsGIbmJOQ5oiP5CGBHW1cSYVS3V
wljgiymSZ/f2+6SV2EWrtV//ZhQ1cRozKJDuNt098LcvlhYE+GDFP7Ju+eRspkNU
ew8iZ26IWIq7DiBGY8QC+OyDTnICiR8Zi2HN1lImkQ50WZAtP7LbBhhQxLfazu3I
XWxokOxmCecKvIfJ5+iaf0nrH2g5Gpqvp6Uvxj/AxyRhl7Gv2bxqnci4GcLZ6NOm
iow7R1v0x/F4b6r+6UKI6UI4Aw3oOZ2zdJ6XWQmky2KFc3my0noRsaOERbftCiwi
Cjm2ZCwqglPgxgYIQDLdBKTVKNZHDw78tbpJpuIwQ+j6wsMVUSbVs/7m5Ztphyl7
9MDnTAwxW/jJCkc65fxry5yyoh226q8k6ePa/C1k62kaZE++b5gcxyhRB3TN49ok
+NKgcpBWWGxjmBEUH2/GRP7S9oMIuxl3ubeHKxpqZzzkIdwaGWgYkEkrI2mri+sK
5VASynIR+JtjWcTdwwVsyCiy6/x9kgSvJ+sNwvSuxNDTIcbNjRy31EZ8OLDYl8lg
+gHD8ceVYwZdKVomczvpWsZNXkKl6d4t+GenEt9WvTq7bIrhRKT+LJSubQaWvMQ4
NxWsjwE3qsp51UnukwMv54R4q2ZEJ+4lIIG14s9UiQ/SLhEvVrpDR8U11VMWyOxo
CuVu6jLgwI/1WGZ1z45gSviYcn6IDJLmowgSyjY2uISBbzRljsSitKTimOv0x0sm
/AgAsChLK3p/eM5b/V6uRS2it7ZmHcezsnwcN+PPvgJp3H2tJoEiwJKvHqzkZOLJ
7/Qr7wadnja3TPsmzI9pnGcu2weLmB9wIuTs1K78GsyrmGrrQWUtWZ0SoLQtuRQr
N4DqlTHEOPGDELWAT2UnWrOI/P+w9N1TvY499qB77D4ju2i84o9xKoL4Qc6J+Omf
nYgC1+dpyazegEWtVSEMXSmZm5YTD92p3+aLt8/X3XMoHxOND7UCnaFiZCzDnf+4
r81bgY9/Rge0MOapocKGKnk+yNXYUONu/eHg3I1Ogi6j6gImQX+sAf5vn5DdysXB
GbclYbRP0x2vncdugL8DDuOtSdN59NbDOd8cJ7g+sgYJJIzmuM78YVHdVCKcHTA9
Jt/+VyUV9GcC0Dr6kJ8VhNp03qJGE0g0c2ZedKE74me6QPv4WYiz6/spC5cWntTc
o3giCILLcfFH6owK337sDHG2VEIUsEAenYl7GcO8QMgYRK0amRHklACBklpLVSFO
1KqvrzR3JUcgr1BsangBiDJbYebyAKzTkjiqjpNvS+g1DQAsQcB+NU/EJMaO9046
/asQBKxLylNkwaIH8CnaYqhBnnNIYAhJJHsJQrJ/CSyEyZbJ/faoh3O5+lk0E+cP
+WvmCMmZX1S36x9lLlwGjRB+e/FOBYdwsAj0iDjyoWgfkttXYA/1fDAFXLM0h4lL
j3rL6BaJCPbcjnrZQKZ0PFKFgOZh757C/d+oJ2GP7SV6rEgWzA9VtYTGuPn3OTHR
ksBULxCPwYbnAM8nWUNkqNwY5oJWuiLNGtGhFCIoxr9kyUTckueoRQwHlcL+WlqG
mBkWH9Ytu7P9TLLHyVTvd/8YSNzCw98yxikwORYH4Bt2iE8I82B7/oQ9kF0THOJt
lEj0nOMXaJEbdVwniLueBg5IMSZ+VOeAjJo2ziEVTViWlKjUjKFJqEKuXKJD+lMJ
WNjSkjYt8AEOEERHsMYZZ7kMqnxBfeG6ZRH/E/JcbBWV75jDBPPSUMeikvC9GH0T
jSz2RBpkmbJFC18PdlKZhic6I26qOUepfTwXO/XKDucIE+VNXOBnYJHOwIwKc/ZN
FWWgUDCrTgZWZszk49PXLRmzOcoCWefUoYNK+/QTD+oCedURO9KpfThpO7NvMwi8
zYJghp4aXBTOZuHX1Nev9Dj8Eq7O2C0MtBzItwB3GVbDO3oh6t0MSww38hoYm2FH
/5yInTGloW67V6qkvglzudlJqjjX37eeq67eKn3ngyAsuUVDrfOvl/WZTi2sP4tp
Qvvu/9pmVwQvwTms9aFoibJdpjxp+imygH8oelB8UfdLVuVzhF7mngeoxOP8VwEA
P89n07acW3J/yke2dgTUvlx7Mu3CfF3pDgFtWBh5zDUVBruUGxMdJ5LnbSlmBuW9
sBZRj8ZlapPv3S3ibKcHKXEUd1yqpOwzzTjZplDPD2rrvYPJjf+lE8bYLY2AJAc5
Vl/nZz/1qDSP7E7hX4ee+LqDmSMDWUy/4EIz9SX9RpmBPmcO9jM3FFVq+mbbg+2q
rGi62W5Tv5CRCbaKkVuLREisxHujy49kueT+d4S7Mewm9w+GYjM2j3fU9pnEpj5a
xKyFc62S4hAl51bQCIoV/5jwVtW0D2WE/khhigx9drKJ7q+AmfqZlZO5xzpBlir2
2txr+lhAd2KE7LbK1qTH3Cz1Nrt5QRVgWDzq+1O45+4AiOdFWu1BI+DAtiZd0sVp
GlnX5+AZAMKGbN8j7NzR+5VJfdL9ZIgDXLSyWgNE24QoVRiNfvJllvk+NuQmiD/C
Kj9Xjd0mJyjXuNTvGxb54QhA50proFuXjaPpE++3Z7FFChg11/eUKxoKLdybx6eh
12jGs35wUKXPOpfmTOncUWnX1v90eiMW/RumRolbEJ4arsVbss0BsqVoJiv5XoJa
EwQtGSrNuCGT0RcVd0FgVpmFultlEfoOx+4FfPOZ5q08SU5MNP+A7DMSgNZyInyQ
V7Q7jFNUHaNIWJN2TqawC41i6yAGl/4bceF/xQ4RQUkoOwLf1UZXlTtTVcaiExRK
6VpJTKOBG1T1jgN0Kn/+4VgCjPfM/Xo7fAq0ig5SJVYxlBdMwbqZd1OpSFmYr2Zp
1ziaAebJhzQvD7nLdVvKd+xXHAay4IeVYOunqzQ0MHxOqc0vl6VdW2mnmNBVhf11
uzP6gWvhEGz82qjAqsDkFY6iPnN3rLxG7CKXBZdRJ/tUHnP7HSgKJrX3MJJ7mPSB
KN5FXTnNKGB5KmupbIDTfV5vKra/w7pUnksuEO39EdRy+FCSYWA+mbazk4+10cNS
zvtUVqTYTM05CRi3Jh+FNnksKQSAuS2jItlP5tXJk+clHiqV9Yz6l19pYipDL46s
qMnuHyYrRMhyCHH4Bwvu6QjTOZDTWOZ62tpvAIlFSZwqR1MwRa5er9KJvrA1Xmm6
kmR6I3+V6e6KLZQA4DTSm254fi/gWwQUaSBVlDDEjH476ufzkwNT4K8aHCv8fAtL
YZC331qTgjrnvgdBsVsj4+LZD7eyhJbKA7+/gCJf8cCqpH2BAql4PsomIMmzsPQt
b5sEMaJKXBnIHYa+8WRNQNrGZCdqVORXo26WOO/n1BONwlmG2DHcGViSwZEGal8W
Obu9DlYGEV0z9cMe1KVGqn7iTMvreaQOYlPksTLL0Y+CcsAlxzOV4t20pfF9olyV
iJRjNw0neEaD5aDcZFzyYTrmk6V67kYxA6yzAqkGeJdbdCGj7TcW5n+3CZ+a001q
XjknL/stvyQHd+VlsKDVWez6GDgDR6ikkUzwWnjTshvXNO++0/QFanWsdcx2LlnX
IWGTUVUHt4Smu/DLm0fOf66aPyrAhn0w6KZKWvpWhLTHaCV285hvTNpY0gwj8hgd
U9CZfXFGblj6Hk57fkvn+//rpTIEKKd84it8rOT9u2nbDjrHyUZ1/TlMqgmC6wiW
yK+2kTsCeIa5lMaKzLLE7kajFyZD/jLJmlfEi/+M5SaDFBn+lV742Yirw04kKO74
IEHn2wUOHNTWB/AepG5LSc8VLjukvQKGbcs0LSi/u3mOQHwWYK0C7tUvYH1zw2kc
QkUak1RRVWWJ8mic7JZa4k3KsM+VS1mhmEcG8xXudKXBg9/z24Uc7Obn6Cnxr3TK
VkD5vZ5GyyC70ZKFrfKWiACt82uSpt6v1eJISlnH87+nHS9xtazSzgv3bz3Sg2//
rhcdOpBNL8ALAxWOFK3jMDzWV8qPDU+YzgVjXvgsnO0BxjDEzeO8YRLagdmSD63O
PjR4Y2h4Pf69B8P/ZXU1NTs4LJmkoDvYNDyqITl6U6k+qNciWpDn0kpTz0PXYVUd
eC2QWwMm0b7TQyXuBWDSQRYaUxFQO4o2vokoLa0o2PRmDQMNtMIK1FJe3F+DukTq
TcXvEFH73eoDJ8Dh4EmTksfnM4uLrU7knPam2YpHJgTyqyTYkuqi/jKLdEIW0BMc
Kvdsl7/IxonXomJ2kYDI5Dxgw1QQerNayuIwkY3EwNKBe/oKXsvam3DzKK64yyAY
l8KzyZ2jQ6qLsdJUMkw0L4q5RbSZkUawnA/2mVZdeO97xU99QRHVXRGM9dAhoYOr
/fVqxPbPtQgFWbONQd8XuXQb/kR/r8G/ndUtcKUXe5CgmMucj59rQGLKyu30S/+F
WfWWCx+/3B2sL8vlt1YQlwTRG5vktUD6CY0p4R78B7Polj9/L71T1S8aoHVxd6hi
/gFw0Cq3Gw+CRfITERvnxsfhVUuNBrFVTMjxa+x4Bq3fEyUqKZ1Japs8WY7dSPka
fox2tMr3qdiTkNchFuv7nJXG6UwRbklW3S6JopNiBUpWq65cmq/uorE74iJJXB0E
g3gt1hwm8ZbA8sJ7tRMIRVXiPTnUWiLydvcT7KDdP/4/5umL1SPRQ2UeWf4JVw1N
m48xKrjz2En9R5CZ3YJq7IA6adG+G4Y7SBRH0OLGcToiJed6uyUhk7FVqo1e1BAP
PSIlgon12Q3GQYCIx4QB3ycyp3VrFvTv52JVsV1rjqOHIuLsZsNZn5MAAeLnhG1S
oWZbTSL54s6RaloTEaFHrSlZUQSM7oVKjP0Wpaekm+0wDdX4TnCOkg9fGv1I6TIk
eQrTfeC0u7UXywI3dcuxXc6aId+tDz6WkSMj4/kdTbXZACXqU9iSwE3Xa/Ii8BrR
ohWOOUKMMj/SLhX2TNCoLdamJSYQ4fYyWWFqyUwlvvxrbSwIrI5iQ8xwGhgamQiF
I3F8ikw8L5cu65a3X9zzmKcgTGj79iBVk6yqVdhFhkpOywaRsYyXkB4BQLPNCsHH
If8cI2wyIMaNkTJy4aoEqjktJNoRcGvo/F6RDWwa0o64o0p6QjVW14FzIwf3YR6A
aFwUrx+UyybOCRaOi/R2uqgBeMbzGVpCzcOVVqzHais5aCpmSqAHOfE3r0Ta4Y8u
4I/BEvG4bP7GeJO6Y44XlbnPWmtvhG7rdjymBxS6Wr/ZK8VfyNS+lB9buTx3O4Zm
OXmfFha9BZ5HN3qfukpLZsH/s7Fzod/XuiGqr4EfyVJSKl2Lcow1xug5gbQ+Cctp
8xNHZYCoNzXbfC7cUcRGEDlfpsAtkuS4021BWKYLwX8/oeCezUwoq0YG8C3AyOF3
tZbWoGa4KEWtVaO5uNaE5WaknhxYbgEmqtsmmPu9twCOaIFTb6Z8TivRQbIS58ch
dn+55Ft7FuC3yyOp1MGXcDlj/8BtN+rgsPAdeQWiAFPOGbAA5Ho46tik8fLV6lu7
0SfUm//6/f9mP9jozBB6NpaYKqbYmoszU/H4x+XQwbD0TbHnKEKsaMIQ8ccmN5tv
AGPHAQ28yb2hjEbG63JWzI2v83bNCNDIRRx/HajoH3sbANDMGbMadr8kXOkTLt+n
i6hMpJNyRofZz5apveXemDlgKfc1sHDk/jhkoF5uyGx6D4dn79QmoFqf2erNo5pK
XgbcuWj0FLpwWXAcUZfYTopxTF8z95Td9b7G3DHsW1bCIfE8xr9imIN1XKkDPAHO
kHJD2C1Zhqee4B1ElrLXl+3JNhjuAhmswojf6W1iN/iSPyrf2cV8bh3opoGfktx+
U4IkbIyk93HiW9Pv/lcIsN4EHA9KKjGEsh7DDnPb3vgMICAnpGuXuBQ0yC20F+D9
sTLmcFPFkEi02SqjT9gFgy9HxpBG/0mfb62GS+MEDs4IOR/4uYu6ywLb9+JeD9NI
KQoiaMMwyFoG4YZtGOM9MfY7r54ef0HiFC8b92fdAzRqbTdxhpKh9/m6QWwu1MP8
gQfz4QlWnl8hTPCFZM2BrAnS06+pFDTIRNl17yfIkuCQ7nlqOWqiamjbFRZrk/7u
v9cwrsj16/6U/sB/WrAEBUUdh91E/vKNq4rTD6OnOcyUEwk3L0t3ZFoIjCvYEOaq
+WlVob07pBazWWcsQ7VHkMIYbJkJUiVAOvzVcgBUR3gnJuXxTwYDZJ/yfjOkMUwP
iVU0xdl23H8y0wI+/ugfG2A9FqMwgGaWYkPb0Xg+hcy8n9mtx/+q6JNRqdLC3RKk
q+JLdlwZECvqRd7IyTh+9gp5s32s+/hGAnBAXJVkpDN00PdTXp6Xu4NcHBFqFmuB
o9GS6Pli0O7jH8FOOWicIbk2+5bO9NdgSmu8aUzuGZWzKwY+RdtDr7W3uGW5cEbD
wLg1k+cYzB7DLsPfOHyK6T4uaBY5m9oKTd62uaPORT1f53vH1Woyp7OmquPiOM7e
f4AbAXVZhTf8oZta6LPxp+2lbVU/BchXyGaDzsLtu0nKsp/RlN1sX0e+FOF0P1Ph
Cj38MjhONmCA/drr+kuOS6Wq9A3Jgf+6tgBFL1BDDlSKvDSpR48ndRqLlNtbcu4G
E5svIdL6PJsoE/gbLCiH2G5GL0N7WFSwS6jiA7wzjvltyBvLfhahYrtlOdFkLBXx
lHMWXJNvfVxke03pvjiO6F54qASUnZPQ5NcWoQJZaYJV2pPvET+q41MD+wYIfizW
0S6Mawn6Bn3MwySDDYRlMgMByHqIRUIioPSuH3KgY1hOX0Lxeed7DrywKRf2iyx3
vunXFNC78qSaH4MT1CFeq96hLQn6B6Ldp5+hjYepMuif+kNAJbq+MUUFKPc63GUs
o0ytEADl7D5kqGOAUcGwMd5QxpMteFVDkrKbrJMSUKLNxLFj3B93jroTXU0go0k+
2hy5tZWNlDTnxPRg2yFT79sxoabzq4FoaCL0fwF6QYIQI9mecFiKvCEp0QMROuQW
LvENHuJblXtmZfnJgDpOHFTG/Y9fNZwq0M1f1I9RkM4aa4qC2L1W1uQYMSZycyqp
CqSPi4xJJfiUNbaH1F4+7obtMguFKFwrTTYQo/d8/i9M6TSYrlyRv7+E9F/8QWCF
yqVqd3fMVQ86jY6c7JvkbtYQ4scnRvaP4YN2kP03ZNY+T77E/16PLbRWE7Cu2XHy
oRl8GqAyQnuuo8xp4rGZAB8g+u19tu8bcGc+kJfOsn3GHohbWRiU9OIlmxfsIOo0
5q8Cgo6YIX8etUtke24t1BToATUOYM7/NZ/xIy/vFFAnEhh9WlLPJXDLuDYjb8+0
tnQ7v1swAWZa0oNx1rZeJn4DmUoHtAP2/dLWtQkjiqdmDxomwn4jYW7xcQkMMGWe
+uP4dOyUCVsmK7rHVlSl5dck/aRlRtxv31VdnR3YHuelEBi+f55EPDPC4zrgRBuX
GVfUKemwt/zMzWqUxGeKu4S9ybqLrqGnqaUmCdDgeGVPB6rZVupaq3xP1fGgUDF4
6xNTnE+ZFfoHTZCdOYVVmdfSjlsFpHP8pLgku3sMscmLJZytgkwycLqgdqjEj028
0ZdedM2Ckh/8DwBeLKXhw/PSSR4cQjJSDC+uA9QWtRIstvAts3/fFv0Fce+218iP
/mO8czSGGAkjLwYtFBbT3ROgiajfVdQ7rOUd2hj+WDgas/Z937M4ZBcwWeflGO2W
M86i/yZAHYQNOmWN5oeSxiosqKCxyhoYWe2QSOuvSag2Ogc48RwMYpB5oVoHfg99
v6PSmNsbfzerOqRCc++sryEcpWPC203UW1Wy/nje3+6uU/sgqOUdO+VmacmuOLSA
vCRXNl5LG921MRHfat0aoEIU3PcnkHZfFVaEhC50+9ILqSeSZAn4p30fTg/Sq6Cc
MhVtehX3e+no/p/rWiY63mX3sfKuI+C5TbaUWcRIzAy1GNvBh8BGoL86JUgTKazW
cWV1j+zVR+T7lgAdD5J0mMv5mZYixOI61/op6mfacdVd7r6TcUAK+1mt0g04fghD
dYpZ7wlqjyd36S5iv916RK82YCh4k/jqoIob+uQlDoeGS3c9rh/mEut+VOgp4+Xa
OMRuPvN5Mo3gfLTVf5FxQ6imsvmri9wjtiQGODVZxvQA1hzLmzbaI5HwGZGtouSg
0wuXrbcCNAfFclRGgq6QrKD4bDdrVow2GIGF3j5U43ZmRBZZAJ/ePZC4Rgb47SO3
T0AWgg84Tot5AA8n/26sOHSzdlFcMkXkZoe09m3LiD531oDaMB5VLe1gWyrqFTgq
AemiMG6afNx3X/qStqGIpHgTkmsjRVsMFIfT6sP71zlVJ+oKJIcLwivU+ykpA5VZ
5qH2/MQerJkpUA+T2jhp+5Pw7YDOjqNQ23N9E55FfHd/kGHoMVOzc0l21ZtThwJB
lsYV5ZGtFPJyCt6/Z2SFw1HFkGzu1Mw7sPcjveKIwIYgsROUcgvCaZdEV23Qe3bA
+1i1Wr3Py5pC6Szf0HbBd0CnH3dZcQITVHhu97vHdakT0hBRF9dp6nL05eGou/i9
hi1l7cVuN1KRH66x0ayQ8jdbAjosi0GocBD0Uur1iF3o9Q9l9R7BuM/GvEo9X34t
vqVTw4FTfctpKClGQNb1nhP4kK4iyKyaRBccIopjNSW8MhhcYaf9x3vZlFVEiTQL
584pB0/NiPaL8SyeyV+1cH9HNXmLSQv5nGAHcKSVBRQnL/GoAXPo4jCXAlpX+L+m
W/oBfJu6BcpvG+vNisvHz0ON6zwYFrAZE6V5op7NSNSCtNF/laWkFPTJrRvalgU8
7wJpvq0kBLtMM6jzF5FQalxOEvC8a3jTUK/xHnpFQXMjrcZKhY8pL0gpHqSxqLBN
6ETOqDbWYXld+/gI9fFGt2cf5SVc1AEFVqICV5fcMdKorW4pLqP8WTZz9goZd6n0
t2Z1ZVkm8VsFZxAPjiQk3wwylwtAey7AXkIDQnhlM4cMAiz+cOv1Ofg+OL4vIyMT
Dq+G2jr+iRgiKKSKa/LVnq5PovVFJeFWxmwTvrM233G7VzMUNY9NzIgJq/UgdKB8
KpLAB+473l1ik/HoJ5aKjPT5BIQeQPtMHrtUgJqf593PZqDw8rbXobT9xUt81uTV
Ry+/4MuCfnJo1tORnJeNhTQHV/54k43vvIriMwV0PYG8C3dJK6PI962ok0P8tFVu
hyyWIK+d1PV+90Ax26lobX+i6hPQ+tsPmhX3yluD6AMztb4LDCvJ0YKxfedxX/FM
uRN/je+RHHN1wv7SbLHD5TMx1ccDrRwkonwWbpJH/0srksM2XNf3gS2afzgF440l
FRgb2kjaFDtVsOaR5xld9ojS0UUmDFLJvcXPiZTqWxXeqAdFCpUKMbovTSQ7JEyp
kxl2UMA1rTPKlxb9Ervs4sXa4TGeyx/E+EdDkPdkwLjkPFVtqKMWdMLhP+4VptJw
Hm8xxcYNMBzGZcH17TMt6uBouA93Zv7ygaVEXrS17d6MugfQ9sxZ9lZgDNQz/CPh
bAT3vnB55g+oiVNJrqStlVud8kPc2k7lhqKAvgJEPVVGPAeBOfT4tHXiixj32Opv
cHb8qdYVmtWdrLp1BfPsM6JABVvVSumjo3fVueHeLAwzMOMTQ34iqS16kqmr+IoW
XHAMFWIvU8vja8w+cPs2uTqUi4iggtNtmT5E/7bhm6H6D1w+i/DM7QR8FwaHArV0
Jfus57w0Yx4j+V6RTiJui0ajM0iFXf9nrNrgLx5ctnh8lwlFdzyP2u6xkEWmkD4S
qMxvb+ai6D3gkxUk+YXXc5GquQJyykkCmt5soyRD2qO+1CyP7rPOiijNpZPJFnT1
asWFhTW4mX8aPpriYZvHIMjAc0b2q7fhQKRL+5zz8MfiNUAhJySGVlGv6QEjOhI4
pu6+Bp8qioolog4VwieQWaIkUIFs50eJR6RS2zYmq3VUw8GQx2vz4nziukLCqSL1
ta4gR5mnalfMuxqYVgUFTW3G4z55l8BVCAs6BjFcmW6xGB5qXZNnts78cJZMBto6
EcpLZu1Ev19+YmGrhfWc7xw3wm2Brhi7Dn+GDuM7ECfBM0G4IWHRy+1gmgxXdXkK
2EEgPO8xugwugB7X4/1+EftL1gDBtKaOpCKDA+fOUsrj79AX6NGTe4IUbL3gmBOn
s2j30mz4FrYiDqkS+OJ5QeEGTPgKloFLxOqX9iu44MKX/vpJYhnNEm0KhgSQRBao
hD3DKPxPEQW6QaU5uDSKqg8xEjL6lxZNlZDqEXQTITAPIBysMy1+tLoUcomczHH1
erlGyrnUvbUyp8v4+cciiq2bInQyoJcjzgXvlDCRqy7mYtqmQ96SQrVubH4C0j/w
dyw4x9rSGX0ejio3DD6F1cbsh0ZwASu6uuK2NDBFF5ZzYZKNun8wOmgn3oXx/Q/H
6rfNwI5e1U176p+mmEkywjaMNdhpcaYvTc0lqlnJ+SWXdfcEMN37BMUyysOyE+w2
gwyACTpvvfTL96kHkuNCR4hM8XCzxyhCuJ+3lwTh03wp5V1tS2NWHcn15GnaxjXV
DQ29H++VuTL44C8ZIZDpgMZhvXExSlDde6VHVCLY1D+LzRn5q13QPzCaF9xw6fLQ
aG5kB2g1QG3SOV03q1tN23sEmMvD2qvU8id9gWRkfRn2EF2rkTcPNrClKEPWujum
RMkH0JvEex/l9j0+HanFP22NjDK4qnjaBeEhay2QpD486i1t3XEFbkoRi4ACihn1
HlpdLOHu94/wEgYHtLsuOnS2NHBqHMd3ySCuXOWogqo3FzlZjnuUD5+wIV0CDgel
2eEEft0ckgpin9gMO72GcBv9g36efjXrbQLE5Ge2JnfkBfP1tO5rpz5EqUKg4YlL
olCqcGqnlOT0UQ+OGDl/jL9wwZqWHlQZij7oDXAVM/qXCR90FjzvCCPV6Q3QSVY9
pA161bpzI9uy+qw+B7g15ozCkIslAfW5NAAGaLOm7hcptDBrdE21Bjgk5eGXINjN
7lrpKs6c6JIOm+RA7MWt5O0lGPkTYawFE+MfRNeyxenjU2dbl9hRDEz/BTBBe66W
DSTrR0LYicEwYmaunDw9jN3vc5xHBi/0u7kGDW2NNSP6afPy1nL1tt0ns2n0mn4Y
sQDc0bVPlO9QhgRxoHlUzK246g/pr58uB9vr0TN1Cr3F/q7rulyf331uSACX3E1w
tTU4GVm/d+u2eGMADAbB3weQf5Oy8N1BI+jm3mbN/42ruj6/yJGAzI/ji7J2ga4M
an8RE//KW0OdlvA8+RGP2HOJefrH0H21FvZqGKx2K9O0h3b2LRCgkfSMq0j4kBfF
Z+F7zI6OlSOmzK4vbMiTixljsfGkxQjFl6PQErhpX3mnmmfN2oEZkFgWrDa8k2pB
x+lj7lRnA+aPLsN9BGXLewi9BQI9ddOGrZPv5GpX+nid7dJG23IFEg5GRBLczWY5
GexN9x0K+iBjoxAQI4gGf0MHObd+jAAfkXQSHZ/WAiJQitkVOKkA9iryFMmPYYhA
sXTgtyDv9DYsoeOv5rn6Puab/3yxkVjVZ0oFalNa68fCGTLuj0rySNf5dtAuJS0w
+P4E0BgCgSBOv9K2Lze9cbI99SkQP5SUBnWqYhHrbCME9zaziTs7FH5HToUzHT7m
6jgLB5TeK/bKARtYEhChaKot+slECpIziyV+cwHFcXFbSrPDNEjORpY0vtm+OVr+
Sb2K3oflL+H87/d+bGj8sT8cmYPyi/9AeCm83ADhWc11dE0Mpv62NTbWhJZwV1qH
bUmHv3SztcVSV2ou7O2vS1pQepJXzZXKzSFHnnt00KFmqfvTpn60r3IluFNuv0mE
6HbdVVhFuRmMJ0qxr7O76VOYRspye5TcIhZNAGz/XvY8D5mPAaceDAhksFULcgJ6
VybC+6Ka3pZ15M+uifwWbosFhpbC+peXzz/4059DgZpFz5l6F6MaLAI20AFIKYP8
eyAUWe9lSXf88dQdcXOXGTWpeE8Yt8m+AGtbpT5aYBXsw4md8j77Mn2PZTQK3KK2
hiGOTzFwYgn3SF82VarurKZiodBqiW7OL6Q8Pe0Dq1pFUvhb7KH5HQhWGpOflr/3
uPEAa4pACAZklSDWWN02HrqB3IXDlAGAX8aXmviC45Uc4cmI/rbHNXeQbG69Fts5
STWAseTfmsVM7TSKPladhseapzyRAnZAaKQM9z4qgcxW08V+udH6T2U6XgQPK3MS
zJUDN7M4nNs1098lFenFfn91mwfVChg9ja+7QaevziZ81dScNcNeh6zoEubJMNFU
LK94RW5sSi+KhXp1PmT2woKeXRfxsai8ga+ggZc9VBwmcr1cILK7PVd+pSnBkYOz
1L8cySt2fJntqVxn61xnUnEHTnOxJrToTHT7HPuHD8vZPwEV2myTWZxSdITEPtEm
3RAgyzJP6gbEVpI5GYalCcYfsYq922fdstharSG2V9oDvQ9NLAGKQS9U++h9rBza
9Bb3PZRx/b7BP4yk4fRH9zbhTj0glUtz1ab2nhsrKk3Jl9vcfwBGpA0PxMYqFM4H
VE7eJZWPCWj/MAwgs35JShF+1xxEbss/hxZsZINgXof8bOHCe1AfSx1nPZZ0TaLU
09VkeMYwLdkD2NK8s5fn8ejDLBXaYsNJN2kkgXAG4Nbe9m1gOqdZn5cC2dRFEDqj
qRGMVNxrNsdCWvRUdkSsTocdD/VBkXIsNvOiEkDflQ3V3sAku/YVOiTiK+f42bPo
zA9H/pxvWXK+q/qCKFMUwHPF265tafiqpXEkvA0GHRkgLAp1wPDsEJsllD9ycFLc
6gutB0DlCGcvdXnYmjEfstA+qn0CVmSuAkqi08kGEfHJ9O3HgaLra4cti54ga3Xz
map/59v71boN60taIcYBHO5w6KYE008YcQHFqzqQcPDaUwsbae9DaSU2C4Rh+t8I
DeQxxEdQNVVMrW1NvuMEB05gi7MlIkFFgVBviQVjJl/OvKDimFCa8Hfb9BP/dkvr
fJ/ksFrrvxTGcjsfvi3jrVvBtJQ8b2lZT11xv9ERVERX4RnS+/OH1k81qXCrPX64
vCyKoFjYdv3HqXi0n9/fPnWBSSnpKVzUEKbVwzKVITT+O9/wiaLcuJ8yUK6L+Moz
SEfmXx54XWCVFx7+SSBZ6GuJ6vXSv5A+Lf8eEvTy4FabjAlM+An5pAy4oiboXC9m
LvVDO5IyNvITtK72DnlI7b8SqH/x0LusXr7oQlkJfikyd/bEPP7IxMm83ZQSkrt9
2q+5S5Fi+Qg+hLUhY68hsaM7StnWhWaLewsphJoOzKN98Mmp41qyiKdEcRYprsN4
DRx0sjDlXi8DIISXU+f+4nWgToPOGpHPzC/zHNT2ZGDCLtbr1TgFoafXHCvNIwx6
Eu3ReG/O0WwfbhGa87DBSRvdxs1luqyxLBIJPC6nrxcw8zkwfsUPLY3vCTPlfL/W
flhbgiWM4xKNHjkTwWF6cCtAOOWU3se4ba3Tt8Q7yyAT8yK2W8kfxaMLlmzanVYL
I52LbUlTY219If1EJbET6HFHfaQv08pDJ8mum0nSfO8LBealuIoQrHQY+KBu8Avn
9FT5vKi3Dc9IoVjulJ62wmHMRoVGUuKE6qrRP3Dlp7WpDmAkAWOm10MnvkoQWaoc
/5cHNRE9m3Ngc7yON/cNzomeCNxq4W5mqVrUCuyIaq76rtgyCGnsU8ImY5S6PQdi
7fCr1tXr6DZRQnFAX0h2WnA42zc/IuHS0t6nVdmjXEB50XuIfQum6H6heCaKYklO
rpbR4IvT1HqXPQK5k6wozpv0hibzyEMHcP2AiQT7RlZJPHh+W6Q6wou0IQhQtyjV
Fkey30tvy0K41Nc2HeRZbKmeTekBGGM1AS/y6OGjr9X5ZWpf9Ha20nd52h7NwX2C
g6oEgQulR/7tQP4lP02lt+pv6SVSEAzz1XqswbRuSIk+9pIDD0jRkgXVllBamQe4
fG+O8UfDHEQB/9uexXS1+I6zsdhtQ3VfYTwJg3XIs+/ciPWMI42Q97eX8AYXxwEF
VDrKkTlDjZMovNSSs0AmbHHI0ttlLc5jjYEpRktIQ2vSSO8EJ2EySONCGFWxSLO6
pSsl8EtcFvRDUsLC3vew0OydeZ3As1D9KGSWZwJYFkiluMRJDx9bvQzSd6hgvds4
hgo3kDsT/3MUNtm0/KvLwSHRYccGaunOWjRJu+nlpwVXRd2AW/uDBxNlJ5oWrW0N
w1Vqu3p6EvCmkvxu5+8y87opoo3hAMnhr70tVaqYNzymXkPJDmbVv5GXw8MjtVVp
7LTFE9P7jBtgqaHSuVlmgLsr28Hty98HjKfHscuegdFXf0UJse7WymLDtQoOLroy
zm4ogBARLve/HxdZIXNmw/V7xoA7KC/2pSCL384vH6rZBfxZ38AAehDqff+cMtpU
zcZanoqSiY/pf5TDeHaLcEbO8jUZP9MROk9oOajJ23KN1gMdWHFCGA1VFJJHctQ9
/SNPoVHD61ouwk8+G6HhE6//nJmYpR7F6iEAfMT/hvjt3RDb5ed9eSJoRKzXxwvf
jEpKJTiCfM7DivKi0+dFQ2/O4Guwr55qRO8zoHmxRW6cGqutE61qiao7naIBMYGg
GQkFSvITTzSVtTvj8DXCPI0Uv5/Go0WeubdV/UAltsyLVQs34PoV/vvOE7bBANkp
j71DMhLLlwR4+Mqv9URUGNVyYFODM5RgDnJDYo01IJkYeDWrhFKTO/Q9PwfHNxU8
5TnmQnOtbw7S3akkv966932IqpPP1/EhQw2zJZ6jtAT278KZZnY83emiTyC36hiB
ZI2/euR/TGO7Z1HB6G9U0suDohhY4vAx1tan2VnPLKRNx1lSI7pfgNc6yk1mOWpA
65LD3qb8gMn31DaxRwJLr+5QG0D86rS7P0f0D0/swdYt3kNjAQB3U6820xUGENIP
LGzheoqdpzQBdvFxv09YN22FDYcZIzGQZmLPTfnECjhF/15TvVu7uBdXeDzNWRdf
3eEwKwR0DO8U74jU2h1F1PE/mcHeUVbZGiDynjIqtQSzl8ivLwGRPZm9InnJCgmE
Cy1q2i54jFYRgxSSXLs8zg0xySxUauYLXfRm3id0YOxP07kO4hs1efrvQY/+yYCW
aAnP9OUgpFSEFlEB8q+53GwugqE/L2J72G21P7ySq8C2HuHRZkGVe01siKpF9eNA
JlQWEcnrNjh2QDsLGVyDS5Yx2AOjfEpFvWVOHkYvBh6LIPIwG6hOkzkMw1YCr2XP
vLm9mH969bCctHDgoZwjjp5eH/nvGj3cpJ4C82pbO+2eSC4Qvg8J/Rb3yNhpGiWG
HLeCjRdaTvKL5SZTbXc9Y7rwOEPxjxTeh7TBh/P878iBbgzqXB1PHb6fatrvdBDL
IQTpJHnNu0JyJ6cxLmUrhn7XuBETvNrZNEPuJuefmB35fdFYn8i3BXkJpPjMgQJE
WQzxEGNq1ZtMtsp+oi3bomeB2abv3MYVCAx1feejGL8SfP5W/Tmbotmp5JD1yYaO
kRZ2Kl3lD2TF0BfCrfIqI+YkVd7mc3/Qy5Z5xbFVYVM5nunle+oLcpLJZ3lJlRrC
dDQ64tovUdI4PDUfsrFTa1q78wEmIIOibLb+UlB9ksU3m67pw5ZkMizsR1jXEKSB
Ouw8MWbG3AQqee9AMMCQ6wgep2wc/V4jX5xVdhjnEF42itMHIe+1nLJNV6U4asF/
y5HHecIggYjvdZDr2b2I+a40NW0J08BI59F5fDFULGVjpIUZjtiNCncR5UThpHWu
xkVr+smb/cP58VPUKqTEdkjgYdwFcdLRdV6Mxn2L+HxQv9jCHEwGq+HPi6nNYXmw
l8vJObe29eVBCsb9Kay5AZGng+4Q+cOxjwCuxD9WzuNLr2ZYXDUXufbmsYzTifjl
MXepY4GRaa0FzPMh1tpIJEzCkTY/cZ6cU3rtZla3ET74NiMhZU4tipi1onrJlost
moh/4aZGxaAb81cPpmY2EvbYXCKwPrdeV7JV1KbKh/tQT3DqvPaLsl7RLcXGRzpM
iywiFMalkYnFT4G9tZdaE3/j5J0tYwJt0pA8u9dm1ECYyNh0LqwUt8OAcJUFSzdm
hTpAgSCNNxLudxAuCZBElJ6ndCvN98GgVvb0ZYe9f2cVTxbr86CtoeZK2JjGU+HN
KekDQwvjRAzp7TD6Vp+9O75gtPnU0eikbZiDla8WT7YIPBP/lc8j9rSyGeEdawOK
myOC9kyOh6L7EKhOKhtUPenjqes/0snuAQ/KgP6O1snncYww+Q0hxYhe8S7y/2dN
77cdoP/kaVJzCg6Npj8AO41N5/2vYIAert9NiiNIgiOK8B5xjsR5w1mkh45Bo9oA
CmEO++wXGKAbhccmoDFOiKwI1yfOi7iIdoPFzfA/+3e/5hJL263Md/apMcnl5As0
Q6SYBEd+iI7mkpuTK6ZScPIlH3dEICH83ou157bl8IlEct7Lk2pz9Hcs9L1cNmWX
5ecM6JqVxERrCbq50ni7nn61bqp7pPQUY00TZ9mIRr8xqSBj7uxiT5hMQojDMfqn
4CU4oBO0Tpx2GDRj/RwfsruZDKm0JM4E0z7juKQuIEvifcXHKhogYjWVGfegNVGl
I0sEdtqhKS0uEmOtHBCpkelWhILcH0w1TA9BaoV7nMy+fG+NS7Z1paj598hHaqTL
StIrLl5DNpUhmaNWmY7cz/8VinwikqTU5jtpV8rmYVU7c9o96LVdcyIucr9SsjHv
Ybizda91/Dztga6SYQjmtG3sen95IqNTAK9B3v68bMt3lzHvZCGUOq5BgZ75Y7WZ
EHHaldntkggzAVY1qLM16+Qx9LgUbY4MuUTNbnP7l5/Z3ayi9DWeQL1c45pfJnDO
cEQsEzXCxgj0BBSW/PuhtJkmJmG6vBa3gqdraihw01hAFgHravB/jukejgNlSq6c
KeVy2B2M+Yr/dBD6LFsLaLfLfdEjGKpQ3aHp4E0TkCqAPyi7ikyqVvvMtSt9O43F
jbxTCygF0i4vBNRkpzI/IzQFftWhigEMKN3suFpSWD2gG7GiJwZ35+S5kzapN4J+
xEUtE+qRHaGBc1wIqMujnbS8nKWB7VOeLgs0Rxe+Pwbwg7ODPzkcceZeut7AVPMY
krYCEJfnDFDFt65N2itbHCDNRIl1nRwlOkODk0tWXRbm5I8yoJUjhfBRVQYtuBGG
p4KBGUYamIn6CjQxPcSPc2HorQl0oP6cAyACT1+NhEbNd4bMoiK4/8wIeSAIuwre
lp8SA/XohPraYy65fBto5SY23zBTX2nw2eBoKvU+R9JnD3xkPuadtQYgC9QS9UEh
7D2H4d1D0LhYh3+83NG+b8fpLwwyLrXGO5Ey3crhBS4O/AYHE23smJf++MK56PbZ
EwUjNfWG7ZoXri/snk5oRIvPLU0sI85+wLD3NrMpeDx3O5scbitdRTcEie25ehuU
0s/wX9lA8R+4tTfzdxFdFZM1b9tJdJol8v5W7KZlJokg7Q8lfZsUO0x1REWLG4ST
0LF7w/96xg/onQyLllDW8ibCsFgt+dU5jHnGrT1tZZEzd+34EgoQXuPVppkpErml
HnSHAgRcMMJoXK1fpwrstcL5hfJLwjZMvJDKnMcBCxMPo+v+hGB/WsYnYUYhwjhU
VOpKijJqRIpYeBqMmlE9wMTYQGhRxYaVg1b1mDmSupYljNkhCyJ1bvOuxnPSf0UE
VHQXBUMAbOX5/d+PHPsjiKCG+lh7bOgc9Cp98TCIdH+j1ZUz2dAGMsWz7kFUthIW
GBLb7LgZ70/gk4GTgksey4fU31nhm/xbjwfzn1zxPnA8RZ9xVOsBnUgFoG8F3aQk
UGcyWtx51hjNtGbg2EhtYRpWhBP2RbHbPhFvtBcMY2ea+wbKYuDKkVPw8Co4tILH
7NVgduIy7NDfaRD5LXigsXIRK9EiwwpPp+pRzfO0MqN5SwNrxSnwSavJmRSKuamb
y2SynibJYw2XqMPkf6CLxqUMFJmsCCFRCbK2HCjoemrrX7h9upYshIJ6df0ynq95
FAJX90L0+HQBDPKwyfyVl/nHYas8SYa5TnDcdsxSEnTD+vdlTtKPNuf1XVa+FK3O
gCzjkKw/iUMWPiXth7HQGjWoQrTNyzjQCDOuiC8nJmihn6UZueWvQ1Wbnf+f++Nf
SUjIezDs8K5T3Mt79Wh4b8RwgOoEZSqetupI+PLOo5WjhvEJyzAKD8mXhQYHcrQ1
TXeIMCsxCQBfs9f2DhLH8X3j2GgTgGRZDBA5tl3yo/n9YIiG++j4NgIencGrPyTT
RFHGQOh7r0uLixzFV8vOajM6/6nbwcrlmQIsZDJkNL8YKs0sTiMUAlljYlKBqjUH
veJ0rqAZRuFew0NQbEXKsSVShbkByQgwU0XBHK9HDni0x/KCZkvlcCBMRUDEdACO
dlPP2NDaKdC9W6LWdZGJ+dokNh0g70JYnC+AD19t8SmlTHLRjBzuVU3tKvfgUGs+
WQ0gRVT4My1QV2ntaxX73NMbMmEXfUaZZprSl591+00nTW98277uuzIF1w3va5JW
vYN/dgpIvQb7kNs/PEfzxflLcFhzCCfG7J5DZCl1Zwe7oRRFYSr3uYEGz5/JpcVc
ANt/jox46HwFOkj/IXkZncnQ3YcNmYSaCf15bmdny2updTnEWgsvBjq76SKSG7LC
X6ZKoYHdb1JXfR5lFkEQ1VbHBND4LM01kaP/X50k/rH8VNDzM+tV1pL2sDITa6qB
bNaUNWtICRJ1W9A/OfG1RaUsgiKvXbl1+vyABaRNFQf78D5/K5UycaP/nOw9YtkW
bFr7FEJm3/cuKkuHcSoywFpPKwKyEqbiAo4U8VOeNQT1JojKZkYQzvdzcuNtyMkS
kixR6k2kjVj3YDGQKD13JZXSyZrNIDeexZ8SfS0IN9Vqn3Hj5cW+8Y/YzYx6x2gZ
o/5Sc01kzzGhWuvD3gb8lNt847kWy0jRISmg64hF1y45Ofpl6imjBiuYjp9+cjEh
yikHeWAN3O4WgRA/08qBnNuOoKJQ+aY9ZtcdXrLaq0hxulhN3DvQT9gBB+MNNuc7
4ixxFhGGUtIr7qe9JNmjP6WUPJO3tcBjB0x+5zK9zGuwL2413XEbmM6ACqvZJFOo
guc/buIMRviwJVJi9PHhjMA6wn1o9JBVHWU9FSn4MkH6LhY9PefBnYRV2im5NbaV
QQ60OX//ATYcLTIwkhu6/jgjlpj9aG7QNhF4u1t5mUyEESXT7GYdPrWRbH2WJRwc
B11f9+3GNvEsUMXYhFjDtEphAu1TuY3YNLPX8qR1FxEBLlXxhNofdhgyk/JyAUdN
ZkXMRntFo7C+ICEruuPsfepZaJgi1T9pY2Y6lPzOp7KoYvl/VcPl0eyoVwF2k9zU
BiiUPDP/E1I6EzG3u0VteVN+DJrbUebazgOA8LGoPA1BKAtRo7MfoPS6JDeR/3HZ
/IE0JxyrwgnWLUEwC3Vao2rttT+ut9swW3SKuAv8ggtbJT2spYXWCHLY2nKxMEJ+
PTbc2QONbmfbwglXYv9Va33+TE08XJ9TvVxWF9E4oiSTXjdCpwX+1iQZolEjWVC9
KB9UoZ2298Nka30LU0tEFmAKDFvseUkCpSOc+1JZ6TQI4HMLUhMmbSe2WCdKhkuq
1lxNJXbE7kxmPeMMDLNzIZ0PI0c+HkI/aC4ynpr47vdedTd8VXVx7uSnbIp8Ah/s
5fd1U9eBD8XSqgUt16aEi91ndg0BdkiJwD04/V6fWteWPt4+sjdjwcJUIw7ioY6C
rsiqPtIN61x4WITqCR7EkwIfGMOzgE1m6JZgCWZ2bS8GEoFdSadYLbMrD5Ahi2Yo
rNe5UGD2akYvh0VPJqjM8yUa2aE4C9QFdNRxXuFk1xKV9FvvISk+zRjcxLgyZaE8
u8cFzGiCBzlgZX3oZSux295mtIntNDy3wRJ8YIntth7FPGOV5YvgVwI2RYUVgUsI
6ipwrmhkebjPi8tfmnHo5oj50OXjqYik3a/vGyHXBuJNX6OaQIUenyd0bZ5DqCr2
hDXkX/GxYflrWck0FWgmphNB8VTuDKaoBpeaDVRSEXYoEqlZHeBrQiTZYP999gCR
7coljnnhfUc/tOXhfz/P7y+N4KRbCVszBygDMWvBAS2krEXRKxhbQrmhjTam8UHc
+ZbJrefXIobmaeFYs0E+mUE7DjFlhuDd8jA1WmmEccKvG5R5k7TvKIFCFRaCKzX4
0DusYKpLtmRN7W/29OyuGppi7A7L+0zCDDDvdh/UceuyXfzNLIFdxmT/tq1cU1E+
39sTFIu/vySv+AHyxxHSQ2kspFhDBICcBu5dlrlib1sD/WIJE9r4ihxCZ5v9qQaI
SOpBr4FK0v0Ihg2+tswgAYa1qlE1Mr93xZblBbrpvfgznHS86kjRk3BqomJJaNFK
9EbsMeL/9W9/Cnz27iEwlW6QD0usgkqPMCbs2fbSkIeBiHc76Ma7iaK0HPGyxoI7
QbVATr39T0UU1AlOBMByINQupQY/zbwX9/WSlSSwFdgPI9o8VWq7jH4M6iGnNY/q
1nn9N3ILCf5XqAEZDzIymi4nlWEDMuX/6LdKHuJlZ3FiAuTido05wIasjWOTlQVU
J4tVGqVn9p2JNbPYFW5TYRWf/+bsIOBu62rci4Rs2ugMq4EqqE6LPGD8FDT3dhHN
6+19RqE/eONVKi4TFdxf4Y3N45q1ZQWc88cV2yUDxihNBsaiZOt2kK3MLy7lQMWL
O/Z7tGoXSLIk3co0dlLqzXbLWRfTpBIfLD0of0bDPO227uTm74QC9BtzYI2syvQ2
tEjlcnG/DsUBA4Ig67OcnGCT5nJZzkfVqIPm4BGrGrLOQFmqweljbHHhTJTG1Uft
E3adCNFtAX4mRBKcje1LTAbmy/igmdcq4gPHSvptSbORDC3a0a2HkCzDI30jLU/B
l0Fz6bHO6Nonpc9qBwV01wB/GDi5IY1rNTwCtL7APf7YIziIK+TpWvwy6DcHhG9H
TdW8/TXmJtI565iGNTGj5Bl6i58rGkTTiRrwRn7sUJjzys+WA/QroEhi6tahgMwb
0hVLFFSYONjaHwxmQ5rpH7O+sSIjnK+LcPxrVObYZDzjJyNLxZ4nnUH1v9j+GRF5
45nMNQwfvJJ+Xhf7pDMoVm+TJI4ie1EtO8jnktmrOqSu8wOjQ/0F2c0NZVisah5m
0dxQcY0Y7dgjgch4I6ZUSaXpBRDq5LHSw7ZhMn0xFFFuxjvueYxt5vM4UMOp/pvy
0pihdZsts9/g1EAG6wbzgwY4VsMmlq9s3GkwtZ0rrOJIglrNBdEx9mtVnJ8Tk3p2
lrSaieWJuS9KqE3ZfFatWVYGflOzvkRANsDOPo9h1fa/P6KfI1fu2fA+3ezAGCin
AIQ7qSMNMRs1+vZDf6f5WHhn5e/lFicNLNvomh8+mP23QcMnJaNPh/7QsvAFnwGD
wZQLIhcCbvHgIZIMAYfNnuan0Tv4526+vtZE75mkCR7/I+wh/fh/9Meu2+kiEL+v
KA2ecQcwqy5xFWdlgWUC4ggwqDhykh5d1zLq5AJ+6zYiJKMzUay9vjctizEc1vC8
B6l9LGB+fic/93GvuvmShPF0Q6AXg7RO1HNM81uQpaXbt/n0B0KuwpM0ycedwr3C
x55l76e4bsWGm5B9a4uzPV41qPi0PZgYdwUdccAeI9We3i7mUEuXra1C3mbRMmve
2Fi46CfjAsSz3Mbi0oQAkhf/mtCdDmCje783LWP/npW9FYy9AGV0iR8VvOXb2Fpo
VYdtbfUpkfHs3Zpt6JPBzT4Cc7tDyT31B2RtA3KLPOsenkKma97Pxaw+lPXkYkQe
93xI20NU7OPKaQJRbh+NhLv6qQuRB5o0rNBxf6U3ciRR7Yu+2r+uoVi+Qs4lJPEc
sPo1CwSVoJtBoK5yeExOQRTYYksb0/gBqgHcjjCTSOpKII+1s+r9ENSod+nX1DBr
krfpJtn/KP0TsZpV0P4OevCNCdig8YTPWgO8j+qI+gyOgHW5KINvp2B69Jga22VZ
OHV2CnHB0fIDakklfRAG4TMaj6RRxHX+0zesXNyNsOAsOmWwQETXvSQLgE0frDIS
vav3fSSeVvkybmXRC88N4MRQbpPkSA0+1NuEpmuOVWo/kJepOoIPsQ5/oNy7jcZe
xOJ8QQS8zi4QAMqbS33nyEQ/dUVWL5ET1h1zkazchlPVgo7kO6OUumYziwT2L94D
hPQwT6wZZR2ouQC1u0XgJTTMRTy/1A8Wnxmylo5KCgWATReL89zIsygXwsapNUe9
lHYCrUdSctFtPPynieCiNgf5USBMm3kWV4YDAzqe8ReMwbG6nnUhzI2Hmhv6HSTb
hRmd2CUERoUq2BbNPQSpld4hYKomIfBQmuhz1JiVXZWSZ7tfrVws38cqjpajD020
3G63J9tCNeW74fehKJWyltMHYVY2RPTw7PxqQJCZN+4Ea28p+Ga3fszIJpjAXzLW
HGN/+7jnX/lxAV4ykncrvuwT5PK1lVUJ5JsrR0dBpZTOWFeBUHHGlSMj3dz0l/cV
10S5YNde/3vkVK2/WPPynTTD+Szyki3WLcDmPgMUI8b4gLG21ZmQbLHzFTU21v9l
uT4KByvww2Zh1D9Ic9OwK3NHeW5p0hBBbvORoClCNzkRdVHAvGJoxFI+zhMDL9xd
xUZ8SqNpE/J+8UVwOkwflGoCEmV3CvPcHhMLFwjgWrYt8tESJD2Qztn1WTmLkg0c
jbZT66CtlMCW50iVo7L8w97MVO+NWf7neRlOMUHQxnLepx9IiXAM8TaMp+jw+Mqz
Xnugi8qOlVgLXVtmUrVv8ZUd8s3En0XoTKKvUAs+aIYI+Wcy1kDiQCO2SFJg8vul
nor2E91ZhB5kmEQBL6GletRwe+J+9Ty0iEMghtRlisie2sbWmmUcchuD7pRssRtX
EKLxgI+/At2tfV47ICAzFPU91GRFChJtv4zfblRiyzT6etmSpldxdI7dlMtVXSpz
vAR7ZWX+80sP4CTIrs7djRPD0nrEUEsZa5XdlCU7Bl90aZ0CB9MXmQQykJLyDjxG
bt6+Bm6Oy/u3PVxSs5ryTt4jLftSEIqgzdX3mQeQw8uI2mcY5kpDz9b8yc9zR6z6
LcblvykBsxl9tiPRvmXiyZ/ayMfciLyEkJ4ECD1S+N8Xe1IWdp2B2octQhCXOW9v
6NM2JKjZX5609bIXpC0kCpZUSbqNJk0xb6/B/lrwMoknXH2r4ecxqfqw6fCVj8HJ
ec5mjrWDlGkrZ493hyv8E5hrvs+nIquMLmNHsfki2FunpHMI4OVdu/R5KyUA5KSQ
izGkt0+Fz4BZauuUW0BBGncWgUcxiCEqCHN+zYolnzCXaszT0gEhyW5JvyKTkOWv
xTuIHjBaMyfdQsT7kHtWp3tSxPe4uNFW0fURZIHxXPSlmxt/H8Dnsh+xrm3kTQDT
CFJxCCJiWKc+Gsx8kYBtfbPyXIGdg4TmEW1BrbA8ZLQILwcW+M2oAGI7dw997SXj
SD1K09uBxsikV4j0/FMO12ovGj7HlkNAZAd/H2jN8MwEjClMbRu00gqtpMBymas4
lL8B2cw19udjQiVVXKMCEQiTt2s+yKwiWq6dFypp9wRX8z2RzgdwC7/x3Ls19UC1
qs8q4t0FmDIapPluWxKlvug+bhkn21chu0cHhu8cjOtiE7xvLg0TwPzwAkrxKJ9a
ThG22NZXJco4b1vkovLPVcsdFAzclYIsy/TwEJNmPdiFOweuWaL+H98Tz2bdJhjC
c21QcJXdSZ8FSdTRKGLNu1z5ttKE/Q7uDTV9SHJ6AdlykjuGAJtCeHsljDCL9nvk
mXA0IuTyYROCDNiz4WatAG767Zhy1lA2uoTtX/SRJGFMgLCp/alSMtzRFSuunceQ
beAfk3vV+KyRGjuIP751R4nkwsQ6IKTAkRCIYPoezIBENbqdHjOdWErR/ozEhgms
RfQ23FXIarJRUzr/ul+R4tggp1AVsrIsnZBS1AleGrvfV5rEdan/D80KlMTP4KO4
gwVTD7rDo6EaTEkie6MnRnwUwu84wNMDbVMlNh6qHqDpfx9OtBnmK0/c8Cjavaxv
V1WHJrHa97cG0TwvjZRsLNlxShY5ICcEc6hfluA5uVBkACcx/RDjK+ShCnt2XvKu
WIPwVJX6+BUnHcksTmItDRXp/OC4GclzmecLC+WiFLOysfS6o3S+MuxtAFhgxTvb
OlTC3Pt/O1fMFj+HscV+nmLZhC1Bht7owR6CkeO0+7oOrgXubSlVhdk1cFnSuRz4
n/1OJ1DpbiZygYClCsrOmujIWZinUGwy/YFLJaIp42FsPVnNN5maUxKq9qGbgkyE
dqV0fPYSaK8BQVmOG23Go5dxjb4myrrSK99d9BcX0/vM7nsbGY1z4UPCMFVFZmHT
REys9ilQv7XCrEjv3RAg63r3Ja/LljXnALSp6bLzpbaiXN7GGFeFcPFA+z7x7QFz
rEUTc3NoCejpwkyplh9q5cyzbPx+IxcdW9TTjUzGqenqJeLl6DqDrPY3CnNvSfvu
F2rCUuo/lWK2ILmeRAfdg194eCoWZSnpoov9pLtGpgjswuKEAUuFGQWEWLik67TI
FvOZCJRPako6WLdCRkBy5VVvALm51kEkdEbqsLXg5KhX5gVVN/06Pd4REkx5nmV6
lwZ/kLhPgm5OPRQgL/QZYM6cmv5mHNZ7lMwfCCLZHRzvhTrKWWGm3DCwnp+Tu5P1
9pR63a9hZ24oO/BsLj/6Xs1xRJv1rwgYqCvgmER6AVSgj1VfbqXcb/+nDHL4ae7d
/3lz+hSJymUJXPgKkqOWn94uGRs9VBee2F2Bwaz0VTX6PBMXYcGoHmd9hK7MPaq6
rx1Su4njl/E8Du1ru+n5K5iuS6qkughdETp8AWjBDEJ2dKzSlSEMrqtrmASnUX2U
cpcL9hyahGko+ZlL6bFscvJsOwNm3KKrfhEzS5Nes2uZhnKADYnIl2aM8ATyH9Ox
LLnf3LY5HYsXssQuKg6IYpGaIlts42JxevNMjR3fD7GPErvAdZ4GLVpuwyzZZn0U
LW7Kxpu5L1pSiwD7AOVWYWYMQYtHRb08cmSHH79sRisgwud9KCinhPmetxhuz6NY
e9M1LyEMAaXaESo3aLN4E2Ss5XeJBOGXPF7yky0mVmyECNko1/6GQgLU8vQ2WKLE
y3Dr2WUg44znoHeP/uvYjRzvoKhoGN6NkYtJmfvVZLFKOc+fLF2WhTQo43yfaMOb
htP8Hi4h5EHCuv+kkkRiMyAEx8sseHbUZpOfv9CyRFtHtidiGp77DMKz8ZF5PwdA
s84l8gO9z0pMtOcOGoTRmS2edla7x7svoLheGCu4up+SSgMiZO1dwaH10jugIKBc
41i0H+P+LDfjV/5Ob+1m9ShLdWaCoZ2kzdar/EyalNInYpTkJmYDnqRg5O6XLUV8
xKwu0ePnqpshBFX/zMCvRB6VwBvlbNwSIFJxhuEmZ+sAYg4QHjOq0WYSymCCqMT/
LLpBARdAexvY2LewcX+vDDMBrqI+Cx4+XI+NUyL89pfov0XHg4r96wJ07CzFwWDA
16AJ+VZoqHBRFZTquFzY8daf/z8IVfOGTWzBNDaxUkbiqKAv7gWQuir1sQmNnseC
SBzKmKp8gwjTdrv4xN+DfM9tikozxBeftxz1N5x/SC3YYfG2zKTkULDRP2fZK38b
tH2LUIJdSTOqKIaIMTzdWW86Z18G1NjOzZMcMMP7S8gpklOCskTnTy8zJ4wDyOae
cLsPMdNPBdzo+o3/fCUsxAAXM8FYNnZCh4+aZrRpj0JyWyEkDxB/F147pue1C96R
xC525tJrZgV8KV/nyYAeXTUr4kMp1FtF7wDisCaL1Kgqg/XLV8eyrTbzUw3VpM2a
8VXkhM24Jk4oGI6gEI4GAbpJtjDXA/Ds5tOpUm2uNTfXy4UeZkhp0evMTWJu3W1C
mD92oHGnm4OH8aRz878X3Ma2EN8EF2uznVkPDNIY/0pZ9gHI/9WVhwKw4QrgUUqY
ucPIK1Nu5F7veqFnFtNaAfc+HrYPsDHBpuRVbwuG1+tlbXKmxjFelpslj4yQXyrB
M61eeoQ9PSBVebIBNh+1CRqbGZb5EfckMs0G8WikwaTMqvd7B3rbxH99YcaAjcDQ
20U1vcgamCr3HMU4HewIUtw50iyFAPXfnBgSfJ8HTJ5PmzA5A03d5bWhC7K2TreP
pvQO8KubnhG8KKRR3gwfy3tgeM1ZaYcXT4u6YQZCZxgvVADCBnfeYmHjhNMwD0PP
NFr+TBmyPEf1wvyV6cpJb6doS1fqdbx/W3nlgIKuW6vHCXrZJ9wqZdCWivYkzWPl
ifaResIDsH9C8sGRO783zZVVvbz8nSamqH970Mybp7S+wkYVu5OlvNdDCAAHw2gJ
y1RLESqMQZdXg3RSqK6RC4YvHTCMpPXBfd6TdM+y0vVsla4Z507oUnwBYdBEbqPV
cvFfCJGB41nhHLaxXg6zgyOtIrMkGeYgrs3TniuypshK30qhDijZLs7nPvxPqGtP
D+JQ2bD+05CpdnzNT1+2gyr+kEjraZnLXCb5J3/gZTD/dcSnrjGbbrHOAYvMZATu
uNJTXaPy6Us2l03pCWp10dW+dXFnuT9ngHJlD8R2jNHJSVRR9fc92SmMHfhBW99m
nQgWCk7P9uuQ5OC3ns2WbYrnuYUeVNQt+nz/u9xoPu01CTHFY26Hbnw9FZVb2W+n
qzfNj/pCvH59s8qS5bpqdHMopZlLjKPcJq1GXZfKXDoqnGd58DEDB2ZdUpvWuy+W
9Wtew0efQRvJL3QDfQZSy/ttGzTEpuTajjEdu66PGQTSRPF5azM19nwQ7nvf4BIR
71UxHs5nnZ5zpND8fP8+mk9dtOAEsy2jeJmWbsDNayJDnawfWInSkNWCnMMwy8z1
6E7C69CyRj1xxC/oq4YJsoyGF3R1pcvSnFb0YD3oKjwCbDJlYgpvEz2FDvUjYGWl
jF3MDCAcZYkNVT2hVH8ZMKu5cGW1lAokkHGTHmACMPZk9/TgscVI/hayIcQIsmWD
kOvBao7JPWvNVcxpY/pXsTBuUikRIXbj0n1U+3qwSjlwcg5+bqSGnucpxAC2Ad0Y
2CeaSIzEsdwo5s5Urbh/eXCjK7wSm72d4nxalAlpC4lTdokAHaJBHZ5mMESmYXiX
h6OfcBTxX3oMaxiMXegpDVo/6xtYNrXfkfR3UeKJ6Qr1Ji6gnD6YCvf1FpOlVfXm
BK8UGCENtlYYaffMPCYeqzrf5f0KSVj5vqY+fnMNFSDhUXJ6h55LvNsqRZPALSVB
dYynwmpmk8IJM0gTnCjoLGf2QddJKtvSzo6JU7oAjJEj0Wnw/vrvOEersimz24yt
Z2FsFvHdzsUmwDVhNHGs0ScUlvPu9uKMqka7wXUwtPXOk6zHye3NsBBcitMNxRfp
BcH+u79vo0GFVQXxXZRpI26IXoKr3LZZbYjPH8fNlcATX7+C30bTQLSVAf6ZDfJV
TT2n12gyE5fReba8TcJdQrwi74YrP8bf9Nwriz1Zk4eiuz00Eo0d/rKSAyqZ+FWL
H338wQ38jV8FZAfPUiObpsmIvyq4xCRblVcviKELCPxx49z+p09O3vP36F/avj0G
otO7skEQdzEwBLOdx3Z0rOGZprRPSNQZ7y6m+9nk/YN4290s5YdadCzuns9usJ6F
kFVACoZznD7PdaZgtDHOXrwvKofmuiNgaGp1TumO76TXGFczCm6eatHP55DPAdW2
eEk/fg9Mfi2AojoOIVbacuQEW2BIRPAK5JuAmr6xHY+jNi3l5HyBkIYBeVbTLZ1f
XctIJdR/fSTOaqAisdYDNH3MsPxWrfCl7/8aZCzhfw2h7BJKI14mf9AbnIJXsCNb
AiP+5hXejTOzpKoKBzIGxIIpbDVsifAsJLYTy5XMrOSuNepjCmGOw55+O0R98m6L
Jof3bsJeVaPa4dqAdn0sqoYDxKl0g8eFNa2x92B5mb3JqH4/gIqMUDtZsA5SMdGB
tKmK9T+X7zVybv4XsawdO4mcFW1GS3q3vSitFT27pLU6WdWHxlzwT5AqL2wRqq+H
U7T0ZOBFZC2RVwy0SMEwxprd9+VEqwF0b/06ze55Nvc2dt0nkYticlxxpQDU7nV5
lZSRFAawzLHVWzagT5pKIApsjoTkwXTt38G3KIKjWT1rONrDy+Zc0t/ysEFqB50M
2ufJmqR+kGt1vXRBOudfsWpMm/6dAk6XsiIBWalJtjc5fn7XZktwN2j12F4R2l7m
fGWWlkZDW24yiY8k0R3mS5tkSkRnBHz5yd0c9/HlRqoQEZH5HKj1IDLOR/Cnyl58
2JEK3tCPd6id9HN0P/SorSCJJGz/R1b3LinKoSw9LKdT9k7D9iks+5aO7nGuuKwa
8YJazRt946DPdG0TcZGwuRcXqlHI6dSU3OHs2V2qiFb6vS7bWVFhIMJKFn0CraU/
R+n2Z32CGfBrsk5dDo9MRQIqxu957L1d3KJxiNp6m1KhPcZCLGpEM2+mI6n/dV9A
51mM3Yy5/bv8S69uElHLoH06uZXGopTTF3lWKfiJy1G458VKtm1KvPAWmKQDq1do
miKlSbI0WlnLHuSQHHwhH/qXkyqt3CkgRac35cVJ8nRfhGFj7Ht+I3QCj4GvLjvl
b4RIvBaZfx9FrAEwSRnxAw9zApu7Cs/F4EZgd+YC9d2Ft+3klML9T1BvtyCXK4hY
lABNhj//ht+aESjPvemYuxnzSV+rWX4CHloRE31Oe8XrYe7Aythom25pb6pEynds
k5gkkWTa/H9SOtfX86vqxrp9jYnpj8axCeZaZaUjM3XuC70+dtT+MNNiiMRlas7n
4gYIL8077EaDbXGtncPq5s2kGWPYLoeyQkQIhomhmjQ1jEkUWsySMhgcf9sVKWtw
k26P+wLru1BGiDwHtbEBnt7gVTPPFZqHTp/ynBU+STjysAEfkY+RN/L7Pd9r6pPv
MBzWZ7QtRwANsEzZRWzrmJaAoTfJ/c+SGAoPUiJ2HdeaIbVzJK3UOujt0ebNebV0
nq8fXEs38sZ9MSewfjCrwHMLswtKGuxak4CS3ZKVjHgbMGN25Wsh1J1AknO5mh1b
VBslWbhvi2H7TXG9W+kWvd+yC9SDm5eAsguyftoCvtAF6vkwrhVTfGW3eBibEQ5e
JegdIbXfV5hCGmI+puQInvH0RUaNsBZoNumrTydujB//fC1gxsZRvmvP0F7F21fc
woY/apDNrXOl4NxxQo3T3kPDdNl/wcGjanCkXOPXY0w7JJxK4U9yZ+nRC7lRekrl
A+Ky7zQKq7EC6vwnp5MqTG2W32NgZFY/m9Fg8AXiYpHTrTAHkFXEGtqiVxuhadmS
kdqYvo9pi9RIRs4a3GcDQjF+7LMtsH2sWb8Mdz8BlHnRTEi6QA9nuLFs82S8gRVU
gw+dDcHLOjcKcj0wK//n2qgGX93wFN2nYTnSadmAAUBAZ5URwrZV2BCq1UOolCII
xbmxbyr8WeGAlyYWevoTkaZt+b8ns/QPMZDAzGhPruVSZZaoXy9ybuEXN14DSUzV
qfNY6txObPV4pQlx+jONgEdyP622NDWJ3pG14odOFyFEi002eSKUXKPvYH1aagpn
nrPnNoSyP7wM+2E5uSoG1xBKNIeBQaEQgxtT2PuWFMxF2RycqfD0OwMoGjQmm+8/
DotkjDqMWZ+G3LymMBncvc04TJJayle9/6HqVMRW1S6I+A7s3k/qdaRqen8GQMaG
5ouyE7cgAXQXtc4LVEiVss4WM+AIFNTf6dJBKpHKIbU7WBsZcTOKhgfOsl95Ygvc
jtFKgFwZ12Ilw4fFRUdICWbCqVgipXnitdXSirbQtQ8ANGuAb35W33LsPitrXlnn
sAdxNDnQ5/n2aVVwRH6S8TVPlRh2LQ0JMuyFoO+HelsliQ9sGQLjdKfYL0yChKe8
gT755VeuvssOGqyA7AkLKtCGiQYGw6aQiZuttMd/BU0mg7Zt62aRPMAHNUJc4XYA
+hFv+1ShGmM6EQU2zO1LBKnR4om5gq9oT/LnJLzDlHvw4WgDggzSUpye/zJJOeLG
xBa6/MBQsmQxi6J7TGOqWnq5GgXEr0DqrQT/UxGcRdKoOPyW+s3vLzDETtOjIKlQ
WVUHtwKQfMmgoylvIt2tQ3mQHKxf4OqLssYYdU+nh0iiNfkBrAuPhAXypcOZ+iu8
oNfiUveS+Bc5brzvLfeAlbKuGQ2IXv1lbYF56qZyyS8sU/t0tTBp0BwnbirrkqJ7
txHu3+pcVJPCatIWdVtfAf/1uvijWAGtOudzI0q0BjGZ+VoAxzM3nG/wfkt2Iv7b
21lhUuWzVVhY1zPnRUmUh3iKeF+EBTGkYi1DGYtq/1E/oYV+L7m4BafIA0VK7Odt
kWdJV43V0O2RvaMiqQo4Ip0kmBDQilw1ePfMVEStiNCS9aZNPpoDszaHPjDv5+Dt
i/u8x6jUwwJ3nkQCpCBfwOB/f8Q1w4gyZOSgAkbzEDwZBbADePEoWPd1ShRszOAR
xKAJp6kkSMLDtiG6syatAZaLKnl3+62tpw0mtzy7633MPlfzqGeBRe5+2CIi00HQ
B9MUyo5QEPyLjuS2f+Y5D5ZU5Xv+OHOAGOQ8lHqHUNKz40AcZn9JlStqBJtQcBGU
kKYcoMkuewiQJn3ny7o1tjz3en/6MrEpDFu3GRsi6oLAVsaDx8aNyN6FZhuI2VW9
egGjMS4pDJ5LSjHP/6V5YBsSn2rbprV4b1OVuGa0dTrzuSyaehjFcN7zEECRRRb7
8xXI6w1ats22p5FfBeyO07lGTi18TL1XR0pwXpvujj2wml5Xm+WKsjM+w6yfMORT
so8HaMHbDyZNY6mUbWoJyRfaHK9Z15SP29EZ3F/mhgtSDxMA1lwzYm6OSruMYvyD
O96te2rFELELsbfi0AAy6va1C1nwdyNE7aqh17IpBFlmQ7hnUPt81/VWKfLs3dD8
rnDTD+NilfNxZhQjp9oOvDBY6AtHcm6I/erVy14qGhJWHOCRYWYY4pFtvM9hkQFu
mAYSaTPRclGk/x3I1fd7OFCbfp3h92kzzQLrskiQzkoVNoJHtpejRtCANXkQT/ry
T25ME0nBkT27vHDR1WJIJWvA7KK3wZbV9pNRPUb/sTjzdI/fn9jSFJ3yGDr7iYlE
Ame7wZfAFOpWiKGU1GSiRiqpbdINOFfwFEUBy9v7GScJhcr2lbag12htLyNiR1UK
GVTP90jTocNp7Up6aF2WGfi4RG7SoeX78gGjquyRLtcCf3LWzNxqbflCiXHhPNKD
K/sB091ekP3De+Wa1thiEK0QDomgGLTKkTUgBSoZRVIvR/C9WBSwWHpZ9GGW/LoV
Y9ag9GXFvkNLkseiuhu/L5CfrOKqUvWxoD761tIKx9Y2fRLJBvVqTzoCF2N5iWVR
mnSU/j0FfMaDnZkDRDRW7PgHxlO/BAiQFMOBWFVxYpdCQHtLcAB/DFTSq95G9ClR
IYn8QbTPH853O0zI2MpcMjEW475S/udqhAsI41MAx8b2xY70rK8040Jy8AlbgT5P
HMgEcaPHmavH84oZdJCGk+nvV3rVjrGWbOqmmvHi01Aq4XqDBtF7al/SWwxRMzAT
Fu0MxduIh0ltFEXzMEot/56xBiiXEHUF83y+bRIdNVbLHLUiBR3VxSC56WMqRZOb
1vq+U82LODX2qXxffa3v9XlYNGufdwd+Oi9KCy5dgPEA0PyirX6n7rdEk5BXaV/b
JcEHIAWSrlu2QIFPnzaKexdDMZmodoWs2y+RyobtnEDh1j1NDveHr3AYiQOqT2Zn
dG86LMxfWeu2zNhvKb/77qRsr1RLwHvTJ9gr+HgWKquYZprc5G0zjSPZ5t538Tln
qwkl98k8DM6lwCaNCfKqmspiCtbvQ88SZ7f8Nc9NArtfgRjdRmdiofvq0bvQWFHE
uZ+9L/YRR4TjLVzWelITxGL7cj0H5sL5vf64JdCdNEXDut9cvP6rgCv/20Hdj2db
bd/jwn9/T+l0o9bAlfQOXAXYr+q3akeBMJ6rHpIyREptDBta2fLYmWkaXmfDxtwM
mao78X13o9noZuEyd83bI0sYxDprCA98agGFd3t754JTP9GNx2Ursw2wYLz8mOJU
fSPR2ZVHIk9ncFU9stYb3YROEmmQD0OTXv+Hu4GDY7hXj/cuny8sCJNG5c8Cg3C3
VmuPJKOMgLOyqCj+KdDPpGYVmXR/D8KS61wS7LdXgalq0Ogcrqq3pXFEOuXU/OK/
98eQAT/IF9cYWWOnyXnTo6Xr5Yn2gzBcL46X+QSezbL7Fx5Gvhg1p4wJOmxE+OCL
ROFmAfcpPeeOQkhNz6T+8hjygyXpEbPcZhkle8v9jItOuBxvETB56LV5mrK4ao9E
MNZcx2PA0YedUd4+uNy7qKG9v10npClDQzVHv6PUZQ67pOLsVIcVdlHexunB9en3
g3aVaF8Voz8lgcPXOrdWzxJv/JHvvZOJ4r6QDqziSZkhBL+IUeeuuS5eUH/rZGdP
0kzqkeY/Jq2OCvAQAO82FtMRQUeogx8XMYEPFNYSu947hKP5WUjUrbQcAMEI5euJ
3C0INakAb0WNLa2K44Mp5wHNc4PcrjsxFh0tnYK4dIa5+HSMb6WpGAVT3NqfSeUi
MHW8DGBqrFXksp5O9jiJuSb0hXN3FSC8c0tyXNIeJqvL9dP2SiUNuvu41Ugb4IQE
6znwcreqCTypocRZgJbVKwgimNmD3PrtDex1jLG/DLPmpErDFBAO6QstMJ/QXhvd
vUeY4he+2zOkDTvnNO+CgGs1mc1qb/J2yWZR+NofUFiiZd/L7yf2z5F2SsU91Xxe
rzGo/SyQKecbIBgROXMhhugAJ1HI5z6L+vlVH4Q0Ml4+kdoRIt+/hRuZ4Ur18kpr
1JuyAZWkYIS86mpgk5BJF5EmKo9/6lMLhhY1L5BVXnljLbAfRsikcGqWXN0PVqUp
0n9Pi92QqqKdAR5E2mVv+I9IconiR5Rr6SJr1YExPOjQKG/U2e2IoGtmxXJJVgwa
jdQ2yvjvjBRmYFoaWx22EPHkPLyXp3X0AaLKND1zLwsIgwmGcDLy385XQpijL1Va
Rt8GSA9dJskADJ6iArenauCRn51GSkBJfwIz186KK6NvaMyHqsUnAz8ISafSQij4
14JD9P0RimBXBNaIg+IOEPhjSDnPgjgRAn18c0wtIZoNXg7z8viAMs+/qBYalUoe
LHZMbx5pIGNAAMKLkRuht7Zdj7skHsNiLy9lVNhTR8K7vnQpEbINaSYlL+4s92kg
IvP+uRDFqwW7ABaE5EyUV3M5YKnBREfQm7/iVh16g3PH0vU5sI2X2ixI5MkFabeO
VqklZprDOgvToQGJxf9PIkq+3kIa7xCIvBhZTWMONUmpbqgdRVAoVYn7839bN2fT
Z6wYpAFHou53xVGmyKRqg8AhO8+qqFr9bUHTHvyUMRmiZZ43t07aG7uv/MUq9m35
Nh6WUhtMWS7Z/SGLFw4AiQDy5V8nd41tt+A2b5X+L0iwTz0CLWuOAnkHJUphpru/
Qf5NYlRkFp62JsGwXd6kl2QgH8HDzi91lYH/Gl1atRIOIAzOo0xbEGJOLRo6ajws
yywiQkGjLjX6MzbysfUvmoDqhnbEaom6LxjPLpnxFeEMLsqukOEJeEbvHhm+Uelo
hO4ccyXEfZ32rELZWFXCZEaoD1pLluRRVuuYZ00ZOJF/2QGVhMNcihXtfBfGUNgY
WN2tmqgRX0cpYMNK7UhRfRjE5UNvGQASxCo+fLPpnseZEUk2WkXCxJ+85hFU1ZAs
ukh84G3dNCRoIMxhTZjgEo3GrFzx0SAaXr4eNNKkIKDCMKuP6nHUgq+JKPSonkXS
o2M9rts5I/QkLYy7QVdc3PoVFx2l8PmN0+s5Y9o6up/4U7P5/XdWMeycF7ESFCTy
I+VvK9JtZtrYLyx3k/8zMFouUz0ut59mWR+r6oNUbL/Ngl4MheMZlf9KuHsvr74I
aQpsPZXqNXJcdgBPKszqev4O0onOdyellY/shzZFomGIfzNmAPQqg4T+YU6y1wBK
m4TmnNZCXPTqNV415dizy/cn/swerRVbvEAmLJMACSluCm9KbV2urmqH3KICQdjj
oAd+PWA0Ik/H3UarIpp8P6LYJ8jmpJt/eXAJAwVC4FDrw7ZYVYgCLVGckmXPTlnz
V7X2L+esfrHEE2/2Jc7ssGykyK+pBnzmXzjY48HEla0sTFTisfhxSguXOEenGWLd
g4MqVRiy2Ncr0I5RIaH2kZ56qX0hR3ECalethL9X0tnEtY8dPuI4HlytHQKX3mJu
flQYVHoHChWdIBVIEUxVfl0MmfXF+zC2ZJA2xb2tBA4uWSjJmL79c2DX7pjOYykF
CN/U+WYWaLWP3H3lvfEP0nLUA4J7jWYXX4XG4zlwrgEF7VPcTcpPEcSdLrlSeiLj
+jz1Q5ki67c7Pljn/mccKLL6j9ilWvyPkeg/7aE66Mdk3McK3N0wWiPXzrI5Zjs0
RbrAbHomtN5LfwxoxUvh5eCNVgouVR+Uh9bzLWijorKqZAbkExu1lOiHG2FTtp02
J90xJexkhd2s02D+QYeJi3s2bve/HGK3ai2RI1hNXp6BBqQX5XzkCp9KYtk6kIEO
SRtlX1yyJqbyYT6PQiaxFJbs/VtdSYVg1sI/ktss3AGOwqtcpmLlBNJa8Q9vP8QZ
ZWBXydmqDAMr11i8SnGu2ZXKUla9e8jJZDDiV6B9acDi+Mx7pTOYgLDEJqAb41Ds
WmRHluqn0gWjwtrkz57i8eyfB74z1Gqga3Y22IUxGq89qsybx9jyESN/TsISqcec
Ntm2SZSAFX69ztFochzl4jinHK14aJ+9ABla4LT83ejKkT1CJZQIQ1TG1w9ORVuE
gIG9s1I4Mu4J341NgWgiA7Kx1IvmbdGRuxB6xlacecWSxco1B19WCgayCRkbCGlK
qU1S+hWeIIy3Pm+7LTtGdRfjw1FQzm7FBYfJHt7zqziIKdLQ+xWQU/PLL99j23nA
RKRvH2hvr0iRw5v3uNUTvuCrILjUjaqdCj03npwcAU+KvKoExOGFnRI8oCEETV3y
BbSMhi+o8Gc+FgWCrNLUXmxDV8qRCsfa8HKdTfRasP7TITwN7tbxiI3o3rmf51DT
WEVJ28Sgmw+JeJ4JrTCGwpNgi5JM1wKOz21mdaeDdC1UsWO/GSECT7CIyUoOqcDt
q4MIAzbMaPlZsRRU9E5NpnjmbVp0RjepWtV4Xg7+xJqd1j4RVeqGG1vSxZBu2kHC
Dba79uPLFc9w4Kn2ldZUawRjyTaiYUK79nCKOGPWjk4q2d2FVaS1pmHzC8rpZFZ/
cGUkx87ZwT21zuWR1wIaaTYBLMJtSjPiA7lhE9B60/afXRUCfG006VMv1XL8iDzV
4D//TbOml2vCJtLKTCRtYfLvjGVxZpEUxMBuDTv7dKX2LApKHpbw1bYZyoRxgVrd
bGANt4FgoDhzT+6mtEZR6qtnJmQ0Z0RWWR45KFuCuoZQxFnu2mv2evS/NpcsJFDj
jl1Wr+gh6g/7w+zZS5egesztEwP0APvoO6rKtJ6JqX05AgUG6cbY/U4PSZrJg/KC
40F4PhRoB+yQ+H0JwTcDLdF9MlPxztMkODvFiTM9oC8RRVKHpHvZe2g+lnTYabTJ
H0E8ZcqCvKexCPCvozFegRH7lbFlDYnAiSMwtI9+yEspv5D8019XYaPcNrtxcPhK
+wjb8dTZuNg7mmVvec2g+AddQDZTWE7V2e+hFZLgJU4QfU2jD0ujlxCMkkReeQve
891MV7YWjw35Y9dbTYUtK1yqzBg0qa0zt0IipWmpPeBYI9DaqoZ2cPq8ETBTeVCs
7qfYGzti1rRlxJJM2ifpuHZwfPPZrg09fkydZ8KWeoeYgU4fnUBtlkD4Fgb1TaL9
weGhDA5PxjV13kO7U5+3lZeQ/Y6Qm3VmErZSxZQoQBr+ozGDRgU0ZGvIMuh7I+Er
Xm4BKks10aS/GaSV56rY8w/lAxpLwamL/HK88egkbs+Xmj+UfsvnozIuXIPUES0a
VBRJTQKH9tVNp8ShFYu+6Buxo4RTXveA8I4ZBR73iMiSWm9fIWSPsqwOAJw2cbw5
l2NK895kXdSYBG45w465N93px/nbLUby/r0+cgaeiPPL+CTBSE/O/bMZpvZ2XvMa
YczTDREMkvUd3qXD4Kt5MmxaN7h43mxtez5w02+MkLycHpmuhaf457H3SLmjfCmF
KQn6WnNf8QXq5aAdUlup3C1Irg7dK8HB1gm/K7XZXKudw2ergvcI6S7Ahh7NoO37
GIGv3CFYQ63Zrxx/3Wwh5VKiSXhYUnz5PCSPIQ7eGwv71XVLUAbWOupqV70+3q8m
8xJeldDlUHgqHZpx7ICOIJtgSbOtDz4+8YGGMg09h2FU6YExtnvOXuEyisQ/N+3M
VgAdDct5LS1Abl41d5JDlo/TuZuo2BP3BCCrAdi5sm5Dk/IJCsJiX+jauqnHvBE8
6om8i38FkLLAXtbEr8FthTcxLVTxR0GZ1kQfT1NN69V1PFM8WRgpPXUTVSZC8WYg
CLOkpyeMEm+7h6zh2LiKi2ldo3EXefO3TUGuP10g7b2McUOkCsXFB3EEKkqPOWVQ
2gUdHsQRaYImwkFpwux839KUPeq5N1u2FQ3nge41NKq76mPXO7mk61JIX91p7LhH
r8hDu8ncDRdne0/YSzVKBqjK9lTnS3rQTV4vO6EEa9fLvHyKm8q0frnFuQo78aRV
Ye73uzxnnyjAqnWeYRba9IZnlEjJNUiCXmjsKBy5cad+LmE5fJTtcwxc+I1yVCc5
3F7nnP9mbC6z3vYJzT3wr64vTJFRyu92CqO3onhh47NTCiQq81ENgfSi3kAoVEDR
t1lAQN/pp2YpwCDG3jgZ8QjDNkP0BzzpEcaf5Wq+DCNQcA4QEVDK3XbH/FgV8rg5
OIGD7MzZJvbaMsMl0xabgxfovC5kSCuLjKwgPOfLqgTg8zEqIc+VyI4DLrAT3VRn
ThZyrYDSSnWVUJf6Km2SOlST8JGuGN+UToR7wFpjVQ6Q5R1+U+1XJWPcmLsZc+kJ
nZ3HFH617mIrViafFt7SdEqIQ5iYqwffT7mSt9Ux3yoRfX75I7ulzikAi/3pCkSG
pyS1wWA6UMANMvxUMpMFibeq5yTP4P5LceDhWzP86s/Cik5fmd8onKw0tn+jwMgT
cZzsHwievY1Y7q5n9q62srsnlXud0Hh+TPpAwKNbiYG4Bxol6B6wqxXIlizUBID8
6lQtQak2HPY3YoveUhNuOD06RwVRW6CpM/LiVMz4NQf5kl6LinGhjZaw/3WYfUOV
hdy49ppLmS5fETiqXYq07HpTYP2e9+yVRI9mJxu0wHhgnqpaA5TthvzJd65649As
rSPp5JCbrlxdKc3uNzWTI6QtqNByqM40KuV+/eXPOykuatMiNvP22ACZhFDGN9iy
0jKpyjlwQv1+5xVvJMGA+b/UuQ2mxKlo4JvLF8DMImL0FZB62Sa4ZeaZUuo6ZR52
LFeM+7USmszksgZJGaRvWj1fHhiJfKUv8Go9DGHAT4NX/T8mlqtEAHzW4HOqTYA2
qJYnOGNgX4ryBt4kwjioH1rhG3DimyJRgPXc6WbFBdqJ+Mu9tgzJrG5nEoELh9QC
PsAZOyJoJZQ9rQa12OTiO477abacZxXXW1F8ZdDIPL5ELOeHsFl3WEPUH29ddwTd
WpV9luMB5bA0NsbwRK10s869F1/EJpxqEvdTiUySnwvfNZAzmNIW9wE8/15XLePW
cFn6hCtOKacm3VQsV2T+Q2AxybqG3SobdpQJb1JVDJWznP9cg7bnkqUqThVfQjbm
spdTvS4H1CQmR98ehbiRr8cgmTH6M2EGZtmoXWCbZHojkrkBrWTWI19Ju/JF17As
I/GmEeJJ1dqlOlelx1XIWUdsXyOnAD/gRhqEN8/7jypkYMsgSs8974aIWEnJkQ91
CgFny2eEvimFo4ooHf2qniw1d0U6mGUE+ZDrJ+cyHlpQgFURBWeeoJBOt3hYqCFd
vlwDnLgcr3BSIrdZ+YBFi/znyaalEiwJl8d80W9IM+Ztt7ix1jI5gZTpF1SvFT5l
WrOqh8mOH5jRLIRdpOwSxKDm5jBpXR7F8N4hC6SljzprCLy6KokUeh+g5lvXlXPv
4A4SGk7nQEtF4qyr2QdSvxMMYLcr5MFUH9Cs4vt3w2G76SHzN+/EdpE5D6+BAxSz
81KmeNH0X3z0rN9Y5AwJtWNkjywhux5Mb0RV5jbi1eQDlFM4VXh77GyajLQ/inSn
f6U3OdXQyv/v2YYD+zZrmeWFsI5NQw9vgYO/S4dpD1PKnQ29SKJZg/fLnqhoT1qI
XQYTaaSNIAHNut+HM75OauowR3zOHr57DFfgFO0sQllpT2Fknx2ab4KVpuwWEBuK
yprNXes6c3dMlQBxLcfSZm449AD4MtWB7o0abCPcN2qvNL069cDYpDtMwOHdlcId
/YOhS9IT1h6KLhiKBbOZdP4XqPP505MTGncC8jP6H2B/oJiY0R4fUnfVO6yJy+Zw
3iXnK6jAp+kT23eWfmYKnYZG/VBmiCvVCzTH06u3VpJvG4vEU2CDz2z5E24YMC6X
nS7+ZjUGyTR+jgMkfwhf8puec75wRHhD7W4haB5Vp0fQIqtK7V4gKWW73tyjAwS6
MYxPf41qSU1UcL+9uWAuISNh27W2PcpOeyvRm/uFaFofQddB4IoAAnuF15VGFrbr
lDCkE6Ylb0xmtl42UCLvwQ9VaJhoU/HVPVplwPQWBG4/IUU/07DAzRuxf8oIslxR
a2b3R6j7SBww0lR22F4zmJS+hoZawEUJ3vtDLd6UsA0OHdTU4tC8YKno7meZphwC
xRPS7BZWwJzKBdWPp7/81t196ufqySn2+cPuzvUXK4VePHvs670MS2wwaS1z4oQB
KCZ29tv9vWw2txQ+LWXsAf5QogasPeA3uFR9geANKgoPt6nH/f7j+VLLBW5O4iQX
bqxXCYW9nfOvX2gYdcu0IzFdYunnXy4GrTQD+O5+YXzPpiCkLtQw3gbpwdzmFrtM
TWgXTZ8vcxPe++6cNBBo1HAlEKvJ2LFq8z4hZ/jBskBj8upSSe1nAxIJZhOVlLGV
/wfQoR07/xGy9aNaiUaoCf8ROqGIqk9XEU1WnWGTGblfGQootJshasRugm9BIP2W
pHaxgxgNPFiNSlG5EMAc63RQOw+rwH9YNFB/Dj4/a+vPcK+2Rb3m3NEReDEbBEdg
Vu4TVmCIVtIa0dlVeG/X1hxQbkEfUJrcGBk2E5WyKm1JEFlfjUfaYGJ/4n+DdPP0
IhU+r73RjGXZrJQPKekMyiwh54SJjc0LSvYw1R32yPHwK3dEJHS2RhKeyd98cMej
BUnZX8+hQdXY4ejPfQQA3d+mQrmfNOxPdR2T1gRNVC28EeqkFv0OMvxo5D7/avGc
f7HnWO9TKKsbb7yBikFlCcmXpgOygavQMCVx9x1ajejAbRZFPTFmdON5p0BWEUQp
zpGKt//G/LpVsK1/DoxZ69Bsr0kk3GhDT0hIJ7i8iOqDAllRgCqPfTf2Ui9JF7h4
wYVpLQ4dNJt9rFAqYpbD17UsUJXvx1m9RV0Vp+5SmoqbC6JkJEh8xt+4EhXNF/YH
/GDWZBtFClDTNnAZi7tJ89U32nXDZnQ7yUQ7bXshLfHjl7JR0Xyn1FWBr+LZaV7Z
zO2SVIJ2ykLmbWhgJuLD2k6eX18XkgXK20eGTgC/maF2vgvQGQihFsi+Ty6L+NeH
J3zxRGDmPf1wHMfO/MwdrFxLeiEPvx5Fzlq1+lOzmxRHqfgKXh7crYgpKvwxCwzD
/YQI4VllJPusSXy7mWX/VIajZexn4HlijXZhKy2R8uiRn2sKfYVdogFWbyN8fvBS
u9akNw1Dj7J8YvcuceA/TzKQgIIzZjNRj7kqFX+MLzPoYxhMbHJgY09+pOfoU81k
HhQXmLle21rQaEWUOK45mocQbPec+1+0nWWQ6ttuFs2Pl9mQ9kv1ZIMsrXh92pmp
j0391K/IONy12k2kooyYpH4N1zCkfgV458FQ1nl0EG2mMP+GaSnfyMOC2Ktmz/dt
zPclVk4BJz1tqqO5yDeIWGQEBjUSs+FVkO2IAc2WFrcaHsJKCzfuJey934cT8hVd
zhxMesFRS7c3PJ17EVa9+M2D1zlwi80ZyKdyd1wlCRdatrWwBY+Xl8fzHEcUcJd1
jL8tP1yWOnrRBDbtFmHpJFy8n4GOWWbpM2Hp+ctZrFgd2femmiG1djoF7wbWX3QN
7FQz4rWeF9pphQwpkWX6i9QNojnUan4OuxU80UZeWZAepex20t2cXn9WuGfNPhSG
frtHkYD/SPhBUF68EBt/M9Dc63yyi9p9vtziRfHaqJJRmnJiFSvUPdEePTF+Plcj
VX91KICex7MmFWyJ5r96muJkPgoNsNPTDLqiwsEOxAwN8iyn9RG6FDGbKNf9gw+y
8F6Ww4hrlXVrd4YGZJsEL6WQsG691AoA1ToY7HOd2FJ3kDWPAn59H9dWuRkIm8rB
mA0LI3AKrDt/6uO1jyLI7unVCaXNOHE5mLLl0hKQwL7MCn4hMfB1iEiS1mWnvl2r
CeAxHiU/FWFDf8c0iTrPjuHBf1EyG0umaRn5UhMaVVQryCTPYDhHghTLrWdtuDqH
rOQdhStanCxEiVn6/qnSC6wxVgS1MPwLVCotYGHG08u9gfFcV4XCde74kQs5Yb2V
nlGYBkRP1mF1erkjkniXtUDQS5/RgL3hUAxflPHc688Bb5Aoiz9Dy+Bbj+u8EJ5a
KvahrbVUPCDb36HUJevqLO4D64PX6HCrJ9tMvl1eaLlKmJhppd13QVNZEo87LM9B
/CWdHIgdHfDfFJqa8V5FqHdzU13Vn2E/EnrLQOZjmBB+FiyjS9dKt61rVidwi8jV
Wi/LtcbnkCVSH5OkwEDOosdq1qIyKRfFNtr30fAfXnlrfDgAonNo4r7xkoyL90mo
lfmZNH0w0v0MIvq0ex0robbvqge63qNytwsoQLJY01atzbRHNkLOFz7V5Dex44N0
Vv1CipwNnK9p1EE+418NCifXfeGr/gw1RJ5lz4fZF79+JwA1WWofh3MQZ9ArZw/T
6o9+LNPoYLEkfhtfoiYM9GIKonAF0CqbZ6W5kqkh7MX1XxlirxLVeo0xiR5U9M/A
vlqYtM6Y14VXUedHva0Ne0qMy1/cqEeZuHCYxZZkecjuCvGzVPT745jcBjTxqLJI
twsQZa+deV4DQSQjSaXzkDRTQF5F274ZQlIlOQTKCpf9xUV0wPheyI6WKg1v+rYu
gU4hUX8sGGDvG3j5Pl5kIJPE5W8d8zNgljg9O9xS1ehfkRovcOMpIXj+y9xYI2kt
ts28o4t3L8LXIQ9dgGtlXX1oRN67jOgahI8j2OU6K1GJORR0NPbRFlnoitGs8N/Y
swjo/17QP0Drk/9Kx3B4s6lcZVhFcU64x/j10j02HaF3WuVkDEr/8hNtYQ4nxBpm
uDv+cPyD6XZgHeRSb1Cqszth7CtoL7DRf4wBFV9ysc8VvWSMFgYq42OFPHHb2t0E
iWK/tsSOj4nGlP7/IyhqYgD7Qf7Da694Go9LaNqgb6Q9ysH2Ls/7nhOmx5zO/s6B
t5B9W3RyN08QebLDF0dLWkQV9oaRXCl1zhA7UCpFESqm8tStB8bTSmp34BkubVSb
Tv6UD8CqxQaXJdQxBDk4JWT9h/PTgLipG84Emc3cP+b9nHo/RYCMh6cfMocTWpVX
KwNhUWVCbbxLq6xxX2QChUW0yhqAeFI0baQXPoEyl8CIc1JphuIHE42HlkhOg8Zv
EbENe8QLm5ZevlrkpoF5OE0/eNGRr41eVY8NqfX/QrRYUnKYN2AdxiOdPQD2gRu5
TAQsWlBluEgkqRBZdshA+JmZOs0FPzMMsF/7N3AoSyqmz9fIXMuqJufF5emVkjxu
+EyCuvHPulHQFE08o7G2TAMKxOxYsQmnMinV2dyAJWCB7TUoUD0PRBIzt72XmZYB
9jFt2DrGRrwH7ig7MjUIuPdcSZbZwJGV/Fubz0z4F6aAwHxA+xrepqiXeIy/yB2U
/eS6iuWKiPTlv2/y9ojWBu4EOToPghB++L3IVpFBD7W4uD1Yj1g3Qx6QMnv1tdhN
GEV/S6BbyhpVEhXZKhayw8s3HRU4mdTRFl3CFLIMdFp2x54JXyb3KPQcPEFaB+pW
sp58mNpsmvc+whwGXO4flr8luouxXjN7c2NJPZbpLCz6TFuGaBltWJPCqC0CTlAe
+Zto+eEmJnrA6mXMAb/utmo9xErqsiA2b39t2uA2ttj3+03q7xA5INh4t6lzL4C6
dE3wlMXy3F4A9vRVT19/NcWLbux+dUA8llu9kLSaSqQUcU4UbQbZikoEAyQIzl0n
ZkAkmEzW2mJyAeWv3SzFEiG4kqv+PN5Qup3Av8uCCvDL1nIXZaeDizVmlikNQlwV
Iq8A4ktx2gFr2Qz8p/N/o3aAGac1LWWBVKOBJwV0HlG/zcT5XxiVl6Wm3w0boIcA
E7YIV5u6KKdXyP/Z0nPN8j6dROJvanulslh1jtcWlxPNDneOJnICoPXl7WzYdUYz
ogXaeqyjl0NqBHUqeusNaOmETZgUoAR+xTaSouxyTLuZWWCYtzYLGA3S26/QQETP
BAxLZ7gBFZGzyqW64jONe8gtPyo8j30NcyLHLfuGrzaLAbvKSwpT3lBr2ZKH3lux
q3CNoGNGVNbx66k8Cq6zpEK0YBjwa5GRJDj+xIhRSE2jd3NQfV8BuAe/aUAwE/o7
6Q9NKgD0atjg6iVLRO31rbLJRMtzj1rA8ermPvVApuuFOuM9r8XbeNKUPTBePkPM
2Pm7z2sUKRk/LPiE1IU6pgovZzB/zn/On7pUeOsNht7+y+N9kvuq7sFm7KlQe0Qz
q2SOyls8fJsWPN7A4Pps9ooyoR5obzORwcUY3d9tfvwZGLoDqOm4mSk9+8AnUsGC
P53J1aeBr+8xjz/GqP8of6ooNOAROWzjMBkRp4V9T8gPdF9isCO0VVSibQwnR53H
Kf3di/4dZpUfdXapfB3ihg9RSGnvdvMUS+JH35UPKTBbob+qf7STT9gQmS1ufbXF
5EY8KobYXlNkQdJ+a+9dMPBjY55IUaczV65vEk37tovlwvga506jkf2rEbPXbf6W
Cs1XD6nPjal4SzzXJ6oJ7VwW+CzkKvG/msIADkCaYRYSYL+ndVtiBCJz2yAemh3M
XyOmG3te1G6e6pMIVeTjzv98DsbJurr8UdE891/cPA12BF/dJiATkNdS2mzd2cnF
Nvxa/8+JkKJq1/i5RAywrpd6h/KOqDy0V/80gKuXJfFbyYdbtai1wz1NsUKKb+5A
R3cICF99dlY/i9Ur43HqOJz4XAB1UL7TWVSDYR0qKYZSlE6vYcs1/iQczD8BisdD
JWJ3pJwP9vy5vKutKeAVMQdoadInRSZwgTfqztr70oQqcoX7TpE/8QsK+PnF68jx
oLPBTb/n4C/UETrYa1/Qw+gZqcPMCTNPzv600Bk7HYAUfE+qQtFptUzk02vLIZfM
Err+iJK5b6Bms8Z5K0+8qwtiULJEwdXcjp5oV8spt2uVkO6yow15sdch9We+WltF
kGEuL/1xOYU+ypjC9Nkf+oYT1gicZKPRZ2fHqc/z8z/zr5qAkl+HL6jd42TpU+nt
D1aSCHzpoPZcX68YzK3gqivSrdAg9fGh7BYe0CdTsT1+bYvI4Z3gBy00xTKlDzqn
wNKw6WCTKIjchFBOaU7Nl0mDvtKV4nXxvxXgvDwwQxdOKVwbIEXREk4vR8W+ZwRl
BWhM/r8T/fT5zjO6ADHiA35UM2EcnhF7X41lJ9RsqZYFDmvzKzuMSHmRyQGRIXpp
BQMw4QuB+94zOSk44X96cpex+o/IPC9dzAhYRbp9zLwukGpCL3WTpdyvV/+AcBUA
aexQyJPxKk5rz2a2WCw1FvfdnjkRiiSXj2rFIuD8DhANceKY1SC/8GeZjLqmh65r
H5g2CMIg/tqCTj1IvomPcoCWTcMhILUBzBvczOpWyqH9Dgfm+ho6Ce1fCx18GW0h
6jf9ayAahz84mBF0enUMabh+cyS6VSIDgdKySMjXZYpJJV5L+wQ4Sdxxi/787pV0
ymoBnCmIethtYo+cPY/wY+287Osf+24KEMqk4UGBt/PDNCvgbmpLSlwtJIvNaWw8
QGXtCPN6+4vhBqHHu64faZRJK7JickGdJvEs9pUhETRUufAehCQBIZyLv3YnDgqL
oFSEHApnISZmmcGn/mWw0mLTvfpIwMTNh7r19KGF0Lkior8Fse7ySG5oRg1KVZbu
xx/lmBEbajfJOVms1YOqjwDmsfm9547xqVlKj18lnCh1KhNb7O3DSRChWVaGMa5Y
fTsNrkqMumRAOSxQNisn5ob9nIk94o7PDNpbknrrMRO4uE8YZXcj7aZLqtE4ROLq
SKSuPr1CnFeNnsnQ1ulWHCefE5LkqSzjudK5y2p/fm1awmNS6JTRWqGcdv9+8xuG
R2ivuxyMYma1G+OjjLuCOxpprh+pTjLztnwBQatbe4a/abF23+rtWIjgVd6QUleo
GeI1XawZMRStFslUmbvwycgJmetSgP0BrtkWVFm823qsSFj//8qzndjSsepr3TIi
jNlTdMpL/vC/gX18vN2dOCudqJ830qfGUMqIZugJFJUVsmwXIQ9D9SosYpnfcQj9
DgoDUvGFj/qZ6Q5Tmhp/epfA+52hRqe5DlfVflz1h8XtEDkSHtN98W+f5LYUFgtN
TwZ1TLrPnbui7DwfLLL332+PR+E4Y/cvGqj/5vvTTGNPMT+XmRd3RFbWi3GuAi1L
a7q/5SuVg59flR1x3NNBNRiIm4rjov16v97GwJrnZIoc4XDeXkxKJqsREekt2I/Z
h56wgrZ0hROJSwwzInHrBvpGoib6h29OtszfAehdDGszRLZwxbG8LYY/R/A14Eub
GE+z7arf3YiT+wcgnkVg3TMOkE6pr3iuyVnhMs3KXTyB7BrXbtvKf0JA+GI8GSZG
p8vw9G/5cvyZxi9hXq/rQZGXaCE8NeZK1PPV33khMYT4GiVlbXy7Hq6wh1iXzX4H
79MFdDU8TyRXAzrumgdJI43ZtppKMsvu25xLAvXxIQlqEwkgTP5fx+1i5wNRmLwz
lzzqO/zAKUaPDFjEVQkhsYD2Xt9fZ/sqyFDT6kD6WPEACLtEUKjNNWdfzvuPOGUy
kzjgQMYg1Pcs4RAd09Sz+a6zydR464DfdsZbGE/GQAQDH/eapwnMKUOfCBzRFNEd
lwwWqsI4P8zA1dOVJASwNDadpZL5fp1sjWnQ5kUZRCPB+SwIuUUa/ItkGvg/Y2Vn
XPf4/GFKXX91JtuNxXLoN2N2dLgzVPAFo9kZ4SDa++zOB2DT5Vdbfqqk6ammjTjO
qfsbyPpmSwGilpQdaO/6gDCLLh3QCZZCBHYtAFV6nOAomk2jNSZJQ50RVlk5m0rB
rK8NkS2etZUQv0O5MJxVbSlm0G/j/w1NrhX9qCXV+bNlPekCrOVJ1RWrsbtOGyz4
o7CHC+3qbQGbQzjuEboEl/WHWqp5K++Y1qdPkN4HfFik7RS1IfIJ5mPAk6CCH5+y
j8EpmYd78maFQurp32IgXLX8MoP3BAmY1SGJFmxGaMbI5ALJfIkun0ibNnYZFfoQ
Z3UGt4vqTFhteSRiJZIrKg9RBWp4xkP5am0YzHmCpCqz1fwklLVzXaPJKPVonxDD
7RvdWIQUXnxvQFBPdaBKdJ0sZf/0ve1m8Voo3aSp2X2HHEPiRobvVgXME6SqJaC2
fD6arnGMgfzzdZwxqe36hW4oZOqf1vVI2t85V8aICU0ONjU+J3kGQxynbKt+td88
hXqX2YBJhKgJgOmjkQtgMZjRCGz16f/TymZ8Km1Zbg9zrQzNHbEJXxik5WpNLzz5
S9d/1l6YGT8zMADCxTJUJdI1BtHVo2bgJsMBgcYWB384TGHjpY+MVnJJiC6LDyWl
eQ14NZZhhhF+wka4wiuyi1VLTEt7N2SBLUdBEI4Wia8M2Zi9a/Ioc4xQOQb1DcEj
GZtsou7oR/EFE21ssuZvskohzbt/hjCJf50FX6WLHlH1ftA4g0Fo9LBEMgg357Y5
UNbG0NkM4Muupzo9Kp3n+2n3poxK9uGtIOFkEZoXF2RMjPqAnvKiCGzPu970DFL8
bCeGsWqDCXvswxy8GDRIsgtgiOmznHMnUuWJ/RZQ843NcpIGse8X+Pg1bpwAUfxN
gxgiBs508JfBzWHAs+JVwm3LaymgjpJuqiAg4cBfPv+o4gWX2FuZsltC5pqyt0zb
Gy2UHQHSNZMwqt86VKEICibCUszQzaPwtOpimca3RQq5Ib32GqgsT8todG+For0Z
dE2KwJkHjCpcBZqrGwzKXJeSxqFR5BMGyubXXj2W9RhP73VMjnegiS3ScddlA3W+
QJJBWiap40Kt1LlCr5mtZYlo9RlJP2V/uL3obIUXlzrXr5ohTB7jeXek5eJ0/5EY
tJjCi7v1KoYOoFj9JT9fdDob/QTomebOam1MdFoauFAfepN5pJ6nOatON5qs0+AT
/4DVGzGL+NR5DuQRbfyo74pR3qh8NCp2Y/u8el/3VhamclMacOXKpDL85wQQiP7Z
n8hHpI6idk2/r+afGs315kRrldIDka70wJOzzJob9gSLeIzKoBTXoMlaItevXVaW
rvIUVDp9UZ/QqwVSt+u1FF7VzN4uk7LrgVzW7cS3ccPlnS5b1QXyaa88WYgNM8jj
PoHA+LngKYsv4HdPUPKl/3yLkv6rqCYaiNi3jYkO5bhHdGlOE6gRQsHLlU58HPzu
s+QPzn/SVt9TTxto6VUthln8bLq/YfwSNcdwTcFQhD6mhSLAsaEW+/+wfzdhyz8o
kd+8QaWIXkVZmoI996hzucdp05snGBMj7JGapYZzBEgViuGQXQ5O7vF5QZHn99kx
Cm8JOd90H8s7GoJ7X14SJNkq2dE68xSmaH39qrzZayA84Ne6uHieR5QgW4AIvrGj
ZJe28T124HqI5QA76ktjyLoxU4qmzbU67A6mh/HXUwLDE/Z1P/v3YyIKcZ6l5odT
OkO4dmmk9P1IO+q9mXBi9POizVKtHIBCGpifLy1c9wBwz9ZD6KgrrTLmY7wCXmA1
bNm1muGtA8o1QulzBlqW9ENxJIwc986CyBXs+HZdc9m0KnWXqx6hg4BXx5EG7Yv1
IVJlBHi5Gs1QV36g0dyto9pwnfeVgJJ6IV8mej6Tfhd1eA3TL97lOU5OgIBgBghT
fXx6A3pSR6AzomXV1iofyoiNhioQBZFZ0RXoK7R7z9PlRC55nRuOKRbwIjrdWIGC
Tdt0BUVR1TpsfRZf0tc4zKNOseJ9cSAqXQQceO3nDYdR3XyTP4n/FRY79GsIo6mb
TAl75+7NFoUXclsyrwQ8eQk71vPIMdVPOetr9e1gfUUKP47rcs5GR6DYgve1b3y1
7XEKnm8Cu+sfgJL/IMyd3zOfGYHhS9UFIa2Kdwu/7syA8g4V6fJt8heYLKkWyHEv
q89LMZAijUikcgFfhPG2xSp/YbEp/p0SifInj/3bwszxPMf9Gi3dXOzTbs64srBu
sn1pLeBi5zqO3Abu1sRtVAeunyCBknZcHQAj8HkUJ43ZKO7j+Um4wv4oOMUlodz9
y6xa5THXEkLXypvHv94/+LmAffSForg9CCH7WzxoDuAmPVzjKV0sxt7n7LrJH0/d
VMm0AfDwSbprpJ+tqqVuOwt//4hRQ/fUwJtPoMJW2or8+Pd/nxYFoIOlpu8+Asj9
hao11HMoRk5s6UQD/MFSG/s447sUFGKpa7IR1ItPliGenbACAn13Ut+e5Dhhj/iz
GAP77N5C9zF1TsNrbJUHCNlvvF5bigutmZyT6pCT7MmghFwbIikfPiJER+XSPu+G
UnUo0IsNgl+uLEgsuLHGsxi2xEURvtymT54bevvrFkkjXMpC9Z5luifAkXmccsXK
JgXoEnBB8hmNl4FD4koE9CNOLgesloyDnNCeYY2Dyl0xJWWsam1PfGSMqDvrYQ1Y
LhmvHkOzHWPpKFXMhkHzBGwo/YnmBkVniSjr1QHjA2ozbmEGoo8wh1wZsS2LwrYc
udTmVonD9eSA45MOwq7iaKIYYtbg7eZM0TXIo7DT4BMzMf5p2ICbaOK5ny7z5urU
P2vbhXuUktrVLWajBaifuldGA7LYaUnYLH88rl7zbbFLbiRQviu5D95V5sbnm4zV
Cz1Tsu8yA6AcnZ/PaTYrnK2sqkkpNIawQmemj8m0T4uscGAwGUvpdoaqJiVwM7k7
TWIxHNOjcp+r0hO4h2624jaanXUJq8UosL32XMKBHxbZMLNDJpcG0dTl408A3ThT
2asmLo3DT8R6zTDkqCnmpM3zKmfFBViYv+oVxbP4nkNrtBT145K0at6appiJsuUw
Pglo8d/AgJbwclyMKwcnBm98w947pQiTrR+1JQPn/1xCZ2ndc5r6dTwGDb6OQQUk
7h23Z+Pe676H5wjLkezIegFgk4DlZ2Tnxj3lIlhBVPx18Qzx/glYh7bYarGedavT
DGEVh/WhwMaB9zhNiOmHMghjHPr8mqrBDa+oa1Py1FjP+oWurjaP6Kdq7wL3HX/I
vHtv9IcmELB33LAC/14wywXihiFeXxnJQHpOQ9+xqd6F7uhT0O5rqBytVN/e1mHD
+kHkawwJ49MFAPBYy6RDrLR0qDrtDDCYDG9xUvYIyo+doT5uDvmVDEe7dQHA1p87
9WWso36K8HjImz3aFHd5U7nJGY2CfSo8NUhNsO2HLpYEO7eKMZPLC4edc7ZkBE92
06CtS4EqZdktWz6soW+G1FRvqtFfaex2zQ8n1S/zl/7w5onOqxO82JVmfHiZ0xaO
XKnkrESbQtXdjwOci163K9rVsffSQs9n7rqDk7Gle6urT5dqSHX+cQDNy3Zi0Dtu
OybWkEtfBAZ2mlM6rIcCqhUN3OuxDyQgEtk1YltFKKC115qAZv3MKx4Dmyd/tzuU
XSJm4pp2C8XS0wwQEP6Uej9lgcxOrlL39y9A4EpLNHriGwJ2k1p1mX6mwoyO0JJq
SFcHy0wTbDNq0o7ChpBhNAKbAmX1c2U30xH1ipVJ64nolNYEf79tHBrpbfteZwDW
aHzn3jAdhrt4ndjds/tucw34drLrnsaNKeCrK8+og2hEPEjV2hGDHSwQ5AxzIzFG
dJ+XX9TOe61FUA5dyqltycROesC8I19isvjmtlA0CR6bMyv6Fa4zf02EwRBBqCOQ
Y4LCc0CvxSpkdJjCoZGzP51LqhdcKrgn59lGIPMxFoGmb98JgIQJg2v2FSVUcfuH
9UwyLyZdZAJyuzS685+J7vtofIWMaNvZyGCrNzpY6fJx5EeI6tzZnLubLOmmLGts
cNfIVddXG5rADMGHFnHxNzY3pPwJT5yVzgS2UfEp0AmgyunRqEPivax7y7lUztbp
DMEl3piqDv02ar/s848oWoLJhTzsv4b89SYeQ3kM+fVQiMyaFit2K7YmhFyVk2/v
tiMeOTuEuPQMc26tblMpiDXPS2+Rq0UBb84tQM3RM2fKgcJLPdPENA3SCQ4IvCqj
73mZ5YI+st7pK+arYgdanIMu/W2p065EcWlQwC8hEGO2A5cgVeCxDNlREb9R5Wqn
+qjHqXhtzmlrwWZa3hUQO25QUOTwOaGncan5+kQg7PW5dPSIX2UFRUIS+GPlL2x0
UWrspFWM+ciHl63VbXtasSNofmPlM4K6+DUaqlemVpbRYl13VPKbYnx3fgzB5JRv
uQlOD3J6WWV+CItd1y2GPjxQ7SLNtt1gbPAYXn2kOIUkDMSEm1MFEN5RALgGbQQ9
teT27YoEXEwmXV8O+Bk+kgkAUD+aqIQOFs+N+z40hABYuTD1lTN43ykauWfAidBb
U3lJko5dKc37NKe1dTbLY4qe1l1DmMnJdB7oA3lAYeygHKyY+ymnSgHA/ZyrYEGp
LXj7ZJsMUeI0l1SSPDScOFKsONP6MKtJDKWNEHPJy5Kcof0Qebldy4u8Mafodix8
v7PVfafpocQJzkK/Yhukldrq6EiZtSpZz9/u/jh3lVyQRF6DhyH0XPNtMY/z12cZ
1irmwr1l2+rcobgebQnOAyQI7kpB40fz7frLOGrMMwF0W25uX9aKkcPfc2XwOsx9
/MFCvkj9g8JMxVffVPk1SsHM8T7nynjGIqwNjaq+XFtFcSlllTWb9xxe1Fbi8NHj
7ht2bQEz9NylEIXop5GCJFXWWxKy2XXL63XlZdWI1VCCE2TCaxL5MfAQMCJU6WfV
/PaLTCdPauBV2/vB06w+0ItJg2lLeUyRdwzXlP0eHihpJAG9LZv3nt4OdkbEp79E
9qBY5BEyAaGuBoDKFCI4osBUp0TylRgyaQLpkZw+geQhpc/PHRniDxpqqi6jc0eX
pIb/zt7oPWq8rAWmahS13xW02SPsq4yHrDfasJ8hGSpl3ETwUCEv3nw/ny22YKM1
6ckzH/jqjX6osu28rEeKelOBgSuXiYiKLMUHu+MJs3CFmOF6snFf/8Onhet04ekF
mL9xUFDEWaG8hTwyPlZVMsvx7P/vipfuM8HAyhqf+FHz853jErJEtUh5qciTWGMh
emn4jJ9JNf85/GTzpf4a5lNRcJa6wRR1rzfkEX/2Qk10sS8ERVRn/TAp1nGH4JIA
pFK9NdKKKq9b4XH0YNa5t7rTD/2OQvUrxZkX1puH9vB3Y35ImasXJJ0oRaFEjx+i
mvQSJXSMXC2uOwM6+K0sayBvYyh270yyxmuVA/1r1kJdJU4QjcBdvibHTWjtjt/U
KiS+41ntz+cNGxYbyzZY5z8nOMKbBvqawZy5blQF6M8FFdmXGPjTY4troFTrtPtn
rgJqeefom9P77InEuvqd3xlrTTJIKczme9Q9O7KpgvWAZd53zr2juVnCCGVCTd7C
U+2iK4VQZUXOo6LADw1lZTwJZHsBWSB38Ksy6s5f1aCX/1Jqdx9/KF7CWBbzfjWF
mHdpY/CEVjiDFUFgllJSxOIgbdCDvQsPBN0K/tOkTLHZfkm1GXwmq/drK2erGczG
wcVbesdosVLtw9n3WsZoyAsdw7yqKFtDrzszXzul7CzVcZh6Qeu6TSKujmbR8Xwg
amVOjJyddRKQwQI3YhTUubyMarRpVvRjpRNAT+CUR4Xn6fmmfaejn9bAZByuSIhp
zEPKmbKhH6S66axnMG7qfffvr+uf2eJqvG80jo3v5Z/NFOnnXHX+s1MlHgOxGh1p
TCVj7uonHENBN3NRcvomHg9D5FdY79yuq8SBPHgVXufpa1E7Cm8Qmud7kHcFCFaH
O8qEw9GHgM0g7oljAiTBdpr+DlaPl2kLAqgahlf5IRjDThqrSqcNeRsQNfVgU1+u
y0og5pLDNRFr01GQYswLA78UC+ow/rvlvY3ZUc2rYa3fV3igXQrB14fEE3qqEsJF
45kFebDAQOjUteztEMJ6X+yljyQ0Gs1gE5wWS51fw9PwY3MbzaU7inqltELk84SX
vhqiGP64UCBzLt8QkTGCsiM1zhBhRlers/90VgXSll3PoqnO6B9VMxzeTXLx55xT
G2GEvSmu+rYutXLT92UHgbhursTjJGRoEK7Cn7q2ZE09AtW533KpyphZBfriNdBi
qVv7luLYVIziy9agGGaJiX3XzDVSeIqC6O+kTHzkcK1M5qmuLY5ZhIIGLqHnYrCJ
fhQA5uH/HfhLQUwcstc8N+xa0JgsU1fck2AYWSlL4VtltA9QGx1c/Ccix2b/oSLg
5a6SV0cSA0obSqhWtRf0S1pkmXriucJz2mW85WFvRKwd/U1/cWmmtaZigo8avLPO
NvJcFfaq41XX7q0/unimooP1s38SLC4NyTC4W19ku8dOm6lFH2JZy/THR8qA9LPP
oeIwOQwS/mEgdn/RwM+dPjZYPL57nUv1ZNOeycAK0teJxV8XNqSXFYyVwTGE77t6
adfdpR0i6WxGHEGr+cW6u9Utiw6Dg1Rg7wf5U30NrQx3i1Odi3/kq58qfQgkri54
aaIiVwb2SYk+hJTnmOnDGABO3muBoEpF+EUndpU8uj19J1ujWd5PEZDJXNQ8GliV
ZpPjddWMmxHYbsBy0oflPPXw8T7IXkkOUslmHYW6RnlKJQag+/RRbaKoeGivD+TL
yc++cSMdXewYga5Xo4isTik93KQYWp1pe6tTUMogaow5moViBVChGJOnP0LarAXg
8k9ViKksaj1N+ETnRAH618shWHVJbqCD0eX+lfCkWp4HmPnebZdhoNuIkWUBmm+Z
3bdjNPLTGIWdSjHCS7m8GWdHi4iDxh59cAfwHrmgDQlj2Q9BWbDupz/LResGIyM/
VznEOmAGLhcMZzID7RczxXELkRVRW2aeYujq8SimZrMQFmthR4BCiRbzfacOo8pN
4SJwNMExEL4Qe1NygX0or9XW/gHSpPnYYr+VXanFwmaVcdE3dughyQyV58T3l5hB
/5W7lSYcdxifsZfYeajrbp+1lkBAyEaiZG33ffu5tDftCvpG4HxH5t+CR35UMiUS
oD8jmO0j1xHwNsto71RlxgUnJeraawN/nSbjgBNBuuocGH0qaXXZcA3qB6V+H94/
cF+9I/kthV8qit2+G8AwFmhFuOOOjFGt0aj5Df6ACwp3L0IH1PU1/82nBZpMW+1V
RuININqiD24cxADpmb1otQ4AQtE0wRUe7S/WYM1MBAKHBLB2P1SNcijUpBAWePqI
no6eVZ3gOEAH9BEUiNnzzsG5BgdYll1q5rRQiDjBj91twDUnBUOMJz7IQVV3ZUGt
cKwCJ0MsvVNCDMoPtcdcQ22rjAMOrf7k5E88s/CxTWLl0Rb6Oh0rBcLjCr+T1qR+
jsNNSJz+A33Z7p2n63HrIvvnJ81SQlFoF9Q07acorCrvA97HbNPD+GR4vNz2rv4m
pWdwgXjkicpAgog2wxdUr1tCYEJkRUpbbK8wZax+ES8/cQU9sGSi9zksMRkBvMKB
M6TPDAji6LqU+B2p7Wu61IpMkbkX1LKKU9HzGX7e8ZvTLWefO2LlvOZeEIa9NUxZ
fTpui1cQpH8e/xh6Nl4XTeeTOBNUnBhky8ogKkujAc5q994zh+SyP6+NCvU/GbmG
mPAW/c2fbmDYjNVvqkyi2zr5WyJZ/UrXwFthGp23x/v1DzlJNAXQwYCD5YY5aJbT
IAQPLHIGLk3hImJ9Vf5O5HDRHdkG+jx7YXezLIP1CI3FVR5wJJU5ZDliFSLLCs+N
U8BMW7NmDAkChpzsSFopHY/lcw9LYBufJA9/K6U422OGaHs3k71MK1nUDBxCdQbd
gFG6U+tmGSQXTdepEA4wQnoO4mUyPfH3+OvFWIoT292fili6YljVavwN12ere1N2
UkVESlrhIIJCRLLHlldN/DnC5XFtKIx4PSMGfTWmUj1+ANvEG0tMilif/la8SeDu
vjsWxjN0/5gosNdi7T52GNjTAGghGeuJ8VsRokfjFdYMBkMo2AEDDnq0AkShHVER
P74HCvtRvF4cuQAIGSLDaDLCEXvP/66uRLPpDQtij2hTvoOtxPliI2tx3bk9pXOL
z3kDhayzX3tGt0JmnfwwZiRFtXo/NLzf15UwGFMrIV4OVo7tHEkNYAg/RxySyVsW
tG8dqwr/0yiU3/fCUPIApBVuZjs097DJ5Ea5HAxAIye77V5/oRUIbBHCx5ZV68nA
rjghozklt3ZGwLmV6uBfDpx9AXmZG3CZAK5jlDyqidiwemuRKjmFnGdJOBoaBuB+
wUCw9DlhTkZPf8F50kVT/fgl6BP6GHyRzUy7hA+wcsTXp9k5vS+hcM4HwB03PBwU
PViHA4vZWUR9P2WzK9Kc616sAX5BIEA2J4jOrLf6tW4ZoTPyZL4uuSzp0+eJEBBG
vaeNsORiP5+2aCwKACWUV8hH6LHiF+ImpnRI+oB0Xp0pAPbNgs8kofBgVpwJxdQP
poSlCfhZKARvyJQVEMceNuGow62a0IcvRbs5N0XouymntYAOBVz7T+dgQanZncka
mhhzsEMWEGlodU8g6egoPXUrlCAUhR9zmV5yWX9jo7LpK/8TMeYs/tGirT4NzHRi
CxWuWWeiysIasxJcwEcB85hJJ7IbfFnK4hHRyETwL/vbu/tcxGZc24KGFcmOKq2I
SqSxAlxZIudPZROHf/GQ5VYz7kpKGd72BAg+M43EIbWdTefr4EJHI2P/Qg5s3BXx
iFs3uoP5isK+V8HdsDeY4Jkg5fbNfNFqyDINGq2e26mfUkYdwWA+Gdp4S5o8kyxB
MUO3Xa40XKSVbCXjBTQZEsWaECZQB8awsPD9nklGBZhFP6QWtYVEF+j40AtrDdnz
Enz0lWWzkwESXjVPibpQKWm8HoPd/epx6NfO6NPSE34RV56F50AU1XGYyKAGhLsz
beJCTr/5kWfoD8oLyrvP2noBc6RlAiZDYLjtjTEgYeJtT+2mmV2yVGJFxojEIps5
4lVkwwLblElnS8zLaRqf3TR0A7zJ2XlodSDFMLHBM1Hx4L9N3n3FUKnDMNq/6jPm
Ncr9IPG79JOMvB+XSzjoV9wzZUmxPv30MD+K4oPVZtI5LlY+FY8beTfRD2DrIhuh
80n1IMhnJVMKvYYjFDRAh8877GIrM3022lGpND+tTogmwd0/h8pmlEj5p7WYgg9v
p7bMMBClXCnVa5jdtLFjXyZAA9VygI2ebF2rEiM1l3B9QlW/EpDCnWRh1u8cW/EV
1Vz6ovySrmVBzHaf8M9IL5BFO2cBL1MgL4+q+nI5dt9KPWtcwKSlA0XvjB/0qnYf
+RI3qtihRjxV8Tl6yo7tfX75/NZD+x9Aphvtiu0tCGfl4wdrPY7OkXsHo4Yoz+o3
Yf90AxOpaT87x2Hofuqi6kAcdVJkX9VWJBjKzPraJEeoUEbBx7VrEZPSxZbmF8Ht
QxeLKfpMLggKy2MwkLeva445FCxXB2gBWGXUWEn/tDlKzPxIRGEIPeRzkDKoVJgc
7mO9+EoF4z8nfrCZea3BmwPWxyWrRyJPV45z2djXhWTSPH974Kc0DARjmjDYxseX
16ACRcUkjEdMngTtz5VGj8qGluBh3I0NR1TAaagL8sMBT9TShrJzX5HKlHZpulfk
u0W6czjbZb5tF25RLIInIoeNpytZ8udCNhi7soMa2XDr6zR9IxJH7j4AzKUt/UjS
37sYipXZoz3A9uHzxPtcI8BimSceadKNRCl0zBt8j8ukGBRwhzRcPGE5IK5/xukY
NbyMD8Ac9SuuZYNKkUNh6Jo6/RsI1Xu/K0AUiqW6pqpQwuOtqRXKtRfV7yMq7qY8
T1r9jLjXw+zsrtNgy2tDdJGyl6K8D8ZEPtm2fVTnEjTiIwbVCwetItfVjyU3PwWL
PdfBYP7rNkPY/ATXLs8hJt/kW9x+CxmRwTBg0F6Kr+KkXKbG1frvbQcq+9WZvUre
YfxIu+5EVgqr/ngyoULa7FTjV3SeVpSqWT0Z4YgYPoueoelxLmQqYTNztVF/nqgQ
bJ9wAVnNFcQf3SKBKfCI1BlTGwJWAUoE6Eg0sRJJDfcp0mnpmhCio2y5EhvnJvqB
JGaSCTe9yyaHcnXiFMzfn+up5OnTzDgx43PtVVT5E0MXEhZWKVcCosU2XjPdEKFw
K5tM3WMgQ9chlKZltOFQOmTes1TPtf41JRBm7Z3HRFPofN5oUX8vLFKe5bcH4yMa
LQyV1hsm2uGhhykrpyE1wDojpP5GB2+tECGmxDfJWg61msnWq9jiEY1ELF5ZJyyz
CWTfs91eNy3vkDv1UAV1tv77H3ixopypr/9Hrd3Q9qWTRIA7wXgnzOGI1jA/qG/n
nZqYTV/N3Fx23oCRYChnXW9mjUK97nwANBf2tROqNBnN9YFP7l1chI8iJUNNMCp4
/FROhdKomQg4fooV6Gs1FtUlhIjxpSIoEWYnYfCWF6I90FbV5WpEd0/snaeDY931
Eju4oc+lzaDUTp+6Ma//AeEFHZF/okLr5u9+tZt6mJa5wT5Bz/Qr6zCKy/71BTfb
A81hrdhzVOSZILHzHdA6VTK/8qAzlSGumKwJy40GFnFRXPKgc0CZAguzMIGFraki
cB08XB+UZrEU9+V3r9/GdMy42H6XfMAQkyUquGNvVEzg6lUTftHhwEFjUR9qny+T
NICa2DbAhGfTtstYMPi+ss4uWsp9Q0MVWCbeDBrKQ0LGgCLT01nDFDIyY8MM+eAp
3/ojjWw+rV79Y2iKQIouaKTLdmbpXI/SiKi76rgR3GjcnDaP8lTorck2jkwTTE3R
owpO9EqOM50Bypzz3uG5gemtSTsSlTORv4ZdNEcCk4HeHe8nXoi90mnEVW4FF42X
QhthonfkCBsYb885BpqrZzLg3qR/41ZEHI+Hvwb09WLtARiLZ45SqRVIXwokoVQH
TZ+nB+aCC1jP11cb+QdYDM7zNx2nUTgcyJ8BGcjB1bk87Vfj7qHt7eSj/5mYB0sf
b5YLa9qr05y0qj+U0zgIkp+j+voBmEjBo4V+eqwi9+Ix50vLieZDrQ3p+e/L4NH5
oiF8XOAjwigSr4x0GQ3Gzqtvm1lz8jgZZ4AXfx+h9hXDZ6kkwTUZKSlktE53sfGP
Hxb4v6Zj2peGpbkT1JD2U7vw9q9urknmAkuTj2pY9p8JdsbLMMgjp5djnaIibUuH
m35kOM8eh83c6BAMG2NchrvqMji737Be76IbjTj7wUs1RbEeKgkacRLiF1R56H0h
lxOmwgaIm/pmBpW/J/hz7bAOXVzCJgzxbolXHPwKhRG/FpL/VIu0sqrKPQVC8efb
0gO1UaTT+K2zlKJ6a8Sn2TX9loBAWR9+U2F5oluQp+URCet+Ud38g6FzeQWO37Mb
sko625WaV46sLu+DEJ7KRRjg9Q6PhvHukqxqzkunLN4uE42O8OHMnuesedvXsbZj
XJQyCdq4MimQrSKtsWyoEcPlpE7zQ5LsmrKiNrRAQ9OmNE0s/tPNTWQWXAuGWZK9
kMthu3UCt6iVq2QiYIWT3LEy2lNZu1C7+Kzq0hwceRzvPLO1PGJgFVM1bjR4K/da
FZoYoBtm5svdX88VqRTIMXYO+l86sQwjzmpAq1ixRUD10JlsdSQSMAth0ygXpRyV
uP+juk04IVWL1cEOdrt2+V1BcYqdeDAMTPkpoDh8VYxv3LLSoh16kZuzZ33p2czA
Y32pZy6hic0YPjKsVz/z7htsPTWCytZMcGdVz48O5OrlBK1m8zK2r6eNfeoSnN09
X/W4SUwONUOEjIzYgYFjdYePj0iIreTSGZYzCn/kp9WGLNDgRGGhoT+tkzc9acvR
ky3EWxmtAXRJgBgRGWmHjZpVGhpTsaUvP8mC02rVEqhgEt0F2knlbVhwbdNE8poi
nPrJykRyQupMpcu2HSQ8t2H2oloqSsYKgAT9CTCrcJcwvkUaX8zRVRHxCeoWaWwB
dPSkqkh+eSmg/6NpEkjjPkhI61a5r+xuyV+Eaul2zzR+5b+wodOixJDQQDdXLkv4
jUh8ivq7lJ0tFmiumtRIuqFzOMHGPFZBjTOlb9elhKHzWTFFf2Ia0tnXJuLs5PWE
CnWWnEOdOcuujtTBV0E3/ZIIC91sMRMsLcH/XqLYdXBD4e6Wer5CErXONiD34rHU
nZRDkqfxUuwYivCKn8OuqPfUnVm/v+MYHr96amZRo2XvqmFTCyV17DcYcOYNNjSN
rYQiv/WdYJTLV7r/ZBJ/7rRlFaXvu0wB9scE/+9wpz1ze3h5sAANEkZI+4Yytj3L
j9w6r67j2GcDMRGgYYVukEAdxPKlAMhM9bzJx+VgA4muGb6DKm3rnLCWSkTTzmeE
68/EIAJyRn5fELnT+sCaxXZLdjyJWI5oiOWMRheBchNh4jM94bxdzv76s/7HV3kM
jD9kVLPjBK1DON3mHjQAkIitJtxKfWEy6QvKAY0mGuN/04bsn3Wpv/ydJpgJXk8l
DjC3LCS4bRHoIdi5VIWGKgCLgNJfTACPLLGIGenXFqca0Q/RtjZcFYa7bzqhxIxL
zHSHf75xVuifp3o3krfwylz/KIHXyc64RDQDvgSicAqZkac/rzL4ChqYwUMXA+JI
9Bg+d89dF9dndj3b8/sbVVrGUUvUJkQLXfigwN89qeMaCbpQenr4BhkmeA1r97pU
vrGIMU8wenKx68+6TMG5PsX20lKyLhjc1r4jBLsf7QUd81zBIhIeSOGk5gCQ2iOx
LiAy1uVixOAIO9jgU2S7CdTbD+6R/usIfm+LEk9Yx5HLNvbaEJc1qBwF3xRxL6pg
kRzTmwd9xA+it19xx9pCXAeM5hm2YOZwB4YVG5h/NWi2q7NWjWmbYIR+llH/6oIS
a/HByc7MH2xWSnIlHODMbzRiWADjEM9KBFf6y9hyibc0o8su+eq/nuRfFFOU6bMX
a03ZJvgiOhP7zFAlJFH2GujYBeAJPPUdUGk9DrkK1DtKb80JZ/GmspbMcosIEuwB
J/R1V6HpyrpONJRHf5Xs7evr3CZIjbC5Bf0whBxP9tyZ/s+M9f/pBdcTzk0cneE7
FscsqXx5rk9kSh7PVYNdMaxjuAFTMbrSYkgDuCIkLpTqbHONNnzA0QEk0OUGH7Gt
SeV3GHBpUxFHInlEnAr8pVvrMWoEo6saJ5OLRUKSveZTsAgFrDegJfzlhuz9EgRA
R37pL0zcgSW3248m7czN4pgMf9a/ML2dIBSvW3E2JPXn/m9UP7XpGVeSqCjf40kO
EYqQ3xVSu0/BKiZqYScZHY/Ypn3kpTk6qOfx66apJas7W84EEB7mQNmd6KlSOTDn
Uo4AM9fraH4t5JrJLf6Um8Opz1Ch/tN6NGaTufeAVf6VuMlLtLXANk/UmloDdpBl
HBkl7UV/zQ544xVad9PLEBuFIMZkLr6b35h3SUdkyYAwKZ7jZlGJ5VKrG657DWQS
y4P1SXEGIkPnSQMvYrjm1/gbhkuEnemwjqHUMnSY3HF6nPGzPLDTN7jn9+ALE1fN
e7EdsQ1o4UQXnH68d/plVST6wq7uHbNYVjosxKgMvx/3wdUE01eLvXyp+owu5HLk
3u0Pzqq8OZFrFtiE1ri3FI5DW0hTEZmr1pr2ln0wJYqAuk0++bhv4FctWk7Ur+7T
HAGaq9nV633NTV08jmgEd9ut+sUqotlu6HMfJfM/Lgyhh5gwPH2QZmOo/CA3s6G1
ur4wOygLYFOgXT6WHvsgDIRaKC6cUcF0BLCbUQYAJmUvO8DPhEukSOjrHKmd0Fsl
+iHxTaozQ8QkgoG4Se51Ya83WgDQRlRVtEE7+BnyUghEmIEi0DMrmbeeBiMRn9Ua
HZ+R9giBIphaA6plZw04PpiKu6pAry1ObYK3nWiAt3fXCSFHBQLCv+bIEZyRwI2t
16aGwpz2luLYZVH6rXh+znyQj8+dGit1exmquRdDuK9bw+5XmIWcnIn5TUfCx31m
zLU9SUs9tPYIYvs05NspX3YnBnGhnyFVe1grdQ9PYqJpf0+6a/jbolDvrlLML/yx
FchE3YBX1/ksnCOLoSQhb+Jp+hSJTopWULZKKunm74TT2ikWCPB5T0/0G6yyUuW5
jE32YNB//Dnu9cS+99CCfHozwGEJo+1S3OPLw6HlltLUiDUnVsTKdcm+O+po1Ipj
2SBIMLg3i7oNcRWCdhoyrExtQ89eM7DIUH6mJenlEN5Phf1u+vghlaTXxiJeuqn0
q0hIon3ULN3lvR1+mMUI0zBDIyCxsmHTH9dlfk2N4aGyDSvLatUPep040xJ8+LFx
Ub831o+xzpSaHWvJFjSa80GPqBI11VUjwOJadWehIVyWhpD6fiDezUSDHkmi5U/0
atdkxmw7nQVYWS0wKFMUFHfPUmDWYgHc8UkXLr9AHqfFdmInMvKz32fQBVSzgvfI
Wz8pFwTKu3jCC4cg3X4L2SYoYgcHVtJ9sl2sYKYlEC9L5IE3RhuYK7SumitGLdBG
/GMfJL1Omj0upfmukZauZcdCjdJOwFfnvn3RCkzMWveo7GrvP8W1O40/XVYlPqFM
Oltzy6ikgN7ZgnF//3nYmJgKT+/Mdjz+w1XCKdrnoWS41abCBkuuVgY60uVKub5/
xoK/qqDBfJYGMu6R8Y2E2Ng0ZAVYII9HEKCk5r4UCxBcPNTAFIK4Y5PxWBua1sO5
LxS3f7mnAwVoX2I5mw1PdaB2J0Opcw3s7QkdcEC56NLYAtHh5SUe5Tbs5KIp+qxg
nhnBzhRfOQ0rQWSL1mIgioerBU6bj3Jo65HA40bvhfMT/nO2k6x+qF86FouxYHiz
GBe352unBTU5IQ7K7bWFS59uO9r3ynGAq6jHTHsZKoTQLKf9RBzPMdBW+SSKzuYi
oIGbeQ74ba5zGIBA+P+PEF5GJ3Qxi0XGbdTay0TPIwYB9DNT7cksl1YHk3sdrSxO
7xzj/8fQ5DSCIhtJqhwexU5TCIve1qx28crFhYyE8qz/QeWAyUjZvNkJNkYALK3q
jcYOnjitib3XZF0quFLE+U4KNePxi/eXkrZnXpg0z+WpNsytfRddNWqXQ9Sep40L
TaYixiT6Tm8xQcqNo93DcVVaRSEQLrd47ZdDnzaS6mkswfKrtQ3oqmHjUjdvKJ+M
QrZ4trtuOM4RNALunaOTqR0+Uw9g+L6GIoCMZWOm5nnOJDWKJfdXdOvtmi1JucXr
vPOK+S0F7hZqxoC0/qxWLhNHzuHyVEIetVQDXMouO9xeh5u4+tkdHC7gi1Dvxfac
0l7DcOJPVixC6hfZjiUhbcVaAkgPbZhDzEdzxhq2BdrOomry71z1tfz3N3v3t9+o
av47yu60ARubw7ha9hHAWjtN2tiozP/OPDyBgMC2XwjA1k++oZALx3ROwEsVXZqn
/h0WNURNkaLfCK3as1A4w0mZT3DvyaVmxYqpXYIRekwZ0nZWNstLRyhN3E/CQeAE
QSpwRNJ951R6XDF4jVt61I9Jn7+Mze2Myxas0zaCBdgRXV2daadFjp1kIrlLeYUE
nbgov6ECip5L5r8NUfhny4HQX5T2fCq754Ng/1umCHgJ7t1tI0H4DP2+sI8eIbdu
uRV4Lzz82vh4YTxDrAeW1CYJWUe5uhT+lK+ZD6NsongLHhMGotteDp/T3r3+qZbP
Nk8YaJw1ucxiLPMHXvquRak9ZzVR6NiipiMpJsXgoCV7dMFLuuA1oIt2QmOZ+cyy
HVvLvSPSy21rjN3Of3L6AUdwnd/iHi3tWh6PvuKxoTXx/bcBTL1657Jp+Gi37dTi
p6fqXnhHPY+COI1csBbOhrKUgPOpeNeeryVaaNDUuLyRKLRmckEtBb029QMBjd0a
Vs4vpXv0WPbmwg3bpvUCAxcZgr8sZlnscxRn4IgiOCuZ3kEH7yEtFPyJTRSaZBJE
2njk3PMDjTRNiRJSfPI6e48v5aJ/VvlpgYovz2m7SQuOrjckjwBPFzGp1mST25ja
ifAe2KnCaY3pm9LFEIMHOFA/QGhKLSjy5mIh0f1RaAnIr6sneHJEYv96R1upimsh
DOSv6+zqT67J9ZoRB+6+znJ4SLBK2cvPgmE9uK7n0sEUUp6eLnDsIxe1drGQpzWG
qjGx8pvWj/AUGSq3if1xK77wym2Ehp0TeQRs5ZnvQ0eCt1bUfWAxXnGpeGXVKxKX
y4xpe5efgikKIO/ntgGikWbPgAj+McdQgF7b3B6QaSvtgS0/NDG4+psgrWWwtF41
yl5b+8eF/Yks5oAnWcIn9GVCfYut32IN7N1MjLf0SPHyy9AFcS0axX1WLu+VY5XQ
ihRHNhFQEyIoedxwgPwS733mbomwww5eo2YPev3eUIlPTHMXFp8uIM+KQx84FDaB
2fDLF92vlZ7AaUeXEVvzRgWTPy6W7d7tYd1VLc+orB+CxhxhGmOZktGH5l6hel/4
fQkKEBo7kor0YcWMqWEdzdREmC4dgrmsarRWgVohcZhZOvez9TEUzqeLeRLUSGuy
RpFCCCUc87F955qfu2g92kMPF7/1hoh/JMSnijd3HX5Nx8GF6PGQsVrpj9b2/c+Q
VYb0TOvn3iJWpLl+bpQjhPYA9nsHjaZEXeEHtCOeLHe72eEU/0V5h3+x/vlqut4L
fLVogvQGXF4X0e7MhrIoWcVylB1iRbYGSB5YQDbcgOEd4raOyr9phXdJTWk5Jcff
JcRZ9Ryaue5jfnY+eYH040mJd38vVJle0Y3IEqJgBXPqMfZsygAG4Yxdb7SvqdFF
NZOcbVvxAVi1yPY1o+rapBmiwFA/rznghyA1HsbItKWjANLSt2WTxG7YP0wUORrN
504ANTrcnriDsjXdwQz6PDxMSVAocH9RmlD3/PW4Khtq3G3W834/l4KN9pcvyQWf
pWUV3Bh0bmFb6ZYft0HF47C8yPb+ZHL6YboAcY8EAxKSJCGpApYsEjCfSUsnpd9+
ccXOkHmPNuLK2BUOf3I4z6o9YsDVVutPwUu5+ho4i9IVhiTjXbRc5ol2qbFjw/ys
3YcvhExeXRXrl5d13msPEpeHIdk932UfIne0XaMJmHE9XK7+YNTbhhq0HHzQ9VCv
Dlq4oTG5Z4jDpK7hnS3TcLB6JJzVWcfm7+R0y3uX8NU3Pubz0/1375w6qHQNWTII
uxNKXfnSSna/4qa9g2z0Smo2+MjcmOeBJehCqWVkHOnnZyTtuiH/I7iHOaAJA/4a
ucRsbMeM46cnhe2jXuQnPSd/DIvzNbnW27u/xNrrEBADHXEA/0CkwtSo8H0QgGFC
bvgiKdWZVgY/dDt93f8JWm3+qbsZGS9gyaDmunRXzNqF95T2TC1aBDXPVU9YE5T8
SokVUOfwDv5yw/zUp+larfeQxRl7xb+0haJrYduCalmL8Cpz2MFGihTGnDu60eEI
y1JQ74Z0WpRUQ+/5KraHBiPyK0H8bYrD3NiLr3+m4S5ZH5Bmah7yo9owYOQMUEI8
P7iFrQ3GS+WrN+QljBMTIImYIG0dsIky6asZ5E7z6uIbyEZpzH6Y17mIUREP0IRi
b2N8lgNquGhUb1j1j46ageuQF8MlYUuIj/uB1KyIMeEtfq4awGfDs7KLp5QlDPvt
sY36fWNBvMgvD4Vts3VmHyUUU7SSqdb9hBIsrk7fHwn3adyGQqhQ+RixuNDjoJlq
lLVWElygeVX1mFnkuea7/NtsEYA9woxG52i6QygTQ9Lel8SkcCDyyHCgH3aabxgW
TVkqDWsEKz42gFI8NKcuZPkp7jGjHp1Z4Fv11wg2auE/BNQaGTTZAXzzvpMePlNB
LZk4zNj2vtPa/x3OfiUj5HfMndCsqz/5AQlIHUOHpuUNyd3qn7DImsRuYyrEeSlL
fR7GJRG2cwhKbPhQjaeCEtMFMXFuijoo8ky7LqXXj6lObJUqI2p1yZl1dzQRLmhp
8ZJ65FpsHVgCwEeCVSwvZDA77zS7ut/ExV9NmM3I76tkhvYd/FeXRcXah9df2Jrb
wa0T1R0DzWzUodjZYKfZ9rT7Fqk6oP8XfAnxakVk4gzpkJBazBpoIx2cAmk4nbQi
r6qwXbqtWOCE0XxM75qSWTlmOA7A4SM6tIDnk0wyBarGHMlQmfrfuBOeLTDjvBKv
0n95sIp+x5isa73gc7/K4cj3T/ArYfWIFkkhcUnMUawe7DqbvRP/bfuUt+VX6tly
ILy+WuJ7rMvRhtDZj5FfPorydbY7Y6Ne7lE+Dwxf1imQrVTs3Vm5RVNhPSJzfmxN
5UkwpWvSgS8q3/l4kSfDe/PC/ihL1eGrgzIkeNsyug9e5beGxquNqNx2Ppu3lVRt
3bf7qdoznrwpqd+QiK6DBtBIoVoj/KBofUr5cYy7gcP9xCdi6YCKES8kJpWs+ai9
TowJKQf8wwu1oPeAd/RDwH6ue/sc5k/AEWkEvkKV7AwWJE9FE8KOP9jh8zL0Y3S3
M22iA5bgwyxewKJlmcd+7iLNHgVvDv4pUtWIoCY5E/31XBrpLiqVP4NJkBq1zYAG
9PgugJ84eOCmYDeULIUzmDhPPeBJiA5rdBagK430htptKUCdD/jALN9jQnzZCb05
VsyTzXdeJHn/Wz1ap85a4hAHzjLwHNGruU8Tk9NXUI0ENlAiIqmJNKiXe9xoJ4ee
EDeeBrWGvFnNixHDpxbS364qj4MvyVhQDMsdbnaawmrFQIQzMwF2zlYC/cHznI8U
0TGDB9XsEe5T5jxDznqgYXf91Fb7uY1BaweHjwMJ7VS2qrOI4EpAAcTSjGjDjGtJ
7wKoAPsTBEuw2JlGQjrXjrlsG5SMWnZEl3cK2fvkDnlxrmg1yzvpGH1LTtqd8e/u
r+C7tET2UUlg3nij6D1iUPkIrzzdAH4uVlpcOaG8YdEW/kOl6ZmlilGmK+9QNMcr
HLw7V8loRRUYquoz/ANyz2uNE1vhj+Kd+V3LKFyVfXnn33HG2oc9PFk4VjxaF/fZ
WvylM5o9zEihVk2tXCs3jQZW74rBkKZveA1wGwOCE1/DiINhgb0iwf+4TTdNUXHQ
lZ6H3+hDi6JGZxsTw97JoC1DxXzWGI0RdVbEXnGTe34NAtyA9aThKXqWpdg6l4Wr
yBj8gYlUOz4ua7k+BGE74BCIF2DNgNtYsgcW4nC6dGJ2FGc2QPo16MJb8h1/dE1o
LVC4iSVGjzgL+IaWcMuv8L90omX+XTU0BJZBXk37MSr2cO5GW/aw2/EXgF6h+aII
VGNouBXi+2VezgsbDY+HNa65KVVB6WdBOGSlRLSwxojQORtishe+yxGxUDZApZXf
U8/EeSp8Bbkfu71tY+I1OlwvUmm4XPi24cfmnnLauoylxjiUssKhTKTDack1ZjkC
+wzaKDOPt6NmaxzOK7XUukTo7ggqF9IPSk95dG/cQPJTWpkewyxCIht3qSaqrfy4
3kvExXWctgVdGeVgrpchj2IMTecpvto47DuFGyTMtpDWgI2l5laSlrMEC1NM9Cg1
rqM1W/oZs/1grpPFUFhmuT0VZl5GezVUM+FzyTlB7Ln2sw4hht5V3KEN/6o4qerB
I37gxT9iFySmvyrSADJhdyG7tU3eeaHliNQXovinID50Tl6cfoZWtVof87Ke0Acw
/vNqzeZsq9NKlQHqQZ3ka9sQmx2GQA/SuS/Ejv4N3FcGKPIq7F2RJ5skMKAM1mmD
XKv1QP6yxYol+ehITUiLDlb8JS0p9R3ljvDaDY2Et1W5pWY+o5KtrWIG233HESfd
8va7S7yoqx3qI8ZQYy2zig3+Xbp8EOqzpQ9BSnEqjDpRt5m/zyRontu15yMcS6cQ
n9QJ+1aZ3Obrna3apVVW8sG/V+IHrsUJuwweWZn5mHwfI6ugSfiZYyVSWLsKDd39
gCJ7N3/4OzqL9XWSGoDhkA7HJEeA6acBpb0uJbCfpKoYHQ45DX+rVMUKIJEElKMC
QTt+Z51lOF68FfEPuh/bdvbsyupdaiUHM6HG66RKlKqTiwy2ANOMPFlJmnKtY8iQ
xKexO16u0pYzsC2B/BWrFCSk/rxwbulzyHbO3YX7zA4x+tIkAYgNjRHzf6ijI3ul
hMb971GOXIuHO2LeONV4HWShabeUgTY07cpUN3GCCsI0S3XXZ5er5wLaIlPm8yiQ
mz/cdB3m6uYuw+tfANUzhftzLxZ0u/NnJp+2dKGrjaKgEce1eMXGGrvWwh8X8rXh
xdjc4+fszf0JFi5DXMWH7yilF/kdaPyM3c7WN616GzdiG+GKs20DqRZKBUsUvEa1
nOVRezr+iiNMgX8T7ZkhogYwICw8fEuTvtXHiDihAubwJohI4lKeKNdTvAuhmjcm
NGKyUSwnv6u+kd39z86FjZeLKnKcE7r7hwXYXcSaeW6rKfjoQpwxW1hy0qcSaFgJ
LVN8Vj5PxvI+NVEjmjIFradIR3AGMjv85BVTi6BLy9Dv0sYADlvcIFweUi+pajqh
6Zj6X9HusUOwWYZaF2B8xf2izX8wg5y66Avf99JzGLguEBVjtmlZcMh8M3rfnodN
VkCO8i1sj3yTzsegDF2PVy7Ps8uXA5u97y2XWKTEqjiqzvpuJjKiFyrlHmT5Sm/Z
uywjbWwFCFx5ZQBVoaYSLWNtYHw4obUhCBHQEsiqliWktQvq0Xe+jYwjAba7KCcU
STbWRhbbto0sPq4OQj9bzEBbrOOiR+pmnvjQXve4HunPPmnowsbCFhP619xE/WK9
dIdTVP7JnMd94eeh3Vsp499JYBAAiZH2c6fwmgFpxjdEW7vW3mzwC47EM/BeIXV+
zrD3HWn0zIUmEbOELN+Ept2jzTKtUShDyqaYL1M/LSpkU9MFx7S+Ve+PIlGsW2se
NlKma995H+oOyRfV76ZFPRKq5J4zsuTBbPk5VTNSka0qCh6jEHiBP0CS8qiiUkBX
ChIIxThbMXaBhcT+xX3L/N7T9j4n63z6xVtKPsdEi0j3JABIaJqCELh0M/Qr/Fdy
UhteD3ACPeAGrgKaSqEIOkkGxAKcvv1NW4XzV96R3T8YPhucMBgJjPpiRXn/zxUS
hBOzvkqwuPq+ruC39zSmGI6GAZpwAZUo230AWFdcTRO5Gqs7O2OGcjSUN8NpAtr0
Pby0QDtoer5H+mVnQDnA/cAlK9StV8iphvM302fH800yWrfb28qoy5mMEzprjCuN
4jTpwoBRLQ6SkBcl4ei8+fcsM9/Wl2Ixen8cs6+d1i956gwGAofqub1fcNoXASWj
sjUo7O02l5ojAkoe6FYvRKFYH10j4LvtJ/LAyDpjLErYPFbD01tGTDuRFWeY+NQH
E+pH7jvps0xkGSKGPud8xnV75G4VjtcgykPyJGsTBiPnGI+c9jnhNZ5piuWiBZSh
DwPK0c68TRH+lGcdsQabrnfQMRlHFhh/O7pZUpuMcL08oHUDu8M4hzBF6vuADFkr
4EeMwdFqVixyJFNtyXyjA+WZnCMcfekTK31qF/OAFmzrKAbSpIVgDIbPWfF2/2VZ
DIN5l50S9h9ImJNpnDVxvhP+6XJRK4UM+mB6miPqf5QJwQEvSRsCQxlROHBp+wVX
4xdJzLYT7qinWpt8AYQEostjRoiXTa82mEbZ2HLw24qPW0tsCVCGmDSMi1+uY+1V
IwYurXmO6SyxBHtNMpTnP91ItCNHuCxKsTXeG5enAPRR1O0AzETPU6xwYG9eFxcx
vFIzxztav4TQ8PwSR5HKkAabTZsEUfksq0/kAUMEtDTsT6946qkaPAT/SuMMrGC8
dyxO6kziTHirN7oh3kBNbv3xOcqulscoqJXIn1O6apDpwMeAYoKNxL6DFvQfi7ta
Y0h+y5pB4U6jUDKsBrd+s0VMrnRNMkLEqXgCrREAWGxRGJUVZIGjHBAkHEVsLJvn
2dVWlsWYTW4KWJZ+gRzHL2vCBSlQLRAxa4rqGAYtpa+Njpxu75osJDVBbR6EifKN
fphppdV8XbsBbAdYM2TAioUNXRnpH6q0VHgtIux4iMzwro94I3UIpc4mqlBgCOao
LojHgrH/H9zp6RnpfQ4X7ZRGeHuT7poEQTn9bGx/hsJM428txNu+rVs0MWQ+F8Om
My/6tMNuH93KGbb+PvnFd63pYCAOu+QHmBwzuypxUasECT1rNHc+I2saQwR+W/lO
GRrHUG+Q/jYRDDx2a1fw8hUugLW8hhM3bYebjHR3j/Ru3VImWBd4B+qMJmnwrIVw
48LITC9Bwv8viEmbcMLrWJ+YtGNaJ4LfCAh9wnqX2Fd7IuU0U+e1h4pVuEW8uzpc
ypJKeE8TjYDZF4oXwoW9aIfAZKI4QiD9lpCGH4IJ1ynRTAVYqVbgXdne0s/ERoF4
/IOF13HVsGN/OnP7ul61go0BqhxusdwCaJzQ6nTtSj7lCe5vXK0hYJEEtFJoZQEm
bLld1grH6onKzXWZDfVk0xYMSud2vY43K5s1IY00mgqSjeUqK2LRTDqAHzhSHJJk
eGEeS0KfhxyiW591Bo5770/u3qIzAOacB8MmV5K6TaTIj/CsN7JpWzyi/HFmbjjk
+NjGU+IyiVNBGp/WVZWc4lpQI6cQrQDiNJpRYH9uoVBVkLpgrjiTV6eB+0h8v6pi
iRCuxOJHIWcnRlzJVV0ho0FU//KaDrtjwiHGojUkeoeb2mlLdigqtddizgjU1lMy
6K+4rfPN8xL13X+Wtbsk+lgIwXjscB7LQfUqiVlmXBZQ7rwOyvxoJRGAbrMzEyGO
EwmrqXrKEnBmPJ6+/l+7wCteVs86qURblr2ozcJ7M89XYonlI3sB9ULDnMCLbrqQ
u4RmarypUERusOGC3304cKb8gQ8fyLifkRn0nmnZscu+oKwNNviFa7nv7FZMCeGb
on3oo1AzrykCou8MYWyQtTyg2I8DpsXS7J0meflin9ylUYmpwWpm42GU2bu/pTiE
YSORH0+ipYQoaTC5Ul4j36f1g9E4PNoNF/dK1dUi0PFZ/3aiSF7A7aZIgIDkaAcK
jM4ckci02YBAn84Xl8jSE5iuDLJtquUPEQ10qxW3WW+qvMqoKQjU7R/Zx5x9KCGM
w4lDjS5f9YsaZdQJq5CiGpdUTmZ7bQx5zQTqeJviPdvBioNXt+dgkOH++4oKNvFJ
udF2CwDuuyUtVe85EaAeBR0Q6TpVl3lygnHAe9JLRKM31B4kmMKoRsgieqgenXl0
JUV3MFoMGh1WXP6ybQRh1Wi32if1Mx5ISLS08jgQ2Esmf+dsTPvC9EsmIqoiHRf+
9H9wxdu9psyJL0ok6lOZGZsqdxOusw9FH2ybrV4VesZhdTwUobbS7X48BCchP2H4
7Rvpu4nlpTVkZaYAbYA9N0LYZh/7gjKYj6FX6t7RXIrnHhwqUTtdMX5Wp1IRMyTA
R3FwAFhSJ8pn1SCaVpZu6C4oa6MgEFuKLmMOt29bpvmGECaSi0EOTgqRWgUIRbE5
nqHPOUqTZLp1xi969bLaGVlGGy1553WJloQvDbXTWzgLEO16ZRrc4xVeUeApsiIJ
CdQJRsdesID6nI8/lbDML7KA1mtuYJcIFVIRQq0M+vkHpXiPpVxcihw5cBgUeG2e
nkKv8dJi/nVwn/iFg5IrpPypem3i3ZnbkvNlM2JeU1aqnS0cMbHqKn2XeOOgDUbI
rrzcMTDdH/CZTnYszV425mj9S8IN2NH5c7dmIZqZ1+5ooDZ2jxTkPdKJceImlI95
o1P8FWVA63xXj9dIW8zChkju6i7Vejoj+yLuHKibcPirhUO5WrqGIVF9Uos1qIDn
G2pngjoiMp1DiF/g+CseEdR5/H6h0wQ+szykRiHZqh/ZnQPn3m0poTKzsN4sFMZ2
kIOIyRZDViW+V9yNJlzC7s7Q8OQypZCU/hhZN9lLa/HJCuV4tmkpAvy87q8+82u8
8oQtPgal0fr925F+lqn1D5mFh4J85pstJP54GPDKbr6s8guTsAT+iJkPXZSP55IJ
E5UE8tBwDtii+Po8iBWaJLJi8ldTJrPmb9NMqjvXasNc8xqNQcOQPO73FsTWFxVX
7cv33IJ1IyKBp0iYRkwseJ8wXOXicMWajAxqPTOyqNOPAdUC0vwbLVVXRSd/XRzb
vAqkrcniSpOE7dE3F8fm84tD78uot+Xf79xr21CBBfphWD+IIAMC9PUi9WiLwzmz
tP/YlM1WHiGW355G5cp8IcL1wr6r7Mp8LjsCAvXZEVwxashegFaku33UQtm/ascS
6l8eq6PywtdSbKkoJKDUnzKMa+AKnGyeU+GaQIRfQtDoSYKTNM9L/bGHJZR2ZDls
F+qE8swe17NM4C9XXm/PmTM3OUqJl0bkSDDPvPJnHIJs9cIrI8n+v8w9AY3weATw
MEn9bkfVhoaoA0INoVoXTroIyerdXzE4TqiN/FuJgAWuEvKLjCCWHkk0RqU7UiGU
nvOrjB2pFPpY/wcvd/WAfGDzfD04SeBs+NxoJGPodKFCQ5fomDe5agSNuGmgB6H7
qt7Mf39EmgNvsmEbmcKdEARFLMsO+Y90ON0irni+6OQ1ZlGJ5b2T+MQzrfq/dD4P
aNA/a4a67zalSnne67TFs3zgKnPVl3VgpBYiWacnMcgwQE9rwRY18gBQbEwsiKcM
/IHUuDjl6KEE1sxo8PCbnjVrf/d8SVnTQPxpj2PKhKkYQ+8on1aCEepWU7bTpRi0
LQRP99ewtGZXhMmo+jBe1qiQsHZuWZzT25Tt51fINTtqoX2aKzSoN3vUyltNVw3h
wMPlLlrmuqRdLbJblvCyOkZV4RLWm+AwlummXk6v5fcObbAfYoXPep4GOOGeDiWm
cclfvi5bqmH4VGWHXEzV3OkFouyKJTAG3n4b8aHj1UzcQkbgWkw7uNVWYTpTvgUu
z0cvuTtlqQjfqIfSQCRfVERUvlJF/zJVUE541z3EmJlIlVQybSFRv+oSRqZpieSS
cosWRRmS9Vmg41xcTZZ4x6XlcNVxTt50krMzn+VanY2c4FKejJpAYKatnq9M5/Eb
C7PykuLecl3F4z1MynYVYtygTUctaUOlorws31sH8CVp5u8oj8h4WQ156uaHqdYz
MaxtdLZFU3w91lOy5HVcTf4Z/tq3YKBqHxyLXDLBlgyvRBKEZU36zfDco6bQr60v
Mp2502RAh/0bwGluzPEfr3N6ztTbf12tB2KOkxCw0atZPFCHuNcPlIZkuCO/+Lib
KS5xRRGrp9GOF4WV88yLwWANWRk+3cAvssKot40MBQfkcuENZ/EW2x+R6vcASncZ
Ch3oG558DDINfoIdOy/HIKkwqGzRRWA4km+14FVVT8dSP20JkxteozyghYW4PBtm
H6GtxMAeXvTUMc/DN2T7Yiag0Uk01nKg08GwLOI8YhnzmLjrb8AIGCWjuXG1cW2n
rUl+aYjalOYToNXZWLsPzFLsdnOpPp5jFaoroZtdWJKYJOYyP1RZDkoe1RnsFcyT
bjSNbQdClSA5av4jPzz7tdAWNtyvN43iHRrS9tJGMJN0zqUkb0ijhR5IHfr4A7WT
wpdlWRbu/5t0ignY6wLPE9F7ZkiVMK70U2o3caPfsPaRz73skSDLExLfKeD1+Ccj
FhHGM5y6YBETHZ+X+4SM4EY7jDCCexvG8MX1AxFER4lvYtVLx2sfSXv/9zaSy1s6
xXQZOYFwKmh+OWo+XgZkSVQVVB+VMv/p2o3qU0dgX64jfLx/1bn5qB0TTM5daKDX
hrap5MraN0NONvoazcOa5prDwn2rLyJtIqQAaejW2nbBsN9x0QHBxc2Y2Ye4FB1k
ROGGPStexayvVKzOlwVikb28rcppjlgNOa0QW993wg89nzS4scYdt0FhrqrUhUh/
yxd/NhV2h72EM65/q+RvdtCr9WD63nrPvh/9GHoJXsrEuqd460Ni2loBJ8TfvEj0
jRpTqyayORSuJ6xlHwtIPzCybR7WQYQTkDdChfY1qYwjdOGb7hhHrqXzI2GQh/Ze
bNQz8m5dU6kCu5MsLGZLL2nr5rgFtd1yxiOrK/76GKLQtzWPssaTMIsBvSDIWzKa
WaZgXb+Ga1wC9CflRLfFHw6XmWeewGvcMOhbcNbWjD9pYOKLv9OwsbDEMePh8ycp
jfte8rlja0ALR+Yx5OJg+sjcJ/ApicnAkJOSkXxSjgQkndpfJq0oVQCjVf62kdEU
80aw3pDRBfMQleAMqHdu1PNtJuSNRPTlWse7W39lYt0tdgFuIs04zOPaCR/X9iLR
Q1ZK0G3pwe/W/Oo/byPohecNO61XuxajfWwVnp4angCxSdUk7fCyFXYOUFi5AA1b
p9QIwpLZ5CRd/gCMfZsssYpwppIZXLdOi9lxZSVafsb1FRruShG2WccHjZc6AIbg
cGoa2us/7FRgrzKE/zGjzehkoKoLWaCaf+pb0mZXhl7u/xXcvYvdPgbvpPJ6o+/z
MQQKqbIrKZDeGqBwj7QGdBBjK6MffTKwWVJZEgjcipMhPd8ZSjUJgfIRoWQ09lIH
fLJj24RrT1Q3im0fqVsfHG5ds0OYbpM4VjLW5tFV9V2l/h+Z61/I8ZAIkgEQkVWc
Z1fvjEDxPPo9NaorhBSyFnm/4cyZNzLzviph8aToHBZYKkt/D26RRNu5n798gwP4
hNxKHkrXzVJCmR6wW9Y6AljtpisD0KpJPOZLo9ORI9exPdr0i6bFyjxaHUDxV83q
r5OGY5iAnb2JtMHDndX0QdXSiMBwgINHo21xB5z7i3yTT5JszfjdrGupr16VwFWV
qI38c1vOPYPO7kaYtVzQwr0ewcoTGO5cF1VPxB3qTyczpF9n03ANnv2uPMyHeZ49
O1mmLXDEcY/v98cP9PcU3i/zoMqWJz+JU4vtFiPe3IFit5ZENZxDElPM5Z0Lh8De
tDuFczdbpwfVL4/Z93KtrI/Xn6RKr35AcAvd+yZqzN+Enbz1si2/TbsqG56ADA77
3ZwGfvNGoU+BysPRB4Epdzx833QCnc9y82FrSGiBdKGpwBs/uFc2JIhq+0sddmW7
WOhkW21sTOArAO06I+u35hgqnKUzjEtipK3RjTG8VhNSJzaDbw7GlO+IfssYZR5M
Uk1zbLgxREBIRSDDq/CfryFkAFSpuhbTB7PrzjL69+rtkmMuPGLUI+bA34qR0raU
d3ovcnZPGY8w9cJxkkot/Bu00h9h3ndAPXQqeqmpD3Bli/DXDn1RZWiVLX7O0GOX
kVJ9CxmMLvKBCQHC1ReKmDylNYf8i/+olD8iqE2gl2KcYa8/Rga9dLia05BzvbOF
QkBF36nl1Sqnrig9HmzfGgDJyzwfNKFyAlK3ZiAExi4uwcfCPX0eCxGtk8SRoGcb
2EgDAXJ6HJnCFMMlucXRPrDwlpPQv7Pmk25zZAnLxcug36Kf7nC9P4AuXURJ2AzW
RxEdmqCJZ/mTCJuf5CwlJ2+C7cyY0Bxjhbh/FVoOZcbolZl0Nw99KjtsbxmY5A4A
w8ZIv0iQ8152UU2xIQZXp4cUa7P2zFRB08TS5cIgxHiDSV5SevsJVBBFtAvj1RRC
HnOdsgtNVd/TQkb6X4cISRMCcd0UWWmADqFokxdNpy2ZxGVGxYBXWEsuj1TmHIAT
xfOpvSYeWeiC71f4MlrZ9RKnyMprMmigbMWpkH0o1Z7QUedMT1BerYnDm+qV2Ljo
SjXxhrK68inLgMNlfP6U/0to7lMymwGJC9G0sl4KJZH/X3a/GsTdurdEKZ7mIcYR
KyY6x1AypMNCGNTHLuXaQqmEAFQK1BTTVlE2eHBz30sq+5+9LSgKodXrepH8FSny
/JKmkj254huUhNXGTSWmIAu7kVTdUhDE3A/qzMBJ3EPcjhrFhCDMwWbPOs9WjaAK
lvoSNL3xrn5udkW8PAQox85b0xhCd2gy3hVaPL0qocjxO2NTnvr9u1vs1Q991sr+
w04f8czSMJaZcfpWbKEIbzi7i00ZhRURYBMU7poI/g6UaPtybGNtuCFkzNHDzfkc
A5l8mnnGYYJXC+ADmLyhewHC3Kyvsb1XfRyMvLyBjOwxyF+G4ExS4X9QNPvcfBh3
39OdooMBiTOQn3cKgk79IUpRp6AWUe5CK24ghQT+dEK2w8zj62j8z9WVHngAfNxm
Tb/1YzbrJW+8qF4K72D/7+zm5JAzd7tX1ijIHNyASFdz44rAKC+EJs+OnIk/KNQ9
touGk2ZVPODLG7quqAx4/hnqfXWU8yyhsDGFvucqlItH55QRIygGZHgO4xoQaSS0
zFkLEbE4T3Cvh044ECYGUOY5XZNlYI3QR6iQrMq472tMTYXIg+LgHUENQwVewOJd
vGQHwxbENcaNq17SyzhMjU/A0YG5Saq0gWQI47cYMa4KoWl8UWHILZAqkX4eb977
iZoNVGD8njpWqLNitIKEiKlzB4VmZknOGTQQJebVmDi+sChQeDG6qK8u2YEcjJIt
FvBTh4YOW10t6rEZ76jIlju6rlaIl+3KvQF+5YAi3I2e/yaUKaH5650gJ0zKtA7c
t3rdur/+xfYrb3xpN0oFI3Fsupwy9ECTbs8JW3Z27JtVcm4Av6IwBFKAuL1XI9lX
dVUQqMixmY/r//HDBy12ZmZuPlBuPsdGJT69etnZPH7X4LM2OInBsIxkCo4q/mCG
E8DRsLp57a2lVUZtDHV5xPAzrmYRiGpOsPI8N0cLujgz6Ek4ScdC4kknff2HE+rT
jvX6tsEadtcxAtDmscGhlk+8sGSu9eAI7Xss57UDJsqRUZaltrAo8i4c5l6i9j/T
U8Shq2qdZwSF0yDpoNtCLcgtNVGu/sHGSokCjbW6ULZJybz46au8pUmnt9G8H+rF
f2fs21FFtmpBMMXJjv+Y7/oqqsahdCqkhsmmdN40UoZr5EO4ikPnZroual+PqJiD
rw00fzKAyGf75fQW6cz9q/kq05lsTkjCV1kSxIEMaAogpx847LPaucw7Tc2t5F0u
eMJSrjJP1BM4772qqWXOS4vy4fyNzSSJAVcz+n7XkNiEJyJcwIj16ihCfbNFZzkb
IyrHWj0jIu8WEONuLVSKeYh3BdFEM7PMlgPdkyI9XESb1tQ/pYsr4YC4Na2m6hzB
WCqejUOE5iv3xBf1TqT8DI+QuwIAg45zavWl2/xUUeDyc6j00vR1aWdl2OdPhvdM
w8HK7LaeF+1+RsFAhgA+bn70YSWyzCEhnIXUCWY/85Weyp0s1jPizh7bM8ODbhl2
8D64R8LQPocL9tOQl+YV+rM6QL1y8gTwxw02p3FnF6oh1sZEL64jG4tBdHEDQueB
/c5VMwSh3yos3QXqng48pyOjRPs302vCr6juXHFNjnIb+4M7hgMDp8vQt0E5wjXs
Z627GNnjU+64SRucpulgfqvx67DmQQ5WqVKaFuTzhiW/zb5drU71QiL6LCpFpyOe
oDHwP694ZUCCPeLPhaGFZvoSZaGpv7s4QQo/r+4+9cN7MHik6kd3Cebp/be7adZH
6OPv1vu55CMfj5dT3j57xlvRy0+DvP6R2kH4wd+dWVDoymTmXLLV3A/oFAqpr5x+
O1srtN/EaK18cpYWELtLYiRHX/njcZD6RbHIUQKz/QnO8nrmYBVmUzoZYLnUqFhC
Q72tT3k0wLr4pT6o81xwddoVQUwsf+Ot1QeX3BWjUS4fQjrKP0y6RV9/HIFO4XjI
UznXWr9j2AAoFA+9ZpDmg48KmLhsF1D0YmqY17jIuG+xtOVclqPE1lm4lFIexyVd
OcDJgDBVa7e6+TSYntqXN2aliB5HCa32mtGNrE7QhMZ2VBzJAS/ycJQlli+WaC5q
eiOD641MVPXef+vVM/tU3xQuh5m/jkPR4pyIAk/TV5eVrxSYSTKZQL/w2bq/NxF5
Bt/mi+4zc2EpIhhSYMXRo7tolMW1stQ5hHP1yk/TcrIPZKnbO40Xuht7qR/cCYkV
aoNKtSbyakqBt2Ux1mzhhkqBqF/U8nsrv5YelAInjJPohEKK5MmI6oERzmnd5rIS
tyZdSFaVB/8R8OoBpJbLxIR0+ug/wJ+fnEQBngn0LqHzbBr4lH4WJCNoowu2720t
3zfc9M//xaEBiZT/VUZC5/Aaj+xd9n85lxpxxYn9LjfYFmo2vydvI7EeHoR36OAP
x/DGORcYX0DWlA3cKhspv9DfeKs96WwmI5PIhh9hWy3o3eQDVzZtZYxXg0N66Hnr
rXC0P3Rlp2lwj4G9H0aWS/IYtjr2wYEtGCg7hGzwQImbILl7HhOh0PBztlgnE/da
I1Nw3iAJSyH8raPCndDzEj1MeHMapZf/m+mag8DuuVqIdMHzDZrlD7In5zpocZh7
8C/1gxXBloPvQq9E29PebKJOpDB3xdxE7BBH+PDOIEflqXTudCIibuYgTcz9TlyQ
tJo9Ci0zsv0U7q+youFp6FVDtVvs2HmugyGDAfU6ndfTPvPQ5U057JU/HnJhWyk9
QXmFyjl31WLHYup/dv4kEeH+nT9cVTa3N10fvLKiwfi/QFTGd9vrtKnSkiP+Xll9
cEbPr17/uNjOdU5Nh1Y5xfheEYoMcDI22PCqb4a35Kfwxjw9l6uWbvVe/uWCF2FU
P+aIl3PZN183JfLSc74QYJQZC659Q2ti0fUYx++BIy9hs6rtrDxuquopey4RYLnH
KHWFXif1mo8J8+RZSuYU0ra/pUIGYTy+VQbv/HRLnt4qKcy+wdfQCZ7mpNXtLHZk
01bAh4sIFwQS263Lmm6Q/HZKlWjWfNUYHw+OKhnsyXG/wIISPW8xMOqDav9bCPXH
BG97FAqBfmrtUU6VsQtdJ0Yd/T2L+WwSalMOS8bezawfo3kvrgT7tii/KSSQhtWI
lGD+Z3kMFrUGNNLQgDgiTeYlsFhH73xQyxAj6SMZB5KBZ7V87EcFhNf82RCCVly7
FGwSZg1meaLoLViFDfdkpT8rnrJm8eQnNblBXGWS3783RTKqOAO9ayzxxaoD7zq7
bZhT1KjrjMoi3jGdU7AuEBaA72jWksAApCpY2KWeVOqVf7AZoVFVMLY5LiJ2Udfd
Ef2YXXscCaqgonmTNSfrDRoGJtCPP8T98jMn0DLPMbzxpcOdi+XXEt2ImjU+G+I7
c7rsgSoMj3WCfjmVV5UDaTyBZH9wGU029cSsXfNqcaAYPNtEnxOkReQvYa7+4HvZ
kQauvaH2CXFsP7/SYvwDQWq4gOMfJ2zttJc7ofYkDkPxlIC6TiZ7eBNzdzABuhBJ
sV6/oozV259Uw3iW4HPHLot4lC5Q5HC8pOXQPT9IRmQyZacOeGz0BAxjE6VbUE+q
Qh5E+f3YzwisQ+VV/KbgXzlWdEUEsQuh+yYQJ8TmxXYqIdIEOwi6FFyTGotPTjAa
bGZegiVrREuBUvtNPNn6YkpNUNIkU36TRXzHNL9LRT2TCRSUZ4M1H2LJ3Tn5I3b9
EeJmeVeCs2W56UY2sONPEAHBf2Ub1rzrnzJlefCEs5eVKdPn+VjxnMe63y5Hzdom
ClIuH7jIvHiyDH9Uysy8K/O/HdYoFybkWtYdOHMyC918Ks42IfR12JlUQaHeYwIM
/CXYppG9aGLGQWGqEXqMdEyqzhi3tHWj/7POliMcQ+PZErzWqUu/AkNqvryBgW+l
dq2Zwrk6GfajWm8LeD7SDT2zYeddZcoxOF1bLpg+gNChXtBowv+jIXQ9Y0i48SPn
hw+AsL82nBY5/u3HzywlfAEpJ/MX8sMs+VtczzkcW9dC2sMAqWwSLFVici+N8Pm1
lA8GmogYZlTbqrcwXEtFtl19AFDxOU1HEIoVScHepIfaFb7lrg53BTAaXiEIDDfx
59sQfV02yajYJfdoU0N5+jGKPkY5dxa5CiVy0a5z7GNjsJrhiBDSjuPpj5ZwW9hY
7s7v2ASMXvaeIpxkuh5cyl8VflFLVJfH8f//fRQPBNUfQmcGBH0fmPY5Mf1UtXXh
aadd0a284b9B1JN2dCvvnz71+rR4EOtVBVn8PK9mpp+kIXBrQJkqevkwIJyI4Yd2
osZfHUOVO/Hz5bhZZ6DuG7Cmi+xl1r2k1umpzas9pBNk4Tq2/2wy622xXh17GB4x
K0bOBCWojHjhKmz08aV800kySA9BOvdfEQaiZfNJD1xfLE2PjFZDfdSgj1/AUeYg
WBO4m1hnf65IJpD5ZglONYKzFmRoGJPb9i6Qrny9YY3Xt5nCCRZSDgFFIHK60NET
Hb/gus5yFEbbNlwYdpeHtAl4EB0eI9h2qpxngIURg7g8JQr1qQbGTqupoY/fJRjz
1yhexjkZxo6RUYC8Sd/+/yuT7lJXyx7i+k2/6FtEaDPM+Nk4sZb+3AdYHFgjBaKh
KooKypDXNy773qSzO1JnDYwTy9zou6CNXmtB3uCmv1+wCo569E4o15wCMQ137mNh
neP6QhTr+CPNY3exdQKgTZG/Ug41EHBEYjUeQ/TW7bMrZ/l6KPAnZJ/ZlkBbnXxM
aMfxbox/6uUSDP6WiKm0mcLnFKTPDwoTs7+eusDFn8WkE6sOru0R9d9BpSih3zqh
2o+NSW2x8mZIkRrJJklJsMD973yfFcjhADNowqkGJZF2xa7Qd8BNz+djN9fAntIl
uHf9fX3Vs72A//X6oycx/SNeKkdEZzxNj+EZIdYc+wiBKF3VASAKjpMCLLb9LoI3
R6wTgNJQQI0l6O8+/XvSAvCw8F47Vm+jVg7p45zvm1+DT63sXBkbnnkBNwDPKp29
nY5DMfLOKs6faeoI5k9bnP3ZiETRAvkr1h4mVIutzihgd7ipEcBdrxkpaoJWNa0h
iHwCfuVmEDbXfMcAY2f5Cb3aoV1SB9CTga9LYPbsDv1QDghiB820MOUrnwT75yxU
rSra7ryNdWx5EULZkLL3CU11wlr41sfPWj18Bq7I7uqftZxzv+VLYEGsvXZfo0SP
YBoH1q4p0OERPPQQObmkr8UYVfHLWvmUn08l2/mp3aCVJBH8NDOgJasU9B5ImZ6R
cHymEeRlhYoRCN3C5ll4nOMFmLPDpj1feyJ6YnGkx2Mkfc0jk54MnnxvDl4+gV6T
PLyjD9VFA+tJSg8TAlmfu19uDqfFtRs/tcQLXnwIwqsMAz6u2g6wpn7coKRI4nVU
tQ/ARIB7cAffW3/n+f9ZCu4i/zpShrNzjuGYbuGpMmklSY4HG8wwkrHhi0IZqKSX
nYd6rpMg6eXg7BxA1t3HlJ9HSkZ3uoBXLepRu4f473wuqCKkbANmX//2jmJ0zJhZ
4UR9aD5+aVy0fL3Nw1lrAyHPNjP/dDXwgZUBt7G5FW+gV+z9bdG43NP48Jjq9PIv
nax6ZOZqA2WFopetk2XJXJXS1S7fOscl6Z3z7M3/OVz3kofr15C1B7LJM+Hm/8+y
G2uTYHBm3B7kKckfzia1p0DjLYZfZcECTm2IOZlJ7FiEADKx98jlE1NyymHkUrMl
6BA5D5sk6HmgK+/HenOXJ5j2xx8LU6AfsYwFlad2FUUCaxDamBjWasBz6TTmxj5l
oI0lOSznUB24si5wYxJVSqZJrnfGIOQenACO7uT4IWGcOx+TS77FjAd54m/Knfi4
8fuUX+kd8z77D9/XUUOgx/clCeG/oD/oqYHzEpTwkP1Kg4n8pGgcpSRjHS+Qo4Pm
Xo4+J3bi+1MoJziFNSXLKHqXdngzc2ZrZDFWjzqyl6z7IFHFCk8KkIqj2/sacBuP
XplqJIkLAdF1b+PbYMT5t1S02jNvHVE2lKvn5O/hsAjXLe1Mv+TmHKET311EFhIP
9OLRwZsShOsJjC9lfsZUdcUul2Axr2kaOVPrMqJTZXmWrBl8Syz4f+5ntDB2lwqe
e8Z8k6pk798srjI0AP4hKE/7FaG/aUVxRtiVNfB6o09uMJlJGtiXnSRcvDOjneCT
aqMCF/Q5JnFIyx1Yhvrl+dwg/c0Ku691SHpvWwoL/0bSHPOvG8DR4E9XZ2IdofwD
OjwyFNTgg+iZX9r1/AMQ+NDUEEppt8SKeRKceangT/Uki6kxreJC1+UJ9/d2otfu
gtpMAAUyyxAXIR7cOS1aHeLyIMqn2KtaE8Lmlj7vffXX8NC2JogU4sP36Prh1irY
Y/8bC42/bD1cJgBRMtSdrj0xym/asNhjbCaItXvYL9xv8WQE5Krz1D0wTlg5qen2
ijKI7ko+uCsYbHBSfGL2huOJkfC8dXxfPQ6pwlzWtRVwtq1Dmz9oaCKIwM2+UBLH
zV0cbBF/EX08cHZC6ztsXj9ZY4GtF1JKDTgP7xsC60NctIjB1XyXg3IYApr8fKjP
rwxLuVJ3pnEBI5Ny4bXPNer46B9WiixY5bLbIL10WdzxCQNzjaA2o6FHKblfFULi
ibDnAJyxlacgBBa9DS31LWFnanNAURRpPztLSoLZRFRMVu6hZbXRoLLFoEyTADC6
JJk7m3Kp7ED0SBUhxAq8x5wPDfVxs5zPk8mc7zaO7AavEl4utZasKV62iL6cLMp5
S8w378ywvpa/KJ6QB0c5if5zlucAIXIfc3+QwbpbPdwPwhpSXmfqNjMPt5+rdaKS
kNaiVKV8ItUY/I9k86HXEDH5c3TwY7/+NQOen0MlVDucGwAyeyZ9mdKV+AfMeCiV
VZ/n/Owr/01/xEn5pkoPS4gB6T1fMJ1h6f5ox/zzLHjNnKTlS4j1tToU7woHu9eK
Wpl2quhNVZWxuA18eUuWGXWDPO9Ue4N8seH0ntG5W50GouJJb4R5pcC9PDl9SaX9
BLwsg9KiYJ5z9wUZTjPrVXoJ71/mc2DPYIH2wZdLt4fgnZg+utrtHf6W9zDdC3KR
wIin/iiHh/M6NmKht3LBQ2n4W1m0voEIz+N/xc9Hl9p5ndDAXoE6ICfyrxBOjiZC
6aIhHxOnBFD0Ob/0MPppYH7/Mye3eGEgCOo8TmxI/5z/VjdcXh+m7Dc9tKI1jXwn
WbJLYIkfDEXaY+2nVHzldqt04o59bRDHzw8kxXna1ux9F/vPvbxIl0KD13fz7Pec
7gKwpmvudM3ycEKyczqwkmfeBKb7O6qlISqGRhczK33DgRz9UzLZAWryVHnOHfow
w+k2a6ZbLX0zJzhXDtOrQPz/aW/iBbl1jHtRSnpY0Xapl3brU6ZRIdAPb6unGjiC
zk46ew4viW5MYu+8/TPC87EJ0L0aEQ04BSvb2C3FsHnI3w/BFz3mRnyf5GlPI0sn
ZdbK5gLQvBL4co0phwodohNgbPXAd8vzxRlxtywaR3W5rIMSaDl6tZNMZSGEAb2S
5QsYgfi7WKrBbF+0wV1u+X1zwRuoLtQ9+0oehgKGrnVI0Ksd1R6xyX0VoMZTSu2e
fzz9iaLVQxIvko8O9WHHrGy5Ue2HUuiQsmRxgsHQ/3KtgKiCabcO/g0dMK+Q8uqL
8NvHcjGfquHUeLZu/CAD9xHZeCg3NRcSNzFZdkmMNfr/CEfO3b/as10/NbCLmY44
wLbxQAr2/b8qKv8eRddbhSWVmDQ+cPI3pQRQWAM/Lq7d3Z/vBPn/s1tlPqxFnQEk
4LIr3GekhR/UEjse/V0dopOWOicccQKJ8qIGXSCv4rrKHsaq+RAoWr1n9IXDS7Ne
QMGmYWQqpuynClYU0TIQLjUiX9HdyotWIQQgnkzrCjwzganUQzfmzDJDc+G1JKVn
xqTZijRsnwYB8cdWTb9gvoZfXvh8I/lZRRPfG7VcWcBrXuwnI41BZhUHYATCWvgv
Yi6bqm1WhuVzZpWx8dwXmE8XosR+nQHjjNGAkYTz2E2YXJqBAPnf1Mwikq+m9Dyp
0TBq6bJcP7NC+ZhGbnISeTURvKcEBTyG1YNjiHS7Eh52Kyi6Z+u+O8fLIVuBnSlq
bWzK/yPkfzT9nYzbc18JordvWd0ZuGLQv9KC7Rc7hqjofTczbFl3jlBo/sBofv4s
00wIXEksqaUKIbN/7mMZz5lrd2E/xm7DQh/aV7T5DKNQHigKDb3IT8Qj7rEZrfRv
jB18DJh0cdBi3x/2kXZNhOnDXsXdYm7xfuOlfPtYHOo1Op+HuJeAFq45xg6Yk1mW
f7ntvGgyZbKXaVJ1DQ3RUF4tXm7uUkPE5DFCYt5q2XKSYMJOts4xzJ7znwBx2LsW
Kvz8B64mmFi12SMyCM3Ko0cxzhUEpPUqfELpfb/3mrzaZxbiS1VtUQJPtrRP/+YR
my+0qHqxnYidfeuv+j+FNPxCOMSBiq1oD3Wn/bkUtMl7ZcA2tUsTEvrajbWkIA5H
MMeZRkKQgNv4cK/zOg0UhWKpnOm2Uyx4ex6Tby9hwmx6mPBzArIwkRnnr60Z7TKO
9lvvc2nBp+1iSJn9P9nYTo3R6lgnxOAJFuHJdhPYMzQTsTWvxUHsi1FbQcpVoGyP
jAqJIG/IIuOzRFASzuWLBBD3KwkRbLqcC+T39GWIeVzxn/UsohOIyR3RQEVlMkXl
D0MqEn/OkkaZAvWx2YZu9KSCpcKDZ+sfAeD/66mxzYA+pxu8O9PmfhrNgUKfrlfL
T2rDeX9UqlhhFTCrwTBeBtGNy8MpM6ugbs3CGWVXrtkz2OUFO+pNdjGwkeSwcX1/
C26OtMN+zJ8CbGLtZXHAwVeuoJ9q0AkDjw6iWaHqgIQ7twpDe0djGfRuRMB/5ozS
BXf1EW6w9H7UZofjJocwA2X5ryQPDy8xqG9JLIQlUAOvczxMpErwYNgakNInyWtn
Fp53GAKFZe2Jr+jmuswF/VFhnb4bOrEdVC1PIgsHxkZhJThHh6RzORfBw7Ca33Fw
T0ZqAR+pINfdYlqBXJbxA+H+7a6/cEeWg/WsJkUuFEJ9AYzlCQLFxNn/BtEp8oaC
jPJrVJh57YZTkG1+og671umcJQSagjVYoqlm19ZoMxXsbGUjGNsh8SpYMkRmOA6v
ZrHea66rtz/GkM3cybha5hZFjzhO6DQ+//btZNRdO6/j4MPavmM+pIKaMOKCTF/C
xq9/Es2Jp840xOQE79QivMjJy1M3nYQwhSqWujBkCftjmcNiZyHndyyi8uu5OE5F
kDpHvRsr0gXth8W1kMToqMBczUigTgYuXKSwJXxReLngPHZK1bNDmXn6nOstsHeB
RfwM7EiF3VyDiGhdKTcZslTC78w1cNHjkXRZkrTn83fXDEZYXz7hKs+tpOUvQ7y3
IrrSLiDigwwRKl8/G7zHgNEsIb6q6jcsGw8SKAuy7ITXLZnJ22qZHPZFiOOQtq4Q
EcncigeBp36MqoabmkdfoSZiNgjVCyfqvoToyehGN7e7ZkLlPABviApn5J2e+Ckk
dfmRalpoa0Ct9ngWAYMMVGX4P6IqFv3136JFhg4lDaqLizU1LXVpzUbe49ArV4Bl
glH+AVoZ9uwkRohjM6e0pA+5+zxAT51a0Nvt/FxRTwsoijV1buC80VVLaFI+7MnA
hsoyEUjwx5exhFLRmspFiLiKc8gtb2L7UJ9LQmz6q0u15PTn9rT6kpvja3Kc7Zb9
kfIBIV2MH2xwWKMriaGHyFkTd/3S5YBLJcclh6i2+Scqebn89DqG6LZd0VQ4hJZ4
bQRsaGEL0SF27nkZq2nublYGu/64e5TW+5jTPATpn3nHxie+FTvCKH++Nedv529A
4Swqh3ECTa3buBnIkDPi2Eir9EHroopz70fSaVbSJg3cINGPvPw9GqT3I6z8Lmgs
OIzw03oWUDfnSXDAmAljzoNSUC5yh5YYZ1yezmw2aYD+b5cJ9p3Z69QymQiPnNji
zHszCWcMWlGumL5OEKiribm35BZDeYBHurgq2WLzAAkVw1Ggnb5FQeYwZOlJYXLI
hkU4+1tgFvf/owBvwcS9tA2HMSBTgBMH1n6nrgEcDI0Lol/Znp8njHO/wCEKUy3i
HWbvKjfzMLbMPcmmfXHv9cOA6NP6WZcwhEBbr1NonkaAS60bTIgdFFA2MJgBBrX5
rIXXxUkNwf2iXbtIDPwFQQ7D05hogU+oBbMNhwPVmxvOns2wvHLOyFQjMfu/htve
IjJc6CDp3Nul0QWnom/6C/P4xPkMMuhkWVt59xXlbq1k0zbjuLCZue8SeoTL5zvn
xFlG7OsTxAH7qVRbtYHK7d+KvBG/ZOeyJ+7t8TT94rUAZe1/L8g39VtYr7evgoth
Edr3x5zbfPuCUJ1M/zF1exJ/BslJ3YGEaXi+B5Pd5vRDRpuPhP8wdgYwZu3FIHJs
Vi/9UPFQpI27MbB3j5lEQCAjQmKIA/xo29EIUsGPGHKAp8w2PhPCA8ZeESpLAfc9
9D6HN17xqvYV7BtZXDMQ3RgkyHbzVVV/oWwIvNmilA/BwigdsR/uaou2qgQxO9qL
QeTbRL3K4RuoDYUW02TEHOd7GJs5kj5dRl9iAk6KLSMqPpN1CQd52V15d3F0CiPS
QjdXlO0N/1Km6nckyEWWP/Mc11Mk4aqGhx/qdrrU8XBExplRSYkviz42A+OO0uxt
16hGPqlvUl21QncA9hl3C4k9n40hQOvQKxy2HBq+OXupVlG/dz7dImP+QXOGPvZh
bqoC7DhZS1EZNS1jRNN3pl2exIom6ypLdRxrDlHoacwkvLFbp1Dzwr6l8jZEPGrM
Om/67FT/XmrxVuAIzrwJByB9egbCyxx1uMNDkQRmZFtA3q4AmJScVDuwQNf/gzh7
WBBOIinH8Qu6axZJXOaETpwu51OAVJZhvNUoahX8qMTjN4L3qgbBNl5vY98byLxu
wUELXAG08i5jMuaz1b0HnF9C8dUTOwnx9cGmyuy+vl8Y7maNd869moQbNw2w9xDq
0ofv81R2tGeYYR7URy7kYWVpK3CfnLOnSddnCZXcn1KtftjLP21lBTCRpR51xkJU
uAhcFW34TMZzIEa2aKEKm6UHWyqFMuWI3dlcIj+oqX7ogyLt3Jt3mJ48MI1EpGEN
kyZAILdhC4pwsVauAmvhDwTSE6PkUoAFZ881fprVisKnCA507fSuyPw8Jv8aodch
f+U3FJOaxmJ2NRM6Uf2h3a2zCzb8vhZTPBMOvYBmluUrC3WL99+/4TeGuml4VkvG
yY/G9a4bOBI4Gu/TPOXu8XPxA/xeQMLBp+p8fZnM5hwDerDr2b5sWz093+yeFEZE
dhaDk3iaTGcyeMQCTkKmgsYmSGcsEXsf2lJi5kPcS+9MUeY3l1Lb12rG/aD2EIM+
OKM8MQPq+bj2/jKJjT1XkTuXDwJzDzTMco0iDd7qL0c938BQNd/YmrOyixL3lFZE
ttUgfoisvZolM6Sb8oInorTzBgBTV/+TKSxNLLkAUzz8FVSXo0Vue6nXnWg6TCwb
XV5in9yYc9gsHzb3iA+FlxrycWWQ0szfNvJCXrhh/0A3QQ3t8UKEn4b7sTE8OzJq
+QKQ6YRWcnOrNlibhhfMlI6DDuNuFpipAqkHcOCVQBWAamI8dHLXzdoqKNnQJ8/M
L5iTZgR55OS+wDX8HY2H2Rmdz5pa/v2REb+cAzSf5DOZ1yk+UtUo5l5FSePbuRqi
zW5gv4+UGl7cOS7jG69/j8LM/UYmIDbDtVNcaQI9mdWjkXYcXmerMIDcuIvIU1u0
nOaPfmkDN7r2HlvFcstH7x+WqAuP9NkXgvR0b37YXlyMbww1DgHET4Buk4YdP05J
r1A0DCKpFdG8AsLsvz0+oovoAt2SwGVx+x6ACk61d+7rqi9nbStVMu1tmssPi0aZ
3g6RZzSXrJ6KMmdMNnGTSDgrlChB5vK17qA6i4Q/Q4t3fjXYLvXfXz3Tgl8VQrfI
WbOqK86RmuhAfLl0I4B31BICZOwV8hCKibDRzqAVXGZDt/RowCFQsxru3QQORroJ
Fw/q3m/MJP2KuLFWvOvF4l4kRJbijrqI56XC/Gsp02oHk80/ycQnC3oN57oSzeFS
7kqFZuh4iZ9HBALKz38RkpkqxuUqCd5bbq5sVZHykmC7E3AmYzp26HmFEDc82Lzd
HJ8kEe3NREkadB2QDw2bo9/kLCZb7S3vG7U4M3C2658WD05q0veCcqL6JwbfmdwF
vPRpa11xGBIh/yGTA86r6FvpXo3CYbehUm7qn42R4EV50ZzH1BkNLiq1dVpPDAKK
zkoATBzeHoIWudkp3cYUBGRqc8xLyvX7VwRTmBC6VESrXF3GU6Eq8F6oN2Xlf5nV
aDtGPvzvssomClQdbqmW63MfYPqPoWJVVjFIMxBK0yqGlK5N3ewR1vLQiPDvICbb
dUutsIUTOtAPs0prDFYUj4V/FSl6nPxxdyt273mw4c94nqvt0pvJYrL+CLsDngan
whYUByPkRxO8W73L3FHEKopuRD3utmNPguEojJu+uEIrqb9/1NextzAOcqmaV1SS
uISBv5pThGDqFJop7NpIOMPzZvHQtPmxEjaVu8avGVZ4zK+BiM1uTlebqh8h3+6B
bxOiI4Rz1pdmRhZQL3oSBNnlX0BDAzRUzK3UAnBYnLKtxKBPAkgYRljebjm3E7Ji
ecR22tOSKEBEdcKcw2lSUXRLsuF8iM9C0L4jNBTKUrCgw1nWzysxMlr8Xu4gFgxV
etHHHEl1am0mPebIR9pxFjkfFlQFFrGPg1YJIyGGA6T96qXour2F5U3ePMYHvijD
Lil+xHTPM4ZYSbbCQ9Nc6vghl+LDSQ6SW9pkvaLUwlDTEOhFs/AX7HZ/XvGITAge
xbUTIAeeh8aFzUwMg3PmPhs3AK+1SN1nWyK24AEBA8+3dWAcXDmzqIpAjzUP9oUY
DAPGqdtHS56yInqotHXS+pEZ39nQ659dDuv+IHYAKVDQVKihRXMW6IPjS89eb6R4
V6CFzXfvxmWkqtg889XuNeYxkY1itnl9YSDbJAQHAsUl4wZqYAQD74QFP2HO4e2z
ZnTeh+bJPPbIIBbvsX1oA5TDK4nucep1QXLmiC/Y37WHCprZW97Tz0NfDghd2nsQ
sB5b1gm0xyixzoSu3LnB1a0pSLfnJ5DkotWaoJ3LfcaaOyGOphP96iqp49v7U2GI
aIEtOKCYit/xsdq//ct8vq0nBrI21Kzyird+6WNkwwDicDtOvnsiu6DialWLD/2H
EV38RmPH4NZazSG8NG9rxSJSysHWAX7x6WjlKT/JKSMSvn/joVRv2WRngv8pGi36
ZvPjA1fLTOG+YgwI4HklY+bt8YnEfOoH3fMw+BkrndpqfM4HVCeRVDd/Kv9JyX/c
vTT4egRWomQUuq+09POWkBS4OaWfQE2AzB6gC230NvRg8wnhBP/e7BTmaMK7578v
127jtpTUQLKS73NHtgii2dcjWX91XvPrWs8T3JUw3Fdt13vHnIpBrHHfoRb3FDNt
B8Bmkiohvuv24t4EXZCPIVg8MpYcCkTk94e4whE01R9Ya1AqqJi7te1EEXktKtpW
jQqBaooLuU91f0AVhZiUw/wTmlv9PVC1PcHUFQ8u6AUwX9vdBlGMJTk2rX9A17er
P3d1gSK36HOnrV0PX1eMmfKGIQ/mv6ctzvrVyDgufyKTLWtKqn6omC40UcFMyKtx
Xhs3l8ltZ4/SWwWuR6elaCVnIQWfZM9L0qk5ohg3ETTyURb61owmXJk84I2wHcSb
CawQm4TgYO/ARuus7VOHakEA+Oc6p89y7laxMb0ElqXSB3uuIkOn8Z4RLGS32XRY
AbmVehAvOaGdw198hPCXqdQIxkI2HN0fyLkST+O1ljgUH9DxKpviZLd2U4OcN89P
fySsLk1NZQ9qkUQ8gq6WepvQ6SJ4Fwkp+CRd0EOAVB75A3ZuIJrAwLfxfqbsxfBW
RlB3K8Hu6XJvUyPmkELFXB4A6IQE6nRv1pvVwAk2FKbgL2o5EBoH1V6A0k2s37Q3
Ciu2PBYkHRGbIaYxjGHRb6Ew2JYsrYoGk+8PSG2mN7yejBqdvXur9OJZKundYjws
2s2NJCdt6duv1QZj7BvwdzAt5Ec/U+x5NgI+hGO/flB5N1TWQKKay69N9ZJlD/6V
QLn2im8//ubz5ZUOwWWzfcx1MMDt3yB2tyw/zgJyaY1qRg51w2YwaxarlGeAsSsX
lOYG4pcGr18W5ma8IaGj0ZbRMiumrjsb+PxWMp64/cah4bpFOYwMMox5c7wgDn7d
gp9C0rhNeg27rCVyhbNW1YIhHMS4+ep5pQuFw8NtyCA2WBxz/7KBGNLdCvM5214L
s5DXjnJTNw1OtbMwqnjQCYrXOuHD3nbnC6MsXrKHQEIn7q4nS+4PxoKaAeHKcv6c
pUIz9fnAORiIKZeRrsQ/vLlTkHw4AZGQF9LVuwvb43vjj6qtbScAjCT5qt7EAhns
wU4VaaBMBzlvHNwzC7ZbGe4Fy505VDNrVuackJsMGCPpRVnBg66Gm6m/VUQVWY9V
zxkPQmpXLAS7ANLGlQJgWO4KAYIKG0ypdzalTAHmURUhRK1PqX+rCO0idxbbfiIo
TpVLjgV/SMtJERZa23jDcUkqGWbpBVyhKRIVK7YDv4WnbyiPj27jYZlWwwPgNVQH
cXzXnAsq0L/D9hYCLb/JrgzH3be8MPwrhoctgyZ/BUh+3D9haHPAgfvxHaoo9u2R
lqASRHhp2+n6q3eqXcKpNF2yCpryKl3IXdUnWuAKKDgjqMbExbSiLtKWTxg65GRR
HdfjHNg5wX0T6zgATVGj1HuUXgG2MbR8/AdEGyX67LJJlVYImN5ytFLtHaRex+iS
U0o6Er4n+VGfuYfOpzTvHKXYzjXZ9krP+Ptez1xrjtGn2KRhKvhCs/sZ9SqQM2F3
RLhiB6u0Th3s3XvLNR1PdLLLb7ppPwksAVRGEhQ/mwo8GRXmlxy6mScQIbVZ6bpj
D+NigmJYkGnxVb8+fOJLYeUmnhnl55+RuRvay1oCLZGbvASnd3uRE9h91pjQ0jz/
NMYw0lBuLbmI6i9de8NQuD2SNTcsqtEB2Z5gyXsiKPcQUDyz9NMPqFhWolYK3M4w
92DU24XgZ7yCYJIFW9cc5MHyHnURHaoaJ+QIwQF9nRY2TTLmHpiEEzTcAWWvQx/v
PFGTG8dqiii5y/clmJFOe/i7ltjIIdf5dLPnt0fdw8ANbWf3xy0ObpHdwJ3KrikP
YL+6IONlRb7IUudklo72l72dprXkcacKwEkOfr7e13ZjxbuHrvZxPGGZ+IvDm0oR
Je0FFbC2J6NQXkRyuOUxmPpz0NY+XQBFsTPwm1T/+QWmYIXVtONCyqUYXdoODKNY
l5RPtXxIr+BLFSFRXDWGH3NvPfLJMvwPWDPrBsFiHXYHvzz6TbeE9EjKFLxmidj9
7RJcoTaE7KZizYblnn8vGwpAbc95jtZkAUMUUWSg6LulhMHTKjehX1kY6jAAt4df
uD4n35dQftyixpD33Sz7K0HZcZDqLZVXfjFFc3bJocZ6qkqixlhYGFcbrulhWyXg
IcGN4zR5i7lMJfdsx1WmrSM0X4Cwy1PkD/e63yF/+xu3lYdhyZGMlhicLrCRSzbY
xFXcyix3CkSMLIMeAsq6uMQde3H+gG/d+coNvRKM08E2qPeWdY+WD2wZsipW+Uq9
HUUR1jx4rWm6cHUX5SGxwTPwwfnDclA69UVUqmhgTw8XuqsXJ/dno427tQN3v5o3
WB8YFvjERF/BM6TuZaq0L9TN3y1HtisnSJc4iIqHpGzuhVGf5H7RtlS+ceZXRS4V
bJ+6q1wv+3v8SBsm8I6qxiApeaZXFjhRyz5kK0kTww55iJZ9fYF4DRjK0bS4mIjd
q/rrx6mPXc0ypqdS/MFdcTt2tg8fHnaQsfPaqN3bEk1MO9eAov1Ui3DuIEz7zuwG
qXR0EIUSgL3No6kkq56R7JS9FzFDK1XEvc/PcdybDIS4aOiyiCD2fIEXKfR5MR4c
lFbwBZjris5MWiad87v9hIf3mK8dfkykULe1jrFW5dqaeQsCukqK35qjNtqPQBBa
8KGL88J1xy/l9Nh/EO+RcfUEpYYSbgtsfoorIWOFOBDQtJ3+rluA/1UP+iOnAbpa
Wpv6Z1mAx1yBt+tm2Wyuy+hf1l5dTf6nSr2CDIe6rmNOA23fl4vqpOKLP8WGY22A
7dCP2JKFe0q9pbtCiQQGDNIITLHAhPS6n0hW9JXh/2R0pAMNPg25zmKjmi30yRXs
vlTkhsGw97ApL6EBEc+h6w85aH5BQ/LA4E/NUtCt7OfaTxR4BfY6Z7xjUDQadW7S
1dLi06/fDSfp0T4v/PwvPZ5ZPMxvxYzWyP0ckvBGvifkA6ethfThJIp1zP+QclTN
5t1W+MGqQ8P8eIX0VyCRU3Fix0ymm2Wf/X7j5Y0uiJordwhvWaM3+wUHJv6KJI9E
mt3WwJ/XrXX05FZGinZSbKFWFH4QGCd5RYmwmw1bPjMBM8ctOcxKqm2195e0G89l
dHrzud4AZjJSACFMqw6WDKru/j7vebjEa1iVLvsS6vjX4UgsK2efN0WkaA9I3C5g
9THU26EGhJ+ZwQY2qUEYTxk90fpqVO153mtA1YaRl5+MKJ8Ovn6Lhh7rIcM46R62
4vckAf0/qyP+77waNY5FCxPDQW2aGpmC1T/acokCAmGE5CU+ixAfvXeeckELWLEK
1vQMgQo8nVnWkcC1jcCNLup1muO+OWRPgdvAw55AgkRCgcc8v4hCjjvrRvs7TTli
3M9aDoAIEILuQFT7p9fzHd2flH/LKnFdXfcpczhj2wI+U06ejzfrp6ogFtkQEwY2
6/9u192FJGfsfFALYxICuUnPCrg7KCoZseJsulqpfJpRBwqsRzM7acyXazWEZMtE
zYVCPcsVpUav4oT8oNI6N4fUxK7fQhZi8yLztTxWDuy7whtePyITi2U5WEfDsBCq
HyQuRGqFxmqvcYubofeiKNObKxqVBDjTd5L708ZkKW4Zz6K0qZQ/DK/gn2FbjhHv
vj/Ak3y7i0lNVJU1g88ZVDEg4KWo7qWeuPCu+YEvBg2A2YONErYjEDsfrWXJ7W7d
dwjUXiz8RcNMt1UkR+j2hlAmeZFtfTds/atbMwn/Vu0sYuzfGKBTAhBRS0pRyg7K
NV3xjsxHXv8fI4vR3sOJdcS9TG3g855s1FeqGQfAeu7MvzwVzEeAUx+nxZok+HH7
/+2xY1WAMP++/oIVEnuIKwrBDR2ZVz2n1xA4vv5mtEM8AxwyxLro7L9+CTPvsOee
GMhi1hsHMidiKsv4KhzqmGAFKeLL6eJsTItxt6wke7yJdPFUhZ3yqi6lKoyar+PL
5fbYgXQVrzs9LawN6SHirjdGlUAgv8Nk3Pd2jIC6qqo2h0YbBdmKQ4+tnY9JYyDg
gUWfUJD7YChfayOLoBsYIsmMI2lMutW4QB3bNGlKgWnMB5nCN0cd4JB3R6TAcEPP
qemrGT6HHUrz3ACEWUhenKE0o9U4xUy6luYjOc8QW24YAyAEXfyvkbJAaemQUqAT
xLSrxpD6Ly1NWiH01fm2ZNXMsh/oA1as0/VbnwneH9MSjtPeX8ZxHh6Jos5r+0fa
EGy+kZUrHop7o4eHs9LKdWSRI9dbP0tGuY+7BWp6IR1WO5I1/n6itlKTbyQeTAzd
WsPdw3oQJC4oJkLhqMPmMNA9tiMkizrEr+q6g09NeFtV6iBZhdEuhtap9+Io6pS9
rqhq687XhiaRAll3lfpqxspto3PYVeAFtX8EokuGdfS/gZmKhLUDFWAg6gpajb7x
Oy5BPMXRurJ1OCLBdcvAfjljGXX6M8F/YvFBOV0I1L6z0iDoxg20yErBINU6kInF
fc6OLKgmlqiJ8puOqVeWiU5MItaFUm8BJWw4mi7JJGNVmJoDOU29XXBnXsBTjc1F
uO5NpSs6Nsgd+P1ffdDrCi2V/5c5hZO5T4TE4Zm32rra1gZ921J0Dvu1Nzsv11z8
oWOGOuDv5elVuZZNcAywgytZaSdt1WXwa19K60amg6aKsJzCBgno+SEHb0QuJYKZ
X6iVisUz6Nqg2D1sLixYBOf9GOLFJbfgFIoGOJq6Tx4N2ZMjIegAIzy3koPuKp56
O+vro/g/XuDBlsKO83tAZ2oQAUdG8nrd1e47xmR2S1s/W8l0tTn52tQwa2uAWmoV
0rQSkM2vaXUMgD2pm+uj/pkYdsrVMTkPhfLP0vadcXSSBcxSqakJZz0v2WBAHpp6
GVoHZNpYNumR73Vx26Y+Aa71M+jCdkJFedaYW7nJkjDDe0t9hKIS8jd6+s0KMdrP
tPjlDCBj0fJeE/c6FHt92E/4smRmjhsNn5s+/sj4aUXRKvg0QgUKTDdyk4TLpIvp
mhgTziA8GvWg4+LPtYlMlBKOKcIfEGY211jALJgzu55tVkmTJ+WC8FLJW42LJ5ji
KbXjvzan1uVVnt1dnJCZx9RD8yl1+57bsYTnrw18PRlyEfmc4omohGRMXIgLLIoH
8R1UG4PQUPtrhuhmVCF2/b1e30rladwyiyX8+p5CFxCvH/5pMiq7e0P1QA0bO4+e
eCLKFP6ceXJPoz+ztyTjTR2M9Ycds9EZmmKanucaAoleF5DKLaSsQpUXxCEzaXYk
Rp1fMbTlJrLVpNTok24lUeGNUT6rgkxbJRwbecKDzvDxd4+ty87wXHPFhVCULu4f
G/swzAD8i+dj6UQEcbY0Q5RwXOsOL3GBeNZS95eAWlD5Y+pHoXu2//qHO41KJXWC
t8jjNKGT/+KleDse3Em8swymeU5E6M/lXpiELUwPM2dUwI1uDXfZw5UH4s3xis/2
KxzH6j+P+xRQy64uCkgQ6+c3LgveE4gTvQ6Zj07UHFIQpfdHBPnMJDoxT0+ia/Q3
az29+BGRJpIohAQ6TS13NtUio1bge1oeLNuNKVxWfIobgXM8QthDt0tna1naqcQo
FtXpzcsug8Tp2m59gF6dJDORa9ETaE99kMFXs+Sx/9/72YZOJxnCnyrSmI4y4+At
hLqukXepz6fIJPRCFuXQxEXK+bg6pNLZ6Vzjf+p/JT2MD2ZF/NSfrHECOxAFzxdn
OnRHZu5jMNUXEmqrry0U6KAmwkyYL8tmdJuM/wVxYJiRqsAaLAYlrr8rJkUeg6q5
x2Um+kISAC9eajaoZPQAH5WyiHgffTG1TfxOZWTwsylsN8/rp3M4xLyR/9A3Nujh
AsoQC0DzsT0Ky8V3BMcuG+LEk1f9AlElDTQTo4BfqD38pGg4IN2cN7P7Q88nrlu2
LwbqkJ8rCy18Rjmj+Iffx4WbKtovNwVtwzfuIfUFUncykftqdoZ005WtiHcR6UCN
RKXAKyn6WO0yStJ9I/eqQsWS8KLlE6XDzkIj252GjjExCYmHrm9YXw5FZNrTK9IY
9TRXcNIUzNLx1PO9BvkyX7q1TFxzqcEoJDmMJxEID4IHCCt24zwVGJLzi+3eUzIV
myjslRX1kvjK3C2DM5pGi+EJHZB5UUlXa1wzMjIw2oziJqXjdoyfXtd6G+jYnGXE
8V6+4+aXh7eBxKKmOR/Ulhxy+WDjMbzZb2Dev0qtUSGC3TSIOh9LuNR/vPVOkQ+K
GZSHsQ2b75Gyr18IOIIo/XCFMdJmeDs193Do6CE2TasH9+yeXyFMFjcwBJrpY38R
TRpTNm/6iQdbXXXLMZnd6iviPEDzzM9vXv1XUECYLG/vswoptyg2kuYLFgZ29a1U
vmRz7ZjfEWyV+T34RWFKt/6BgbX6vwHfAp2bczwAfvhTFVxdcBvhkh8PS2fBK0SC
SButQYgvlkVYVrhd7hfszj9pGUKDaVTCQJ38JJL6QUubbtBVNhUqZ+yjvvoll+Pd
vxt1g57yCYqN5I16DVaNgZuNFCvbc1m+8k3Lluqbx3FvBWuE6zRLgMA8xeVhZdDr
Ir8ye8kPYVR6/q9SNO1CETzN9OEuhH+pUJwfa93DmJBjYDgjk7CjntY/kz9npbKL
23eNvZn2dJR6ldNxyMizhfQ27HN0v9gHn+uzh7DExkL+wyn/vqv30hmqEUSeDpGs
5rvekEX1HZi3d9lzZEyFe/LTL+/pAH8TyQS78T/mWpCE8lGKoghIZfRtfoDdK54n
qJPmiNOtCJHSS26ypOd+ykUdrz0t0sg3Bzt1/TD5OfI8AgpS8DoKzaawySAYmLGt
Fx7kHZTVgJJ/WOXJhugasGtRU36L0Mi40tFqV1cBXApg6LheS3Gd9KW+yjPq9dMI
xjOaUD8M6lKKa+Sfj97qlAyLMl7GjALB77abEik6EK0nZC4pVbuyT2L6eScdQ4Fd
PIZLe9gZM99jH3WAzhJwkp+pexCzULOUcicSa3n78YTWigCfTv84cOFf8MjAgOsy
k150GdUzRUUWO3leVq3iEqk4tixbeFepUgcNAxDaAua6XqUzAMx8cDnvEBnEpvFD
kWl6v2DOVSl8Slwp9vE2ngydo4oti7LGyf5zN5BOAf6TGkWPbwakcH+u93Sx0W8p
9iNZMz3B6/mBqlg7uPgftIDgdv1poGY8QIUhZDhBveMloJ16tjwcRUUSjfTfszTt
k6ZWhtoMJhKxuaEUQ96JFdLLm2BAT4BRq4J8YnxPipdGrey5YJzZb9N0/I77VGan
eL7KNB+75ZqvK8S+XN0pFkDmUutUi9qi2UhJ1irzecL6Vec7yFxq9WITW+8aP63Y
BuRTsjNeBmxShrKl2T1Tu0MskHGdkPpGiXpFfetOm9pFBLT3vL4I60SD4P2zQ0P9
v8bnyN1rvy3z20+40i2stv4eK6ChcCEIwbQdtL+6Erbs39ZeR+3B1WdqLY8l2WWh
4SF8LrOVQG+NIQ9MA8CG7x3HKSM9RzTNeodi/uQ675tpbx6ruCMEGqXLaPGsOmcU
7y6I0MrjZWgyCLamkh+izFayYrg3bdCNpJ9WCkSSNOUGsfv3wyJ+bOLKapBb2Ca4
W3pzeAVUDZkZl+isQ5RdaMaRpvefO16WCUOL+A2ffgNMf9c92FY/diX7Kt2qGuEZ
DD4My8zKIneRnnIZ6TNcz6rildNSozAA7PtopYVlQjCceIdRiqnFLH35qgmHcIdI
dmGoTHd6lwx6k86cpkF+Fii3p4z917BgNr/Zsj3l2HHA2IUBVG0WcQ6v7Pgqz/YM
wmIBgmDJrlcRI/8NEaFeOPLU0NwDTDF0hhRufu5hpOOGE1GpnFaSJrGRlJN9mg4V
L4Qc2uPKBGfhaeCX+h2JDYHWOAfKp0LhCogb+xsvrX89vXSzE6ETcE6CBrkqy20V
htq2mjppFGvPUcoFSQ1xR0KLAuym/cMg1T1B7kQjKdn0uSF89/M/0502QTd37/X1
iHt+dXSolPGQNFnT5yD4F78XT1vFT7H3QazNM1jyVUvXLWAOjGnZrVf1UwaAnvX2
SZQ/ef563ppGfhyl7hpqxKYSL6xqEGD1l9BuvOp3W2aA63ifUq5SRNmC6d5UOuaQ
QjYKR+CnPIxQcrPDKWk2729M5LYr+5fj1xbKbWyjQIClwA8uSE032Y5s3YFnFNZG
8mg6DfCeA0AvAEElvrnXJVaIcbvq4X1SRY0FMBNNuXmwxSjD4sgdbzpFh5EkWb4d
E5WKr6YKK3QZxdrd2Wbr8VVnPZ9PULBeHSB+BH0RgFe3bgUe694NlSPIsonH+X1q
zCexnOBlwEVqe7TJtXaPhT/RoFxBWjohIY/sjHKpdaE5N4tSeU0Ohpz7ikRtM5jc
h4VVts0CuoBeoodgzF7UHk8QcJMWi1Du6nkuEDtMfpVaYvGO7DNz1BKRgHC/7RVW
Ad3nGtTegDFOchnJFIAXbVZRJT7KOYPxJ0lv/YY+2EVHQBACG9WETv2Fb51AbDJK
vI4L/CuD3P8jNWKAOjYTyu+fbCfaAOvYZ30mrNsHLvdKIPL8infvLuPQjlalSwOS
peMJhSCsk45RGFJXyAgMLV1tJxxnDVu/c/yRo5Nx77LLO7haLaGK44a+IBf0YFjL
e28wM8ZbTEG/A49D7lRrJ3AEiop/2A5iVemYfWi7ZjHMNenZKn3idMVU+mQofo9S
VXDRKaC7HbCXrlRJeNsbuDmPtlD8/+fjw4x/xc3K9+/KP/Qk1mDu77jkwxcfCiW9
YdpdgW46PTdURO+2Tv0RYyQkCgk17GXQNUmngv8eLnPiL+9Tq1wZ7xH7nE9eHM4i
FlVQnXN9lQBB0iJQIgzv5ebk8XMkW1YAjjorkP9cly7YL/nhc6erHQBZSxlJCZBI
K39tbwNwlpa18v4VGphaFN1AFopUvlGH6kv+Rf3vRixBUu4rd4/9436rbIKKG4xa
zbjurNkw0St3fY0FWvXqAiAczCrm8fp9uGRra3UdbnFwZNAgliub0QaWHiYJKX2c
hKKfHXqBQbk/hUZHhtp/qg+eh+It6ZxjIVUZIZUff99RxYNVhZn1f61vMM6j0JcO
e/+6WsYfWaNH6KtpXCe4JouWZYAFYfQDphsWWEj12atqllexrYjXo0MRYd1mjECN
/HhELnrr+oueMgT2dCH+gj4StSKE3LhqxK3AS5KuAyc//c2CcojYbpeGUIgndBQS
9+1NPhj6dxhwrH6SxmsuTosUjH8j7cjJW8eG0OGch7y3gcRjWHI5LC/Ve7CanZqZ
J3V5MoLakgjSinPmI9bMniVFS3mhjV+1GTZxbi0Dv9K62hOL4QybivtFcWhJpgn2
IBCJUlVoDkSk+yNsHJdnbgtH5/dVq6qp15/ftID/S+9qqitxX4QlicmQC8ZSY8eY
VMS8ae74z3VlZN40qt2q8DnKXq5jFZyIlEMSgpAJ1eIwXdzAiw8TDlZCP6pO+CtG
V/RrqKqUs8A1OBSHxcg/jSL6dHFuW5e6jXp1SEmvBeG/g5sw4zZ3XY5a6wV4v6LV
T4oab/jzME0f8da86igRZ9m5/rjMR4JZv2dgZFTEkDVCHEkFut5wtUCNdtj5WrMI
xQF68DHKfkEm8uY72k3a/5w0uBxDY71IBJoPQPYfjRZ3JC4W9W4It0EsIMgxgqwB
Cviz77cuIeQy0PQ/wisunn8d5zeFL8+mDM1Y7lqasAXh05pLj3UtsU0ZZ5oCRt79
oHywOu3v/HQ2M3q0ACBdC89/gXZ9kHUquDRDB9qFxtoLve0Sb8UYcWLoobElU68H
A9bFVnOB1B5tVvMmpNlog67HeB+voKGzGsL1MeDAGxG9GuOnJwxSMowRUWweW2oh
NpNieu7liaNOMMkZ4/Et3VJOH/30h7FIw+YP9O4N20yc9XFN6TfoDljn005mQlKz
bMkuXNgCn2qz5OqUTIa92V/N0f6TFu22/3Dmgtfz8X+O1Bpf/uHqc1G0cmSOzQcH
hHhoOK1+EYYWEdDa1bPhxuIbUM7/pODMAI6xTrgT1pPz8bLyAI2HwurmjAV4Nzk4
MVaMXTf3XZoS8W654y9IDjSgUjALEbeFVXr3BVHLGHbUn+xd24SSoZi9PHjNf71m
NJm3FaS5cn6EWV2zX1BHyZ+6bYuwKXs+MT84IWoJZo8w1xH3+Fh3kiPAEklqHeFv
eOc5dqPPMIn4Z7zHhu4KgUVQYXMOM+dZzWgMCbPMy44H/SM2M4Mx/Lcu3EfHdxmA
DBly2uh0f5IZ1GGySaDhFJ10vni3Pv6appEaHd4cPyTmm/bgBvpcqTsaahbUhCOF
4qufUqm3dmLOsKEIqHSi3WdRWDoAnIpt9tWNp5zBKNwLB6UT7fHVwUVqG9yYspuQ
r3sPkQjLg/BLt0zwWUjKHn8JJAu5+N8KdQbVhIUMHp2ud26AzQQOs4CFzhn3kcNs
/4H7BWdcy0erc3FrBnzb4p7/tMJyM1Mc4shBvSnIB3YBZXiua+8izCl+VxV8Rj0q
N/xcDw3yMhPF8yv+6cZJD6PWQlQXDoZTrcXI9JonKJZAMqm3Fg+CO4nj5rmyqAMH
aaKagc28U3q8l0+Y5uWD0Ji28egKZC6+PYhT8a5GGoTn3A7u2UTTQTcrIaVramsP
VMN7wvm1GPViLUcGAYKtRwhsV/0iHEF2DZ9H7A1wFCNWxmeslVEP5vMHIs29BmX6
ihaohMlJvBIO90CMEWeyQ3mpFSXAPch0mJxHxsFueLrvl6YrrINmREctfTroMWqq
FGFPgCaEmsLgqmxFlIk90DlsfEVbS7l+XC8ZF5kEhOoDuOT8B5cM5ind+p38BnMf
topzTSKHRZnAHTVcyUYkF2eeS29Ok9a73k/sfQHt96Dt8d8BHA6Ntq2e0XB1CCsC
0x5i4AMF2kSuwtvCHFWQfhatiZlv0UOsG3OtatUWHbTndQNWIme8LxL2q1OzweWq
GOSPY82lc/gVyHXGBUxqhfaym4zbFa8aetfzPg26u/YbssXA+t7EYX4oZzp6CGqA
thgy5nSSfLuu47B6y8iIqmCAsWv30o2dl2/5HnUqY0Ue1Nkhqp8bjb+rFqdWDxBd
t8HUCmqyq7/PZZLXp8Ug6ewelgzxVZeHO4IL0tyy8uGTflZ2Guf77f8IrL6dsMOw
uYgJ3w4tT8WPmJ+7ZOLaNNDHg0ayTqKUJOpC3AQs9u2uUcC8ZwPIhqUeDdDoxGix
XF+xAs62mg6zJZ5B3XLTGcR0DRCcLXPTevvAafZdH9T62/0UQjmJVWHNSR1XdHU0
S7uGEPRCUBeCetPeBwsg3WF7eeml8mAcKviCDDwDKLbGSdb8cGcMpa1X2muU+7Gb
5u0YQiMR22lGbBAu7QTPLXcYcLe6CD6MJ3+FaT/qYgd4/NEf1BPWU24CEKdMIIqp
irMnTNClanM74VF+bc8B+JmP00hbzriLWxSa1PIpCaOItoIL/vinFviufkcjtT67
wx60WAxUhtQ3GXbyptBjTCKzivkCHKCNh7vDtjTF+hmBRrya2AUG1+bTn1HB3zCQ
3ZTbi5DjxzwgAxzNrwzHRQYyj/jqBC6TFfX2oWbkhMxpMPqXdfWAGMzEn6LCKE4D
qxx+AgEcb2hC9bNhkRj8PUDnGMEPTaTM3of/KfDBXmvTT6P8MhU3fPZYqK9P+TBM
4xLnA5NsTz2/pRcwDqXZk3hL9izB1ftbRSJEWnYCSFUpdcyQg3BC6d0bSqJ4vD6A
arEeG5FrTG04jjEFxc2aif+Ztx72phUa6eI2cx99Ww8yyPhYd792+yIY6w6g1CmM
Q4LNr+3X44WAVIb9Y4SR6eEC0ridt4kioCTVhn5rCrqvHjXXTQBaVydk8d5y2cNQ
Vdz2PPf+cwaNITdnseurXGBvzIMkarr0ziMluU5Mv4FuAmdKauh54Bd4WxZkGR4j
AjinbPbEjmbdoYJDkf1Vs8u//T/fmXdUl8h964k66Xj+3m7rD+KEZ2GX1q1ITfqR
qT08SZJFD2jcivFoPAHZuNSoZuPpPkFuYDCIFkgLGM/xftD3+Q7zLWmLuvuWHUJB
QUhsntQsQmjlH4X5YXHFsdAEOtkLv7t1NxT0UtMIXERmZJxkgFn6+F4OLUZRGYWG
0cCiBcIny/ns+V/Wu2+wIqBlS8PR1VGBwTVfqYB3tG873HwupMSH8g+V+clhldVW
qTjJsoUipcUHtKfiGjfwxqzdPKBgo9WqEvpAwUDrgMVQrryX4vvchuLpUdAnoH98
rF7EHlKSp/Lh1FmIUSDA43DDZGRPsATWAEZL5cvGF4cVTAZD6iMyvxEWMYlcsiL/
7cA2sjOFt8PQ0vei3c+iAqhinRtIreVBx8eNFnIVbNnQPzVJn6ZRF9k4klTSWgmV
3XMELG5lB7jgJXECu21LbTYJ7vNCzRGz4KKoUXi3oSaJUsA22O2LqELrSxsfRq7Y
LjKZaGyhndQV4SFbVS0utrqWfT7989tvAjS6k79NodKuqiqxCP3gJD/PFfnzqtu2
8Ke1wr1ZwjznPLaaFlOoSJm6JnH4wtdJLB4WzwcpbFTI46OGbOk+gUbaPCgLaOiz
BLAHMPYHewdgN1UdRvRAyGbtJi3hHtXeSCg8Y+FeeEZ9Aqcuh4UHcjJHVwkAf6eM
W/Q+UUDehLyEVOkdwzeHJSty2xn036fj/OIE8zP+0W/9VqGAi0J0iF9B7ktoR7x9
BUvrVmM5jy5WZSobCegsr5IDGTJNABgEmZZsQZbDQkk7xsH5wPDYkueT7n1VRRcM
VxRZwnrrS8GcoD31n67k8jxPDoOYckuns4QNLY5Iw9Vq0Y/yQmIhcWAZB6UGGp1Q
QSm2Cqj4Oxn+NxsA0AHq9H33NIOgH/KJYx1CVYhopsEmXMFNz5H69bKOwZ9NtR3G
1OGHI9NUfCSFlk4+dXS5pcSW3F78ThmOcf4C6vxbx9eIvIfx3BiEnwdXmAnlSOIq
9eCCHq+8j8rs+tblnyK10dCrpTBgKMZYP1RQ9Lcm+WUa1AUmPc5hs38wZFRmtVxk
BRmqtQeDEEye16jLDTJhQwsEMeRPihqfp0pvJnD+2r50rJowhGzF9FRyC2l7PFHU
04Uya1TMEpBTgtEdVxgcbtNDKPl5QHvsQoIpiDh3d/5NKscijzDmydwoc7+D83E7
+b4AzLGxlePhLexn+5Ipf0IvEe8+D5TKeu0i4A1iP01fnuAdTE4zogsw48dNXrY8
8RLQsbEiuuUu8bYI/PYDMahjF7ZOE++f7YXzWcGKS8pJLkMz7iG2ZYXa5AWXxjj+
5EF1ta+UOD+DGv+22K+XWlOdGkIvyCFfRsZDvTyUZ4p2+o7O3CxhOWyviA8DmAQO
ryfZTY+Lk7sWQmWvvismIAclAnlznLanpPD9vLBJ5R9pnpp2I/XB6fWAYYhjtHIV
64VB5Gc2sKNHEREUiqCz3uDQdlN/b0wOXmasJeSwGu89PMcbv6P+INW1akaYJHXm
nlKj+okF8eCWZYi4g22uYotyhWO3C2L2wEwrHHLJ1PrnIVjWESeeqR/j3eLndvDk
CH2nXkQsL0Kl6eAk11dwKlhvID+8XI/VbgK+TPbOHordiOn1dY1wQ2SF/9LdDXDl
EKVATyTv7WzV6/6NegcXkUJpZrkk70EgoFrvWVZpRsnBlLXiEgjHEOLiXSqImfDw
lUVWgMBVCcntgqVr7RYrJiUET9KbWTHnNiis5/ng1u4Wr8k3a2+4TD1dqfTE9Tl9
1Mvt+GCMl8BuEncBilYfHStO3qI9noA/Q/ZNMmxsUtTFMb3bAEMaaPC4jGUr5dkT
I+bpDFFXzZOTZEbq/9V9WTP5JmXQNw6ayhlS2aoPYG9uqEK+i9PCOg3hmVQt1Zmo
Vmp5ljAaFTj5sYKGcetmq+bWGYUsLdoixKk+OcLu57DmJ6EzzfRtXxGvrZyxXcFS
POJg0sWA9/NrUUCDohcXxjyAYq0dDsMQlEnCNx4lkx1Kph0sqYGXd5dSRJx96rZy
vgZkq3LQUtBb0ULUOKxiUjTE+tdkhBGqZcuUumkL4wWEoxsBf4MLasw5v6NDAlGK
SI8E/NdrppSDP6YFMZSmS2cVKIGgJ+Wv8ZYx/HVCjy5vvvZsczV1x37XN6PHSl0w
2CBMZkN+hwg55U9mXLkulQmBZ2vSCc6q9prtnWQKeWgILrubJyWX+uK5GyoS1l+s
drX4O9oP4Q0DI0rAihBSEZNAU/YdKj6f6mq8fAFHYa8spdMIKic9kfMt0hYj1dOo
GmM/SSqj56JyQeR/Rrl0XbNK8FiX2x59dPZWH8PdD3dUBeoNl0bGrXsvwytllZ/F
ZOMBkbDpNUhLLIns8+9/prYKWyDYELZd2zaTJJ49J45dnPd57/7d4c41n/Bra9iE
P9jFRTsaD1zFhaUR+GwO+WOUs5O6oQHtlP6FiSnumpPXMYATLMRILJyne49SFGJT
O89f6bV18E5wyGCGxSAfOvFtfUS3Y8ShTlc5mckj2Gq8xWzwS8i9g2e6nosPHo2+
H1doVZMddxPSX4b/8i7ogVibxWCWa774wII55TTUPrEgIcykUuPspzs5JbbQf5hW
9NVGiMBwncsZ6oOe9PsJM66uaN/cLYMvUtiVPnyyKkNHcDwFbjwYfWMBwI9qgOEc
zOcYPTxq0k1qHBeq4UUY5SZL2qmq7QxKut5TNt28HpS1EhONyGbCk1ieQBhtWJrr
xuBCmklGHQnqA9WF5mCarDKO0zsL07Eh+HflKRWI5QB+fRE3Iu1U0J3KBcxcxpFz
xFQBvET69QbxFdj5Mz5TMSZa3Pywo7Y3yw5hjJRIc5dIccyvKYyi6tHmR8gUgcBt
YxPoQBUg6wFsmNJUbNQvgZDCkHJDE7NnpAhOd4QTcpFvOX5wSaAonmkvuOOPBUgE
CtQOoREgitFKQQJkizxWWYzkc5bmFrPrbPasZXfKrlnpfTThjG6qNCS5I0A/R2qg
qATfGmVo7E/iU/0fdYMpJheQIPIEpLzZPNAU6d7FqcqmrXJ2MgNuwUCOBqC1OmOt
j1tTd2LpZsOEXHaIqe8felEet1LrCgnbNVzIsFAqAs73JIWDkm64qETh6znhNLyP
WL1ldRvAXj08xxOZommk12GiqzZFSZkh6eF5zKYH6EyYjGbyByg08LO/CLGISMbU
dNpvuPlj5LrWBJsFJooPA+vrNq9ZIUzFGd16jUzoQCIg9StTgxjvTBeCEE3PBFQb
+OOXIGd027QuOdKBWCj9DWuPdHPYWBOpYIEG4XZ5TdhH3WVIkrZWpGRR9MLNBalD
bnlt0hrw66rq2FOfLkS8wA013TX987HxJ69YMT+OixtMbA1RYcGkaVCyhzVtkEXG
s0Ya4++tGCODu65PuhLq90YZhH5Vsh8q1YKHDPhZV5AKpqThLkraYbKjwCJca4rj
H8UahJvMX4sFnANgjFkKmloxwlzDpUmM5X2yMthAFwbH4qAY1kJqmNIg3iN77Uhe
SrwdgicYVMdQYpsccB07XoaOpe3DoZeDV+SHHiXOWMaQUcVmo4RrKjnemjRBSiV6
nvO+E7aE51t6YEImHw6/VyMrVyHKUsuaHPf5uVyDcHRoSp/wkiuov+PsWFmZLbs8
cGIkZFdOh69rjTYDjc4TMJMZPqsa/b4MdSZzc/YXMPMv7y3Ln0AqKoF/rm1Ih7OY
DMIicobP4N3WkJUvVQouS7pw0mIngHHDQSDAbgov8DiBmk9J03TScIMmhU6qwP4a
IjvvRydY6eckkd4o9pRa1L3Y0TRKGfMhIpoMf/i0lXzZrtKDJJgN1zkgG4TneSYb
VWj5lOnjEDhcExK3oRH6vGEy0JbkhB0dsd3S+YSshtC6afkGCW7ej0YlFsfmOvai
by9vcEif4kRPEp/CaVa/W0w2xgUbbA/AdbU9hPfcnPaarDEOsW9rjYI318wwYFIu
TJfQWiZ85hSPJoeDuubmBwPXluqq5tWz/ogJxKbVJBeLm3R10VIIf8WKsDFrgFEe
Da3Kfb4qrT61T6E2aB2weo2DWRdgIySqtw3NX82JK3Zs3bYATMxTmy7h3pOiv7X5
QGQwkrqXTBynoFz66Lezm/FeLFkbKLvQXZksoMqJ+L2l9t3ORHruLfU8eyVfWpGo
r/t6alUTPKqNdG/bMzXUTa5jI8MVE5ysqM1jSuRoFeddzgotW9O3qS+OSbP4L4uE
fLQ4yRT4EfnQXGJdm0+5ziZXC4s5y/h6AVEI3g/HpSSIDdeDBfJz3k+6GQFdTyYI
7bLtplLXsgGhQVhEihTyYNqsC7mb5dojhUcK3NvxhkhYC2c/srRfQy/e9yhGLCEG
CbL8wty1e0wl81YzcC2wpCGXkZ5xjKubabb6QZc2aW1sv5M1LNkmd9CyFTYupQO9
BC8g+8c0OaK7gGZbbpSac6Yir3Srhyf8yhOQi34ZryAzonyQkT9R/aXXD8/g1eDr
/7ZwixmZFsCVhKWgwrQaZ6FDTeJDFEFslGu5VFJNyoiFv5c891vGnR9Q+EgvBlfK
lQkPP20/ssQKEz/G7IcGxfie6PUC3mDvlpbK9lc6K8Pr1/Y1P/aNYVHLJazP+AEj
ZSvzBd5Qn7TB+9XkQEDQwSjspJSrFjOG5ZCDPdHnj6yK2XHRVkJ/RFR+42FGm3uG
tYfsOdInu9ymeb1NBysr5PFVFcMjVJyUyRvUbjoksornBaMlc7YvS0ecD1eQ9IGd
vFS9cNLC//0zuor49+xXe9Dpg6O+1uRrOVSYqIOrv4qY3H7JVviCyc8dSqCz4q/H
tMMBcIRV7tejXY6kBGKNylx8WKs4zk0bnsuQ+5FS0o2KulKen/z6v9O+Hmr0XmN3
GQHy/D2ZTDjbBZWp5a2fWZ3DA8thSWvQsg9lJc8ipi2XYEWC+Sbm/Ee1PRhlape3
FiQABcoui1KticefYdLUYteBEpIxwWZLTLw9NpK4HMGZmcchiThcv49OLFmZvyo7
RIMqwA3hqmIpcHYs6dZ8TSCrYZCji/2We0QyF0n+Wp9XuABh1jZkoHtMAeQsrEPf
xou7dX4nHlkYIH/8uh8zS1QjbxzNFwI3S0qmYkS3OCWMvgjFxGqwrXcuH4pVCRkI
01zs/eMVQiya1Fvh4m9HlPTkeaMdnwz36ErWT/bcJsH45kHflO+d9A5pmuusebek
VUyDWDV+I/IFi2UgpDU4dL9J8HumEwTLDwnJIb+XdGJjUagZhEXkr7TklskokNWk
4d5gSIInLBVBbcQL0PqJcGFKq4YVfMUWvNNOv2CHn7Nvpw4KnzvrVItnC7MukVEM
z30/DaCMjIneyM0aWQFWVhloFSEHOnjiDIYVfelvMs6LscOWR4E1QZhMhO+eucIp
YEjNrIovAUb4oRHMC0KgjovDqxNisOzYIYp6Qi9sCpsONgGCcxVXO0sZed3Yl8h2
vnJrVGuVifioRWO8ZJadnkThcjdXIb7EwlSr7RUxb8llHhZq+2vYVp9G7EQccgJJ
AmU5TaqDIYD+Zx9SWzNZhGWveBB14tBvoJ2cgxlhZC9QPDa4Ii05BBbCIFZiMYYs
3CK3sDh7+ltMUZABEh27+Fe/lGArDwoEpz8fa7bzwIDcPnzXS5Mbn2OVl1fYSvDg
i/pyeLmzgumV3LFxAEDE5PGJctJsENKRIBc9j492nbnTGmS4VJK1fyYPWqqVNqaG
4cHmdmrhOeEomswO+WD2VrS5NxDsGXwuaXNvhbaAA0d4/Hv/pw9sKts/sG5+48Y6
3RTI7ASFA5TVf6KxrHBmfYVfCQ6muS3igTVJg3NGvZSjHOLYmZIptq5VH+pRPCQ5
6MetbId3X/juGSggUAhl7ePkD1u86PENaew86Q3gU30VumX5KT/lF/dPKjL+g7QK
5fWnkm8QnvkhhQPs6TTWi1nCYvNu58h4Ar56bW8m/F4nrblwIrWAbyzD4tsdayTG
hq9dCublFOhmbqEimMm3oAtQQIHq/4PYvoepOVuu7TMr8OWXWYnP/vUqiWAmqh8E
wThRp9r2eqO3jDXh61OPzUcfDOM1J5WOPC+Y5jrEagdYzIsvgof0TwCZReUR0/7z
eiLB2DmWkfZo7tB/qDCu0M3k/IxHJ5jJ8BbasTqys39nxhfVn14d/FflIY6zMFIM
bHhfdthNGkYW68fsuQY4pwA+C+5JpT48eRHWFZACKnBvQHzRvk8rQ5/+jsenaZOP
QORG6utgYhWM6mcUdpfCvuGj5YiHHRiaaftTjWh8ykfrBGW3iM5T249lRPDt79Gg
P2/iP9IxUOcEEVWVS3O4rpKnRg/ZUHRLkhHtesh1S9TYipSHJS5L5wgZuMeXNQ8h
h7WmXW20NSB5IXxA/tZUrTpedNPG9UUr+iZX42td+cW68nHVSL7oG3WsrSTNMF58
s4+pS3nlqicauE4Yr2SPljsXcOBMg4PtyQSCInPvvWPHX9/t7w/+gqk4sW4Ei0SF
tC33u8fNUGo/uivp2U9FhiVUi7QW5ln92YHlrc+m2JfJTRjdBQJ01885iQVCxFtw
zjkNO1Zr2z1xDwb1OW5lBhdRQyDup8wWjZjsuhlt4WSwlacN+pFrt9mfjpkKsq56
EZYCUy5r0fLOzkBjzDx2xWOElTKUw5iL71j+9ZVcHfZb0iATobaG0FgXM2zhMX28
yaaJD53R5HTT7AO6wGJ2wkK0K7uSTZQyWY2eo6qlzg4F1DZ/ETKCyoqx26jHAqjn
mtqEQwavuiIGU9uhGhvzJviY1+BYkhHN0XidGRXUtbUqmLjW2w7ALB7vsjZN+rEL
7zzlr5dMWYBoYJDBmzAyD1o33syJkwfNT6zextUNCdO8GSqe/3mUuS2UT5u9vmwY
kCRMsymSaQ1hlruCHxbwGFeozzb7Jfb+gw/k/RVm3qz8cJi59zdXKTv/AO7qAbbw
aZDCvtLuZWhjjIU+x7xKSAsKCGzg0jDQWZEH+k6SDzJftyG/J6QEwnyjvwl2rRgf
EPaPW5oNnQtCuh0Slpg0aFSoAIf8yQLVYB0rz+x9cgVg9CYQBk9lHRlzJoV8XeBh
tvAAtto2ntBnZ7dFk2B1fSqo/6/6ldyQOvWHxM+Cq01QKNEsNMCyUJJjPSbrKwQ8
dIcVZi6y/LKZzHNKpbYWwGHsRxscpnpv5ha6Z7zZ3jnPrcktV9OR6VaDVLLHcuL5
ognrhvi4r9QoQ3nzASxTFCcyqY1WinvIJa6Kvj/yFlXtAbI0MEoCAtAXX8zhCofp
nK+LrF6NWizWCzevX2wW4s8KOvdpqMC6y9lprZJ69Wjlfdm/U9wsKVVF0quGxdZ+
PVSFmMKTx0iaNVXBzWoWVX6/PmiiO0drkJN0Fa5eNeNHsE+O6XWeBPK6xn8eiUtj
mOmsEjMp/mTK/8c2gy9sNvTs0GxZXh/7HyBPpSlqB4Z+CkJ4WMxRye6M5KMIvHiN
q4YnxDRrApCqNrDogTfBbd++b10tp8A9i3QkLskOd6dqvxyy6PEPKjG6iGv0qJQ4
9lbDDQS2+jQlAABr3a3Y4l4Rz8qTdYHSL6fHBDCBR5SeGsuf/8UJIxWt1HKajSep
xfMOT08n37wTMuVRlnS/1mGaUGp8Eh8wu0C4mqYH6hAR9qGBWepfrUZGzMaiTbxH
VdgYVePFxBY0vna/SiBnXpXGcsXXL3ViTFHnAesgq9wAd42YyyUbfl7t16BX+wHi
eqvQewjb705vsuanfYwQvk7w1ABMo3ktd15nP0+f0NvfGlH0nYQyeoURtuNjVMz4
Hagz+jXduD/pIg1eYAkHFRTSkIlOqOXHZA3+fuqCElDQwIQqwGKuI/XzChxdolWf
RSnzhVwH5WS1VkwUCJEVpyc+2Q5qm7OVl3VxYhl1nFX/qGbKOtqzubnGTP0p5Xdc
crL2u5Vb/gsyS3ZDlEHF81DvTkbGWDjwYgObKS++R9l6K+zPbQREx+eFgw6pOANl
D6E8flMBYKlXzZCyq3/k5eB97hAWph8/vtdXLPbJ7pDmfe8bJBlm/RqHtk7ZDGHG
XMUuQ1PRRMEMwJ47YafL0zACDjmStY0y5JajdTUxWI9car26AHZjX4Yz3Zbf8dZi
3JJSk6QuIxee1K2HqKI1pwhfUTok1TGlmnmoaO5BuV6B+oBg5BAk6JtYpLYvSl5s
zcTvczcBAAtdXfdVVS49boRZPFr/ycDmwBySwYoezs+eFdHc0UWTNhrwNSlaWV/2
MjHOl3X72OpcpDd2hku1asR6jSNpdxcGFdszk2oHVyNpHw1qgjFu/UgIxiru/Gs+
zlh220Rq8MGnwIAI/1FvN2IX7XXHp8K1xgaCQqPqA+gNCAs3kux8wgHGIq7d26if
lMEolYmk3f/NU2lAlLYtY8ehWQ56u/uNylquFoUaoHEI7f0rURNAUjEmZPlEQ0Mw
PhZ2u/UVZNT7Jngpkn9v3lo+zarqZFD63503I26Ry/C9GkRyXze9D4Z2BwYgalJ6
dcOMhNkUcE4H7OmOjuL+X2qFaU4sJCf7ku+RaJnhkbb5M4d/OCqmbeq7nKOleA55
XBB4qWRHOVICmqZY4UXY7PIfHSV3SU60m6oSk1lU2zOERhtyQW9IW/0vv1/xrPHy
LDXg4flBXtn1N57awuurBKDfKNE83LywxxwpuqxB6nOD18/rY6KQUJ9Ig/jJfQzz
csvhH0UBESuHATbhJ/igIqAcljJD5orILv+AcVZ4/jy7T25NlHvUzB7rj01ZwRGd
OskwiRibMHiDWBuhIHPkVDHGwEVdIBYT3jHPPy/YCuTMIqup4IbOZ0uNRsD+jnIP
R2mo53uuYUq3B9bdACtjyr3zY9TDD05vkPgaBH/5hh2wj0PyMO9oOJFwSVklP30k
TDC2D8t+Gkprgewad3pTz6P5u0VBdmn3uTReUhk7lzatrTP9BZr8KfYhAYg9BI8h
150yQmqWfPaVEaTzY+oZ6B885+Zu/w3vGpt6Yvw1OibF6L75+S3BMfl+/XDPJy8j
t2IB4fkMU0E46zxPTvlGPkPOqmmeKrMAPjyAX1E47UQn8Zjshm327hDLIDjx05Is
Gv85ixGv+kpaaS/ndUd9HF26K0y4WgEc7en2rF8vNAQ4xG+3OaGuxS6tQwFAgxpd
vIzJwRCJvMM68ZxxPW7Uwg6bS80GvTnGq733svcUPveW6wS3FPPMR5SIR49bBals
mTD8FVgTJgJG/CV9qOaPkEHudWRrIL6xEoNFTRsSd0vED/YpimX6lSL2MX/BYdOX
YgfYFjNoCPtTMnoA943hZhEr7oQGME/rwCtbuOIuzQfytE7VZW72jnqp6LP589xA
xGiX0ovVD9zqtatzxHAGEzce7bPTh9JY5YzR93DtdBGXMoxgADC0gsmccHyKYoLR
o6zw4j9XBE/B02bG49+mq05F2j70jhPhBBdjU8rgo7vVq/HMqwLkbcYtNtrix1GV
Bg2rp8UBoJjjIUzm/7erH6FSRS287GECGhbaMLEC8gCu6/PVX0Pt1iuIO46j1l8D
68rsTR0lBf1ClLL+Yf6Jum3Tx41aNMw5s5PIIKniusI3FQmywhwQ9t/m3W2XLMN0
WWdo1BMlx0MXudFAeDu4eEcSMpzlkYcalwLlNpLVS0UW2CekvCdq5NqERPXcLd7l
JTR+04n2n4UOyL+exupo1AqiurXQB1GP0Dh2mMkNSYJNs+FgyHlZ+LYuAXX2CJ5a
DT7Kqvhi9NWorAJrVcZ6AtpQbpL5OfkuK3eFRaqixbpI9hfnKvMoYlpwI4hktjyF
3+MFMucgMMgg6rDmX5TFXfIs4ORdpurJDaW7zZN6HV1BrZZtcCcdjVF8coEObAqS
oiKv7OQu8hAI0Wvo4CfoYxh/hiFHmelGMH1vo0hdi+vLzE5aoDV++QCeEblVNEQN
fehQvERi2RfvfmK2X2qrxS3n4TyHL7QJupEJ7sY0vCChVKTWp6qhyZfLinV/WrOd
fuTJxRVFxX3ScerxkUgEwbfjjLjMDi82Ue4mLxBL7jxIcSEqk0AYAdVqQh6kI3Wp
aXfhMgQVadyZ01Zk9u1VuE6lMO9gpX0efn5e+0g4TEoZmBZ7v04b96ivx84sxgV4
3O33b1xazYunuJXRSTQfYxhY6VifN6vp1zWQKmh4/nDX/wDhqabh8mPNC5qwTuhv
Kbm2i/64LuV2gZEWS1SL/5VWQR1cdBvEWtLRARB9kLG8FBHTrIv392xslhmkE5eP
XGUaezokzND4XoV+On7yPhtpIPxyQ2gOs8yMYI0qQ192HkYzF/H2cw0y/I9Q0YqD
lDU6TilpEU/1rAcGdt93smKQfeWmUpD7tSL/pryxTm4k4aY3gGfjowDhmpGGPrM2
UXNs1ESSY/11DQeeEAg5EXGIXo8qbAME5jYhL+Wcs0b+3kjXDjgQBLICLxW6Jq4B
cKhdf2y3SkyBbTzAlDohbVNandyq51HWSAsosP5wNyM7AgsPEjX+O+gs1Tp0m3vL
6N7RkGz4Xbb2PyBCZqjw4T46OgTQ2XJuRBl3oF3XlxgH8DE0DqAvi4dv+wRQQtgq
pOF+kavB3cMDBHdumE75grajfAKVwiMFeXWy9+V1tQtYHopx7k8otk7t3p/n2Mk1
Z4xJ8KancL/0SbQ8H5jTGueZaNI/zD0DZs4BC50DjD+IjK+kjNTS4UnBt6oEA0ns
sa51zV1vzpEHmn09PETMRk3VaGW5YodP7F2dvdMCTiJ2+tCeB5A6Qn6qjyJSJYdl
7/TSwwIt4zPPZRHf5JC1996mHCVFmHry2svwRG2DR6SL76z1RDM6JEm8zxV4fAuw
ZzOLuQ7A2bc9L7tus+0ZM2EkgFAtSHkj+p9OGn6fD8D/6C/Og6CWqUF6AVYmYZQn
+HSf66WF2jkCTbAmUHUjtbzZLaY1cmOzMeQimGkxxjA5JOmwHzVG7MByd7SKK3L7
4cKa725L/6CIpbvXutCP/fOIikI7tgb6Du18kKRx36XCQWUt15GJIgEyqi7Wnzgr
auV6qooqfjOn1obBhJ5uESP69l8bOo9AVOwgIQFfvuN+vqT+ih0eTcHWEDZzyuwx
L3g8k6pcjlYzMWe+zblbAo09BFAyaEcBti1ARGdNNYgUwcHzvmQm7VP10g6YgTZ4
kg7icHbpDaH80tS9JAOKuC5lBL4DM+qiu8bb7h8GzBQf+ajXDxMrxHMaTwLmAZKE
f+ATURD/MXh5u/6sBLTsKzIicB7CLJawH9QafIl5uY+mAEo19adiQImO5au46iX3
7GjDbcXyYenbpXNymL7PDNFlqJaSIhLqaJXimpZXpwLnp/u8/NoL4bwvMUmodj7F
PiKbaSUITMGmp9LLajUCHozn38BCZCf6aEf5ZVZBs1ovOcj6XL+PjFwHhC3MIXws
a3Wh+2LWK8os/C/0FepXUwn6soKB5fhA9waILUfdKgNz5lXMLt6syQnPYSBaxGlZ
Ebp5oQHOt8L+tg0PuR9jGkdxgxYmtiomo3E06ewVnOd0eHroclxiXI6Y/N2fauM+
GxdvHLgq27lSS84Sz13xxDMQnepdmSsZ5WOKey7uS9sTPBYVx4wqc/HPobOUo9k/
qJihFkisoAZpkUdYO00nw2HrdIqY5ls+coulweDDRWGfsHW7lC6lCohCBsvn1IMD
DnOH74BI2ZO0d3bQVNd+qn9atj1twuYZN7vLcGF2yY86o2unIiXcz+3G/Ns1H9FD
fIwYJO5LC9xXjI94zu2YtyFamMCZ2QbjP76L/5m2ppWu9Ehw2Q2PyUQbXWEBAv6+
bzYQ+IySGxTa+AbvmgCnsrTdW96wSecVVud9pkR/CXxNNypF3G6Mz1+1eH62nAde
DbwtrYW20KsI7SrPNnP854lslu+qa3uERWP+g2rocf8zAYQb7avkGCaLM2jI/mWN
EjxxL3nKfIxvqhavoZlnoAjufD+4DaqzWxBSY8lByuddiu3Xt9DwraRfPIq6+nFo
9LMCqJDFiPUya5/kFgZCeAkaPTJBBD77GheU4WhSOsNM+G6Vyi+/iLQ7D4bB+QOb
HdRKAeaq0eQiuc2LPegOSh0cgwjayxHs7Jun4OAcaqpttOjepq0sOVCkOXCcAInJ
q9tW3b3SBLMNCrvfaQB4DZONqkzDBF1CB732p6hqqWvxpx0P78fFpmLB3KQGsM7O
7q0kVUHbU+2yDWk7hSf3idRGpOm1C8nSPdqwWec/6JehXDtymtupVlkTV/WiPMBi
ryMLKwWMRpGZE8l4RGrQ2OgJCin0Qf5UxYn0daDvy5321BdG5oCb8LtN7J+tyfMU
ZDPOAGcBY61TWqkgqtkk2EuTSBsooxsg6VoOhChhO9jvYhO4fdXdHM0015o8aSvS
ml8R972lsZLjJ8PeLdHzjP7Cl60SPCPyss7EpJ4k8AOySqx77JT9V1fdFHrHGB6y
kASVIEiD5w4tCgEzTKE6m1nT1roixVwqiQ05sPUsnZxuWix/u7sC/K2AftZTNMe5
0dDTF3qWbY/vAxLwrGZcCa05f2VNcnAdn8KFczRYKcezQs+9amMLsyzBO0ENcbQH
lrYKSzJkvW39q52emMCaS83NI42MOcha8n75jbtxlFxGaGxrJNeitRtfV2a5kV7M
621mh6A/M8wXklKUwaoxlYL2QvxEAPhfXhcZ83XFeSGSzCnEVVT0WOrmVw+xXstY
1m2DAzEhut1Iv3zlyHD9xF6y1lGD5ywFERPKbF/Hve2Xdns7M7WixZeaPGBcUeVL
9I2/7YQP2nD+yxb38VWcY/o9bPir+M+mGk4olICwswfyxM2CKP/LV1UT5QYTFUDS
IqPsNsW6JDZjXTEV7qVFFQF2tLkFZ/aYTDMcJIpkByixCUD8PZhh2pCZWV89CUX/
59uyiFV5NjyCjuut4ZAVeV2w4PVjYHHbBpg++TdMlTzOrUUVUrDW+1VoNCVTfwj+
y5HhxyFyQcOLdpjhTrhAoBvBV9McCRogLs7vlbrPqXstkWyEjjdKTptcASbOjruz
5ZQlnslFjdB/BjE0TkSQQw2/oJh59OzdlmkKn08LagKIfLK1QhqctG0zrvuqZ1hi
h9e4yRZ+T6e4UBqSLwEvX7eypOpWRddY26oISNPvTM3aXFzWVQirY19w4JpAOzx2
KewENW+kJ2+T1Vty6TFu+B11HUQvr4v3I/EU9I88tWDzsuE228naR1d2rMMYtzDr
76GoqrfLm0ZdQ/vu4whfNJz3+qLpOja25j1HxXdzgoNQ8sq1NBCsgksIcFNgBMBl
PyZg8tT61r1KIeVnV/bTDylkI0CVV0M6VDkV2l0M61Lj4OKsnZXuKgv/P8DP3khD
c84jnYP3Ae8h0s4g0UukXnLoKtdJ2O604F4Sl5HVo/6wFjhAfcWrQZAK6gjHC5Tz
OMEBXhz7GfCQ1pHR5LXZ9RPpN/knMYCphwhiKzHIlUcZnOSoSu+B7C0G9LMNNqaH
8D1r9OSUT9Xpvay5LA1ilxOBwpk88dgD1QwIxGMNQG4DEZnFdreQUt9UTaR24UsZ
vT5TwALSymWoaH5XPNKHL0tPGTKZFUZ3yfeEfxyYzEaAEvY5v08bdTRvnX9vUgmE
fPJIl96yxAFIkPQDAnZhv94n2SnyKi37pAdDaiileps0ekh9ZnK1foauGvxyCh8X
m4KL3fCWxq3DDp0azIhs4vNsV8xAevFmRShIJcb3BK/I7spqEP0Ac+BJN9U6RjYO
4fyGG2MrTMS7ykd5ffs7xTE22ALZ3nzBatNF/lzJmG0yqV00e6tZq3Wxc35H6JZK
Dj0GcYMixgiN+wr2XwMCDUJkrbjjmaQOfSYNxyBuPWRH7N4OAZ7AjPPrRiepXMb0
0YuvpBM0uJhnwOda3zQPURmOroQk28yu5THmDe/6Z8mTdCoY+Vh5Pn/D1mh+zG8s
q7mnhhGDNAm38l68mACzxtzyccaA7xu55wIjL9cg15iXhjxea+SZVQBEb1Phlnzt
7SWN0VX3pK4Zl56I+iYg9QaYETznkItVJ+T16FuIn2X2r3ArDBazwJPJXm9x3U5p
jE7WoEdjMUrWTr8VFn4dEYPXaKXlNZlqZC3b5692PJfkxGbLAeucGBXokUaOqX4f
seXVb7ydIH0A1aVyXsZKB3XKXw+cyjeyAAscS8gQ8T6/2lQLyF6ZGaqMxwVAlwrg
Ji8BTSeRk//5yvdB2xWN9BD51gob6zmjSpFCWMjbjXu17zGisBqvpsDiRgxgodsg
BW74tjkQa9kJDAItfI3luyYXmvkFQImBXobwhme+z3YMk4nNFirkIzFVDMb4Ruh7
yfEjCekXkAC65skQIUmGrT0V3ChtqWpLdbbaWbwfc6UebU4IM8lcrQTu8pnwKxed
onNOBY+5ilk/bjoFIfNeuiBq+AU1yDM4PXYIhp5wNveGDYX/+V9nBET54mAu1ZPk
5zZ932KpCacKuvP2Y6EAL4c7aohOipFrJeKr9RhZbrg3T8hqsRQrnrKjixP67rH7
eoGnUTk0PMZpJw+WsaQNw8A6tRygY7RfRhK84JjTuKZ/b8Pqvz0fKLAbCrMwQnrH
oiy68W7o9jQbqEFrM/TDQUvD2TrJo/Us7OvPNOyNiYzE0EpgZqEPV82qZlmPVDHl
b6ki8GFjRv2Q/hHDbVy2Jyw3E3IQbq1qY7uvonRnExFgOWEIG2eMB/NZYE5uRKlb
PmLmAFUVcwOaKg43XCc6LSHBB7X2PSLTbaiROmK68Y23LJ1rgAQoU9jEAapbHzQC
cN0kIp34KFybOLSRQyEol2/pKEjShKb2EB/4uIHH/4lEc+Y/JGPwoOGrvd4VLXNF
U3rgn5ba9OIgsF9F70tpXy922B0bSGVq9iN+t8A+iACbkiYVUcfflWJsaBctpZvy
47vIXYoP//JQwp9AGRtRxfuFyYx8HD/hVrWq4qglCsbwrpRmaMVhL5MJUfYSC7+M
JqxhZ3TGqBtJmjuNbvOE9J+vGZgK2ozoTwifR60rqoryv/lDmLUrqcZuBwZ3TWPd
PIWZKlqG4SvH5PBlz5vbnerTjmw+fZ45Zs64+YaZtyZ3i2nR+Z4DjYXW+dxw9KVC
eFU9/vJDmRVXT/TC32yfmCKlWkuS/yXM2M1lsnsPPCXLTBAUHBtPIxjGvnyRyGEA
Mzr7UGSkmNqz4YvzPwSUjn5OUnHt6IwD0bDhM/+frtbQBaIIoub3J70yZvo2MuSM
rJk8J0XIFo5cIq82UpLazb7nwbnFkAAUOCJbQv17Zb35gzmVAL36JtThJHyn6hwC
mVAHLSspkS4ZhTCZgRKaMicZcmFad16q8gogYBa9BaQhvFdVqGPcniYe/5MXCuTb
uZFoBU5b/Us+Y3cdEaXo0EcQoESxyB+goTS80qNwx+mPq/Vh3FGMPqKHOSzMkyHf
QPU0ykT0qseUCVeLGfQnC1FQoTjFvX0y9/BMJfkDdxncSs041ntJabbQrp4Hcmp5
veiU7eJcMnvFZXmySfhgm6igmM0BGeLi2KeJ7M/RQm43gwvyDfJ+iPNsSzuVJ9Oe
mVm0ry6xPfpR7DmQ+/IGiU1neGgnM6/X8w6D6i+XngRth44dGp+rU2kiWuMExFIT
XjuFKfsHEr9qKQ8dKDgKx+CX1GLYfZOFbhgcfioe2e5xs01Nj7u3kyktvQOAlJ+s
AugB1v0H511Ve+Kmdz72ZyMuh9/v15lvRSFC02RP8Pi53V5YzoqWdD0e4+Ujbhwr
EmfqwXHLG0aXHng+gpQT5RxoqGUuN6CTMKgG2oMeds7WW23jWwr7u5RSijOy4CQc
oRr2RAYTz9DbEWw4T5YdYn9woiODU/YhB+19ah1gyVNlsf+h8n59OuRnK5TVgyQ1
txwNLt/PZg2+mtusQt+tNLWZzL2Jx44kHXmGSk9NyNROMi8pzdiavWRJvPEDgbzo
VtsHuGfWU7l0iCa4fRdNmhBEtBQPUvLc0gYKc3QV1nA5pJXrKRtTxEWTGgmjqOXp
mJo+QwpALriDQJDeXAOvfweevADNuILLj+LehAkQA+mes5NIMuiHP+NN3EK4yGtR
iWc5KiQcnzY8+EUCnsI8fp9ty9bWsZa2Ud+QO4W7M4fCIUNNncpWQCS3SO3JO6+n
7qypuL/w7eNuB7iTQ7QmQalkWPHILZ6gcmqzovbFY1Sc/YXfq4Am/1tsY6U22GBZ
LFXUW+2mNgnALSm83ELHDy2l8cFtTmAKB8SKQUiTE27eC39pT6jSvGvIfWKURvFi
Ru2AvwRP2AaKkPWd+Dl6fqiTH6flySx4/SLTOxLf8GHHVN1HjF7U+bBd1V8vUPlH
oj1cLHO9uwfzCjKTFoZB3YupKQC0dn+5u1fuk3xxBn8FK+/vJaW31E/ti69bWgNR
Cd0ypgr9fIySr1UhVhZf56ZV8/OwfmqghTcvm7TncSl4H4pfYKl8PFoP9XPVNHh/
HT+03sI+No/yUiN/5cWRCVmLgDRuONljJx0ArfHvqTgwrq80W7wIIJ5kwTYoy4WR
g6+BE4Qx5uchV3FwVT6f31/82muyIUBljCfIfQVujH4QyjSoRyTSAeUoul1OEKNm
JFJurhCXTqm9ed1QuFAIQZdcfJ8TyPVcD1wAgih41tULChuR8LHn6tZ1fMViZM4m
sUpLsRgJ9T/QvOhE3hQqrZwAt+SWEctykSWPHK7OMqtYQCv2Jrljw+hLthOaSQdT
zQiJhyB9/z2pPi9JGW8xYZDPf+9ygbqHBaFzgQKiLiH1bIwQBU/8u/WoqBnaHMpa
t/44yBur7K4KlPZ+vROYv95CMfu76RSbKkKMoLUeFNa61DbRWqKitc7/zdD7vF2x
snjvzf/4okGJDIUU/239ofvhSLnxF1DtYPL7d9SZgtTluY4qy//9IxER4p967Y4O
saBkWdHywAHSh/V0scUydXtfqCE/nSFrXxssq8NOmvPz0Oqq4WSIg6xrKJQYzlKB
hzLmG/8zUF3KffiU0Jm9dc3IwfZci56BQCwvUbBwrsBbeS3TYdoei21VIzW3m0Sx
S37dvEZEUCfHqUGePPv4rm8y7Uq4bEqLn4J8GABjNhZLeI8lERJ9GoByRuV5jLKe
HXWN4ppAhITALya2VneNPXmr0mwRsy2rcvNhVBmvBd5PMPh47LxtaFuEwSTj+ZeG
xVeIwAZtZ5e4nA67PBw8ujsaAqTpT4TIZMsLYg9ApU9+ZxkMTmh3+Qq/ZKIJ8qdo
Yl5VfqfI4UB8RgMpH4RyiEi+lof8rYg3z9p4GDU4mYlKE6THWCJjXrL5xV4NLAJ8
Wz7Xu6A+i/3tzOXUycl1E+HVkKwvCtE3QDj/rpaAYqLzVghf6JEOn5REqxEw/MEJ
m6+Gkpx7CGh2otTD8fciSeWVVOVgznywheeeCWCSgQ3VdH0pUJgHC+G9s9swpw4T
PT9zql4xjIrXKPURH01oduxxzz8GocWMGaIqcxKBTyG7mu4+NL+jjcQYWERazLQ5
uaGQlX9Xqv+Km69PbT9pDLnhNwA9VMBNDnQ354w23ikH+CyA42UtD/xJabUOZkED
C6sk2BCehjOXkuCjn9iZk2rOkvN9INvvZ6lEjPts7sKDgvJpz5digAf4K4wbxuUZ
kUywRJ2wYnt6D+8YJ3oD0sGxsOzItGt0D2lbRYA7Q2uSj1aBfZ94aMDi4oPuNORa
F5PrJN6P2egfeStH3BjuscJ24ltz9MYpkcubq5562zaGqpmGSJBqCgKLpJsSAcdV
8e9me22HCnw7D8KgV30tFZgY5euSbQtLZUVypalPiWU4eN7H69b4+QvtfncvIe4u
doR/SzjgU5QANeYcC9M/49VA3SLdUDGP+hksZKJc3iw4aClT8WBtXvVEmAbYMrc+
JVfAH9YTrNTNvOY+mIDw+mx6STzwXtChlhoIdUN6OqRGlQbA86CAhrxLrIbF58z9
C7wFeERauV900MIQHZZHquW68lRsYa0pyvfILQILWROtpRb3icQ865+U7in0bzDe
uodbaBT7cPgcqsaticJdrBcNWj4fluHGjeBRWWqh/LVutwKO9C/XjzJhmfTJAi6f
XdCKwKkQTw5gbSeg2jYJ6GPwZxkGnbB3cgch5nSQj3DfixbckgHfeQmpImN7SOUt
jA81u/ipskZ8H4sE+lHss0FrrAX5x3rnVCtDtbZhVkkOwLvfBZMT546wZDDdF9GO
Uz27VhGjBrTK+xPbjF+zZr0XOjjhl/b3c62qgxHHwagj5nA7jA0IYtHwm+1SGtZI
dzrO2qE/nlhkcTDqAgFCllyLRQzAk6m1febOAMjcx7I3uA46GrQBeFTtLPr1lPIw
HDTacEwL7KZgtcw6JIj16Nk/J9O7w0YT7oFd/e2uNiIF+xHW8qF1DOB2+yJw+G5d
sppAToyMfyZaB22D3cAjSF+GoIhwpBuzehnxmiYz2TIw/0M21vnmuhoAurVDOY3H
UAnAh64D7cVJs4pyj4QD9Wx7dXPb3T68zBcdge3+fwFZ3YPNwZFhaIU4sn52AS+E
qXzFV5Jz1WoxM5SnQiWUlizpeti8kCuiCc2SO+S+Ff0Q3I4eu4f71Y4nP1QCgRUY
1crVnb6ADojJz2aI1bvi9UPbngQHgbgqcRsuEQa7Bb4Kn+xKpLxcgJYX6oG687p4
FcQk+6Sc5IdzQGS07DeyFZTLavBQVVazI/orKGQWHCbjsAWFB58OOk4AgLCipz+C
Sgd2DupJS90QFCkzZiO+eSrDbzhW7j7UdZBfTm2CeSpL7yTHDy+57GMBhszLfxJH
MbBv4L7FdW/ggqG3peNhRNyRrqikX1OYJNObNZecIjBX2E80SSY9h1Nf+RiOHfoD
TY9lSFOODJJ81q2t82icgMOOJm7WMBI3xmBSnLOmIILblyV7uLfS79/Qd1JKw409
YVAQ3yx/GxVcmxcn3WfWC2SmMpItjvlzKYOrR7BsvYvbGq46HBUdUBtU20Ae7lrD
Dgb1apSvuCS0o+mDnAs37GhY92van9P59paXabK55mcYk8+bLM2fobyGicuFDWyb
+k+BWQxu1UXHHS9pd3yJ5iKs2YfXnmGTP95AOy+ahi5uIg61A2T71f0KsRDYnllg
or1pTAwwUTZPNUQw3dbNtSsG0YzlWdri/ZqS/j8CmJRuoGopX+EWWVHh9pNSYizF
hjBt5oQ3ayQu/qt0gRxX248gdlEy14CYloCq/xH1tmRSbqLhejWj0zFIZr3x/n9D
AqIf0H0O46c8rCQ8idyYr2kzn0S+oEaJV1/nihm4bGXJS2/vDwQ0mIPYPEU6r766
AR52tc2PoKUYbkEzWKd8W+h5sdbcWzuRB65vh7BB4YXF+ihzbYdVKrboAmHbCZf3
q+NssAVWVvcqbUJkLUyXDDjBuwD43w41CQV8oLpqRusHkonsdU7/nvAIrutDHle/
MG/xWqAwevAHKWBmLSGL0/bNWvUEuA9VD25BTwosgIivBtPfYi2UMl2OAHEb1LML
YVDq//C0Sb9+Jtb3qa9zHbFCsEwl8cyTdnDDiPn+UTsUIr5oG/gvmasPXGkg7+GH
SDJ5sBnH4rJw/JALrtMTbdbRtUTHhXypuATR1/UVoePNSChw1mG3Ox+m1zSDdQV7
CTCLWlvURr8xbu0+JNXwAlW0HZi1AaD2FDyrA7osV5ILAEoekOiwY0OxdVpFExt3
coabvFUIClbLFCoYl+NvAmFugPZW9o4SjbQhCG7yTJCEhvesjibtT9F99wueNWlv
yOV+CgMliywb2Yn1+omXyHJSqRsmaHO0elrPz3mfLImMUuoSPjweqetNZX1PSm8t
mm2WD5SJYCRBp6JBnKf2aniVf6ihIWrzXTOgSX2+FUSVDgSsBjZdnnpwCsnfBUpc
1WXmfzJqvOHI9ciBSl8QIjrtwE8Me2l7p6TIz7JuLNhLczssB7VNcueFF2wccQjd
0XJIF8SPUfVrus4fDXXsLu0B6KvCUrO1hHFU8XDiDsGzVshImRZAbXyVK+KFGrxF
EtDrmCL2BAQTAENr5kqhzJFeaZX+mSVu3n48KBXMxyJWCtsXaw/gqgbKj1ApX7/C
ffNdAZwDwXh86wfBAoJqQNsqOGw7xBAb20h5pN9mTlRoZVKWYSaibbTWI8+F/1WF
rSyZWUazQZVXZX83h1ZNu11M+QC0eyFRrOWojzA0RNEmgBMJEbUhfh6CEq/wLEiW
qlLuUIAoEp1QZEvwQEhBx/1hmfW6e9te4motJk7s1iuVlximAYpiany2h5hFUoVL
0D9Ivo/T4YsfAMUX8p9OELwcM9d1ajIaY16WqpGl/l4MTc6PGARa0rn8F/nP2/54
RoYEzWBCJQoeNYYxTkbsPuqJtfPhlMgjHcBhvlKYGoNDr3EUJnS/Vgy6anX/VANK
uZ5KHM2KPjrZTxALXfzuBijuNiwyb5EuxfVM3Bla3GpGeUBMSpDZ8esBy1fEjGiZ
d3bZHdIt7YlCvsULTYI6gaeX95D8fFezbCSHynHzkWSjJ7IcW1fzK23pRW7LtAPM
ggqjixixfFIxilfLm/S0V9/UEFhlNc7bdhYSxIfq7HKBsFVeWRhGahRIhXKQpVHx
fsemwM606bP840ov+LvCkdqwj9JxFpnpcZxls8orGMpBFe643yzG4zpBJHKB5lvg
Du8tQqiaIkA57sP4YFkInAWIW8O0u5/n73DCWSi5cr/GHwX4Sg8NElyjrpGKRt0I
C+KS+o6mWLinAjZ+ONjZx9ap/9tJVjoBI1+w5CzVNGbatSyVBdJYEtjR8RYeNy81
N9FGQ1wQZV/J0B4lnHln+eMlkNjjcs5ZRpsNtYHXvCKM522xYVQbHF7vsNVKeLCl
tVZiCpe0trTjWxeIxEgGePtAvbNbPVnmcvkryy5V7Otk2oU2YIvXJcb0nXLe/DIJ
Jrc5/9JApo7bEPLNySXnL9dkif+35ukm2jQMVLvVJXGksHC0sBiTnId7pXZb92Hg
K1ckhYc5CBgXsMwlQRezvQvc37E7ukFHrRtEvCzfo7OQ0OKKvVTckR1cK3IU2XMt
EK2U2Zi3Jczh8emtyXLXeJrBRJ8WxLTL9g5ugO9KwDjVulVMDjokCNI+a3UNjD8U
dYIfDYYbuFHD3zgT5jPbfiuK/Jq0hPnjfuJm1qOa3Lk54jBWKpvEnIKKxjbwyJcd
WeaCEZzEVTALx3C3XhO3jH7ah8bRpf8Lcr88iu20v8tP6IMctufKbpuu/KJd+fr8
gbh4Se1hxipIBT313U234FOPq9G/XKK3qRKw42EJbsp1SyviuCHmpzXAfdiMevGf
nsbNTcnvaN+c052YqnzUgd2/PzFOsnQNXDPcpnhh0XUIJmLh6BhlShVPpI15WcIR
n6BVg+9UCN9Z+cZfNQstZfeNOWiSr6PAfG2RSQ+8C0u6wnS6WEulpilCh7teNuLj
U6F6gdz5zRVejdPeOzSemQqNBYZWbhvj8mF15fhkP6BxhxGZBH6eDF1WKo/UCVwV
OuAeaIUN3+tTqdBzmd+9lD9deFH38fnPw9KIxKUwdl0O660bf6MQhRVXn0PlpXoW
p0Hu6/EA4fb4gsgFlttXm/Hp9ysE+tAR/KHcbDI7q0WSWyP2ocA5IulkZbF0Hphr
ym4t5qIarBQJIf26c0jdNVeVm/OP5QHYvWKV61MnLbD2YPV7eC+fxIotv05Eexgq
vFqEM3oVecrWYOmknlcefInJYzz+Vn1+kUivsnLURjwVez7QSwRSzw0e3fQICY4N
yTOvQyluLrh47gN87QEkWHvHerO95fMzIqUIPcYw6F1FcpnMTifFcBEPEu7uj7FV
o8Y4RXojyl1FKs0SqY/XIuviXfs+ZT23TUnRTktW/zVeOjbUmfU8ph+pynxIgZPA
j/Hd3J/gtihgKzw3s2oEbclU+1ESx+Mx9ap/uqq6/MO0iKqbhmEa4mXeL2CWGCE6
aS5q/UzqeamfMdFBxs1UcL08uJx1yWC4b4kYLMud/0pSQQkvrqzvN+cJhi4dlhdS
Hje48y2cVSf4Ja3MZDtTbsE4H5N8i+nnIMKW1o0d6CwGl1joJRXzoStEW6gJXZzD
k4jhy0mRIX7dNIAyItKOJpMbA9i5XdGLvw5hI1Dvx1easgx5hhv6GKpjnfrS+a9X
4dC2e7k+qwDhFI3Zmahy+xkvQzfg694qSwx3+w5uBHTn+WrpAgFlYAqX9+Zal3rj
bvIIvsEgf7q/WW6tUJHA7pSmnmL0qFWgwbOImosQ3OQi8jqqndxkTPhoLTJ5nHYC
dH6OFxS2k58Wddu1DLXm4spcjiQ+tV9fS0vkGd/8JgAzsMwJeSkuGkYtY1lHKsZw
UBcJc7kDinHEPAMLeZfU6wKWl12WvAOVP+XTMy7Z0bkvZ5isxO+Xrg+B42yT7OPB
23B1T11c3qcO1lOzRSv3O9NKhpxnNyoDlHSCyS6N274H8liIPbgQCC02KP3dpMil
wyZkkdDx3kzFrDXL+jFM7H2lxKVfIbhCkzeN4B1ZFVQkv0JX1wfrg6/iI5R1SIw4
dPK61zdIxAps0yp8S5a+lB9XYs2nkr/UHTkpoUNZfsIgTjtZrIArTsW6TRWDkNZn
61TpyBCxuu0oXA4WHbdYp56WD+Dceo/plrruh8EIuPVemdCYEQnuRmpZw8+zKUFu
DHKur1zqwxoIE364GNEIisvSZuZ4G+LSd8zC44Ckja2a2eG1rMwcSk/6TyhDbOcG
3N9Hq9WqOwmuViicsB3AxHuyShe7SA5gfJsRCCdVmi14soYvmLNWXr9nuZOqwuon
N7IXVnUZNZ8v8zmRWf+TraAxhaoJhsS4pwLjvKqE3e2L6DykcSEgkq+HK1SmPtro
dkXaPrM+zgGG8m5HBwfSB1qCETHKzT79Kg+qEodGt4cqAkCTLgHLn+3pSGLWQcnc
U6yFopv144T1Elp8r1x4GjWVq834zT3gnNsiNdVzU6jN7bQGKZb2QSAw4JnihBuQ
meGVCvdSPk74t7k4UPZTNzKNItiQdjxtZ6hm2vUawtCGpj87oBAFbDl4oePyVz1w
pmvWdeBhamaBY5Nx8AsbaTJy0GaF35HdKeVf/KI0D0MxFm0idgfT9geOGZxWceKI
shjE1CN6n3F3kHnzcb1BgNM9hK09DJTMACKTLwp4XJGkJWtMBfeeEXK0hXkfqJ6Z
PMaXg28C8U2eForLQbMJQZCA7n1K38ZzmIqY1Dznqj6E81rnB0aOpOnUTzSVODMB
LvWbfhCl2hkpbESPUFevE5USpd51B9WOinCrKqdz2peYsc/N8iWzkOxHWsZtPBt/
tjhbw+wDDf+CYtyMasFe7e/1EX7fQOeZAuDGKsNeVnEDsOHx23K3qp9qfOEZMT0/
p1aROrPWViBTaYWk5J1oY2oRjukQGHC3pE63dgKLr5ncxaINDMhYfLyA7e9Zz58q
LG8+G4MT9yXoFhjrYF2QGVEBoy4JnTc2F989W2xHf2haKV0/0IVGdrqn7FQQ8Lwy
NSKVhCHPMIDNGTTJKoDS5mxn+GiIuKyDIunWbcOVM0QWQHgTpgpXruUOZcVjepA0
9qurMlil/Ow6pzV07NMdKQBbc6qBC7HMsBOxJ1CcqXPfI1jZnZYBX2Zy18ajST9s
4pZUCHIuX+j9Db4QeHFAOeWcB8+17AKFykLEB7lqozQJVuFkYilHCYq+BLQ2w80B
UIB8JqyBCcqMEqZrtOPD3h/yq48Vyth/7/w3D++cmdVD0CchJdQu6i+8Qr721g8V
nZ4ZxSrwsQxkUwOGi1HAJPgCWeUriJV+12NPlRWnwqkiSt0bAIxX5FZ+KI+kB8MA
8DqlQEOooo5hwZ4oat3mdevtgU/rnD8JSBt8C3YRmw6+jTl1+8XL4MmPDatM0YtQ
4qTJPDOc+aY5X24K7gKfkr9H86NI7nH/rtiuBV0VFXS0QPTKgHfsLIV87Yab+cIp
p0ump0MGaR7FrT+KXuiVyqtpnyOl91SaG/nJhNzJ/txVGOU3UMImtsIo8eDcp2zT
TEXiNrrVT+sFmlKJCVe83nuu44mRaA6lFLay1q10iA58TxC8xZLcNZlyLL+oh8Mr
TbbrowWRWPzNJJ0/JqIylscl3nuIt6qaY6sz8To+jRZA+NeLAuiJCE81KSCnWdXQ
WoeWgVCTbcMYaES5k2FDM/Bg8iBYtTvD+mWh3cKNbCeriBdxAafqpE+ZRQK9O6Dz
FDgI70meVYFCIyoevpwLWJFow8WAwxoNCfRs/MT1S+5/4wlWOqKDkE1pBd8Wbgcn
r8xjJaZBWbksMIKKG1+qldx2zGPXPtO+7OZ5uOikYOlQ3a0xFnfkY77yZS49CiCl
dObz7dgBby0VDSmP2C8sEWXLnNs2vv/1xVYvWj/OJ/eTweHCQPPc0n8E5eXOVBVd
F4bl0VSaGZZMcypvqJQDZfS6i+koa2CxOOGRN47HyragDq4Aotk5Y6MDAJx/Mp96
30diENQwesRxsta6+wcWuP8BaHbc/DYuOpdLUW92u4V3ybSqIz9ivUwFpcGhjF8B
SLTaGLL5uJOWinK92bajvgNiBybwsHgVoVR0iU/ILzAoFFs0EIXmGF5Ys6tlG8nt
pQt3CEspMRQFqL7zYdH0GK8B6bfyLyHksl1P81Mg9kpapwbooG3hmrJFgqr2OUtB
YJaatHEhUTIbqgnLlqet/KLxlUSwXNDTj0gLrWPWhedNK9Oq5likI83MMlCeUG1V
ChkpIqSsRNIB/YgMG5J+lgfoY0lwTV8kXQfdg7nqWc/ppeVW2EW9yaZEyCWQGFHN
0Cd+TgZxU1Rza/DrBBt5Y1RdK3x8onstM4yQLIx74UmbNyAMknqr/BddhrPuojIZ
Xn1fhIOSowoJo+tYKuEPyP5t7Pj4mQRsQd3IS33UgejFstZiaVelt/9Z0k+aMZ0h
3FA10HkzBDcbTntyc5ozktavcq5KnnsWFKWN5Z6EUt9wP6dIhnZA89kkrbRWqpCk
WKCUn3Yjq0Gke3Wy0zDYVghL7ATB7sbBK7w1ZYOejcmRUMTjbxkNhpPd9ECxGc8t
k6ytOTUK20vAjim+kzy/9hUsjVfrC0fzu8cL5BOX2piCtAR/wlfEwyJyiUOqNVED
wmynDt+UUZVGm9M6XA8X/Mw53Vyhv2VzSXAaxvnuEbhsJZo/KLLGimZ1wvNmHV2K
79coVyP8MdbqAvnEiyDC7VQomdDQ0D9fDKEmRsIHPnHki+BsyCZSAziIRqxeZ1bk
tIzP3JUnEwOX7g5WRqsfymH0cSauYxU5h0LcCFT8WoawO4EDLLTxwQcpKldi91jC
21lc372Eg5IMEleN9FoVYw1LpY6U6WGdc5PTrTMs0/x1fc64Rma/SanO2g0Xc78m
LeeyeID9saOEBlAWXH8mlxeKpGMg1oa9KkhlRgS/PQp2g5LlawKCUW2poCW124HW
Z81oT5YcVI5qMGQC2axvowC4aoEF4olPD9GGgj/PNqeLJwIKzBr1n71381VF9n0L
5EAe5Hd+1RyYkscZgYS9MN3dT25FewkdxO/0aG9bSUnj/QoiFnsR6G480m1gKV/y
Aoc+sVL/R2lWvL8m0crV3M8V9HNMMuIkZnYPoOWRpKwuYMAYQy70YtChhJRD3A+l
mCgqapxvq7FjtflizlVegCbaIc3gRyt03nJWSta0b9fmSzIIwp/xg9KC9eWBB5QS
7mF0MfEm56hapwo7N0/YIAxli6/V9+7tJvohjd9/S9G06ziGF8xI8hA2ACEjapCw
wCI/Nhg0SJts+XliKec4lhjigpRo9XSgPNEGzJxVh9YfC1VAW9VLNPQWUFb75QHX
PJLbU1l5mp44G6ZlB1VTvyph+r9uq63Mlgu5PBcYp2ZZ3fap/Hhd5IZgNsA51Xjn
Qyvqc4C4MPz6Pu5lImwIatV6YPR2lOSfQZLrQHjtFnuYr1sjdT6LVeml+MJpHZJC
MT9TvWKNvo7OrjyloK6LI81j5hu9C4o22qyAuGsIfy743h3/zX7rD6NVOc4QwZAI
ptRxGsQCKnC8pfyeQUWMy2OXTmcsbPDPQ8fwfj4S7qjqLJR6XPc8Oma+SxREsTYY
t8EjVUBOsbvCiCPBpgRzKaKABx0D5GrAEnFuwkK7k9KaHaegkEoXgUKp9PZi4mkV
m7qidVj/eDugi1Sd79IXGP8izoxgoV9598sM5AdBFzgXy/gMEv/JQdEnx4i/7/Jl
CmCyrgSjNubb2jVTBp2MsH4LEsygre4RsUQPOF+Betm4JXXYEfVbr5KY+fbjtC2a
UmhtYuKQ1AI7mcvdx9kkXddKGo9Ngvub/KPH5NTRlBMvVjWMkbajkuLrBPuHQKyP
H7qVOzeMlzjseJy6m4kZv2zBGf172+bDdBY40cvS1wbtFprR9JXAdXcNOpnj9euA
gSeCB2QT4UTZwkGNqtXPBYcMVaFco+QMQoGLPelA2ofqMPAc54gFaUDQ8nbzDHVw
n/p69HQCdQI1sJ/+eMJrPw3v7j/uXrcE39x6yPIT55FBKpfnNiKomAhu2NkTRvfi
fW6mnfLhoKTRL1LqKMch2jt0qTJl8Q87yDiveqkzCA8+8Tztd+B9RW6YfPgSD5iq
H+UBQz15GeXCCIF1UoGGUOh8qm88sFWAR2Zv5DJfKHxesp7Ira7IZ7n/OFjaq0CH
0fyH02Zpy1s7snLTjtfPtL/1syn7avNknMV1zVAQf5dL5nTxwX9RCEA5ht8HkwlW
XBLpZPDipHQOUYx+cth/7EfYsVjxwCJ3R7a4dOlG3gZdOaP3+LFtxh3jhlF6Utth
i+Jup5nE0OFSeZcT3fLW0HbimaJSTfofIrthzrgo0akJMydVFCTDhgXC7QibpiiJ
ODv1174sVjbt/CQpUAkfaab5RoDm0q7JZ9b6jafGa8FsR63INiTQJsxFHsyyes4u
/I7rvCgXpVs86nhAZnyswbu7rwfyqAJsch0E3lHF+HbP4atgojwYCj6ac06rXI7M
BveqtRigiae3KsHQamG1UgFfW8JMoKEmxY+X+va3TJKisPJh/nouxGG0y+vtA/z8
FftehGyxB+KUWWi77A8zbQH2LuEXq4Icrm7qj32+9NlfAF5ganngEY3trMJRfZ54
aEclFL7cu5LUFHOrvZB7iMPAksIRpm0mgmbEireOZqBLGaEqgQQY5okQtvXtxo6v
ZdaeNkEltkIUVah4mGV7Co1aWmvsxfEr1X7eLo85Qdr3+kAs+9e+lXSuiuJwcn02
e1gj+8xxEduoj5VEy/nUx0/mJcgH3V/dkCdq51WRLQfOrdQZ2iE5+0LXvnDHsG0h
5xNqZVzdNk+Rr9PXAjY4Wcd2F004eLSL4QN89foCTXTKi3HxAcqrdEp891CTn5rG
4OZ3xlETUZxuxGUPKO8/5ugfFkope3Qvq2AsqGQyJJ2X3d3bl7eRi1T4SegPAOkt
92G0kHlBAu2e5cOeGrRsilut0yoD6TBG4LvG//5xyRFA83Su8ORnvqnvrFePd5+/
G9kWsFPtpmDY2WPPCoB+Ul6vrq6uEI11Ije5Kmg/g2RiEBqJ3YP82i8GQ84f7NlM
lZU/TXUp/HY+f5Q04PhUh+VPBlVhGWDDqREvm/QDexZBOJz0mVGEXfFMT6/zx4nc
yukmteUXJclG2oyx1nIdR3pteT6MwfIqA4hQ8T3wfOj/ZS00R1TqvX3Z1eCoEwzM
wNFErUNAAFE6c9ZTOvpNI3f1d21fS4hBw7pVqdw38w2y4CB+ewf855e4wrVCeVCg
pDIkzbMEBwqo4vbGqkCiJOhNh8tpMpyKaXVezXierQL6vRIgcjsYfopCIzylUAqH
SfQ9urqGQ99bnuOjz3U8LGSTZda7cz99wTa1x+GlzgamhnGVCBRecqaakbavEcVy
X8ZhEXi3Y/jGWg3YXvvkJ3YhsIUdwUh4/Hx4ifeGLDbKr/2aA1MlHhTiupzi41Rj
nvYvp5a4YA9JU3wolW108taFyZgU6nl7Li21tV+ORIH6NsGyChpkoReqQO/nPtwg
JJpgHYJZiZ2MFZ6lBcMQuTC9xwyTuP6xcLPrSvIUNDogpEuIgw7RTPSPIcTQjUdZ
mmLp1puevsWdNfVt76LpIfz72nx2Hz4uz/x12DqV5lwHenNVIBpyo2Sn5hDqPSQr
XViV4jrhsKOe1SKXg5Iy11JxbjYv85wrCEn+S6VRTXpIw5IOvK+Sc2uoUImUA5sQ
CLPXjZQVYdUMOpEmAnG7TApZR3bhZ4cRhGaalJ1yTG0wmz01pzPuvG48i9P1sl1S
vd6yC7WzmaU2k9CdIXX6meGf5PmdaHc/gnzTJHWBGh/AD50+/aKkJ+gQfIjdT5xZ
ydqnhz1qCQjZAiAe7hCUk1/vNwifUyo6GqxEwiYfYn/MoEcTjAMWhhoEVMTZoTkp
xBbj4d/D+J1PKJAc7Hi2EY8ziAqgFGeTE/HjsVuiFTwSBtqM4PfvTdA/1b5cZgJ9
83TCEjN8ZpWjcOmVxxjPaGFMNL2w9qfqBXh4mUESB85Cg4OLXSPxVLcZrJMYmYsZ
CWYxuOQ8Iv4XFI93nEYLwFvKUkxuKCoJwBWtPOXQS9zJkAWX25ApQcgBR2tMQ1ph
j7ljcXbd76ii1RD5BjwFEe4LsNFuLHDdaXutQDUdpf2FFfhWU4SvujKiOgIKhvTH
0LtdC1I5K59XfI2/0/posZGauQ3pIizjjFtvHyPTs8hVEd3X7f968X0GjwJ86rWd
RL25sttOQK4yoKglA0XQgYzRgWagu26lE/4+HmJXLRWP5tXnb6xj8NLiPVzl7Xkb
S8n1xyL6gNQ6t7bia4dQJNcen81kct5/16I5CC55Uoco7A2UdlpH3dryAyxDBx6F
vjTJZxK0ColLqvS2c7lEpyDUnkwM8l5jnJLEgvM7vw2EyMNwkZPDIFkbBv9okWUi
orROXuzvkYX1h0A3JatpAngJJBdc72w02Htg0GLkUeeTluChA97i5nsUfD6j7Rj0
XJYaqlfXLHI/Uv4i+qinREwd/nAlgbI7WKba+67pvX9uuAOY8v4y+X+J9uSCbiQk
/AH0mL4lx7t4vJEQUvZ4NdJ1XfVklfqM0r6jcJYTjA9wyDSAspVQ68oDjJ6NU4z5
Hcmx/3khlXq3a37IJMF/rK56RLcbtTVmoLVklVSM84eg1frMuoDwDcfO8yJf2xjO
1xGYcn+agSw1TDzuZ32NB2a5865RdSD7t/0qlFkCbWfABOGl62lX+vbQ3P9v5578
cleV+VBNwplnw54lBbO+VF1ZYP4xW4d2BPkokoXP7XDtJ0XCO63IssRWAP+2hUgH
VYxT463X1m8ZbNZC8Kt/CBdydN4gjxL9Ns2HBaT3n7WfOYookNsrBY6tK0IKz7B5
/ZAR+NFpTKguu0IPLwJLCYFp31pD5VvIN2KDPf5hVrVc+gYqUtfMp6SyjqZU+SW9
IGkBWFkY53xzwdRWL4EAoJ0NLMlFE+7tTblvvKGXpO3v+kjzO6vigTG1hborgOQl
monFYdX0y3sT7F5eV5wJBX9raLD1DJNyO553KiZ/9jbJzP2dzVLMlsM90ys9Y3Vg
AMiKDTI0xVbFBrqCco31DHWHBkDTZn2UT+x98hHV2JAr01dFqJKRpNhPSxAVvk9Q
azEexLHebrRpWxpXqA2gHK52BA7LUFtktsc4PJmySjRBRU82hOTLm50jZf58AaRP
NMraU9+iL2zWDfgeu7h77ybZdUUMCjrCspbaG4iAnXnxslBezyqaBHOxoKc4mW0C
DXlFMLxT63WLINmB4P6tnXRxdvykq5hehfYODnOX8A14pXVH+XtUXTEZwyb3QnGK
A9uGJADnsN56zGJ5DdSJqDIvcGmSF2z6oQRG4bvhCArbGTq+oT8oXfFBkROu3bCX
BDlI5MjK5XiRtEFRAztLf/KAAqE8AplZSCZbiRH2Z6Pf9HIJEO5YyXUxLhHw5+di
FXjhwb462//9y/a/c4O7az5E1KYK8I2GiQ9J5Kv7v8Xz1+HywcaHCWG+V4do70mo
aBN+dvg+ldYM6UkFfkSrYndgFVfW44tUKE0TI3mp2zxjmVJh/zbnMh8HvU82dxzI
fhpEFmDr0s5loNkAa7oaGCXrXE+xQy83HjyqhnXwdmpRcUwihTMh9ZoBCgcCqeK1
nucBch3ReaJiHehyW5e4/T3NeDL78RE5rYJWIxPr6THkSND3lMYVJhzdNqUxCmD9
HexdpywqWZOPcMTI+1CKNwqddD+8GqWT6s0FvBQDLDk5j6Q/Ot2/yP+mLtRcYXyZ
TrkBTerXrmzxKLSwquAaqrWb71s+E3soSCI9aN+PMeY3lbeNKA5LBZ30pWD9j0Aw
wLtgGoEdn8zLqTyDE2huEjWPrzX8Ep1zR+110flbvqI4AX23SRTKyhWGbHM7WXma
z39BwXJd7JgsRbQQrsV5IreoIFicg+tm4KVpmRhDHZ1EFMM090igE+vIVa9Sr8BY
sQDa+7gQAyw1ReOt6wPHBwMUMGqzkZHaT0kFSgSF59UqNjJmLk1g/h0AzR2YDhlU
/9BCP9rO/5hkCQXgoaa/FopbCnQL+6y646TJsmIAcrakVP9NnNYexM/PijtLRohu
SpkEqhXhtLDL73BD1QQz6JdsNGbSLylBYynDevJd7GabeA6izJtr62bBlogTAljO
IIViN2UDu3SHLMUAaRN9Wmj5EKD2AFdJCBkPMnTu/8Tn3XBCUmiwZG1Na9Rz+If4
hteSfL3YiywgFc2W6QGgjTrCL/Zh3f4pCNxT/HZFjXFFkFj46kYsVSPJwCu7KFAx
XHGiMa8Tc4hFj9ZQVxadNi6D2pMHoiyrMcMM0/98Yh5oJN4ywouOSl2ZbaoujMg5
7uLHDfaXdFsdBgPfVgSlafYAvUzYY0xMpT2wtxnfHVwvYibyri32jK7meKLAvdOC
Qoe3413QeC1B5I/9/HO5Si1kVHORbySA0nrOIAErk9G9ypccqvfE+HwE6NBhGHlR
ZTIKy0gT/t5cBgpHgVj87Al5QSMkU1u+DTHkIOo5dapiOPYZ0XDdTuexV6LOZRD1
r+imPjtdqSdtCR22tIYwHv3qJQ9H3vcTPRw8c2xDwhCyukYWbDNw/baEUvxRIULk
aK2KLiYDyszAdZe1J6ajg67GMJ+o6ltkULcG1QdFf6a4+lR9bFiSBeZ75I/9eTaG
jO26LWtbstcJaeMlxsY67XVQV6hAaicfHTzvwC1Q1iIMn7UfDlhiBeoW7/b7XreH
O/ylJ3hCqlJV5bfyAFDdDAWlD3BeWcrbwcyFK6ibbWWdY5W99tYhRCfczvKIto2n
j4e9FqsjtFEhX4y2UsuahTqE3dXdwI8J7pAiluLrCEyLvsQGmqHr2yfBQYqc26c9
p7jTjlIH6ryshRylfyK4QsVHhz1jR81yFXnYMIua7mt18/CKl0kZrNKMPFd3wcTq
lUC13tSJFJwExUZT4XjdlTjUFerBMP2RNQmciOAoquVzuPxmQ4jj3tELTjlwgdOa
35FU22xDQcAJhR0z1I2yhNVtIKCbND8dX/CC0DZJDxHgpm+dKqZQvXXBSsahkReE
qugRIYOoTmJcQGlUQDcGucfEEMclB7+hR8YmAM8o6TxZPTvMYIFa/lUkuos6+hez
6J1fHBk45Wxg0Bmva/SKdjncUU+typilCu+R0ladzKOXUj/w4YwAJBRe8vl+VF3h
EkY31YRvwflLk5fai2rXGwgafxguhWgECDZaITanjbYb1IlgcG32njzbhKFJU6Pn
e7Khm/BUQqRZsk7cs4zWsewtWIaq0luQoYQPuMfgxACDapbZddD0OlHKy8Nr0QOL
BC3jLxB8ar0Ddvg7welhnJqD/6+z3jGoZNpeGvqCjEW5mhYV6hLXGa4gkKRbUU1P
BBEqzAtaUAmv4mdgHXbD+315tLugolASMWmctcZI2jBTQHUsShOSCeYqq6vxKcMG
3sUF/dMXGieV93jb07ZcolHfm8R9gMxX0XXfY78IHgVSJwtyvzAUQljzhnM/TkZ1
JG+wyzngDAgVOl2R8uA8PacE+g205jV/5GqXhYQFham8j4cVZlvKT3DHMBb0zjaS
T0CV17Lx5CYS5xkviPisbqAJrjPX+dRzmv68kiuS5bBWgCr95Kc+qSjEs4w0F4I7
Zx58J6MGIap/rNgKzsDYzcHN3ClQkQVpvs7MWnSTAQETI7lQwtDISMEHN6Qyawzz
Aac6wiNbTEzOi9D8jKafc/6n+JFE9Rcu2qWj1QVxdn/xzDfour/GmxrIiUO5LrUz
Jb1HrS3I6ZtzJpKo3gtrJ+m/T5gpRoEd/HUr+n6nwdP+mm6ko2UQuIxfwqruWgS4
nX1FRW2Z06z0DUMDZOmI1RBBlMfu3/eN2AbGpodwc6+uh8IcUycdHhl302o5eX+c
E6FsPN8BtIS/AqJ7Q8fBLVg+5znz85zRdnYr9zjOlLBswbSCjxI3Qk78WuFwDikX
L1PZYIRw/2Fo4uTBfk7fgjBncVNZCTdtGZ9BWJxcwUjzZeS2gWveRHL73BcUa2Sn
DHYiFtt3gZ9UlU45a3oyqd8HIv3N4jQc4XzPL1a8Crya9PpW460kCXq8HpK4miEx
UO5ffGKm/rPW3dAiI4AYtC5+wIni76EAVbSvUtCQuufQuxnjI4PJGetdLwf4/p7P
sLCtHpJXgIh+UTC9wsgHhNlMbwLRQNc6KNlaKmpWNTc8Y7alLOFnPPQau802QibB
kyZMC8r3b6sJizkIEIrZ0UN39/oR88LNAKXO5WwhFZbuLA4R7PG5IC37wRANksfD
46Z1WtJw/rDkyr2tLL8w+MrKJ+YarNFLmP98pWUt0+yG71bWwr9wR/sWVG99SlqB
cvo0HEQo+oDRIJMDDB8TvaHTofSI6RpEq+PVzLUpza95aqRU3+TraPTURrB3VdQI
ta0IaPVu+Va9GaLX2V4lTJ7/6e07+PlbZAEjx/YLIIAm1PAit4IcIbMMFH9Boi0F
vowCL9NLjU/0fCus+ITAUrw4x29evs/0DWIEhH0klkCdvXlBNtf5nbovunaDDGcj
BlL8l0H0vk2DeC4q9+xX1aN1sZo8SQLKMdbvdKq1fNlu2bfhgxgSNISfNIYcxdpt
ESQvTqmRSwowbFMDV8n7LsQWxq8CFfUworI/4EKRLXUK+v5Tnaew1wBT9zH+ZZNE
puC/8ByEW71rgblX4ZHz5n3JKjcViUqRnK//9vnzXB+Mqj7gOn7HIzH8DkSEjKgN
bVl60A1iwE4Xdp247UM+uzEjxIF8c9HbN6PoIBYfWwiRUDfaG94PrNkWg6UZDh78
WWml29RM7KWkvmU3xj8mS7qIOt5ohJhqZ3VdfgoAqLLpEYIuOFbB0eiT1ddxtKTz
jHJqlK2dariwEqvNtLBbH9l5iS2hlRofo7YsJoxJkuXuuhpRYdjMAxNDCdpR3Qur
e4fMNWAA4yp+AbxCXmo6pem+XacUMGpkabnU2kszIXo4RynimgeqNUNJOBhKxM0E
1aPRLul4xpf+sCUSpV77Uw3U+0WcyvSOmNRsXrxis7g58DnCZhmOM7I0sIQ1OSxz
5qC4Ph1jXi8hYQk3U340i4q6oNYxcVm2b8AKWB92+Fv+ig34zeF3xwtvz3dOyf+s
T0yzYBu0MSlpkUM8QOD2Q7jKaauWELQmZcpAnIrFeS+VIll884mLMHJp4wiqrIUF
HnERQ9zjkbmBTc1uNBHIihLG9mlUFolAiRRw4soeBle0j5eT7KqJ3CTis0USL89+
HaVcQUQTwYoWcdiAebRc6MX/AryVQ5eq3qFOi3a+Rc5rqb15zs2IptJuCuQLVxvw
lLA2XNkX6ZFQtXDQNjTLRfR/Me0JqtO2+vo8zazjWm2Cklp02mMcAIaKRzedhTV+
bVitrDk/Yka2ODQ7bybbQ3cPdcoafnSbwBjvaDxaNe2fv3Onj9Ru5s5OV6J4BmKq
5EqxqYIdB0H/0gqNztJasg0V69/+aNgGjC2mCl81yUf9R6W9xmmfDAxZcj6P2l5s
eLQCcRbisKisqQPHevCJxq9cfhoZrnAvFVqb8opgkgHywVEaeisjJaHGIzYRV+cX
T3P6skFKIMW//xBwchik72fdhibrAmxTSPGu1Xy4XaZkCFnGL+xZpUY62TitW4UP
luBmbN5NkvTrTC+rXexCnd6z3Mlo5IEfS+SN2AA/0bUa/dZrWMNzQXvEBYeylLVZ
QFiEW+kfh8w0y9C2lS72Xyfg+7rW/7z/Ob8Ctth5ayl5wN3t4/AfEzOjo8Avh9px
Ztd7U+p2qO+/oQksezkP06cquhYSWZuWVgTPO8NUAkeQCHjgIqrBbGwFYWj5XH4V
qPbpqbByhxOG/+Ui3ohdiX9Sgs2KbFxhvpyqzi0UBhM2vMD6Dn4zg92KSiUqZIjE
rnmVLeD7vEg/rNGMGe5Kt/MHzVIXfzx13204f4Kau/lcfCRCyLP3ySOtfZZIr2i1
vfR9ASMK5gSXCfKKKWWhtEOje7lozm2KRXcfBDYDRGCHkWqsiij5RNIrMoG1A7n0
9ICPQrcxXp6ZCGUqtz6EYCmONj58dm6pLj+0AT3Xkb5vnWP/kdr5KnwXsKGj9P/3
p27q+Kzv6QU3J3qr9Lmwt29Xpicu2Bef82LIXTXsCdD+K3ky9ffN70kNVqFf09ok
c/kz4fsL48DmY8hTymc93J4vpajAFM9B93K4mWkgmWy3msCjmXfGw+CKZfgtdr4S
0UOb5wm1I/sC/yrkuMkT7AXS6xavPOoFGpMk+y4hjFE4w9NsKGS/dd9RWZYtRAVC
HeSTvX3xLEF1RfYNiVWLzu/VgymDwPuQVx4QjEAaQlnNfmDo/rjK4LoasVuzSYy3
DQBTS7tgQxvH5IyKJP8WF8cFbiZwo2cx/bg5cSQ0CdQ2u6ndlsv2OW5XuTi4wthD
wwFD5tDv9mYnWWComaJnOiYX9J6AHFNIq1TaSqd0xjU5UHWDYfXs0oJi9QbtLXdn
a+bGGmhELkefq78mnjOG4Yl6gayBSipm+zjO4TASXAbpKGkXMxhAHvEw6Z+zwGA1
+rci1wB3WFvf/zb/hm6VWQXz84WzydCZL+OOOMx5OE2twgks+VJ5dt6sB3ZNj0W0
0etnP5IdqBC5LK0exdi/kHTiAITM80blTH9c4yiephFRHwsvBH5dbaFHeRIA2hAv
/mGSF2FXFA4QdWoWVf8RhT0bGwc4ydWN1j8D5iKTfjNUCbfQnw5M8fD0gqMUx3FC
70M+TSvQ5rbBU/GaHPDcFc7/DolbDD7ZDJNduQL6tn4dAvPtaShz2BFXnAXPopyL
rqCaSUJiwbTQIwtQoXeGrNpcSF70e0nsdAg/pZmslKtAt0zOudwttwpDpZyf8jct
EOWEBplwCMXbkyg+nlj1ddtfiDR6D1VHjTZDo7LyOH2VE8KJfajCDrMd4ZljiPsK
GY1XLoW9cC4MHWiSJsGADlj+eEWEvswUfjheng/oehDYkd5izEgXzsAr1KLM0DKu
CXZI1mFmXvW7oEclByVP2O2N+63ankQiWPIknNLPf0E5SfP9juytrfh4OcbAI1A1
1wxWgpHHpkq4AlXIR3xsh7kejOtj0sk199ozh9nqqXEyC8dQbGNea+lMW1DqjJgm
LDRalHchfUsnMmj+WiXATRA1QLi8A8vFKzrVU/jy98+aQ2frPajDb7wOfs5RFdee
EpVI1WCUaiXENn5Wt6HLJGJjYOB1kVJq4Ucq2UFe3cl1m+GT5dWDidffYHpD+Z87
ZVGAJpwTv06F1j+1G81GEaYWOMD+obTHtiV4mGSDqovg+TAPBL2b5l50HrSaUwBg
p9lANBGxWmk3ZTS8VxWcK4hvUiCWazp7a6qeCg3P0/bU3SH75MPE84nv5A9QtMRf
e8YUdmVuX5IkRrnQc6gfXvk/XecTaNtVLR+gHQDpIAmKakwtmUreXrzR0pdziAR8
jrWFgstj1aX/G1BFBfbg4KeNiV+0it3T1P3Xrn1Uct3J+FT5ogqVaBLujzZO22Zc
paB3fZHUPmm127dsSERECGWPiTd3X92zOdCJrfNXacuAeVSqsRbi04YZEenAY/0r
46wyd9ItWAV/UFKQW3NmpUK1OJsZuwEpZd7WtIOxd20SooEkjZXb8oM8ih0FlaL+
Cstf7Ynb+VXg3ulXxJevSE/gURLqCPgDgmZM91rKuTzlc1gnvOYH97t8Xc/uBHbT
7iJhI9WXFUXRVa4UETkD7DhO3yStTvhZIg0MG0oyMDMQKTT5AXSI+5UFQ5bAd3HN
1h8DzFxYtG5FN056/FvyN3gKFEqiwr0BgwqKUlCEDEZQGIhwandepqEG4XL0uNgq
rUvWmHx+Hddx7L1G3hZGt7/foFdpbxd+HfyQqWSIudOAWvWpBuSrVA5L+PKcLOi2
I/uWNntxUWzD5EkZGJJ5QacVHTHcX1kZsJdyc0rzEyZteDgWug+nnlyYOHGcTQ3P
uja1Qq4R5FGg5cfRINdaHuiIFLHAtOPi2BQETt2wrppBDxHmrCOF5JcerIwxwb/k
uRurzbBoq7YlpkHawGEGhGEhtDUJuO/tfxRioi5l0cbn+GSJKqb0M8TJU9nMX2TL
kodlv1Kxd3c2KHSpOTEzfgLyBbAjLpJQjVrA0zIJO8Kv2Np/61SKmFrIcJnTJZff
dX5E2RuZ5L6v22eGaSujTbqDYtqiev8CT8UAigdBawuCBNs32Id2lGiNeoz0V7cB
gnP5sv6XeFYvQDXw/rmlNPiXesp7xvvsCa6bePs82xRb7nC3w45PeySAvoEvzkwn
USa/S34oC9q96WwW9WRa7dRboawroqvduC+LIopoHcCAXzr7b1+W9a6CTZsq2WYn
wpAUJP1EGvIbDUMveJmmwWZYQuMu7Dtbo9gB2Dx/6VJ2nkkS2w+RLu2Pl3v+//em
NxvI+vAdBSmWOqXeQyZ2nH4ifI5+BZqfbZ8IKOkBDRxsqAlmw+LZj/pejiebALvd
piNg4+YByvn4y4zRZuUUkhEE0tkM7R46XcN+IYX5M41gSPUSu346ycb7+7fOfmbf
my0OKuWA+1tUsVwzOiCLzMKs/QAC0vtUfbNsR7i2804q63hHNnnyDT8zx/BPrB5J
S9HcfBudsp0K55zkO+1Vus3u40mSEfEdwt6xzlUdGZVK+hHAZqz/VL0urYGwVuql
+CEZ/m1fZx6QKYbkkKj+YAItBxiP5of/BEFnzxfgKZ1R4HSOUGWBhkp1YAeefnZS
gvfNrXYZ40grYrgalbjC1TFiKwqPm8+I+wsslPaCYOXlAY+A0ZfKnOOdDtrLsK6i
dIDZ/0WHugYLHNXp2LHvSs4nzOFoWiEU+vyjVSW4ucaK363w/dCzVN076UlBrVEE
UPEyRUs9W6Q0GaQ/8KeGFDQV+cbEK94I4dUo6QIBqO1SuuYcF2nYxQ0BzW1Oget+
00eHfFbHAQI+53CJupAjZhqaY0FrAmNuW2FwN51H/+BpD+QXy2I8a+1ZTvXwTaLB
WcTaQ+amybqtsb2KeNnZJKuQWcSXURZWyLEU33h9MGvggvsioVTdviX1uJeci74i
tUCPYWKzgFSMkUh73rjxeGpPhr4MJYPaF3I6UhjsBImxwr9RvgZr0CliZ8fmZU4W
E/cqzKleLsu+q2TSOKrhXgTPTwMTzNovBRal7ER5+Zpi9HPrF0SsP9yJ+7fZjV8/
VwvywR136Xd5c0T27+EPG7979NZzofrTP/jE1q1ysN3jxxbOAQELSz45NVCDlSkc
PeXNQgkdGTw49/F/Z0GzcQxhfSehfGJDL8/cSzbW/KhFxtGU2Y8xZgO9FCgp5X4u
IlxhZUfhi/ECooXNr6fjRW7CCcRLA8+pp3eRR3/5LnbxK53WGkRJLX4eet3tqobF
/5HdcNuHpfv50YiiTBtY10eoS8Ix2yYxSeEFlPN/BMuW/I6ellJ6FA5piUqwNZeT
3M4D2YYThAx9B9i8RvJKBCgQYHFJaQTv4U7NUdkb0JSpS/VzOX8SPtmCpUcOzSE5
sEs/dtTOwI9vuMSH5L2qj7rUDHOoV8Wh1o8pq+ijphGTtSR6DgNUPfhBbyJdKdZU
OZPvGc4lpffbvajhlgL+eYNV8NypTCMvV8/B2OU0zGecRwWIIEkk9u28uYylP/Io
SgnR1beOTDf3KTpOcKQvjP+9XnLWxVYzud+gwCc0g6HEpLoQEZBQWWWqoPyj/53v
CZ1WZzfJrf5aa9IlICDG0lQjPqpoLWoZCgRTU/rxuZo+srEpGJOC1X+KTk29sbDd
FSDhN6c+CQElZyOmP1Ca9veS1jYFAttI0nbEj91XF273oGnahdIbv581xXyDZ87s
lXik8+JDncEyXPZENvFdZI+DCKL4NwaJdNV71yR3E1ULBEsjuCUS4kmCdKkOuq4n
IgY7W2wu4CEbA/ep/YS0tAffy6fCgeLGYMWwxgJeUhegmjMB3ij0uYqZQJDjN5lt
lb4kqAShMpSaY4Zl2ZoS9yDj5qTQzCJJAXNMUKGRjCcMTczIjbKcI6iJuLjxGKVR
7181hC1NnrQU9NZU2q57MUYASN4YY4Ymb9aW2usl5Pl0RuQJGrE7L89DUrgdsFpq
VCLNPs05Wqch5mkX5hZgeKp80ZdIYH0oSx9gmNasq1GIn5Bj+Fsq9FnFCYpbyEbJ
OsACzKbIH1Ry3EE3YajioPRDUzzX5xkA+50PGWa4X4Ikp2JdX/kLzSpqOI818SFa
kOP8i79YNE73yXMG/PKfu6QqYFc1g5EmW7WyidS1j/urQmchBvG8FKngrk/DqiG7
0t3xVtF2cdny8Wq/89UDAtjarUVHGxbjIxfgvekiOB2mDP/jnZ2yQEHnlGgNphDm
eYNPKy0OfiurvNAMCLpK/kv43hT93nVyYfaEcmr4u4N9QEnacJ09FUj+A4KPbExb
GLJqCO5YmNWmAKVyeZlZDK03p2ep2AjLw5TGupTDAM3d+L68LwUVgoR+AQ39POwC
AaJz98pwPWVAk/0Wxd/AV7BM3gaBgJbvur8p522DZzzemhB5zAa+ujkB9OumqVM0
M7okOd9/MICrSs8/TjoX0+ot5UAxDlEJ5TVRwuorDcXHC8pc8oVHCA2Te3MHMw8W
fJy8uqeY7TlVC3qhjF7F5rOe0jiiIbhHIwpFRGv0C6YVCM3CK5waqmoPNozkLatL
fiRpG0BYcoU2ENo88igerx55np/A+2NEZpWZ2XTkZkzebq1W0Ze1Fl8lt+K2shki
blTjkKzD+ueWB8lw65Fb7LoMARl3MpoOtF658epO5mm2gndF9ZyCQBxiasLlUEgL
/gxmcDvIxwbaC5S5rjN9WY3+FIJPYOTAGswCU9ogBBIERe2rHge9QRYNh7p2qS94
KLTzi6ER6f5u4ECnuGMOmNaOSekt36obCwnBAgHHvu6hp9QFEToSI+AxKMw5kMP2
QjWnElhnpILR8M4u+Mg2dFfzU5d8rc1P7hT2fxzCwPy6sfO36bri5rWlC6dUAaSS
2y4beNJHsB41JfkUpESegc5oTHNcgUxfVjsP8CYldHlWiKrz+AlSNzDU8Ixrte6S
tLr4+Kpk+Nk4J62fOmxKi9Cf11XM4RA3xnUA5mxeLUpqJJVWqUp69Al7D8OZW3lB
6qLAhcIUNsCFvC3pLerjE2LE0hP4xnYxbvSnJUE/P6J3SpxiAD18npxMqh7sjgFd
ax/ysCOwH/E0RLgGQYvnZ2QrjnGVOuk0m1c1XAoFqUV37jkM6hUGlGWfBIHkFeWj
+f8aS/W5cYn00Wz25uK02CTZ5zRBH+peUgP6XOBH6RHw8whtuJ1dK9XwbinPPUyC
MmnGEYzWziKY+m5V+8+zDsuCNy1BKt2DQnPxaZQ2lwM8Yv4dOpE84gCJ88KkVPnM
D7NB5C0EcSRYwYOzjlg2T5O3klfSesDvrSuRWl6f/Qz2MFos9nkCgSMws/uJQ6wq
a4t1RYXe5LugfjRqtNuNe4H6xiP/jk9H3hyr1Cgvjy6uqiqwsNTg+Z5FwjHVdann
cPa5x02mhK3HpLeIJaNQDToNLylOScr5Y00jiDUZfLdtnzndUSrJPAW8bi/uEvPZ
kDcovGo+HRtOPjskSFHL0zPOh/FfVsWAN7LG68Dl8oma3+4eDhPuaegT4h/+2EpI
nXODYnlhC5GIcDkoxmtR0PS2PwUCeq/dB3iT2Inz2wbA5YVA+kDY0Yi0KuIYXghD
2MlZW/b+gRpbeHnyJCncKuDAT+9GcL9paFBEOUe+sg80rmCnbmft8G0MbH0luzwe
mkiKm6+vQuQxp53WRv+4HD8HHShr3wZRmDAHjqlFWe5aWV2wZ9fx8aYqYOgeZgEa
VW4LfVPWwcYRebMj42H+qHTyTJW0Xhy87AvxPzqJkKmwii7MkzUtZkf5pDBmnHwN
S6nabq1r+LMiEL16kSxMpmu6MerVbq431U43FyzOl+JHMyws1TyIAYSJE2c4jZMR
q4cKMk43Jy3OJze5aD6j2IhFAty8XKTPUPOhOqBIHjjI4BRBaXqjp3OfeeH7/cpK
mO8SdYWRBL1Rw8gvFctUMghvXz7UWa8pGzgU77NgRf5Y28MlPw7yU0eaJ3fSWmJe
QH3eJJOgj7upB6cQcVCBt+x9AGUUiCyvQAvr7XW08ATf0jblUp/QKeJptC2hhGAe
nTB7efOf7xqm2TCo5GqaFk5xwS1GcGS9oyM8qrydSQYcaCEM+MmU3wFHwD9gg1DJ
la3VAW2Xe44GtBfgY+FtY4GBLAoXIGF9R9MuNt5fh298FfXM3kr8HI79T73I/WqI
gI0jNVf9G+mXbKbyEZG6yyRBcYNG5rx1Dn4KpRrfF525iCWMw8OtsnWeIYvI5HGD
xJA7S7g7qxbP2fVejDp6qgGadbOAm0VJCZPbToUKCbtkc5RqQiAjpo5uBLN7fe8N
bCjSmUqlfNdxFGq+bOfG2CSY3Ja4B8sZdB5EAEc3YxyK+7zqMoA5GBzndYEiVnoW
E2nWC2aTZN6gTWEKQ07qt6EyYvgUId01/btsgpl2TBn5D74f1ee+ZxQbO6cg/fZb
5wqni2RNbr38XDw4dG+gHCmjVjnn96TUcBFh5PwL1YZL/f0trYSPOQnYt5w3aDdi
TUSWEAe9yFzWtN7kNlJmSK/kjueDfPHjvaWaaX/LBEO/u0nSf7Cq6tBXCjgE4Nra
HWs4RQWKbP0oPh0Ulla5uGk5yNARmd92TcpSQUVPTxSJkqkjy8sGQh51b+R+Ijm/
nZetVvrXX2DFot6a434aixFZILZ5YCUXtojwSVK3nL23VO1eq9x14SqIc44VyVvC
VZWU2ej/gS8HVHX/v6QBHPUzo/aZl0P0I4vYNobSy2dPoqqzs4eF2TBwPLL3Fln2
jpPr5TqVrD1cDr42r7i2YpFBcdY0bTavJTz+mAVWsCui+3Z/0cA8e6lDM5uH7dCS
czTn/X9MMnhmk2Py6QfC3ezvchYpi+49Ng0pt6oNF/KLlrTVpAfWwky0NtNBoGmZ
IeG9vtwKDrnIdbgnez+9JaaKs+dJh89ZGBFX2PCkefgSa7drnEy9GfgEqNVs0WiK
pgnRUoHwnRZ/m2j58EurampoOWV28KGHo7JxQGALBBDyKYlnyiLyI77olHjVPTcg
QKkuj07fcg2QVXwU+0aKg5+mgWmyor6PFj4R77CpqvsD0JofphsAYm97K8l7cNOC
2b21e/MWzfyoGGBok7QRMsNnq/CLITtmeHSrDcFlEIS2YOO0u/9KQhT1C2COHlYR
sQ2i+EGd9B0JDCDYT1FClrxcXOLoQpoNdQhvKb3exj1SoJg8mspSkzCTHRNS7xca
/BnaDv5LSU1fYlNYzRjGZ5Q7kMGY/7i3PBhe6BlA8TxDAaQzIIYMuH+ICvbCA5ZA
qyvcg12Xak3jbRSKuEPOpCsa7ETnpN+Lyou3RQsAtq47oKXL6oxILKxotB6QUXNj
CGzrvOGh0Z5jjXaVMhsPVNuT07AEV/hARk+Cy9rtO7o/dLpkcYldWtQGnxfmgix7
D6Rl5qqHJJnwQkXdOpBsyjyrRAmsfiExArA8sRhlV83WKvhhLi94IWvrRm3+qIC1
b7m171q5qBVFlHvKdE34DG8CY11AWkzGEjfHd5swQAdk2/bXEZhxpuIQf6pCCQkq
YE1yj4SaEavU9hvQa4q1/9P0cFDNZQubX1LIilQs3R/S43SjSCTyBGAtJv0sTLF3
yXZoZL4ny22kqZYOuS4b0Jmnsh5pdrm0DcmxtfMwLYrPWhD8vmuCRsqUGQhaxY4N
sMBGpx/oq8zGDf7geEgkdyLZFy3HLiZZdjokKTc9llhWczsjAxl8NDH/FAHlvRvn
khLxWEA/dWW/vhnG1QwQ4ODQFIl0Wm5l1yvVtMzk8igmdpfhrk2cUs+zc17wZv4/
PtwAkmjG+hD9S8uwNpLoDpCploWTlFddKzBzwN4deRHeUKeQijRhb8hmwbZuROh6
n382RP3NWgwFUoG53XIK0Oi6qpDzL9gP0507igMN29DM/cZpwi+I0Cm7HCqZnLlC
8DI2D+Tc3eqcA37fmbJKNrHtVxBmtRddHXvfqgxbaavRPKKaCF4WjgFGtwgeCdLt
6c8wcmoP3zzduVGQt9+pSlyDaQrLxZa8NHozwdSEGEePyo1+F6kdshFXlTS76Ph9
hrHB8rd+snMeWgv0LQ0thaGBiRApjtFovSDyrauo5S3TCXPf2E6+ZVz0bgW10E0C
lAZsUFb48yWutsQM2y/GKNjQVIl2JlUP37PWrI0wx7ohywkqh3nprd+MDnrrb6tV
sSnMBvT4sSb6qPBVrcqZzbN/CMFgLL6hafaQ1+2+Gx5/IL6GpLSCGgcpjk2oOrVo
sO4ylFI7mHOTgxwFk6rpdfUhNQTT67wouM6CaVxDTqnmzesZ2XuoxAfZRDGn74Pb
cKHm1mFDk5aD2/oqVoxI6n/ye6e5r4iA+TSEhtGlyrGt8Cbb92LqqT8lcDtYOtoy
9TNQ0nBx2BiC8EGzxPHCw0OkC55zlk+7sUvzvgPDQM/y18vDSpX+3ELtSdWrO8m4
mmrSkK33Ec8LA6bgtt2o2yrL2thYpfFIo5HaWPzQiih4GryBTXxrOOp8PjHDP2DA
OlYVJTOv3bRZldEDqpxAj4n9gFqg3hRsHPnvVzpUInViC8nHyyK5Rq4kDna09KRm
/fspkSYADKk+uefdMTrnvu00Y3/E0sy1WFEHJLqyp2Mp1Q2DS8ChtLDIZcDW+fY5
QabdMkWGk8dxaZOxgOdPcf7LBXqc4GXsFHTtPtaYMiD9s/ymAhyCBRwfL5OIEruH
qBhpp4Qdj6JEmY2lDpSdBKuDP+pgUekrFMl/1sGUEgaQPQrrz4Jb5a3NVZsmXGZI
x1KiR41jA0LOpee1EBA5ARf8rLqnLMwb7V1dOalPPGGOFAKE6aUxNK4++Rf9lBk1
MSX1geIzXwmcrhYHZegkkmQr4+Ix0rIytBUeo4MWH1C1ihal2rLUkn2PFAugZjbC
74tTMLHmZvobFZfGEyDuKtGsl/9k0bf7h795iWuda2kiDRDAQcisK4VYp+nmOvP0
iClUGSP48V099x0CQGwJNuDwJiX3LKewksVt3cvDe112ytjKqYgeFL8dWDNRAoXY
aphYwiQShFhKNehPQ9XL5o/XcRHEnYmyqAPs+Ark6Zf+JXgiBH4/ZGSntx82jf0T
xOi8Y60ItMGkxZLpNyw8uDhiGkPkyz/3LVCvktfYus3tFrIX1hrzj5Zryk5TP8ug
meUnC0nMTf8IRR8rA1b642Gell/BJKUgEPcsxsj+SAgaljfXsFJbb+GD9OqjGDqJ
lW7x0/yfDWy931mUuYbPJym1Lcyw0wQpJBoM3pby7NSsc5EFHcwBt1RT+kXpGjfT
t8N2ZQZzf/eHQgC3UGDPuF7uiU0fp4D4uG/CP8pUvOnXTmrnDENTDZGGj6uYrwFZ
h6VH8+IypoRD5GTamM/YPgduhubCvQ/1wXtTlLsiTtMfkc8PYnsxFIXTWIU90eaF
pJ3SgQdpatvx5wYZ5ZpTabTptb4AhW4+UjLBuzhWqf4K90P4y6dfljp2s9DVFR4A
7lSRmba02EXHhkHULLZq/72qZZlcY7GSumZsVo7lUCSMdgS584kJeaZJuJFMOjtw
jk6XWOUbYv53Rg7BZpHR77YlyReBgSvXzpMUWu87LhAA/3g6ydzZdXwGqVnKsUSX
6h0tkOGfIHkol02txxD86n3HwVDYeMCpHVQGhgLWQC89Xs8YYwL8s0dUW3leR4Bs
XWllkzQ+/03jGwbJMPA+GRo5FgTqwu3YwYRVoVW0j3Nf9UUd5QDiHI0Gk/5H4bTe
rcBSdRrGiLyi7HqQMR2z76RB8oLVtb5sckovwNdSNIr2uwKzQqovjKBufxH4p3kG
lN6ZlSVv9HrkpnoflEZvJbfwiKmQvDLVCzIF/CWl+x7yle4/iOjOzILnhyeu1P03
bCQXDtNBKvntRAxnmBJxAdnIREzGG169dmwLlgNEjuTAlj4kZQRGf9MMnDCrJFa0
hRGrYYXjFXIYOAd234FmHyg7yf5x0WkXb1b3JrU1bramGzE84IJn2l3p+gj65OWL
/xx32OLmoq/yYH1uMteQNKx06+pbPfO1ZiRnRF+WC7/FbImX1KawfpJxMcGQHmNP
t08Glxmp2yM5Kga1D9WAzJBp0NQ7abVK0E1fTFp5SdahLG6f7fUrkMb7w90RGQWi
iFzxQs0gZk8ek9PcfWzfyShJU4fQ6Ih4DohwMshAi+/nXv3TIQQcbzjHXktfNtV3
l59tM2SVG99xKv/pMVu6uKfghBxwygjany3W17gPwCf7ByR6yLcl8WzcpGOjh1EL
MxnaTq/O3HlEBy3BVPq2SX4v+aWUWjLfsrX17JVrR54HMooJq8UrZyb3GSPidMBz
HneWEeTNbBgA9NS2TfdXgEatvTJ1hcGVCq8er3AYd+Y6CGbigwNWa77G9aGYDmGl
Q9H80iNNbBr06U3s+a990HlodIg+SbS3ObiylY5dtrGtZBQn6MukfGs3mA/KwjAC
650ufFHs4tsVc0bfblxUTL6Btm5pEvRmi5VaUBvx79/J8TyP1S3+TSuRWAGNGf0m
gNyv1CjM5IFMbpEDddRoHnWKGtBtnDnWJGU4d80Cam8Y1zsePnA10NC3TjH7s/Jp
s4FMPOlDLrsP+TB+wlBNMkapBM3W3LWCzeeHlr39FyAGa7SSJO6Aju1LbsUHZgkm
QudWAbxbtjWQTTodCYrmQYcZZ02KdHdvCFkbwIjJ3Zq9s9bqd4ODxCusWwXaVH6G
6T7pjiOVHUlZTF/s5W5F840IwPBHC4ci6oJRGnzYevII70B2K6JyKaQoTeg/gV/p
hWHk3sVg0p4xeYhaGlnwOmMQ0atqkr04Oi1uMf5nGHpBU0PeMr2dlQ8fnUdTJlKy
i9Ug7XZMFxu5kxsvIH9A1PovUHBV3kRTWSm3K12cK8Mv8zUAnt5wnD9RXexbucpW
zaXY+TP+Z1w6yConJGV0Yj/pVcmnRPPIE5c3Rly71s4v0FxOYIt+W+ZhYtj5EMjn
cWI3xKpvL94I4AWH9NgRamRCIBp9ybGYufTUMhOcStKhduMkIkiCGwwHHsfr4pel
qDEcHUAoi/XjpJx76+KjeRSP0rhPDseFq1PfPD9qahUEsIlddB5uWDq4qq5vzFM1
tfU+VLUMCWUBmV0hWK2ljsT29tskG7oXy2S26mNjKXuDLBiCJzyoQeNqviGDj6Sv
BTs4lwhuPFW6UPSofz6vucf2jY/6BiqBKg4LOvuc13QxcRmD/xWMZENz3bD9+6mJ
RT0I4P5lUKPAlF7cAY6B/dOqR96brhN1xg31ytuycs0W7wUh6pX3G9M/7dV54OgY
drQxv7mCiEal73h7uichtFfll20x39CtPx5GHc8e7VkqKCl28V+L9nLQtTLoWXlL
0fEY4Oivw+iyKMcPZcDsQdq7MKoKszm05NEped0nHwHN3lKo8qPLKLHNF9dK6sfe
rdXxxVmeRnD9u+iUqTm8u6fyC2UhdPbUuFJ1RPwr1QpUjq6SroK283o9y6hCTb/E
0qwCzA5k/aKpcjh5M4FreiG39IChku/+2J7449K7/uZSYMzlCz09CnEf/Hzi+G44
+NRJox3IrFO9Ej8k6w46e/MhzLVMjrHJgfJGjVq1duKr9aNouKYv0xoNufxak9Id
S2GSYtNw2tkWBnadhQDnIc++vX1BGfl5SvhIkt+WpM83nk0WClJPQeMIwJLmjpv7
P2L6GC341oBNz4+Z1eDrxP03LN9hHGSJBghgmna4mR4DBR8DYQgFZAvf8LWrxuHz
Z+SAG6oBv1KvQVOP1pjvlpD3qZVS0Yc//290jVxXXZjS/5UxAasY1YHRMQIZVk1u
MyDN7rKun11gwFWktmkmGV0gxCaWyrABKGeU9Hd0IscINCNo2XRI8lAYwCJnrj2o
1amG4oWNVtjyuY233ajCPeoyURYryAsWbQt7ze6cVbg+oA8hFyRN3QzWGTp8GoHu
5e1aSFcgY2AMajRfAUdjTRKMod0l85F5wirMAUMI6j4dXkijr/jwrJ7dNuAKA1Lu
5JsLrEf+MMYFVAxQJnP1jt3cWfVGBAB5x4rp3s+gETI6rctQlXizN8/1BV2v0Y7y
HtEWDgNPidyd+btK08eBobSEcOnJXH+WFK6vZAvZcmEV7cSyjEDJUIz2Lq3VdiWC
u11/xnIR71sFD/KL6BpJE1O+Sqrf0FrLxq+oah+7ec8z1md7kC1chQg5ucmOXeO0
2m4kydasgU93MvJykSWhzex6kHyvKVtNvQxzUNvicYtLvNU1kUQiyRVCeYKlGPRZ
DDaNMpCvjw6kLIK7j8DKZm8O7P5Vw72VecIMShdRgMkGoPr3N7/45SgqwF5AK/xZ
T+si9J8mKqazmPoiXwJSDJoCBP1T3lM8fBZLKg0FhonBNUaX80QLl+CeXNYdsC25
631saZ9pzxDyTPB18jwm6qDDKz6keeqpAiYZeh8ATEuqvlkLTjunWLc66m5YCGKa
THwEvC5iOz6nf1FDG0nuNEtII0Jr6UZ8DgFxcdANwSpnEfm6V+loUaKDkLwQBYVz
m5RCpVGEsjArQ6rysi8uHQB5c4v1pA4zxHHJCWzBek1Gus7EO+WUVmKX67+xyreD
dx88CHorYzi4XGfVdzjAqRySDVWY40/uErbd61ujkYJAHrU0GnlLExfC+IrJePI8
Ucvas1irEHdlx6o7yDm/ReKpIZ5pTEvNIReR0NgZlQAzau2hsx/BW0ekrPYrD75y
bI2yoUWkpotVa+uyzfkQkGgAGdM/3/brtQXU/glR/BmQo2rtXohAQNvG5vD0yV9f
eCbtKnpch6XGo8JFWHigJvuPgNt+aJyTEECsECJjeH3RckJ6I0K18tdK9oJBHc/D
FIk/eWbpY/ubIl7L6RoDzO+choLo/T8m+PB1RVfTPC6Q0p5BaEsdEBGkVAdhXK36
dkpNEc35tqBe5Xu8JqDvDiA74p04PGDq6gvfoUR+qRwNRY/k1zZrze7Y2Z6H3X+p
7bfAZlijgHEoSwPXWP/2gbZmR23sr0xZUzmzolYTnDv9K3+cBVvXudwRxyDRauAv
qyiCxKziRhG5tfGpqY1s4SzXc5vJ+TXfFsd/Jm+sKwLIaTFYPis9ng2xLj+tgmlQ
FWLWThfN32CrkoC+74vaLdhV3d5ry7Dt4eBBsOareEfj6cwAA9z95u3py4z7QaQ3
CcnPeeELoDj31KgY7uisSw/G28TZIn3ELAjlthL2+RVTdrDsdzZEvYcI6YzsyqWo
JAQJ6qRbx7dU9GDoOihjs8MCepP0dSnMTUdzfwx4qC3ZEW1xxUErD00K4qadYn76
LjKLz9jRHJvPktuUeGyKmohrG/22VxvSCNmNhAEWBaOorH3begBMX4XRvl/Pei2V
Uy5WOZfsXPWDb7j8qEKsB4H5hjn9OaVnFW3X2EZj9mOoc1HMGuc7eFWbtO9J61hG
PJXBde4S19xowU3whWR3BPoKhZrzOcBC/djjQYRKrwcG2xZ5Ud9TNu+yH1YQ9RQN
Ao8jEpnuIPOGEExuDgf15BEY9N0JUAwLQQz6ZdnPadQawt+QqiUA6U7FBvi5eqKe
yjm8KhDClscoK1KC+TGCPAPGZmExn2tHONPaegcgU+73+766t+WENZ3F4jA1q4PO
67HZSv7VSKZr3jPxfT17byH4qZhn3Jgp4rV5prw9YA8y/z2pvXO/VLbI6LEcU5Pa
1vYx2En1twF2nkigq/ACAY1Vi6nGonHhRTgDRUtNQl1OqaulZSez9uR0Y0dqr6Rc
Z+wmPvfgdjyyeL/eW3rK8R/FJkxY4yRK6v/CZwbRHAvTPfomfW8WxS53lz3+yrBf
RaCs7oXwoIDLTZahzne13bo9st1MZ7rmwZ+giyOMMMIW8hG+q4zXbvCLVuE4hKoF
K3sk2o35Cj1WMcdCjB2n/B5tlgr21Vbx5meBJbD3tqGTdTJljq/n5INwm0DZiN1H
x7aRUw7gfYfOsEsKOMzvzU857R+GMuyDyzsmMS2CsVFwRiObt0Kr2Dwaq1WtRtYp
RHFiFOJTzTsXDYumQiql6l7OkzbfEDs9y/b1t7v36S06OMp/kIjwdM9MDJ0MyLTI
GNx8DMvo6qr2wrCt4RAwG40hinbmRoNEwIssyVxjfRnMkeqe5Dvs10AaWTyJgB2Y
K5FFnVSOSwbn3MtJDpPYSwbK7W08ueszocE9LPIYAZUVG7rWUg/4shfKvf7cP68T
ngX7/lCRDgZBjeV0gRPAdHPELN+tEAfQ8UyI2TZBZbZm0L6QeY5gyRWgwqXaGZKn
R+dwjgPCK+ifRl/xEJBnYX4jztgMqD9IgDGBkiNcIYMsvuu2UzQZvdwWJE/xvV4j
SlP1FX3TWQP5sHLGWKGzoG+OGRnIAMYzlqDvENaKJSp9YcEXXA5zhCoLgrLhtnp+
30MJD0ta0UbOqnge/EXET/99SoCaI1s0wgYz3T88zJpKi+gziKvyBn+vRtIWb8YT
bLiKmNJgbOoMB99YF4hKKppGI+quOjs3nU8jTpwztq6xZ1AUvnyy4zgxwTXywsQk
2UW37U+mlzt+1fVK3Rqnxo046cJ2SjXt/9u7PpIfxu+0Q/6LkLTzQKvw0mybd5Wu
9jQAKaRZ4RznssMIVPnFViDE+sjcx+jhKspHicmG04hRTK4S1xCvcNHgG1aHWhGE
l2PgbBnioMUGyjLPs3KrtRY6c4Oqy3SOlWpI5W1I9J5/uccYKHqxIWyLbVoLkZPR
0GfOhv1gnNx0JEbxqlKBrJ2LJbS6iUgTOq653pAKkfj/d6oFZqBtNqpAlufKLYHx
TFSXLhtDKCg5lJgUAgmfz06YbnfwgGeepk7ELjzx+CNEuxHk5y58tOTRb5pnDvQm
U1NXTk8zgQuxyv3bZCgAMkF0VdLtBsEZGT1UyBypkmztn6HXBKWIskW4FSyEn8M3
T+8f9jDJ6jTEENcA2aA30dnIsp/aaTwNinbBKdulei4FpsxhAEKtgJFCd2sOp6MB
BU61qy0Ygw66j4hV7lzjNO3iazM8M4SMrMeyLdoxad8NSLwgS4C1nh9rebwQl/pi
XPXYSL85qqV5LVizyOaR0bhNkfs0tPUcGzmpnsSQWpUolGv5s05xGJRQUUnSd2ay
ZB7l+cxud3H89yNRuJv9hNWiYTyGf7pzytpaWKrPlVQWWSL9ASjEbhN5zHP0iDPm
DLIOeNxQkfL8CG7p9S8GIBhw4BLVKEhc/spjOe/fddmasNP7AqK9/PelF7Q9VY5q
/5bKrZT+CihoVnebDJ0qxtjS/9WUUgKykAeftWv1TYJrCPclUG02rJa52MlwE/ro
vcLurX0polsvIDpnWf5ekQNlrjL+/UUgTurInn9NEui8d797C83zE9xszJURfFF/
Kdm8NxvNsf7flNhG5mdqjURZfWcsp28TXXvaewqOV9Knp7oVVZS3kljLjWi4yp0X
88NF4hVr6990V2ZURc/2o95PjUnn7SiwIOuCptYtn9hPj/xbuXf7Svj88q/kn3U+
64qJ3L4qbjQIlthsR45ISLsBdFXvsfE317mTj7KFes5C7MqW92krzlWu7GZTF6u/
AgxrxVTY8xfXHNYBSGhzfS1Z0Zi39lbaZVZsM3nUpHzGgLsPyDrWsec5p3sLPq4g
5tsUsYy1F19fJcAsJBuqtFwUTxkaV1THgxygcoJkX0y7UAxImOcOKLz0Ug/CpUMy
wbLl3zJnqG5m4E0TGkHTKEXsV6Kl0ov99TO7rcZCXiJ5wY/82do2NoxMqpHHcQzQ
oaGE5O7eWweSiJHjNQoEqRcn+KhPRF3BbTw8V37oZbUUIZ0KTp3dT1Zb4TfvYvR9
8I/0/td9xKm02zkX5kRPh/f+3nN59KoxGGqcllLBGUQUCq0zmOYPNtKr3kYW39xn
ihYS15yI01s6udXdapVryBvUWVjHCGFoowk/wAGSHg7u2iMjmTDzPJaq6d8S2EGB
9jCGrm8Tvm0EleWFYnN7xLMlRrRNtUVDNa7U6a3LoshnRUVCJ39QYGy9F24hbQVW
z7JJL3D3mQNDOI7nQYWyCiCd4xKQXG1Nvqj842n2r6yzmNn0PLamGv+CqQrgRRsw
puUWYVVXZGL+mnz7UwP+iS11g5zCzia4zxViT+TVVGAo2KGhgrzDTL4yNNL/CRSV
EBGHMd7jN+TXHZ3zASIL4RznaWNXqxuddcufiCqjPKi5Rf/F7LeEyk/bMidHx4U7
JJuo0UdoSqr/IkB/AUNPjzuh9yDXzEY15Kcw4QO4Af4zAZBSRSYTH1mqa5rL1hyo
EHWN1tzHy14Nng+TNdobJrIa5/B361VJwmekGQdJEWxutYqfE62AJG9MX2MJl0vY
q3HniL1xGC8aerw0NYOom5f9sX01UAEXXWGaiZFWZlKMgMMcFJMN8ZTG4IfpElXB
ixz9GuebD9hcunD6ZDXogpnpkSigvcQTckZqxba0cbzGkrjm3nfl9a2Jk7u5TIwv
0D11kzd/6aho5aw837YaNFuKy621xl+89cWDit63oYG58/4mn+4aMjzz3qPUVdyp
Adx+aSwbvOkr6280xAIG6++bAjwV5VhabVxsw/7m/n1SbcK931lRmQEB0CPFMVx/
Q0VERsgroUGlffs6RfWkFXO90rmvOkzL74pcAof7H/YiZX0yGvTwvDqRInh+bKfk
v0mSQMwE/jvvVIQcx0r2TZHkSSdAWJ2VDY3y8qBYBfnB4ZbBQjZWSeAgUa+PBL6r
+4WlIPnwLfT+LXFlhLvs5kBHw82dFD4oYdAkcRJV1J4jDHoHmPPYxp5JSJ1LgtWB
Z0c4y2vCYnj67QyFDo+ademR1ddtCEH8JmDE9dWvwLeKtFHcADYrE6vXhzcNam9G
jR0H4afGWmbmaTboU5J9vWOb5DvdaepJd1BYlWnRzFOU1D5wVkjKECOsEkYhryAi
MoXXRYgnAPyjdt2FPe2E7p4QrXfpMOyAKb2xLzZhHeIQFDRvMXkzYvagSr1ooXxu
8flUh9abmgGaIIk+t/HKe+gdkXnVK9vMYpOMbVvZBJi1uk+ioBXGD6/by9SSCVYj
1nQATTU1Mbj+1/IsQ/4MDHsesPmv7m3qzsKhv+Z1HlnHv0PsRWNwBvafHqXLhmp0
yNk2jDPhjrmOEApEKWIKn6rUcYP3YKZRS6XpDTzXY7rsm5QHf0L5Ku8xXL0uFwmp
mhuxoSbOG70kXCnRwaJPHNCj8ysnynuGnHrmGGypmI+ibpVWUgOBmVluc+lbXETm
hzx3L3LQEhH+2P6Nac92t1iOlOL9ovsTZ+aRA/GiDwM/ny9BMAjvGMkKSfi6PoFq
MCnJ3vvX/jIYlG7YVa9adIXJnaf7tvD7YZH7BrTkweZbVr+EzZUVl4S2ftwzKnGB
lXdHWcSqmX7jd63mZH9WSynvSE2Bu0vEtWOR47xZwl56RPbiQurBdeGpSvfaYicP
xUma6QPhHFT2TfWJI+UGH8XYnU+pWPNSek0bDnbMUsko8OAN+QkoSJgJeDXzwaPx
s1vWy2cbfhHWiOil6Aj+OVgtr6V4q71hCNOdSiiczaTHRvzTRocnx3eBvKapnAKm
3p/tYUCxUpXQZzZmR3sTIqe7obcvIFmvDuOoME04amtusNQGiEgO0vWefKsFeeKk
/bFfV2RzMVuLYT8XnMrUmDjShy+sX8Qx+Pe+rWRvX+7bJ6SUbTerhkGBRQu1ttEe
ayxUOTkxkxb2B5bPzk/m8enc0gwmrOaPeigJQPYlhZ3hDLp10zPggdF/fvrHCrmK
3MoDnqjWnjEkKo+8VkPdo5EDVi6slEiSaCSmCPMHPUqv9aVCTYuUXYkdq1zqAfcy
kyEH2TsfhBle3kk2Cd/u4XkjUMCVJbqBgx3QBMv7nRxk+YN5qgpzhdXw6brOwY0g
rla73mH3hJowtBQzH7c+C8f52/oagePQ9aIm/QCrPBVi272aaK1VjNm2rl6o+z06
YIi6+mpyrpvyIB8n62DquBEcHv2N6nqv3ZYclMZHaSvMPfsOAaDifW8JV4+JIDgL
mSQZHw4ycriZ0G79xVE8XYBZurhm3eSqTUTlgw5xW/a+r4MANtXw2ljR11FicQoO
GZ77WjCoxg/uu2akuDjfwUjbE5Gjb/iJygxqdBCPXmS7zUF4swCOCW1zGWeebKPn
Bufz3LHkX/lV2QKzvXDkz1Pyyf+EcXXoxHFNU3SAHBVbjzcKNSv3sq3KH2mrS5+A
5zcT+rspuQyGpYi8Uf4aeINcpBcBGss91hIZKh9buswCzDPLh9YQZpijRo6jOE9t
tBO99F3sfDKWBx7eIT7buD8g88Nu9zfh/u+38b5K5DEMxR4deWI//ZjCthi3cx2c
E6fTY9ED3zGLpg+aFLDSKUN/vHKZTOIh2om0G7V+3xpk3J3SGIqC2DV/2tO/A0kB
MSn+kfInoWG2auKY82QLxlBGk4uvgb+0+zkkPsNWt3rk+udH11w5Y8G3GllB1C23
+CGzrc8YYvGLqbU9U/TmGFK7idiHudi70AIqtIi0nVySoQueOqEiYK8CBOVn3ivW
/1kttGn1MUsJTxhXJcqgu6W1LWEsuEbWV6t79PHn6IWvaYb9jyAprFk9sEzaHSXE
3vBXBHzPcLo/MTecx19iAoVtUKAKaV3dqSV2ibzL26Qh6cvkJvfdoxQ4nLn6iceX
5bBmycudVfVe770DldzYwiVghIjWCxwUUC9QwNEtIXnajeECwQ1jxlVf0GzaZP9g
JlkZnVQabzzaMHWzFlQVXN5N5KwTS8SxQSdtFgFRBr+eHkO9QYe0jYW5CwhUgk6o
zcZxqbzdeXBf25gu5rYsha7951pgvnAI9enRFPoKfIZK1AAcxZJRvVPiPu1U+8/z
+siAEL6vf/nVllPJX0Ud9Akthb183oWpo+GbK5Uu9FpaMiimbrLK7k12taJH8m7H
Q6Gg/gMc9uW5VyOhpIGkTCQY+yFcInePvpXsQuUr0GSfkMlwtpYoGXpEfK8Zdt6Z
3o71rGe56xbJlbwBBMtaeqTM+WeAiLDrX21oAVPkcVLqp9ee5LwPmPbtGg71UnPW
YRBOniweQuHnFuLDJlcsstZ6Vur36cAp2tSDSOSfANmgGhwt6L+vmAi0LKGv01O5
2oQD2+8GzSqDofIq7RIdiiYSe6wH5QkzcR5JTahY26b/5MkKezBX0DqPX/iZqVzL
KZ3khtyqISjJo8uuAw3fCAW7YvX2+IWIlQ0LdGBbpz6RwWcX1xRa2ts/PKWxTz91
hfoSRD5MFazsMXrTmGdxzJQiYObFQVFFuYNP//1aT5q9kG6kRmWmqnIo2+jwRAEv
zZjJNZo/ze1uxadUKNc/yr28WyNqueURX570QTl6ZxKc1B/sRDROAl2YaMeZWp3z
+mU9woyqyxjoMOZSqOIVMRDqiIzEAxek0nAhmcihzjzJIMuKBmAWZdw0S+0amerQ
xawTU/MEoQUUEVpvv9+I1WLhWsSdOD9znJlDfEhBkAEMV5VRR/4OO/CCS71ROlNX
NWqCoec2y5a4qLQj1Y6QsCrfNQzxUTf3Tt9u1d+jdQsxN5HS8hQB4ttSqwN/oY90
toOcGhd/mXYSv4AZrOFA8jZTK3MTgiZ8xb/ajS6RqPutGUvll6Kl49VXfCECrcb+
VsgkKMQiFdJA0wixtAHD8cPoUqv+uxzttM4pLdgtplR2GvkJbFeZwqZrwZHyqMkv
1RjXMZg0bMxoBjtsFWIArAyNs/wq35W7OjC7ILpYd2Qz2E+PU6uJy34RiPN/vGyC
b06cPVYQGN6fps3Aj3FpMatCe3bkIlL7xj0AxoIOwRipl3tpaGdbpcpnRkYeW2U7
z6AA58Z+S6WKocXaicaqUb5x8G9GqT3z8MRmnKdJIQT4Wm/TPrnyerhK/iivEA1r
OvDKtlUpSrvTfMKxwYpxK1Vtz6DEIsT/dWD3r7xXR+3k6KRa4klyoXRWDB8QfWwo
mcIu4MX6D87R8kmOhPRoQWAnPKRNmbFAisT0fhdGokXtcM8//hIwd08+P+OaRF4G
ua72JVm1sJIf4r9Wn9G0n1HWReW7U4a/9jNGhi0pe2DCebEuzRKai/UEL9SPo1c5
9NKpRsGgzph498DnZmYG6G0lwcfp1U9sxU713FcZyj0IchabAPiBU4xjTlNNwkhh
YLyCNJfyqNNvMaYxo93MOzR3kTk64FP8o0CCpjCTtFXEwhovGplYaeJ3btzF0lGX
2zpkY7pLmSALLxT4+bH8aNCJGJqvc3GMW/am6363v3hm4lCSswR2Ylu3SOP9CJbX
iDt5T5+ryUtFfvn8Y/rvkSVwiZ0zFJgsUTLwWLEwEANmghKVzOkv/sKflAQjfRKU
C1ItozbUPqpiXD2lNS0PVTrUs25F7o6yFzh25XAZAl+KLSCL7WIUnp6qaqj5x7zl
11I3bkpeXYkOXb36xXrDUZJz7y/gEdyuObeGWdD+sT8LteQEFVdtGdg0Z4PM7eMK
LNkkDJSHUi2XvLWkjq7nUw4welBQtMRXRIqtul45vCglh+ADkwMQupKa9ZRd+OAi
Nz/Vj/zAwcvJDTxXwVBTBhIuCj6A5sEjUmMNyEmCatebLRaupSf4gYtXArCrKboX
Qdt1RtIWPgGw8douTrtbMRtKkLKOv6Jkn0Zy39YIW4xczIbh8YmPe/zgvFhVIPj1
Zh7yNycyokJj2kFqIUuJGE/j3q+Kob1oCaVcPlNXnAZ40RRxgL84M2cMVQ4DSvYq
Zd1nEVLsCD5qbI1ztZt9hO6DtGrx3o5uHFIbcrSMsx89JTcoN5CH955BJaVj0C5e
hm+jXgi/GrAKomx/cGxX/1Xt1VSpigiEEv7dO6j9PhrTkC4PM0QbVKivaHSG6kY2
ZS3d3uYdKHahQLo9DemHQKGWK0Osvfb0ASlCVhZlc8NZIGcfPGwqxc9FdpqmbohV
BUfI6wNNWNRwGuzp6f3ap9EZ0NDaXchbhKHwDz/DI8uaE4KxYvYdbyBsrVt1dAxL
8vOqTKVEorx/ADCkoSTLVIepOJWMZ1bRPa8KJzL5QuyW5WMTmZ/6rHDj8SsZ0sGO
9JIXzcR7p7gUQCb+PuBYeAkFO8k91NtliOzpWbCsjeIul5IlfsbyUY5ZHAORToYu
BgMYWEaGaomc9aC1c+n48lOQdMBDDBYTpJPYi0kppJERVTWUo/0ebzjv2cTQTkmt
YIOKPJJs18c3pmiZNRFExr2VTWLcSYwRE+cr81NMbDAMG0cjzEmnmI9CwICUwkh7
i4djIgSq7HLpF7uBZUrtmnSo/KYfe8TgDbBNDsMaB0GmVqmkXiBGEyJ8aP7oIRVM
nydaljLg7roAcgnZL0zfhznFATIyyrT609G1nBgCkM60mryyZbWW8RwoNEcrWSww
eWr99ihywx8D6S77Kk0GS9zURDUAPRVX+ry+n7GwqDHJljdKYYK/zBGFl37L0mkd
FYmyOZt338XII0oHqmmP05NyQ8wERTrSbCuTE39yy5nwkZGvbFCeaL5/pDSPWuqW
YI6NRigvDA6zbU8ucrlWkjqJDf3LWQ/1AABQxovJg4towye+ie7jusSYnXvxbsXz
v1EOu3V5U4mGFbtUn8ut7WBcgqzRyxGQ7QYywLqLc+BM/IK89b1W0JZ3ktQcafsA
3OBelq5/TfBBIAErOKxv3lmP68OjUfNaPjds0QHH5LSynwZfvj5favcEduMDY20f
iXqIctwDNmcFSyYxjhx/n5pvD3DHLTPbFvFmgAXlv/DmFWotBxNks2iq85AQzSPc
42mc1UCjlTusdBKCAo1vTjzumWAghYXIhGAuUHl9KT72CWZvGX+Ndr2dPL4DeQVH
hG0bi/Ip/cJkY6rL0Bq4mdJA2qePXxARIP5b/1dFWpEA9ghZkd4mQRBzAJueCBGt
1cJ7vY2aXAv6oiPa6Rs/6aT0jrV5ohhU0dqMVOEhtB1Gq/lfRXwWAa8eJxlXuFC4
+vKd6QzFvURy5jlq16mZX+SBziJbs6cmuDxJrdJhkBBJwV7lVFE2/mgYwFBMb6bj
HgN8lD8MGXDQAMmxRHG79FJ7ZAeADH16A7lYhDPRWzuE7v3mDH5N0sAXW+oj5z3r
LUt1ylfVArQZpuKxLIa0aS9I0UYIFD1/ConKccMabqMSiqzD7621ubfU6OkVmDL2
f/jRTfCq4AsC9aO28lj8U+6+ek4/luf41WAtKL3Ys+YV2MszVjxlsevSXLyLGO/W
iNN4dVgBSt/W4PleHxoALredBq4oEONgdwMWo2MnahqbCJZ7a1VfvMLZhKZqBxvq
hMeASOb3hAt2JQSwKwVyhN3jRJ0IosE0R41+j+hjlVnKNWrkQmUttnaFzuT8W0zK
GKii2cu7/Db+ymZLWRkOIYHP54eWnJp8dQv4kH5VW97nCT5SghVk1p8tNH+qVgFs
La+LG01gyav6craGCFjbpdG14HG193ubn2fx2OYON6TFtikEqWvOlNZ1iyphzbTA
nKfZ/m1sgDpjWztNHNdn89iNugNiOxmXLubuuvAWBKG7c0/BvnyXcsfnolRhn+CN
OS1vFV+0UPP5yzTbR766O0cAnyHBRkVUa3nunuOjmEepDnf/eR1Kg/uqbUA71nl8
UnMiZcikbdDGFr1xzmPr5GZa+vYVXhU//Be0Lik0tPIjhZRTTiGXdDK7dM6wBNYS
ciTFCfcPGQ0uyVYD3jql8h44/PsyAFW0LMmaf6Butcqu7xWMTbt4S8v/wFc3MyT8
c7Yc2Gu+hYvngB1oGS0K1UHgnB+vGcJqKp0Aw8oK6C96xw/SJm7bB/Kt+ZjY7K1W
tMbxFsWXT55Xwgq2W9C/XzTwN2VedUDA2kX/7U76dtXNOGwUlfjz6XHgQ3UE87rF
0Gbq8MSY/neRjzEBjJa01mEkAjSWIOzzlIkUAaLBP4U6gksz91jzIhT2fwZpxvJ2
bN4XwWwhlNE8C2KBoHZEdj6V9sXIPXDIkpqnvnkhhjrUkQFlLJ5BgYdVU/p6C1OU
BwW0xNo+Sc/rraUAJErXC/Z2uYMMNJMIC84/OXGhqUDXh7eZtpQfrY0HgyyPfpV0
ID6U3pqXR8vmX9aHubpOkB3+kn4fI5ZpYXzNJXligbk2omPi3z7A0WmgNFQGVvMM
By/oGMe9v3UY8qEx+oI/crxu9YRIj8l5weowykc8+RmbkF1R2AVfC6w6FzJSXwOW
koB2nzZyPhj78TLquetIFq5awWMUmA40BYSf6WmT9FigCk15qePm0zp60ora3lVg
JiMC5XCQMgSOuxezInCr1SA9VdrxrVGYKeGjtiP0G0OUIkQ1jUGtXL8nHcwRoOv3
+aVKh7Z+3fwVUGlmelZcZ7EH/LuE043tcyuePKu2U/MIc8aI8vFH5NjG5rn8WXOv
b11FoJFE+RwS0JllpcaRYJqUrmaEj1RXNMzFXlJRw8IEgjeBqj+dHQZuOWz74SwO
CFkKTawWc0aTYK0pV2tdBrLjOZ3y4TyDzULfTZddnQdA9Z3mJUFE4L5R4s+X3lob
nBFIeLGgqldTMdbUKU3PfMyy/QyQob5XP5Umx8J+Vrzc41qy+XExppnrJ4HwpDsO
9zY3d37fm89MBHsFr3eqyILvVtdSgIF/sJCq9ZaCpZ9e421NpdteDKbGw6Mjm10A
mzBTJiqydqPfo0p36qKFdd6y21QYscjnOJ/qzfiMoZR0Pwzk4k56mneX7g4WJEDy
+Ugksh13Kgzjdk8cfCRURcFChrzGz57bHZkwdvGIslBehoNpjH66YNqHVqgvZZS9
Z8MAwHAepF25/TT14PnIXXuS6TwNbRbUFEqy3+nnBpvFkTRIrdbntWu0jO6aXNl+
dH8SG7HuHKG/t/34bPqjCFsQVWzwWrutilyvyqdh6zOAghIvD++CBNBCdUHpLM3t
TCAv3UpH5+6PuYNXpuOrnlnfYVOg+hvgOsFj2K/moakOAnDfTEK6pSMkgpK8ds1J
EZcVQJzCQmgRwW5m7L2fLvqaz0RWZvUbdX44ryvcuMvILsXXmEjZ6SEKr6VN0hdE
QmY6uhkfdA0X4X7O4rHZIxPg2lHUzzFvU2oe4SUozf0yiIK3h2OoBJi1C4uAvqIe
J6AKaPCAuNzYZkgAbKUsiw7ZsfxC0Wsx8Hb4J3JmWr0wKkmHlv8s69/xTuf125Gm
/M8fKs3oWvbk2MGuPWdNsg9R5pV0gsXKSbUCE80s65lMmDBrNP8Y7BaJWbFUJy6k
bm/aOb+2PBh7Olz5uCnzfOka5jPxreWEJQh9wZuOTJ6ubIZgUUy+unZOsJpSValI
2UmZwRnKoGFyUXoelSLN/3bwY64qBJrxRGMjLpiaT3/qMH5jHrZ9UCJnIVIWJ3qk
mjfEvHqSWQONMkjVYBzBMP8AJb1WqTaRsHi6Cu9QmJpYfyW3gY3e8wYq2TI9lxcV
nuw7ltzlmtsECTXDo4i8qZVyejKy7Ze0p/JGSXrKfOvEcqEPlkxjDiMSOFw8LohT
u2cH7C8uxvleVzeEWSlAR16CmUnlCMVZuUw2SE1stVzTmWEzjJOWBHnt59xwj5Su
MXEw+zJhs/7Gq5/q0ejaGl84nWZSByABjUpigsf2DVCQpYc2F6SHC9xO/SDPSVrt
1l4awIs36s5lnWUq8rYdXicfpgnlLLO1JYIneD6VV7Rco6lCuXrylezGGyyreXcP
qpgicAWRQb72aU4/UmMbvOLelEMuPe1SkGbbGBw+5WpfIT3F6VLHz2nhkbyh+who
rWrlYKFD4/ze8Do+Bc0L4W1OH0lOa4UcPHBCIGuiBjozdzbN816GBjlAYNKDOT4i
po5wL8ifzLH51BoFmUHd1lqueK2tC/YrM4BYU4s5HbPa0tLGtd5se1IbCoS/bPM1
XPq0iVf1j8ycq1tsMmLrmRXYNPNQjL4VPGGWQrL/4/lpnumhpiwQEpcTLo0DmQgL
Dfjn/4X79++8a/vDfL1SS+D4blW6A10hg3K7YhfGoIPDu7BEIo032rprmTgVemMc
R6T0FXAhBMoMKjrCUnk7Bk/VJoJVn6JlnYMUK62I0HT/igYhPcyJiJk4khK3R8lD
VNDUkUQISoICaMQFIUnpHCaWSMytdds+FQa3sYIHCGs1/yL3vfZRJiK2BIiNssv5
s/44hcjtIxChLv2L7wTCu/PM7TwGDtJRYqQReOU+iWxsl6P4W67v7Q+epSt/fHM2
1yxZCdGZ3zcmdyww3oVt/uyAO6BD4On9Xbnecm+LC3gnXuNV/HWCNR22naxwCilT
VALzblZUgtl/WPsDtuoLN+HiepUevLzyr0l66n5Z8LGkeynSsdFriVAwlpKYtiGc
9X/YFU8DsUFmKQZdkeI7Pre377EpnFawL9ssRUPQkrpCW6u4fGPJ3MU/iyJxxcP1
D6/vvLF8eCLfazgug9qiu1TtYY+cx8pHFWNFr51SC7QfxOSU8kBLAlmxRMd+Q4ft
A/mHU4sAGXXirPC5FEmvI+uXkt8BOs4We8LOOIO+tA74asaP8MMm1jCIGSaQXBQk
fxwGTd9NDXnanBM9+ZzHDPoAxFyklyfPSTizJGJQLqK12YQpZJ1iLp/c+KW3BRe3
tMgv7OfNjPOPdseOQe/II9tGwzRIDv0sJada6Drs0WEJoWOTh/ts9wYf6FxQhi38
seY/nJI77rSurBpetC+nWjoA020AbtAs1rmpsuoW5bBh3GihTJ7knO3putXbYl93
IPNsQlC9kLVp2MUfLCcEewq5x24PCDD34MKdJ42sNzlniEUBqhnJmugTCxlLKi1t
HeHfb8fYOjsfDYCscEqr5M0DUnmIqO55XOnOwq0sIVh8VIpUb2OIMJhdWs6pnDc7
lYpV8DHk0z99TPrR/j2g8OKt1oIxbGTTjXcGcmWpWKZqn5rG1bKuM0wtFBY+XAPU
Ts8lLe0S09TgGw6wGa0RQKJ5o9xBXkgNYDd4VRcSTjOAluxVdKkcfvj9Ra9Ed+MB
Exf/GS6B3NTY2ESaJeQu8GMB8q3hwvG/dWSUvxPWdnhdulpUMCdwy7dS0F8zczyO
zidPxLAppywsIA0QbMVDuetk33q6ERuSbYin0ueOwflOcUUZMVEpFnU3xLD/w2+Z
cDUkKGodJpnEnbNpXOTYBCOgFv1HbiagPsv7Y+jL2TNu4DvO5chXPVnTzTe9fTk8
t5XdbY0rfE/qC1MnNHWdfHaa5sohgRbCceIvWHJvr1Dn4M0zaLTGwIxGEvqQ+GPP
M0dCc/hE7tCe1r6DyadkBCrPBu3lVflMkwY2vme8HFyCQ+3nskyMf9PgmAR1Y4NP
O/dBywQUyeVeHNlm1y1G40AI4qGg/9ioyrFXg/cav6yaoJHXGyu9uOTeUD1kE0Wg
o+wAVF4NG3F9aYgcm3BOgNaJ/Cqp/WXEMS5tIGdGkcxN5U4xTYlt0sJHCo+jpbIo
yCQfND417cd8IXVMtGM7earqs4WMw2ua5jJn+QQdvGzTufUV1ZHm9dOXUytf3YFs
KA7FD6gvxWCOwshvXx8C/cquo5/rD2cBsvevjJ6BtcTruzbKqgO8i2UTT0BCLrvF
lTqHc03rapNQcFTExq9O6nTmVbvSj7cf5wUVyqqaqvVdtwCMUuesxQ2v7znHYFOJ
RYsGnyPYb1YfzdhU1aA2GXGXDHy0P3zVvV2+ZGGnk48rzzQlkFSbM+0XCO2jF+eu
frV3a1C+fMrkKpBm4zU68CcYfBEQo5+88rR7h139l+pFSeZQwkjZN917E6leJYPz
QlG4DE6VgtdPQ5z6WjomT1hEYeA5jOrdhrfsfwr+f9QDAe2tCe1+D06hu8Ec0D3O
+nF+2wFbpzyohlFGXGE0kEGiGjXpQwlwh0b52M4SHrGcymYJx/n14D2SyECKTkM/
J4vzN1hSDeaBw+DpkbCnUak517n6iiPbN0tsKf+WfPPNrpxF+vBnmLh7Z4Ss8V+Q
CfSVJGptex/siQRxmPBXaMsgzZ5smtJbeDp7nI5hLGTqvyIYDDNcw7jWNEnBx6s7
eCFNh2yspgDJQ8tyYxoBqdKqXTDqJ8jz/6s0igvGP1VjdALE4SGiEpF7w54MkiTX
EyG3qrof+j/U3rTsmG0bLH35T6H3Vgoon+gJoV9aFIdgD6U/HQ9gy1/HyEiLPY2w
gXFRXZzkV6Xp6DhFFLscl7Cq04IeQYpP/2a7dVSKauo3PtCAHqdTLaELdVwXsB+p
8wxDO+y+q3u5qVWpDg0YZAfNtDhYRxI2Bw8ghFr1fWgfV+UUqc71d/IwTneQJrep
6DEWYOh4yk5cisZoMUKwowoKNr46Jxu77yngLEKYSwrw1o35lVeeHoXRvE2+D7c4
AV/YOw/P2hX6wL7cohN0V/sED110fLWGFa8UYYoraloaGc0OtQD5Hk13YkTyfUpp
zatBAS774g4yj7usp8w7HhwkZ3pHhPKkNbq5yCMgwW5pbx/eP1Fn6HlpmKiMZbEk
YBO9u+5q1KhbvrFWf8LCoAfYHIEptuODVXz4YV9Iu4EPNJQbtW483NBS+m3xxwNL
ovCd6zjfdLze88n+nihKE6Bi7Q5gbAQYWbzysGq8DE2yu8m/rARP7PlSwg/UqdH2
k1GgddyZbdkcDckGPSdpd6PjKqPTw1nnuEbtPgzbsKPtk0DzOl8FeUimB2rUibd4
jObFXGdE5qHoX8p4cX8Y0D7HDhYiGF64eIDS4gnv6b5gbU706IaBC2ORCIpQjdfj
L8grPgJYK/Yrzd5EJYRUvQSvAjit/SNKZT9UICtpW2K81u4Q5nbJTMCZkOWGi8an
Ne9KKc+5gYMjCCbPAbDlFyaulX51YKdESbMqjSKEovPJWACSNTt7UIVCJNydJ1AX
lbkU2GRm0TZQfxoWy/oq0n4j9K/ZaHrzjfjKPIXmHSFIbz+DNprznJ94E13XRvh2
6A88Qy82zLEMBB01E8vFmTM9drfx+II43pyUSaZNmJVc6hK1Bj1xiXq3+P2trckp
SVtEEcQwMQ927GqQHtTolghj8BzwJOat8vsq0ZMTFZtYBy4v0mlpWDAWfKbM9GQ3
R3rur7m+4ulRw3LtMxTaKnJt6cZ9ZGfucRd2aHSfoI9HYeNpmZ1/Gb9A5dsSYD4R
E00Aj8leYIrdL0cyvALtEUoUDKhnxSLMGvg0+CYtUTT22LjzA0TnFIIMvWHN6Jbk
jNbdL3LTxMpOQTTTCBJ14EQ2iRdLl5jjXquZDNQyo77eoRxittklF3VoS+Rre4G0
feNGtLc2CslHfiFWORcWClshL/YKc8owHhUwM9M1rQuj9ZCh+9uObtKzvhoaBJ50
mKKZIT+3VYXwYhNXwjjoy5hdJwsPkWOqONlFACfldVa1xNl3NETj63ozRKzc1PYW
0QeFsVP9hrPfRvg32JTYoIYDLaAnRCjKVIMb6Da0iCsgX3Ei89kuK08F0scIBhLZ
974VzRiNRGwHfOlL8pbhNodXNQNedLC3GugwWjgTiqT1cBbHSLap0Aj2sg6eZd6Z
PXBjmWSMOxXz0Mo8rcxPojkpy6xrywctR6mhneeUE1bRaI7Tq4y0hBKHldms5bp0
ovXdGwDHIeul+nlkXGplmUQ2xyE4CbppFM0A+bO10v+mTsQJtrsR0o3sL38rCJ1Z
Xvj8sjcoo17V6yaSLcgT5fWcijel116ABDNuyHAUvFxB39AXyZ3rxL2uxM74aM/v
pJ7a6z5UHsDuH+y9/wxpycb777slxI8RFlcTmih4G97SNGzMbnInGGIMPpCYG2wP
9tF4hejvWVFoDZPKx6/9cyiEJG/bT12S173B6Qds2nJZCm2sGi3KsqhkEjd8IfTE
+sTaKkO5RY6bl6LfsvHRNWVjvxsmWpMn/O0cfEv2muzJ33ORs0KPBuWSFfXwT+Nw
jdt0HB0nMO8MH7t2jZdO7euzmyXU6+WQG3PknJlRyf5wB/siZcG4V3xlr9/J2uxc
zdBOMailBXSdPzKs4dmmzSgbzBQm/3BepsfPeJbxV37BLRB/qbPeSocGCn1mhhnf
aVeNRVGVb9HuhuMd0JZsdVbWPapAt901JQUpYmx2W4ZNwkKmXaHfOzzcCYQB9jLA
NKrpGrqlIga7V1Sudcbrcn/rGxQOzRV5Lf0N+U4jI/Sh6XWJKzJ2s8zPbpzvTClp
5OenKCeFVcO408mEHv68OcWSJyf0qGK9PUpB0gvgYNjGGbpfECNK2rW7quZiQ4EL
EENQACmm05qPb8fYi8T14/2UV+ko6XH/LPC3fsibUIigzfdQhYLnjuWF7YJGLx1+
wYCVVGs9RFddCeDYhEdsCaRfi1a/EllDn6Vcg2FKswWY1IpTkJCRBrsgtslxM3AM
9iZ8t7PTf2DteouM+jrld0wfFIiujjJ2erSwbFYJeKLc7ZZBvYhucYGR3jMXZKsF
KLlgfDKJ3RogiWc5m5B2WcReAGaZKKOpdCkmcK7T62dQ6RaBdv5BAoMh7LpIZuGt
2ls6huQP9Zt3jD3XbfN5bVw3FntNAmRCCfv4vrNLgZHEbIiXMtFnfv5Hao5wq+N0
oxWpyl3h0tjSZCFG8+ujznBIIWChDJ29Ca9zjoSZUxUNOdfJjbO6IsEXfuDvWDpv
Dhv8xwbJcaMDMO9kaOjm3K+QgIQxi7TaOFwlHZS0FLkLrYiJILLFhRaa4oNh7pT+
/dT64zUK6ScETZkK4TAFQAHQzvcI82hhMJee0ajdSU9Kvb/dW9/FOMzzw2pX3W5c
0/3KSPX/YokLviEmVtt8ZJl+KvqIbb/ZlbZbQKkXDx0oZ8pErboDlxcX+NCs4gJa
BVApU0g7CIEO2mQq0TYb/vmoPDSH2RFutXdIheCi+x+WlQUQQ2DCUUexWPPw8s2y
MzMcMOTH33J1AfFRo4m46Oz/pr+RPu3JPG4pCnhzUkCr9PTtmlDGCqOFq+x7EyH7
YcXYx6ey1jzI5GdH2dA+Rq0iqMeYMbiHIMLywc3q5EJrXLKe2dzQH9DOWvNrVKQD
bJFKsxN838eSDBewQgnkqCo2/8lveBroJfxY4HIFFTbwW8axMjoG7Cx1am/79VpG
xsmF4oftmDQ2U4DW4sXfHy2IQ+vF0tcNBjEMHN1zBvS5tgJ0NVtyuIFYMR6HREQ7
p3d6t3F84rnqHaS3cr3i07dxqItlvmL0VHBhkHQbdP1YPKrNeKipQeWlVcQjRUG2
Hyw/UkdOBTxJJ92y+HmMnYraKTaRbP3ekEsxwD5R5REv2gWEoOt0yeYSLrXEj4Uf
cf7BQ/Km6zMVjJArFa5vOPtGTSHkY6WCztNA01IdHu32UvwI348U/TtGjmYvX0jo
t0Rd04Q+sMRAVFvxJUoW+s7pM+DUEmimVZh/5nnejtw62aHUSIDBDL9t8yeCYqvY
rB5OtiC1WPhAWLtCMaCVNd56t6RkzzBsQcWwZ23aI5HbBRKq10Tf05PZ8IRk0dmN
lpGhHMjd8Kx6u3lbDjM0M7oAdas1X+Mrp9bFF+yq+koDToSt3kUe18X307RVG7pv
xkvCwjIsNjIujJ6RprkrrheFgwJ2OKwwd8LnpWG7/61iGQqTcJt20HZ3v0JD5Mc9
E/NUX2a6r/u/Iy/c0yxptfyv0kl+3t7Q2QXcG3buRwPkB4Fw7DnlkJ40+Sbdp3fZ
dBxYDFgOzbcvy7WbloWP6VbrWN5bESXi3z3DyjpWd/El2YfHI3z8+uQxCZQSm1Lb
hBEyzLvVpuYFap4wu5gvFcwLP8P5YDE5GBztj1oYKa9zVw3KFnhWBEZMgquk+iVX
YKWRAMWYzC5V/wJtLjiFa5x3fJ4+n5qdcSVflC+Nd3ZelKnp//9tsGQzlBb/qLsk
0W2SfjIYsrOtLqIkMXNGDRAap7+07nYAQkHtgDXFoCRT9Qc/wO3IsP7miQoPpk98
bH8PxktRKFWHh99iXvgwMbaw8Yxr3jEE5IW2OMl/JFVGkuw7H62jSAkVsxUnUZFr
Owl2xNIqirEyg7me/kLdq2D19MzKBttshEpAP27lKkA5qRmJ21TDkJAkt1RgDSPo
JJWG+ax3Uhk0DVvGRakMy4pDxWQziEreonlaArtU0rbQOskBOBHja/VnwXCjdpR3
Mg5OaYMV0HmlIC5eH4Yeav8qwFY0Uk8O9kCz87QegPCq2upt1hcdEAiD8g0Dfxfx
VtChbJX7UQ116OdbK4cOPl1EKGaHwVvE9X77jeVXwGrdDWxrFjNgfDPGchU+v9z+
1tB80md/rs9j76nXU6NeUw1Yln+N03AGLCVQ/s2fLC3ULn1HJI1sDsORPJInzB+z
QAtbGnE4H28CwQIqNRPcZuNYCSjea/4haIgjRCJutXs8JQq9XXgh/sOAcVm5qPYH
JSf8wYpJZHLoL+yzR2VKsOJbtj4tnxWtMzTvP5z57T2PlPg+T/3KZSY+Vpq2X4nN
ElNeeRkDo8PQYLgpQmHip4fDV7ZPiCXRB7cr+IiHNJugUCxqWWDMt76oqz7j3bwU
P7FucIYThSskhYTrMAXfdAKHCzL9z2GZrIu7zfeRLnJM077FMeAnnNtJPBLWt1HM
wx+2Jbo5gipjHgttMjfISPJBI60fqSmOKy8dSgA9z4E2e/V1oQBK68L2WwBbP77/
Mt2w9Ig/MPDitsA75TI2Jhse9/lniSdNPoWAnvrYW4/7FjGecud1L/+uM8GuThkn
u3xSgd+50UvW9t1tKB53fQj/1LPjxuvneYp24VCYub6ID5kjU/Q0z5Qobi+nWu47
3pGCdYflNyDLce2B8b2gySXnKmM8oe5LTt9Pe4JENh8Y5N5tV6qWR2C5rVFC93YC
30l+wSdk/e1Ph8LKzqmjhQ15imYyVI00BMTUpfKFGggq9NWZU4f2n7PHuqDU9BXO
61XQLMTkLeoENdiNEHmlzaP+3yqVzcf0EDtU6n3hkueEvTtKhlYjqCDcF+Pjf/D8
YMESn5ViVgUdxfqxhTtCYuTdQzlXnWXmtsCK8U/Da55BMCyRksS/DOo61v1NESag
5jijI1DDz5LxS3xGwSyJZzy4hBnqRKJ9mDXHywVdPwIIxzI2z0iV+IodqNLPFWGv
b1WP4ApEBbZLfwovnTY7K1shG05F6eXAM0nJS6Qpa3xuTeaaN5o7v1shP270T0pB
dBgSP5AVyQXUl+FyMkvnUe0B79m3rugtf0tzAEs+l1ljO/H9BLu0vUOUtAfWcgPk
qYV98GCml+eRlPAQ+tSraA+f4hJa46AGMMF15fi+wuuVyf+CSJBfil//yHavfiJ0
J+c27mVEbs07S+3ZFXP+KNOUPpNO7M08mcXbS7tKrr/o3UBodRfJLcStIl97qVJx
C2HHTDUbKQCfZi3K85zkr0OJ9kAGE1fzpUa0mclX5cpNWPnbvenpYl215ehBUxBO
68jtX8PKNBeUmn/UlreClpXXx1GVZ3W/8LWnD46YL/RU+rf+heoPZrYDOay28Dvj
Dh3XpqTlyPwgmVFnxmB11yst9VBxBORY7J9ZvZX9/VP2xm9NCzWsh6aQ2isYt05q
/rWtasAFwxBVtsB2VDvubuDoCnSVuk4pS7OJy9eBC99awn3p/NLi4LQuvt/ADJgp
ouDHKGlF4XACTeLugdfc7NL7SlagkYIRqJrXI4YbR9YBEPdEQ38VOdVfzCBf/gcn
U67OGdvN2uiAWLWcFCtsBHZBXlsjPRR4MZuzYyqpxKbUwicAhr7gAbKJDruS+L9X
yjzdIpjOyM1ZkvpFLneeKdhvmBUwZYGT+i0nKri+GnK+b1P1oM50CGHfrEr/q6GW
63Uh+GHOfUvGVb69zi9Ofnu1MU1HnS/fvHaUxh0ZMBYxQQiJuugARFmlzyvEqWUT
UiEKtorAKgqTrlxv2csG8FfIyvnkkDe6negLJbk6R/khd0PBu3mM57dzFLzQrZzZ
gLFcZMRGdEqHbtiuWSnLuYT1eNW//3eJaoIzCbzkVwTTMVJHEAH/VpQc3pa/NbGm
yzm1hW8xe65Sjag30jU/IuBRzLyHh3qzrQYEw7TE4gmGy1W4PktLofVz7wzf2ZPd
V3UChKI6aZ2e3FShV9p78OlJESbgI9XHvSmOpBEOJHUm4M4QUv62SDddvC4spO7l
JfHqz3VNbg8xstWqSdmgXuda0dxS1UCqkG504Mbtt7/a8+sGTjg4d1dYO+iy2LdJ
xYmcqufBjkxChoEkREZX/Gi5lZjQconNZl/6IOcJ0NF5TzdotINDcU3UUvzvCPDp
DrRHOnRa0PI7XMbzl41DAFlpM0JGikr9Iq/eQWHqTGehuh8fTfXAuJcXaMruaMRZ
bWz0aRowmzNF84isJ0l+ehlWyYA4sarghS0UkrdAk3KU8hQ83XRqJ4BJJXc7lBtj
g8k3f0wR4+xSVpWF2rGOnmgobieEyCYRZLXnCzXtBEYk/9JenkpSO0S3lFw153tk
trqk08zECpv4lWvPrwz4w9Zo0OPaEPwnU6QME3OlPtUqU9fG2foXJzANYKbAfh/y
vUPQjipRX2OKaQpBRGZDN2CD0QKcnuBT15FoFjhlUirjpHwI9Y+ZiA/CKGe5uova
YGAEKZBUlYNx4gvEy8Lmtu/fIgGeU35XLtmcugBhl6zchpzSn+VEpzfUshut+HhH
9giQvPOleKEP5xOwTuzQeiVGDASyZbLpAWPGaTJ1/9KexcRe4w0QstOBZJIaHo8t
hUnghAEZh/i82Z4ZLew3p4bYhbjw/5EdUDfZwya1kmgRbRe8d2lYAYMHQFIOtfGh
i0Obl+4ZQoV2wCnEDJwAtcIx/Mz2JVnY3XhoP3mLamWo4F2if3BW6bZ0GAkYjyCE
hQJL31penO8TKB7aN3iOYehVDBmO2Y52k2jAunC8g9mLKwnv9cqDjlQLDCIfeYc6
ehSmviy+ZhbLUWdOSiGXQAFvejmNYqFnx+IxyMDWxYAv+LhneMsD+cYy4jUOoFjC
DWrnajdZ3Ugsp+PZ9rDLgmqoEDRThvDL6qj953lMgG6r9IcmAp5JzxVafHJ315aQ
sDcVVABBsVnAN83E7wAf+WvTnQoybqDtY9NlW0qoGCtuxlvf6OFbfuG9KMi0ngLz
w1JUC7hsuVesWO13NQ0e9JXmq8AfoJqwLSPTyAi/Xsd6/GMaST1XZnc52lUS6pew
09i3nMY/dBowSeSJF4gT22UvHG9HZVjRC1TpdM/0HDS46t6465CoH6MNIOlQLC25
VAcKXJvZF04kFzYt0KCK3Ifzj3IsDIiOWt1Mm8hCmCRZ24m3h/BMAP7i8Gj3PcVu
d1S60D1C8SRRJUJuAMz2RV42TN4Qniu7ZCkc8iLx8D4GS+D93y8BW9jchUjt0GYs
4P2Z6pR6TA+Vfv8xhS/8TXefE5aokBzP5BZWcFu4rs+OOF7xkn2eRVeOEIvS4c37
ubZfG/oWzkahQ0L1qrSZ3vl8I1KdWSx5BYu53EUGshhUOvp8jBUn8QR5ef2hBCt3
PwvPMzzd5YPd77ygaZx7vr7NRl6Cyg3IrT22sNnbyUMiNC4Dls96eZbwqUbgORYl
Ui3GK3p3NMFL9i4sInSBgL6jhXmAYTkJ2LZZyl0qVX4pZF0zOfp5fnDbfRckBYrc
rQQIynsbpb9nU6v7xhpoMS1ZtQLZiEsKW7ZauFdG55JY46BLRDllqiipXk4a4mDv
9WBJdwgK4pGvVTMQGXyVuVbTXU1omxh4ZFxbPPfOFX9Nx0kq9aPc7LB+XQWYuF5n
oBIcG/F138M0C9Xi7aY6OQoJL6lpI+Il/ITdXki2fDgCkG61SnOTJr4LOdCaCar4
ssYQ63Rnx3DU5LkKjZwOWIngnLW25UHFFf88r8mK5nCFKYkLkBJZSyUXnUpL42qD
fZUEOd+uLnNX22sd24tnQb2o03lUbUe4jDFcMNLouPbE3u7hFEOP9ChNVSYIPV3e
lzVbNIlB207TaFdTCmz16DfdMLWCn+oLNs3HxxStU5N+RtHXXU8aeuSStT2yM6iQ
lOH8hQTwIUy7AdtKq0OMDmiva2T/UpcUVHxHcbtZy8iD1feVhi/BrfKIIiP4t5kP
uk8NjXLPlNKdqIMtMD0mriLbvxMPdkkP7Ip5CYQMCx3ncRD6sQkp7auHEdvlOz6U
1EmCyv2i5AtHnJaiWdwXjbX7NEOhnVV7WY2fVPYInmcXdFilnwvrlPBZ5X7VOBrO
gncVriYE2xHJKTe5YnmzXKKXjMJYbZxQn/pRSf29Jq61K4KhOltSetV7TjRwMdyo
BZJncQskTGwWuMM9kIyDx7MA6LQHYNOJuIeonyaxFN8o52KVo6M0U/ee28LP67g/
TZEGjRLmRvkaGelfVQQVRLkQU6yxmWiqNJwJG6ZCBvt9XawBBIjGRNpX4SfvR/Zo
/1ybultaiSX+izLHZGPawy4b5BHZ8XhZ/fDJxiK200FcuRMaUqzCk/DiF6RtD8IU
4a462beaa3Yj6au59xou68CCXQERDa5PBAJYaGru9mIUr9beblroBBG7OfwSSt9Y
6pm6hMYbtwGQf0QZ1sSGQ/gIjO8rueA9R23mJ/MYTzgBhfnROcM1vznVyjrfJNob
BHzi43ElOM5LNZJOIYf6qmYujcCI62zL0bQ61pzuLjJextAIe5MhlCy6Z/HwRMw1
XzgyZXlv64WT5MfFQJQwH2XkQxsTM9+X76dNM8kkcjhVbeIYuxXmF+l2SD6T+Hlo
HlJ6tISvJa2nWSCbcH/7Ye5wg7toD9ktwuROmZ5EiIA6rJy3l1XTLxUjlrl3+joc
uKmSQu1qFGZnagOdjVKqW5si+SL31IP6YSyAgkHqh1xu6MlgDB0yNjpOs5kdlmoV
kV420/e0scBokeBSiuMRrWSFYvUceXqmmQelhHIPU41a8d7kdAJR8HTtkWiRKXXr
zMb/Bf2G29C6ycQpYpBJhT/Tcrb91M+Oauh85FmgQhNRaaFMdR5pBvIGnbGGWVTP
hrjvh7wogrw7cYr8P6TQuxe83hcLV+ByHzbxwC8cAiGgwdE8fNC1q9GJl6OF/3Wr
/QB7JRTor7DYx97hC+tgi0gYHnGB3nL5Vd75QDUSXc5PW9cb8RNYleUNJsjTL6AH
KAHDEAFLh6Td9V/i74y9s4AfDy7LBP8uw186fyuadIVad4iqXo0Ple1dPvu4QY3/
kzIqZkFTpczHun0PEAfMmIMr9CIs3ltN/8JP8oDSb3sXjAy1aWBvF6JXF3OwfDDq
17EX5oXymnowQ1bZFL5OSW2nWQHhpbowLTU29+TyQjiwuIx26Vg+78AC2ruqfIYA
pZ4eTx644NLSIDu0nMqdHvFc3Ey5wQD+3gxfvVTsx/Ri9We4z8T+Ad1Xj/envFRy
JwjHCVaHWEGgMX0Je8WNkJEjampaXknvU2Z2C4i/Uc79V8wBP2Ocv4w2O3/keZE/
5FSzOVdtD3M3Spc1pb+1vvSxN6YVrs8es6FMMv9mxApKYV2o74EEflkmXZrRm8PD
jOQOg5Wvlxu/ZiWCtSwYa6551OzMBIuzqFEcs5Fpg2CiV7bNQYHMQunSd8Pnrb2d
mRQe1qPUfafkGhB7ma89TVWYqho9fDu1i1QLkOeA4H84R/Ee7Bx1SkhQleoEhTLY
1gAPN3Bg6Nh69SggWgRnJtkHokbEHrHRwRWLgW4d1ussIRmvLkldFqX+cxmpL95z
o7AH5rFa98p/GI/hKNuUTcn8npsJOTM6VbiOO1J2tntdJ6bxJmCuxz+idmVYPeOu
5Y/mA8AwGFH/xL+zScwyc6apDD+scRPPgx/KiVL1O/VllvgEGkEN0u7dcIQLazj6
VkCnllAqntuX0GM0iPXVszw6hcz8T/+nPWlYPDZEvNFDcrjVrvpKHwVo6GCsNH++
2zgfLOjQWKg/S0yZhI1PhZuHa7KQDLQYn8LH9Cumoav8YxfPEbYZsAF+Pea03qJ/
2YqeDUeHfbZ2ocEIFN9YbtDOb2N3QlobiXrzOxuNmdnZONynqEb2AwLN2ftUM15K
MJ9foFJ/QG/hCWOM+JUyn4nG/qproTNaDS/Rmz4rlEVAbEuSqZyEw77oZK2TSCLp
uzMbPiZluz609f+MehR+kiKWGcnSGDl+XJkFYEDJba+p/3kqqkKnNZo2XxVuOLGg
RdYOSOvxTtwjf0aoaI3GTViOSL2lUpBYgzEgKvQEAQ+A+txpOkkWlrsdAkGkzEiE
qlYV8NhrGvPm+aJQJ3mbw6MMNlPnaqxyKht/kOzV0XX2KYZ/gM5McKxQz30fKgMw
2Fy6F3mYsxGIJkbihP9Ff9OJPkRtFiONeDSFZrtGXbaX+cmDdynwgS4hyYD+5fHk
uWrcWTm7WaG6FWh+6oZuCPqzLVBn4bR7RqTwbBfANf5DD1mB3vyGTpR/Uous4JdP
Hlod8KVaI7SZ5qXEhxxM494oKVaeFZnJJrCdE/9CN1gr0UgAGHxEygZWzS//xm7X
kSC/Tbo5ie/eFpAM/MFZZMz6fsVu6A8CnTbwYe4lt/eVXjw5fljAnlLAiyKy6I+c
g6513/CRz6pmblqs0Xq4zwUAU5N1SIF3xCZPaZvJmHeGwNmxgCTVhmchiHn1ykbv
NqNkMY7tpW0CrGr39hVMwkahbBsHVFURaPLsCTU51RWnqjBakIg1lqe1i4Cemb85
yCgPo89iQ2nKa/9ssFGp8E1oNUBmUU46Acf8j+faY6Sggtkj8VxFlfJMjja3NZ/n
ebn9kS95BiKFQtTyRO1LYdRoqNnrR1DwQL/Hh8kVJg2tdkXG9NJMeGb2jLx7yO0q
4dlH9/lBzPG0pEW02mIqb1UdG1MQ75XQh3jJYRrnXmODJaqxCgk5N0EwWJh3162s
Zhc82cso7p0L2jIYWI3zyPbuRfnzPjrkAYBSuLmiwIXXRf5Z4yz/PSnIMV8FxbxX
PkjblZREyckZdQHoSYrbh8trw8NR7wXugFHEnBKPnUG+E42zXFRva5OitF6FGRqx
Fh8SlSiHhYNDB8fsfqeSl6l/1eK99zouI+rTB5em7m0QnlCcb69uI70fNuptb14W
fuSugl2FVpVBp+Wg1k+ptObr/VevJybINRt3rP9jqysBpLe36PnUdFjTudS6QKo2
4aN/blnqJ05Teb5T9IzbOtofs6fWNknCQw2JX6UrM8n1EVtbVZgKaFoHcD5GvLxo
b4z+RGi0Td8XtfO8GrofBOW5xtfZZ6kjBrhqr2e4KFs4fnJcGm3UKKdKE+ynZRB1
7tXQWXIpUfiYJ/PQqIYvmClkg2+uRKuWsm4Mu1ur66pNRtTLE3buPzCpp7Hnn1tv
tYH1XMqMrjGzX+pxZDmpXXrBbkt3Epnthf/PhNCzIJV0VlI/8DJBcZR4t4Br94nF
y4C9npHG1sGe8d19W4ctAq8Rc8KXACB4I5/MYvyHS3kDJ9NNJ5Au5YG9yr+WeFV7
qVixpv0w4Ok455TzxIVIpOkGiOxM2Eyzr8foGg1yJoFmlR0Lu5ZE0gNOqo4DCjz6
GMYXcPbYwjOxTvx5syCZ5eN+O4YnE3jQvoLRVnC6Wtn1yOaw6yWUO/w6d0E5BcPy
1nf1wMYxPjcgB7YYHHJtPdMd1exZZ1i/fH39pcdiQAgjqzQWJSbLeH+qaar0HtN6
aRN9k+KHpk+rbMPkALOhwd/sQI9qY0wFgkLVoi7Sw/tiq5NXQia6yfOeRtYlbqps
fYYP+7CefB732DF3svff8VhGqnvdGFo8PsKZd0NbC8gua/AeJ6rz9AKG13gl8wRg
pRpEsD+rD6SQiYeMqlwW7jCnWnmBnIp4OMQpwxz54OjKeAHJMCQLK0IfQtz7ujHe
jlgZ2FjwawJinsIj80JBvmnbvQpjTMX8Nh4Rb2eUW3SM+q2rpvAUePVbdhEzmQIA
CuUDa16lx8yRGP7tIC7ltbPrybH6HxhlNpFHWhGRqRxj4ccCRYyOwSzDCaOzkaGO
shvaUi03mXGT1kh1Hrb3pTOPuoSlh85SIyWRK9z5o5cMFZHpAFcgOvtPvz47sOaO
aKTYYR2mPakmHvdERntzcdWfPbqQQaUQNZ8DqPh8xMHI4IKDzMcHz7M7N84eRGpQ
/v/OnbV/E9U1k1F/DjAK91/djP144hcDAVHZSXftDK0/JTP8hF4tNKoKyK5mcPU5
T7XQE7C/4smBQXH6nYykM+Dh6HKH+Xlu96BTcUY2QbjcCcrb9LAJLG/Cn/6RJc+Z
cBrp3LZIujFMwGpezOW4iw1LTBr1MSgViLgyNcYV2f6tCt079G/QoqJXFY4jOQsv
ruka3mZIHpJM7yIaUtta/CrIc44NybVUNN94U922DYL9ZtzTZAvCfJEeWgNgHjXD
zLIxtmHyoKi5TS8Q0kLtUWDYzQzQKAUJjIgJBPcDV34LgO1U3vj6AN2eNz1KJvx+
Ur0mSZeddOcAVHYW+Vy4ujjHa1Vi2tEzQrr4gf85AyQt9ohnthWQe0qT1xcu1nI7
ahWsOlCAsB6YGODZypDc0sYnD+CjNxYmO0qD1iQEXiPe391I+cvzP+RfHxs8IkhI
nZeH1ewLR3cL7qRugSMsMxiiVZKt1sxWRE7DccjfKA4aZZcRqW5m3PAeZJyVO4cc
yuDHs6RvQzcP5DHab0EmBxGXuF6ifaey3T9kvD2wP/yv1Eq/pST2NYAvPU8jGmWu
t7eXgbHXNn37eHvLu+lZhr+MqRKIZI8Y+iKlXewiRz02YrkLT2YfafHnF8tOkA5+
4AbEUuZg6wRuMq/Pb61I3I7fY+xXDUANZQt8nF8zDp7Xj6CfVA4mfH5yN21ogywj
jkTamEtHIgwQj/Ab0iVejnOqdI3nMBEx/PvgZ9QJnczOJJXuoLxTO10+lGDNTn6w
rZhB9StMyR9Vzim7YsLZ30D2eeyAZSPDBAWPAUXK50ocDBcjHAZg8mmbEXMkjnCM
+dfKk08qGpVvtWdIxDXjg0A1YQLaafYpPDQ/bXcl8cIrcJ9Kl8lOvCqit8pk7pBr
Tgy5Xa0XO4fdGCQ8nGpJqqX1mcDxc1RJ2yvHgdNkZN1tSagLLWgoSdC+tv52PQW1
YykqQ8X91hxyXUcUtUxwUjA/1LK35NivNUg/gKfd2YUIJSYsxPMScA6UeRMsGxyJ
CGUkkY/1/suQzEr0/l3mCzP+1ajaSoUX4DF9fszt8gcWxSQ99g7IYKmifNXcUnDe
zZvTOLSLNYzEArrxZdZmNnGF5slLQp7eBvvu0dyqI3QcDqXjcHIjwIdtG8qY404b
hGWwgwq6cNYEdF1xVbiRXltQJ4D1x78B7OF7cA5FXznlW3R1yIDgD82F54hTdUDX
lZOGZvD3o5XPVmsMCFCh6+YBk1WhlygdUcM39Q+h0uqiDkyzZpMPZJ4OM6g4Z+Gl
VXzPiyzCxpGeXa1dFu/cFsCBN3z9FhUF8/JqhxxX43Hkxa8aXVKkO2wlGJvOAOZF
TGahyQBQfMJINwGVdZgqAtRY2yQR05GWwAw/EK1s6DgMHshsCFgTjgxnbjDb3l/5
57cPJUYxokXFBpjTs4MMiuuAwai62uZxnRij8upOGLHc6jFk591F2wQVXMEBbrzY
8yYyY7ZP0h1hzjBSZ4MnMVhqHi1oTrl6ko1IInkncbe74+FYNVWpPfHYUMB526Vk
eEq/AmS7xpuKiKxp9vHo60ZV+H4cCT+Hrlte535UrtXPayi4n0Iw9SgazWVqdTDy
rZI0C7+ErLZUYSNttl+z3AdhjP8SqQbDtyR+hUgvR2JqflC5e0m5pDNKeUbMFaya
OHWyUOHP9SWn8GYaDzcyA+oDWpd3w0lrv9Wcf0oHVq+XVma/LU3N+fwPrYTcKNLA
foBKtriRtCwzCQxj+F7b5e75NRokGkdlfLjpkCmh/PAspXgAC/FJx26hB67iMHRB
ncnozf5mGX8oZ8j+0zeZjuz+taeoxw5fbBu+NSlCn6vueQLN/QpHPW6Y7Wm0P8ub
i8NflLcb0vwCPd/numc9IMSAd94AH9dMRp6ZYjcgUnajUqIznItwtCz6d0Gu/KgQ
aqU4zypLT25nmAXzGcT6yaBqKngeQSw2aSwIJaTWYEFSmahggso1A3GaBL2Cy4hA
eUIOiBrBGzeV31ScWzvw4w6xHtzpYUh3RxEWb7YBWUPdTUJqnPeq0glfFl/QTmzK
yMU+d5KudR9rQSMt3XDPhwguuPBQ56wlN5/wnvPpybssus9l1qIRT7XBD5dEp3nC
/EGb8XZMMTBtLf8EU0Q/6D8jMYjAdihhHhuVW88NZr1xcudpS6ojY3/LZpIUdQZc
342cjwhZhLj0IU5Z+/+sv8S6E1fPKL2MaNag0mVW3IsIlTKLBjtRxrnQfff6Lm08
atO/r7asT4va5M4f5wAU01+69EqA/ZctKNpZLq8YR3F8seo6Q4zqTbKr+B9cpqUy
KcxBWEznM8SE3uZoeuAJarBeEoglDJyiXHrXD7tDtzvUQWfN/xXWGZaSZUD+GW+b
gM3Yb3TRaAe6txme0bwUSzhZyBy1ueTiRkEhFlPJPw1k/QbMSZCMUHcFPiyHH/i4
eWaNNL2+TYWdvhEe/v0vfwHBspefCW0MEfIGBs61XdqlHKcd5p60Vj4XztIh6Jnu
3o7e7OR7pYDM2BcRo6oxjmOQvF6l8OtibeEOTn92FxOLUhOjC/QoEzMPKu8WYu6g
kiYolLx6hcUIFUhMWfkjSfHkGH9srHRKOqJRwtONHAmff6nCiMu3YZra/VR/kUjd
oTeSr2J1zJsXHKRVbkWQvncrV4JsaemfVr8jufuc85EseoK1otQ4dwjmI0dF+LO7
HDLmIMOoz0tTEapX3w6Ag/mqHjiklGlsfyFW2Lyoxi/NJTX6t3CcuyyFvXZfLRnK
UHkSFwJmK+aDXkeUbfnxFguExX9bYd8Baak6+qO/ZtQSztxJhL6PDS9ygN6c7cjP
2KJ7jy0Mr1376zAf0gWRtMzvFqHUPNxcRBQMM4tuEqQ64fS9OkrwC0jwpg1u7rrm
Mi6fxAfVkTlsuLnr9d3yQ+gN5TKFIiAfziXZCzUMxke8u3rJawQq43YWaj5HnfH9
2U6Vcj9SiOA+FvY98Xvk38nB03YLZfm/XV5TlgGRuShQ8mHylB2AemOhIm/F/o/Y
I5RwiIWPyxy56cQoJlS3vLzElvXzOfwyuajWZbdhERmaltPshnr8ndhMTGWiwcFd
VzxieWbCO2zmvlu3R8f5cYc0deYBFVwpIE8Ozj9WuDhwc8kSghfgr6ovVl3ttsw8
JNEmz1VpllekdSx9btpJSVMJhelZN86ap3ZFSPnVSgfCn5R0Mf9eonz1TmkS0xVf
xOrtVbU3g5+xxJpmoqFe7EiHXbMVg4jpxTrXnZAtWp5oLyhRh3eSuMl0jViXRslZ
iVRPhhnY4OKhpkBJnoTvF0eObREC8iuHku68E7pcpZoHhqswEGHHuS9cE+KQB8d/
yvuHDhxSDZ7XYdiu6T0PZXv3sPouhhlQRJM4BdcpLf4pJ9vgMGiR+4o+mRR/BuUp
TzPa7WxZQltdEmukuI2Tcj//B4tycGkKwHWl0f9g3ZC9/mfJncUd6sEFutG1FFYs
WIuRxCOKBCfoK/ZEEA5T/xp09vAO1GwyukTQMtpfM5qxHofSfFzAkVPH1mzl9se1
CjDu0U/qjorVvGVIaZOgEPCqwRcLd3Slw15KtQ5HfPI5rQ4hR3IMO+z9ugFFjA9q
84Z8loAN1WxD6l9dslshcl87L7IxOGfzk/fbBmMJJ02xzGDW91ywv30SLFr8qUYd
MfZdah3jAaAjhTNfDWxjpm1dLxDkbxFdqEOdBpcbk3j2KZE4oBXsqHxrAF5OFvLe
A3YARwl9DXUEJicg89iXOPLjqUw62bYTgSUMXOPpt0vWwdJ4piUaEPgVX2U+Z36K
6o3tV91utOsFYvm98Cj1zKSGIQcElTaaTzkzt9iJYDJbzHONq/tEg3r8fm5PJIV4
2QBV1WPs91p8KZRCePTXsU+R1iuE04uTVFgiGeGBGV4EpyAt65UhSooPe+/kfbzg
wIQkFnpIFL/QRnlsO3yzLbTyNKzeZiouNQ5JT83b0CexZ7mIF79oycdJO7iyIi1g
YMA+Qo4LR4G4K/BS9qI6SJNuZQdEtabTz+YLAjPRhjEk5crisnHn62psn8GR+/da
6RQ5pCUd86JZcCjqjlbpvbwo8DJRDhS6WZqgF5z+u0K9Wdk+SXekPYC93v2wMd0M
f0tuxXk0Dap/7iZFcZXkj2Pilv4hnBhW7mHsHILbDnv//ZezTrCnZ6uBrl/SBxwU
QLbB862cBMWds2JOsHcWhmgTV7JBWiWATCTYXmuGYjtcjPGUem6XnMbVLlr82dGR
x/q+SC0mBAXUZtl+QT0qxfuWV7rCDvNyx8HszEFeUnlOJFCWIX+drzrbCZGYmZOR
3cX9NQVp15O270jq/eyLfXzay+4igb148B8i7aAFCqL1swODtTWTmzQIU/c9vz3Y
hxQbXpTcjuj35IcV/OtlCRo4xmzU5KDmoKWGPInqlYx4Nxs6R41dY76phEYEZIPj
+uClbgsAavl9pH5i0FUU/mNmRTZxfma122L1gr1sXtGXWKO7Ch1isyJgzk+zUINn
NZ4bgEzKDXLRytqOmv6TF+Wvzmo0gYvxL21RfYg7E9TJle5u4qHUEwzJsB6FWAM6
GFT/2DoY0MT/9rsQjKaXFAUnrzrvWxBA5dXAKVYaUHWxC7FxEkSRa68gCF07D/FS
QXAwFc7HEXVfGGanf7beZqmnD4rpdWxZYsKa1/VLNAyivihfDK86BlGLPq700VQa
EvtGbSYhsG9fBsse0f4GGSJE5SkVBssfjThGCGlkwFkOCTRab6e0TluoGjJw/YUW
m15/T4qQVarU9Tsob4QCRN30Lp+vawRhYUlqskz5i6XfxxY5O3HsJ9LpbOvmvbSX
GpwCg6rNP6jSCDIBV4NubPOOr6TFKgz4k+N0cf6RCK5IHvylsFhhEj4BHHddo7HE
whaHTkU154E5y/lMwEkXyRf4IqpssijN5/vGPw4YorpOzI25JKVTNuDYdfuox8wU
dfK9N0xnTsZa/mHAZVU/VKRypE/lqF2lHp6wKFw1EBkP/kHseQ0FMPaYjNS+mXsr
fGm+jTNVNJ9VDAYdqHI8bfNSdJ7H5sdgjTfgVMeUTc73Q4KzqaEtQh3f9/xEGbvp
UH4ofta9ySNLxCLma4Um/HcAEEIYBrEjBC8I8EgdzRH2qeRbrC4PPw+w3B8WblNE
CljhnFH0C6trKOKgwvofaWywwqxmmTTHSqdMkqB6iW1mm1umG/WSiQRptjf9SgUI
ZRo38BDkUNQCmhWOqzIPO7bZdsDCaysr+P0yeXL5Z4Io9qP/yUnKfGGGT3Hsg0Vp
P77oUaA2JvNMpuxKqkB3o23xuxFSMW6sDxZEiHayEiOkwRy+sEhAK3K3dbZtelKE
UyodamB8YIuy75RdgQmDuiHN432GomudlRFHCbj9sAgyCcyHMDs6eXtjmCEk0OaT
oOqscE5SrhQu2b3PNM8BqazyZD9/vENJ/SgVq9GItjwRIC3En/s0Q44/5QL8Kqxo
WHrGx6u2PEAjHPsWykYCUgzAoS1j4rdzT2wECEeX8iLfHjbqZ8qqzYS8A4BwsZm+
Sb+iF58+N13v+TuWFlYbyzPsEd+xCL2zrkDMzepgotb4dHSrPwYFW/ussJC5JlOQ
uuJZU1m8gNxTYabFWOWwQCYTDKXPZndCbhJzdOdel2+mIZMldTQTkbPdnFy7crYd
E1ocyBF1EXtvKN7oYbHPTDoNO9WShtc5q8/Tw/pBxf6b+zUq5Rwv+oDy6Zvcf8SQ
1yOxK4M7GAbZF2eXNMaU8eiFKgD1jkVXZgYsG80qrgjcI3b3kg0rxFKZgS4DQ7jQ
11W9GlRLe0nrYgvGIXnS6pVig+vPuyYjggHZwUkQlHS6OEciJQStP7QWMAz/xh0N
COUb/qmE5khxa6H16zvXX6kjRPxIi3HHcrx3nTkrFKkuEI8187H3jdDDsMPMaOhS
bfiTQVO5fzq5HvIJbc93bi1d7TYOsqsdzbEAsLL5+0ENrBlAWWH4CSZB1VT+VDkW
IZXQw2Plq6q3KvzJtkj2Oau8xuOrX/50a4U3lD7A9x4Y0aneYJsujl8xcMsJPsth
6oR0jgTDc1qIlnnmuTOJHZSFBssihBTju/5+zt/BvyCUpxyx1Arg0pokGB65U+lD
7XQA6cTswh6tM3wQZHE1ACsraD4RBaOb0AinQRxK4qwfANtpX5QQkqjmGO5Q2KLa
1aiRb4mwBa+PLnRDc53enkeDg2mWKQ0yupgUa+vTW24+09QBLdApdV2Z67d+Mthy
oXHQyS51WWObgthEt39WixBXhes6M1QJSEeyiEc5h9/TdCFrYeuXjPwXj67wuSKe
lbHp8Um4dkPr3tkYyDDrN7f7RPVRZe8J1WEmt78V5RsYErL5tI4Vh6dy+WMNLkJp
USLGdU3ewaCsmcRRRtak+YAkR2fXsdcXuE9tDee9szEVPXC94iKYedZz/vaPwAQq
JgVxn7FhPq19SkJ0OyYAqeyM1P2FvQCUJACkxQorIqBdoZtv1Cg7sVuJ9qm9CWx0
qq4s6ZB25Df6mb7+NBKlDDcjpcq9qvxs/54VDS260Nv1KqSHlYFT+kZyXyFZw9a6
S2yOb3FWLP9CEHRjabI2pGyv9FPqXZyASTaj+4a285x0sI0ypf4DtuUFwmveHHhh
iakf5neK2Oh2qNIuO6sTjJXj8WXMAMD94dXxPUdprV3ihdPA5UPgmZtOJFA/yO/A
eop9PsQHHBGDD/Rwq1f6mZ6B5y28MRCTylC3K1a8Yvepbq+zo18b2+LP1kKeV20z
Gc+d2seZgzY3H6NKvcjNB36F/SwIt8F6pko2Mu3nFXYCc9rWLdRM6Kih5zWbr0hH
0G2veves73iExWCeiT/rLYdE9Uw0WNc1xqyUHlgssY8NzqaGaWyBRQhwnVFWUorB
qG7erkoz/KOF54IiXUUIbDddXXRJP2OPuUWna/VP0S9466Kc1RKU3p00m+Y6/NVp
m8uYCJLdOPGSaYKX7+uCGBC0oW6fB0+lUHewBUPZgamWFIin78Qkzw11dTuz9lLn
B8lRPC1bpk1nNBy8j6vh6QfZYYPpr8A+f/DrRnF/QDm+NdvABYJbvw60c9CAwnbq
F5cYe2nCSFsor4RbApvgIu9DT1fjiUm/FzLpEIi8jaK9uqdbMeZsCVZleFta3+7r
Zm1/kct+LYQldBQ2R9u6rqRWd8Mo3iOIfQaZ130ctT0IsA35YyEV5dQzjwKgzflF
I249V3vOG8jmgPBNbchpaS7K5VPFyGFkVwDJUNnV+p2hkXfUpwOEa4ByNkQfyQYg
CsTTUPDhftngbY3MmlUOeimdj4rkTM/+uZHzOarFnErHE1alVwp7FsTrGO4rMyrU
hlTdQtk2VWGEjeB0nXNOjCf3iFS69jJ3UUtJZstYJVlB4HBjLY3YCVl1UZjTSCJv
F6GI+3P6icRyfvejFIBJ5+ZKiEg6R4FdonbSZUhgVNX0O2bYZWEYxGUO2/+e+Ssi
uNqriy/vDajGt0bOiGKtsSc8fq7cP+Il28/cWvsuqCxswIPf5ciMa4lrMc/w6zLS
x+mbLvWTsurtVlUK2jHwt8h0lE63uY9TyvGkl9vvuBrAGsuHM99a83b8+bP0dKl6
/jSY7d0iAEkF+Y4CJx1DUkjUqvHFDHzIrqStNoezFr3uxO9G7LyE6q3p5Y3Ely4Z
xybaUum4HykmIEBao5+D8rdsSBwoyCbjyTK98n44maBXrW8xsacGIj+DCwYaefeO
otmEDgXckgTLJpyrt8/UFbX6EOzLbM83XXyGpKzZaEFR8l/7b2fjLltpxls7XZPs
K/VpfBLRP+yothBwA+QWernMJ5fxrfRKX95PoINKKWuTgKtEVFhxJAL8GqvfI3dT
ZgiqfOHGJLO3dAcIT1o1AiJN9GiAUGpeO4S71jM5nf9bX3i6gnXMf84/A69yYHNH
TmnbeoexfSNEQQyxiuKP8pTO4nsEUbvMci6LLrKwzJIMWWshf/e4pQMkjBK1B6ZB
Bexa3cM8QMROYSiGwE+pjW3IMzsIDB/0ia/Fvxia6U/SjVg/mwvFQl/XRk72yMXK
mTbZ+8tOBrGcEy42ncVwmfXCWX62nXPsgNV/IxkE3ZzdpZjV4reQK7GrIavCwNQe
7YEolemY6/73MwIxqaBcrrKOdd9E+TtdH9KLWH2B3EQ838jyc4YZln9EvHW6M4wU
aH/HjGTXgqu4wK6w/lIx1+ZG/Setn2D3afh7flQ+Vgl2Me57jHvOGz1BEdUCrWjA
aYgF0fuAZ7EnBchDz0iDSJV3NWYOlTdoJIIdUPIARLYFlNhozWUrfDXwZSQbKTim
P0TkfpBowF0WctJ8nm94CxBCi+6uK7WwZ0t0BlhiQQq8o6u5RUB21aXg740R+hgY
dXk+3SO/y7GmpIjZtXNU3GLyBnAigvjbHGO9uBH9WyEQAl4BijSRTMKGx3m/DCPj
nH6A5FeOi+Ath0OBthhDmqp7CyxB7pC5TePN/AeiCKjSUAroBb9XTwuSl/2+MdA8
JkeFN+uewcf5wDTaA3zUECEM8WTDvqdWYkWRg35PPvPr9rob/GSCxI2NetxAhuRh
6vggX6UHjATNHWAZ0s2FlwV+AGNu3AIQ6bTe3iGnUWJ9u20l86z2tGRwHeNgv3br
mLFL+162pY5uAcqF5gYGsSvFOz3aAUGTMSpqCf84sXXh64Nn32S8kGyAE4I9yIvB
P0+QGjcCRx2aPhk98nQECwaXzCzTgTcpfKhQXgzlr2UlztvHI1IBPGWt/+DGJeLa
AoxL5ti9zgF4OvWPJEXuJEQy6lfhj6zWfL//6IUwpqk5LrFHxGWXX6S+5f6izwed
ibqKIJ1OYWDHiuI7kVcqRCbAWXZmG2dtieGbfdHJYKaX8bXYx3e6s17/cJbwYrKf
p+yA+HLf5UvoDUYAekTVmFQ68XIXx2Rhns6dlkypLDzg7FzpYZIi3AZ2UqlKYtly
LZa+LRGinKNDk8z8PiI7V/E+0/uFQuqI2T1tRvwc+4Xjcmv7trc4I3/mpq3ep7aO
MEVqyvS8QXZIbCf3i60RtwE1oCm4yV+clcqVDhqI1rA3PriUD0NyWb3X8S+mXrCc
gz54PkdMCncEuCAsnmd7jJ26M5Mr2+cqFOqjJRBkMd5T/qfqPQ6e5/FXS+Mt0n8v
DYyFmjAhhlzPsiReLztAFxI24ZV34eg2IqETsSe84MrUyN0OJ/z8i2b7XhoMPv3q
zdjccCnxIqOnEJ0tj8e2p8KU1lKyl82O0exIzWPgQVaA8FQ7/Y25xMVVtdFtrP5g
0WwqG9M+EIfNGENXC8RJRb/SnU7xH3Tmdx/c04ToSsn3u4nYLJjgRWw9levpOSfZ
YKzwGL8MWF0DT9fCfU9jyfbzyGuUud4pS6h/hNMUz0BgHbsmKwFSWKv/YXAHTcDb
nXw8o1KJeBQ3KjD9S74qhY7qbOdnVyOGrhkARoIA0tK0jNVOi5nyi4Qni9RQmpoU
aKxYSIV/X6dqGziUmoeImCDm9f0vIamvd7S5K9A/5mzXVD7e02T2mbdRf3NBzjIG
uA5Ze7GQ4FaROxOOCXvJ7aG1/+2Imdx7jM+2qAlEccH5Bfu0+oOZDj6KiAzuFyis
XNsYNmBy7+vfDKSTdLEOwYFByZ6vJyRJHfiao9N8D34MNK0wky1GH9v2RDy005tu
hs9lvb5LECiufI9M0ZXIVCrqia0LTjCNWYfQArWtLMJxLjP5M2EClFuwD3AXimq5
D6Embu7ZKRUshrXfjadp6+LrWvto7yxyDinORcMu9VEX5Gw/5wSdl14Cqdadi9hY
SxqqhsXGDA/NO0J0PyYY3vKSId0804WUW9wOak3aoLSWdBOyuGNMIU0UTOT5QeWB
MLFr1gkJXFYiN3LP//4knLp1kUlAAxOpFQ1cnTic8Mi4rTF2epn/icuYxGeYo3P0
esDp8pGj2UXe9V6fhp2qH/70p+kHIlg0WkzY+2b2mNQp3M0uPbsETZ+fLcNbCZL9
r3JOw47YfaPBwhjvW1lCLWW2swl+6RW4ASTk4kPSpHUgv/s9rFh6sM2+hN2X6aAX
hUSbAhzr9qgYKUk6rxaf10oHxTW+gWop+JBM7AoTc/BmBDEQUzNfmI+ECz/eFkIW
/L/+gaad+8oYwplieE9QYq+U4YXbXg0zZWQ23kzk8PHNE3UI7Iyi3SKo94ZIrq2O
IHkO5bm9mUPD3rw0VW6BFxWAbUOEgk6yhGHtl2idjD7C/jbyCArOdJjReME+32RJ
hVtXdisj34OhtaCMxjQneTbjEe/97sfaSwPVhg3BtxVCmP3ZMF68eHwQG84BuEAa
reow/1/09vtEUBJA+mEaK9DutgaawBr1BURbu/htrDVo2gAl0bP0S+l2Vm9CufBT
bLtoBcuNO19cP26mVtZff2NxNnpaWRNL+Sb+ZvS2t9HDPkIBmim2MoLUJWk+rONP
9LrcSU095tQtqogdgJpDPTWFUC2MwPD1sBe2GeDyCDRoGLzobKejK5P9Bn1EAMEG
JNNZMqgDiWy7X0ZlFIub/M59e2MOK7idvX9yPJiYAdqEEaU17JbiFdDTDjz3jhWl
n/Nvgu8S8sQtz0esNae+tfPbgFuZWr2SoYZPyylZGEYXZx6IydWR8QJ7Oejj2T6p
nC+sZEuj/OUrhGQjjZax4cxBQb1wmAb35R8oFk7/8bzIeGKHOqXhRVdofyll42wB
WZXnP3jFITxH21CXkuAT6zLnX5Q6CCZi7FEd75MtIMcxPjePKb6pyJcvGc8Jgsft
2fYT5h2FwCEk3BaFqPWChZKhuq4nRuENmhUyP2YHFSiAn8+0VcWTvGsbLz+BZUay
3cAikC5YhyyIZZ6rZSS8yRFTbcgVroGYZxzJeKug/ptaPK2Til5UJBbLgHi5T+TV
XBZ0GyJ9b+inRhPSAZ16+cIQkcNTcQ6XuHLVIFQeoO7HcQgGkzyNqjPcIZMza9am
VK1AjwrTEOeH52z9lbXpBsxUQOzeEkyDRojIUQBzJUP1nCPzqcmLCwNxLmS4pbrw
rbEwSw7DZJ54eQjEhdSpahHflPLpH1ZwIY0T/UlGD5P5szYF1NZSripTBf+V6kEI
yEGQQWDLbjrYXtE4naU7+mfXeq/kbPvHgtxXTWGmcvXLYJWvfMZ0QxX26MhLQFYh
gmS4SBEoYb+SGJt+SMOTKRz1sh6RVI0GJx9T/lLTOuYJJXt8EXuLA45WC4KGZlGT
x+z7tyClV62NLKlGxLG6OPDQKwAJLz/vN64k7lptuOTyHGFmRmfjGOgQzb85UpsX
aIztH2D1fgina02UfP3p0fuYtZl4b0ImcV1IHVJFfABLHRd6ucVUzsylPZBoND/Q
5VHXEIgJyE/SgDiug/Xg2I6bZBWA56H4T8w7FE7xNF++GP7g1JHJIB1fqW8GoEeu
m4xgTGx8bDO/p4RaS4oP0XT2HVsgnoXH/oViV5CfNjdTG0W722IaqeitS8MK/WZ/
BD0dJktUnqc3ow5GTMSrpcYVvIEGo9FAdwXHUEViK4pfJk1OorhfW0e+zLhkJV3B
pc3arjpvGM54Zr7ZxDpbpIMAp30yGKDIj5nJ9dD+px7yhLr+V+tzN6eJJAVAQhFb
u79NlX2Lxg5mVw/EGri61MCaqdUs//7flhLCcU9eIcAHPtzfm7L2dsvkbUS8ChOE
R7jqGC6ydg/Ve7sje2tdR5ao8KNAayUoiB5AVW9fk+vkS7p80AdX1GAtHOSsITf1
sySp2DFHuiDq7RniYT2Yt+Gw4tIqjIsZD7pDxfUV8+fZX+/b4EDEYPeyzye7UAIb
2NmBtmoItThshKFusinigJTwZw2kbS6izL4luwiCBEM5M3Y05e6tsTJDyR65CIWi
Jc9Cy7Z4SGPuSfeqig7ymIkgfR3wWxC4959agOifV6LC7k+Xg1MTOvU1EA5JuWW+
eQEkmxVpMot1YxgFMavzCXIOz4FdOHprhe/NQfgx1B9muik1aEX39s0eoKW3O7mQ
O91u96uZqzyMUBWi8nGcDfFl6q+3le2FEkKEVv2Gj4LymaTks1pGUGOZ9Z+jbtFp
3SA+Ik87CZ0A0M6kqL3TeTlOiBG3ox29+OflKE/nCo7Gkr5aNGbmomuiMbHnVdf4
M0o3OdqCfK8pS4aFGAoMI33nyW1SPZQ5B32o1fpM1Ikw1OrcvumSlQp05Y9p8alW
7daDSCO+/1Cae6kesOEfanC7odMOah6xIzWX78YTYfbo82jewaYKeXQ4CRlBBTap
Js2iSNREquLbJajv2kMqtOOrC0yT8nWWKG4PhU0W+CGqOVZlUUeVBWP/0HZE1TFA
a7geDG8iOPL5U6FAGbAJx2PdR4VlVE5yQKSkMc4CkefxQzTSu7cYbJis1zDqw7hV
mc6sNubRZoJhZAp4ptdTWKypYjEUtyOEG68A95pJBnfhxBKGzh6wFFhaNkeHyCOD
SHm0JkbFx2cS4rulQaTXQ9zmbFd7BrCBa6z/l6xn9U8Y/r7GbF0WZ4ptavhkygy9
VRkuB7dIyY/TAH9i36RXqXdaQXu6dm9Xt/AbZCl5puO6eFZgvJIf0Jj+13H0Cfi6
t0O9SEU/0+xgngPANLrCZ61uvvBUJBSl97f1+7RzsDJ22azm8A+QvJd1jqJqsjGh
lfbPfraLeSD1k9BLlgB+MWqHmdSv5ACLVqbnF9HZRswKbv58EeEuD5F/wExZrx17
wxTluCWEdF19YsPwG7obE71lUrxMjPreG6kPil6yf5KmrxATFy43TzT+FaVZVl9X
Xbv1y9PC8aSBtFp0FbBR/bsGpFrE8808o8hE0iN9Gm3QcWo5ChNtrdqqJyGPEUaY
G8OwnJVz4Z1qPKXhpSjKOus1qM/LoHxOsclmBuYVmfBp0TD647MZhZEE0l1PxnE6
z0eU0yw1Zr/02Y/he1Rv7OMljrruMK7kll8rCsdSTwQasFAVAjm/7K8X44bmRZyE
UHRBma8Al3m7MYpt95jYn7asmkd8BH8B0jCCf7vB30X2EYPtfPPFLl5SkFF9SIks
QjmmAJWk+fSj8iAKHtn3xN+pxlHflB6tNJ0aZmGGloLnbkyX6wtl7EuMkoHW1Pfr
7K5+Ozs8PZg0a6zVN4Pv7GS17s7Wi87YgDMuagsLwBuqA8ayiN8qdpbDiRzh+O59
63caZhl95F5+HwmGRjwxsarFwWOk/0R4wakkIi8S+8XSRCA2i+T+hgBZUsT8JECm
SqI6k+6K26Gk/YNkU13gBX4TGA3EP1+rAXi0/cC2DU7btJ1PNUK4GxWBMNv7Cq/G
HZ+yZACP+akFA94WOgfWgOOzDrvwQKoESSoO0D9HygeBNZ/3Ax83ATX/yJPAGSQO
C8nLrExK6esvroqG47o3qJPFFs+DTdU2A5+Z1Ap71nMaXBW/hXcccP5zzMb8V1T6
GOYonM99kGF6xvWSH9eA7DjOzi/WQ/I9YFmwV3nToqlfK6vdK1LYKiwRcn4o9cZr
+qhgp/VP7mwB+uQN8Z2q3C95rxaly9WRiT1rjNvG+lsyOldxLfu9DtaV0XRd19Xm
eXKVzacSnO9tZ5lVhTP0E0PT/mm3Ys24NL5yHWgUKAAQowdaLE/AFuNZ2g71Gm6B
kT2jmQZTFwJaHb/0y2cXTesJaFg6nAwh+Y4XHcWNdRvkXK6HUHYKUdPXpGopqKWy
A+jVxirCwB1IgPycM9Kp1CaN4U+gIalXQ/kbkpFAQ/I85/kfNfGU87gojRmFZwN4
sZM0i66/ZYBqQXFdCMwQXZEjYglI8Lz8CmdLvjW3WHHgRE3U06mSeoQS5YxwSq41
V/XT4Az+R5E+SOSyfBwpGLweTtfx3Sx16JfZNfkdGwhVN+zACFmixUKqw43jgEMn
q43RV+E3oPxde44vviHbtkLq7tvJsqYcMaVs+729ui5tJxi5CNXfCj5lPZzFTQ8D
xNCIIQO77Emue/cZTMCVlLDwRJeJRyBWFhwtlLr4WWp224cj1Bfh7czdeUYux9zD
yru64DPTCwplzVgnuvHsREPBXGHbNlpESq8N4xF5B4Fgws8b2s4I65PHAh4fTvQY
k9xwCgL+GQP49YE7+7N3oyGIb5Upes3PEIhOktW/yY+u/HTSIs3cR3l+6b+lVqj5
G7TMkT3C2laDyQ2a+9BR9T1Bo5ADkXXuphM2dHnyH1dpw5sEO3K0oApMxKMlhWWK
KYEpR2nGuq0YZ4mdsOmzjSA+3EACYQNkOcH8xzpqRtfO1SvmwzYEZcglCX2QnG2c
qRKaepFopkt5c/Dw+u5mV5cjB79eTOxXKPB89QyiXCqv4LSW1672QvPM+6zn3oWp
u7lNvbgnl2dy8UPSOgYh3C+odwZXbt4+r4SxIRmFU16U4Ia36jg7+a2IM4zjjdx1
bnEL3BJmkmUXjxvm+8ssxhJ0dtVg4m5EYmrZqP8ASa1RGXwYlgca/iMbcVK/aUp3
ah/p1404WvsPmJ7cVqXuGDdk2jSYpSt5TfpyN+gdelwwo6boaFv7mbv7aniR4tS3
nfoVza3x9Ckq0xCrabSxfdFkV7HMRDeAOwjoNt6okQjdFSl16fpBKnBc1Q9C3LA7
oysesfnyje8egAMOGghUZa/cW68Fgke/H6KSWNy86SOOQwTQh5jaNhUJRk3an4nH
E3MCnRXQ2et4IK0qzFJvuePY0NC94Ji1A5IZvfJJa9/Nkwacaco0R+sU/CRxHpxY
kublepTlr7IUTAuGFQzugo4gGr05WzKz5I/TBRGtxj/0bA6enRmBIENnW9Wkfo80
jJ5sUxPWMvK7AqPFbCSuzjaSOwLF1SpHGGb+NXGXJ2+gAzho/bszuwYCelSqenk8
jrzcSxLqqiQcXihWXg3JVPBfQl8HH5pC+6r2WTG2PhmZjeKfSBPoICFGf2SaEZwO
pla9dStr+Ex8s4qu+8vmg5V2EDsLFj+C9rTmEFH9Dhr1LdERjyvkJtaxtW5D8Ywe
bdoge7tzM6aLvZS6gdmGp0v6Fy43Go8pAY37j2AjhcQGzIdHRxG2x+3ANvA43vTb
l5/qjoRYadYravASqM51WanFDsKy01GPTsnhwIcrxOiQNAU5mKD11ZVf/5EaObWL
aqbCJzDrFyfIlRNI+drCLpnqmEz1xIBX7aRABZYajglX2KItiXAVzdew+Wo1Eq4a
6PnNT5SnK+4drw7JdoBrN2vlgfEbaRZiLuQfA8XlqhkCLZpUOGCh/mS2x3DjFWOq
w8Qgunf2n4OI763FlAArXj5OJitDmV63Np6Kgnkr3Z1wqi02GgIoWAQilNK81err
2BC6WqSXPBHL6vuc4mbbO7T6qw3EnMCDb20lx3JGBzuAPcUOvRVqUSxWgFGHwbE1
FuC2Onp7hGVK2MRyqj127m5euVRJW/ApMKAh4+itkwMr1rz5XfiG1IQvHzUx+pnK
VxRv3YQcNJJLa4P3ROfadYcINyvMWKRQFz+CKmHwvuogltl5KGdZZM2rALIfoWxo
WPahTgQwzJ/rjcNmDsNNnpfbRojiVlp9+vTF7O59AS/IOUBiGbzfkGytQtkIcgWv
ZZg1HT/oa94mtAhvQZq5ep17wZs+Q+0OhRvRy9uHvNIQ97/1XyIlA2UAExkIb4Kt
FFE2zGf0V3r/+vMnB9ciStq37XSWrxnLZr7vIlTYkWr3so0jJt1mGM3RpikC1Iny
3VA+0Zosza2CbHro1RGuftmN+c6RGifG+dLBNfl8TP6e34OR1vOishzQmskNtQpm
MnGICBMe8TFTO8fLsgWmVDusKeGLwQMoEK0mlQ/9/2PRgbwp1qB+B36OYCDlenxG
L1uX77NR9mbGvjuKrgTbJsNZUaBFsCaQvvUmsKRSTTb7MYySI/0GqJvWOH9eHZgb
SUKmLc82lzBEid72SYYBWJdHc8TywZpsvEfAwuDFxlo+4FfzcFiBdAZAKCIJdeqx
vHiAjOG3MBSW9xWNkmOVqoB4pqyC3q34syAvh29fTjiCJ0Yul42NIt0vGAgltI4k
g9z74f01SKgelj4k58XfREoxvViaoA2JnqgACr+/18gmVMQZ/1JI4f2X68eNE84k
CroD8puP/NPPcQflnoJ4/Km1Xhr/LisxqHzijLFAPwwiT8EhcguMqDd+hHSzNJz8
dKOHIkJSGs6GkeEt0+2rYftyrZyC9VS7UBw/LcIAmkCZHiU8ag0AAnuZk6L13x4F
c/tMhAOK7aR0bDWBtVXlsgO3N05oMrh1WFL09TQdgKCVWUBtQ9+tXIbZEsWjo+bk
K3WcCf7TF59prKdsm+Nqk8M55SGKRfidTH8zAT7UF3vHg7/MSCFCyLqfrawmUHk6
zbIH1WWJKtqTvHoOLwGIrN10MKpEZKJJAIv/JxCuYxwtYOBd9BkU7g/up6ej4Qbz
4nzxafEAMKSAq70L3D9sJXkQalfEcUTmXiBRPqKjrElB9ysZXKXw0IFc8QKZ4D7A
kWXfIuSj3qU7yNjR3vvdlNHgTbVD7pzIr/5kI91zoPs3RtLEBse3KgJCtAaP1cG0
tsj5d/PXUEpHXGk8N8pTufKYOtThxCOKpbz+NBM/QSRJsYK7K8yUyyYrVGxd0po4
Xs+WVxLp9QHgqCyWQ9RM8dZ9a/XRzu0DcrYO+eDl8Av9ilvwqDCe5HrRUw9YhWUT
jtkgVJfGwTViNI1iuKLNyDusnnVtzrvI8pCdrYYXqQe5KSieH6vD9h+SfBWkDhFO
1py40uqbx8MF6RAO0Yv234dnrGL/bsUehhbq1lf8lxglBiX0IZqeCRE6ZAIo7UGY
dTVnxVGIOhTniulI9yyjb/XJF3I1qUsHThV2wlwvj7ERshMgKZNe3A4svezZpBZL
pU9MWlY/sDZhX9FF3MHxhBOctjmFh2Cz5JNPh0xh/yTT4ZhFULgA5UGVbfcw1Onk
10T/WZsQbeKrxNO1TxzTBJkgl8g8FcjSTSpEXkcYSJNbPo1yFXji8ToujlGGHRQb
wJCBhP5xsvzqVVOARA6yhM5WcXMsrgO2ljwvE5i5s3zPaO6ioVqLX30F1tJ15Pz7
9MBtU1MrohW0f6fsh6GBBOq3pOnXASui1czVncoW9RCk0kzxk/SWWTC6rnmW/sHn
r7rx8kyQdWY3/D2y4AHmSslSHDvTPT6R4WoNKQZnCTzCX/KXkLzLmqwKcpjmNGX7
aYGUYJt0I0YSfyXjV+1oa78+ZIl5Qfh8IKbczg/Ckrb5J5KcUVYvo9M6zZDG4fzY
jpb0yfgziouWYtdR1L1ME0xQPlwEsUEKH/sKXEqERz21xw2gWi63R7tavPlUNV9G
BqhrO9d2R3QcEMryPfTH/SvtGpXRIK8gOX1hDOJ3Fza8NJdpCIc3KTx5UgxEqRiH
BvoA4V9Ys4Q2Y8kmuPN84q/NG7ERrT8lCGUWhHtZ5SoPuQjoFxZJHkHrYBBq6rR4
hYFYMLspmdFG30lNAGeHma6nkOnZyn0V/yLjhDWkuKW5dI2PQ5kSMrWM93ulceOl
FA2WPE7T2KCoZvfjgE7FImv/Nu7W2ZQeTauOaLf6qNx+ELflVcoHalIyZk9ujMij
r2GMQnO4I8s5QFqNtHfzDQPXnm7uAlmrFs8PrlAVh67ob5p+JzYWSBkLUfrV2VZI
6KbpbimnrwRTkePn5GMBggXkuawENNZCFwd+t+BdV3e8U9qA5sqAs7H0mXWfwNhZ
LbZyRTf2+dDUM6lLZzddba7tyH92AZLlGUmiPZT+cB9pGg1/yvqtBHAv6PUoGrH6
oUwilOFY61GZjNO53vmruiEbE3/JppKVZa1b0hfCjGOv3qdb+i9oxjbVPBlmNEk3
2OxHgLul70BOFHJTcBO7oJ9foqkYxIivAFQBccqBqdcnDW9tkyTR4en+1UE2BxRz
5V4kfgy9GJMUL+4WRlwwGV/23fd5DiqK4zbHl368vuFZrelQz2a7MtD0FtozuoAt
htJnb8Ay5gRO4pd5uYZMyCqsgyHvC19oQJBbdU4HgjAZt+Nosw4jrtNzPNBy+iuB
Bar/J0Gu7/ZKC+hxl88R9tzY7kWjE3hE117+ske2XMOSzIF5BvYVZcssWh8vzuR1
rEuJFRjH3p1Fm1vt3ZtgUuemkX9x8Ykw5TYSaYkq3+nt5iL9aKgmkopjh+x45dDr
OtmewX0IJnLjcPcPAGM2BDIC0ybFP/WaHXWP1/qZm6ZUQx/d02MQAw+KTvAWFrTC
2Im8ahQKPVwnsB3Wt6K8a3uUICbtsDcb20wYkfS50x0nfwGRJJQHpTZJQUP0LCNe
kZ4easp/WRGPGLc4yN9zwqV2Fd44d7UXjyldUhdqXuMH4Y3cDM+nZlRPi+USvnGh
Rpwh6qX5ian1lk72Fi6cqbTTaOXGBNWfROaWBrLrVbroTPSAPVdq2aiFit3IKVtm
TGflvmvSgUbFCjPSBdwQyGfJeSctiE6z4uP7LSEk+P/63Y3DT6LLxO5bDHAUNmqV
dkmu1OB2xJfb2hFD788MuSqZ6sBdEysZ3IVk70B/zAAVmI1euw3t+g8tSIgSr8VK
WdnB2J2+Mu7eNiQ6DuzH6+qziMA2AbhrVMKVPSjjp6dm95vG6z/TYyyMTawXxx0S
KtFCnc8oNxOMaTJtM9V0RC9/CLkGLOhBJeSLy4sq2iCNLkIScRvxMtIadVbhVRDU
AjC4gclJRCzvLtKfz7FMkfTnBzKHbd0PpveQCWx/VngnY1YkT9bjAPEZ+LtGxuPY
MEVgsryiaHrQPFn9EYjWtXpQdMHrZjyymdR6usy7HzUu28DUGvjA/EFs6BrsMOdx
l6xhwPLGpSyqv+bHVaptcsSOJSVbqnIaGW2C6ctnlLFRmDDpVIwCLK+SnPS2ufCY
B3LL5GbSk38tTB06n3R6qIkdOPcp9+0gU8zmUsVs4Cb1jr3vOI1zxD2kOxXnEgR9
agVrXwoYgRrk1jye5FO4Tlyy575O1jTuh+hKn9OKMyAUhejDZkT6gJT9RYBI33ut
XCBN7w6ubnAullaTqD5K1+Qd2+APzhModecSBxpUhbz91VuwDZkElFWZUg6HV1AM
0wAL/8yjqwDmoGIocGM88r+uiA5EgVs71DBIGsJ1pZCDXH0J2O+/uZRAD9YEI+aI
l9uzMpllGhjuoEMv5Wcla+HJisdtTqyFVF63VZJQYxYMwDdNfVMWpmGbWXzE0jCL
01efC81BkTVceAZsXCuuIP26TCRpb5rx7yGM2CDXhnz4SOLpoItersi2gzSa586L
bNo9suWEqjET7shkBAv/cNkyyHmFG/WepF1MOsXHK2mnhb90zbB4JPgAvNZslOCg
UxeNlSQNaDeK2o0y4Gv5VSvopYpXMBvOVf/nDCq2q4HhCWaDpBMWOMY8R5FvcayY
47FajVv9YcX9zLqXcEqnSpLrYwxFUV7NjrU2tBvhrCLtljqWVOeAxFb75PXlRQnF
wqFwoW9JuDpvT4KhISvvT64n4tULuN5j/t+tjFaAn4ZuyqRPgR9gBLM8t4vHLwpc
4Y5hGXx3hCLx/VBbubQfmPr1A9y9h3BW3NdgBn4UOkDsw10S7x86yysuAk/gDACR
qXWjqdHfIlTMtALJlQlmIsmcep4W19dSnO8E0DyUQMUtV6Banxvx9CUupIBGp/Io
AfBrea0Ouyix078AZssh4VbGUk7idE/CGY1Nr7eGbVcnk/xbRFXeAsRivic6dErr
FMm2m/txVKrypGGZgzh4uc6z9nrQNWvVbfpTBTdD6XLzlMjuj9mdmRqFrC2UT4kh
B6+Dt/jyYObttuJitMrvZbEYovUA5ESqC1F0nQ7c1+m64ZoLYRetZNYDR/IDwPbu
Ct0HlHTx4S/1UPhnRlmfftRpngDiYWXBUYqAfQD5jv6m/RKhR7WtHg87zygjr6vh
K8jsYVZac01Q2BphyKVbsIndl+oECZzub1FMIONlE93LoAtuQdVQh0EJohBfcc1X
TfbFCYVz5asKQV5k9lylfXbQw/8OKGiXsxnrgX85NhCqwiAiaMljqzUsNNjr3opy
jt2bzPibCDgTShhRuyIEozZmwar1y2QA2kwb8FJ+62SaIAqIfpVgyVRBxXoGS+13
lvvdWpeHXinjsRNd/tK3OftYR4E0PH9dpZNkqp87eyuY+Rq1NF4dHEZjBdpUlbrx
7JiGBsZ+ONS5F4xM+1bt4GqC66JiMI0aZ3P8iPAxP2j05cfYlT0wHzL7e0PAmfZi
FTP18SNKtGj2kq0SOl8kGuG7WLsGeZTZmrbL2H/olqjI3mUJokltZVWPqWnB3aAW
IUzqImKGaCScsqDq4K+YWLV+SP1wI8WGn83d9pdqNLEg+GwD9sWI/2H5PiS8iQt2
q8xn4P+4kGjmVFUUCIPdQ78Uv3m8mMMPUvfMSH9qTN4VEqKfdEG5iurMvNgAXXkE
Cowm64cOQ/WJTqXoUCHjtVl3ldMQ8tbQGo2yPweTUswwfZxnrDSrGVFXphv8+va6
2/Cq/l2oi0dYpJ8y94bYLgetIlFzwiNjYPnjKU8AdSRHowI9gbw8kO3jiWgY2DbC
ZYG/VQTmFOmNDSj2I1AXnOrngZ8WaXR8MmYkCZTSDjYdkxK9nVG4EHtAIgc/ofzm
rx32UGp2sbx0Im4DpkVaZcfM4xq6MyZGmzNmIb9FoqfwMgs+EN8O6GsRUA70Rd4w
V+vxjVQUTlbloesgm/N91eUdHeEl73iOXkaxf2s9Vyg8/kBouHpp/CPchSqaC4Xb
OkUMhBGHRd6fkaCWUgeGOz+WfAt8cHyMTOBsB5wdPzNbwl5HDvxAKOqoRiZ5zh27
FzlUyELMPfFDNKNwvUXsXtCm7N9QPu2GKRVA6npYg1+sNm6ZMV3HTSN43kFujnUF
0SZ22JaSq6m8VOfBHYd5qJMsgDhKssoZS6tOCwL9yLWzgGCEY0tm1GkIzUedLe1F
Zz/gc8WotkBDSoUw5rouQa7r2G3K40UOmD8/jN3hirIMuVBp9KubVrUFpBscZiTU
5MICu4SJecLjsKk2kt8pFg4qrCiXQMN24qIovV1FOgEBCylzZBJ3CedWsTO/0xH5
RPxhCswEd37PJbowrC5texN9SI+72TDrglhGhTxnaoS7yQchbc/iweY2Pa/zGqf7
5aH2OPai6t3GtGrps84WDE+PWAHhNOLveUwuZtk9ZVVSlp1rEprJGUw3pNqzq7u9
Udgp8PY0WjLJZpfSNEBEVAVebs/0Z5KIpc+D5yjgjlLKLYecYjAN7MpoyqybrW0C
5TRwNO/bgXk5j8PgCSKQ+5IxFNk1N8y4wDzQ8qiysslnCuH8PiC6li0xoaIOHYra
ZqRSTesn7+OmiyWpx69UvhieEpQ+27/pAcXteZwCenhrgPAeCOR6zUudPHVoH3jj
S12HltNuEb/Od1U/mewQEwI2EiNTXQKfE4L9AMQfTQ0kw4pcv5fTRT218PDrnD65
eBuwsj7nv8VAmy0wH9MgFsQShYAeIwfg/v1KNNGinFdF9mNOG3MJwARLPivvJNOp
i0thDQk9oeGxCQPk2xYN5arkDPnAGmjkhqq5qFt9NkLnYc4mub2CNSjXCSAr29wu
SrLbviXiwvWFxta/x6GGR4kvqVbr5UZS8MUgwkunlhjtg08YPX6RfApBGP9Z1P52
b3xNycc8MRR2I7Ac5SbdZTh9yz78/3sa9nBjYxuD2mX8yk6NgqLSKDkwPNPYb508
dYjwDAvap7NhFBAV8uaFG8WlrbKtW1rF2VLS8yDZIrlxtA5nGrHhSspGPQfpTdLq
HKIt05vu1Nl3Zh+CTbvOHm1VXlAOhH670g3qUXkzB7r8HzMazLkvxhKUXhIG/8MA
Tygffs8wzpfRk59BGfk6JSGN9lnqIvhgyrQatZ4js4P9WKFUJLE3rhCTpZuDWJ6b
Kg3L3gYOOiMgss9j3QezQqWiCrK32IF0/jXlC2eUnCBDQQPdEdRsMqcCoBgD+fiU
QBlPsUb5O7cqinUZM//E6ZpxQXYyLBCpJJ46aZMWdMa4xOwmiX0seJmSmfKAqn9p
tkq8vwsFTBj3I6vWaNSpEEMZL/6hmlehAmTmmZrslLPWMZife6g0/6TkDNta14An
2LCrzpxpgYwDS+EYW3cvAD+hmiR1hz68c4zI9XUXWluJvIvL1ILpkIqae04jFisQ
+Czr2Fg809ccxSxjqGxf5jKGkNh/MACRWuJHUcNvQlzGAWvU5uKS5BUuh3Hk2NuG
nHTTzkjdTI+HhtMFK8OZ6Z0Tp3qTPHVS7b59TsuffV3zGGedGeCEehglFack1zLU
Fy/H+sdegt3hi86JJVd/m7kJJti1qHuflQl80G8EEU4mlO9lmp7vBGyZyP24AnuS
Rc5ZdsprBUUIWpCXCJ1BXa/79wMrmF/f3Zz+aI5UJBqfdhPmjLdg4PCa4uqA+jLg
hXuoHTZ6eoUQRd/H1m/v4lXLRxD2WyfKTN5h2gHBFxyWSg3TGpqjoXf25lN1jSTA
K1/Vrd0mYZkWwgD4n/R7R+c6U4n2Hd4Ap/BFHTA51l8bawAFRZS3D+O/cg2Uaw/W
pr5rEe8WMbLY8LAA8t88EMKGP8bq/ZVCx5P2jbJYpB8wKdibBwl7jrAw5Rke2I2K
RnxSXOnzWuRdM//4rwcQ0YpFMByMoJCDn2wt5C4RJIeZ89CGYli6TU7t1esz0J++
zyq6evG1YI8ceXbqHla+ntMVbOjhIubHkRU3KJPxL7ZukWaGCe9Y4TZHQM3Nz6iu
GI8injheJp0M/rF7xqQZjopIhSEHRVUO4C+r7OrsrARnWPDsAwmEzZQkUKUm5xmt
hfpaBWsjaC1GjE4Ua0fLxRFu3nmEkg7i6b70Lc+DxW+/57FaZQo5yBjLRKzj4Klo
Zrp1dVjP0k0h702YO1Zkog+y8MOX6tdKRlBjJDWoAICgubrBs3Il8kGhB4xmXQGc
d//ya1Zy3OxESz1CsYOuTojfvSOViu0C27xU2f6fFnq7kIZyPFdcJ4nIomZK1vTa
sU5aann19yH92s11nBYvaM7rTN4k63YP0WtKQmcpuYwhaSOe1lbmtGS4TA4lVVkU
CiBHZoxNOwVuK94rGxsRwW87vDbuzSyM33bxDqRfwA1tas2hnkbY7b8J6FKFGJc9
6juW1Zhg6oxSwKLMXMK4FWCaQWipwQiTecfsSkr8bkSfF/fkkdLO+ggw5JY0SRb1
vN8L8CRLheXAHNOQ/T8nqwKQTBnV1jjoxRG/bAhT2XVvHr9GLqRQxJHdl+0PtfjG
/EddhGuTSIitEZLC0GwLYCG2lR57BZ3BvYQk51wBmZ3uudOMqvrpgM1KS0XtLlF8
sqXsoXQX8Nc63ScXCxl7OfyHZvjHTsb4Bmsx72fZ67joybVnYN3hPCkyf/mZ2mO7
vf3jBRlnrqnM5s/cDOBXHX3lSykmr3FIpvHLGAztHJk882rz72Tu47HZsrRf/hr8
1wmC5kbzM4O0ZTO1G5uaF5vh9/+m/D0l5/b3IBZjKphAIFZgiA6D3gjQgdmuoMdu
XePYE5vUj65DG+HoIjy0mFg78lp4Z2tAgrhKGH56qQA/nYHCGhtGCfnBNa+s1CXY
0qPydGZlLA72zYGTekXJbltz/RI9eIzUqovojM30M/tvGb0Y5BxMbVrbmNFKmg0X
XhnrA6mX5CB5koWDmXZDO5m97mQROPQSAIsXGAZ2a4SljccXl7t0rhSd2+JQZgfx
p6vO17DyLWH7Y1kbFAiCWDwmKZ5OIh0+VtBlhd//QNfjhGcW3+Yur4XXOzrPy99n
zzOGHiCBCIT9ZNi3fadY16UcXiZO4c6INtW347N5zc62enAuVMN0PNFj6hNQUrUk
mUh5eji0j9e+YFkhSCCk+F2Ll9F3OWXsKWbRSZsFTUSSYkK1ssOOS53ji9GvweUm
Giy8QVtkZrmtjlz2AR12o/waGAOe5SLAeT0EVujM018Obq/leMscAvSWDzimLd22
D7UaEH5YFbCxrxQYOkAljGPPzXZ4D8oRYBpEIA081FYRxmTxdNovSXLUOwDyXIvn
0X9++HbyQ0rFNL/iYjoBIMhJz1PuhTRIOpk/qjAc6YQMAKuq4dvDHH681NYPKuqo
/JVNft2N6t953WZS+EFsPEKvnr1ZVxgSmNV1xhQI0V5SFYIn80FevjgDtp7s69mG
oMCtZyHyJwst1RAG/05iJyyGRD0M9MRK4r9Ct+Sv2lsGg2AFKPU/ou/SvwqAuObd
jpzgeYZbp8ilb3bi+Szd8yiO2XQdslh4fySMK9EYL/7kztq8KLRGiQNv0bOYVDM1
Mz6ijMOGlaDKctUz/15E3YZbrqiEMiW5620Y/tbzV1hMmVdvVsbk/1rPIf1Tx89B
v+4mG0sxKTQPpDSdhcqfSxAbnV/ZivwgDaPACwul9gfaWP2r8JTs1LTz83NpTtwl
ifAlPbJh7owD7Ym0nKJyYTAZN9aEigE+8sZfRpHQfvnCHjmxhAD2nJ0OPLbQOo/8
Ddc4BiuW0ElR+4G715pOBfzZu8KyCV5sp0yPLIBd1ew+JsaLNE/HPtTfQcNMKTuy
GZYFb4oiksZCLyK9ezA8e+BxFOUTEjh8OB2U4bR6CuqQo0tEn6Htg0T+7AtLs0ML
pYozsnYMwgauxDIdFwGv9DBWpnQ+rnXnwOevBhrY739tC1sJyke7hsi2OjWlhVoQ
Zx4mNmut+OX3xfGFn1K8H8QlZoRLnvP2kYUV23SC1jTuR1X8lMv4o7dBHporAlFG
Kb4ZLSz18EYxSLev4AUp0UoIMpcd3iUf2NhM/RCJO+QDatz//6AR1AptXX8TTVTo
sz3l0FO21gXcEKG1o5ozt7HaubIgdrpe0NUlNeVc2DjCb6c60KfZbjMpGO6f2KV3
BMcVxSzgaLPTkCKtfg3WXO7lVTlO6OKQ7pjLHR4g+krNvnJImguGeULRovqh8Y55
1/66ewkZmwr54/nupnd0l2mlSAX8MvvMD9cpe0TdR+hx3udHZUhUcr59SYDQn5cX
PxX94qzM2tOrJ/eOst0N+H9vxIyHuJ9Mmau8ttunpJu5Qc8S1q2+k+yTjs/eCK+r
8a71K6ySVVHSGVmf2exUr/xMDUYlu/9Tj5I8OlphTdiCZbp5niNEAqSTDcGpBUrj
HlymXOqeZFLpK4PEc5miF6QJupjfd8akzSRJjt/eo9kbc/2MMwJmFygotpbzvNzk
Hcttt40yuTWvla7d3UoYzUoHCgzvCUhEO8aoMEhQSnXpYAnNTpGoT9nmhiQ8iM7l
fKKNV9RBqMUUrRG9y76vkah3iGiVvbcZHzlLDqihlG/PNrZuLd8C78o+MFHJhD9m
7OM8ZZjBgKbrYHSgZLaWkvSpFSCjzDrhMxW47GwBeVQCrwRUOjkofFL2Dd2ASuPd
RMDOzfb68YLNMZrNUoJQNOijGygg/frnrB3MN2MO5yMtJDBprnncgwi/VAY+/uJ9
ZwgaoHyDd9V8so29rd8s/JDNk0TidQcAxX6k1tQ51xxVuoBYxLo+21J7l+Kh/tTc
grcm7FlY6bQ1ed2pXTnTTMBlH9/J5nYmJU5HISKmlREB33AA75D/W0/eYoiglI2g
ARiJ3ZYpRlhrTgMUHpsJm4aEjgblmYe7dIKZWJaxSuhLD0XrBEVV2P897x36CO9h
0Hzj/tiZskboNxPF57Fkuc4H/6PQVYyQP0jO8c3s72vI/rvGOefE3cGYsdcY92b+
YAgM4qy0q73fdVbt41lUQxRk6lIKoMEANuGZWwslqkNHHkqCjjCXr3aucB54DYTo
vY6nVNuL8KZKedDwmJUBx2rqBR7Jtue7xObSHT9I2R1YVkrvl2+V1X5FvCS5oHGT
QfY5igM/BxOhRcSWGwEdsnH4DJQLSAcgcWACoEN9J0fJnszfqL6WVAhWwyidHn2O
RahxwBh0Os1R90lE5LNCkXTwnGa3b5bvqOzm6guj/Kf78dAm0oGN+R4ODXMZ6cLN
ajYfbmI/uoFy0hsKmJ8EV1z/zTDOul0TaBgu4rOQF2fIhhvN+XATkjiTqlpwpnkR
T+Bs+LhzL8yckuCzyx6o8WtI5CufJV72w8WNVVTY72yFimZW168xc0yU1icSNv2/
PuKKXFyU4RjaU80jgs6eAo1gzaVnXDoiSw3rDgvxf7wIWiTthy42KvJRrCo0D0Zn
7I9ZapJ+w0lZL2+6VOY3pRywA/NXZyQkLVwhDvQwA4FkUhF8nOMXOKszdgIdEN1m
6ZaCOpaixO2BMREtnW51WBu90CrXyigCSBaZ4YTFeKNxCb4EA8G/68uk4RDnp3UK
jCPQKk4mz46g9BNfl2S3WSs8e0FQEqrlAarxo05cM9uKs713KtbyzfoRZAZlIanI
OAPP05y/I++wqgkg/FD8frRLckOW9Dsh0a1hUdQ08dd6g0hAsu+U7Eu8olmAMFhr
xxmOeihKci1iZjoXKbu7KZL8K4pMI32Kt42Xt6ZCjrk173HBQbM4MUhBw77Kc2C/
quA0Pr0Y1D0dAOo0GvJVozrDSJ8+2KtsAc9kcgJt5R2idfSA1CMBw0HXxIX/E3bL
fgjtIR6jzVzNGEODzfjQhjNd/HxSIn93tcI2XZCmIhpU/ad4HpkLijw+VWSNe8VR
qpMVQnsDvcBwbgUHJsBRXl0MyawfKXamET0dkRlH5b4sOeCu7hbSb9gONabUGLSc
Jmnj4DXRuSB542te/fEyvHkb5n4APkatNd7VH9yUS9SK9m5C7ZwrGhVlQGV2f8Sm
6zph5V7hAvjIGC181tGzhr8LRQCJayiqgX/FqVHeDtznrUmcgvgmkum48WYsgy2a
OGo8ux1kL/hcNUVV6xX6b4O0boyaFwqLOJRDBA9Zg/Et0ndx6ikdtKEXxPIcRuTe
N4Nu7eaRXiW9lmUohF5CfTja3mBxYuEB3S7J2VnxLvb/7y6msR/5UHz4pVkkRF7W
ACP+NGxJD3kXEGAAAO0DuT6ERBzji1iOFCY1B9SPe1+mYEHTZIvx8B/reEKaXvvA
wLOVqeVH/GpVVxtHkqIKrF1m+TFoywiPFk3L+DdAZVoqxdjEaH/k49mA3DfsEx28
nv8MTbN8gS/H+zYFehtl5Dyf7RU3TNBCGo+UDNQI/0TUlpIssGAOh5U2ceweyrEl
wTNCfEdZMrp/dKc5tCcXKfxPUSJEaii0/LaXjnUy/EB8gVPwHcu4EmQ6fDGrfCT6
9+cFjX1ysmVHAz0XXq8E7Ll5Wy+8Ic8lPI0HJP6CosQKI54V6d4h6zRqSs/dHPbD
Q2E2bPjqn0n/NHEv1j6w5KT1XW+GT50FZp17dZ9DoNsbwk89Ty+NsZnzYblSWsya
CghvUu9s5s1wK8rlRx12qgF2snYG27jiessEi1n5cjspZzX7vIHYJQwizM9FZfr0
MUj/yLzu05XS/ZztK5G/9h1BLQeoe86hbUdpOH1qo33xkVYQ4ti1zzak+QJFc/mb
WiA8gWMUm8ytmXy9IxKqGd5DYMuwS63DMT1XvGi/HU+5yCQZIGylxEhW50ddmjru
HmOkSvWnfWlZ5ScPpC3haAdhjCzAFP3Z659X4mLqj9qThVNsZ2SjoIadzbO4qQjD
wle0Tlfmc/JBS/p/gSHeVaoKSVKWEl2CErGY3dvsrW9IgEqLE6FUuh0+4QFWvlC7
qhV9my5FDT9Mu2SGRRnyUNQpaXg2/fnYH5gtIy5MePSNa2DN15j4D4yhVew+tQOR
B55SLmoT6q/uea49yV4DKENX+iurE36sgqD9lNC63/H2BeML2DXMBFV70TGJ6fUb
cG1a0zoSZJWt20HVx66sg5jAVBk74Q/0yuVtQQVQ9tbQejYNCNbdyQhTNfOmYlFk
XPs/fPFlUL+H5cCTWNG7HWPJ2BRoMFRJ4k/yc77W3pv/P+4rzitQdaivw0iHhic7
2y48zM51sciGEPOI2moJo7CHpKbs1N0vnMHUEhdNu8LbIy1wQS0UyaLh5erfh4GT
dRzrvTVAtmrcZm/htChVTaW0l9IxvXSIULxk3vGd0j3BchYOIA19lSagSmCBgVnW
8O0oToBSropXsLK45d9UCkQfqlbRtpjDKCoUJbWKBPedz5U76lumn6/uBMcN0RWM
0dsener3XTS5iXoipdgKsfS1yn0Z2bwVTFzDDBloArLfAh1Jg6ACXcLPLf5xCoBg
xLZ3qLic3rrjkz1cLC8aZ+pMMKfA0H7YHMTFGo3XRkOfoe05Px0Htc3YMOrftpCA
QLlCr7f5+wxxG3Qp33JQ9bzwUGQOgT0lZH/7t08fE5p+pzPQGA23hiLnzL7Yz40u
8aBsm8ZlBk6wv5f62tlpIboAt3bf5eC3wdygIUyMWdEaTNYIoCmJOIlnhw6tmNT1
J4FMpG0GNOYQ9cYX/QvC+JvT/9GLzbqSmZPLncEu660q7iWIbNRH7xF8ChTkzFbq
eFM+5IcNoCc+fjkGZU06ne0uFzAoxHZ2VW3paO0wVEVQTY0VFKjf1miEdPpzAh+M
HgPnVR1MyTamuK8JaaPI5xefFT1q8Si/YkriZnJcTHXeRO5rw5UIkXrDXecJ8Sgu
czWpAR9b6SqDnIMdo8rTdfFEK2QyEWSEJAN/0Ph7QUbkVIzk8goJgTZSLRhqCtTs
5NY06c4YtMO5tnjp7qddri+ZySq5O5n+HjluF5ZGGOlR9dCU/2a3kLLxiCXtZH6/
Jm8QE/33z2aketUw/wpcXG8czSIxywhOsl8Sc/cievNzjROHEgfaxS27njk1YpBR
01vDXdkDSF1GJKPis5XJB2sV2wNVjN92qBO2BLAynRuLaFqR3Qrifgm16QcGFMzH
gbfw5VFZ1bPOcygDYJHJtrOH/QRLWaX3sg9C/4zH6ompB1yg4tc74zMPOYMpv3GS
wd0JLvvmElJzVAituLJxEjcORWD6xiCtPMt+BIyFfk8Tbowq9uG7HXE0C9KTB+ml
atM6l4MTiTiLzlPR1+rSvITIWGTZ4vnC61ZPFSo/oGyCE+LwiP9zglLwHxEDFBsR
fi065pkP7IXs6xaicrbcW/dnPyV0R5GiopAhhYih4d/b9mLlSWKY8r9oe0Cfw/WR
IHzHbik+xwMrgFvOFUV+KlLNM/jv9U+6DAtA+qrWdJqxRY1slnOCCWZy51Nm6cAK
IRgY8sSRHaTC1p0Zb0wEt5rICjypQFJPWfLPA8BVOfrQ+YgMP0lsQBsKhhawj7y3
AvU1/2TO21FhKzxjB4JtvXWDaMgD153vh5Ne4f5QuT6/mZq/pHujU+jpupdmxrmA
lD2smRVxJVyxNW+EwAPH5mQLIwNKiUUBpfEH6veNFp+YDIeZbitEzi5SnpAUEf+C
O+MviVPw0gUEjlMM0ZvkX8iTAyQLyYfiZBEpASMAPxtAAyOrIcISgcVOab7Nw297
MBNKeRbIKv85HWd4mOzeagJ0cTAoXjIfBjK3FZZuYqpJDq2oflaHzORCFHutyZfh
N6oNbBFpJ7AiQZDmV4mGy8BWCD3nSIYCpzyPcOB1TttgH87JhaiwhI06GBaEooKt
Jjmuod67DF6L+dz2rzeS2skJpA0oJsDjPNLiIRdtLCGfxA1dMcKx5bJzWy84xXkp
KUfdPi+jvYVgRijeYxU8GZnIFVpK3sv2DmFZ4t8HwaHZGzEGW9ZSf+uF2xuW76hv
3MKnBtfWK6klWcHR6rwQ9aebYILZpp5qY2pQQKy/uu9ghXUO924kRMAhCcgX7ngB
w/5f+9sGcsLNo2Em9HGK305RYX7BJutn9bPE5v2fmu5BcghdHd6g8GOfHwjLLe4g
+hDQOH2sZ3yrmElU7GZmKuigJNsXVpgtKhWDd+ss9yYqp2K8Y5hG36Riaq4M9iVq
e2Y3E/t4rPUoVDJEDNgcRDp6XzGeJY2LvWYtWtM5GP4XnkhfSWe6hWd4n09JAI/v
Y7GM2Ww6GnoA20qEChGT10mHWjON4IDIq42Sdom9DmO5cy+MKY2ivCPawsfZlg5z
364Y4qJ3o23kvsTgiJFMiCU0WnbopO62gzTZ7XCCjWEHU5W/zluqiz38594G7seR
q4lkFo7A3d4ubwfwrFpfCncLYrndSJZjAlD9C/hJaaD0K+YcIozaQsIV4PgaH0IU
taC0CbiwTGyR7LY+DVpq6QjOtTG1u2bdvl7ZwI4/HohtqYf4gqVt4R4okELJY0oH
bleQHm7Z1qtOcLalKGAJXeEgkidv02n7iF3q5G4KTSvHBODdfaGI5gBCZBaReBn5
Spo7IjxuE9SLcCUBjlOZzzjHt0VlArtYqIXJY60r+QOaVVEozqOdxK0B+N07nl+/
dkohyD5+/ZURFG5L/yyfdui/mYmw3kTT+XiK/Ut4gAb9dcpVeirtlOnIyXqc7iUS
HncXYfjTcJgovUnbmLdzkjsk9wLWZNbSIyu1jy5HOfjrt99ZScNe9a2oL5+yvBzp
QhxSrZA4XQq02lLmWxssESjgeP6zw2CJR8fNpDNvArdD0VR7+DpcSXoFE0M7R1pN
V90bbLVge3IM5A1DjZViuxny9sNuao8U5v1J5kepW4ETLfsIkfsbgkPMh4IkXEID
HUle7VGytUhNcpIM3xLCOi29vf34iE95hhD0UJM7jG0yzzjkA1UZ9Sq3xgr/8n7g
xJ5WnUIBnzYBVqqjsFd1BydXcE+oBjMU08w8qiDFUVJiDy4PY3cWndHqD+PAcSfz
bC7G5SB0l0bV2LUsAChhL1arjMTZZK/zhZobEMsEeRNtQegKbANamaiRJpSk9T6l
uz9kW3ELLWfvzFzWjSHp2MaocOKUWk7ndazEZobXtTvlk18WFP0rCaJw6CvjmUlU
8JGOktbqLGFRYwDMwGN5vp3ygrpKucRevSpbyriEIGYV+15yWfbA9f4EwzFo08WJ
n3jcO/bjuRTW1IVxwFka56VP1/H906qY3uRw20573cEsEkzF07W27K0yXU2cGv2t
PXWQCc/yIk8d2GIGNkLORA40uxu5nvlMjSqJRv3qPnqVMHpK2bI+UdypnrFslEeV
rldpU/hSuNrcGn5tHb8V5JiXvKZ2RzbGwC/1oZcW8jW5DzmZDHmY4jDwEiBhV/c3
oruoi6Ua2vw56FIy6lXKZic6tSVL+Ts40GayXF5mFB74VqbIVq4Y/ZLj61eB90MY
VrsR/qyKTl/VnsAp68ttK87IgCeldl1Z1W50tLNCt+6ogl0kcty3kFIgB75qQDj6
0m26FgSumrOCc+1t4UZ/sw48jubCqb+FDw35yWU4XqFK27kgm48FmOE41tnPAUR0
Cn9KA3dH9ljPDBI648W0naHp3uLXzOJC8W4wmI5f5pwpAQe/XcpUPH47iJ0TuQxl
pMcYYxBzTrBphQsZbCbg6jG8jij6DcVULj/ohoP93Dv3/orkzhtXMxvqizhDJV3m
i5n9PdPfbxKfBF5QayL+ic6SM+ECv+8m7Mifq1GerlDDgScmDNBEJkWK27+CvHBe
sUBezOLlKDgpPuNUn3//tuB5cPjc0e5qRIzMk438FbHWbJnE3FvGyd3nyG5IQVvY
ExPDTq0eEakEqOMs0yIkjZvANIqvyiRTCEpgsh6V2ns1uEfM+zIg5trgzoCPWQ1w
VqE8A0KqyarV+TXfa4jjncTChQaERAZjnh5Xcr9W/A5SKnORFXcTKdNGqJiyMQ/n
eHjzUxoFpneqnT5PtljS5Gvns+Qp0QLSWowuzS6ZQqHERz3xk9JmcL5NvMtSFUBD
0MGJgSd5gTfHwSJyH6njwUnpnRYZARJDS1DJxNg4H+l+E45N6e0zvIbddvcwiiCB
bezOpJ0Hf+0cbEXIdJ+o9ZfNdJAIcOKC78tswTSRVBHTCyr1GjvOsnMURm/iCwcx
vQZYhRCCQj4imMdJ7hb6DZrMSQYybdL8luLxyLP4yzzP8EsQz/RyLLqc2GZ14Elz
SzIF3utlQl5qtNM6KQ3EccqdQNMW4MGoh9ZUNu8yPHmqysqDwopOS1F1jpB19/VH
MkjKTc6+b47xDNhwX+KkYEEONQxnUbtDfoLclipb7r+s5FanM7WTLgQJJ6Cpy1Gp
IvjzgCYniIhKcXcrpwd8u0aqlg+Dqgkb3hvyBBOWenNCQ7taksCWielkCpOt3drI
Sz4dOFLE73sbHZJc7BwS+igBTTDMVTo3ylAk2+Te3aUEss5kCqSzSSHIOhScxgz1
rjb/mzL0EEafyj/1XQs9h+r+EYZQmoNHOeW0T1VdTKtiZVxUyV38vnDbvlrHp/Sp
GhrNAA5tRtcuumm3UG94Ppm21sK9w1wKFlDhev890+s2qczlsxaT4BvgEsKXzVyE
wQ6qLP3JX/deFIBdzFUoTcj3W4Vff1vxoiYyGTs5KoBS9PhaBvf5HYLRLdJq/2E4
XEELlgsE8j/GP6QA9LWaEQi3AkO2AV3dtaljXPu7lx/RYREnWAA5uc4+QTpzktxs
VhUCuIzvxzhamVjm489XndIn9r3lFrw/ph8MBjbe/yjkQ7SeK2t8duWaQcam838U
/2o3OTS9jmHFF/rSygeiOzEtZKGJke2/BiwpePQKkraw+AWtpwE4YRFTWcUE+BZM
KspKpBxfAAmi3Z/5iURsqjJE8Plk9IOGLoEItT11N0xUg/A4H8tMxBqQI5NvvHWV
2GIthf12QiH+fg2IBhlmHd911MjDH29bQUdRW1Sn43mTXIZSHIpsLEN7eht5CUOK
8Zzh5lBOlge3w2Nb+EXtMSPgldAQN9uO3QjS8C/nINVCiI4YzfFxqWeOJi+jcmCj
KSuGgpAv5If8Maxvd7BLCgNXR7GVSeByWBpTSRNCMuTQfWkXaUtaaXX4Pk1ZYm0w
YBsQCxVyw+ZIylZYVviQhf2n2F/GW9bpElCrL1mt95bOD0Mathkwq0BdTyYTotVY
KTs2xABeo9z/cpwItLdLQSryKMFKppXqIevUtauIkLFVarE2ro4HBvdCVn73F+Gq
vAQLPQImcZJrA+Olnpp+BXrnLukopOtnqIdRrQYt7fH/ERT1SreVK0vhGf79zP4D
bIltZW1JlS73e7Fn31b6N3pFeJ4xoYzWw2kA3hGBf34t/r90pDO6QUSCM58ziBui
5feppTbIjyQLqeHiRyr5S1hzjjKcJJaNXjO4N4rf7fSx33ThdIAXCQk+NPzScYYR
KvfJHkdeb5Se1bHc1eidVDmvLfo8s79X9Z14fTBHw2hSo8Z0QjYNVJSSMbsJGRgF
zsU813vjHCFuto7DkVx/J4y+PFFWVojMWjRJNCjax4HEzfYyGTRV+sE/Hp+oRn56
qzQkZqLpXKVabV/pGIAPtAEZJlNjy+C9Os92f90qUVPFvmlQnekFxsFyVB6jMsOY
V7RSaMbkbu87vXlVBfT1hsMHErKaMpepGL06/1H0kQNXd03TNIPo2cWFxkVMHL+/
zqZumVSxy74jwnF162eMmR9PcBdcsjNRBkUsyWbBot8uN+vq6uHxIuzQwchSpY+s
v+Q391dFrAXZuf8gsZFpZ3tJi6aS3pHfNMnUw+dMxSmolRBsHzcGR1CP2pSXhgPQ
KSUlmP4Ms7OAC3C8ObwuxGD885Y+qeND5kcoby8NSQNXg7Iocv3EmCL1+fkWBxid
5+JoQjjwrP50aXPFcUuoaRDWiYDodUAr4CDO8hIfXdu2j4nbqoAAIVFkUrOMdWEt
Dx1c1lziEr5i9TVv/zKeKYn49/gswSUMQMTH2j+hSuxzEvrPy8qRk169CsYeorJB
3qxU7go0oVGilIT1YfA0x1ekeUNcNArjbiFLCKPdk00x3A52mOaiXaE4IFwGO+l/
ilAD6VgtHEWMV0nktGUK8wix4nA+ejhHYYzTvPcta+8ucWS/uSpxl5WLwXKgRWs1
kJC3prCPF8yKJV59lx+U9iZI4O6b0FKmuSWmrxT0ANsOeiexD7IOMcI83XvFJWLs
f2WEzKZ820QJX8Nbd6HwbSp0MRv/yN2EQDHlolXtfNM9KUFlnrijxnXMQIUtD8rW
mu6wgkQaUMm2KaMQFnDlnH/terYAfMzTN35KPLJN91QUUV6pR0EPhQEG86sWu9x0
PaBjpHKq+urjaVxvCm7JdpUVEYJoI3cFxYy0pl4tbnfRxCzuXNjqcProW92ed7JJ
DFJYKpWXpI01Fo4fvkJR3+O91CFUtOXLaD1z1emXwiFJb2h6PdhLZbABOGmaz5Dv
CT+6geOe1ITtM3BbyRGCPcghCfpMHS+CR739AuDl+/A1MUXsqbmbgJkhhQiJvaRB
mpzej2elQIM2tRDnBAqlKKCkxgJpjqTY6OeEjD+bb1nWvZWZ0/F1qY+xz0QH2wsR
R1aHokgFdj1jyykk6yBr0M5RSinP6fwIQRygXEuHOglZT6sESuLhguMgJ1rJA5Q7
ToLFUZ3YIjERNIV9L3ZrHpu/KKww1futJDLLSzfnSX8hQLXVfDXtTd/87OhPDpaN
Jvrllh7Jp3tE4/ahSfwsCnZjo2aOAQPaaw8DM7xdfd8zdG3JjeUbIVaJ+bN/MDkX
v+6N8Hv2fFzflHtRr6zTO+NEEkTbg2XbVgatUMSZmf/3eJWbxYVTodBcUvMKiRiw
zWwGEuuvR1GnHl0fubPpnRare4VHKVtejBjRGPkihzFXw8ji8/aloBwgIU83pv0E
ukZTkDrNpz59gSvdC/lQXu56dcNDtqGI41b4aL9rkLPIBzRST1A5oWoaI57QAORv
/ylcajEuYudvuk8uugh2eJGSb1ZDGx24S5al88OYxsXBzZyRcUndki++wj0+Nqsl
KS13VI7xxvzc5ud2QXLqAXmL/sGQM7VOiBGs9qa6b7bqIa/vRQL7SD4iS8LDC+5f
UkwHBFRFuwcBd7cEgQu1lq8Cerr++GEWHnnlmck3E9e9zdA+rBkMLILlZa4nwJg6
YOllWIcs9GdAvlMDDu+Q9ZXALeCGj6YVWdcqOS78u7YsGYa6uXxFJgr1Xw3PXyao
6MG6/PIEktVeCSYec7e3e7rguERUS6oHKON4QG2+uydVu8IYHAVxu0fKi7ngtNZq
7Rb9l5bzuXGZjtcIu8Y+8wmAfRhYmg8jMgbQT+9zprZpMzDXu2GbWpnUMj35+56i
xPxiqQFMieklyShuIcG+RYBwOQ0RWkkSFGLOSkYHpykLuqeCQepYYZ+AAKWxhFRQ
cnoo4bwDpwIWuP3GIiCl5mNMK5e4xosLPV+qOjN1Xp5Amg90AQpzfDAG8/azO1mW
zvuJdV9vQ8hK0r+aCz2DyAF0Nk4CNW8gDAtXH8t7up9yUUAYdzE71HxsudgNdpxK
B9fTSZUcslD97ds1xah6hEbVRSK3JbFFIwdW/dy9JnObSiOYKbNGEdJnUDcGNd23
v31PxtQoMBpsRcSI40nQ+QFpdXwKN3/YryIYo2JOkM8L649kpiX2XMXnZzltuUpf
f5MTOVDi0n6Jo7WFj3eJRk27ET1cOkfwdV05XkGcBC0paepJE+AkUH6yvdNno7uh
K9qlLUN7IS8tvWtK+y4qINPBH3+5iTedSQ1EzO/yR3Y40Iw2nOJVbLNk1CwYr7Tk
EC6+ZANfYQOTCSJ1vEFDjlQMsl60fIgOWX/QsfUMKE3Srfg/j7wW/MnNJO4n7FRI
ygu1iuE51RPBpefJ6/F6Fnivd2wY1tdQQtsvIiotuTQ/Hl4IhIzg1vha1n0HxFRJ
8EwPUJOI/2CXvgfYC9AoxfhqhYNfz+3fnp7Nq+PZTU4h5UgpyjnTpJGwHsYakNI3
teW1T7XwhEY+LAQWSDaYoSC0ymROhzT+j3mMQf1EUBu62/lpJa4aukDmAR1r7YEp
YiqG1d0ld8KYYQzpBe93JIgzhMXaFdtkQQzwaLiP8xPhAUaBfLLMwJaShPhbpHik
qTHGAXM/uPVp3k4GQZy36uenv7pkeycYAzzgSWtCN2JVMkUWHA9O0LZ95ghfI6SS
EB7ozoqadzzomGjvyFNId1jbtMf/DWqvaeBJh33x9uYZ8IKbzAjjj5BeSzBMX00q
PmsrvRNuYlIkB+wbCJkjFQHELIq/SLcQQEcWq3m7dBhrsBe2rBf4iCYZLXmmfumy
vfu1KW9fgiKE4DKvpTD5oXjnCktHuu4wlyoCWcQ+CxEWZ3GOBHPwj9WYZVXmsoBh
KF78SB/LXq1Api4r2WosSr19E7yWyMe5VCjgVtnAK1STFQkwgqha9cuV1PmvrOvZ
J3LDGr3yET6G5fw1WbJZPiBRJykaMBDqGwuBJtwlgtCQNBcs+z5ZW4oK4ufRil2t
jq8Jjd5WXrOwJ9e9RVY2xO1K4k5B+p/fxpMREIq1Uk5/hZ9O6/cDp4JKNRIeakLX
s9WTVIuCKisoSnwIhhk+3N+N2bkNT88xZ2BvnQN5US5hSvITrlSwANbF+gTQj+kd
kjW++88TYT4xLJgk4nDEp7zVy4j/66KHAK4J/G9V0NgJbwIohd7mJDSNOUZLEIGp
MCuJ9/If4fL4utiruBmLVjcxAxMNJ/Odfmf7WNYs/j3shbKv3xLA8rs6QZmyqN9H
M/btdOuYTbEpQ3v/KXJoWrLiLzb92VDzSw1N2G49grWw93Qe0uVkBx+fVPPi6Fa5
f3M7S7E0wMXDux8Czh9xH5j9PeIalvgU+r21kJM85bi9ZTSOVLSst2o1CjzZM6UG
ZPV+OLUixHMZiP4ALM56WpZpQTldUg8A+/z4ohLDcsRUhOrXToC5x9Nv36nAJjyy
I1mABbc4YlUANw91E7zoFPvUwF7BAYUo2omW0C0bjfQcgmiLzd9LFRJfBQYzpOvl
xpWT4sHztoSbAJISqQRXSetX04JbFtgyT7OI+I3s2LiVyFrtE8ZnxSo9D9OX4dww
49zwWfDkULkEIlCv/xzmjlRanRKZQz+ViGi7NFurewjnVt/33xkxdR9ROQXJSwt8
o+IvD3bYWrmI08k5SGJHVcjPPSHXNfNG++m62HBA4tSwzWIwdmqwQJ4kN0XLiagK
1aJThRT7pvJ1fSB0NsIs8pdhteoWgFXX5oqiDhoq2q/rcXnHEW9onTl7UJxkOYkG
mc6H6LxEU24nvLmjYncJHtYDal64/08m9Tl8eZthbsQrGbF1WBVGoVDTPsjc4yDd
XbbQGRD65tK5k+MefYb6wgfGY8e6PaZQaIUrrY75dhTWm5wxu8gBV7ZZi4JEi66p
IOw3ikx0xqYzpp9jDrTmH7bsD2hot/ZdgxXPvW57yA7Ex4jedjzaf77ZPty8S+0W
u7xRy692oKK7Bx4R3mSJgk0Px0DMYZGzfLLp8xQzX6f3+ru5rtGuLgGRHeUiSvzg
kRLCWe23Ey9nb1CTsRSaPqUD9ENY156rrNtxtNkgZCWptcYBMaGXMoSV/knI/LTm
CD1b0Hik6r8+ZrQ6QJ0272zQrVw9/6nLwjnGkPT0OlESXKkQRBzOTCZECLrqBCJO
uOpjGSjUw1KkpwswsiqmAaVhv4bgml5lm3mW/9RQgPiW0OsJLYDGIx2/rdAeBu0M
3e7yTEZju92mC7H51Yv8y839Jg3XJrtIFV9lJlaGcLPPlRhT3Dt1DtlYmp/Bgq9A
fJS2Mkg90xHyv2DQMYoZaMXEZvnDSHdIwujIyjtaF/4+m7Kh3QMR6CS9AL1DiuUE
3mL1pKXVUBmjy9QhrjsqjtkjeQnxKvrhueg77GN7qv/8V6gEnkZl25c+SWFghCp7
gTj9O3ftbjiWYtgMsZGwRsK7wyXczeCPmyLnHHYP2lMuRjQ7YuM82bWWy0DW8LSJ
G6OkJTTUGizgNQDSuiG7fNX8HILwqnrqNw7vSMHxIspf3wndts567/FlA8jPvKkN
zNIVOdLtIpdiHDaE5yRrcPT1FZSwiZCqZHMpWi9ILWN7KsL+6cy84z8K2nZbWBoo
y113iITubpMmQwcfzfhIaU6MZc7+oB0U5x3EtuM6wJ0uwYO4dNW1S7t7Apyqno0d
C3pm8fN6JgM5s1LrjCcJ+UMcdcdHRoJDypUGkV53a8FrOfkspb8uVXDInMi10qg9
6QEuwUUlavLwfEHzNYtJ8zRdYnFagCMuE0YwWaqg5hczGIuZqKppxiWFi2w+QJEZ
UCdX1wQfeDKdjnN5ClNya/Orbp+fcy8RiroDPDvzAkuj+Wfw3RaY9YTQzNxFz2uX
ca6og2lYwr5I0iHOFg2Y8A9pFntYTfwM/emcH3jR6FgIve5JiqhDh32vj0WeUQaB
NjkapgLQtvI15H1vV/67SvFAZ+6JlACg8NqyXaOAf4PvJgPqhKNey4rUWgJaMOBl
0PTuesBfAxlvubVA5niZH6gXfpmiyRF/+viruIXpeFiWTXibcDNYMexFA69fGP0r
LHcynRSte6Xqtq54lWvXiKbEPXkvdJNdPq36KJSGRJh1eW23njOE+icowEgbRRro
sfelQ6Nj0W32kMyfXdava5zeN7IwCaQ9a+9R8DNDU1gfqAF7KIbO9smMFu62Afyj
apxfIkqxM8vVL/wcuv82a0d+AKm9ksx8hOTyJD9C36r5MoHDR62Etv8h+fvGjV3P
eB12yVrVNDPp1Is/+ORJ9mJAxbsP5IzCYkW2fQHLj6OJMvAWHGl6yaLjM5UyfI7f
82szOkk2kok95MOgheI/L6fX3ISUncBRs3pSwwb/9lUoM8c55SCAAOSdYiO4+/Xb
pPY9XWlUsNe1TgT41HzMbo9YIp9+S2zCSSUa31XgJ/sT5Yx7NNJxf68Iv/ksLaYR
p5nP/riHMMLI3xIlxYUEprZxMaSAsCaRslYx1e7rLD2i9NyYczLIY1PWcOG/D3Xp
ecpvsWJ0mlSawnJLwMnK33+fv23qS7mw+9qSfTW/y3EdFdkEh+UMHgN1Ml0Z7Emj
guP/QZSoRFug+s1pQOiAovwIFCRYLW7RZThZ/fev0fxV0uwA+urxqo24YeNMMoPA
zpz5Cu5DTpuGnz4f1LxOXrm8Lf2BO+anWpuo6lZBkJX8NjPrHt4dHSuQq3sH4vYi
iBEPo62okVvq4EZ13AR6s5pZA5NYF4lDthICvO6cu5T3ajqkutF9uxJ14kpBVL68
3ClJInXrTk68/b9fSFZsH4XI+Sz3S28Zz63gcBhizFbziUCjVlkRorS2WzcmWZb/
0nNID6BW1kySvXUvAG4KxPrT8d1JdIi6P20t4kXDfevoDqagJs47dXrawJEgTZFK
ugBhPMedwuBBZN7aiUgpj1q3vrICD8FBGFHml4C54WHjrtHOTiVbDlAMcigk2J8M
psGGnUBRayhgF5wqZQBupYX5p1MniEVxfJspXqflr58c/1S2EyEOEEZv+IijRsSC
rgcjoBMg3ioTcdUwY62vYLtlhiPUvqV4Qv2IkhKn1Hepi+qGpYZCn7chldJMgZ5M
Uvsl+xkC4nuU1zYiVl5nw/Vvp4ccA8hQsSe7PwLyUlehXankHfb2v2Tf/J4pK0L2
czmHz27aOPqwBYtB0GBu4yTVR6yxPRypWQfli2OZrRkB4Ajlb/1saRn4Wbxmz9qv
ZKPpUmPzlUPCfYDRIY9xxiywNwrUdF9K00nxRIlz4eCW15PH/ZfGr0bosCwzjFpp
ayo8RPPoKL5WToiYMuG4mLlFq7cD4N3D/gZWFiQFxCpW4pawGhkAD395RYMC5lLl
BYNtNbSBUTaM3svHNsHAZJ1C6P3+kgRF64WVOmiJS7G6gWpkDlU8j+hU7XBfwHQq
7dru4D2B1l8bqAHp7SdsPcrqZF+dAm5zbuiVKydxAiLImHcPoW8GSi55bL6HpClO
bdTmyWe5o0vc4SIuGkuxwjuDgKsx6C9L3if7nNh4qMi1X1pOhr9Tadf1Czjh+ltQ
vJ970tRDXfL1kmdBco8PQZG0lIppskk1b3a8evv6hQiZ06fjo3+D/ZT1Gl0xYNRa
z3jE49f5fCj7m17hMnxn979GxY306tb75g4XC5yaZuIpMbwfeOplYdXCRvh2QESy
K2myO4oqbbj0FT5CzH4xXKt37ZaDq2ZRpiJBADciUrow6p7xjJ2pnVt+TF/hUqwD
hrpWIIaS9uuRuUNrCN9vt3gqPwW7RSY5K7oGmyXAwycYNlOmcA0EHeI+9wXlbilp
fnFT/hDEQoklqERcnvwGHNUL4Sc1BlIH/FE/JXZpPwpJ8lbOzxUfh2FqPPOIyudB
MVgbsqBSc8I2xTb+R3rVklWR6kGwX5nwef/GCCCKpYOhnovL1vpr2z1JwY9Rm94b
3CW6jqRRlIJl6k7DjCDCyOfZzh6eibvEH7Uxqb4FPRrRMSHMwZUAwid2SK+Np21+
L15mGdbAN9YElFn4LiIylg9gAA1ed7ChSxLQMdendHIiV/t2NYSyOyosJOnxARuB
4WeXKcZ8QptsehyZPICa3GrPnzbLVN+Wl43e6svcp3lkWqQNaSytj2KiFIuw88YP
HhPkh0i1DR+oxRIi/zr8j8qoyAtZkHdU8SY7kTRJKPyx6AGa7jeymDiObeekTMQh
CbemfR/WqGOj12tzXISk95HAhVs6GbAUMo4e768mdBzMKUZLGS7o2bOH8kG2P6ZE
/4+CkYMYpcot0el5IT4OIRzGk53x7ZZcghfm1mkWr1UQyzYcSeu1/b6IwqCNNimo
3L3meL4DED6heb7nQ69oJOxzvzJGSZXwurEJPLCF3Z9WLCqvLtBFup34iEQRhFRB
BPpa/fLwXDlmLq8xD2mrk9fFbW+0/nQCmSiCyoCYCoBEMJjZuoOIEjG844zDstvE
eE8NjXSsAbnOdrSXTB5kGRnaNe93q1+mrSZFpthoD+3Wcrijbi50ZiRbBVBpZJoB
/jll5nUorIWmhAAYeMow48SyBe7W32ms/ZOq5Jl5x6e9f/P/1ZWXQBlQ9NgkzGqf
srKcE4UFiGeX3qEsLooRlNOMugo5LAdiyYUUPE32uppdKKX3v83Gduhq3PJ20WNF
k5PW/LI7gFFQdoNxtwp+LEhGOTSr6d5ABa+vKq7V5K+9/8ul8V5WljQBB/XbfByI
GsUUJUgPMFMXBtSmERFI8PUOuQWiZtKuauwbCXTbCBz1XWU3qGcpYS7bkctcelZl
RBFLhPDNfptQeuiGJqpO+zmHDvUJIH2o8P9LPbXsbSBUQu4ZYZ9FIeQeJSnDk5nQ
AyT8WjY7gEsBVmFD/a58ot5DsA4hrqH8SwKU/sMl8w3FiQBFBmOhDuA7/inzgo2E
lb8sw7JmmdZ47IzmP4/CIAKDXJJEc6tWf+fltGNu0N5PTXi7KgXFsD9oF701/7SM
AgRXI/+OSfxyP/uUnkkDkF2/rquI85zO8KHoykAwK7T90BGFxZ1yw8ui1f/1ZJnM
bov15TWMXNDRyFYXKnbhltm7f13g6+CXKzchjRhGEuvJ1Q30pXSxzVcsmZjHpRiG
o/yfpUUZOu8gD/u9ZOnENqOurv9GE2+tzkw14bGeYdaFnjkZtQHcRkL529X3ibAF
+kAamSXrAThXVkZYEyXE7nuNAxWpipwYVNcMeRrrkLwuaYOvy3Vp2PaGFsZGioYA
iNyBhrmBtZXkyOrcdfoifMwRmoDVXePN0o6LUkCWlkfQVL49KOvDrI8u8H0YAiIe
jw3RQ3v9XbyhKt0r9lgXo93ktDOX+AujEk/vdH7JUelIB26gsVfQ+Heb6sK3unRR
tTlrT+vnOiWusubTWfV5EIf1AL5LEEjpB/koUW2zZuToBgaacKqk9gmdvf/eje5H
C67OPJupY/bDwacpJN8A/Z4DHesbm8vGXSbuERZTn88byBLSvSPCqt2uYkettVnG
cGbHwRQFCxtcP1HLHxc6hbmgUrPoXgxvJVJ5NBfecA5X3ArdNIlThqEnUCzr+M/T
QtRy98/sZoIXd7EWyWe70nJwu4L1AZXn4LhbD7Df9SK77W9X/9tQUJcZrQAIavLd
8OMZcPhS0ewhv68UOQ6HAiyNNaXJF1VoZKnOsit56SY2EWYFretH68i5roNTGoaS
eVCHt9abFXR1a0AxxjOoinlVsyFctHOONsGrt/XlwmXD59jpIrzMAvTwxZPbRh0p
rOHLTwbLmyc9SBBNEQFITlWRrJJeY3LPJH345MRIqIlGcII1sG48reMCiPjSkz6E
VRcLRuVaN7c/UN2wjUTHSmou5RriKlvNc/NRydJ7uib++JHSitD7wGAP2+yK4A0w
iBRvAt5F9DRp8QjdE3SKceSoQns81oCybOOFPGnqEGrgQl2fgp27ieX4WjLGCigh
e3nj98AUFvwL580JXKOvoAmLRAqXoVvatGYakYOTptZ38qBurHOu+O171JjNttRW
CMF0IBUbnRVP9Z+QSmQQTPiSihHRCFXY/cUTgKNDWJ4WpYynShQNww/BCXEFvM+0
ojU0VIaIFVmZLGM5XE+/PgadE1aPGzSemWJnD+dWgvhuidAfZ50026DpsgJnzfvx
juwYu9L2CNg6vFxxLUW82nCh77CXT2wD3reIfol9CSJBwromXj2jZ4O71C9y4YVw
8B7zsx5yoaMV6isynXI2qxTHCd1P+IKUQhhzHUMq2tjgAB4aaY5uisdl6v3SVeDY
53Yye6yiGFCm9js84/H9kDjs92gF/ipMw6s8qO82nWPt89W/50iFtcKLZECDZHBx
qT5PvZ9WbRukt38yf30z7ZV4SDlvGW+z7PmxCmlAOjYt9m/tY+wX2U/sC+w3nNHz
f1k61ZbEKO6pj6MyfgjSW9uFKm28yn6f10Dwe9OgwBXyVHau6kI0iZLzQdH9nxGH
Nvr1f5zmNN0TQNed0I8L0B/103BvHzzClLwQXete9SQR8IY7zWamNvZDzE+/jVoy
RlVi/ftmi/lDczUR+C5iV4rb6rIW6oFfHohtr77Eq0F131iBGfA5TFh1l7ambTYN
QNg1gPBSFS8ZVqPWew5lD4CYdvwRPpFqgZQLkprgKqhkpx4KwANp7+sELka6ffoo
ara5B6BSmNLZ/rxhyZO7+U9MHc3xOQeRqGtRfyWBQWvmn95/oBaPU1k2ZMm767z/
iQpj0m4bbLHk9j0PI9WLYo2csghwx774auzHcvvxa7yFlt63grqklSk2EzffU+ps
lGAFKYmVcy2c308KHjr8GAoMSFj29XCoIBNhW1sPPNghqsS2YFAYP5rIoMgBvhvZ
Ntgb36UPPYUVhp5U6miU/MW9rCV9E3Wsc7JVkYxPH2vGYpCJxwI4rQQDU26Xn8q+
AhVZXZH68ugj9HjSfEE8wK7pqFLu9qjtVPXPFLtjmRzdhTbOWuq1iiO8HKcyUQUY
vKhoJCVu2MyRzFjVq5xNyb06EtbkeCSLJB6PSJCqtn7zzZIVPlGn+lElqz1nwLOv
sFoNmLaFAUT6Nb3zsuvrDUOeAlOsUIHt4x/eFbDKsLZ5rG4eOAebWTxymW2ATj49
uO7YsKMxWR4iFjXc0GYvcW49qYXfUGAI5jOsh2lMAodEPY6mRXM5U+2jbxFhArKD
fj6oHu/RFp20f1PA41HyL7JWH8WZH6j4G+FoqSb2qeB61a+fxS+n5uIIPKzujhb1
knP4gRiRl1LXkMfiM2CmQB0Bjod3RBvbMRQpX4ko41opdV4edK9NmRAPffRfobkv
XdjH+bGuO2/AzgyeRGadWkcc773qUBnnT9VId+XP13pq6Ei1Qsrj48pwCIYcV2u9
2FntJ6abGabF42n9gFA14DIeNhA0L57zmvf5vs8ljtjHJXbc/9PdLc2YkM5OT7Sn
hG6Q3gkLw3DFy+eYQm/HFFd0522M+b1mrwux2GyIQFnQy9WK/9yE4uwMi9TBYnJi
K5enOS1wB9dBovUom5JMQfwrxrBGE5pmLSArYLDWiZVDP909rFjxnkoZcFodzY68
Uu+IP9eOPMOLZoBoQiyXatVxeyoLwkRFitO4h/w76auHALMxIcY6uyCaknzGAvqY
5jLopA5IXd8o9ZCRuHG4E0fIXAkDHq3y7WqkgZPp+MHU2+AJ4QJS/Wvj9RWPWAi3
VP5gYAudK4UF2UZy9YrHIUBNqA4dmYUKkRGW1Br/rTAdkvJf7tLcppq/5Yfv2iJx
leZH6LX2TGzCdoSZEtjuziuq6lnE0WCt+7cfZq+dZ78VQo3fLp6rB3tscm27sU8d
TKISaEpbnQDMTTM3WTYSzzAn5uf9HNqDvHJsZznI0tKX5jIXcDUWQFH3ktM1uliq
FDpqJhUtTxVqwGuZHypnJ6U42Gq9i3XGxM3oVPNz9V6ZoQqJPGW4WxpTKtu6d9G3
4K+EkNzbIa4zIr9Ur7cLkO0pjttWBYS6hADmNvnw8+8wngwjo8Te2F/OXn30127C
5LbieExahCsYBoQkgZ6qRdF/0i8PTkxk18XWY7eKZIlCMeiwpNw+Edbg/kw0yrfI
PsncWVQRw6NTFPBVIbkx8BIUB55yRTsFt/OPzXIHjb978ykyFLVc6SLqQbfUBu0Z
mgEav7sKPHHc6LwCG6JWa8fRqztoSdo+ff1qYh2QM1EkHzuOnkOUxWFSmM34nUX9
810e0y/4VkKvZxC//6nu1mAfbpWvF5OPXCbUuMeljEej98za9w4VKLLchYVdrxyL
tcaBf5F0KUcTsPQGtpoL4h1OBZ9lB71RAeX9zQCwUuXovRHdcbn3Xi61W0Jv+hqg
yBivwaOMOuhhMYAOJGdckK8D2++k5216Tk5/ikArH7EGKWRE6qKj+Bf9f/1RCwXA
VnssHzM5sl9N0MqZLxmUY4DCZUF6SEwe/0zUWNItTaRRxRaqERfrhilHl0cTdqx9
K/4VtG8O6dFqL/o/oKQqlulBagmMS43R8EHLEVfu8NNlQaX2mke4Jce81TPhTN50
wfutwXqdrDX9+RzDxqClnT/enB/w4N7z5CsrM1smKWa9mr0G2Qq5AKuT9GYuCOtI
0Hh99izgRoTlybMnEeL2rqbnhokv7XI/W9638TF1vr0dF4fZW6SEnl7U60GBkPGO
S+OihIcHrJiNgwGXys6rLQhfZ/F1SP4Vts/UwC3kFtRvjEFOIGQeIrNw0IF3XLYf
mq5frr6dLZ5a3AozRlAziNHk5UkmU7WrIqXfRTr8wDmSNB8Xnbd1VQ2llATnao8T
qgiyietYO0b/4NuVw8tZYGpKcyphki8YxPWnCB9+ZrgVc0fVwCAF997Vbo6cLKki
QnjzsP7v+PZ05Kjp4cJkypVzj7j+zTBBAPVz8xtAmXW1K40ncI1iiyvR1BvrmPyM
lE5OXQb9709sL7RV+GyUeYh4R80zT83wVAIzzXJ74RLJPrKUe3RprAgW8O/OhbEt
p1rfzAeLP8vvOOqX+G+DAQGiAhUGdXvMh9DO5fAkkZ9V2+Pn3SGb8LhRk/PZjUNc
uDY7js7lI0CW4sxKZrS+DQqDMnHZxSiYgoorwj0C7yxEukY5PPB/s1QLkIhhVDB2
mLAdJf1DmA/Yozhr0TuCOi6WyMWu/4NmQ6P6avfMpiWJSNZqii2tIJUi00ZdKoIp
C+N6iLvFzJG6PTvmXEisnoPYfYVYxM/ih5d0Gx+29s6mMAlqaARX3waki5nTJrzF
sArLu00Ija7/ksxxvkZ0RnBXlCnSf5262f0pHFAbtsfmYDV/v9R8XeO4zz1cESeb
480MKr9FV+FzitNcBLW0Nb+38eoK37aGlND4G/OQ3mDxS/gHa4LbBbp3MbBvUirT
Glrla5sdJwuzny2apf+XZcKPSkucgbV1+dcEg5rDS76buVUZJrTTatNSoFwL1P+/
g8AZdyyq0aCLsB0HYlhcyuOWqz1DviQxea80YmEynKyuVd2gSJewq2TUZgCd8cOC
EdiPqLqEuwdld4wR65CXV5heVYNrX4QcTs52Nkh0BfKYTx66Tn86PKCjAGneyNTn
1tG1mLdJqOTg60MvhKmobw1KnZXpdoBDdsZ9pWtiyFf/wqRcdfYnRED5KatZpOWi
HiKu4SmCc0r8c50a9FV1s9A/9PRdcuG4mye/e6kWYC5ZJ7loOBrwsL7FlhVcKHZP
BGtkLFCsXg9hUJktZL1B0MUc01fIC2x83TuxY5PTKSrBZFCTIhlhPNnBfAKPXCDd
20u/J8W2qpXQIe7xsCcpkP+1J1V1/N4JcakoiGUVFC1ngAdaG1lfZFa5pJPO5cWt
ymDLscY3KOLl76NAWaeZq1GH2k4QFQXJ49//vyfFLpoRrTR3UsRuR5J3nWDWU4L+
bSMpudDDUjzb9fbLHzvCAklHvZ/0xAyvLo3Np1E9yUmY3SSs9nXlMUwOkXoa4whL
MUeCHqb4QeKYgIsjVSH2Uq23tWM+Q0uZPGP1jtsp5FuGAMTqMQtg5Fy7Plzh/F68
N6Zx1XdNi9gXgE0LOx7XyUZ07O0k29WR5wcYNwHHjhfrm5c2P1eYt1fQZLChT16+
BcArPI1Fl+41E6Oh5oDcSfLoE3J/yoMY9SyREbsm+IPTNmQFggNAFkUYdSaqhy1j
KdBD7lXU+Rzc4KKMT+FAI464+jl2CUr368Zg7Ibgq+QUWmB8BfDs1KqcpDb4fN4i
h3jF+YTNa3/LVpjPlj/QJgTz128fCPUulvyEf830UTg9KDrea3evLzF3sKn67nwj
LX4VfDH1QBQ8CzeWnWOhZT6JFmwcuNEqhGYr6vhPz9uM/VGMlEDHlXpTwUSvKxD/
Z8LODtVGdylJa/9b4qIrA8KLCpyzneIZPts55jHvIU5djlvGduDS7TG2HgBvAdYL
FEI72WBbqmwyyJxW3Ff9PY+izMgdtFXOBCOe+LwHfMU1Hg09Kf65xaL7YNeRuqlX
KIJMVlESoQSzs3VyN8D5r5rb+UJghYSObxJsRjIOD6EQkADqcDhiL0K3b8WWjo+x
r+3JEe+8XFyltJdwaJoUVGIBJYsoaPuV0XIegtAbXYNRezQHFS4sUUYWU60RlqFu
XH+ckww7tYtBVzRYeae8guN7enDuQ6zWSgB++Lax7cPzC9ZAapyYtmNNbCOqXM/s
fpoHnnpXF+VZnqSr2cPvtVzAyaFk+oK67vQAsmtAd93suJoB2Njv0crK6xyFZfql
PtEbwXZ40CP5P/xQGFvtWhW3vogcV66jr4ljKdU81iA8hpABRkyYh7QT7bnlb7uD
+KLEA3lcIutENaLNg8HGcOAqqUPa0x/2SnmxAL9scjhIp7f1/jLVMuUiJ42TzkxN
Dd+WDrYWbkvN6KPIOrZC20HK1u2SO0qKH6i5Cn2yI7gH84CsWELp8jCBHmdY7g64
K6EvAuDk5mRQG6Lana73zHBQz3TEAD/zLh60gH5CxK/R7r3YY1oG5ltahQ7/3v6Q
BCy3mtIt+Zv0Ry36PMbSOeiGvAqDU5b5DgUxsOBJTgnQZoaRbDpOWltXl8Dw9KUh
0pC7fyTaFy0Az1Vi6bz4hFSRUxacmGr2gSMrZ1jEBUzJI8XQo8yg/vU/RiicDCaE
r7AMUWWaw5wqHMDk4DtmXOZhaOIqG+4yrrUtUbLQPN3CMHZsCuChfo3saJZBItlT
N3jzrU7BydaPPuOFkS4/RkNZY9/6vavNJlVXtEkXXRrkuj/L9Gqs/q90EY3Rtxat
bSg6azLreBu8rC1jDMB6h9ibbPIw8I+UMGkdjlWT/wtwLYvOAPrMPdSX98i3il2r
2T3vNe0qr+/N62nT/Bq7XNf9ivkbxZdAhW13rpleTsyrf8j2aV4GJTOXd2h7wX0I
Pk4BhT+jkKzf2xVF+ZvtjilfEiKVPAjxyIukbAzrq+4E79sFIP6uJlMifOFB6UOb
Y5+RgwhJNkKUs4OMk8/RCW02xkxp9wkJ8m225fHI1GBsplM3ZkhMpX/C2QLfw5Lo
pDG/45NM5N/Vs/gVOW5JWi+rHUQnTuVAQkAT6h+MgYFMnoiMfvNiQHOyKNHlBvff
7HMxJh42GqVtszTaLqAsi8Wej70j1NnpccbEEOoeRnJGvqpxlKCQ98+F6aBm+uiN
18oXZ6BR/h9pMYXe3qkJvp/I7mtVDZtdCSQQjxSIhM8faIQ2kFseBoYiYUtFTbk8
POkRHz1TzCSLhVphdCFKJqIXQPxum2UBSQS312O3itSpkrttO2laSGsKRNpOPHKZ
FkoNReGi+jGEbFmtmz1W1O3WU+s/hC8qQ9HIB4buw19X3hpZ5x1E6CrgngVXkKzU
X7EGN7yfPF4zBjtfOS6+CLgQhlfMAY4UAi2VPzIqEWsLU76EyfLTzpCcFhSZytx8
NFuspGcKhavT+asHt4zA+N8JM3c0HufUr/yjJlNrrKMbdA4URCYZywBCFC+Cmada
n4FTyxey79KGb0NYn0zeWX6DP4oiVcwnpBhayfKEPwyNZy7oJc0f5YnlAEx4Qt+h
rTc14OUVNOfNhr6wESU0DRH+yR/7OybZ4ccgja1bMJ7AkTi/A5OCoTDtVObT5g76
a17pDFldqfV39RBwEt2pQla4mdoC7cut3P26fBxXRekVAbzA63ZXzUV9SXddSEYy
2JEkyXzfrkniT1LE0r/lFyKVtDjlTdCUeD/9Nwh6kboA4n01dfZO9GJZrOx0GUaB
bV/3pCdQA1LVxDKmn5B/THvZCb0wgTfrDK30nkL+EcgfNwFv+bXXSOeoAytsRePN
B3KfFDY44Mt1i6AqTn9bRtiLO4odUIP1mYbR72H7wiGnq4B87XrwmheMpQU6uiUJ
33yVGY+6EWMjTepu+SaktnpIoa8u3/1pq94A9kzF1tW1f53RCymnRnGLKbbY27K9
QqCMsIwNKbLiBEb5zFtPDaydsAh2sdTle8T58JT8oMXvg3QTiAp1uypC4/Wsanu3
strMPJN8OzRdK4/ueneLWiHTqrCX4CCug0Pt5YuTzT07Zn/Tkt3866AdLtc/LpvO
EvpjasqB5YeIfCx/JxIcdOhsXh8J/twAMg1LcuLtayM5z+id/KPr0wIJRhbxK4vv
cYuNWffUVG4oIBaha4ZaNzlPqxuLRzfowq73v+uWS/AFlB3FsEaZG4FGOVc3FBjn
aNBYVidFtv3IcXjuhjzCQpUkr74gWvwZMgj9+0gfs76AAp0O4+4ts36GKvkI+fLz
rFqzUAqTkywhG5OAqK5avFzK+fdCzopVjUD7lUthVxm92KGm4aar9/099e2NaWg3
Lw6H45rg1UYsxe19DTonOjf8z8jr0M8CCfs/x6feZVTALdSKmaw4uEdctWHYhM0I
rnzRKyc2RGq2CCnBLsvLkIX8tbhJKh0em83na2OFVwTN1FfRcklrelni5k9exocl
CItHrlhojGw5Svpe8YIZPz/uk5APJ0cHxwCP4BPAgYN8CzSKVGlL5ezkE9kNGYtc
mOBQrwtWsNrbHvfQutGr9/0+NDgC9LGi7+0z1D7wghRoVkPd76vv2uadMFlXS21e
LApQx9Gx0O9bp77XT4rd3aYG+TonFkrXZWPzT1F4WuDryYAQUsczo14s7EQcUpoX
IpyJtpSgDFCCMXpJeb8jzZdbqyRk4ly6DZ0bT01H8xzyqM7PUOiFf/7D2Rsj1NAf
wFhHYSqpOgHeq6qlOl/bmBSoRKCB5tV94GNn44Xa+uT1Vwh7erAK0UgmmTuawdMx
c+p7xoduf3bKtKqSqg10N6eoGF7G6qu29hFNicM7cD0ojPEbDAL/V4hwFVilZ0U2
psyt2H9RXbiuWRhEKi5PewPSs++vSccALgGp9RH9Ss0H4Zga8avMGWmbn4nQBYji
cJDNFL8ZKrN/NFV91atJk/COyFW9zUuwr8IXSaXQLsNKO06/I12qVERMLIhoeFE9
B/htVeelXs2gvMiiQMCitCzT0h5y2w7YeU5R1dTv4oQev8illMdRmKE1s49OIAfM
4UcRkebWySzgJ2OWoqG1Gwg64AiYy/9p3dEEA5uaFX3elbStgEt6tQ2g31F7Z8Db
VwzfjVK6z7C+L73V/Na1O0mIejQWrYrN56ZbcsDi92UZul+UShv27Zj3ETsQgcDP
7zoyDk2iHi6a5r1QcC/RNsW134ghuKG0gXhv/rd1lJfsZ5z5yq/FMiy+gIpLluuF
QBzUadJno56pMnVYZsn/4wR06a3qvgE2Vp5h9UPHMP++KmW3ddYBs4Yij15kykE4
Ffe6729aPx5Z+3YjBOYde8QmdpbnNv7OQhoqzJ+7qsjNE8wlQPjpQd/1bQhE0QD6
SmYhdS/ASW9OjSI3Oh3WbhdcfOuRmSAdgU+jZz8z1xKrhDQ0MLFP7KbYhWB2N4z1
pGyIfUncZKMx2hcnC4M7tOSyeXqTutW7/JHArvCMvEyg+TcBz+0Ky/l70uHMxHaE
35Gq8mhBkmWaQdJpnem86UOstueVWJF8awRO8TgMgeXfgX9nxcFg3yXQ2lECUfcM
8Mpe1kP6DL/fpMaiwBL55xmQLyYhFMbgbccaaFdxSDMOTZwMzwUAQ8kJ/wZj4DNm
6AphyTgVrDetnBf8UK8Vzy7P42RBev0WMFd3Ry5ccqq2L6YxQmfEWXzmu5JP/8oo
MiSUhEiV8DHj98JuRLrJ2kBCUpItMS+4jvYRpF6yXRRAjhnalUW8yZ2jVTFg466n
fefN8T9WxzAJo1BlXINj11h2muoqBVw4tqHTaUvxqcQ42zzXGL5WapPL/hwghE+T
bD/VQdAf0eGO78lzep8H5KLj4l4Ens7DhMZJEXzhON4cIOTq1HiXzsF7gZ69M9Kj
KP6rLCnX2pqe8o+sZ6b03bROdt2nUURczMgTl13ztAeOsClWk0DhLgzYd8CUkbZM
pO9a04aet6BXaZPrHkTXvECOeUckB5Y6PRCzDe0cBK8tr8PkyH+gGWVHbYnn4hS9
iIkhhiM5vnr/fk2eRKGVh88LNf2873smp5EEkc0Dk7Ao0WKVwSNnG4139kz3hpiD
Amyg68wR7Xwro2BNgFREqljKG2COO0knB2TtjNY7vzk9uLozhYax1cqtx2s9wpAR
hG26veh6c/Z1lXu1zZ5CbZOTbEvuxRRl8KoAGLTUaPVoCrbEqViIWshB2WvEBPix
FnleS11Cjoix/crwlJRSJZHP5GJ6s5XGz3VUWSsu4Lc1NoqVfhKEFu5urBo1cpor
cOiCFguRGJONyO3XjdnpkJX922l40/ZkdVFwB2D4eYfEVrk5DVMDbWl8kreEITbn
OIVW76lOzpli8GBRv+6SJoMkiQX+/d5Zq7ImkhKplg6HQiDymjQK/pdiG3uSx7Zk
iFDkdvSm1oDeWa4EB8nWnUp8HJkaWdiyBqzhK63/uqGytUbnuYWmkbTszmP7ZZN9
3uLnHnYb4Nvyt4cPMqtePsfMHxRtiOq1WKHecIjvqTchoyJncT8J/uRO35wfGcn+
p3UBDOaGUoap+4bZcMsuId+3Z/ZayAm7mawmRIEY9t8szFm9u2k8TYL3+OBuefYp
fREb76I2XeITDicnj6hHSH09kwDUIWVt/ntl+XVhcELzZd7DE3L9he+8eZESk56o
nBm6QGQpBvIidzkCiyN9h0kDAIEBGXt3EFmAHqTAt5yXJskqvjeXPm9wnHeZOBZn
sb+AiPad+sCZTPJ479JXk4XkXjEG+wqp0+3cow/+9DeQKGCBtWj8LLrWg9VWOrUX
D/O8IIizOMdxKfCHxS1SlVezYgDKNO2ovpcGTFbMYJAaCo7JiwAi0NxE/JTnRlEA
mx1z1dXfjKVdIaiDE//XPgbjicGK4n4qvj1mp1x6HSBgPBYdA2smDtTPeJQrGDBs
6qSZcn2Znp73NIFEXp71hIFlD8WvzdcuRBnpjNapTKKHBIod/c6knyYdjBqFctQA
JkSg/OrbZehL7bTfKjxOMtX7wXVmCTuzWpDA92ZdgcPNweadpx7l8BrzufN56d3N
y3SwSycfgXOQEBFjCkPoAbUuxcKn8ND3YfyJErnzlUjMok8MAkNqS59k6X04RPvo
bk5DWGHHsU8mqR8e06T5j0NT8BhTaIvjFTZkCiJXg0BbUYO3ims1V0S/dPGrBJjf
BuoqU3NjzeCRcBP6jN+JUGNEKI8fLfBO63P2X9YAJhetJWS+LIeQ9JKkde4pWePj
pUUMUf6ewIMSJFU6oLhlAxu9lf+dmXPQIf/B1DbYTzaJkMrW/JA42bjUzfR329zE
z1/Y0whNZr06ZQCcyJHps1/0+WbjUY9555LJlsmcqu0K0/8Fpj0WgiILfa9Uh0n6
LrwtpyTjuv89dYlymRIXJz21W5PZUKKUoHNwVLzfMy4nz5rawdBPviD40JQt9n3I
COFly114pA/yrGl6n1qPkzmQoPLQf5jUOQLrCXpJJVkOiNLJzckzrujRBex/7Z6z
OM109CjY4lxIRq8rfxS/lgEWUIBEL+GywkPdSGkwyq9McD2VfyDOqzeRFzH5T2vz
G7g874Uozh6Aat5jV0hAk/5eF+n+DNkp/Zrgu2Yn71z4YDj1vZlL5RaKJQRWQH+f
83GO+efhiDbCWU4ep3ikzb6BeKQPB62OzqiWspRJxtQaI6J+aVTDHMZlBwh/MaHj
cHJc6GZyhi2ZXosHK9td+sMfXKOFeszz6bGi0Cg4mjJ0fD5Gxa84aIC4rfDXm2Mi
y6aaJjuhH2kUN/1Qk+/ilrUZR7f09dTj5Q52DR+OjEwfcafVzpvwcuHtKdfsCnKY
PUUNkhJ9waLnq5ogCsHR0ACxuv/h5LVTkM5fsoPpfwsC4j1HZWHuJypDQhTvx3Uv
XCzvMUaLU6eFhArw3SHM0T+Q0HdkXrjMJ4StgEjs9wAwmpOeQcYM8Rd96tclq1+h
oryPyOI6k1itiX7dsi2y1rG/ma9l2MoIXiLGvo7OKWj52CkPd3sr7pfggtdQyV9O
kl6PiFJk0KfUX75EK6nzu5BpP5bC6shBgiFDUYvgoQmRt321gw1OKOFF76Dhz0QF
5N/dqt+SACnmZEXGbZI+KqTsrLUJuPxhb/si6u+wzKc+MRTz9j/tOi0pS1wbk/Nx
tLoB6gt6XjNCFAgGs2HbDFupFrCDBCGmM19P2ktaq8cvxFh+Au5pOiQ35UqBlKIg
c+jlHuOfeijlN29wPuaW9gsoheOEPZaUVyr9B/nIhYhAkAu006op5nxGGkfNmX6i
DpRRs2/mx5B2xXWO6V1lYPllK8xy26vN7X61LzgJeYXNK/YlaMNj7MpXI44uPeEg
g0Udaj2kUhm/Qo5P/otcygYBFWds97O+UohVJD16xEMAxusvblANWGODRtz/UMeE
IDP/V0+bbNpTzbID3VK5eWr/W6gulD12+40YeFJEatuUacptLmAjH2amQSOuDW7K
DE/d7idF26AYaUWjKbBlbBZGinSyWwHBuaskpXtWjDFJ08Zzq74Qfmmy/D5/TUsE
DhHZON7mR7FtG29c0mKLABNvfjGIpKJ92hg2IRaCta7DdkIz91Sna/oyskXmqZTJ
FgEg5Cgb8cBVzVOkPh4ufk7JOUWF8nBuULs6qLUiUfcrqOeClMqsBheDSkMGtLPZ
8pCHKaLz4bW13l0sl6YG7uX4baAm76CiTga1nRUVfZKFs6FXl/PiTJm9qy02qT5Q
lyJHowpuYNXcP+R9h0BxYZZJFwZer5Gv50jcY4PM2H2Wt3PP0AsR3WtTNxdbV85M
wFr3qn5XIjqnvJsiH9Fi5UrygtPbf9Cbqndt9Vp/kARivfk6o8n1CDa133LH1Eqn
70xelFNybSf5YsKo744sOkZ4A58G1/LVghv3tiBCduZVOUUmGoc1X1ubWZ3Vr5nr
1C76Q6lMJwnAfm+c2e/KkGym1kBErykapgbNLGBoD7keEaWpVdXUg1FGd0sFCeRK
dDcgOcdSW6VgftpNSuZHuVj/sZYmNBFuE30PTNm5s4FofMUYTbhWsaWAwv7XvU6N
UNzvulDPBUDigVlkJJVcdRhQ0mnIKMqBYaexNdzu9sNGy4wUeW4x7QS+7F9o/ONH
AmjoPxM/TFZ3mGVLxInonZ/Y3OIXd4LwKOAtxiwZbDu0w2Bmm2mlcUlTR3g7bBqQ
36vL9KWlW02fWgRgeHoRsVI8wAeQxiG8uWdlXOzrvbgSIW0NiOKQayC2CvT8+SUJ
Y/tC8a1MGXOszWrOkKzdj4tfW8+0ZROsn/ykBuaB2f3FvQUu8RZy4RxByqPX8MWY
qwY/87yzYuja3kPEy465njqjvu2dy4GDqVcRmMLLrU+aUGlYCNFD+MsWgTXGESTK
p0rypoe31OA4z2DRrQxJ01eLnUOMnvyj5gNKQPXWkboa83rm1yxOrTkz47MSg8bd
q3LDYN163DO46S3ZXup/DhqI5tsMgnSVBi+/AI7gSgy5xL3BnQNYPBLaY1WAApRe
v4ZoAhooc2eQAeqrgepTdfl9ylok/ogh+ZyL1rCfKG8b/JIg96vf8cl6aUhF2GXA
zNO7A112iazFeM/jizTBEI+duO0d0XKhnFeR4rmMTO7rTa75UBwSowkEk3LUQkB+
SusA8+Vq7FXkoPDW/g1N9J7o5mixM/t7RMD7C5d0wClvC1r+ZiRNiK1+K6jv9PjD
EURIhYa8gD8FTgJjO2L/nVHy9PRm8A9T1KezaYldQVob2/ocpiju6NH8iZ2cBw2r
Agr34e8Fw5TEgtjRJz/ARlwOWPXEzQJzrPV8D6P6fuj+61MRRx6nRtpgmVE1M7db
71xitNPM9583AdsDermn7f8+klnfLzPHCUVr3XCZvEfX3QOW8+DrdMGXMS+pJ/SB
DCXktTYynaKkyGzdDqUoTyv3hT4Ac98hqSpAiYbxkvhdRR2vkZ5V8N7V0HrQxBMw
OUICLc8Scbda5CGB1xiv1Twa/f0FtnK/fM7/ZyeE9ZYkWdp6yuDdZBFsFZuNodGx
qBtPBvpD64cX0wyGd7nx/UFItInjPLOHwlhlRWWA1rSvwcQIzg/QNlILbXwtoaGX
X8BiRTU5UPRpYzZiQHrIQ7OtuuNhPDfxfuuykVB75Zh3NE+0CnmVdBdOGDtTtARL
pL5st6AxyNLVWw45QOiagsh2E7QhmNSVUNVeYjV7tgdk5fc+/xg/pRiY2kPe6UeU
XyMKPGiS7jXEsNnq5vsLrBvcKqcCNmJZ3BZoXitglxjrer5dTgM1gC79KhUlfb3s
iAwQ+446FQRohvVWxZynZ8AegbN/kdgLEtCFZAKKRSSlxbwt80u3Gw/8+GBM3ohy
zXo88FblM8+SvaQIgKoGSSD0lBwJzRAUxuYThiHwLvGvqZEkK1nZKxqOvuND3/+e
LAkbwjmglBosg1eOs/L7GZWZD1dBdz8+N8+dvpBsDN4CweP3W7AgGSgpPfUSnwBV
06Xc7aNuLLS29PUP/9/M7W4K7+zIqr6/oRz1P9aeEkoEuyJz+WewZaU0Egp2PV1u
byFYzDdWpZDo9yl+1+nV7IlBjyh8GB/NKiWcE08qmnph9ChIsoNh0Iggon//AJzp
/v9tBGjosVCw6RCijFBDVtaqhTd09grkCPJ2QLmdJmMHsoWIJfNZFgylWnrnrpj3
uUP/1pe7T4LU0rdhDKA37xpElaXDOvlEOu3eEmS7Otfp3yD7/GYjBydhQ+ZsI8nt
AKT2Q8eoFF0UQJGuG0kkMF6ra9j2OaIdPMr0I0Afn0GeBpJUVL8eVIkeEDTS2CCe
ar724Mfg+7EtzcjP1x+L68Gug6i0D9seYnquhOp/FUgsq9vF0ZFE2MWsO3eSyGDk
b9gOOllxw6xGWXkMvgotV1yGxzuPIsCnxb6xuK1AkplaXFIgHNxf4AKIWk20LVK4
IRRa3WV6l3NGUSSPUXDMBWxfDQO3uB8EtXHYoI7ocGbsrS9UfMMm2qWoBS3aSgeB
O0rXRa4Fg367NTdXC8Sy/6ROYkLMWZ+giMXXOOV19y9x3ix4dnIBYNnKTS7RULBV
R579pGHhMUlVAvXsO5o8383kL8+QXLv2hzveq6L1p+AyXNJD5rDZ5AgECp0ptcPX
AzwBBIKypg41kq1Rfuhg7vdpc+zS2DZVm0r2FRfV17tvLIJJ+/hBoeJhpgxM/pbX
0uQydHf/5ZBUgDUOMxXauC+23Xi08PWTG+FF7ky/gvRliY308zvjiY7Dq41pfVMf
Hd+kYmAoTamAGAz3DtOT+OviYSVVa2eIIlo+uC5PoL+mZ5M2Luvbi22rj3ut20ay
bDvFk7aDtdBHhCxzlbFzSTKvWLh0CgKDgt6eGITtC2v0ctiI2h0dyLJCwXUJMv8g
vjDBb7UeZBdCzpG3hWuuPyU6OfkVYaUtSUvjllHbTdDhkk2JkQamZD0OgH2XT6tE
5Xymbly1W88XXMd6LdazF3bOdQRqG6iAWGFrdKFc2PfmAcPHISKMa+Cob6d/CYeM
2mz9KQBD4FBv9ly99CEPnGqA/MTWdKzcURbCoguZtsd1QJh8J25shFHGYlqzjZwN
uY8sYUNnefZpPDd5v6stzInGw2qX1IB7HcExvH9zdAg9GzsKToJP8wSslpfOO3wZ
SVJFdK9YKbsTSrM6miGbjX1owXzKwqYszkN9SzrvG6HO96xxURpXpG/iafjSFiLx
g13TzJmI8/BYfwZ4YXlibMcS+qvJAdUbKzNyZibnRvWuAlEEVlyIE2x4EiCTan83
WNzhrLvGDcmYf+k2sY0C40VQfMzaC98YRESeJluUAbeLbcq3RZv0WmPH6A/gY84V
ZPr9bUbJIrTdaz+e6Ah3O8xbFRVKOxI3yxFNmEk8IcY5anUhDLOs3K4f/oHBp6Hn
GFO3q7v0aBWsEbmZs1ADRaneRup99iHrleuM9vpyd1hKXFFywBV/MPSgVgvpACLZ
F/kbQGiu3E0Gk2VLP1XQMjskPvzkr3Q4kJ6bB4v2wSNtop9fFMNHvvi6B0gbKiSi
nPukNDs3L0rxlPOJFsX8KQm10QNr3gJn4nqKrofjKyYnsWcrkqjYoR52jmIxvqK3
fsf6u76F3hrXwC5r3RMbUHFKBgC9rmTpKeazPa+0BosaoSKUnIchiMy7EaUBQ72N
mxip83C2kthRwLiCjE4/iOCksF2TNnZYKhOc7Q2iOzP/HRldgR+RHgid036J5IWg
QXRTCWD6BpAO2HdG5fks4YbMqObyMbDPTqfOafgLFh0R10/Y2OqzeU9mBY/SiSbo
1R0WbNshcTCUBHP/8DfahipjaLekXjp5NQSwZUk4K1D1I24ORxl3DgQUCgiETfUx
K3xMuDLYLAM2pQk+cjzdVbd1gG03KvRHRG/++bDKzI0bsnM/ocvQR5wqicVtCZFF
auTBkfxoosuT2j4qHMWkWgTfLWvafU6XadAzkrlbwJRgqPa9q98HsCpn6YQIRYu1
oWihLH5aQA28m8QNvz09jYiT9tTMuTcSHI062M0HVGBxWXiqoahgSuPeOEsVqL3f
fwa/NNNLi39TFcyQghURwQL5U7lHEe2KC/75z6nM1j+wIoPscqSQGxJBk70DgWgh
jTG/jwekC2DVmUTSm3vsNxdoXFB8oXkQdAVcP1ump4qeasWdh49OYT1gy5J3aybt
hvh+MnJg7V5aZc+pSPa9zaO/vY9Pw0LBShv1LsUe0czhPE83lRgFFZpLBMPG5eR+
OFSkIOFib/Ku0y433q5msamqkkzavd/SrY0lBsfxIYTNvrBgVx0qILoZke3mQ51z
68p3Bdic581N4RbYgaHaUc0HW1z/V617DJ3vTJkHIu9G8gNLYVct5P5KS/RpatpF
V5qoLB7ikBEH5ceUAgiF3YaDYj7Fn+GznNN2GOu+a2PKg/lVI2JXXsM0XMWrJAqT
eeCnUoyzNf0vq4yj6ekD7gNNCf4Cps5cxqdrVc6TQvwRh27yCmRlMTCOfvTq1ovl
Et13/Mlvz/+jlzgFZ4TmEfO+CeRpzo9IrnkJOKiLICrXCj7krGryyULZKcy+XJcr
LU3rRYAqLLdXnhR6k9LwXevC2vd+TP70UuE14PQ0u707czVxSDnr5T+9/Bslhhmy
1msdnOd/SfJCXL0r+zBc1taqHUbWyjqeTjOrRLL18RVxDDfYLCpcSv2Njw8c/5pE
3dTtIHog8ksZp8/UOE8uftbEoEpYec4lyK1KcDsnM26+9JFiGvAc4K1W7yuZK2iF
3WQzzHbaKsa4vjSdYvLCpekeGeV0PKaPKH7zVDAMHxvLtxS0B5Tx4qDV9abPgVpZ
doy1Y9XD2ttzmp8/M0nVOguezgPXcKzwW7UGnprYEtSxdGCDJdKA8j6Q12qQ44OW
r/3Bh3W1HrbOvtSOuhLdrulKJ6mTkP2AcIJJ4wXMA5VrcZSLjbzk1YyYOG9dFELq
pRq7H8SqiYC33BdU8KG6Ouym0NEJ1mdqVknn1S8Tq1t9Fynee5VRinLdON8ECAG5
u8SUoXCB2y0JTig0ZEB6yAVBkX+jXtTXZahbbGD2voH4J/Ug2Lw8qzQgIgOD45AB
QHlne09m8JkbJdqbgD3Ohq+11s0G9XmX3q9MzaSdSkhGp8BLyuUYOpDUIty2SOqv
CPBiRQBS4xam/hbIgu3I4D5Tf06xEuUuuWYpaw7EAeJ4+tEy6Lsp7LoOszi/nZ+Z
LTeRrwtWCgGqS5YBACdtGgQ09n5cNoQuEbcohMPk4XDoNUl+U94pFXX6bKFh+895
B4t0fYxX+7Bce49xgP8JPSpB5r5rL8nS5RqclLilyW0e4D6X7KygkRBpuSW69II6
d0zLWM/GYy4uKS2GFUV39Bz42nUBaPciy/wTuoKgE7pMKOCF6DhPrgk8+u8g275M
hObUbHWx1qmHlU94XNhfSgcMGb0peIOIqCDB3JatYYhha9dra4ph72fRm9pR2uH0
sUcD6LuIEHY+6m9vXzTdz4IEHiQRD+SFezXPf6iiVw1Oqooz0wY+k+cQsL5oVo02
i61JzQjbpY/K+gykElUi0Bc1bz3MSU7FgDbx6XZo8RJsKFufr8DWqmB5ZsGWlT3q
jTzWFPvKJMWFH8L7Up5ja2I1flDnYo1KmKANwJF0+Ak/iZ7DMWnQhqY5CRzpn2lP
28QTpIno9s9Km/82RO7nsp06sgf+3boy398uEKcJF43lCY8cYVP3dFl7/XcIP2Xe
UMOg+xMaRoz0pyhYlgZeffnuWhzjDuCPflWfLnIymA8lOFfXieiEMQCSmhFIp/Ia
+LZ/aO/1D6PtJXq/w6i9t+PTszyP8i+0+n/RXX6hf9nwgyr3i7K+mGOjmA2JxiCk
Q2OM1rnIq8jm15b4PPlmDdnh1C9yNal0NIEZ+aW4eqVuFT8Ogkt0qnJ2EDvSWAcN
vuh76Y8Pif0ROOINWMOk9+kIz6HAo5U9RprVvFPXUkKqFofGq5xXD1WjTVkmPCKG
w25RU/HqT//dYxTEwe+qU1eW5h5A5hB0aKxDbJx2A2PczE5De4/EyJNiPIhCt+Pc
KD4aHcypEt7elKGnQcp7GLjfypzqZ4wLp+tVUYnDtPVmUNgaYt2nrTreZP1Qfikk
fA8jULNaZygf5Ou7sO3Qr8dtZfSGKYy9wzRnTm5QjWjoGjmnxSrR9dxj3SH8q69Q
N7tBgp/YNfo3GAeNhLFmjzWrJwR7C3PfT8Kc0O5nPmhDE9AfTJePZcG/Ea/8uu2F
1qVIuy58xGtGu+5XP9TAcfTAFtmSc6GXN6IGzrmf3L/Jv04Xzear9r7oZxw/67/u
cBcUsMMKDlfFSkHG6oiyWLsSPn8Ykb+RiVpeaUzEHPpSPu/yz+QhEJs9KLuIll1h
fpukCBmdVU30UZ741VaHdM101vND7/6Jt+LklfWMWZk8khnLd6f1BFQWnY/7MB1L
OM4sdSyzrbdA55RGLqxtmvOZgueIRY9zPPz3Omu8e5xKBz9Mhip0LsuhmokWMfrl
sbxURTBT9MoBkEYyGywpJ7uqhU6RugwFHNX55d+rdgfzjtrJWsnw3Qdz9hB4JdOA
bswIh/+Z/+fRqSO9rNopbYN6/bn3xwumRp9r0aj47z7xd+t+2vsCBukzUf5NFA6K
LLXHDkgjiSOkx/HHyfxblkbMID9s1NehT2nNvasJQw1aSYp2tKkiwkm8Qt6aPx+z
zIg3tl3Bh3MdfimOKguvs/qi+het6MDbkimuue74heWVvNQ0k+PGIxpSI9W2RkLg
yOFeEpldhoyfu1fPmK63niR8T8hv/IarDzBZNzx/YgoP6BB5rXSAMK8Tem7ydPeC
Kix0pcyHIJRXsVvvTrIt0HGu1cILBEb/PfVzF2K3DjzF97I2r9Rb3Wj+FyTjrw/F
dwVkzPsGjM5nHgNmqC8kkbMrZEvk+YRfBUop+nz052Kgvy+kNrt4my9/dTTEA7st
j6dL7KhONwlr96ajAREAR8it445gRGEgqe61SqlCeOFkJPshUGi8K8Vp4/2kQyYo
12dMAhRIPlg7V4hYEmuUnqlSrTUAMzBnxGnO6EGtSrc0vAr3ZOnNIjZCpKSzQnt0
CnQei6h1SAK+pPkpaG2YQ4LptnmwFnKKz/n8yS3Is7iNBkVZOaRV8S3/4XcT0Jpl
oYLK/x1Rj0bZ3KVjLprHfvdww1YxisGZAxxu8dhBAacQubiX/rQk6HbKfZXTrk0z
RFGAihjF/hCXAj0AP/iQslFljF1PnNTe3sglyW/qxu6uh8vVwVU/j6kCsrGDDyXq
ifaGnkl/3lLrHMAtrg6KuHfbASeivSaH0zpsXCBdSrbKzIHXlsw5cBnsArEXW7QD
L8XJ+ZjpCV0c7cnzBINOqYyuwUriILEH492IRsJroMIr0uLDH/pRsB1+g9yiecmz
9cjh8WfrkPKP5ItGHekSSYX98FL350+nU3Xat4qPZ49ISt+9AxyLQgVTbLmQ5UkF
gSR3/+oj83eoliE2TTQRY0nVNtmtPUfBqZ5lWsxqmEUJ4lYuvuFvpjC7BTxF1ut5
PCqV1gmrExkCytKluMbCsVOfz2xy4pbbU9KzxohQetpq2E1yz2o6lljEpgEk+byn
JduJh3nsIAmrlsJz4K+hXeeRXGqzHte01SEpu2hxy78RN2ONSqZ9qlRXT62scARG
0QMXZ78/CrFV7Uoa68YiEjWULZPKRrNf/IbDrHeG/7RbfJi3c2hIn7XNZ3sJ7BfX
cWdSIe1W6vhd11VWEbj8zV8o1kIK8FWclG6sttlBng85/4RvM9XEdUKTw1v7vime
uYEmYO17QgoS7PzU53jVRxN+1tOHKEsRHz5RWNLZ5Nk0tNHC8zw5I4BMz3emi5vr
z7LAnMxsDC/94utM6uYNBhOA/gpePUFzjj6FN2F8rs02yP2+oGtVXANC7WYoiLnq
M9iAxdD7WoZVl7G6ip5BnIVkUX9/X9K8+xbFjdveTSdskIcpr8VqwWkZvDfvVc2A
nviQMV8CR3BzMfNG94cvpu0A8/5rJleHzXCujrf4bnVZTRHWM3mjIOABtbeYCXN2
elGc7b8JgO/0YxGX8684CHOKwFo6YZi3hS6gJHZGyjTcDn9cmuFuG0y9gUBFgRQE
jETeoMtD4UEHKLM4n4YK390fWH0CxPjIwjF15fh4BVzYdG1fwig84zGku2I3c2LB
2jeFWWixNjAv7diH5huH28p6M99cS8OCpIPDPkifTscylqVkfZSfMXSzXo9VtxXW
E1AJnOAc5VPXPzPhP6fiFeXRTpw6MGI/VyuK6ZYz+OokcteOFWptUH3OY0O/h3DC
LwmTjAsO6w69rjv2WmOcQESBu/Rn8m2H9beQTCm6P/YG5SB7za0P7Bl1rY/fT4XW
jCAx8nihAkKm9+7ma48vsQYKLma0B3TP3uLSfjdLZWTqTLJYDCKvzcK3HwMR5P6K
ZpATpcjeTckFvF9VwGKQ0lBOXyR/s6Zn6OOU9A0haLiLOBYvmdYJ0g2Gt+ftqi7i
sO1QWI4uhpwq/AkrWM/wUwHCSkQsSp/gre2I283egTSzNyDajd3Mpz3DsQrK/C2i
ecH9Ux1GYeGYf8vH8HxpGGejAwXau79+f3PQB4+1/BAo0/moYWPsotPljrghIUiU
IaHP0AMXM81S9zE2O/cei10193kkU5n6WXcCulz2f+HnHeVWWpah43NpkZXyHwAv
c2DL0Y5KiareOEu2OidKeQx+vD7+yJVFNqkRhqH6+zVA4TmHyS4uJFaOqEj7QG0k
arOIrHn8lF5OPMVIetEBFuQFp3Gx1MY38sbw5J1oe7lYaY8RqPFwW369w5vUEwkh
XRjiR5BfR+VljuSUbIF0eyG8ZozNl99JmKfwNH2QPlc3KSpf1/sGVzPDr5UOdstb
/IGVqB5pm/5HUXWKpI+Q/PxFvfkPjGVuGCmqLcqngcP6USM08Xl5qNJjkHeZ6x+1
aV3ViYMjWq7xKib+YWT0jROsE+T1Eu5nSin6fb6Uwk96wSjPjX4HeDLCHrepxlgU
v+6HbXL21q8kSo2JMy0/0EZX7d3V5DcLOQZ04JcKGlDaJq3wC+hja5ix6hElwm9m
soIjS0qJyG8qnPaADbFMowddLBdslRZ1ozzqgpGCz8rmgXpubz6w0BjjGzG+ppLW
REMS9/KorWydmRCmIARFht4p2T93idtyhlq3gWS6nuZBVPCU85w5g3OyuPLzsOri
lX6tU3LuhPYzrcQzEaFT08o3D32bc23bADENQUwLllFZHyWaHJL4sw7jLUzNrJPu
RYTHED/QDrEuHb6kL0ZBReNygMYQp59WV4REXK7rFwB4eDdzNKxmQj/erJoqC1qU
ojgeXWv6f6aeoRL1DMH57K38CWvU+amYVhKoqyI2OrIrv3rfrCwWz5XIldfr+Wwu
gO5O84DMBVgbMLsxS3/ylXdJDiPcQYub2UNJp2rWrKOYbZKmlftIqFLUUNAparHx
YKYVK9RYKm9c/SR3zPRKGXT/fZWK2GpxmjKVmw7kxEofphTiX51H0tmbkOEwsXZ6
xGm6SMyUGAGm21NrkW0a26sIAQ/cN9htatOn/CbkGoR8wOVw1cqZGaZ5ABkPzgW/
xZjYFRM2xNfdQAuT4AaaIPbQNo3v5Q32boF0q0lHq/PJDvARItqv4XnrkHm4Jq1z
Iebgadv0LtVbJKY0uOKrR9TLVilX0U0YBT8sVRNXbgzFhinQJcn+PhUQBqB9Tr5i
6pcEvTLBm6nXkIRrAqBJO5NQ4lq1ZgNo6IiPuOP20uaiWSogTiqrwgG9UNDdCnfn
Jmg7+VZ7frMMJZe2euav7wJrtId4H52AcLGS1WS9R5OinvnqUHkXiPFAqTsbUtj3
igLyWXOeol43b8ZjChcUmm5gQw5acygOms7eNw9D+GNPt3uh16QdbsCCfws/0TDR
MhP8R/RtnLiodbLH76RnWigNW71sYUOTYXZfcVb38CxLgdHrxaWsNW1qAqkHreG4
KwuBlxEyB7SCfG95cVCDryRuKAVZm0EqupUufUzsHZ6LBWlOJbP5q8C+ZBs5vApU
C2ricGfiPwM8PG55zM3L/cjAdaXT9/Ttj9GqXC7x7hp+mkdAhrmychx4fx+ubTpq
6IgAy+DCli4IWzLi0dcLxtEWQfcwAApy9ndLpL1In31Eu4NpcG5NjZKdDF57B1Jx
MQyfpjsPnkGbFXGw0OS7ipbkh5z7vX42Nqd6N5aoMOWxa6FSFFQNopTBHH9gMxlT
9Qxsj9CHgnlwZbtHEr4Ltll+RlW6/LSYwsicWcuG7isof6RqpTw0ElISSvLzBc//
BPbW/DySPsTI5c3NZzQY5aE+88QfdoXK2t7uoL0O+OckB8oSsBuOMmw/JUFiUSaL
jWtIwFMTH/7Mn9eeJ1bYbqTqonaJ1XCLE4IsdoFQEJQv4wNGHlSIROfhmkwDo42Y
1evmwvPjAiSYrwgLR8JRin1e8Voyz+fWWRBz8yA0aznEYlhIsC05s1Uu0PAfQkl6
48CJ/f92ji+Pec/DgvurTfWDWM+zFsZRRmgn7uLqqkjETebg9T9lDRQDbhj/v9UL
50HQPRdcIiyd5LW6olqfubz14Avqr8NMemBOB+OsJjZlVVqTzab2+ru3OZVeLo+9
AoIz/Rewg1tZZHSSosgmcH9OWbQYCyo7++bTZLMSj/tRM82HK+U0vbJnS4S/wy23
/fA9QpjgfJPExRdFEvKwT3CUMePrcmsLWTe9slsSbluXq+7FqDu+HQj8nwy/+sTM
iWONBcaalPaZPwbrjYmBBzHwvGlwONFpAwpTe3RiEk011uTbIGzzbOc2Juotw9wt
/4PiYfnUFqi63K5/9U5gmOT3k0GxqvlC83lp86TZiPxcDWgdBdK4PijdWPMKlCNX
8swskcCEAgqIDVhJ3btEFrkGFCX3Nj7qYZ2qzpOv+o8lsCs9EQaHbD4KrNt6ssJC
dzU/rQInNo7S5qmRiyiAv6f3KcoyUQb1bHBYtPCXAwmkuGRqFQJsntAxsIiyi2S6
dabeqVGJfufijD4xiYsnA70M4pNsWbQQquagm9uraEMMJT8ztbgqqwUu/uTJd9RC
xVjneoOx2dIUXERszIBPBW2pvxKre2XnUjU8IVZcDj/HYAs2AINjK9lnBb98GFVE
Ck5GhCOJOgPmLqxwPV+lHd/VyePc/Mi5yxmBoFmhxbKu7y5cpNj/i7+VD4SZqBU0
kgJ7fyFXHBidopJrHJKf+20fBRLnyYngtHRi3HqMa6pFYcWTqHyNHdGDZAZplJHo
TDXXSiIPxbOQtwOx88XVQj+HqdbAj4YQRGp60htpGJxGZOnDAE8W3+7xhFgV6dvC
B43oebJMobKE9fillsXT/BmpEVTPjcbJ13eJMIauFW8dg2xdokTp/st1yU2QTbOg
zj9BzoV3CiMj+7vtO9NvMLoIvU1PY2Op9DxRGskm44E3LV4T9AdfjJ+HyhiKfd9J
er1g5BBYZiOkJ0Eu68bxYH5ycY9hRtrOyi4LG4j2Tu1WJb1X5Tc3itpPpEr99an8
qdVuhQqZHARLVCaA2Ar/xFLoqO01bDmgiUTR1WWE6hh4Qdbf/dgRZsi/YhDPoZyo
SOq0sm+21Q24ZMNMe6cv3SqP5SrlyCpb52YVESoGr9z+xMsyyEKm0rQ4cTSAMIIi
koDol70Lg/zkZlPYPOjCLTqHson+rd7gZh3I/ev5FP9wI9kOHnhNZuy4Pfytbrpl
pF0uiJp/q9QUAAQNwuTaXAXNqxKkxWoQMUgzcEdIYy4vIn9iJrSRr1bNGE8+AZui
+o0jTj0Lw2une316X3SWRbKQJzy1atZiq8dZrPVgWGlijQrbNSAtvrmhobGeJL92
gdsj7Z9dDueheENCf900re8It3of2VRqgVIRb+2lnNNSo7xQUG3zUdbkdtv5kRYM
7TKIVVXJUuY3MSI+/uGARYPsPRYY7/DLgzossKiFeovQNM/s/5fEbZVNF96oDifO
M4yZtj7/ClUumHBvq5qcf1o3YBrWUwK9qFwhVLPkSPJ/ixtIjGAY17I6JWWgnXuT
ZfUYhEHYI7pK3wsW3K6ytUnGmHTyMMUmmWldgJrmTMsVwP7XVSnHGj7ydWEGtaw3
sdetQFDxtInmPuRB0rjgG5CPl76whqWvSRthmRmymZSDCDqIXw63eUKDeAwB4oQM
1H8ZeRzZnTzoMqAvRiYDOC2yli/tBbwxzuAAWZD5rKFsXw3nhj5nA9xA0Xw354cU
MSH+LV9sFmtF/dhAQNpk06h5a6diRnQrOwfCW1e6OQysqFNpYqDDunO9EsQCrWpN
8XcTGDDh4PTRrFWoU5oV03tM3YXd1/nIkFZ88/b5oeYb25IFkrZPtdGe/54qj6eD
BavTPE1qkfEN9IqeKssJsKm32VCAzVD060th6J/arm7mbjoZ/0rdb9gBWclTGXsc
KrbjCTNZui+Dsp0DAlJK+Rtut7iYgb4fYFl+EAEjF1iink7wxGCDC4O6vdLeO1e8
tjd8OC9UOxmQF8m6/FOC8B1D/OH/H6FSsqLOHRDjEWxXrkQJr/e6+SBU+thZJAPn
yRWyfX1GR9cL8WBqC7eD6fXY/52bobJ5Kw69DCqatji5YJYJ6mVvZh0oVCD7bQfR
rHCl7RjfbInVcUitHdd04CBF3EPT/FUO7eRWCmv5AMF/6HIrbHlQ9g6xiMGkCWQ7
MkhK7Hhr4ACdRkIZCIhw64ppAIHor/MMcHc5L4IdT7VtovXopEy7YmCx7B5NBdix
yjIpAdXISvS0jgg0OAwkW+ZXgS74kUB5eZxB+BUp0LmE2D/thXCFnWCVQkH7mOdv
Ffsfe8daqdcYSD//asfH3Bq0iYDKta3Zhm91IhQkttwgIDP6wq0I3UDX48mWKpB4
fOY3ReykjWaME7pk8NnBWuJSLpvcqJFQaVFTIMop4DxQLsXbarOvfzoS8NdmoVl9
90c5vD1c5TULpcTGi1Kd8Jr6u2FwVPG4U+xy6KpcJBW2uB9J9O6XlzY+2vcD0o+K
cMqYxqDyDb+AqCv+hTBj8d2KUffkfTTywwJjfbdRib0s9efbjiF0jyXTMKdiSg2y
5+ZUQawxARgoM6PIliDhesKd/ga474sesertaPEHiSBjoDsmX6eaLUZ/e2uB3+4S
QJujG+G/K0pX8Ii7F9Kf4yUGXhSsy7+myruJN/GA6s97TksWD9Uxmh4F3ZM0j7gC
FXmuJxtZwvd6c9Xv7r3uencsv6L2E5BparVYrKkQCA0LDN8mZoq57qJ9xt4yN1mx
i2RxhZUmrOjy52hGqe0kb+80WNi+nozh3lDEt9zxC36nguJX6EClfZgTnJ7VKFA+
v/jv9zG6QV8oQOFy4eXjoMF+I33zqNCIyQxtMO1i20oHAfxXyMNkga0pNwQqzh0z
GIsCleCqDNgjBuqyx8oe00lHJTJ5Tdn8lNUbIDE0rF0qmyiQPEOz+qtP9p2+8rtm
zONxuY6dkk4Nq1O+Mm3ee2GI8Sw4MfJ3UXkjkertYCrYh1FyAc1FNccKZcDV+iFG
wCtixin+NomX39YhIJm+2KOFWHqKuV9mTcm8brlwilPbffILnx9HqLUMJncCoG3D
Ka0Vbtmo4+Z/O35YYaAIJnRSlMT1OUT3DI2i+ZMxCvPiik7CV/wD1vHQKq1k0DOM
5z8GZWoSatUjs4H5b62WYMFk3uO2GEQcXImW7eww0hYCUhtq/qSDdEaYPRZ3Ohk9
az/qeOLBAN5hTp7aZ/WS4Wn0k6IFEsHCl7D7J8n+meswppBhDZ26g4E/7I6beGwl
7H1urt5TZKxUDMcVHAbZkCoOGUvdUXz9bDW2zjWbZ7o8J+ZEKHmWxITihbXnFkau
6xB86k9loPeHF1I6NrqoM5pgEjEfd3hVsVaGMSJxkncJbwhvT6J/vBuz9m5mnOqw
KDKmMGbcI+Etd6LycpLiR+nU1132lyjCLFDM7bDaNnNtsauW3MOad0CxrLBK6RYU
R4w4tZ9Wv5tjq9UQ+7G2yPPgSQiJA1CzFNYrXFCzcKbc1sGFq8QxsLhmBGB4VzuN
6en/zziD0boWtXhsiL/7B+9FEL0+DuaPUiuYBdD9QkTPMhRnWDev1DsYLsCe2vYA
9ePOzDybKtZv/rbCQMXY2pG3jYA2BumhoHSyBgjh89BybCz1uKJmL5CevffUL+7b
fTSx6/Ec/eBboWYqg4XbWIqB9M5RMgXieANZsc90nIXMgeja+fQZ+WxGYWV9WkDi
UaaMlCxaTaQKTurBzwSqcDkPubLSmAiAaEi2ozsqZVtonFhV3FLv+v45A+cz+D8I
rPXxCtoCjP737vTyQDxNSQxGTQvGpQUEglNssrzJkeamYPxmEK4SORaJJ/O4fFs8
uee/HvBaMCzw3DwFUo8PQI8h9vApDN74f4hAEi1OEqadBHs8Lqt6kwVIDfpo677v
eyhPVZqF7F+FM6V3kEFuR2t4jzeVnftkO2LtymouZxqrtz+uakdjRprI8qF29xeY
EJmR0Vjxg0VD3MWIpdhWD1p5yd3R0LNFFcTclcAihvg31NuuCQGTw79TDbHwgFhU
nGfQFskJ9imwvnDumAqgFtCjo/rg0WAai5mWOYJkCwPb+HYxCHQA17PDG36e1SNZ
i94RTeKDR0ojUkT5zUAUO0BRviyCD8+z9sf79E9r2Q1ywH0FE6jRX3uoLttIRys1
Djnm3AvwQv2ZWeR8wVp/n+mbnFjrngsa6Hdi9nqbH9FcgVLcX8j6+qLBPkFAHtum
lW/eVgFQbJkDJRCb11miW1xeapWzDduUm+CdImhk8FJ26vQEgcyuqVV61Q2zgLl8
X6b1NM14SKbzA214PLipdycJ7O7biCSft1h08ue2laYK4uKL1KEz1wa3zJC/y1Mb
ZRWzAcSvVAL3kxX0WCVgaVrilVpnkMSJKh4Lm0nToMK6//XfHuvdJXgUQkcR1Q93
aRQmT2n4lDB4kqOk0mvy8xfRWCDaczL70LE61GX+1LWA9kymjDauFYy5wDDE+uUo
a47pL4hN5Dq+gglvFPZz2AxQfZ8XtFQVh/PwLl+QyzriUJHtPufFESIcRC8cpyHb
GiU5TIQbZnOjy7JPO2EqvTism02NYiFKkpfVeLiaRVr8aM7rwyzUWmge/WmEb91i
v4EV4TO3Sd1lk3aVAUDuuTNCkPjY3lCP1U/+YTR/fXWzOylVHs/7D/MXBEEv9OrM
5LA1INgS88bfBVfK2iDh/Nd9I7QauzmiAAueJESo3elKoj84SE3+lfd7KPWA+XGZ
wZtg5HzUqhRWQW4DXXhXoDkVAkwLWfAbSWNXhTYfFeBIEB3pw+Ua2XfULu4c+atZ
5g/YsFQzRRKXb2ne1itFG77WdUSHRgHsA6wnUxfxtJT7IjzTApHYsVHbBUA4CREj
rr/UCZyXqozJ0tXu4iN8MokLz8rZfc4P4U3BSrFG2Fjs32x/8yteF8In3nV7B5/B
eZ9cCJYy30sDunS3yz0Y+TyY8irspNfB5kIEQ1THaQSLVawZJVGWF5Ie4S9RbQdy
53qyqQom1gsBnwHLtqIx6VnJXTF/vcPgIqnJ7nIkeYfOPcBCsp8X5Vc1cU3Pgu7x
TYZk2hkYvApkpVCWTJIERhCXUnIU5tuuXqkkGYw/eIH02Xi21ZB815ZBPGy47O+O
Es5ELT/tYhYOkbXueLdQkME+D/6M1kPxmIvUSVqwTSOecaPlwAMYUa9uVEDYbp5M
cMj1G8BJqSnetv91eNUXzK8oAgCcfFRccTzBgp8xoSmhm5od00qxzgMogCM9pIwX
yPkBQ0KaZKWA/E/FRaMATp453D1umTdviQV12DnEC5qVAMs6pz9Um8Cv29yAmYen
xV4LWq86Tn9ZSLZgx498z040Mg6i3BXY6475AK5aNEZwA08xETV6XJMJJbp2I/n4
MWK7Lg1JOFlQO/ex1YbzNO+au/7gTC9ChDeESUW8pXflqr/6+PrCLF+nEfDhSNlK
Wq5LLlGTudohZSDN74AMHz82uEOpFSauOiZZ5bGLZYHnY9ChTiiSe6+IEG02DpTV
sXaXUIR6NXOblbfXkl8+rvSZdXwB52FNVfqPaHWPAFzNIWPBV0oTmLVBeZpTyy65
CxtVFAv40U+nL4x6AMQjezfN4uBFWGm8X+EV3rfL728el8wUbLuMazkCDGunXcHh
Ji2qHkxNySxQAoiBchxBZ4gGDPq0kcxcVScb1YlwPBYhaVP8yXReQXCNVNIFjW1J
JFMTkZJorLd7fqpYVw5133LUPL16lDIK4+b6MZNeOfFA8LcQHYcf2rZBfEb7XS1Z
AwtLHjdzMnMrsRRZQoCcGVToYui2FYoyFnRBnUNtnqp9o2mtO+iIbyhayJDM06e+
X8FPY4NADQ582wTShh2QreYNwQCLpJi3DKsqs+3G4XOcYSlmcDfL7IO5to7v/IWT
gXyd+YJZu78LIYJ6MuaU6TI7okbq1P+7tp1/wuzVNg4lXlQcEOtFB9gqxSS1yOPe
lStaqxanCWoiJPiEqX9vGy29LxHP/Yi87LF6er8XjAmo3fqv+A7QaSndF5bD5tmj
y26E0u8oFGIZl1b0mEzk6jngkNmy5cNzBRi62tEogMh1aNFnW/vVT6bfKz0J+xI/
m7Jev+Zfvga1zRuQzK7LtSj5zCC2Ojb22cri9FoeD24Nc9YNL+VYRD2a9RT53rub
mpDnTBdNLsTygdr9J4cSEldfG6iPpHs9zBpIL/cTbLpRFs7cYNUK/9+z/CPF+8ip
MvECgrKeHwsRF/kGqdVPtfP0EPZ6QPyMunxOriVMUHBHkUzVmz2Dh1bkSXhRCmzQ
jhx4OGi9bsd92UoFH7Lx6dulrRHYLthKbyzZ2ky4WUOg/4XEKBhXUNZoZ+CmJmNg
fg+YUQEKtvLZ4PPOKIMDlCQLsJdo5F409JpzL130ykbZn/P+yH+WLOOqPMBTWBPT
bUYFAcst5CIqe/8ePNIZdNuRdY5qCRslDHkJFLZ04hW8HR0pBJWxe47bXsjICng2
jctFmrut/rWP7Sy2AOd/7Fcp0s/8UFj5/kkY/6uzJMSQRLyAO9E4bEgtm9xdUFib
rebEuWI6eyQ8PLOd3TTjv/dRGg80aN37KrORISbEemxkOqe+brFvrs6FTa6RdIIZ
Z2Mh/Ho8g3q4kRRFasvzsp404AuPQbMaoAC8qibhvnTEYuJsMMButuAri/bAeO7I
XNqQzpk4gp+O4O3z5WSsdiBum9/TANVE7/PdzxYpKWCU69gN1xcEbJG14nPgGggF
I90H+8Opqak5/vNMmv2JSvZTuHcn1xIWEI3RL802W1nXND6LXUHzoRSZE5r145NV
ejg98Ue2XZStN2uSovJVoTOWNqcaXcaeg8Z+Osx3r4bv+1kCdnsPZjo+6tCNWDek
2ReOFuvobePb8DnCt/0xt0BXlsd8yJd7bRGQCeoXUkz0vAp8J/hePcMDLMoRd/4k
ZI+MlrcFSSBa+HHH+QhLnf70kgX+5Bmb5HY1OUPqAIqyD1fnjFYHOebns8MIrfPF
pHQddCvx+1LF3NHrPyPk2mYnngjabgFIRTnDxbbl5JVkslySi4i3AXnO1A8jUC2z
phU8vmhLwvYhgUZ7OgNw4jUlPvhLaXUbDQmSfPK4nlhcpNlOZOY7IrvR9iJxcxJ/
FGQ1U+GrRNqJTrMe9OGnZ49Xr0hZtWGaUNPdlJERbl7/n+H9oGuPl4IHvViahmUY
yrjUxUXVHs6vEIIGAKV5MYQ4JAmuschE+I2t0ix/FOjT9XZt35cqcM7dmIqryDKX
WJQixTMP6AJ7KFDJYedXTLtfyhN2Fj1DuOxpkV9h6vVUALX6CZpTsjTbkPQysEMc
K0vkbQTD1C7d+fcTH9Xo4IieSpRrkF9w62ARH7FiQDhppM4C20aQE3fQsyd8iJN4
PM07h/ZUcOwZ5hU72BbEN2vk8fx1m8GqbVBYinJgngUxn1HTJJyof7SwUFLaP3vX
ChetGEK9q0A2QMvnctArZFJ0nubxYJy5KOVeqBka1iXkg/igp7c3EUQsH9iXYjAJ
ye/Qa2QxUemxoXsPw5JjFjSA7+HiXmPa32CBD2YPgzthfAHFRg/x8na23DJLtDPf
fNqVdK/UuqU/+SVWvFG+ZTC5xN7//+oUDOBjUovLBP0Kl0hB8pbrutCkKef12IjN
KFEIEGRuEQWHZcUgpYMCcHtBnK67vFhp2BfobdW5isSya2q+ZuxH2455YEX7Atuo
6gTzqCNrnfTvxB4y4E4Z33vIrvOaHIPTN+oMUOW2hNvBuxnNG0F0C8YgrYlmqsEU
6jAuB8l5SSW2G7vuW/gAny3DYep+vLI1brp4Xe/jvsfVsxWHxWhx7KYqhvrLLuSX
bjyeUNUgmySwlxmraT9Q+TuP7vXuw8Ig6E02QJE7R033/l+aSjb1qJVFQB0RR4DG
jQiNfBuc2uftulrj1jrdryLWSlQe6JNJMTSVKn/Hc8EaBtKmDnNOB3p2xBqgseGA
3aPrFcQvjjJflpNgZPmZFJKIdlxR+2vGIclyZ4/oM1kRbOb8eg51dxr3iTzvlCVh
93tyB4rRMQwo/9DzWum9m18y9px8u9Cn8TOPFgVxVHS0iQW7ogJU0EweLjbzEJ0c
6i/mgpGjKXn7kJKWeI9cTFbghHpMIyk2/Ms/0k3/tu//sMoZSKJo1B2xewrWpWXK
rYnsW/0YsbO1xUa+gK8E2ass38bu9Xjr1wOeK0UQdqvz98L1ndLAF65Dg5e6QO3M
7jsyI15if//3fda18iRJged3BCtkJORuk2pppZXktQpfo043Xm8njFjDXKhcG2oj
uP9vdrCDgK0aWZb0eW1XV3MuYb0OgnXnRzDf0ttQKt7X65H9il2giQQXXfJiipp4
vg+x47sOYAVRyf7cKiwjldeWxYUYU4WGRYxQwfb9vlihVFaFAORbZH+jwDfRUboB
gyl3b3PBlSZyQI1kEb8te2oZJCEfcq3/bGqGxH+j7N6BLbhND0rkzDc1mKeBlZKm
Ep3wTnFV6bLGrRFhk+cdfC64Ij6EJZMwheLGVz7FNbdZFJmsz7r+cJ4JnRADbLgE
c2Aj8j/ydwI0QBEw8aoNEbte46TrrzMGOfFSQ6HX/kk7NMhrGh64mrtVY8BF2haP
LYNo+gNJv/b0+YhWQbiN1AUUJ0l75/kdd0UR0FMLIU/lTVRlOaWhYV1rXrvb3clX
4u/Br2U2LA9Dy8HFdyPogWmIDURNITTUy2ptIjHTS5mWN5zaWEoKBShiQgRnwGM/
rDN2ZEKtqa82dgrJhkwpe/S4Ycxc78aq3oO01+oWAqbmkpTXuGRDaE2yVFEteKuk
Ojqtd5e9nOdqS3JlBDI7FR+tbk1SjF/YQTfBT8NwqwP7GC81XoGiij9ByjogHMJo
8QXimDkWZEsspa02jJ5PiFWdJR/3m9GF6XslsfTDMeDafHaetG/34VeUpKX3yORh
bHrZkxzU6R0Mehe6JgvqGrRFlEp19M41SM2j7uIWVobYcYx7eOY1FhJFGxcGWAh1
PidOx3KP6bZJ9x0W3wI7zLwhie/os4eNnGND4PSlYMymyjn4yHELpr4fV8DNAxI1
+NBJm8MGO0h8Q5qPlc9NzgsGjP9kbmpAKVDHei1kaqUKr1pdxLNmTWHh5fh6eWpH
/ZBnpLFnXDVu0FekCtUw33RgPoxG+FcWzzWg9HlMy8Nqy4UuswfjhJhjIt2Xsa0E
42+Kgc3QoFTnTgXJJ5ZM76qSR/nvKTnE4JkH1Oz9Ih2Cl7JPxJ4tu/czHIxAM1Q4
seeltfO7f+1mHdi5RpcJmv3tfIJ8+zX0PSkWrPVwIm2zbsX3puND5dW6s+ZnrYOv
35vn90dNO1qW16aasBNBmzXwvkfur9SQ/hRU2BK1/juNGiQgblub26D2FCvluQg8
WWomJ/hh+Q5BJ6RuQ4c1UeZ/F3kNb37eDqnwK8ENtkO0s+WeNkXYPvMS3oXl7SJy
lIU4IMwHUG3HzIOIPuTtyp6Xj4c3jdu/PpHmn1HxIpGFopzdmPkAwyZu8nWA37/n
98eYKzaU9Dp6dFibygJJlSG+At1Ln5YJdryO6yVahXUL3PCSS94fkF8miADwRyAd
nfTVJ1Xcau8+87m5GtifHkjk8MARPkY7zAAW6lKrSm6j81LPMcLXEEavdgUg7PSH
iyW7DWFsS219GyNo/yqnOfP3tim/WVF+5ulHYHnMMoed1m3VjO2Gx2YrHMa77Rup
KynLP0VLAwpBuLWIaBLEKO0B/oZWQhHfToknKBqjkSFnI5mTVKAMlGojPUZzMmyf
iCUGqPHpFGTpWhYekN6mHqNUSgvJZ0mior2tl7Qp+dJu1lgzWNUe4+VFy8oSagdu
xM7qYxanORLEHK0iBx9khP6TPl68iEFrYplimTtrUGPhTbfPp8LttqtZsC8v0neA
f86EXK8b4FoFl7eAql+bd57kK9Kh6vdSJQye4Y2QvAEfp39l/lsxZlLF0RPmTmOL
e8tp1ZECy/VPOXI7zZW6EENrc4FCity6SNZvDCz/jljdswmU1oa8G6lbDCBlKQ22
hCEyTyKRe6wiQApXRs337duevktOZbZL7xi6jQNraYM6CxoiJUg8pB4H3YIXx2GS
J5tDvjOlKlokd3MbQIWDNVEgZK5Btsn367lPKPMjCCeq9xrGCy5Osun0Y44P773k
reVlT6NplMuG8JH8QL3vH8r32aAFaebi2Zz8VeOnX3KT6SR56bbNiUD49tyezF7/
L5AuOEleW8M9Cq4s+eiu0wuX8bs+dHHF3PBP9uGpxiVgo/cqGiKROIvJNMdAgj5h
/PCog0H6kYISR9dd5aNc8vXJIkgjBdmAJS6YQm2egcUyaEs+JcAClykAzxeyhjRZ
jJmJOdC/bGAkjS4lbWklnTH7rgZIzVcLu7yi87FuFwGno9n0YfYg+om1Ty/2y/Ru
Pe+qbPKUOIVB61Llmk1Rt0J5yCLW7ghiwukLr6yP8ltjdGsLkex+kUu4mU6KkFWp
4aVe+JqUhEDuOovTq8iilnOqinjuLxlXVh99zKkNDu5dACD86gqvIHH9DnWqQvQA
zDi+3AKu11p3OL33lXqWlGGuIKuOWlY8baY09iC3PppLonl27hbMrlmlupLOCju5
vo4ogfkp64G4zczeKoR/rB1bWcRQNpngN6ECkOyH7Yb8ENgSuiDJ/4caAUQYOMPl
BR9vw6QJdde+2Kc6yy1fg+FQqI2voQlbGSTsPocrnMo9tWPj1rEZ01vvP18QkfNR
VzFZwaYDZnFUx35cIGwDUz55Y+CDLRNj1rmRP9tHAtdmucEaj5ykfzVddtsBsDSL
TLXl68M32IvAkDzUy4NraYe+McyEML+T7DgRF77s28ipy35g2ePeVi/ACCIPUAbz
cmoZrdVjE9GHCnxIXeWDAwYVLkIwiX8Je9R4xxc6CzIJlnEHxZdnWhhFuhgSTWf4
BVjzJlp7tTkoLCPbpweiUcenGKxmDSixBQi5zk8nPYViEzNRG382XDsGOWBaOgEW
ewEEjI2jbsKr4iHtnwipmiRc+XsP2T39O+wxRm1xL+0N0mPrsPNUzFku/psyouIm
mu10InarMmRcA25oNx7VAPPVrwM+iDVqC0Q9X5HGeV3yVBPbhALbFHfhIC/vQ+ra
PmXtAIlrfX8oQ+wJzNFKwzqjSQ27PDV7qpSWXh9MYFlu+QTrmPBIpLFjcU3IVlDY
3EDh35Bdcn9vA+dqmlp0q+QCUnDbZr/QyVHp0mX7UONtqsb3D3DOEDe2hZ3tf8xK
dG9dNzfIHVihvL3gQxGcvxgo1g7wn1nTLNtMYVQoybaSj/tqSsfUYQjM7sD7t/7N
5pwG9kJt2VGirbrQJIJ0MiY46326Kdf1lFltp03mO4qXHsN4OegRuMtcMQ/B7RvK
njzOtrEqHzrMvBIPDsFcCgTYTA+Up5jAZxa9R7J+ssSGMBlNh9SOg0z3fOjP0j4g
ecWqASVdXOAmS/MYMXyMgkiWzcqL7UFxm7s1wm1eseWSzEPBIF2AsUqGcmhi/uk4
pu+Or+KvpBaW6I+9pWA8vZ1uXaB8fNnlCCBkotfqN1uIhKaTVK5wdPejCDQX1tt1
R7DGTDHM+krWhZOKpfOdelOo78QNv5fczxOYSCr2D4219rotUnbhkwJCGeJroYwl
q95xesoGJTcllZK2TvheAHtoKCeiKA8XeObIvmegda+svuNYjJVtfbR5u20yroIx
z5ybWLQkxjk4PMYLJr+v9SyJHqqsA7ob75Ons85dA5WXTd9r9OFeM29fUwn3KMdO
KqqbkxTOyK+GhcvZZsMd5+smNJEC7n+cJypFyvArjaMwjyMCfpBeo35F5INXC4yk
VrreS3aQIN747GpTRLyfxnHlSABxq1UY+DGQzYfLHLaCQGPU+SlNfX7YPv0n11ws
RZGbdtPRQVARVkvHOlO5mFVjYX7Cfk1+u5cul56majzyxrtACV0sBmAc/J+iuvKH
p3/18ltPITHg5rGjBuKB59pf/g7ZXeMP6/KnVxBt9KnYQh56hYVw8vE2O/m5Ibet
mEZt19vMJCCzSoBYAfomXrv7KpIAkm1dCI+wEncF8Y55C+msNnc7aLe3NsdKFBW5
tmTfHuqfphWWnf64OnkZ0g6zjtk5YJS7VZPwraSd18YpVINFce9c1gpk1kpGxXfa
BPAmqoEfiiHHPtJt9912q+INki0wPct3A2bzGHoW3mcbWuZWQanCw187cHazCM7D
/Mr5ithRvU4bpefkxAuH6VTdflEEiT/oIgEFbFxTLif0q8GwGSRUKjuC5tcl4ERA
e1ea7aJy4B+CMPltOW5vqxlqMsJPXU8wPDZ4RuR2tcXPO+orUBPCAcpnJZlqFD5y
Dgw0jQFV+cEQkI3PZbNRJVL43FdJ4p+peVcN9p1R789arQ8uH08iGtNeSVn1m4zE
WLpEY24x5BemM7Xqg4378CJ+zFlNsugoxpTglCIg+dt3d3tPtI7pXGlBIiFYBldU
g2aGf9QOtsDE5zoPwCD6Y3jZu27ruOSXt8svagXwtUs3NdMYXqrou4XqusMgMBU+
a+GQMRj8IrNbuKPX+CDSf+xk4oiimpfOfRZYlnFtT42iXfx4FJuqaLzMRWQCTHR3
bxnMnpEZNRh8YBOeRWWKNFG87csaW4Pl2MlWxyQ00vrGQBxDyRrzb0IjCFt/WsLc
aFLjXch2JIyB7DP0fT6oPJm1BR8vyK5sCxPgWFn+iZH3IdFb+8scMbhlMApt9h7L
YLti/QUCbyrP/zzIQJ59Qmbk3As0PIl3cUBoMfM62goLAqGZksLRpMPxCmTn8Yrt
1lBD613vz4yvi5LoDAq9tBiVUA+XqZlHScYt/f/6Lkb4sr9i6UOKvu21p0Vh+v0V
rxtR8SlUc+Eh5/E0RAf6j8Q0AhB5v2LjmVEHmPxTMZMTm7XkoRFd6n9cnIDzmImj
6Gn1bdIpBlxzhUaSzZU8Yi+nGS8y5YOT3QGiwbchUib2XCDj93q6KfPUtErAxj5E
+3rFcjcQDs4GtPx/A5ijnXGtWfRFvl18dNyzGUq0ARqyRlMRXpNr5kaeyTTnOUrj
WY10aQSndrCRFk6d1LTMEQHE23E/bk2iMntxXk4IsljEJ3GmYFXymTRuMaFEnjYY
hnEJpBqK6L0bGfN7wMrIgXhpqvhMvmhkwfhd5gKNM3iOVT/kwUOHg0sqz23dr6SR
prCF5ZNTeUwluNk++hoPvy7j8b5quv23v/ymYi21bZ6oCBez6Pse/HER5J0zRiqk
l4sMi8RZYBOq4Am63D2isxcIkVYp02IHE1le+RKdIqKdBDvwK58C3rsGCgxXyY/+
t2HvitY0z2tVt7NOXSVrRrXYeLsBejmW2E82mqIjMbvFuG8QwWr93QV2lXFrAviW
9puWHHBUazxcXqL4mY2Suo39osBk9Nh4bUJ230AqZep5lxPOXJ/BvXq7LdibRnS0
5OQjjFlvVb7zyH0Cp+1aoaOgJ8XJAyAZx/xVOIxzPsfjIMKXwdB4ssfC/UK1va5K
NRqbdMx0jTE2tOBKZ9LmppT4fynVos86HJACbyZiDqjrBASk7MZAsmkdidXDMSml
xfgcmPNQ8i5M9vqlbUkhIUvan/hF5AWIrhDhWfWazsFdM43v1V/Y02wqslfEDUlI
dV7YNuY9sM/2sTQOl7f0FQg/vxlHG00XEhXRUKWdzYbDPzzWVbuJ5rEq1rXNRHpc
o0uOyoQV9WTF+9A78lYK9z7gsJG5IaAalid6CJDHsb9maZCoQBHwIqeWL+3fLF8x
wQKWBjtitEiASvmsj0/x749vkMbDnNtHwEfuiLJL2yUJi+5vqozlaRsmg37uzGLn
kS50CkABHXFmtvar7ocGcaNJfjAIpRglmrUBlqMe4P0O3egFXxvou9YjdAft/Uy5
TndBeq16LLH6QSU2jTOCtVhmrPmJ9DeCqzo2XsmKPNADtxgIFgB3n15EF01R3QeF
TGvX+ZGYPTuEdZiOpWjiJ56Y0kgZgofWPWYVJ3DA5pn8sCIQB9TM9m6eVQulGzWf
QGHQOvcdcjlIlbukhywWCkhMA/JihzAiS8pe6SKRrtsVMTRd50GJRspHcEQmMlfV
IJoXraSeguU+rT+MUNHuJMUtXPfe2u9QyrzuXaQkLFpT8mKKYysI6H545V+z9cVj
4V+iNHa8tSgw5aiIo/PhqcU1SehX4HKAhCBMhcdHh2yjTSxJePn0Q5EhYibdfYsq
KV4c4qf2K3J7DxCVLk/EGOqwyG7hjV52dHjy83fRiVIa0r3eYWIIP1lGOCsiwns9
TSCiZpcJ2w5RwSz1PPrEDYxKy+SwilLuzbC9ksLCJkZkoX+EWlU3xOiV9BhH+SGS
+cOPVF2Ok0GNoisr/jfsAaslETQGXdSHbJhsh+/3JBq9j4PjR1SYSgclYVF74xa/
9buLth1Aomhdb1OnoETz4bqNMDbaode9iFxsIwUyC4C8bIiNZHbqdw1Lr0lU32bZ
uDg05kf9fc9tFxDJq5FjzChHINJCm+NE60sVKiLTg2iiobJ53lgoHWFYn5EA4lUc
ZmyqrVJKu1vdr2uC8iFZvdck5XZRVsJu7sgB549nSAQAcFX3EyP1UNlbFu3xgZ+E
IVC8LUuLrgPccevC64RyRb+FWWClU4U9JA8X5DXHI1EMt0plseKg/lNDGlGf5geB
sQMOMCIcUzsYQYWr2Nz8NzzAx+YN70m3JXoOFqKXWf1ANMDbPHz7fSdjKczHPuGK
1nmO8adj84uciE0EgsHlbHet5kf62hgGDahGhqpT8xPa1D0iCUMk0dr1sUSZX2Ik
95/gQ1S34AgbSNgfR/ukon+BVemxGhMTb1ROQJY/E9efRHI1pRVRUAAXUnuVtYzT
Fn9SU8bVyg3z7WYC6w7ivIdtVdH2vp3d2ejMmmjtzI/iWwYxXj67+uJYDiQzH7vJ
NXwXQN8446iB1lvrzvylt0Wfn/IPqtQw4hHlbJveozLDEgqmv7yt/ft2b0FuTsNm
aOPG9gDty0iYFIe05GwToDE2us3BwyaM5k7HAXfiWLcOqfeevrByZ5y4t4x78mV2
4NfMSmmd5j4XBf/J+UHU5tp9p7Ga5VEclj5tARcjj9GAOJDjhTzQa5cCyBVxsWiw
B6XWhgwL5IAugCpfQ22gCdxDGH43kVj9ilVUqGhLkGPdPm5CJwN76aHxmwDF3Skl
OBvAdHceu5WJ8/VX+OBuobU+L9w0/HYX+kpDujeTleWDra0pFt/2yNlfxRHN5LW0
ypnfrhaYeVViRf00TRZ8n/KCe7vjQnAR/GGHMo73AfL3aPiP7WlkHdZG3hlbGf9e
T6T7SnJDuWINUj5qwRqMHeR3GlMwY0cDcyeP+6K7kVRPWHRJcxfHLgoK4jCqM56q
UBHilppfGS+z3tJ4VBhvblWlTlaTQeREfih0sTXMqNnmPqWVPFy10EN1/gmXq08/
bRjh8C1sDiy2IXImV920Ie8l1nmhoRkiEaKmvVhBn0A1/8BNNAdG3A4eAcEZqVA3
03E9iFahdSyYfHUoqh7HjpvHmmjLzlCsw+/9dA9QBrKEIx8hOWOXT4jkz+O6OQra
kofayh3jgnamTaT8YcOI+EwLMnJ1UBUMU4rxKy+yUfAv35vs6MKd6+j4Uhw5UexT
3K6Theq+k0hURLC4dtMmvyQY4AqBsamJ/wiiUkqjPjAO5bDBFy2n2pMluEejyzjr
0bsV4x6nkTogZrU8HIPXMtZ6dZn+Rrx+q87HlEfGDruTiB7++y8+4QgDSDtIxPGO
3Xxcj6Ae5GEY+7tYaNhukoYQN/OYntAj+xXTYeroEUuD1q1sllOC3LHzZZMyhKGl
n9CTFyDMI3gsd/UPTa8Suc1GXQ2kJdAeEC0dJT8ZVFQcldPgiP4moDhuwYjG+EyX
solNjQ5inPNSKVaXChan0QR0dTTykmGs0K5vsNZPuaPXxpGfRen7CkcMObUPb1li
TZGuVxxCtRya4kuRn+27KyWp24UEuQ8zC6llDdJlVmZOKcMZcgpS2d4rM4tZQGDi
VMvPLEb+lAC9gG6HR/DkuGNPfYSrmwnJzIGFKjcx33wLiVTwodJpw+CwAG0IoLhB
E7sS9Rzakr5fmTz5hIRsOQHSammqUUe+jeqAYdwqvnsZgw3EysblvENr9KULWRjI
bANzm/5FaPp3XFCszp7TA1KRoZc2EUW92nzKDAIkLnZ2zbhIh9EHFXRzTsLj7bBV
RPgO/GYhf+kXu+cPKbHp943ntHd3zJY4koK+dnJa12EZDZy5rDG4T3OdZ29bZYgj
jAfivwXi8ARcIcyZ8votrlOyDSoc2E9wqfU34DO6emFeVBhEh6n7qVSj4ZwKJGuH
bRSLhzlJImPM4Wmq7SdLRzqgDqkhUwcoeF14MjNB2HZXMC47I9MgQL6PSpQ15Kjr
h1bIhGAtBkhnkNUZ30G8YVHPX7j41x4NYZIn+PgDknTnyiCQIILHM5aa5HimDvGW
bTcuZwvQyg0eT8musKMuTGvztfSi71FgA6YBx4jvVA+XciqWtlWobGQNrGFM9S6Y
C1qf7fMUllpoNanIjeFFj6N4ch33X0b8nrAQywIUcanhlVCDPrMEqLcsflbl57Mb
fqz2/4QgEdRJ/IB/Es9k+ENv1uMldRr2TQ0jAkNdqTlG9wL3wG4kRHdHM5mmSYPF
NmliZ+X+8XaJLBFwVOrerjOJ/OtgjBuLH96t+hYMRO8E4FyeTfoOYBVYFv5Ld6bv
nN8PsxPAtQ+8E75sYnDYQ4tyr0tcokiyouVTQeFyldPxZxziJhTsnEtMUyY7Vitr
CbEVlWwd9EJoYo4wjSGTZR8gl6oPb14s4IWoWMNU4SxsUkJbmSKMjwMcLLDyZUSY
lO3c4zGCi5a0KimYzaRmbEPSce3W1IttvJpGiOboeDiqg3XFdslPUXGQp7ahWla1
IGXN6gTUxQGYSGSgyu+280aJ1pJuYJpvf5RlaLEnxYlivjaOGZLzO3XUL/kFX32E
l2zCoEcSCdu5/OJMXPaZgKV1Dii/j8qMiWBjRLMSDt4bHOaZRVJYddI+SURMnyGG
Rohg88PPPl8QP9kOVIl2JDx/sAoRbCfxwEjGakXmhfcNE1ADNW35RHhjbLf4oYHy
EcZ321cYxa7iLwz+eM0+gbL8r/V67j7+wLeDQU/uI38sRKL4kZn0NxM8jigtIQem
oB1XesseutazOTpSLDOS/FJoJz0j8dCeRv2EFJlyrwjXshBCKfUhO2becmJHn+tP
b4SDGLYn4KIO2t/UXDExh1yyj9fbJO5kPVWuRmdkKe8X31EYCXYrPSXgKTWvjWjf
Ce418lxG/N7kVRAoizKFizm7MXQ3X/9G45ipe4yE/VacaMXvbP6RuKFNLm0iwgw7
ytg/8+6UQXofZ3VC2ujiS40shSO0UI9EVB5qI9ee2hPQMiVz4rPwI1omHadxXNVS
Q0Wfj3pEQV2uIMIu2Nemq8ZYhi8qQ5TT7qhi73qJd7ZQGwYPSXs/PkGElWeL1Daf
tzF0w4Pn6djLc/glr8lKFzAf3pkgDI97SJraY1qPD4V7Yu1BX8ai+j9mKSm7tMpF
zhw3xjwcN7Nu86QQJ38Jyf6MJPrhzhynr8j4iJ+ZT/3MfrnMUoZ1rjC/btQI9w01
fNS0w3rd+slEmt+J7pRNfGTWIlNYfv8rIB8RBZb1axog9fX13Dh+BQ6QlQGYgXVs
OJwomevCYyj0XFz37RFyfXPEt6zaYigqLezyND46O3Gt+B6x3L65Lbu/Uk/alUXN
AUz44zld5SWmcpOae+dRGsC/dYE2q2GWCe+S1I6z/qvPzx+oT19mzEZTFS/miPG4
lJfOBY+3LffXefBcJtT6sFObuomE51zFj9cKfr5fbUEKJcKYtXY6RPcgf+MET45F
OLRfNii9mGWdZ7a0CbOPMDLWckLtOpgtZSuIH1d8UAnXBvfYxGnCmtWFnCMbSeNG
/yvTIAHTNhsuaRRKxQMKRmH69TBXir46O/abzny/mGoHktr+PZJVjAFqBqoy6OUB
bonLaNOVxvPB76UqHVj8dCjC2eb18gEPGJWR8xJb5jMV4OIj773VXViKbzcgfcBM
K2xXmsh2aeeHlI93S50RtPxKgn82mQpFMfMU1B5bzDSOJlrNY3oX5OIKAD+d6gG3
pmtNGzBcwrI14YFCsslPrP0TdJOBD49vJ0ot17GhdkdIhhyEh8qMpxvepgywM9i3
04wwFKcGaNCTxlPQkBrftFIaxjSSJ87jLOSgn385xC3objLBbOtw2wDfSkr+eQT6
SEpZ0sDYRaNPRLwWiz28wI+z+InD1tcgyaS6rSkjkiuslb2QBwrNdM1RqrKeSaH0
Fy0B7H0bNas/25hzUJvJ3lL82t6OEuAWFfXve/MEv6v5uRmaHKv4+wUIzTmj3Tyt
eI6gpP9No9wJhbED5iIfsA0+9MDNEnWJbxulptb7rQb8EApYiA/xvPZgX8lMECjh
kwBWuc3EbK2Hbd3Pj3yC7CDtIsFTbvVs5/S4BvnuryaF284IUxg+s/pRncQnD4qJ
PD5HwS9rwFBvwwAYD+r9M3lMC1CYdZMnVTzWkegJGGL/dr7VJnqMf5kG5shXudvR
nJorJauVk+qc6yfXjmfklIwqaAW6WbzxWKVzQtLuPsyPrtR7XBfNvigiJJvy00ds
d/Y7TUosMOU01EHS563c+dL76723XzlmqGx8Mq8ZhYPg+VRflkn1VWJuNhVO0fDD
abDASU8zzfqdnx7GSc2xF/9RFrfBIi2JBppBBJ1en/a/4W1hKre7FgUMr2vcxDg0
CYqUCpAWLXbCYcDULSH4qcZDLQigd7w4Gt4uIqptySUfk4P5i3GhNivtJg/EF+b0
oDpMR7P1eQ156KP64ThBG8TiLkMddix867J+cNxrwLUCVjKl3c3UV+KdOsTv82Sd
HdjAcSRN+vnLQQqzK5w28uRW/Z8KiiohrEVZgjg1yQa/LtGZhY80x6XCmwR6XnD/
qMpfsBPVyEaLoSoV72hlCovqDVIYHfzXxYLvY0g56IcEcZBQEY/i18rTXXCcABmt
nD/nfc2Enja6wYkddF4XJdh/81Ii0iw31lProiy0AbtElBiYiJFhjEGZ2Z9S/6TY
1mrTZLDr5KkEf0Uf07rHRgK0egP8+3sQ9yGW5G7r72NtMbzp0hoV62Faj1UEd9rQ
6jFHNN1Rn4I5XW0XHmRtCTPD9gpX3d7BdzMXFQXuG/VHKov6udsLcc5mFrN5dccD
aF/lzuFMu6mJaSHB397+1l4KCjozyogPYfcvWDB6leKQQBJwwauhB/8AxtDpgWOY
Ln4gu2Oe5zhCSN4/3Z2qA+P0k9ztomWpih26Q18g1M3QmnqGDn4BUFmJrnoYYjdA
7b4x1BE/0KFh7sqQy5J0dmjRapEg1YGEO/Oy6phVUL0LkKvD25E+bsp4UV/KvkMm
hSkBMQ3BvNZdfE7X+ac803rVWiSKE3ik/riGt07vyQr29UBjthZdgXcrrZEdTMoA
nCPS45VVOyWUJBAanrXyd/QBDyX1FMQfjFNVlZY935XOj/IBaZKRvAKkCoafluI9
HQWi4VBZCN4xapzSFK5SyMrg+kgXL1wuQZTRIIzDt4xz+OmnpnpKsMve90+CMuDw
lUE+lMJWKEWnM6xPQyug0hz/bkilbwemWWDWQJAwFDf/xHR8Twg/nCoM1HLTvexD
59JWXicpeDuX1erV5xYJJsAYD+WKo1wQ2lwzAcxFiXabo6MBPglP0T5ZE7rTTagf
pJ8jYBPfxtKyxUpAMSnnRVYXwD4jP01aR44nryb0qNbJ8/HVtvnqhUGzCFZzNwnK
fmoate8dI7Li4He1YkZITSDYDjCF6f2/UYltVXrcW2fC8/raE66Ytn5sA33m6WYu
sJlNKt5F1OrG9mPH7x6Dc8RjnUQZRwS/SBDc+4StfftHqPJqjB/pwUSOU80un/2G
Icm6Mdsa83U+UJbdrvbFUk3q4T/dlHzluX/BQO+7SLRTNqrnS8IWstZmSASoaK+7
bi5/calx9DMzF2b+5iTMZOmsTGxAO4Dw+LKHGidi488OSBsfemJ/Xt9URbWOqiXP
v/2E1Z1x5DVsJ2yMLHodLN7+0tw+8aL9lXx5WmEc8LTcar40uhQPe1iZ/iF/RISh
31A5zNil2ARSe64IEWx42t5S7xkUXX3rk8/WhYb6faV6VREKPWYNKy9V1XwOLLH4
R49JapP57f4K8GkkAigYlPvTICq9v3wiPE4UODV9g/LGM7ThdDGVgLwX425imEoG
fOtyGri/VxPP6aPJEQIMt55X3ee9mMs/Ouh7Ic8PtukfzS1J7Qm+/9otJi+ml+1O
CpwEQasMnuFzRtA9/elmGeHA7WPl2P5nkMveCv5OMHN51i56CrjSpWTuXVlc89aY
BLJfEcqhnHgf6qErsiyoyz1NfJlU9C60mMTkTNnaZOk7jcajrzTT7JFd1+f68/sy
aBstzNHYeJ4m0Bpzb6xjvTjYEmOhspFg0PQ0XLFYF9s0lEKoUvVrs9NeL1S0owqL
Q62PGDTLHgUDW1T6cKLtqzcHCno45m1nsbr4+3qhNicnicIREsH4W59yUmz3FuyH
Z1B83NW1P+LlfxW1rgYGjHX80RUWI+7M61OhCsgDm2/3FlUZ3Rc8qvDsH+93gxHh
FkzAh2VuZAFdRs4TEgz6bFV8oCeCDp67zE8dSZa4/OqcN61lavpKe48OEtIaS0me
0nIlGMgdKIUP0DyzO9mawT8Z9UvPfLIqN3dn+p9ijiU6NWjheF8xqHTtedHOnqQJ
tSgTCnIdP+hnPRj9eF3qagvRW7SSYWBnYfWhktylRKk8cqB1P83m1W/5Jr6Ru5s7
4BEYV/wgnPxbgrckgie95iqJl4x/xsiUFrNEbbDm3DT9F7CYoIceyrCF6F5z39Of
dLgEynNCRzbU/o5ZvVNbTbQQ92btDeRjWI/95rmqfWxEWKOhiWkdxhiZUpXFnfDi
VVQM3TxeCCxySl1MuXWaCVgQnFuzJPRueSFbRumcbVy34fYiqrJVKODIjx/7W1Im
7iKxE+3/Vd7kgQ7+6AarB5ZG1wxCjnuFK09XIDBVzbYASzvt5ZdjmjhGo9OGAw5a
FQFucJM2NGlTrsKkS0LHzwHsdpicCV8LwIajHHy1kA+fiIYiC+975ftAd7Fg8TiW
gX8kErWmUEbuMFKRe1zEM/cYgI+zR+sTplHnMUW9DijBwYKK/uwj0DQE4UNbMI3k
ho/VU57uOMUi80X64iLSKILgIQM3aS17nLtqJShtAQmkJR1oHoBoFHu6ubmS/sKI
re1fEOXALbVRGWOJYw+mxj8h5rOW2ny45J/b+DW7A0gPQSWD31FUwDQJ+KXbAfbK
OE6RbEXKuODrW23F03dG1ezLOVltfZYacD3HlBgs68bD5Z1F26eceIS0XFCWDXGv
J+F3v0t9j79+YSGYBEJxqQNwhEVyn+t7mQm0V0c6pTHSdtEzrPuQet8/07Gn/9BZ
iMc08mkjN6HXNbI3hTOtet5Hbx2Wjl6GQSYf8Z0L0rnyAVz1uEjlzPI3laVEbB/X
/X3kmumHGw3JMadjnYem5f4Pq70LhvFxsAaaO439M/6rMTSxuLHqKf0EN+UR+EzV
zmQcBQw08fCsyiBAba/OZxUFbX+FmMZcrpIR4BYtKcC/foBpuVCpODn65nYsO/Ca
7ob3JwRW2LpE7TTvBPzdvo4nZJeJU4+zhgzgTxIOIoOnBgqR9NE179a1zqAY1fGw
CxISNiFXUcwGzKss/cvjoKgZrtwaGI4VczwkpfcRynL52F+KMb9EsPic0/IIr0Tm
ONToX3j4AuVUOQf6OT7EdUs8zQav9Vm3NRTmSeLEhi4XbeWkN9hztuvfYNY3ZRhg
uTa9ufj0qnHVrUInPUVf0sgq+zcpacMG0eVzsofb9f0bylMZ+sBpP+EPVPw89fcX
/JW+duqDsC69NoL3PJlyL/HglHkTdEWC7XCndANxOkfAq1wptpAAutnqid8CFIer
foamuPoNMZLEMG/cnxYQTi0R4P+LKIH6527QHP4x1W/alU+bOCYnq+LNc/88bk7h
DSErUuFMazq0dyoSFv2nuzUmgfRJ249szAsw/VTme/P6nFzUbhgTpVqN7XjZpa2A
cyrczDOPmP8rhFtGgRn3Lsbilqa8tSWIYYg7yS2i7ardEm20wYWfAvWPIVBAGDT6
yZqpfBJg4GT7rp6UlfS9KvUUSvmu/dYwqydl53Er+E7clBZF30gsbnJRj6v2toLF
i/PpxJlr/e2au5mRd0GrnRXGWln4WLM+OuEIh+2wNnEYoY1k+bZ8AdycF9Ur8poy
NTB4yc2kPqwFZsh7jXnQ9VrscsdGUSV5kyTLqmFQ5e1Mmwr/4+1WxWW4PeimXJGr
hNhoxLnvgviMOt9A6bXmA+p9RQGysbyKptacEQxd8nX1E1McahcqnsHmSRrgtwFL
a3KzdsmuWD84jX1n+L4R+XEH+xXroC6A0/bXIGMiNSu8ELsVFJG8H+YJofA3O24g
ojf7TKfalg1NgJLtAMgRmWntt3cEhqf7xLRxBF229gW9phi6tJguKNQ0mHRL1NtG
bn5WSCFhwgJ5nnhYTf4n8QNm+KBllkLm+5hntm/F3ZVM6z4le8RyGSJNk5Y+6h1t
HgT5wpucYQlUXdpiQMa8KNFQe1/s1KVF4eYcL6Gvswivz3T7QPB8SH6H5JN1MR2a
seWRMgvqGQOIGA86Xhp2t8cm3aVE5BcxLTn1wemgHVb3jkyU1RlOZIFr0HAjDwyE
6BeZg5NbmSznsx9YQZDwLMdzDQQLx7bzF0tb68m3WnuutMgdNgi9HGEXeuCwl3SV
xuwtWTL07guIGob69Sf8XGEmdXVFLjDgFIiLrtOfAJze1UChQeWTw7/e5LOagn7+
Z+qu84astp6Plv1xYOtgGhbkIvCvdtUX0m8pfsbDK3BQ2wb3Sg2HiOFT8ck5Fk/n
ktr9lOrZ+D0DoS21ohGfj5uI1HArn2YdtXHjLOqP1PtrhlJjXWbrJM52ECwnYnJE
lzrZ3bJaV+d3q2zXYTl6HsAlww5KLL40OEpdmfiH8S4ZJlfxSPxs70RG+HwDoGOo
r8lq3qywEXeEZTm57YY0vwMHrK92W426c57L0kPAyP18Ed1XodazWnvYxp7z/QBW
J9UOTaA9MGQzFrvLv0118P59x1ZZ7tD3VGhTXjr88CKCPhZN6YHYA1QRVD/xK4UA
meE/iKtFYCxKZUbDFKUmgAK6nvF/mgdMin4O686oH015xR0D2uaWZCVsj8ru9d95
n6wfFSseTRvrKF9X/nDQkWBAq1L+tLLeeQIEBeX6V+XAXYgWuIBkTgfp8U8/cEjl
uevs/vvAzCSIPut5lYFr448TjXX2bdF9dYtwNGwiJ53DSzj6JU2QICur8airt1PO
N06jMNNWrxv5HaWd1vpC81aEU/Zi5BzAaQ0yvaBnHsHnOY0DdSJ/wQxzQzEb7TF3
wv1pQlIqq+BwsatsrKN2lrdWm0GQlE5Hk6eTw4UeScGi/pAYkb5icfDf808Ryi4U
5UoEsu5vbtcfznhOR3gXJmuor1NNo0zdXuKeMy/Nvcb+a2nVisIhvairICb92yN5
+ceYugEgolndfm1xcuhvoCHC4CAG2GFMaMN1rVuwFzjsMcf2qQ1WwxTZawbfjTwp
Na+NMKV/HACEbnpn5fQ4a/KiwQTOD4cQkjzR6cJsPztE/y4/zN8zqOJ52Ufm5mMn
EgUUSXXfY/TXXwtYUGkkUgx6LM2syr5vcYTUEpWVgXmOi4zTJpXafuK/rXJsRl2T
IzIK2P4pRgi07/czhw4lj5K/H6lH2X9Yyqqah2vUnpBOjqeW8sqOWwREgf+b7bmm
WcyCb3Dc6xp3d13pWK0VemIvS9Am92Ug8L4GX0SJQLmWitFXBEVVwweZ6x2X7j6H
lfv2KiAAzYQGpgrt0vuG5HmWnZwZ+2hEpkKAxIbQJRhTs9En4IzhoUl4uxAf8HWm
BpICyS4EUu4BnN7E3IHUzO9ub0N+nUu1Kcwkx0TzNrZkNjxmB7U0Qtor6HPNJEBN
gLZPmpY8SuorqxJt2g8XWc/6gNmu/uIIs6ATAlF0hRDE5+XZXo8v43/pvOmMOYOb
t3cZN9xucJw+n5Z3NXeXazZRFmjJ6vd79UwV/83n9YnW53Gbruej5XvcjQk2Qx1F
FWUl2YBKHO6voKwE1FdFpocovGNvO6MyURixp5439k8vW25OTujBFRTbXC1SciTG
xyv+p7fDk/OUUv7lu7N5vg/rg4E9kKhBaQ7/m/Z4X8yrffizPq3bzZc87D/Zlc/L
choj7evIUTKgHlsfcv7kj1cGlDWtTxPOqCCJrZ/YGr/49fUREuz8/lQKcvU182s5
qiDZdQpG10wwIvous51dUt5lKgrRspdKK4UReL+45sEp/16/+VscUDFOITLoRUyx
2mu2KmTTKAGo4vM7h+rxJIvQYWm3RGEIoz8PlMs8jcdImJ7QAS7+/WwkMcL0DlDI
RTmA++UlWvZ2QfFXqAvj1VQlFZnfVMrNnNlGPNqU32ebc4j/Z02aOYKaEswNUuAV
YxzPYbCrstnFj39jV5IeuLt6n1QgU0nbE5uBZizqD2N1rFPrz+0bnunYzms5zbvr
Du18iSlfstn8C2HRvKa0HOvOdIHquF0HdBHsId0jfDDGRE/15MsEy2yug7gRgshY
djEQ+LzyCE7gn4I24Bw0SgWUfD9bzAZ5Fqd3uv4uG5nWUzqi8C/V5kG7i10RMc5G
zUn1Tc49zs1RXBVCmsE/0ZLylyfO8sTGXqXnHBWfrGPi6aipLAGZJcS9LW6ZLe/s
QPNtnRC85v//C/JI+rwoo77TGrTNXecrbjSYRvoP57wIseyvCtRuO17lhbQVWxFb
buXIF/ApYiV467hUfxeZPiY0IcJAkLE6UgS4AMsL5NIRH01GSORZbOFZ0JkTlxSa
fqDRxRD+ppFlX6xJ1N81fbFmm4C7ucrUHQFphLZLYy33ViD8aLgr4qV1zAdIXyKP
3kgCorqQYYUtolITVEVKKQu8/EaCn6OsFylUXyNtRaTsJCU17oUfgOkxpBgkNedw
8zUfUlGEzt3qVeODWiXnQzsFxd70Kh1NKEuIWHYeeQIDXOvAD4SxolzruPAT2dvs
LIZhS8+8bQvibhy+NQpn2B+sZpqugdjbagrILpYjAHtiYC8Ve3rm55MdiP/gp9gf
EP46hCNnWGfzCE8dy8nWmE4Krm+OkNwmg3lwLQS4HJUCXq3xbhQSXBs3coi6YMTc
PwNpxH48P6t+TFXe/p/u7p/pDUCF2A7lMNfHCU2VqWpByiw7yFTCNAjmEVH7L0zM
XuAtAQwBCsmvzHXzDaSaT8PHHQvkPnDH1CAJe0ZeXBUXbNl0XJ0IaGbOYw69GB7n
diWMEDeZtKKIS+xA1ezML1Wjr8SSPQ1kgi2qZrqDSSiiMEAQxJC4Q88Y4TTFmMVX
4BpaL2jeEGI/pqiJBZSZL1kxxtIJA5CstRptt18XgQGXx4skWDsgT2vzuYs/okPB
lCVM+tbx1vlyk1VZhdVNRGOlcU3/Mp5iUMLKHtAvYg/kqJ0dnd1689kCoNiTcr6b
m+MiA5ayAS6benL+dDFqYegbV5hK1ef8SWQeYVRaCZ2H9q1ssFF/Aaqead0ceHe6
EnffO4ZNMUV0wN8VRO9qXBVZpvdZ8wMB8e0ddC8TTKySZitzi5BWEl61/Thot9VP
dZdf6uAusp7poUIuikL7LfVEpmVozSCgRrfU/nxEizucyFDg/MZgmJqcs5Z/42Ax
KM1m0d1rgCLNmA3kXZuL9tER5zJ3xmWo/9+AVFoBdHZQBmel3j1g0ItXYs3oSde2
n+Q71iLEZ8DsO6W/x5X9Udn70X4Hc6TvwQOxVZYP8zuNxau9VQC3gOLTex+/gVDO
qzt1I+gQ8ZyQk3Gs4PAPowKZdu/J0RNoECEGzhbUD1XDDE954djRL/nRdy0nUpre
AfqmCPCg+RznoQEQcViSsfXXnJRKENuv7DouNm/CBSqxCPLh8hZPI8LqK/LTDazV
x2vM//Vig4rHTPxUuRFBhq0q39pjQ72yfPkHDLHdbsP5YIcUrfbxEVSMyxFPnrYB
DwlEyaMyHk/X8sVV8uTN2ilMAB43XjQiWIexSBYgVnppVI2nbuTuQhUlB9o4Xhyd
CcxcVFkjYefbCMM8OdDT1SPMi226zSn0HdRnmYLkcaIePaLuleCL3iCA9MydAGS0
RmT92IWSy6CFTNqPOFRV4+Jx0Qfj/UJWHPmL5M4y+OS2kfMF0QhayO1so/4pUWWT
cdEy1RRQc8uSonIPQEBsyULIk3rW9GJNFgvqWK2ONloAs+nP6NitDK1KnCEl8E1m
vKwMHJXE+s0iAfaJ6QX4Sr53mAaEn1Bts0FmejGBzIx6TP7DTlIIZMQU9a8n1o5J
l3ZkM/tzTIjGxN0pLJdfyEQYroCvPZGWwRcu/IddYkHtdNpic5xCQw6rOdNP15Qn
Y7YwzzXk06HmOZLzqX0BtbZfB4BNsCVU/0KWm9LSGELUehR0WLSr9OzZnLJqj3/e
i82IXgxC8eEvIUmQHBX/76JL2wRkBpmW2FYmHRzcPY87eYZCDj4caGZ39dQuHlJx
AwR6DUEBxNWax+fcsk4Mpd44Sms4u7FNVe9KTBIrLcGSU8GmpkmloesPRHUFK6kG
GMG0q6vV2+xqHtZ3FQpuYxkOujbpD6f7aHlNu9CAVyV1EeduZjvFGVi8Y54yJ4HU
m2D9RFr6rUyL4OqWmlYujo0xoQUTi1z5utoEUQaLXaz0T3ABI9Z4Lk+425nffblA
rusOjGRasMeefBXk3aZI7VOw1wEer3lkdpejoL7sJpfQInu3jnXqwV1MeSD5/Jws
lcDvaHuwqV5FTQNYMEOeNPK6TIUM2xLYMgAOg0AtU9w7QEcuLMCzfYvI8Ca/pXBe
F0WbQACLJcGpXjzz3UUxPylbNCiWKMU/r45MLXxkPNWQfMS4iCIQ2bT3DWySnICC
bW8n3P3SUuGEsrtoTLLFoL23vWmub22sWrraLQl+1RghanuGrIcK92tfYc3ZyF+K
qfs7sZpOIgHD9ECPkquHAIhXgE2bttYaB/L/crJ/DtE6zzgpP/uf55syrNhB5IH+
45DmhlUDbxIL977XcqWxumIn927vsuH4ub4RwCm0NEihuKBPY/qH4m5cqMgaW6OK
a54wWXfcP5QDyt5tc8oeiKxjQcXnzm4cur9azpeCFJ9mDLRiyArBKkGAt5W6d9Bd
pgweE6YgBxBMqK8MNR38HityraAb8r9q+4rHbPpm7SLxpwkEZVAilEH0XJ2RSkki
qE9Hz4SONdVPJUhnuDaC4M1OOmwU98SsaBRzbuNnhQM797fcSObdWj2su8ZoNzp2
Dk8cF2zqAF89hsXVRO6UYNkkimkEYE/hkMIQF+IGY3XifEUrfEZx8eL+9clRMSpa
2Bgqqlv70c+GPCESFod6+o2aYqtkOb7e/gEsuITpJYZf2n7MrqhveNV/4pKwcV+A
ekqpAuog0L3fVYc3iTykKK5NN2xDpCa2sivKnyxE7Zv+NlDZlTC4RM+4mj/BUGYK
cmVuGIZ5vjMIO9ESTfIZVXGP0N81PZgclyvACwUa1dWxSqezVF4e6yDaxp9e9ZyS
7xkAhMOcFIXyuUV+JXODnwQN089BSQJseQoZqGiOIwEkhYzO21+EOE5pmllJaVjF
0Hpp/3dIcFwhQIvXqrWyV9Tf7ZVccdqBu2hX5u+J8XaRNcmEVikc4s3V8uRkkuwR
KdzPrRIvjsaJt+G5gLIoNTGwrdI2rS8LYAyKNVL+gI3VAE2Nu01CqxNTaPVpWPHv
pXUW3oLv9aKwfluWHV9hFqQqsYlWw48WkAXu7JU5CoxYV10bofCl34ZfE0PRJva2
n3/cQY3QNgjuDzEiLKLTvQFOo2ev1xGr7uVwi8z//Euvnc6kMFIZusyH+dXLWAd+
KFi0+I6G+2zle/7mivKUu/fZfG3GReXq1tKHvXIdn7FqXloyYLAeCSkTQniCLQiQ
lfK0CmX9F7GLIIP3kopS4JeR6uwhjmEiWZKkiqiGsEoID9B3vzderP3t9NOV2ILA
oDZvjxoumB/DNX2vncB2ONDKkqUjWnT+NT5/kHgRUDTfsRmqjKBLAPQ9hpIJq+Mf
MsxgxOuSlpWqJVAuENEZn6wYmST5qmSmpqODb13s80P7PkeWOi0F929D3/BYTS6d
uAyK96V2kqtLvhcd9yMAysLhLX1gxUTzK1uZ4MytauHtiGz4Wirrnw0YdU5T2gjc
Il0xhHXUTBTyajtqAKoc77EtKyzNomag2sR7QkGkwxYlrMxqIbMrPH7bcBrPwZFZ
lKKOuLNZuMmqbKL3Uyh4RcoEczswA9zDuH99Z8vSSdyYMByevfY9VqocZ/D9U4/Q
dIRANDjehaG4qHPy8piMitEjgJ12n2ChhtAoNxAss9XGqtq5UEIo/qRHYlINyg2r
P3r2tLlamzzdfqNzy1AV1NrhWNKAUIqjr7drPos2Sr8ekDlDk/Bor0mKLldXfXYp
OeZYKjchPSrYg2yjzG3eQ+z1KUv87pdtYmuNAfzDPrn5rNky1ZAtKdYc7hnIRS3C
YHEuQ84ZY0zJcwnE4ljHs4mxrhe8L8CcUTb7N1QE4+C8cDmwoeSgjz6ehEUVSl11
0/O72jfGypupnox31UnD5ezIWxxmDwDgMcfVfanRuKH5GFmzzs/uGmt6VcNm5WJS
21DMktAWuoyJk9hFtqnQhIcHR0Q/1pujXXp4duLvwAtsAS1RgZXQqz+mVy9eOFHx
Jb12mWy13wDpcHT9uv8K2HMTqtxKG4SfVMpLHZgTx4iN9MYAVGi9scn6paC1knZE
ExMkm7gAIcUhRVDxxZeynEgFBjOSRvTrjOTlubB/NNn2JsjkMHNLW+67C5n9pAfJ
iXvGz8y4U2Mu815YQvFMPGIhu3jUyZwPLlGyPWZRGwn2yJOy7uuonQofyVngJxzN
5If6EVybHt5l3CQoPv1jxi64o3WdqoLaaegAEevUnybeVOWwjg3Y0S/YqWSNVEqd
w3mFZzw6NUnKgQB7RNidtuKhfhQwbpYyGDytjAYJhdQGYiyTm2XDC55LYGiB9RAA
T54DNVMQ9IvtcZK8GVWNGCEmbUeNit1jG6Mp6TwZkG3zUeeZHTUrDIfsndt9XDAi
PkAa3xewloK+OkMJfp03l2D1qOPNAiSE77s6otxxBZ26hTM4IO9L48hrKBO67fOv
x9dZBoj1KqkdjFsiYR87SFcnW1exysZwaKuNqYK++h94h8OryulUrfFYDK893F8S
oKyTy597WwWKY6pMP1Ybpjedr3Th77qKAQO7aYs/9zBfyABj+kqToMSw3G2tTp3j
Eiyb6ANXMne3IwgZEn/FGE6hpbI9b+7NrF0u34s97uMg1e1MChejS92kpwyhxCyl
w+kRSVoKMGDS7cmoKd3DzEDBxAf5hja5c+8fIMPDojfqnikiQQH5dZavmD9Ac/gu
ZTX8ySRLaiWUrblVgtflGgll5O2tX9CTAtxIw8N6044kUBUoxITZhG8Zl8VDkN+6
Lks5R7CUG9NsSXTI0xUNU/NbfKqFHTCBgY2669Ekv65ngMoizqNXk/NAvd8fOQ9g
dh4j/V/PDYcZB8ldfaWQbuvMzKoT5wGvpGYwWOQ/qQxjJBcBJF0UxGt7CPzmlcU3
f0ueG73nUm62m2ADjAaQWd9Hhn/8uNa319q48RvfRs9OH4OaU8YFjs3QkYi8pb2p
apkrAvlhJ8SBDjUWVaxB1xFAjMd1QMHRP3ZSXKh7WqxzNkD6yToGJ8tna5U6RSfp
iijo/xvcK0qrvHQ6b6vBPI2bYZJEaHLwuSrhJY5HitWgJoAq3KBGzp6EfCfQJtqP
WFDPiU3cYcXSYRkPebuoixV9KKqlhL8nOF83HJkRYKe2DT/ruFkfBNbq95NMZ6qG
EpewQaio07UxxG7fnTI678nDa7E4Adk576gvjd5vI0JIttMy3+uGw+tQAt2bMUMB
/ltpvtCcrbaSFnJCYoOyqw2CEYttIMuinm+DdyatWmLS3zZQldaRphe7Z96REkNW
qKmUcA9YXQex0BSTey2dvAQqsWigEOcgZze+xHbGtEcXcab8TyegMqhPjpp3QN1p
KmuQDsk57vtTeOX5BG+7IArYWQD2k9f4tRvJlEGUwyJahGPJo7rTWtg6n+wcH7bS
WJpVmN8HhJSlZ1Exz9Ugh6P6n3n8fO0Sd5GMmxnlGzpu4RIPyGzHY7WNKlLgtWSq
EX0iKZWjclW/IT7OR3OuR7dNxhT1igpiAbOt4r6pg9xUAaIt7HQPYLYSfrEqdxA/
b7I22BRK56FM/fbkoffyrpaTgSdQI6uX8v0OIr0+nphw1RBE2Ux1VeiXxvQudX85
z2g+3tdhrvL10Vxzfcs9mY03IxD0aoYvnWjPThDGOIIn8O2YqwtOvrZWfHTSyNG7
BbQ4xo9rclp5Bg/K1nyvo10/YS0Pdk8rtEqC2f7Vlbo98TvdwRBLIOx0qMTUHBlv
8ngMW4kKzPkyJdcS6ZhCijo/x9T0Pka53D3s+r7wXIZ2ym3do8rvDVVqotluu/cm
7hkTkFkRU5VpR/IOtSxJIHRo0gMHVllA0ldhmnv42Koyurjn2iXdlI+FuF8pmlch
A1AYmtTXeoSji3gaYDqduvUsHIABR+Q05S6QVdTpOV4hchwhQ+QeXeCH/Swcl4H4
lPX/UzRMXCo1pHwMc+i/EJstTCAtfJ/0HKQiDpJ+9wbo0VdhwBU9z9NgKL6V6BaJ
zxDBAWM5VjUDhpc3YgiHHuFaPKyMV05PSOaFhqKB8G1ctpYTZHjHDOnEOCXIhW+c
Z4/IbH31zMHd4tBEXGEf9tCy8dtpSknM3jmyhj4flTBSAUa93q/qcNxcGdoGmNxl
stSoBG8ZETXHm6WfmXWdaoHDwFIlU+0eEVzs6wh1FufK4eSSOPDQ2EkaagdFkbPK
PVeYpX32fn4wNPWMjW1JHNw/q9EQWI6jMqyxareE1Is8jaHPAS2JaAhDVEwypNf1
wNQXWrLfYvLMfDlReHYlRGn/t7uqUl9AnSbvxCMirOLm00x4+i3NAn/FHCkX0ult
+LCPj2tnUwR9HwYGfFg9v5bcVNUGUyK5tC9FXFMy45f7Mw7l54kKRtBW2uC3815Y
Wu7Rp7DKxp3rS0HTZFrfyAnTxyqoSibZE8QbE0BI92yHy89hv+fcAiqmRmRgIUH2
/n732LONv1+BAhJgkY50NS+j83DFcsI1LJAhYu/AehKKSlE4jH7bkBZVaiSwqw5J
8GkkzV/TvcZyyGlFbC/SFt/fseKetCXCfaUFvMlcWEt8UaCvh3VzzPYLpacyuibC
JeL1PGqdotkBbZ0As9rvX6UYRL7yMX8D7Is/7XKeejk/8Bja2HXk6RuRmxxb7pgY
AcIbhNW5gVgLFMNlf5d7lAAchHyLvHQ478f0k+fU0ZoL9nI0Cq+b3ulHs9cjR5rE
WuZyLPDuDcz24E4dt+2B6xUfsFbNHY8xSp2kLkvMgSnXL+GdFzFWDZsivCnJ+bwO
M1Z4vfYfWVGg+piR23kLPsM4oN4OKoonQABMgWZCxAgjzqdehLTLZeaws0bHRRFV
beyiDeYtH4ALc5EC1Z7FA1TdFxVFg8Oy465zKOnqNLOLxVLP+1JSLxQgFBDq+sYD
qnIfE8Erq4Qc0S2bsQHkke+bk2jtDpDvOX62G3EQvs49a/z+tbfQyBou4i5PLhqD
Q9TP9DzVpE/032vIYi4Tw7chv2BksHo5yz7H7Kew5SjCk7919QDNlANenQwLrJn3
lZNvtHNqydEbGLtPbkgIDqbtznaLiNH/HEe7WXSFeb2CATdr63tOAbQNw554YdPg
MSLEGF140BPBcOVMUTjaRK6n+M3QtQAPY3df6Uqp6Aynv6il9E5DFBFQvuyGhQcZ
ISKADmx7bR3V1R+veYmuAB0OPhkJHbYkgy8srzxCcPdN6dyuvkmV4TCSVVuZjElA
qowMaqFa9djKKL6P4qm8i+K18Kixm7Pf8p+BGoq44vROyCtpdajEWUUjNA3UiY2N
hmY+YDRveN4fndQR7eQ+8Yk/FySkytL5BpCElFBKL/ueVrui65lYfFHLmxk4R2vr
m0mJsLfplA/DYkVFXC8o15QO3tDfPmA7ccEmt8g6LUtTb9SYJDCe72EcPX1b7N+w
AGP+fw5taxM2S23KqyNbfiADzI0I3XLQdWck7zy1c3hQitPKC0wXhtPIEsxRl7Oj
WKk+gCzGcwEWeVpGbaqi71YYnJwJfKjqXN6vhsfl4HriUGJLwhaSuy8I39UFOfKE
uL7f2tB/bhDrt/mMkKyKUPfIwiEiB+zJDNRkRAolvkptf8ECpUb2sxSSVCL7qKo2
kLRwhdUQlmPgsEyFTb5mu8/mW13KP8vfrfTeHQwX5vxMCcumLWk27vngV0qNNSE2
38cUWVMBH+lPFH5uOGCOU8z+fT65zMukhjvcIifI6midCiP4iZ5TcxUiEH2dcqi3
MqNw6+8Fi1dzn2SqQ/WSpMYS9H/KuTxavb5e4Ylw35DNJaKAYU8RsVPP2lgK3Smr
kiOX8jlSLRPrhMU1gedE7EhUBMH2pKNwFgjuu/qXsjJq7D6LukMh+oVkKlRog2J5
dhRXj9ag97NmYysckR9+fAeS+gruaIzdDY/Coo/k7A1KNTR5d/KRCQH1pYyZ8YTl
468cEVjEbDOiX+IzV+4AJvaKDW/CjuSjP2fVB2594tcgqkFTkCSc8fU7ioJVtpWk
yJqfR8pQC0N8nrSIuMM4Pi6jBeXUBZONVY8GU6nKCTab0VntkGHDlxbxGZbP09DM
2IlnuxmL1kpzBKxdHmirfxdNqCANHvCRA74Zt3trtYNttKndobF9zsSNQ/ItTXhz
fu7v3NHAfnTY9Rl3QdCcoQBtOc86H08VoE1tGVRWDDf0KsxsOsEq3ApcAl45sOeZ
ljxmEEg0gESCxDk8WXjqlly2cY7UT7Meg2mMplAJPCqsBaNuKpa7yO7OvtZWzBAK
2rbjlQJ6TL66s4A8NVcZl5shFmYEIbvSKf7vBE4lvaHNaRVIpl1mYAC3+y9EJISW
qDq3254gLbhezKTYEM23mz6GdZMcBELJeBIrPzqgIZi3H9DHgu+4l3PZvalcI1vL
fiKQDSgTDIJr5bvbU0sJH/yQGS/e1CGhEzfxJ+2dIr+/24VUuHT+6TWJfEOsuRqk
kXxWrYfeK3laFVQh4dc+OwJLcmIr3vVVVXSLkulG9JOboVKOtZYqemIuAW1Eeb6i
KeRavq4uRvo4IbYb9G0KJpk1VVP5f4OwHK686l4/V2g2nuz6bhZFUYrXcRQY6dwQ
My/Re/+h1xCaMzqNxL4G9JoC6SZazXtYph2QnqiU/XE0IVPs6GYv4/GIN+JbDk8g
qJ3pX1wwzViPn4j6ITTuUGgbo/r8o/h/hdPom7YDTirCy4WHa3hk6y8XuXc7rg+0
t/X9IDAPNpEuxuWjgPs02PSKlTyOxoaymxugDOgiRAsNuuDYqbaytVaEMh2yi5x4
IstzTM+1WSUtwk1z7Re/wZrVhuRc4PPPcjCOX+BxGyOazpEECOg4cKlRv9mxACha
qCs3SQcMQBamiOpYmyZQQR1Ca1FZHOcj+KuN6zJ/L+N3Ko3Hz451nNEN5xZjgCRV
10weCxRpHqd2l52sxZUMdKDdJ7kzGtPBk/3ArPmTmpGZhCezcbBIQdTWtiWuqzyb
F0oI7wQnjHUNgjjU0gIf6wAI0O+XvmHnrTsGohxhgdHhxDA5dG+1qeS/BCfy7Ac3
lIlwiobhnIoFmRswqmu+y6vqU0dH45pS+XM+HqGuMbRfyiAcN3/jBh8RBBB//uoJ
NGsq2sFsjDzLf8xwIHpO54e1yKVVCF0q+m4WlWc5N35wyNNa8RW9SZTmCsJOCf+e
ho08dJ6tWaotCkKzYNTchF3tGaOrpY9BmeY9yJbbEVrhy3ZM9Ju67ftRNGJeV4Jt
PVXnTkoQKwEj92o3Lc29vSklSengsuUeER53UK+bVld7BArdwk+S5S26ylOweCwB
ZEOoPLVrV15T88tENf6cpd36uHasJPDMeWWFIdWMhHkka0if/L8177+7wTtssmwG
dV/9GmltEDdvuCT1nyrWTNgjqffqrGgDfa887shgjV7XuHLYc13g58TK2Pq8oVyk
kECkasvHyT7sR3HOSneIMkmGolI3ne1fH3KpKrakHP9r4Xz8w19rCODeKdPrMz1z
Q/8gCRr+G5N/UuCMXahsdFkQDHeJ5bb44bZ7p3EhREL26m5SnFIk6JVy60/24tWs
dSZjgst4Twf/fbJ/Pd5gU0afKIAi4t1oZzTXfhY4rBJjrCslB/EsweErRC5QHaub
epXQgqTYiRzaklgddc6inQs1AlIle8oknjcJmysOANzagyVFnLd1zR5JUrdupb8R
d+lI3fuqM1/5zkzANf0aZygO7qNCw6nBr+xSeoM3hKVVs2CYe6opM29tgeAEvI7c
rzXgtOmL6TCT/HLrt4IRVTfpwLqL5Zqmfjt5pxFoxRaln1ERV6x/yr8ryeSkTSUP
jTaYTI57OvhnuDlAkGoMVEvyG4fjJ75vIGkxaOaXnIh/s5Xfuaa0IyLVhiGRzKOP
p/PuF+fGquPkcD/KjRU34kFBIMK/WRcrboKE8cd3llMdTac9JOp3XYcyw8VynNs5
mkwpmnHCsFNKfnH7upo+maLPkxIQLqtrvHnxP40501GfDozZbqw21AQSt2klLuL6
091UcPXP9o+k8CFO5oPP6A0PcTCl8bPHtljKlXmMLNSyDyeffpCOuPVYkkm6TPQJ
sLXtZXlp2vfMFSMeXaTUesrC8m8uftOJ4Te1yPIxeLFxbWKjeyQw3K4w5pbl4/od
EiVchM1o2Z4TJjWXISmd3boqPueEZvdlWUyMBiLHyrKR0wEaGefGJGmXFs/2SWHN
UJuzers+AID5XoTd4oXhMJXygZ+GAgq9xs2/9HvWm9qsEFScUga2BV7aMmQ57pYq
6ACyUnENU410HHO2VvgrZecbqA/nG/62XcuAY0rKz2nHwyqT9BTycHO4YFkUqnFB
EYSmtrEjcNTAZQgUgGqy9Ds5ytfVZGVj/f70GafBZxKJj5Vu/bZBvwIxaaZh0Jpe
LmvPPpMmpi3LtcmgmQ0yL2fEeM+8GGzl79Tg04jvkVc6vjnbfAC/5kwSN/jPZa6K
IJUDMwYlc/dTvAjkFoQDUYjqAIQXbhPIZowmEIuSLlWdhQbjOQ98RBEJ75s0SeRg
m4g3CGOK/9walHlCrprNNVEZLYrgArMUxFq/iVJMu76ocI6hTFwmwQgB7qUA6PRt
YC2M0LiR8XhhNcKHw6qnOtM7pmB8wMVc1Z5e79iaeyP5QJSHi1NkDuem+sHUdbGh
wPbL8lLH0J6nQzJJtgdPYPp1CKxYiUAo1NHhtchvcXDFEIF/2haKPsN6nrv3dOol
cIBfX/3mSA+D3AMTja63/Wmrr74eP07X6p3fz/NAJ3rZztptY3VM/LWE57Nh52eT
7l1MFyahkGEudavNPJxwzGJl6o04bw3nBa8lmAqUbPhzA604vQ2p3xetxkkX/kLp
9M79HJbNebZZkQKzVtgwzU67zkt3q51T3Ku8aSRwi44WoywjB+wRmEl2yQWNKB1f
v8mVi3TSsHtgXdRNXHeapTgzl61dw9OTSo4PLfX9lGFHUDygVr2nEgL8Xqb30ojn
G6uKAVOYKUcG98rX1rplLQb9c8kyez4bPuG+D67ABLoQKgdqotWCgtm/QJNe+tbX
/IFlTz3ZVrA66qVr7dAZ6yWNo/WY1lTlStQxXjR7fpYwDmYheRvwDKWs+N+MVrWE
+mpQKjyHDxoEYlcPswHBI54gwlpoAdNknn9LwJeeoDeV89hKeIvTe1QW98fgIafM
R0gngHoTqoR3R2on5HRfwMKc/izOuMTtD+gwOa2tg/ZNdrAigcTL3pLn2jghLqmJ
TwZBa+Am3sqIYgPCBdc4k5ZZxVdSkPaMmrY5WzMdW/cJ1oQEla8AHTAReYewpN/6
Fd9rEUUwIBacIVlYIM15qizwMu9CepnmedyIRz5bz0F3cgx/Hm3EccvZyMVBWm/P
yC/LkD0F6NEiSztYbiKeXWOdcaJPM9egAgMvSJe2zMbGHuXjWjkb/qyQkI17BdfD
QBucnl8fxwNnCKtVk9ZVwFbzCtnDbRLJ6XufFBqV1CGyxaE1chX9rQkMok1Hd+6L
xNm7BBtgCNoNyvgVauV78ZWiiRznv/1dQqVD8qIEuceio5Y/Ro6y4iX9knib9oaI
+0XzrYrAEddWReXemVtDab7VOM2RdLzMhf6fPCH2Pe3HI6Qa6/INX64iESPkjNgS
MZVD2rez9m0DZVb1arU+lZ+I0ybYXP0sTIpSdpDqrmGKNVhPEJBks4Sxd7njbwPT
yjnkAuGwH//GnjDk0BKzVuTmDAo4fOVi0qSUJbymTRJcWwqTotQpqkuq8s+IFyDn
+SlpvvV4lk9AeEUWQDDLMRA0DpK79IxV3jcat5iMfBeznRJw2HNgDndbPif8y8kY
trZu5tMFA9XqFYBVM3dYCDhAO/nFj4VFqIBbpr35UfcqoPUqxAdHA2BB6aTjTe+r
1NQtJqhizXfByznwgITy4lsBU+bky/lPuWsWxuXjH3zdvBPu9SPkMlB6J1KW4rxG
TwkcQST9egEPvdvPLGbU1vGXJune9idW/OcrnyHiO+DHKWC6oKLqk9z5TupHjqFH
Z5uBvQC0davYrjggLSXolaQTisiJFahfAHpftTLLQl1XLYiZcasNzhZspmqUIZgX
cwhFwBNuSTPqr7DQsX9x5fppbrbbBYv0mZNj/fVUgTf8rKL8jPpaOtDUrkAxu7g3
YGtqpybqMyF3/mAf3cOnligkTIO8W4kAGCBE+J1DmfcdLSzDjziCQCEdFen3MZ0I
KM4nzmQPvn0dbunY7szoaxVoyKDXg5xbJskCQ3LLEdy9DrlCK6esetDxiSv8R2ri
dv4WAjLi5wU5dkqeKnftDZA0tBUTcVzZV3ro7KPsCYqGHfWCDivY9T9l2mqrEdp7
aAEFeCD9QTV2OmNAIC7DNcNP/3+WtubpJj4ppb5JswRwmJacEb8tvzLckrT2BmkC
EKL/2/1DK8tzNk3gQWjqTtow85+Lg0v0mqlC/Y4WBoiQI71KXhZx8BMdtLXKW6bY
HjGIVP+OtyRrcCUSm3pPayfnFB+Ml5bUA7eOgne4c39aOijwZ2k0K2S75xoZTDlE
iEHgz1LvZyaSwyZrt0CU0uolvkjVi6kGhWvLiZ6U+RMznv1zGiK5LhPuvfgBOgRr
oBO3whwDtjKoDlExCGiGoNV0IEjL8xUHDbKBlO6fa0CMv26V1lUpZpiPfe0RmtF/
DZMIBhltGDZBoy/zcU1tQRLAEbYQ7yeYk0jdvcUMw2AjwScrM7aOrqTUB8O9O8ah
xJf/9NBB6kgcwVM3uqe84DrAYudF6Owg1pR3TBlVzocS2WSOz+gCx4cvS30CvfEL
q7C9P8XuIkrvsISUgX/NLFTv8RMLrFp13A1d/tncUl/zNDY+nS+hkO3yipQ6h3oC
yDAYPRg3rJuGIPeNnQi14D8LfLsIALwsh2D0THeBw6hL1XDO1BQh4QAGlLTCJjqz
r4TfTAJlklOcF2ktgUtq9frB3HKVes1imqNV5msIK8PRCYnQN6b9/YRkVgGeYsCt
/3L7cSgQHtuhagGJybWIvG5FsBvDcSK41wq2VAo36DbB109rh2cQglN52tWYxL0L
ysN6uvv0gBDmshDiLG1oJnNOpwD8Xqus+PqD6/spdbR/f6DcPdBw/Wy0UFcL79PT
BHT5+x+yvo2dw1C0Ulu12ZosksOFQ3mc6ECqygxdsv9oG3ucNwgNiZbZYOkBsX0t
G/aM+rPWMVdzsBpFzNYwJzOkc+8nhOqaVPOy6GLJfOdBG2O9Wm8v9SxPMCpIZQtG
Tg0di/ZWxr+AoUeIAa5P+FiXEUL1/gwCT68Mxt8qqskW9aMgYAKQqgxGQJcU8h8O
iyLXfnTyGnVaHQK9tWHhWRt0Jdl1WolWHb+bRCErQxX+y/kRDwe6TBxocoBI3WO4
sNu88hMDgkxKiRMV6s//DqwwrO8IHmN8SnlU1OA7j7q8Y0WysiBRFQQw55IFdKgx
f5y0R3LyQaBR6nlYqpgoOD2Vk4/XonWLI5KEIkJ8NfnPcJrZupEjz9zuW8HxUDSl
qtjYwTWyEOIpBnuKSxc4DVvUI9V3ns5oWmnG3h0v3rV83Tn24sPqahCX5iiqaRAf
l2Fhwaa7MxJzdtcLjkPF3t7il6o9tdupeSwZPmr42tlwXad2LmU+cMNAGkboaJ4f
z8djtKxNxxOik8kpIDIzQWiAdfqXHG76uxzcCQvmN+Poo556NIlQCK2h4WhryIg+
ram1tPClzVHT6yCYWI15sKU6VeAr1336RuMqLMEEP8cKW74IPUiJWFem2e/OSI1d
opHBrAvbkgfu9UJlrygQTFlTH9lFt+W7h7rgUG5qo3AAChOS3Sst75NHxK1LMFzZ
66fC2H8haIR4/km6821a1Wq9q1+SqBXbPwdS6b9eJEaFrskA9Tj0VkISoaF2zYpb
KGgf6I5CD+FgQIJSbwAVQFsn2xDFvDCE7O1qwJcFBe6XSloOc7KVOcbpBSjKeNw2
sZ5jH5oMQRWrVoD1/wqNmVm+clnUu39qWQIRcGuDpIgBHYjpvOEFbPV2EvD0RhwB
o5Jw1APsNBVnefKlrImi6xbrmRkVJMo9ddeu8YsOgXWn7R+HFVCV0exhwt3UwPar
GAZPeJ1/hQj/Kon9/Oz463RCTXxJEO4OjhNdvfrx+k+Ftb+l70I0ZTkXWsKrWxsQ
3BZUqMdncvCjf6En7np9k7eCCR/4WeVydARyBJSSlnX8qPQIHLvTAidZnpzM+g62
hvHz0LR49fl3v+MzGe45s+sfYbys+igCDUkLPx7gwuuHqjo2hFnSVd79LMWArrPg
CukAC3HyS8J+CpaeyStEfbx/VV0z0QjvQOgwULeKmofhx24HbP1WKNIZ2+hVUOOo
xCQ/QePpahBBjr8kKxZF5CbJ4cB938aLxw/Zelcm8VGpe2KptZFEAir2jN3PXLKk
zd2ttPTQ4XtVmvckXwERmg1xkouO7WGVCBisy+OKsAgCjTzDmjNcHgX2CBIESQ4U
0+rzZZe5U1JubikuQnkYDjhIkzI6nsDgi1yUlBPx1CSpu9j8SkXhFIYvwUHUyqgS
6v+XBn8vVHODJ/rBDjo2wAks+RbWgbz3dKsIC5qhYUQBMAdsTSqqVi5iYNYfyEat
WwTRflLVTEfgkPj6SwtWI8cFjdlK6O96EhStbiyX26I6EaYjjDXshrc2sH9ID2rZ
N6IfQqqHd4S5mxjKhmsPXY8zEezKby81HwBpZxmI3eLwcqsh4KbkNSn7+bVjGOHq
Qj5nOBjp2oXDZlK/0kmKd3iEbHFBABZoTaIhawC+BmLB4y6YQmSff6/20jO/U1s7
TEqtGb8MWM5yfTzY3OFSlItuLK9Xc8aXu0eAAcUQqXD9tgRQBuMz9zb2iGGoY6Gg
p1wtNcJbuiba47jZBckWd+D3FjTXe6g0MOIxFhimp3Es9jgsuEH41RiRrsZNJQvE
a0MbOvybfywav47yJzSc1qVMa4pARSqafjp6++JDZc1uqMBCrnYvstI3UnXudZDE
kzcWYJYtnKlg7lTRvcyiTASiE5kWvoNsFNDjX8pfwMCmzufqKUpKT8/1fahTMVMJ
cj9UWGE91emMadUVSKgQ+IuBUGN3B/cPsuy3DNFPS1J9iquCWPKMWMQoXX6OLAxm
t8U8wgk4So9MyrgTMbCyGQpk3Bq97oUGQY/HhfmSEGjCYZZzOAeSePsZVCMC2bCy
ViqgMakBNy7fOiBHyYR0sbjSkBAFkFaN7Hbw+vsdNoY84SXA7dhNpc+rENY/MsLg
0UomPHR4f/gWtKFh5PZNCqxtjFbk54cfNDskd4m+GROIRjTgjR0NIkA41QwbOtv4
1e51ctV9HZxVtRssMTEREzer9oCI89hISZY98ckYYpqJ95nP7Cojk20XTUOSo9ge
Wseu8b+D/5HY9SDUkGek1UUBvnXZ0JgNjsqF8qBSjeKpcpBOcOWWzDR36DifAP2b
b0n1ZjUYNMI1xNrjE1tC0cbtWNES/kOda7AYUijYztNlXaEonTNtQ8fS3oIv9M8f
SONmLPLPiPyWfmXeOHojVkAv0qOmM3Njo9t6KseKAj9QxywppRAEotwZB3WsUK3R
4Ksfz109MUTAKbbKYxVkFmLSeVaDXlK4gHvmu5cNTHYIDCVUdSjGp35lEXm4ni3s
pVzfatNepcflI/oCIXXBzAyiXgk5KLHbt0X4H7pAXbk+CmC/pA8AWVSdmsPFq4jb
isYYXWqzaPTRLihq637XeVhd1GdccnFc/bT6Q6RNaGRhiOtmJfAr++Wpj29uFNiV
CJ5rCE6tFHKLv+Ze2fcrGjcYcas1G6ULEYg9mb4T7QwMxj+/Cnv3F9qufa1zBKsH
bu2ALsTyV49APcpF2dctpUXkFy8YzaldBee1OdBE+Ie6sEVvwWCHvZo3lu1rLpcX
sTCYjghq4TfSQDN54hZ57GGf4vmq5J2Krypm9bt+b94MkDIPkGPwPW1Dizu3FafX
FNyBKXzAoAgwMWwJ1v/QwFBOrxzSvYKiFUZ8dABzfOmprrOtc+GWEs9eJy3X3HEb
AmVMrzwY9rh/pdw29OuqR1acpqEc9q8ZN7+t1L2Ijs1RQL+eRE2yU5UQQEgbYXA0
WjL/GpP1CE6OEvHjut0Up+GOO5bqAVy8lPOgDcBNqI3H0GcON4megZfkJcN7pKBg
Lix4u+GN4N6mGMV7U9ftamm8wA2V6qnQ8B132d6epj5i/HB/eI2IHdsrVjHkjEH0
+gXR3X9BGewD5RlOOBg19eIkkbXKnWflAcif1FkRE2M4t7BR2I/2QTAvLJYblAz/
Dw23LHMh2XXS8IDEMn2j5K4IadofEjxLRsdP38Bmo75ObuTVodlk6A7V1wNEWWvA
aw0fRz4gHXK1bFWx8wQ70SKabXblIPwVt95n6fxEj7qm8giEe/Mk1supMeprbzwk
S/2n3ZS61KF9PHBNdMgMLVj5/V7J9xxJC0O7Bru8mITn8DWOp6D608tLIEVRvdVH
tVbe1Zpqqap4iQpl0rC83WGrODQzPg9swxpMwlPOE/E1/FXbQwjiiWEm6tgYRU00
NQOTtScUWq8gZw+VYbjuhf8gms6BN4P5CukUPFwiTWsOimOtTpsKr6QnlJ9JplPn
SMmZulVdHpgO40kxRFKbWqE9T8YEh2GqNX+jaFRi6E5pgSzS7p8BDr6eqrrHIVDi
aBzdmcKLsnOWeB30TWEQQQzBjsaWiRTBQGV21JZ8FIiBlmilvGj+dqqEXyglMiRX
lUSgki8GWu8TJxha4pL7ENsZJ29ZzwA3c2LTp/wzBYmxL2n9PIjWAUk37N/MyXKn
MnGEOHavgHEmV8oHcKYUkHlZCY14eQjY1GB2wyeBqIwU2ithtR92TLPBQ8K3vLDK
iZ9AG/0C7Yz5cOMIE4kdgdgp3dBe7UfXjVNuLcP7w2Gmh/afFyOIFiM+NW/TFmhI
YtffgdvcUQUDhhsJbk8+7/M2DuwhX/5aaictciNqX1hOY0IKQUIKNO76Wb7li8gy
9hWYdm2ga4VMCEOKT3e7d+ob3RRU1t1iof3wugbU9VNREUEcLs+9mil5b5Ig8PGC
dbq4Z9au5wa91TKKZl1+dUSPkwuzixAQJV2s4DOrb8IRBRNqah6E7UoKlGVjsjcc
wt8dz36+SlWtkrQqh5en4zuv/2/bl8iHWcjWqt+y9kavgx75tNf7pq4dMruOSgKS
uRn2qcD/vUC3oDRcNSKrGXUoWkDdjQqVY67Pf9yTvGfeADrehg87NceqmCQFIAqY
mFp7CCMq9Gv004zx0IVD7JjjcVzhnvZGatu4kY0Q5LV9dhUjmljxZO5ZmuoXXOz4
LSrYd41sX1WZvINuWW3H64PFdWIAHKZWAXhOu98zo273wt6ACV/7pn+fEeUkC9uW
+M9y3xbNOwlqT44bdqHAqRe40JCD4JyvV36sv2cOLqdwjobXcduD4YFBdARM6oQJ
p6FCmUmWtVkViw6068IacG9xUx6fzPQKpcRIX5ki7Sq6z/9yaE84tglVi2zgDjnD
d8GV8/HZt41JNZL/x+027w0wxhfLM7cyiSZ7SGc/htXm8eUfC/z3OcdeHMVYqkA3
cMnSq4GSnkwIfMboRtTADbfE4+VPJYyn8KWE91UfgV3TfrjIi7tvZAnq6akEVv6l
1L9aCRvh+GAsv9rqUvXOk8GJnlMWbXDYdDpGDYDgF6zWDn+XMvMoLeUVKAGBrwsI
EDXdNKbBbQqGOWDmZinQ4jALzZzuHblRSt19fll/Q7AaJev2lig+rD+KudvqDxHy
u+LGVijmF/g0nuROIqov7zvhk1mo0vEVzNTZyPsKtrG9uhY9bML9H3rvqNMtBDnT
kk2soLOEILRpcugu4+KXGmB4DgOFKkKK98B86qnit33sQky5AuKEpnbvtZIJJk7v
OBOWDliqdHtOrvYSm8ojWBa7a177ZsLK4AfRermxCcAN4zQ+C6QG8KbE3a7hKXSQ
aCLfT/yEutn+0ACfzOaUfq/KB2wf7UqsxuoJbXb4i6jmqETfmQodRYM/PtCte36Z
1QuNnguDPWZKKDfjW6HbrPYh7zHk8C6kShvp1iBQmQ4WKGuSlvC1y5noVg2lg8zT
3Lf7i4wVaArN3tb1Ka5EpCvmSMrRao+oquabGyECFFZDUkf2kJTsSFO8bGPd5EIR
yjUwD3+59e+FZPwLSOM35o+k+gyfGLYg0PknS22ZfLzG+fmQY9sRgaZIiTRLC0AR
g9qGac9QFPMN6P0+eH1hdedhUYCD0P/CAmMb57OMmdf0e4tzh7F/xbO6L0PI5bsX
lpwu0aT/dHeBy0MCfRMb2GZKzJigU1oTKsXQqXdPQcrkvTC3BDzRK84BOV6d0BZG
kLv99pEdLNXBF70oZaq6Xq/5rs3osKTTP8d4PyIVpi58tnTARIpHfGlVNJMnEN/Q
krzqzj0YMxzBzeQaEv+ZZ87W4tpU1GmZ/AU+5BbieCudzAVcZCe9wLrKxA9JhxP/
CyyEpxYGUp1DCw2fe2C/HQfQ+/7Pk4xxJOWdeEQWkk4eXeivLNH3KjDDgG3ZMTNG
U/0SNsMNZj79Ft1pjnYW46A7z+lpdHmjrOiZyk3TOkM5i1xpIwXUvsBcR55V1RpR
3u4URLZHxjIjcQw2UE2IxCe2ralVi+ZxtCFBxRqmedumb5btyV6tSmp1Vnn0Nu47
b35Mm15tB1Mp3sr/6JM7kgv2rYpCsCif1q5Bz/+nUq9VCYTQJJ35ck8ojopOIVTU
+dH+eBpnoRuKOOxzluaDWbNry7hYx9sOmIBJVTfEsnvw7O9T4hOfekSBr5ZK5hZj
0+0xDJFkzWruTnqY3K0IGTVB7DLBqJBWXC2pzX/C+VZzb9wwz4njTOtgYpNI1Top
y7kJ+KJZa2ecyqgX6xsHIKddIv+qTPwXPElkjMdJ8fXCPHMgreFmU1bruSQ5We3y
3UU20Rvm9Sc5/oZKsHRgYpyrZ2+R85lepORYucZWGJpK8Tdk/rDUeyg6ulDd8SCr
9jwlO9t1r2qQqrU0R3KH+zmRDRDnQ3OvMCaj9dXMkawNZRVTxwNHNlciwsiSkZ5f
e4caMQN4gXgzbK6aY32svDswmctaKsDZWfcduhm8aY/JrC2C/Zm6pn66WtiSI1HW
EmHmNEuJk6+JPwu9XrNjSVPaiw+NFox1gC4CnH+2wl+RaDdFrFUe+jfg/fWjYCWm
2oqcbY1cPAAupi3ECl+etcUwTavcqylGY+84eQh4K2gXDKlc5C096WIcWTKL7qB6
7OVLEoLbGiR/c9wbffmslsXKoh3BK8FZJbzwP5L79T0oSmAY3eNgE8T7DOoWUSjn
oou9qbr8HIvVmA0cUIpXkEXH9xnLQfBH6dyoKewLiyo92IxA5/uOy3rk6yCxAiSn
fEMadcafXDKvV6NJ8hWp1TZlo9rO6G3t+yxBhTHptvtooOe10UVEurZZaexdv1no
Ijfi+dx+pmypOoRC3XINGCs0Vpj1FuAul6ieszLN937OR0zFrQCLTmwcK5moahC0
DBjQ8Fbec+8CIQcmeLWx0ZHD4+GPf5LGzx0rL9RlsINxBxFWbqPje4beD0KutA5z
dHLSfYTtcK6kziYQflkxZt/9ghlEOfZrBOe6rv9/dwEkW9RRVu2W0jlhGbi6+VD6
suEkdgEUsv8+hzg7Nu2h9J7dA0h9qtjbiHoJDeaF51xSDOmhjylhEXUvgf4yPaAF
yaKg51tgkuw5YYaiEfVMVkF5dOZCL0K6vxzKImddRpGravbL9xds8ApCoXasvet9
NKtmbecv9tJ5YEjeLPGwNj5yMQawjyEn+R3758BEiy1lzCVsiYU4LcGzOle1dzD9
8FCkZEtwK+iBB+NC7C5IdZM5f5MNkVFcjczVWI+LcUjBsKLBhNxecw7EI5QMa7VK
k60ZehGifnIyQdZx7Bx5GmMFZPRinWn4T6kxmDeRfbKEA5adFvbuwYpviUztcpws
LDnUymHqmhW73h/iv3UPs2kABKR/EXewQRfDHV3/yMJVb7tG2WBy60TJxQc47g2R
E14eDeVrfc5S6gEABRocZXRZbr5kfy4jrQj0S3XSoqmAYlCcvp22Q4OSih2P4AJn
Nk16P0L2fNgYFuslDb9EG/m9p4NtWcUCoZYACiOnAfLnVxHc3qUeGCPFh9sDcE4x
dRs+Q9FHzat6dSSrbiJyPBX7nXrMkeWnhCd7Zu/6fSBVG5CD75KUHg2DE/SCIIAS
Wyg89aV7yPABalp8V2t+jt/c949qjSbESHyuxS4mMZ+7RJq4XZCyfaNFRDtw8iSh
ACQnQDFOZQj91nVzadYkrlgxVdCGmhzWH7RHXxQeb5OKvgqhEfyvoPlIqtdVRiJ6
tBJspzWZSw4db/VzlLxBWjErA4LsVfBxXzExYZGrGPboeEPTHE7nHZvUd4Ee4PMz
MUrCBFacKfUEyDFKAVp98ZWcXPtNSRHf5kFcANLoqRXeDOiBOZ8uXzpgS0QhM48e
J+iITTr8gQhy1+gdnwFDw1frsF4A4axj9s29hBu7WoFQD7p7kEetdlm8XjrNDot3
opkFObHZNv7KXy33jJ5iBrtwkPtkscG2A+YxHT/DOtdUJshQ2YbwWz5fk0uAjnfG
9ClnoNwFiTdTvJA+9mBz7MHtHnQzw/RO3ISL5k8R4WZUX2tIZjb9btJ8D658EO9B
+CHB/apOH3hgUxpCt6am40hgYPw3e7pGBnsM6CYve0JIjFULfiF1N3DKtU6jmElY
6sECZKuEnvDAUiRCRhhVtCJGy5g5GhmS24miX8a7BZ26AfQX5z1MbdI8qjEUo6J+
HgMGNRnmpLKIObHX3ZX5DanJjh8IrWKrEgMwnDAwWticxWWmjLJh/ANwtXBk+KVU
obvTgYbNdxirbqbgwuG2OS4nmmgGA59MtiXHFXSoEjFxlA7GTNA0vM22o7lFnRcB
S+YEbOXk4n5yeVT96z9L2nBlc95hZ9hm8IpQjHTGItE+ACNxzqvdgthGzldZjsRq
oJGMn/COOCTxYjngZ0A2wbUpk4TSC7nL00dYa05agqEWPk/W8jZdHdbnSr7nuB7o
D0zCU4jmB69G5F2yo6F2btaUNL59UChlUUdDKb4M8VZgoSV+HAsacDEEQziqhM5w
8rFR+ErL6ZAbSeCjBDtHbVF3UVBvhPrWaIc3ybfekhRKpTQuF/8LmRDNvZ+GN3jT
icOlQwy1etEOiyW06dPutjzgeflJl26fo/Hk09hz3H+SOqbIBjq28yEtiT3Tre+R
z/dtdhNGEC9AlbxhrAYeR6YV6SuOh64oHS0xEkfZ9fNqW12BmJ+rpiwVnPW8suBY
Emy0ZIhKo+t7yMMFUnbz7091Io4fPLU6p4MUIcZYEeU4hBqhtz/Q7YuCTACwChxD
VeGEarHCGaAnwI4OVshQdG5Dnb4ZqlSvk9E/zOspA3ugytjy9gc0JLRcS2MdXu6s
SzD8C6yxEY0rYvndqbzjiTihzMQVOk1VlgDdDVeytivwzJJ1eNH3CsQmQAVRr67X
eeYP+6D5a7VXSGd5vYHrc1rsm3P7jg/iI4xpSNCtw1gw1F8Y0MHMYAhx0Eixe+cT
9Lqdz+vyttl0czmnyhbAxpg0FC/+g5HP6LekfJ53e/fMPCQB2TMvOvSEoSteqiS3
R2rPypQG/2rSwrWhNswZ2e1bbZR8lKmYm9fmwGrMwhd4dWIg0FYa8MUI6BYVhWKn
llW4tZn7FQdTEsdeMY2Syp221+3XbmTfVkQ0JsbjS4HmfAEzvxpUC9AWfsfIqmem
1GYFUR9IhgmADo77o5mBVfZOLsu01XhA5MTFLhyebkHd5xdjpTTBmzdPzNF9gKJK
G0xC6MfnTTRlJtIapugXPJZ/jEfQcck2ieoYxk3qxsxVYURpnhpLMz5rABO1RZAY
miUQ8I3hhBQbkt5LiWAkPC44Kk4NVpys/qaXaR15+4UjYCX596z+GO0E1OvC01T5
pPdvWBywLXSOWltkMTn09jHn9AhCWibW651kmXwLgA/khGMYzW3jEJS04Fl92Ofa
PKxmkzX3Qcdr/FJbEcjp6PxAv/c4MY+ZCl4wcQHeTZoqPXF8WlS4xITg4b0o5c83
5eEnt+oPYoSOr/sqOTm66ciW/4LmH9Vtv+P1sUeGFhLSJKRWnwwz+l/fEFmO/7S3
T/a8Wsswyk3SI44hdw1CnHLnCx+mg+9aUEuo+MjanlNMDGWDHm5fPtFbY7wIRNYe
RFKTqKSgVHwe/w0G8aawp4ttTH70cXnpl5MwsOpPP8nBJO1EO5CdPCsBvRVS42Iw
dUB415hEnyLnjxJQxFYZFrKnF+zb6irKPl3C/x7W4uJOXn6IxT8WzT4rQlOTMZZj
SaHqmV3rfqWHTGr7q+ti/M7JcmxhSH5F/Hk3QAs0KaY2HPeZFAIPbPOKTzJGB+iF
u+TBJFq4JHnY9ZUsCMieebEHXPOf9+RkNUPq6dnBx3qJxXeRQe5Zr0+IQnkpajj/
Cm0c2GE+U0Zrl8tT2YDrgpJ6tvP9ZabMYJl6roJUY3Bx6PFXSLLJOc03yg3DRyDQ
PyWscjaf9+2ozFeZSuboO4KNH8KsNJDaMvoHMQpt0tWHTBOJCJj/yEkLWU0BD0UU
3yE255GDIlQ6jxxnqCu76ONPPaiz8FW95m7CgcKlsiFMoGNQVd2exRgjX4YzQ/pL
SCYNsgh2JXEq5nEYu4tg8yvmeheN1214hohbxP1UMjOEA+nhAwLWNmCQLHZv5Mxf
+an6TXzCuvxLQlhwEmMoZrc2lOoNt7WkH7AgEDuYrksAbIuUnDKof3rnad58eRXU
RHtXPf2tb94dRVzzfR9kHig4+CQch58LWfQHge4OljOiSCyFZVCpOSkxAdk8S2mL
q9gQpme17IArYi/bl9El6ItGA67Q8trokTQm50VBJmZwcxTTAk0ggzX7GG+fq1D9
7Twx1F5D2DjA6lXIE2Zt9FRCoE+6b0YX8A2IFk7L8IUuE7n0IOfLL8j8AGs4zAuw
NNT+LBtbBAJRrhuWgcU6ltM4ceWXJpeRhCRHC5qs0i/lQ6waIhzm7jIV3xL/fyWq
VC09Oumuu4vkKF8LPbLIOuyUhdzHVExsNNAwR3M6anUfesUuYEHL/IfThfH8CcLJ
RXxvtv4RMQmbqinaHCKgzUMS3iKjrA828kElOoMuqrMGgNMyJNGFcOf4trwpNsJ8
F3qDbwM0FPNJYYnVt0UVZN35sackxM3v3iILVNM2OhS27ytkZcNY8UbuU7l8FWoE
YgAhMRMmjBsvukG4x6PBOXd5o2NOVbkLy1Yl2Pljsgy7JTl2g+XMvEaPLPNvYpYE
e2077xKaB3dcp8vfxhpU26/7QJ2DrPJPdimE/G1bwvXUu0v69H9RZL8i0en6PjOr
qiMpzJydNF9k3XgVRHYPKC6cI7Adl8uMRd4yXUu4VHt/wrcse572Nzdf0m46SUfu
EjytvRWHtBc8cOWJfzwdIfAqf7eHkMgcIA0CFYCHRtsPZWuvqRsoM2TaX3PzkkHl
St4iqmXhfFnDubAohNfEEYa2QIw5lQQq+omMPRNdXrOPUHZsZVbZDZgY9EXL0INC
HB8hKiUtuPEvqKSEKVDMJfMdNBv8wf25yz/ViGju6cvTxwh6KYjT9fKrFSXtgqh1
xGUYL3AYXgshC0i/ndlc5xAKHE7maKYJEfSPDu3dEVRNjYrTxhjb4Hd4zu5Idnf1
ZBoel/7K6sYC6HTHIGmfgOgU4Y4pa36oYyW3xFTB8vRMBrVawZJAlUDqXgNIk10S
QPyl56Sv6FIeSBzGyA7IK/k4Y7tv7cHtCwO4TW310guSGfl5U5RzwJMIUgr78Os0
E/9L8+cvMHBfMrNIpAo9Fwa52PmvPfTDVvAOL60YssJpKDkcgXUm6CZ3Aaq4OxK/
8HaSxlLODx3742axBNwguCPsDrs25+h0fMNnkj26xP/lLwBOjVtaAthdZECl5BVc
RG34myGTZ/Kq5v62zU5z40Eavq+nESJ1B+VDBc7GUnTSbRScHvmzSas/4TtT+23j
JpgRHN/c6mxDUr+xcg7y0zEW02ZKMubULnr7/fHydG0JGjD4uEKqVVIS1DZmnTyF
23KNsvIjLay8tcx8fbnkRCiuWO+wcMba6jncHJXnRwtJLTJhLQpEXncHRF7xjE5v
xwnnf82QniKyTHxtEuRXTevHA6jz4HkRTq2Clt4ulKtIZsN/NXqWMh2j5Est1Oy5
wE0Xtw/E1w1+p9BB9a0Qi8WJimo5/atXd7HSWtOORA41wuM3iufCoP3pq0FlWyjw
4H+2tUBJ/Z2DqsKP46Uprr89lncvT8FpM6pCiA1ZCSjrgcQepKmpZcotbHSNEoFV
3l0x/Tm/u5wLN9F0HwjQvV6Ln/5UGXrOUmcL3ZMqUXtiWm1kJZbsbqJQliDd6uq7
gy6X9dviNSIdCYK3rIAQxuCOFC0z6Xemq3dVnFAa+H4OjEcVArUyeDV+qs94ncVZ
N/9NfpK7JlkzjWYMk0xQ2fnRa5nvU9syJxorMZ0JHyH7HZo7k2f3YA037xsi+5HD
RBhx5hE2CvktTJ1ykHmvUT3JFJ2Z1+Xr9/CtyPvuJpKgvZPbNyHMhK4AtOCwua6z
LT5zhU+IyIXexiqXinl9caCeWKzc+0ax1+jP+b2np4yVip67/TeaP0EOHXnQFP/j
Ih0iSXO6eAg7Q05mHWswY4x0yWq7FJ+0IkH1ZOlmS4cScKIzV6ACNYtM0uYyRA1A
CBAs0fxWyahDjkktjr4LOLdkahHjkpAYlc0gl2WYGrjPzfRCx6HT95c4HWI/4I5s
U78QWe7hFovbrHf/AS/JrR5PgqnGbgGWg3Y3TbNZmGadoMc8DtMUQC+DHoJLSWax
599qp17sYujPOGG7HNKz5DC26O4y84Q4ypU9LTMkgiFWMMalFz+NPQw1f+eqm3b0
JwntykoY1rgYvBphSXhUN4M2v+NBkWAayPj1G3r6OKj7WHEheqvL9cmStVijY2Aj
dAQPnu7+3VyH8n94PRYzSBsgR29IRm9s7meR+5VxXKZoqh/YPDGGlifK3FIEmgr9
q3ag+1B23pscUnAkl8BF+45veC6H91y4VWioarSlcBmvPPOc8FiPv0rfa++iCbKz
QYx7qFTPFGCOdGy9t2bC+J7iAld2aTifBF21K93vClkOZdYgeikqlUK68nmtNyB9
naqEDur5n7hOwoXol2j9fVDIW5pD/nKRZJ3vdBHsw58mE7NuzFlNOSCZcGmkg3cx
fSYBeyiMGZ2pYbydtxksbSmZnk55OdIUoFwx/cLsHADXNh8IECVhVsFAcyxbg0bu
YtJC0mfC2my1e808wmCP6Q2Uaf040O/PNzghJqQRWTXd7r/rk+ATA7T9gf+P08RL
+HQ5OoezdxqRj/mSwnWU71NaVG8Mex0MNxkwUGyyjMT5cSn7OVuO5oizsP5yyHy/
4bF4mkAjU56KUkioNIjb/Msi4hLSgoUFQEb5CywwzPg8iadMSDuZo6AZdKIe+JYQ
iyUgjB19u62RSjeTRhYuGM+f1a9ZIDBnHTtohDgdr0oUNe3sYkhgIFtHA0vEyFXC
mGETqwwh7zDt7iSzw/00ie0SsJZhCGtznnwFUVF8HAGnCwsJ2D6BkSwoJ7A+YsVs
zn1e6+sJru1es1aos0/joCbjM/tx+7DrhvtyynOJBFFjFUuVmJezfqQPyTuEq1n9
qknUOzJ1baBCcjDQm9Wf15SSdQq0oXenafatPX7y8xv0T3VrlhwvkdLYwoSDNwf6
EC1BMex9JTzUNVO+naxgYW9377O2xc+912CSC9Npx3wWSGF0SjtR5Kvy2F4FqF2d
UlRYx28tRydPXjaNQTlQsZy0LjC0r2r4wXNYBX35Oqzov4Vgb2R3ckAulENblspN
Cxc6kRMjsD9vwl4D1IF1QWeXspskODSBetbBheZUcD7+ixs0HacwFF9JgXo3lIXC
Ut86Cw8rEhFQzVdjrLpkbh9XgtiPM0Dhm7nDE5oO6ihnfIDa6zrP0wUmFb0qzuEH
0ZoLeNlSlT1EEo5ZMIoZLchXbdEO8pbk+K08D9HuqzYEJ+YN7iwHn5MHZB2qnvIA
jYVlRb/bywN/7h94Tv0wznQPCEukjB3fQa27TzkrrldNyXtUmQFPdRCCU/5iX+GX
5ECnWB66j61FPmoA+xX9EcB3WTQ/l0rw/E+8nQDUuyLKU30Z9npmrjDOz4N9NMjJ
pdBW/J7KhqLQtJGELoyom4TSENQ7mvEMoN/iS5XACMhxl5a8DLPXFTsWDQyg72tR
0xdp9jpGWFYieFNrypl2QUYmnPhAKScU/Ab65buHlbX2NY0eOJphEaS/gU9aTl8N
K/hN6BfWoa+nh1BCVBZrvKGST7nKdrh8avQlRugGsf+YSq5X3AQfQs3C7GQwKLoe
195h0thMIrbWW9U/3M4/pS0/HVl0+M17FcJyOM6JlecDojUpAEVtL7L53RHwklvw
QK/Qdg9CrLq60ZSdTTgV7hy67DqQslQ6ZsA/ixHAGD3fRQEO/IU570xNM8z29VIy
jBWUndf/d/fdytNFfKS/s9PMIhtxW24dzW2TXfEopZt2ccTO7ubFpFRBIKJcDbA5
Rls13B790VOoces5xV2v15ncbSFumUhhLvHvKxyQNbltiBOuJGF6rgmtoBblj/y3
eexfh5WSiVurhtN72CK2AKTh9afwkxcyzNIej1EFuhn5QzTuOhBYrzpxjlE4G3o+
VYAZn519IygdVfwY1RfFB+Enc9KiSF0Ch3vZheVN0z3k7cV3q1oiGkeHP8pweQI/
Mq/qHRM4j838Q4WFRadVfo7vC/2BYfMapjmK0TDUn9n78olMSCiQkKIUPkAbCO2F
8+DsEdl65yhQS7NYnO+lPTOxYLxOtYUnojtZtIYt7k8LNFO5UupY6/WWMT9MR41H
3X5YKKvB4uz6W+CgzwHqESoZsAd8JDvutwPPwzEHnPhIZtRGjbb1gCRM1Hl11MxU
SiDUZgrLkEq/j3qIMkYqlfIDJ6ebSmLq6IPi/iXG+/YRB2dRZEqPN+ig1sXCQ+Rb
oci5Cm3QwgyTRxQux2oE1iQnHwNgCGM/+H4fUzK76xf3TuqS17saCNWjwvWgQI5Q
Z3p/5DqQSeer4El16E6wNnPECP1thM1TmzvLrosyedTdZcMhVrCHDNz3GZlG0VJQ
p5FOpS35B+/yCMD+7iQQ9iTRQfvzjIUWV98cK9gTrFEfPxjI8YPnBpx1VmzYv7m9
6gfeNQtJYIZ4353Ac7+CsHwIgHCS82NYfOi0fwN2zH5mWD23O+P9JhEqlGm9EEVS
IVxKhVH4dV3LGGiYlffJ3mmpubOOEuxAqDfBMsmAfzyueIpKxHGU2ktYBMzkWoVN
dP3GmVzwtluPAYzmnAzEHIIa1OJtEHLP5LE4PHwQsGpRDRj/8Csi5xqzVNc/W4iP
pO71UQB16cIpClBO4UxXsg6x8R/aZZjdBk+mtZUwplNGtapPMY/OFkXUZs0xO5EK
hssAboVlmxKa9RpnDsN0XcO06WQQlaQRSV7/9g8W04KzGjP088ptK9DeyjbUEkL2
CZ2pp1eUWExJk6wt0mt/Drk5dI9R0jPY5m1wu1yqm6hAYJOlsh6RIePBt8bFAavt
78Kha3QdFuml3Ng8j16W7n4j/aABaKmzGXsLXpkSVOnvjc4KVAtpvu/xg8+INIA8
wQDban4jUUKEshCEfO/8YuIT59ZR5chd2N2QWwwJyRsXnJSrLhZJt3LAD5bqo2MQ
zTgxM3IHCoT92gowCLUAOJgzQ30o60cS8eP2U9a3kWWJqp2enYoJ0otbfKW2lW6y
MyerV6RNufGroBZ/jvVYze5hcNR0ozNUYaLOvlNEQWi2awCMifS2DFdvDHH4j9ii
aPQCiphki7jNw+p0AxlX7HY8RcqmoA7Xq4o+4Zht3WLecnGn8Eyd100CH6COy2PT
ID3Bh/UudquU/jH5cbqHToEf8mXqsvd+XvoZIofu5SPoGj1e2BoSPUc6MzRG/eU9
itbyd/7qEaJCG5Nk+x87o06UrkfDt1xCyzYUHq9t7k48vkDd//cKtFNld4YAFewy
tGyWscfpVVDNi6O2LS6KMgfybnP5TMt29vpt23bqoc0NSW4uZ+d+Ff9JmC1cV1wO
Yc/VgoAneE/yQqmvFcD+GTLlCkwTTtJauKEfFKX31yqaP25TzlTTy6Xl16bW1ttV
eVkXv2K+JlJ8GSxwsqM+6uS0waR5HaUW4NEri5nIW43rbS425Cau1l2+ZrdvUc+S
grv/3wI/Gv4j5Azitr7ZPjFWCx9SW14pPvPIwnU/FasRGlPBJ9wPD5rjpsQt3m2D
T6gX/Kv7f4UrpaiqoGlhuQyZ1om8XSp5Q27QneGlj2aA9KEmqtOa0M9hbFnAhXnP
dcamm4s0e1RNCYw/5RebdMFGSyVxEB6JLpjITPUmI2SAg/3w8k+YpC5w4MpBQBu2
O3TTQCrXhxDaf6mKyO523Ro0+pKH+53sXS271JR5tg0VR6skvZEKbhOVfvYVPapl
AFlauFYUYQYI0y0FuYDbuI2Ruh4dLd+GgtSKapqUYZ94rqWG4LSQYWXbhSTElfAm
vAbRDNRoOcSu4/u+aT/d/savwBPHS97ph6AtHNCZ2nFJGHXvaz9DBErODTAozEbE
b/8BQ3n3+2MXx5vGBKS1q+LHDoz4+KlVYXV/2b9j9nmUo6DnLA0RzNF7z11jPUhb
gcd4VlkyPK0MkD7pDHkyFIV7Luv57sxNqApM1T9FGcn39wHrrCJAp6VJqEyBZb8o
JRPGSCeIoayksak1wgRuZ8jsPcaS+1pzShVQ4VNUKGSoD/plarACaf7+JxCC4fGY
ExzH9D4hxnQorPptOx2KKXyswGfPQjagpXxm3t6o7mURX9mSq1J+YHeRr3Y5kX5E
eHB1RV2RI4gn1PC+f8OmhwH5+0fY3AUu0rO0Xs7HAEXVxUpc5UsZXSh7GRZKBVgC
MJ0j/7syP9U6RflU+s7ONP47HIVrD3X3JdJ56BX0LPm0izcQasa0NRNCRK1nBVWO
vjc1mzWABPGWK41EYGY3ipuQ2qoZV1P5PMWqIuEAUyx5j4ugvtnz1EIQyEHNAChn
clNEhEeMTkO93JMEljPHycG0OScXSW1Ho/ActvX1+WzJIJFdlnAY2Y1E+VAAGSjG
4DDoXR9XOPHEBeXZgndOKH/FKLwc1JOD6mjxIWgThHNB4IHIhMBl+V8s+ttyWJMO
CxYLw/5f4zE50tDKdHhPVkjETb4b6zO0ixy4iaXXJDv85hyMbsqjPXaz+VVEW7+O
YHja3nYA2FtbE6f2rhtadepaEQSAgJWTE/yJunuNZi52pT8P8FCWCzOs+W8Zlca6
sSruPXS5ugLlTQ7VhXYKTuDTAf9uujVsnqtBFwR5eQNw7tt2r9OY/4DfU6bS1AAQ
+XXOQjV4yaqVkqi/mCasfJ+Y6eBp8eyBqdP2Enyrh5J9VFOPZAEUnsy2CuJ8rIJH
s++fEZa6cH/BVgKzbS6Vfg5lrGEEi1Kt6LV7H9o1+uiisFLtXYlGS1UZWcx5ZTqd
Wge6juAvXSyAqz4wHGxkbMPWDGrGq8rvRaqNKclEmUKvvC0vD7f5aSXpksGCi1NG
59pMGevkGcsG3Sg34CacjwSsQaXXwZHgfyZ+ReIocYhPmui8WWQDTqKY5c945RVo
QFCZ/+51lKPh5m9KJalAIS52F9SRGtPinpOr3MnoGEXWX3VYR9ggaErF2xbxL8lj
Ei7Z2fKlBKsYFtmZXwl7+/6HmSVr0kCZ31gZLxfWPha513UJxR1nOKgXcR+DQioY
HZiIKUFOzM9Hu6VyBb7nyD8aid7UsrWz+cwwbhEMmo0j0x3OpcXjQ95ZiUrEPLBo
0oBvdfFC2sjIYcxyn5aZ3KUv5e2JfA2QVV+DLN3yjA6DVZP0Ak9EAjsmmCkpcnOn
+snwmgZ+sGlfm3+4N5ufwY9jyEBDOAzE9Y78AsbdAUvc1BPaCw64JrYfhnpE6xYR
gS14bYLChK/VjsUIRDmBguA2VsxTlvdYUtmJSnM5ao0T9RLUNBZnQg6MEg+VBp0J
SUTCPAU8cxzMtX3eP38nY9+TpDVwhLNRDZIKnSdkOVnK+q3tAjZNjAo7RSdyLa2E
5losJ/DE4kF8JoRr64YtLds1FsWxg9DH7WEiCZm5R3aqDHMJj0cWUJbXpPYfsfuO
8RKzB2pvt+SFL+WUz8YaVGQf7p3mDVjOZwLdHehzxK3MPg/TsrDzTX4O4zHdA1+T
JvynZTj7nGrZA3OxDbDTtXb30CEHiMbgsc9VmDTd9edo0lgervjeYf0Kj+7mWBOU
zfS/F/GXmiH4BJapdQhvBdR4qgQnKWBuJmwDABX3gAVxkZzQFJ2EdpHPhzY5FXCV
MWiNNXfjYqM9aUEHhWDrdpVy/LmVI5EacrImg3veBWp6hADIOVVaFL0TPB+zhnw1
tGIrKIN6Mt+MJQeB/6CKahSI4HfmNDPigwn7UitxPFi8XAZvMvcrPKYdhR3Ulj5Y
9t5F4dlMESgkTr3ypjcy6TdX+AxcFdXhXa7Zr5IJuf5CWxtfqak1icyKYR1dbBAn
+OujleuSymax7POaIwRAdMJ6DtjeCf6hjTyKVPIkA/6MHLRpbDS4OzlPRRgM/SDu
AvvzL6YUV76Hl+Hs3p5rK8AopRC20UrBXO/8A98F0vcYFjWymA8eACworYnDQ1k7
Qo1GxishZrzOtWiMlJS5NaIGb3oFcP0OqP9BLP/Fc6n2UJNdJEEtNerraQm+GzqG
GHQ2DA95ErfpDtsBbnF+VkopUXg8unBH8v3rCqWS8MgaTZhEsT78t9OISMK7W4ip
Ueq7ABm5scmrPu0bZuD0yAmZOtpNKkyjnt5RYrVNKMQTquNiwtm8OTpHakrdyqsg
E6+KcLAXVS8wwCGedlj/7uDNi8K+OoVsW699DwJFbdWb2/p9rANqw5o2PNr7Xbqi
hR2zHhfn5AnWioAsy/TGo3eaLcQlQg9cr4IZnyDEY+S/GOc1u1If2Iea/h9f3daL
UDRp/V/yTzb9oS8ccA+8k+HtEh82HRMJti7tHPcI0TFMtEm/Rg0KIHyOpJMGMjPN
9pr55Zoehryu+LGbJYCMRdDlZXHDvNftFjlsjhEx7KQ1okwtXRi+7B3dslHw9V0N
Y1VL/AkQK3BSCUlN4SsBMRcI4DOj6IA5bLE9wk7r61ms0+jrgIlT7Aa8xAjEiji0
6zzEtD7POzFtIGtvdad57CpFl18RXflpLc9flm3S6fssodoFGVj/0S3mrHBublAe
c857CrfqQSrjeDR6gHgThP8ns5KRNeBTYZazpLKvfydW1guv/WRa62vLis0rntOc
JWpcZ5eSZVspqjzf7CBRtpE/ocznCFETQBlqi8i2SCfAYNuSyGRFp4Wb5J4jRjWu
xlmEDaUQIjEOCRNkw3A5fb0cbUF4cC5OqZnh42iappngoTzfAVNAHHbcZb8rp1fE
VT2KwZ3ntzcKmYnSLDuXGBiKHfOllsMOmPGR7UdH7FhgvQm/IkYYi4paACYXP6oP
lOiV7peYUiWBAvtyewC3UTroOeNbn2JMf0eaHwcU1wju2qD2dfexIOjwp6ic6+cK
0Qwiaoh5N5d+WPWI9EDEOj9SQfdXS4WH0prjjRVkWc1XhU2yYHYWRPWRW3J+AT+K
1KNFfxlGjIZbWF4Yi8j0V7oD+Sj81La6vviQJWtTm5UY6FVYbNsmkluYmqtRC/lD
rOWRFK9JKM3tLiUct422B2+QKDsmf+tmKj+EGbSQOhDl04zaUbDABuNFi5a+w9dp
0XrEGR2GodvSLsM6e+XhTEqW44UQNxaFCMNxSHp/YPl+1yUbDMzJwVJFc8iHuzuv
1IcqxS+qBnL1V5/svmO4kL4JCR3/FkXMQBKxQZ3tTQI2w5QjS3NWroO/fRuR/1C7
r4+aaUap8GW+hPjgnPrCZAnbwqhWqV55BXvU/y8VehUw3yxmuvW8FeXUWDbglvld
tIpseKVyJ9hytphQFL3tR/qjmYk9k6ByA7FJc4HsOcq+asBrbpIq3pFapg1M5MsD
6HIOIlUWoV/pU7ceX2xrkFWruiH8e4zc54eMit6XyDeehkqGSZKkypL0t/7D5+ZA
NUym1qZ3KO/a+9C4k3zosgbU4SwiOh+CbZ9A36sTMQ+Id5o/xkf0nSQFAewzgkch
pBj2vXy0WP2vHmTnwhv2d6Hr7mIqcGcc8C3vmUjD2EMzQSTjXGjUFMDV8165ovA3
Z6GIQ6SQ5AY3hDofMTdh9aSF3j1ISBgNHEVLDyRdCIxanaeynIOQegmbY6hKwBgw
d/ee1sO4vP5ZnvmQNb2cY5y7KcR7lHC9DTJUwpKlGKHBdmidCn/EHCTKxwHV3Myu
gA55rJGgeFXXLldV8xLwi3OCYM0v8pu0eD2LFl9hcCE+Msw/zVSVSKe7qUN6Vjyh
+rOuCYOFxqCQ8eeRmKgNSTSq6BknKo8yyGoQdh+seHakat4hvX6/nvvLZnT1dlTz
KI+QgvfHEkZS5RYRJpGRt1YWdGw49eKnllBCW3urPJTgSX3BcUX//T/jtVEt/Mpl
nrYJpllQ3eNN2k2mot0aQRvRyx5oYDcac1nJakn7IagynA4xEmzRLJG4A+wQvrK+
bBy62TQr0QVZGQsYlCfqPVp+z1d9JFPZAX8MuBXhoQmputSU0S1WY+SFhNdqN4Qn
W4RH8nouBWNVeni+/lvbWgtSCq2z3Kz6dzzKySzyhwK2qdtcyRlVSfv60v0e/lU9
kjV1kHOU2SPwrMojaLJAgriOnuH+lolysCiSzDrYfXLUVuC3LMrXEXJy5Bp3Zlcs
CpbmpDiFVnct8O6PkaZu/TRMXyncMb8A1muS/PN12Ggw3+xCEyRxLw4oaExU5uGc
zys6zUUpkVa/cNXCdimAWz+uroBhk/oVwb0py902jo+wHrZeW3bsi+G+ID9Q+je0
yuC2mFoDp399irBOGChCvXPjG+ZsobpF4RA9b7u61zTyffEkis/uO5V0xzeD9ipx
bnDR+NP+uALLl238lWuWqgqcafXjcFJJ+tGoVE0mKijvQmszpticR9EvdBTT4lqK
dPyPqMHhkm8IbT+U9eJxbflL9YUAefQMiOsnO1i3eaXFjJnxL0zJpY5QK/Lsc8EA
b4iZwMHJfNJXuq0+Ph4iIgyWuU7Aow2Sxho03DSpK9LmW4NQRJx1e+g2aI3U0D5m
BHioc3+SDp2G+pHnzZnjUYueSA/DFue2u4acJSqt0H/OlXmv0sYNbtBb611Or5xA
+BRXn5ux7S7ff75T+aNVwfNasszFVeSizGdfuIGvrUEA7PQpQlwAFo0bR90vVVeE
MGnhLnvqbwvZzr8aCnVUwMcxPbwPWqpWa0kByWAdl9MXiE2Sjw2coBSneYTePmqS
22AARe3O18dwyU5llvfxlwZwq0q07FXzKrG3mcl9Ep/WdwoylVnB7UnCASOkgm+a
+Mlm8hfmfERgF0WsAyQ1bLMvCr555j/g3MwK431faKy5dY4cNPhgd7v2JzsPRPxO
RPhCdKtye4zf7VD1FCFfCFGZCIkitOM6YgU6t/73tso3+eKYO2eW9vYgzc9n04ZH
8B/4YlC2B9kQ+11sDfq4UJnG9OgFU3AQfb+mj6chgw3WYDRAGoHNiEWgWzs+nb3D
wVYRj5eoO6DGswIHChgjKb75pHo/BmGcvZwWHIqlvQRKHNxGfJsud2oiVzwTxxEG
HPJiXBvjxQjFqJ7Pd/tQuQYXunHUOZMdhNylibcl8Y7IIT1R9VEfrzaY3h7eoo25
BHg/jrE5vIqtszJD8FJm28zhEWhN6BLBX+UaYotMdW1gA8aXPq9B4NXFaxVwr55b
zp14Frc9XZEXq73VzkgSjT9qVIu5xliOdH2NngFngNQk4ZXrOi1i5u8382sm0cio
aK5ti4Cf1n8xA/Z6it6SQSNFIg3QbrSs7owu9s0E0WFvVEDLun5r9zY7oksgr/qT
u7UGa7YgSNM52WtzqLp7kbv73ZQhJgj7VQsfmwF1RUxgo7PItARs0NYh6e6eHdHj
3cwric39rFhrGPacEI5/dLrNUCVKCWJ8OzkrfmgwUCN9OmJRDeLKj+LyRCtp3vWV
ZX74XLb/U7HlP25BlSXEjk9oI8mT7SGWd6NzqiZRh/UusBXMw2Fyfs60qvjXhePz
vDI12DhDZXeOJKUPErnXv1n3W2Xp53TbWqQF9eRNxe9VqO6LoobZrcq+G9FZzPDK
7iwPBOZl4gdDaIgUiWPrMfpCiM/vB6yi8F/iy6nVy1aHg0Y1JrAAYYDd4DYBdwEv
lrr6wDu8Or1XpQVcGbDNtWOIuYEFd0hO9KR3h3+JlXAexi04IDMPC+etjFzIjOOO
/N/kacNYfA2sdBi6WNyM5wZ8qCOFOJkXPLI4dd9hYw6d6lF+89HxczcuvWRkOjvd
tdv/DMwUlUZ8labDVC3d1SaWx7Z7eiiW6lswoUNMRdNMEiWg92U44z5U+1AkIkfv
6lhgPO2Ol05V/F0mmdE6wKMKzsBYN1bYOohNY9P4cwqd5TItQqpNb8tQzJz9XF22
gBCXlNK3S0msqNxYbUSZpGESXwg44VDQKvDfU9TebI54OTCxA8DQPtHV/4MMw66R
JfbNzIBuwb8J6/P4ogOKQZutzJtWeMRem0XXG+f5iY2EwUDHFAxIBD35vtcIRtKV
X6wyZCNL6wOOjQ//c4zv96izstV0l++7S4a03T8vQlnBgWgIWicXqLVkEQub9/Vo
Mc3V21LlZbJVro2PbKDSEFu2kmdQ334XNFirAppDO9M4T3hAH3YuUso/ChPVBe52
YIKm8NweI1f2ufzH+BhtGP8jijxSGiS40uRBoSqcrA/aBtqwEdoe/TWbQI30sJ+M
hgpZSufz81HJzTUoj+kCAfRnR0fugVk0zEUJLVmuXUO5QJ9LJIVUZ9k3FwDT4EvY
aMd+4VKF8ZnJXyJsITUs739eZFWepABrWFSGU5cPAj4RUlB5UROKdI3GqldqTEjN
L/mlIZ2YSSzTqXyDFiPipcW1f7jtPySa5ibm6LuJ/T8Js8eq2GNSvi9KL3ObtQyH
dgUFRIstZHx+XE05Abp1TrbZbNUmlnnZOj3tEyEOJX0XKz4doAxUxypry0ZcYf/D
eii9T7iqzSmG8MXWsUd8XhGwKf4ZUeur4YeCS2rcXkJjNX95Yk3u1choGfwg3FxX
If8YprzgJjFVZJgj2a9R0S0R6LW7JBcnG1ATEKUssG7lzS1WVfu8e5bpoRIIai+c
VZLQz15IMlrZS+zsiexGPUV32+3n718cvK36AEpalZ1S24MYyCsVHn7r7NG7N/Oa
WVNCFuP4mx+tVPsdjXIZiXScLw55t1AvVNK4GNRuHo3tNsuD1hsbl1S18yx4+VAM
SR41aoQTJg3wiKo4LAjHDKTZEQ+O51YlVauNl4Zx8CRa2q8j+UgAZrxaOYPMStQB
sM35vKO7XKvB3ev0PoaQqE6gZE26gyYv+BFmytoUN2st1iuxC8izydyeddHOvlaE
6FKe+vncKECV/tefLqJ2jjzKISyUEWOEj5HR3U5+dNVxcoTrxbUlL1IBGTLwsBE7
Tybc8kQbKsx/8KdnoHGQClglVF51eVPU0nYmwvKeZdlNAsJ4luE+9OvQmsf6vmbv
SFIZt0u8NPO+c+3IrmSCfKVz/SYe5MmDHSAxW+vPexQJnKUiLfCCU5MvXYvbYc27
IYFYAiGWsXVRlsBqn4/NONyV+RFIf2lo87/7/eq5COolQfWzyxvveIR/jcObYbzd
bT9ThEG0ehbC8rsyLLGYpCCwkL4p1yB7I8Sm87iYoyQxEkl6HJgDR4Z+573EqRJI
qTnHU6NXygLzggHBNocfE69E5lq795NePCxECGKdwnlc/uUp7mCFvPCWrrNGX3KM
q3R13diXpZ3IRUEpJDvDfDBMK4FY8SkaYrxP7y5SGxZLgAfXOv/0f5yQq6G5J+Yz
pna5+VH2DYGOt4Emb0SkfATIzEjvOtb0xlgKpE8NeIEgrH9U9baNawn+xb8HE2LH
D/v5f2a32rs9ehE1LDoqzR+wHQ1op/WwCT28xGzXZD+xfTfL9lPCmh2lzJe4AMSf
6SjBwsq3r6EEw6A2Fl8nCpttO6EjToyNWuGSb0vuJWjqsD6kmzVurYNn1SAHmOLY
UIIm6WIKSw9tdcHlHaqSNkV0jxSUV8b3Hsulm2GEOcCZMS2Jottc7PAWFlH3U60R
RtUqvkSDRwa/7r205zFXua+4IswBCtxH0v0tUCQsU2CyZ+HHZ4BuGbSFBe99RpUk
PeNJukb5+zu8xOqYMiqZTu17fMPEy8PB9R9v0sShKcQ86dnsAETePfUkT/AGfh+G
mmrJCp2V5GbqT/lfOEfDa9q0l5caIMAihgBPG+42Ees1sMrXov+Pcxvx9XRTctcf
TPzQWNrQ8KjuB1Ce/JHZqMncN5/s/I0X1UkeIX8Jt+JWKwrUxFhJT8aIWAmX7s+w
QYzWwrvRP2YPhOKuyspEbb0+mEZzVhl4yIl5+x4ILU7C0iuha4Hh5qpawafO5Y9L
A+dMI1NGFOtumVuUKQZhR1le3/csTFtwu/F2X0n7q84ZWyKBc3Z6Ai3UdbY/pSbr
9zc2DB9b3v9Eo03ilpE0su5Fm8at3TDmsre7RVPHk/XTyN9iHF3TJkuYrCv91kw5
tvKE5E2mbhc+mVMyaRHdJpNNtc3JWsK3wUvUZYITxGRkvT11dz4auamglRkS+nq2
hIZwj7JlzVVjRT46Vs96BQ8R+9V0fuofV66oWE1+z1VQJOOZ4PvqawEaRwJITTXG
TTV2Kd4YGuX8CAZ3jpiPmSlC8DmGf7TYABRBMpE0MY6FawijIMk4DOhi/hzAZL2X
Oz2ryenyf3kaPQ+hLr0JXlt7rxjml0f7tKjOf++CHd3FO0krbjh8MpsFCNofLU79
EEq+hqnG25l272unZS0VaY1kGMdD6v7HnbnVPNnTG0mc+FEOtOo0WmA5ZtxDMeeU
OHt99Cb5kIlOS4hAvt+NNc5LmODO88Ql07D331n7XSmZk1s9ZVIo4Bv/apEso6V5
69Z9tEgmwKyA5OJ3XJ2uqc+mbKQjOlhvT3j5TE/umU2If+jkhmWpsSmJz4qYfURY
KtbeSA3RNpxUXeYGT6sP9hFkHArSZy2bSXC2VxeV1JGwZir8M7GRsl9nhFa79yUL
Iu30XqB/0EoVi75a+vnnU81oKDRRZWdqd+dwTOXmxGDE+CU9Z//bQzN7tkOC21c2
MvokbWXkXWfrW6a84E4Yr89KLBfGLuyGQ28YlsAxDEt2ofKWuXys9VV1VznfmU3d
zXIlGVZJw/B5c/2zmOVX8uXpwL+WmzCJ9VHUtSp0tmDNEYGEffthJrg8Wrw1BQVE
bT15bMPk09H7qvNtLsJyM7BdQWS3QOReC+6b2rIHwNCgJDxjj72x2+hvbwXkyffx
NJfIO9DZXzf4N2ds9uoczlXTEEjlj7ixcMYyV1RljnA7Qg4vYteMfW5+0hexoN22
kVjD2Lt4eQlBPgNOeX1BTDhYBRulDxAA6MD1Vhg+HIV/rZmcalSAYvSfaLZqUj6I
boncodqp3lgQZEGn1t8ukrXByFV/OU8dTtAuz8wWiDbAnLuNnCzNodkkqEObaM+6
ttm1/fQlSxd1moOJ5Crl9iYVV3saH0xQ1ENXAphHsIkzDzSx3FLA4yjLxGXMoDGl
YTxxqFzqRK+xsxmRIgypcrNBsOclG95DpK77VV8YTiBrlcprBHkbG2DNsebmdENS
uvwqryihZyTy/YT+1VnnmZR/+LY7gmYFOQByUkdgBt/kilsiG+wC808hVjNhwYYp
FYNwrtlxMdOhQqfXVf6PFvIwnsyb23N+umf7TUMrYL43ijLPcuuMQKIfjNjGhsii
r+43Q4PudDAiFm1PXuL/WDKmfShidFj4p7WhDb3YrRrOH+kuoyMRdtEvaYEyD+vW
x21q7d5wFJJ0fomi/YiEnlVCdX4jXwq8SzGKZ5ehTVdre8UxSB6Y8/LSwKEpoG0B
BDnu8klxuZdXEGgPIWTHiiVMM/etv1GfCp+xKFqljRypQXWDr69yyL362443lTcN
QDh/xwSSUAIQePqAiaqzSHXswUaUAxgmB9VeBKb8K+fv3x5C8qXUEmeZszJVCy0s
lqWz9cjGINJxhK+Bsnb7KVysz6Me+1AjJ9qv1wMZ5sPDr4WpVcFBBemDNFzCJNgy
yU4gtWGWxscA8ZYWEaRBUAn7p1cxaNHjxOkLWR+LOH735YocW9H0KPb5nlvonIDS
oZdr8/sX6nRd6I9P3ZDo62+wVO1oq6Jr2LzEAaKh+Zc+EQvH3Bik9GZSI+ZTAusa
WkGxQbOJnIViRD79WmZMQ6jxKmU9NlxM2PK6npD+UgZABGp5o3W9II8+C6WU8eiw
r725pfFtSjMOswrnNWX80N6oYrdM7c1/Ez99gwy6JpX//Pwo97idJrbUJE8bmC6V
IZEDb5kBmpJxoX5L0b+n2+YrATPm7kU/OVT+MmXSoZ9MT38ez9/lmVN1bTYHgbGh
PUm9tp0KrPaxhHUDLxpphXqGi46fMZDx5En3RI3XrsveshfRnJD3q/gyOYEmBTyM
j1Ilv/Y3uZIOCje31Vas2P+w8DXcxXwTLXtMFTYiD2+e0GSH1cCmFLICig4j/IQ3
IFz+3ZyW8YD0yenvJzKofG80K++hgW5dlPntpfcZRU5aUSHjvr+JHFY+yPF3FsIT
InctGEWBtKb/iv1vVz62ksVKkQhuqFXzVsO7/yqL26N3V9DZ11gfeRwb3NQF3Yps
Nb9WcUXwVrx9amyiW1YqWMxvYF8IoCucI/Eo06rpccGx9zR/toZfQvD3u0pmlMwD
/cOo3Z+Zk4m0rQpkyUZ+LrwhCeBIJboK3Q3yQeUlpcinVT4Xm5HqihyRMnh54fmQ
9ovinSX+SGRkncligRsKHsZDKqzs8JKA4k1Wm8e7EFJkvXgCP0sJuN8rWXETKWOf
y/9SBmapsMBooF/tSk08kIgaoZTQxtkVId4FHRgb5A5FPsIwB+fjGg5IalXuB08T
nXgCm4vslxoDxI6TY2cz52Qnf6P/J07AxeKuWO+NUQ1VmU0wj4Lczsh/gNDG2rJw
sB59ERfeu9afs3qT7ZrlckLE4aqmdUZiaxB4mfYblFhyIGML9zgAAj4iFpYXM/mV
QNdg/MRHTW25lqIJqC5DxqiBlir4/uYPdcT31qeXvih086m4/thVEBGfZ5qbmj0V
bZNZatxlt3Kf095wXaHSVE2yE16gjNalyhRZWMr8ig2c7rD8HNzKL0XUEtRd+BJ/
OPYx6b/i35O0ox3nfKqgrf0ZND2v/TEE9u3A4HYfh1FI0VdMrlKC7Ujeh7gW00Yo
vUuwoDJ4CdCoWG0GselSax5l3DoQuVvko31Dc2rCS4bVjYcrG8Z3x7+yFiebzGCP
3eyCGXWrso/EAv0Sw4Armvje5/H4cNQRonOcCif55kBFD3nfUkAkxZ34gKssHcMy
emj/x7SfFeZw0lQVJJbdVF4i5bhjebQ0vSVlIk8s5fZbPQw5nTwIk1qrGmR+Nw5C
aAt84mXJ7jXY0pCLdjzc+faJMx0s2+WfUZKGM3wLdHMMnJEEm3cyRw3CC/3DHBWp
fooxPc5K3CbpTMxzS5G1sVzytJjBF8+ANncTPbEmZnugLHNpu3wJ0GWlQOMhHGQM
MVrQvpWytje2rsz9fiVVBNsfriMLKSwGOtiN0z/2u3wrwyRPLfcmZDnt8EOA03Qg
RnnQvmqQbORmIN6H6oxI/5UZ7GgAxFcN343w6AkIM2Mb+47QZ1svNLBKH80LMArX
guXpcRUlYeTeiKnJ6eQ6vegEE3tJQFrjGzyMIKyokTSDPYO7bwz9jcIeqGWmPpAc
IKyWYS++9Zscg1WypOep4Ofj6yxeMdPqdT8hvdOIsAoEbwMnu5LfV2jHYthbLrsr
W87JWBlHdjpqTOgjptxuwvyJg7zBBygu/KUFrz14iakxrZ0XKPHPkHBvzlktvVKM
f6cNYoAqR6omtuu6g8swUUWE1wjn+aFHpyB42f3U+hnDDftvVYHeS8b0lER2fWnK
mHiRwnM4ObmQE976kgeFt2d0DmTlTjCAU/AP5IfaY/pSfwk/Qbb+eJ/NfucbFzdO
zGXnNqbrLBTju2S11LTmIvhmflGI68gx7Axr4RlwwYd4eAilB2VdXEpcavMxDdBE
o2lT6sW86YMLqEYp9ONtx456QwbJs2zxsXHCfh/NfsfiQc3wG0jMyoXUDA1r6C+v
O6Cdw21mxOIL7tIpgsXEpq+6LBUgUlPtNhHMxdhuV0BnfJGcAqgiOd8+UArUPbqy
edXhdWD3A/NyC7I6Q11uf+yFuxu+qXyur9I4xpxufWHdMnuaGNxdGi+KqCXp6qEx
k/NPsBNDkYD8T6naUWwKYuJnyVNHcCaQhkBYSoZNeqXk2Q8AbSyF4XeVsEavpvVV
NsyCnbNQ7VhgCTiNg668KYg0gmmFhAIFh4WGF9X4NnwkeQ76KW572/6loBSID8Xv
Gz4xy9sxA6clkXSy9l+OTSF5QGigfWui/+cER2Ckw6od6gDkF6/d8K81i1mVqvxh
yjmjtB6Ih6RAw40GcecJd3Zmruf5u30cOYT7x2l00mxXymsSncqlAOLPpTln+qWL
eQqgok4DfljxJw5LL33527iQyqrb1tNamaDv/A+vDsvcd9EPoXCIXSUwBsCbfCLG
9e2oNXpazQFIQab8i7AN2PEX17kAR/6VO58ajEKUCtdF3jQlYYphjJBo5FKjX2Yn
UHEqb4dD4iJ++7pJHgPdfrXq6q2CwAfHZ9CsRPQP+UcQI44kDmZ1L3DS21e1dv/B
2eBEzHRY2Z+UMQVNIX+Ri6seGYmfqqf0uViQ/l2Oa9NgJwDJCS8b6Ll6RvrSQwTH
1HGRNLK46GSNmjuL3W0r7+7qRivpFRAF1DsOf5UlTboI68Xt2aDfRBeHxXSW+1zA
5ZIqTg3oHzSUKbNVSnRlCnXJ1TVkNXVqgiusvQIs7vf/xorPDLTqzn7g6TG/VKwe
dOfNZwL1htnsSw16+llOnGBuQowNbzI0xBmqG1N45nBqz9uj/kyMrMnK4758Ya3h
SIynoPF0ZZLCs30Izgc9yXbjh18a5d59uB3aof4CDZGQJoclXPiqHsUEy6WrR9DI
2XLOkBhukbo3GfWEwcLJjrYoQw9Zth6zrFVprEjhWj2r05lXedlwwrcZTFFzgGmm
i+6HasU9ZrNCgx7txwrLfJTnZN+wFnDyTUW5ZwTg8mTBfYcLE4KiYjvTUrjaui1m
ot3op+4evdltcK2QP74j6exGM92Qehhk9YV7xLmFPFxlSxqz0AXHT4Y/ZxcI94fx
Ix6b6gNH2+qSvPPeVKojdKQ0C1pFPzhvUmtJZYo1Tt/gtxfe7Ktm2L0c00brZJuj
cBwH/vSIa1ADHqOJ87CaA4EwBbznxWEYgC/t4zkSHJWN47bxVyzurUp60r/IAkfl
flLHZS1dLd2IldoUTxKMxqxTHP51BbxgUr/XsZiQYuzgP3GmN0NUow7uGIcN1+JR
HeNhHqoI5wue5QvH55jzlHD5QlL7FDO7XHcixFzv3g/w5H2OPg5PrfDRuclz01CM
qVuQW6NRqcdM/OJTxt6fg7zg8JJwjinbMKMXPUtYnLkrni/rM0AsQYYzx76o00LE
pN+/weAnnBjlJxcx5b6UeWGL1LdjNN6qy50xf6Mb/Ow+r0l0gvKuxBImXne8LMTs
JWvkYdPVAb2DkD0unwk0EdJDI943BZmzGywRyhbNT8GOjiT6doPjeXVSJo4+qeKs
0+Aw+caipIaZxTpvJAugvnoIqeWMkjb6b70Un6D6iM7yGc3jl09DOEoTbkkA5pzf
mFXhyX5hmbpsv77lUen3B5X942iBjQN4pOBYPG38sZrGg4hpcp3SLMuj30XHwtu7
CLA8rqmg3gg/3nLIgfIbhIkqc+EqCU/jCjS+4aI4lItl8HIJ4YExs7h3FtVmkCXG
rMXcETz6IsoLTPI99zystcal7ocfEMBR04t728t4YEKJi8ZAgh88VBHXhL3YGN8v
S9jy7QnvG9ssJlNf8MnoN733k0HOSeE1HvE05IARO6VRAFxt+FP+S/ynioGOYqgR
Ki6Dz9RbSjkDaLjNJRP8hOlVKazga2eSC9DJLY0D6OYeXoU3Rn45vgmB5hEfdFUk
7WSylpdVyq6aHsm1OyK/+ThJ/1fbPU5wjNG4CQfPHSoWafb1u7xEXSHDG2oYhZzW
kBefnsNXrX/bCCrDwSNUD24M7kum2ELey6df+t69SPwd+7tksqtWGcd9XVzdVQ9p
6uafRsz9Re4vQMVDRL5SBjOfY0Mw+sv8mYb+AZSm7QOrid3Mng4qV/MJtk1IxoW5
6Nqy/+OnTr4/Z+M0UWrDCcNA23MQ0JP6ntcO5k6fmpF7Ss8vsxIXl7z+L5udAtCg
YgFUcueBK7Ba9rx/UbxUeLlPg9+zIiTpFLi1/4tmFMLVfNwBIwTjhNef+/kLTQgE
wGiuoSDVK586FiQ/xhePoVzqWG8kmbtJHmKhN6Ln4z5dO6AvDT0fm57g9N0BfrfX
YCq+1UZmzCn2jcnqhnJuTTVgHIjdQNwDhjALu0BYA0ublyHMO1KV1d4KuclSMQSE
ZBZ/6aHQLDnthXFtyiLNWwrQqQDhEG9INEa8CIeuUGtqzM2dtWcDFKY8aVoC+JXx
ntPnTG1+4IIGy7TJ/baWxwuOHS7bDgLpGcU7A7gLszniu1JSwPIe8khP7Flfl0GV
p309GmyMuvHU97lh6sF4bRkpY6/aPsadU57AFiqt8LJsKCEoo2Tv0McGtdlfq3fi
d9iVWiEqQ1CoaLzgf79VDFtR3UVu81Oy1o5znSjKmHW6pZ7BZx1ChZDGR/k+gjX5
phTUR+YjHojLvEskhNNh+fzOTej9ZhLdXI9LHelAbhsVTHTBd8MK+vTB0Jphk6kE
d8OimCH00jSSvzNamXWzuFpAALzgA+eN8m25zP9kGrssslCcB+nn3Re2OElO72BL
o+1GcEbymVRxrRBE1gTBLojB3arCrS4ZyYbr0d6D3Ao+8RCooGpl2/JpOVLQk25C
UxCtvlCqiDaXB62iLeLzw4irJHE5w1JMii4jE8ofSyBcbXPmUDITR2eCT/3LQOvv
Np8df5WqnE9HbLSpgRf6BBre2ITi8atyMcKc+cbS1eyZDSQvjHPhZkQwpyJKO1UC
/+dvmtd0rJpOJodDtukTI0QcoqyzzFe77e2P743Gy5B/OW4zz9aMEQwAo1bishv1
lP8OikHHYh4rUyxPf5oLaoY8/IUw3skXD8bM/jwAG4VgiBTxnU+JgMBfjWN0HB0/
0jy4amYH+JhqO0U0aj8MioMx/zPlzyNz0AzA3tKn29StVvnZBGQpQF92AYZicaDH
7EOXWIaNitRSx9x8UdHUxWO57vieXtHzJWdWK6OiNc4Sm/hbZsJIK+1auyeY74+P
6I+QqOsuzARuAlFqAsBjdX9/5u4hh6cU/lRhfCUsLmoD+Chp+Z4DfrYTC7vpCEDp
BSYTBTK2PUTjDc8OTdFdFbvh01YewYuBdLK3jsCwKbibzWd1ewmRD5q4uudPy/5g
H3fxaL+yMOREyVpy8YcVuFBDhCeTYFrKTbcdXSGWVm920EM6iXE8V7AaAC4XVXJ5
hHqB4TpQd4i/hI4foXM3lZRvXPxBzTZylYKHSa0n7CPEvuF6ekNJSkRKrIsT0r1R
Liz+XUIPG1qHnukUEYUH1m/Trp7nEO7M+A425osu5Tzli7HdKvNV4XV9D+THvVUa
jB+LG/adRF7fGXMut5KtqSGagEAqbNYkPxUcB6wRxdY2wlls/GGJamL0jss4uump
WCfF4Zou2fZ322jEXTnPK3YmNW4V9ubLht/dBH0Syokoey6LM32XhOkCYMPjMy00
VwLcBlXMQ560VZYAUwgHL8nkE18FNB4R8utjRySreUyedmYi7XXzmPFzMyT0Z1BG
W7AFn3qj7D3PJ9g1XgHRyj1LyJ98/S/g3Gi5ZIMUmYzZFBUluMrD56U9UDN6jBUi
sOMkx+bkJF70eVE6/NWFLeQm9NRRYJXPVzaCjLfnNY3LQOhDkWeKDpIqEIyA62et
a+JietmqWCgn7KT/5VbnvhdsDX9ZAYaeillC8BeGzw6pOgbxZ6gHIALEm4K/Ejry
AljIBQe4XSebgs2Z8d495ovrf4Zqoj4lObnxWEg+mhWDoduY6Jax+/gMHh0/ws0y
RGPEFyqvVgDn5WaMl5y6bZkCeVDYVFSVmU2gnuA7Z5NBU6wbNqdPMqX2mgCRW6t3
UZcNWx2Lz09ci+s/l3UuSJ31+5YkIIY8NdVyJns8+nZdSINRYIV740MGHSOPZt3y
YRI4umAB2zqH1te1a71oUCiocf0b4bFWZIv+s6ecyVz+rG8Ll3ZclChFMpaiOQM7
q5NRXvvHFktL1tKx+SV63v0dC3Ve6YFgBP+3VRWvDykWPelLxB6Q07ZZ0HsjkAAo
lxtyEi1usPmFXfysME9byKXTyhcQo6MbuGztCVJGKdWgZfFC+FQqz4tZJrSVqJDp
vkFX+bOuyF+8dRbysi6OzesKmJa0ZAXUlz+fEpyvX2ZfSwwYP0PeTmqROcWjg+99
nXtEgSz43egr2IHXJuok3i8ghbrnrOsKModTdr60p5KKj8CllbapOuEgS/LXrjI2
Em0cjHPYjfc6Fvvv6ncIkJfN3PeUtj2+LYybUfH+NZa0aAF/qGe7vsaOXQ8NoyPX
kXWLkIpvjBBacZeILYAPUmg8yhOkp/hI3ZI2GioTDo8aqpYeIuuY2usNFgWd2Wbx
HJ0cWyRsNfaEptS3C6a38Mhw1G9TTfZLStxukuzAXwcYzb/OcAcJbBTZ9xIQKRan
nSQyD1QV1fKzYMPxYBS6WnszuFq6Xd3cL8ofOdh/C/2qo4O7UFZ9AzxncFZoiSVB
Sp/gmyQYYgm2QqRIp8XfW6tQYlLc1vXxt7/twF+mouzf/pqFOm5QMGrkhQUD7DPM
Z+HhZlV86gqrOnPNzbB16EMmdUuS3ABCTIONA7rJvTm+sInDF7xRRDchkQdy16rn
DJGQSG8Kv1vyIyMIve88w0XZC3AksRbs7xjANEZZAOed6Tfmhu0l5/hQyU/ggj35
YFgcTE7c/MIuiE0CMzsHDvCHqMmWaNeFPKlYMUQImwcdeouKI0LBZmlcjYES941s
jmqejWvuLBVSmHGcaCqsGWQsBRFw5DEYFrDpWwJS2u3MP3GbhlfxfjbiBpFhouzs
7o9rem5lFHs/UTnirUDFsMKvJD1VbstrEZnvaxIEyjaQQmIPVkACxIY0MyZvShE1
pw1rKdjRxMA+nNo6ED0xXjhwrDJ7SCS0YFTFJ2DUr5ybG7bZEp1h9paY8UzheoM9
CZV0eyzrQw+NsWA6HUIOrgL7eLR1oZHMfwFTvwaEkvtTIX6dAqRDPDD4QWFf3aEZ
TRNEnoZGtEh9gqtLdVI+f5/lC1ZliNcW6XAZHUD25hxz0LEj2vFleldLrBNyGwjt
r87KqBLfFzFizKCvL7BNQ+gwCJxtz8pl/vl1/4rq15BkthAqr0HHbeLton38Mq6c
BzhRBXKYIdRUgjRJCAYeWF0nlgqwuYwoNqa2fuI/UOfBwwGISNb7kV63v9/7HtMm
IsJ6T1Krs+kTUqzto5LKEGQfUv7GXlLbXyDf0h+mo371sl/OPfl4jfAIo/I5RGGU
n9zr+ZStGmzhQiVApyIeELy72dJVZkK0G09Q83XRDV4w4yZcm7jun2hyQxVY7Q66
OJM4VioXqTYAzinQx/9q7jHRqYcldwu9BzdTObUQsjErDidVZEAra8Qghjzefwx5
gjQRQh9vBcAo7dW59usXtOdvZahaMFduZV76RB6chcRnDSOtGxImoEgYaF5n5ouZ
Fa5OazOiNbyNxdnGCvrcqwV8f587zhldBLYKGeiNveKuPzW0pQ4ClLX2kfocB5c6
UTv+NepkADUNobxcrWi8wTe+3vlNbpIPIjmxDcGSVTa0cPXCQl1GIyI46YB6d+yi
apA0Ml99uVHbgo4vQlnoJqqSSrrOZnu14Yo20rmjePeyCgfl0Q3ofNJh2newDflI
hzcD9/sZVMCgjMnddMx3Zwj2S9HWXpEofV+DvtXFQfCvH4HEFcD03KNdr5wXXV9H
mvd6tg0fhSg8QUguHVywNBDwQImxI8ZIRPjLTqpviipzDEzRSOIlEDwVRJP+CXuL
1TQxB9VvnpfurYcFXtW4/ykof9pEUVcB5uA00cTjHOTyb/3Y7Ptwu1lh7dm7RafZ
xlCwDvWeCsXWEyG8+mwEHEP/F75BG12Eschdkh2aWS8tS/ZW9GhH9EdJIZ8Kvhey
jzsxffMd/OzgcVyllyrEMKa1xu2rjGDlD5jzkTtxIKhZ/6iP0zRlrai4WUOf/0/X
xW1excECwNn2rwnIixODEPSCdLBpvGBf4WHCiQSf6Kb9bBoXduyWc2i/6qsrLgQp
Dr/vJ4pL4wmAOOPW/9lKwrXfWJLFF7ozFw7yDCSjESEqxQ4vQsuRUAJi/myKaOne
bFW17uW6u4h86XBF+GOxaZpXpdfNmlyonFK6WL4MUFSq92k/2W8TFu1fMNjuHRp1
lofdCnbIbtVmqE42HPBkTF/KCuJrDZ5Eq6eG5jZQHgMPN9wY7nYZkWMHdg7g3/HE
CY+5j0pOpG3blurrfR+ncQFAQC+ynGMx1jmDenxFnfot09HrhzhjKlZRmTPnszFh
LG6pCSDt2r2m10cRe6KbdLLhn5h/fKMjU9ZE9jHQOGVU7lTf7fzMSv50Tow0HXpL
LqGzzGnLl68ld6IOk0ohmn04hkOT/J7UGbwuBYmrWx5t9CLwUBWghFRSHublCIBo
CbGDfsUbVRdT4iNx7MDWmV30AAb41Ck3BKnH2+pFfR9AXYH2m0ExHgU1Xmx2AdvE
sIMFh+DMTbVs9CcJ1YRu6yMYXc5EXeyit2E6FA3r3Q/pMabQCzLSaUe801Gh+00k
1Fiy9mXw+kBlXPxFcgkb3HAdf++KCGiXFxq96BZ9xrptTAsp8pMmKTjvbqvM7Tnw
/y6R4n1U9tAK9bzMLAHBPQad6fUyXmkDZEp1QdlKzz3oQp7/L/HWLz5NLrNcgE1E
RRPnHFnrx69z7SEi8dzysRD756kyxNkp3P+t/OBm1lQPEb+BzDO1iZTiUkXNbC8m
ilIO2v8E2Z6hj9G97qzby/ylpbUO4HUpMwJqgBFAAibE1P1QuFd7sbDwcKDZqcgT
RlitrwbxdxQjBbh8w8GAPjsvdnu9n6zkOs/0lPbn4MWf8gCsSWT+havhVpclgTpz
x7wsxIUyYHr69lfkVAOPFiaXRRVO2u7Anecn86ljzeZoZidpMxKh8vyGakGhmaGI
vJW15vs2ERFBqZVOY37qqThnTizyWq0OIFnzDOWn8LPhOjgBNJ2GGph4hoP1Z9wy
yDnDdMs3vLpvU1r6T64sX2Qm2lOCYdfvQEdhoQdNQCT6dmFhGoxo6RkwCh+oPXFv
oEr3gP+TepcRYjEuPTHJ4wg/Qo4CsbanTMFxeizWywyGD1VwJrHd6KnW7J1TM53C
rQGy/hlyvDcNTmVQNSYZN0qF+rJROVBFc+44lYa9mBvk8Hgc94CFjxLkUfmvy5HJ
2Q2YLYurzQR//EmdizeHc35djE/Z2amcG495050HGL3s8bfAwR/G5gA3xhgsW2xz
OvTruSC4xTQBEsWppPXYyETMQ7ut3cdYaNcYO2wyj6eD23lS1yXn/qmwdI1HGjEu
0Y3iNyv1g6Yv9LuuGITrCqtB4gWLLyxOw9fVRoNMp30QkbDFAwpUb1ahnzq16Eou
jfMm1gDmPMMDhxZQ5jtLMnoiVCTrzI2Ug5VcCoeBThrMV1fP2PZ1IMdNcAW2deeA
dK6fCA8dJXOA8o0S9hXtdls6ut/2hsYFR8WjQIsF5PEeU/0baFjvPL018sqjnAeh
bldJR6M7p1FrMokGJv1yygKvlCQVpXKNrARs95pulxSQsZoHYzsvLQxcWj3joDtU
zDa8gof3tdBlWguJ57Uj//ctlfBlusO/OZU3i7oOSlu6UvqZDRUsnYv8ywypajQ7
8mBrAZA0mCNa4f+sjWwyeYKL4KkGQnyK0ayxrIeARA+eMF8b70OcE2gDhZM/Uy1D
psl0HsmyJfAGIMQcEHGwgsce6yjnC9KrovKnt3YogWCpjmcLMq+vEQKaUh9wPSzt
MYmwurRdGykqoATaGkfaQ3iC3uf5MkAnOOxr1fhtQRDqPVi9W9znXmPZLcKGgX9s
lnKCvif16p8hVefu+PMJRcMeiaExSGO019++WNFb6JKhuNahsHSJt2FyRFb8u5IC
owLzfBT+JFEPjw2oU4JAm66ZXEHRkQFjhWy3NMK4WiRlPKmITXOQiAb8Hm7/Dcec
Cy7eX2L8jrVPmJI20Y48mT1FT+t9Dfi6KGDeCbi/S7cJsz9NXRyntf5SUT5wkOE3
yyMPBiyerAfo25pIE5yZ/MgQtykBB3KtsxbOIU1Y70s2iB9HCQmu6Jhj31543kwS
pb4QJf868Mra7/r0Ko+7mVilqeqN78VNclgYs5iDbW3k7m3jGpEEVi5RU4ky8x+P
0m/4vdsm8zCrE0z8Pm77j5oD8kxSeEkpBK/AOI0zQXQNaXbmysF5DKWq7OvY2wiD
/dPkB1Wi+N7ilZB0jqEfqcfPXBHGsqb3+2q9/LtB9OrnzCNpLOwFMevayr7PB9tb
VRrBM2ktBNLkVL0bhjsonQSAjgGlOtascte8Ntu4StzEtrq8X1j9nElxQMBiTGZi
rikfDYOf6zYmf3ouEfj5rSgv0brtXo3Pbsx2gJ1DirVHTFAerjee8zU821ynJmeJ
M9ip7fDHNqa+ErTxAmyf7xulEYv1ds8tlwqm2w0iZpM4aZmeUamel74q0ClGkC4C
ErlLri5XLlEdnI4lnB6I/TJ2VcnYqLeCbwhIUWG0gt+yf5LGSteGZjNWoQK+XoUg
NLpSwKW7pRXQ1tQUmMF9nAbJBbyZGFSVoLUi1C9PmKIppSuOATgZZo+hPwCKIeJO
JOjXhxE/X1fDXsyqxUke3ciDALZsgjw7YMhzcGVfpGzYbtfmdL7B5TaH2dDrtDZ6
Exs8ofbNtzi2QpItvE70h9pv9b55EsFHiL4n+gT20JpJsukJxcoajvqXga3TQB/o
o6nVeIf2gM4nyUK3Wkl3HPcbuuJI+GIt9psejzJrx1LxLW/WjkP31cDOO4ouivYC
HeJfADg52U11NU64NkxsoesFaEY99N48CvAUoZd6319t2y3ccCic8GcmaNinPW2O
U66xc7QSocAaCaB9zY6HIouFF23C9mO4hgN1LNGoW7XdXX1O4ssQjRRaBTGP0gA/
X2GZnOf3a5TKHO9CoH5+VpIX7L+AShffFpKE3Wz5ymgyMx2jcbEUBubEqzLwcV/i
/gDmYp5IazDeuAMaxldd1NWzerkxX7I8AYhX/HyXiOb1AOxNVCQsTGqbayArHVxB
QUvf1LTJ6LWSNS8ViGZocnFuxVJKPKWRnu1jPyQ92X9hmUmRpTANK8/6tuSIBrwR
FtIivRIyvZ//+0jAssEIhraqsp8W6LEwnxEzaivhJjWB3eW/8cZt8jN3BmDnX/4f
2B+9VTkZK/17nXaSfEqc1I+GWQ1l5cLpZjaWq0iywFxSDE9DfKzu3UsftMd1iR/j
VKJB/jLxiJZkzdgDR4PBK5qfyYYx5s0kvhY2YtTY56D9h80InCm/bQS4xD5GZEBj
xjqdLQPE/CbjrJye6nemDldT7B/cl9SxEm3oxYnXlgzWUz5ayzLmx94cN38imzNi
/8r2tOO5apS3fwhYE1a2n6MbxHyGtpx339bIg+XEtFAUgf8jdykqYbqNd/YeqjU8
5kJqR9/dYAbWPs7XW3Z2pYAuOSdBPvLB5U0BDJa+Zql7i0x0I8yArNGSBEvjsqL5
ugK8wHijcW6fpulrzH2Vcksy7OgANRYVfDOWux0KrCt2ho565YQfxVUEFWkOwGlq
58qpgyzgudStt14Yd6mhWMrFwHSy5CrhQQCNI8CfpRzBdZtaNYw0SyivawmFrN/O
Gqqo9VYu17YZEVZoH3YeTqJWdgDFMKjD2sGs1/zch75t6o72ZS2DDmxpFFO5KiqK
Vgkse0/u5GL35Ixa+DT8z7yRYBLNQ+Ar9krhsu08o4hZvAZrlvxIScUVjYCU0s5V
vNgBlNeagTFb5+m1dzzMXpl1bdGDyL7isMwuxHVbL8Lci8MDh7FKsl07Ebqr9a4J
pto2fT1iBugMSF/k9UehtgS3ZeQCvCXFMUc2nzMYhXmwSl6sWoNWzfxOtp89Xne6
GF0D9mRN1V6MQ9RfgvBYh2nKhIj6tNxA6s1yvK24NWdyFWbLpjnx0PB0vhknDghH
WqMtgKd1a/fkreNsEd6YyyZ0Na/CbucjJPZXvYIrCLzNR8iKtj37lbauaUbI8H7E
m7nSP8RzVS2ZzJ4z8mEKqGrwKfe7A8ldcz2osZRraqZvyS1i4WhpsyVDo+7aFIbU
gzS00Uw4jI6ON6pFNxKbfVD+bunuGcLwuAlJ8eynkLo3nnA8D0U8lzD4x8s1QkE6
tnh64Og+w4hsNOyTUFJJpAzOkoYOe/4Skn7ujY9wpVroiHN+S+TQcc7QJGu6ZIHt
4B3fARwrfB74isVstk6gjSQWRrwf7C7i+k/H5u/R0Fs0XITDlXS5DpDWT35gpdzX
fiAlfCDFoR40z1gpXINY6Td4t9yb+RyaNQ0UDmnZ7RkVs78ViblYlpIzDPzqYU/E
l+uYxT6P7fg89IhiWi0FNp8smqTXdlsbKa10AiOUcBbqvsyTG3Etfytiv2QVjVnW
yjQCYq5L6WQni4KiQPoJQnV4rKyYBooRoCL4EKLw9ADz38M+DxIUdJ2a4q9H6jO8
sviYQ0ByobzDjRJHfiudN3nyF+oh7mlu9gIV8Hvci/cF5PEHH5aMRlUpVW5tcxfT
62y31kMmWm27/ZwnOjg5lJ7mZcblkOyMzC2JA4ZlcbPWStNROCZrGPPv36iZbb7C
OFZBYR9ecmsgMwxRtCQW4ntu0HTetwPodMFWAQNfk579mimu+14Y8A4r0Vc0Kllf
RdFlRUXpUAISBtlik1Snv9hCaxL59LqL0lohq5hZ4mxeScd42GtWQVq44NNggq8R
wFLF02TPnSOwHi01+eUGb/G0K0wTjmotTtlnN9XGzQOs+w3NR3GS8TxH3UYlKdYq
7yH/PAEWUSJ7OhsRSaCl1vlshymufY1C7pv9fymMK9Uyd51E1YI0fTEHRpV6M/sB
0AMGoDE3jGcVNnmDjVImcWgUzLGTUKM4+liWVh/GvMapuxnXFdqGQbJCg5qAaNGs
a5q0oN3mmoomPyYLOAzi5D5H3TRoTHii9tcFOzHjShuwp1vHAZvy88M+QZJP/DZY
vh6eaHMzwEWV/kO/bVFrQQVw5Kof0TIiHSnljOORcfvB+ZsfgfLxRJIcmnNIjasP
o1HG4pNNAVZmEUw1cZvAZAPQ2zo/fBadUZjpJgxh/E0kt4msyhNFEriJisHW1MiH
3mLON7UkXGOd9QGUBGg1mFl+OE1YJGXRsro1vVZDle1bsfxPC7Fd/kbFG96rwmWn
6H6oyxyBa+sCCfiFGuAd/zgq8AGRvxim9kSBng87PngX6MenOD9mb/L3fJhLU1K8
Wb8nyeKjotobmUvTLUN3U2HpV8gpSiUF/6TkISyzVkkhf8lr2Opu5LR1IbkjKp0H
L2SZonKAFGds3eAuFwHxxlMmMS+6OssdL8/pIRFsuS9brXD+WRan+VJg/TDwuErr
wrUFCclq4jNxTdr3K52jbDs9T0yieR6hJGiw+wYT2daRKJyyYN/LnRxlgzkQK66o
E+Wsp5787nWUDQwo7nfx/HCeGvWKKXH4WUcgSPgV1U5j3PykRFENelc1w5s0OA1r
YabfG4ib2p4eAAit/ipl1hH/jQ0OgQOD2o/GGHfQ/QMSdXxDg6BBEHOzTAV2fk4L
yn7ngfoWCW7vHSbeWXtwHLf2RDw+wfoVHFsxxb7JjvpzhjJEZs1O69Ojzs3VrpYU
5kfCmjDBAVqVtH2x2M+B93n2RhlWPZrgVqs/M49ms2you/Nm2/nZtnHDAmjaMwd1
ny/WZzmJ2r9MLW61U0VmA7lu3JpAa5sVo0Rau2SpucPQflbF71eT42ZlCf3zYT7Z
gQlXupaoiHMolu6aKN/2f7VrEuamRoaoUhTci88PpYjto+WcQK4V4p0wAZhp8EoA
Jl+lsL+PrPZBhJoAWpdsFMi24k2WV+eLyrTe16NJrAfn18Je4i8jQGuU+eQ68/2y
s+CkAeikn8D7oLXNUxPcUkYdPeQU0bhoOiYpBX/M+TbyqtKwy5nt78U0tuQInIwm
fX835j7AVAoR5cMHXjGxOd0VC3+IU9HUOVXwU6O6f25sswkP3m8SMbbA/xyPEbBS
Dwwgb562Mja0d0BdqAcG2DPiWP5eoFNd2jTTy/iIYiGsKC5gSEK+0drX528C3Krq
Ja0se9RFF/cnh2ET7jIFeN4GBtiTWS7aoDtrg05n1a1Yz7Gq8lGaF7QrwQBKI2R2
nyQYlVr/2/nvxtV0z5R/e8rdVqYF73yl+BJ3SxUsRWSaf9Awp3ErgSmbfFEE9imu
EN5K0O35jmQhfwyOI9+Mhzlfi1d1oFFF+fejQQCwfJyJIH+tNVGr3hZkZEMPS1Q6
3feiGB8BxcSa9XPz5v2Tro32IOjAlT7LYsU7MFTcXMerk/JTGINeMmU/eV9bf46g
pNN/fUxZh+hnF8wkMxLdmLtV0FqFbsAh/3Qnx1Mv8SBQcriuRQISZlB9dhT1D6Uh
KUyfkSqnRyw6upaN2RoOCh0nJl/3siZsHQwPW8bUr5S5zB76F65jiklPcaILSC8O
Oc851/MNBOAmihDO2XcnJ9ttB0/+9MuEDzHBUHGAbyLZYOrpzo+5CbzoTKLMWkHJ
J1J2R7Vxjj3OOhsgNErrSG2klfHapG1R9Z/gzpd48zV1EFWszxG7MaDafoVcZ5a7
96tdjgqGpL07WQbsE9u01L+9BTsy5WFY2h/SzE/W5Qgz3cWh9OgWSt6UUkmevO9q
4EloJetEGg6FiB1cFcge/QfkFk2Ehxf0+uD+ktU0/QOPp7yMNhnhW5/X/UHzULbm
dUuWYtKDiKOu5g+OQ1MQ8V0h39hTSL6Uv8hXr2PahBuWlDpp+PosUgg9GjBrefdf
oLJniYA3IQr2QKuI7vF2xnheXrfHBW5bwZAPm9A8uz7Z9+7/USPBs0SnvjEdkCly
XOlr2J0JQSoRrYP6dNjAe8dB8OkJ256eiizEj2X2nipPAfUaVXcM42xQX9cMt1dF
Os7SLgZcoYPNHjTV0k5kT0jtSnn1e9TTanDPkJ4NEUgU7O+WmuRRdoNA+B5k4SFn
N5nHSnrlbTmlSklk4MlNA0NTHsyNX49gRSTrS9egZuwzTznHHUMHTXZXc7gugGrT
DoW4HTDxNaZuHeb4fnERRnup1mHrbJHhhLBLQbC9uPMEWLXLCMt6N7Vt4/EknZQ+
eVS3h/Xu0nzNnoc1bauRWjKfn0Qv+UzQa1QYH2RT3H1nMaiaTeOMkhpiHi0+ryse
P5THXJJivqGSQtUpT+jvbbnw+X5vhpezsY931JtGlEz0r0xxbQIrrh+1mvEhojoe
uE2Ev2FFBIZGidAXdcCuJ3985cO1YQ2SGbfWhLJe+ckUSkNaf6qhq5oo4CkHaYad
anXQzSr9kxMmmfs5OlvyOSMOOamRSo9ZcL7F1ahWWIZz0QZFo+quUfTAU8gsYBAU
2RJ4fj0ANbFNENo2xqSH0YMOzWUOHfV61ZE7LNv7oKfG4iLDChLW9VMDAmRSc8MN
8HLDS5O26VOPsOvRF6H3wBqgVdw1U9WlctryI05CN/z4MS6qIgmZVPfR1YBgvAFn
CUTFvj8lvymF5HlbBfzkdovn6mMMCx1EYS9TE2C+d9SgHdM2SqnDG1IWxGTiYque
Fuw3PrPOFB3fN7+hf67bDAu7tFJxIdSpZbQ5/GwL2XdlKUxfLtWknmTUXWS5DOJ5
dX9oEzNaGO16EeKDw7wDDHwT7eXwo1M009rkAqaoi141ItaWUZ81hMgQTkdRna3e
Si8b45pHUg9ihaQNNkzQ+Xh0qPJ09AhiJzYB1J5oJwi/jDwktwpX2njgZe2r4mUX
ruAToSciKQdHHFlgf2+0V96YLuuEW5a1QChp80LS5OhFadABgyzi8S3OwxD9LTxV
mp/kNrex9fwuplzhcdX6Q7xxMC3wa1vWd0snS1Hodg0qu6UjVU6J1xm6fAhBUKKQ
8MzB95JVtPjptY9eNArmGE/lazTof8agifzBYWDF1QUVFfowAo1UNnNel5di6tQ0
YgHqfgssmgr56T5aZf/yGlTu+1lF0LckyHUm33odzliakml3GuX94EP85BsJfkQn
z6zgSjU8+mWElw9jG61zkeKqeNpvBZWPIoX9uKb3pOp23ufxPLCLq5tuiBoOSMXl
GT1uG7lx+y7+wSDIpHjzjuVdzJ4/Myc3RnOsej5h3Ama0A9+arrkBgmjZUhL1gza
DOpQPOiwOMU9YCMQByy/wnOZI1E+t5nI4KDgNMriX0eTJ5qiUX523qjRdrXsTU2O
m5heF/do/gA0djf3ucUO8ncJn82KKaGLpPKtWGYjRSAtiNziHUsbXz3rlk9V1N4Y
Y3tlIh67BTEjJ5lOrITEZyPtYm819jPJMqn61zMijA7JGRTNOhTrFfN0+E4/XQki
RUmVVxBCNUcIiYCRL65lPHDYXciGDivEJo4+tjkljZKRR9jJT/G3ooQOZkQsQ+/V
8CuXx737HBHur9kXh9eKpqsajgAsGHi2/6Nhe6YYd4YcBWCa3FTeBx4VZ+Ze80sD
OCUEodiTho8GN9iCfobFLq+BujrHliVfYUPGoqmYqHd67AASBDX/Xq9qHyDvgM8j
M5jwUW9vTp3k4GxSEm5vLM8NnBOFYz74fjNFl9rf9HC0Kr9eNCQVEn+FUI4F80nH
lXFRK8vm0lMGxmfsYsPESnIf4fwRGIxx9pOEbJyPBBzndqfTVXueTGrLhNabPBeT
Qc2I4S9IFncZ4TW7DDUxcCklQsB4bRocOFMtjI4j+QnwRDtcLPSbd6gyiy4bHuUL
pG8+UBoPbWGPbcEJFxb4GeSRPz0EthAY3Px08SYUjVsuqW19zeevYrPRXTfEJKxK
fsdguOFouyvgzFz4Cdx2e2H4I7A3uuLt/kXUtZfFF7yMPsIUGV6JhnDEHI1MKKxl
XiVXGIcSzioy1uLDj54KPzU21TMRPSKhYSS0rMpFfdCjcgUJbrk3b2UOBG5zFCBb
aqmbq3MFqlHC2CRaD0nXTTiFUrTaoGChW+ZwzI79zhfNSRj/LKMrCcukEVf9qFVw
EYAla04mcCNQQFcCPBzcXFHmasiKhZ9Oqyqdjx3R3fSLovhW1UpEgtRmEKWMN9aN
aLLuY+eRoUKFJxKOx14XtEi8i4HNAGhS94cAD2oDeq0wdTLZur2uM5UEhvktFU9G
KjODDdsuSJbbAeCLw21HnsWQRJQd44DTnanPc6cwA66FeOnLv8xhFOBkBFlIDqsR
dbcKPRWW4Lg8L3bOu2jgIlm73rm7Jpfsw+eI41eOUcbBYryAWAGYaY+qeaBvsst8
I1V0OFRNrj5yO1/d8jYgqbaestdnkMe5Ln6zHalR3rcQuopMq0fpxUGQSf5uQKd1
GfxpG/NOg4XVlpmLMEBhGd5rw2XIi70If3HShAq21wbBI7buVj+0wEG9ASwvOFa/
jwWL5TdmuWjSHea6Xn8P2W1EgXUmv2X8+r2PGEYihDCdSt32nGah+TqOmkZ0H/6P
JvGOebWKO/RmaqAMlRz5wTw/bzjfdZHd0tt0FQrCHOXAv/Z54cuVQ+0J1yIWDh1J
sCwZE5GjjurlFO9boNcICJkCGIxA8ww8HWak1h3axbvSboCBQs4ZEFmFJCA2/Vqf
0+1FwMm1rxL3XV/tLn71+aVZPXRbw0lxmMwbSJidcIpUaHcrmk52KDe4JT6ynpYN
YzoglHLr7pTa2xHsDQNGqUOa1GE3RzlIBhn9KA7u/hqC+UkD8V/tZ18abOQQEKgR
uriv65hEpAdeUN5et67fDwIE5v0TF9fe3x1ee/QyMKDnrELWcfWF0fZbQuzLTUM6
Mnz+bL2xjzOJEq6963nDYSxSPsOK8iQDIYgn/CqzUjcYsu/M3H8g3+DBXIfejJ3d
1c6DRpgGDu8kQehCXhoBBggktdH4qQc/lLSO2zRg3P4NAcjc7yElM/dkOxKxh6ak
Xg+DelglkbCi4ABjYVxxRR/pM3nE/b/rGzCDnQfwoiMGCGOQhPb2HvbUYNZq6VQB
P6X4H33bEpYsRZPO4+URKbEPjTpkHyRu5H75GxcmxX0OnO1wfeG6YnI4RzveKP6P
hM8VjTHKFNT4reliKsdX0vypI7Z1XnuW4IvBOxYvVeo6X0tioagdSyyVAb4uYSrU
KBS1JKh5xeKxv5uTzJEBYjBpxG9D9Pl1Y03JkRMt+HxqoaCHa5sK8Om1WlwHTsXU
KfNhqLJetLbzQlvrVqsGl9f6iq+IP+Gm4qpRjatxoXd2eY50ZkcEd0Yt8cP9TN49
deAc7uIiu3IKBuXO6KxXUBysIheUbDCy9NbVreuzhdGoL5+2LdRIg9VVraawNSYN
LRkx0gi8M5xQXhANYjlsvpXKrNcZTid5/Pv/zpG6j/e8byyMGU0apdbCZm2Uf253
jjwymkRh6e6f8ejwHxItClazN9j1YPgeoS+WIyPiKqw5u6sa5CTFzxyo8cX8zO8h
mltFb2eWzJd8knHBcBalGkn6NYWE7kTH813XdBa4uzEPPw8waW9wiJFGJ9yJEfi+
HqJDCiUz5FVnpDL1E+iUaldhItnbprzQpg4/jtYmZsvzUy3bjC+ApCEdijLWZCcG
C/dtGJijtP+L9kzkKPahukeI0m9cF7IPToc5uqn4wJeJiXyX/jWJ0qa+RytxH3hV
TH1aFWEoLKyYjQkSD6y3paQDebvexJ13U+ZPDBYqQ1nFtimSbhS4W/gdu2lC6R/A
ulUVyQbT0b/twdbTRBayOJvyMKTZhJ7LCLy/NsAuf3ZA4EOopHsOk2VO0b1DmvVT
FQBz3SSsPEs+eauGodfCa0Yz0sAPeLWVvB+IJXIg+GlAtxAWaaOjvLkzBBUTQajs
1QlxmlHTPDpxhyRHlLb4FoprzIdmawkmzfH+ZbJe7XcedXFS+aNDOIPstL/Xci0k
MzovCERotg1fqyxYfJOFoHsXR/ak8jOoyDZ8xxdyvtnNlnjvZYKwf+oIb84JQZy6
YYoLHolp0J5TGJ7IT8kemRnEjHpqFDj5SvVbo3seLDyI1HDtSWav1DVeOYNH85gQ
1w5l627ThvvG3iB1GufvDitx+S9vFNcAd4BYG2wJ/2Yi+bhKbD+sWZDaep07FHTU
+yluNMHXziECxOGRy2TyWUMqadRSJSscDJtZLsCyL3i2hEjAKbYw1z9vdKX1u9dJ
E6v7a/n9isU95Kn7cpUh8hpQ7H4JtyHyuKgHca6FsfevVUGHypWuDGr6uRkELHO7
9lOBeyyOQq795x011PIKDYdquaC5/+I4+6+a9B52RrCOePmLl5UqLjhyxem/bK4e
NWkkZ2vBrpKwQXYX5dDZZDkMIrWVtALmKrttgF8H3jnaQGg+VibyYivJ1pmHni7S
mIXVrW8ALPTa544bL92eUCK1pju2ec2uRKvvJDULzzaUWt8VZOzbYTMcWSZCJf6f
YLzYbYav5h8HX0pC5JohJkFngD6rubYuC0wMzoU8pd335V1ZTeEGXGFC/PyhN1Ef
VJWHwwdKGktENvCfk/MM7v08Onh5yKXEFEi94TpPpvULQ8YuRCosj+bEtCdtDyFF
qIlnhXT4IZ2+QcFnV8qYp9D3teZM+9IIvyleEof6VH+EiEBPkPRqfxjeBgstBrvA
2X7iIBaGSFwZQb2G2fzEmyz2nQ0YvR8HLLBItJjOHAFlT/bmp1IVTA6/SF0+l51B
si8FoEgOTPJPx9ryO8yOMSa4KppXaa0w4T+OkUTPeLApktph51nN+p67J5BPs+VP
MhyMwBWUZW6/NeJjZfbBTWbOlw9RMctH+Z+em7xaIkyiDYJ9yGdnbB+uEEEHVHTS
aM6KBvlL3VrDeYDQbDi8qBd9LyE6dC8cJAvsC7+sDUoyN32FMSaCfYeTb02Qlr/2
BmOh95krCmK8JnNFtP6ajpmNGZkL/jI/FOTZeF1QYjPEVfEXqJa8zWdh32cb1Ynp
+4dhxMKkYq/wdCj3e8hkOpGY8TXwf5Exj2/6wdSSflp16p2i1rvb3IPSLRl2djAP
hjKGmk6VpAgA/cSTp3Icawj79DB8u7S6nuIQ2d9RGChbVFRragIxTvtJ5V+V/jW0
g67NIqma2UsKIEL90+PxBrVrctjOAOiWuPwnCpBmqLfMUQ3lSHcT9z4LW4VLV2lO
6ThIZPyg4SwTMcjySp66KznjOQp8VI8nKJRjsQnruf7NHzDH87LAvnIyQKeQakSA
z+WgBuD8lNQZJrS65Td5xT2MKEXtFxEy3cVhm8uNPtCEuAxY3fRfL1Zc5Mkxv9yc
mZoS40pPh2OO7y6v7X5b+LvZ+kQx3DGP+juU5xYA61UWHKV4uDhRA/UEmRUl+N2Z
dwaThLklRUD/PVpNQjsJ19JAnT52MdWdoCG2DuzK5yns3IfrbGpzyeqX6dzmNw1a
NhQDwaUz+TvuY4/1FAsPDw6hmWz1hy+RTCo+gj61uVNCrG2syHEFUqXQreXOny3o
2s0sRgfgx+OXLOZcTilWtMbPPx8o7WV4q91x6kd0gEPUtGTQtbbPhAoJMiLmkrkz
cps6MwhIoH5DxuDfEst6Rf4IFs/KKx+V8nvjtjbs6HOkB6eSKHRK20TSHNs+ECKk
X3S76h18tO9MTQHgOe0DZpvkfddRsMhNz+0/mbs2ojkxxP4n8fwDuvf6FdrvsRwx
wVYgVSE3GIzvvMY1l4vTO9c2BUVmgOUW9vNhm7EN+pQ1XICDceIFhgolC3Pi+IX8
PFnFF/1S/snjnMp+NqAYA5OEiE+jR2G2hturZAtBJEbOh8fo/hrI6rcU3igTWXEo
II0tL/D+/0T0/5GFtgQ90S+H7GHTwkspcwB7QOSau0gS76BEyBfB9QqImipqbExq
z4JkwMyrWg5XfRXWCMRExngT/GQyoG+G7QYhWVPS7XfxpqXUJbanMsXqjUEFQRIX
iwb3dInhIQdBA/SDlTS1IW5upfHT/uLcIMjRDAsSKMEl1S+3l/nNQtH+TEhOIB1z
UcI34TrvWgERvswSfS58HPqAUixz3MuSoPh2mKo7Y9P7MWx1JfXqsjQkLFEQGfH1
M25aDXkbAkNZOF7dYvQbrwLvFceU5JT3ThtUi7wjOI7mnkU7CiRwYqzve14P1HeB
YClsd8lH2JGGPZvQnTDVykGu+xfS+R/nNTcgWyOApfq/DZsdv6tgHIcETQ22CqDR
XEj7O14wLCVYwAcx3abGQRgLFzMKL9w4HOX+vlvsesLLGgrXz4Q3RjFz9g2yALxe
jWtSxgqnmnjFnUcM02wjU2fncPcX/qlLGjK/S59S/GM6koYRnzymU9jMwJotfk0k
9ef85RSigXjel7um8CgFOxvQjInl/mFgFsVTYFdd4Y9yv4lx6HpiYItkPbsnI5Ex
A4P72QHyi+ov4Y53eb0PgmxleyfdSmlmCdrc4DBsmvNpraxM+4iexGiAg5c9Fk/p
bM6tTdIn1vMfP4HpOKGQ0qe5TqaL+1gfR+kH8Cd3ODnV2SNTheIOQXBWPP5uv9zu
GyBe8LpIFmvWrJuFJRAn/6Y9EVT53EqM/dsaqyydBjaBectPIaepDFPqT3lZw28n
RuASV5GczXSeJpSMPBZh7mt71CmY04q69koWaTTpRx9yaNKwguBGHbzCYywTWQk2
vqJ0viroaLlK77Q5oWkKh6W+nKWSQA1VbS3uXyUgaHx+kicAXQ1bToiucIrYMBDj
1cZXFk5nd6B2k6DfVgxjEtHo6LlXJugLBGwOatEKjeKvlwx0VR91KS02TSCaLY9z
fnC/FJ8z66AvgACkXK1lcj6lWNai/zArq7g3J01QB/ChVg7SgJ/LfHElzzUyHp6i
mk9InQ7p/pa/VOPgA8nCVYPe8D0yUWUK/yZyHdHJVyXn+3BeZOeyTwHuZaJsgqh5
Fd9nAHTWIDQbXNinwJKvNdc151XzEwaKQYVqX2Kjd8Ly53/6KSc/AKOfUubKYo7q
q/rQCbPkVPMS4DJkEoyfIZpjvEouErVPVL0rH+xZfoiGQTKoajNhoH7YWj7mLxuA
ve7w9GHpM7Kv4RrhFibMLYEUB1DDOevxTnVHtSKRHcslg3j0OaOS60AtptxGdB/3
FH1WXlQ10tPUw3oLMEV6usf9m6r+xeczS1xVOMsDIzIDuVrmt5AgkcyUh/OTac2V
0bS3GqLshcVz/agsxEikOs7Nyb3jF+LowrXfXun4OzZm3jcN6S+NSG/iWDsQ99UB
rGEjWb0ld25VdBXyG4mKZXYI3YNUMhzLD/oBP1gsb2e2d2wyjKgImye8870UiUV/
AID/e1u/LynG/1teQsKzf2jy79kXbxjEIf4NfQP2RNjrLfEaKNbSoTjShl/QY55R
1n7bRmX4xmPW+OYXIHMhTXplvtxUBfaZEXRjXcCfcftarGdsbgKt3aUqjb5xWQmE
4QiK4nrZGe1HhNQb74vvRK+PvodOBBESqL68NjH+F8VEGZqvEqkntiH8n9ranUS8
hRjY8rPhSPPWyyql9lG1zGticCTD+KHGKAWCgQGRsDZl63/lEtbK94Sa9U+4LgJi
X15otQ3fG9Ai/h/6ZXnsNFBYEwxDWUI9JSgbTXWP17ObA9dJENJP4OKGaAMAdQdm
asgNs0rjXVySVsN3nzGO+zdEiYDg/vmw5J2a6c4UGguF3BWbpB5KWL0CEiDMnrN+
6bSTImwP1pBSdQ/huvRQAj6s6RWjdeKYuCwAnpNtIA241nyV2TfT+7LazUfYyki9
wIjtBFJJH3CutYmsB1oaYU/zjJFliYhTR6glfSpniHcJVNVUyF6tmJo3VrcyFeyd
6dlKnH1mSSHyIHXq70ZDuMvfkaA8XUy2340tYb7cMVbuwD4TMv8wAb6Sp+ip+y9O
U+vWFPJL/lCmSbwPIfKJdc0Uz+v5fk74JgmP/OlcR/K+Lw5g/zPcp0ajiehJIVbS
TGvy+/nnQ/pLXNSyW7w5aomNAZbG/v/7ABuSqlOsVbeqK0RW5Pn4zje6ZIBvTNh5
HHgeFkGp2obFRlaHd/LkP9TRsEpyFQf10onSHDORbBfI8AU2cNNnOIQ5m0DWtgj6
1/Tu4fANtzKmqtiLahQ9eGM8W28bZ3S1YcWhZlW4sffi2aw5PeqSlSf71JXCVi2d
QHN1bv+bSpwB5z9YB2Hjc7Ry9EAS5Rm3Br0mjosdhqbuYlwvasazBE1G0Kgypyum
xtNnVANcEHSflByvvVfFOsdSGyALBP9mqTJjPgHezWNN6ke0iN/V1con+mFkAO4B
oHOFds+JXhCf9MgmGZGpXKBRoDKgtSd3ZA4uf1CusoofC5ujHpeiPlTWeFShVxvG
cG21BpZys9g25KJRVBijY85f7nv7JGGFSILuRkLnwYAxVAbOFRIKcFKVjcDkL+Ih
b/MTrCItOO0YnhX2zRVySkkQOAn1b2QG8y5VDX1fH4giaFKtA1RJPb0mQ0Hzrwrq
DpwDt/oW34k7iGXVXdO+zHwM9kxTEQi7v7drVXYy2bbgSqfr4qbMBMVnwp+5EsFt
b5ywMXgfb1miQ1EEX0DDFP0OGxIZumK/FZZKA6EOkqfIrSE41TQ6kPwohL0vT+0G
OYrScbWA4nYhfnwkIqgoaZPeT52cUQdxNHx6+7TDvHZmY/GIkeIwwmRxB0/UNMLV
FwcD10TyWMaocZSXrWJdaEo7zja9s9sQadb29cHrSa/MEEY5RoSasC7HO8BzTj8U
3JrDo+t56rWjhayaQP0cbhKzVf9/HK4szgDFlj6f+2tXc18537E+weiN/P+8RHWM
TyHpq8hD4OTlgLKPPjKaoXpK7/tZssFZmSoIo3odhEx1PS/hOTR5Ioy1Gfg6YT9j
LCj/hIx6BVQZEWCHDHCERufoOmQmkdiiyhrZJFIpFHPGDWt0M8trVCsGUaCBefhG
saHZWHM8Jui7fHV9VCmUOduB5TVI5M0OjkQIPhuA7obZJBCTcraeqx/oltxlIWAg
uYq5nwfyTjsK1vwBsuX/hk0ucdnZqwGoxKE9j5dyFWbUUrCPaFmTJYFt/PKKiIsk
+rYf8lP9i1QhomYaotuoVtO2M84S5ySIIkg1RejxbKgRsptro6Q26JZcwEn7T9zt
nDcyuyp/WLUHRrYqVptoca8Dt+aER4ctx3ECkv5AKbovhqO9Yk5+na/wFulBddgI
owW5STkob7tL6hpiiTXxjFPP/uq31GYgAiiqND28nnidefRzZSYUNr6P5TnAM5aS
9A8L63/fylHNhbtCNaVqwJCsVUgylwb4yCCR2a8DL9rOLLRLRO7iiniTVsn1cU6j
WwAvKMo5+sTgKd3IpfOEtz8fQTVmnvwT1VV8h4uu0QEPp06vb6QP5ys58n7Uq1Pc
+6HbaOCQwMI8HK9k6KLxe0D5NLHHH6hbwXYIPHc7aZP1c8T2RG1gwz389GHZ2r/V
VgLLqtbIwkSBd55zuTwO0I0yBJ4twLEGRh8jq63A/VCL3LbHNMoI9fxg6V9GWlXH
oJbrIuflQJ8dHxlNFufFiWwukzFGZhp2BTa0f5FGgA2VeaWoeVrIlSWYCon3wMhc
duEaoAWIkAKD9m4xQdC9ZCBXfeqCiqB116c3J5kOElbXV3xYUGYWT3z8kYLJQt6Y
WQqJVGex7GIdMD7QzSsqxTDP3z/FEAAa5hd4BDqAyBMOQqkSKD9SVxyrNzjWz3IV
WT8l7uyYjSt5HyDVmjsAYlDLbv50LWXK9ZGCYAyOeJO17fHiXk4nqGRBSmY5jaB8
vBx1W8KkebmZbvdkMCyfMhhCLtNZWK/LjGZudRCkGSybJ8ZoURZFyDjV4l6tLlkE
KtBxJj1NWOwnktjgdyOBNrRmFKfDmy5OjVBqPlmXlRTGGSx+d17lzFUGbKLPSNZl
SUXY6611CrxCabYxfNvWGcB+0XBEXQmhMGlpZy7rMk/MCSb4JHXenMaIPJQrkCMj
58WxStVx3DjgvmypnHEgajfSQEYtA1cBFU0v0cevg9/vtCY4gAUta8eck78z5V0/
RPILTyDFL7Pdw9GDkJg4VuhwDgfzmSpaefhxunBO6UB/Y8zLR3lPmVDCeH1gmt5a
BW9BVf8KGoAvJR4To+dkJq542D6Kuapa8FkNXkvM35UZuZevEjH5HWja2Uh/e/ev
HJpK+eUNpIFzN1X1duulib7n+/kjNIgGGdCCBkJRpJWGd6FG5uH+umr9eYhuPg6n
4bgpYJ73ykptW4hl2tVTCm9lhuuJa3xj1n1Wx7sd3cZqEM8jjkeR3KI1fhHtAEf/
qZK9DHf8m9XpPY5Te+LVDdVrKnUTKgiec4s0K6yOM3HyIXMP1F+wGcQ1FYK8D8bm
VeurxaHu8EzpG6Ax5oITj8mNi6FnHyZJd3v80d4oh0u8YnKTD5+z55gNqjFJe7Wn
ryfhllQ9EQBHhs867Aycd2xjd3+heEBrz08ed0AOPmpz0+xr8mXRb+b11UjdK3R5
M66slASJPHvXMVbvjSoNin9NLrldF6WmfOTE4IfQTUBOsrYaMFu68GLLKTFiL9SW
Wr/ETp8Vk3OOsYbObg1mCdlb3n6QB+M6pgM+oS5rHy5Buz2V4ZOR6+CNo8aiwFSV
dVdiyD2f3ZayfGZ7ZXOnc6hcaGbANVCo1xRq6Y1xeWpG5M3x+5AgrUw9+fsyKtGN
hZK7I3WhdJdWDXvZyFT92XRIKDnX1TEJCyn2vvQ8MmAHhIh8yjM2wVm7oR5eEVZl
y2IVTSDNQ7pdzijlr/9Mg/+nSUS7lW5EtuxHKqgvcKwSEZj3/Dz4zsg3I5tvEK7E
bgG2IayqB4ZHS61T7/IvX+btcHLaqtO5y2wEtpNiRwHVfG/zlZwUKc6Ohl6wFt3m
wx19aFRvWrf/rZZ5BDOlRmF9RlOaXbYOe9b8yooKHBY/YL+5v1zsTyYwCxBi17dS
B4CpGfjw/nzqFSH5aet2sB7DhbSFMSrhgGKSmZYVnouHrUHtMbXFOAd/H+w7iQlK
RfyK4K3jZuObdCLoWN4XDTObLvHLXMb+KVbYt6U+Ot+XDG5Zfn/ios5jGrRt4/vw
VhlFg1pjA17YxYy1fC/GNvdqsU1IyBGT5DkdEJM7ZPDTGu4lCQSl0V7qVwoNkeUz
AGztrq1DIsuNt5MuGBr58Przg2zZUDRkpvnR0zizcNEt12uRE7Z5pIqGLcLx5PS2
CFeXTwNkIqdZM5+4v6x5VDmxrAxso0Frn45mrczOLNEdd1hOPUS7Lp8rVfXVwb4i
/95Cw58qQ8Iqamtk6WcAmmhzy8JCNcRJfA/6w3G6SPxwfc3qij8WyKXUqBquruxe
9rRfAQT0Y0jcpppFGomKrWK/CLPgLotmugH2jxesFPvLYrzfyaRdoUEriONO/z+a
44X/HUixuYCUG0c6uSDBJ8xyds/8j08Utz2KwFpJoGyVZpVNiiP9C4+NgdU1GWUW
/gnflNNw6sSV3nZWCmtGoI+6zrrN+obIyA+184lhMfppTDNshu33qnQqC6Vx8ThQ
goGusyYrKegCUJGCcRyUzjdPiajbBWXdSX4RcLoNwSc3oCkbQ0H/rUsX4Z0pEf4M
ATn4av6XVlKdvZuNbhoeMCOFzC9aPcI9iRGgoo/vWEIqDtUtrrgX9U4Ht96z0w2H
CJ//vMYDjEyXUbnbc/gW8gugYZT1IvK1IFtpHM9H7riBR8QXwoaWhO+/MadytwCl
+6UYz91n5kZtuqTlJc6JT5yuLEbe9GWAtOzlMkI0RETMfLN3I5yYyEEhYtk4a0Ln
KbMTpO6sa66Z03o/1wJBG6XDghfT7zuZoDS3VrXbqhUm8LfjS2hZ8ooxShpO3c+9
dkfwcKOxeEvHOb5keACzK1U7pj/KwkGSsBnw64fuaRb3iYDO0S4zt4AkZxWVF1eB
3viphDZw8qU8vJClDByKj5USnPax2J80lDmOJEVrGokhNYXGI8K0ey/RUiaxRHe+
GdZpR7/iPvpMFU9D12n60DQ9mqFMfnp8PDkKyqlDkpWHrOJsQQ8EPe3FLa/H/zhK
NK7nxx3dFpDpiDC8hZIRuz3yNpW11qfxGxYnD1LNgmGQkKGBbk1RYDRryEE2t8m7
MW+8HPO23b9A6ekrtUiX1MNF7afdu9ZU6lXaUSkFX/bJuvZHMKpJ8sldQhTU9n8R
t/7u9f9RPD5MLGfbnlOvsEiXFvCGHNPC8h270RwNZht6MLrjlF/jYusUDwuxKukp
0zOQRic4NFh0Az95Wblucs2/J/DFCN0V24CmRRVlQqBZP7l+MVl7i9AR5QT/cS55
mH/VgWfjzCQIigKVmKBUAaZwkBgQvOMGJPBUiQKSuXxs7AMdHxU7m6l1mJuPiD9s
CnHJdvXo2HMW7P3K5vnrEU4gGSIEnOQ+mxD89SmJgtVkeML8T4SMfmkk7nzRxE/y
4lZKcWvpH0xywpmU2Dm8eoCkXIlTf03emI1d2IHkZoWIv9wWtnOS+wCQzD21QmIN
OMIwpny/YzLmWv3TQ7eHxb78MD7vKmcc2klhw7V7CtonK0AozIEs/ttlP/4NAsg4
h0WmV3qhDittodxgkeA0I8CvGC1bPLJOaqqOy+ZmGs9/meuX6aqdoI3k25x5sRWN
ZMMg5aAOGyhXqnW0kn+ZSRcowuwECmgTFVW8U4RSoZSOACfyYoXvm4IsRrwD6w15
nYfuA8nteiDnudHgNXzR2Mv4qdEankUQ+ZlTVE2AxjdiSvIADtXGfpKWK20Y3iZB
gLat4RsVZPGAOy2Ef0XdDhYpRZfks5URJVRpiDQmDYAwnMID/Ymr7iLNyJkY0ZhS
EzLLxHwHdEdnHFEXWcj3Mhdx7Yjn/ApTIYb2ebNpX1EssPQf/l27YSrzKIYmvoCN
RugRmzdJZQ6jBYWVZfu7aoLHMIPYAaGp8D0S2nrF9dDPWRvlOBCID9v7bKMF/VPb
hgKoIxh9AMNfD+Yg0woKZ4Mu+zg6X+0pV6o9yiPgpkh6crVxLnDTsQnZfu7VRN80
zrW2CG7x8KTZ1pD0sD5Yw2hyd7VEMp60Kkh1V6HuYsAoc8i8iYoxDBV1wYwdlumg
JxPI+jYbPwyH2L6Au44rC61NXhjwjFvIH5CSmJzddtAbDQd120oJ7g8y/eeorBfJ
lBKWAaCHhM0BtfHx5ntC46jCEVWw9hfjMOqDZ8cxdyi8BZWbdSih4xP1VqZtTxrD
GUYxE6VZvt6Yg1WgJFC7Ep8sK1kYh5wASrdKHkjPBGf1lDSp4VvyJF0afbLSbHKw
GxEO8rU2WNLWRY5gV2/ADYqbuV3KBOJvmHK4dBHahYV2faaY7rjvJtpf4Jl6goqd
z+qNivbj9YYMiEeGAmw/cgLH/9rfbL+9yfrh7/ljp/EbGSd9I7oaSs51LDuw5Tq7
2RGRY3WkJjEU9invi6rPBF4I2tAT4NeBgH47IkEs+7203EbAQO2bX5bVfcH5WgvH
8Hsw/ywrLbKk53WT27bhgkmij0vnlsc08OqrZzLVdY63Py9wMt7VT/VU2f5YthjJ
NDDaZ6zAmuOK7osyRmt/D37zD1ThjmXe5/AXRtl/3hkOwowIUy16MQHYMhH6AS5k
Ibn+nnqnE8l4rYc9Jgf5UEPkSmQzr7GjhDm5nmn9kknsy2esVWDZ83ZmX3ArpnwD
bzst/TwBkHBP4lHfzWs7kZBRidR6Xz/lII5dvorvzU3pwKsB0NCob46fihnWaGRG
5QzSDTxIjKlfYtva/Y8KjocgCERkhq9zprQsGYU9UuzCCuj4fBY/S8ewSUEo2kfk
DOBz7c0JsMZx/DJlfHZapdB7Agx44TJLte++MtuGT5Z99pxtN5RLmQIJNg/J3obu
JVRW0cLLh1sECjsQsj7d5raODG6tf6fLY5itYCy/Vhhz4H+kLy8CDiSdP2r3Aml3
wnmlZApZ8lXyobQlQ8wI15Rws+DzwiY/E7TwySF6ZqWQVXdmaJiOyWXfviocuVHM
kEOBMyDw3LvXR/dZnRHuY3vZzmRwZ0O0QBMw0VjPv/rc+H+PzeqAF/qNax4Iq9Rd
7+/Kj7jZ6TlE60Fje1ZsL+a8rDXjRtA1GAM4GdfrYWNL42QsCpwSbvv8+OOdnwLX
gLT13kTENvVSQZPHcBUPS1YRGsIfO/LYEuYVRMiZSFwZvVWjhY7z4IG/IZJ38Y1j
gqTQPo4LmNUjdAGUkkSCZTfEWigv0A/zXWC2E+TyD7vSryOQjbiaO6nW+PByTxz6
CJfZYElCKe+ps/Pgc9ihFoNhE6hs/yYlhuy0Rez7Z/8pWjY0DdzemWCdRkPcqd9r
kHwAaRf9IS0bBesGvAD8FaWdgdKLT61iffEYeizIXVY1rTcYTkVvyVrePWNpJiWh
CPQrsxQlwh4w3G2NdeqPsmPlSjYd0oMFBa8dqbfhKoOozvH3gYf9a7Pi7n36AGfd
CTv8E4Jrg441OELVJTE8AR3ApPAuwFXZdIhrFyu39yZfVTesfVPDWJMq8OaMqush
BY9OScXSGVk4zU8mOaYsGiCfhzbcPmcgtySEnldedzTlOS0abNVe1UFTUShK0M6m
aMoellsyMcPma/bIB6Uz9kBg6Jinp3FR1IK/C2526boR922+BWafMWVLabA0B/go
U3/b6HuHY+NNnT6QUJBNJAYVUDkGIv4ltAjr7UbiRxtGePqIuOro4jza0hgSteWY
e9ufPmuJApX5RNWCNYJ671RV4PNqJ3l4UJ2PqmkODUR5DfQuCgAF7V125XcORuqJ
jZ8zhq3hKppwdQyyKq23h2Jof2+8hzUtsodExflBtiGu7T/w6+nxfC4gU8N2nA3v
ssildHnJkuzFrHW/TEe/Vw2gec5MK8Rv+fpTBZk9XDJ7A5t09Ez4eJ5bRTfu9pe/
3AyFwk6D3vW49fLVVyX4XbkkO/K1UjQ1b7jboY9ovxf0VtZn0FQcLMed/LwkNhnC
d/Xx1xpMQ9LE5Q6gNcBzgkE1p+G8eOWfXTtnlCHlxpuLewR49ZcjkTVFY29hKdIh
xbjzUJqHQPNd5ymqhXmfWUzvh5wCvjhyhYjxNkG4K0P6RJJJzNDWXTSD0/mzfPUB
eaZMpjkRvd3OYLIY+4vLvcdskKgxjgPDdzereZqoFhW4br3WqblU+YHVdmnVZtyS
xg6puccRWnU1vdhrLfl+ORVSC1OjB8r0y0q7U0yeyHZorZ7fWGaVXldWdwYssZa9
bbAXC25jStdUzZb12lh59eQBcc1CpTpHcYwcl8FxZ7PfcYs152wOt5f8hAWMXclN
6vHP9zTTM0n1A5e52g6TNtjOUHnT51/cIr+2xS1/57mhbpIW+X3MD198ttNH46ZP
Xq8XaQW+eIn2++exnmCXVe40O/LO0Jg48LRQuWzZPayxZwsmweYdUAIBy28GMz2k
8QcRJxGe75S8N8IYE5uDFOxK78tRYuXuAzYZyB2HO30umlhRJv/tLlKq+pKc3s3e
vWb8hY/xg2lpQFo1ZaBhyqwJfo2GXmYR36Qt7q5xSC13OviYQPKnpTmVfjDfI7yH
KrHOPNw+g07Bv7qCXt2Hwc0l3Tp8GZ+GMCWVWlYt7QeX25iYIyDwAwM6mwiN30rz
d98wij1P4nqkTckLOBVvW9miJ8WtBMSP9ZpyfoUttycU3vmOXFj+gGmcROJdyBwX
EMswKfsLntw+m1mMQd5b7KAln4ITmdJljJE62W81wzeAWethizHdEqTiQ0jNXccb
33w6KStiqdBtSV4RKgueMvFnyJtcU2JvGOB+HIuIaX4dpCLxSs1MKPrSb5LMibO/
XIy6AUfZJdRAOyvLWdOLPou1GS6VefXcCAD4iBSKeDida1V7dqaXseWKEwh1oMvT
OY69l8AvEuhR9tfEcUeq8KHppumUSh/bhy+v9eNa1V6XjEuvHOzXiF3Qfet3/joy
QsQekUEVB+IJulSThWypHz06uy3hQKpIYXCO2hPMO/vDdW/Rc7iwb+KnTUhVV3YF
JYsCZagqjZI0eD3PZWixHgt7RjmhD2exvbkjBCTIQ1avnwn/ayq5OTiCn2tl6/vr
iOnBjgXal9W41RpWIp9jhruCAlM4O/F8/At+m21jGF4tB0fUjiZdUqW9xchAOlf8
KyC3Qr6Zo64441qIHKq7owtwz6x8T92+M/Rm8fytfHdcCuRDSoe9RBnoKiO1To0C
ZCX1EN5eOSIjlV40Ym4CnAnNEN6YjnwbQkHimlRl2YIUrKz8U6Wss9igtjyTcDud
1qsj9nhKOGr2YrK3pN325KpVFmKWZ7ROBqEolWlHRn2qDJEEWIrnT54m8oDwoUcY
uxUKEOCq7l6IlJMoWujF2t8Rs5MIO4zVtgEAjACctFf6jgOtNe5O9OEw8o0Pj90u
hyx+CP/Ff+RZEkAnMFnhy88TNvu7T377NxFVQqAZVChDgrFDO2GlTG6WJEXGnCqM
YpZpT6p57l7xPkWaAvSMQ/MWG2y2+abzA7xTnLMrqZL1ldjaPjZLBR19AWEMjyWN
hwntoo/UsvfTpQ4vrUKrTi4lE3ytGmEXiCdilWXWuNEw7bbG1z8zh8uOiP2C1MqK
i2OTGujQI14c/QC8Erk6NRyxk5Njy8ctUfqn+/JeJSfi8+25decuU7XzkY2C7NJS
0foyYJ4LhBWCngGFG/p8hI5hLGr8HIiU6UWYoGWQZhCpHK5EJNDs+sTv6pFw/jzw
biDPbqAMDqLz57lZw4eERR4PElSUq5GKciW3wHprswIeZvo593A8XmZniVkrtBmz
Gu1cwv194PrUQpdnSWKA6RWN+eFrnSGShk6WLPIMXM/hco9baLUoOqDOH2bP98jX
hVH+sZ6ydcYpGqI0uc9wgtswN94Nr+OtUV6LSVgarFyT1an8ST8Hp48Wn6fD1M0H
ZPyycV+QYfnq9ZFfkeEUt0Cv8hlBUbU8fNmIoOVn3lSCt6zz9AfXfe7TzyAw2FXM
53LW7xORvm8tRDvWvQimJSYAtS0xmLnTHpCtBT2d2UK9k9B3fWp5UjvUE8DPG9eq
YOiva1OvnBuNk/JAzzUoFjtfps24u5l3a0lt/V9TQipEFy4GzdTvRHd4im5+Oc/K
Fpquk8zhN1b3S/yeB7l1r6+dOo7JRvzGTYjCpf4KNHrz8vEmg0ttWtX4//dxU1sY
J8hCpvrpeSsj4oU59w0uofPvd2ia0G+Ij194NI6FhKv4YGIIVSdVsKgpuUtM5bNX
V+wIx/qW+770vgA/U8T8X1uTE1k5HFsAAIw/N8S5xr9QgAtLFjJDjb8wL0XZUYRL
+6G0wWFCEIE9nS5jd3zMmaiX0UbpFy/AUCl/awbzYtGAuLaPe/7VCsbf86DJEIy8
Kgs1sG1QKBoCgGetDv+9FmmIE84IyvxPODu9phn0Ej6pWpoG887jrRgENQJjoQcH
dzv+OBt8jEJAc6BKbFmY2RwdWEpNXDBkm0JRov5UanLjv5mXAhEOxHNABvwQhIx8
P52zdgOX7/WdtOOebFxlCDgzf/vW5Bu+E/OFAu4+n+9W1leTRbxNq5phv3KHLhra
RlB/j3b7f4PYX+zCE106gULPBuFuN5yJGz0oNlz3yoBNayEVFnKleA20j9T0K2bn
RemXTDjYA7ZNKRxsTqGTUH10p1dzTOVjUH5sGaC20hhEo8nto41IYOEVZma4Yf+0
p1n6zTJUM1n5Px3Opcy3wP48+Fk7cKcwfhedEIgsEprzTESy5M6pIusOzBzOQiCg
aSvMFU6n0IRFAGEvUXPu0oWHulozDbCvFXkspXj4qUd7MU+6nlfuL3CmPxy0vvWm
GqZ/wPt1XegZo/YmK4HuO7JGDArnvlvtBnb9lg4bGD3C3vHLMvM4MPP5eGCA0Atm
H1bAg9NA4UJu0dtODmo8oixnRJeZ13Zo18NruHduWrK+LyAcxMHScNScJUEXk1/n
3VpKYo1uRQRQt2IWs3Hm85hFJLzCS8u3udVZNee1oEA2LKwybZ7ZFukxuGbODru4
qEbnxEyQPQlNPN2U9BXyuV4IB0WDmxRk2DrOmw0WRG8GWdbQssM8ZlWL1/jsy9u0
9KKHYGkodKSxw3RiEBolCkuVD2IE78WOr8RWl4n+cFOwSKnb6rfDX1y4wxH1Ap2m
vOS+sUeDLxtptcMQ48UAZEzIO7nfRcmgrCzuoIEVxdypFFpGltH4rGwGwBIFnf7T
pXLWEz/ICaaSZtxcoPJuFhVX+IHCDAODddliD0jFMGaZTRfPg8h8ekXbg+a36aGA
JglfHwgKSp7N7n0Ebnc0NaUCyqLyDywR41AI5wcB3pXI2MiWcRQuU/e3ZW9ZE5pb
oBeaM8zwu0sCIDTNqw8o7HWo+WsxaqMK7UzRJ7Sgq4EWKs+J8Cb6eq+Wad1MW8+U
cPx4TWuVdQiaztS8mJm9tzuxe/E+a+p+/PNWVzyAUIpFVZ5P3RjLK8ZjOmf6naK7
atRBB4KwgQ+L29g5+ITX80Wm2sbXPM95/2/HSPtFmlDgLEyp1o3aXrnirtZPXzar
IT5jxvT8twORF5STbylVAkIEZeoVWdYSiY7zP42rJttHO4dJnKfgJ41BUjyiEgl7
xMM1KRhSBRUFGr8WOqfBUibDVdVVKfbq/hT4Zzw9df4etS75eqCoVYiXUB839hsM
2ENeCfOyzQbtOXyOpgn0f7zk3P5HKBn6rwVlYm8CWqi0e+Nyp6iUlnVLgPRKqPlL
kPIM1e5KaQRZC9Bof9CCQwj3c+Bl2KNfEROSH2i4drQEwPdsSFS85p83D1HW8kXp
Jd/AoqqJZ+3OiIX1xFWC2nf9AC+PFfbYD9TPdqKm1bGiQ65BlMf4PyBeZHA9w5Ry
Z50M8E7lqP/+KJVYC0/6f+duRBj7gKg+e3A1qnJ9zy2s5D4L3zPKzecmx0uBK1aY
wV6N694Q1jtgjEkGm23DqMD1JEdAek76RUP6n2syzabD7I+jFjxisWCcSWhMkAM9
2POLFYfsW+ZvGLkOcfVdJ7uMbpNJS5ocqgLKciFMfM9VoUSULJLBraZ5kb9lXruK
3cXr9SBUEkVcFSuHBZi9dxowhl7usknF0yfGl3EA2hKJoBG7oOcDTa1XqOvH0tgX
PrYkDOJ1a4PBYg45GK3VrScCMBWaclknN8W3eR/RQKaOfHyVsRBLM7MEj+pUUCun
wYficLlwfb1pjdPADuSM5vBYKb4B7KbCF+3Wl8qADEkhwAPs5eox0rq9xOyX1dBw
ybu/T9rhvgIW/0WvkF5ewu0sdGYBR8JNObnAqGpQvJskvZdWIeCWprHprtsC4G56
cZnKdgXTxhVTBnQQTvmONuQiL9fs33TV+PkAXnVvW2rpH8/dwUeucg96lXcSp22z
a7CKYze6/6oMbnQ/On3cn8LYHFq8tSWyIxxPpOUTRYrYuDi26fy2+hWyFZtRV1r/
2Tp9GOq/2AxY3RqBmoKRHea3Lp0NYsRokUcwdaf2fvLZF2Jofz8TKMGO/GyhnlTg
wK4Bdn+e7dyI3I3rmtH+5Y7IVqahVBEdRnNo63zP1K/0eEinA80YHqkSGpuEkNKn
fjrU4pzkG4f/Pmsxxk8MwRoqRKmuRUpzEYkuFazZqAo6Q1Q5KfID0xjTJhUCnFD3
el5iu2GjlSX+8ElrpUYRacBN9s8bBe20OqTtyXBcsHGEu4dBSsIVfbKmJsgPSRIC
c4x9Z1iRwadvDrDc2gSXNZaBpU/TXSDlmTfSQG5eYJFvr4bNLL3Sn32vlaRahjXV
mLoPo1Oh9GPXzL6HiVWu2FdMNFxKpjcoSlFGc4pvr7GUh9Yi61v7gqP8/poxH/s1
mbd6vOq7HyCV8t7MzX1iQRnL1inypYiQQTpuV/YSerY69vZi7obv8qdIM5Jr5fTr
iR2l/7C2E98u0u3x2g17/GrKW7W7QC6ttxQkZR0lt5NqMdAX+5LBbqOEUwQMU7tW
0RAewNrOE8s5Bs9uaulGaXsD62MkNewUD9zBQDpWjkXk4CF7HSla8r8xfJ+emfcL
7XvRv50Q7RfbfnSJ0sUeoBg78QSQWKJNJK3+KfHd8ENLSMFa71zj+sLOvoKOBCuU
EhDnkQKIS3zWvX0J7UYohjZSL47KdNKR1iAMpQMRuyzUHnTheEhuGhfD9+TQRIK9
Shdlv1zGVWlODJ5B/VhuEYL5j4SUEA++TNKc8C8sa60EAfPxzzJxerzXRrhbolXu
WMdRzumIFPG5BaHr27nC4nfxbQxO4tFghN2otvzPgGu6P1lFz4Og7zuGkN8hDuls
Pb5R8DFv7xLlne7ofKxEbD22xxZ3r2DYVaKngCk6MjaXw0pCvB+6oR92yDKqwqZq
Psvk2tAYEPFW/GOr5iPC7WgfgPq5LxB0v7WipPDsMnQm8qRXax7rSzKK963kmL7K
Rh8RK6ySYQd130d8RR7tcuzwL+TRplZXRSQrrB4t/imVH0I/ZbXlNm+v3WB89ldL
sZpI80or6FBU/mm4Z6nx9Fq8ldNTJBzWi64p7nbIWF1HEc2TVgjNcWWk5kNN13PJ
bCJfkpXTZhbK1goqlzMGG4wZV7iIcxors8/luyDcoRtfPgQ8aVz2c9xcrbuxrFbX
44g2iH+pTRo9dXwdClNaUbLMlzZNHI99ZpnwGHLPhPn2zjVIafOtLDwomx0Dmnl0
DEeM0tB66GgUOpQgzAVwQUWl2pz9SG6/uENJNt+I6IibjWiiZOBDF7foUUBY3Gc4
0TaDXcB/cf2xAPeRt1z3bo9At7y9iN+33mG540Tf8CqcHh0dkVRr2t6nSU+uvYLN
rFUeXws4mvMw746YKgQlV/Ie+cwo5cjTOthObZwteSeIDhMtySTT/KjcA6TlJL3S
mUSx0+JsJ25lEvNOVmriOIEi2HNxvvGzIVDYbor8Nb/cDTz3TDct5JUf70FiA3L+
DFTlexZB3/t1gzDU8VBKK8yje3xE2Xm9meKyfum89Jg4ub5+ynZhDoxS7dt/cesN
stUxg55L75Ytkb9Th+021RhMdNm5sgDK+4Oe5g7imsR/qaOb1pq4JONuqmp/Cb7R
ERqpQgb6828OZDhozMChdTv95AAVb/EGQn0Mm+o4mRFwC2j0riazWjmb/4JJS0+f
Y/0ikZjCebNxWrJoBtnezL7wIxd40r4o5pH/5hd/c+TYBgyfYKgrGU8irp0+OmEh
RiC8ff4nKFeU8PJfqmvn/nDxqYna9tb2Q7IeDJSVYdLNNaUKlWKYsNAMzM/IeFVk
I1A2DRsa8C5k4/3VwemKOuX6IREwQK0ElDaAmylEiC6KJcECKgl5mqZ+VwldNdvV
II3rFuM5wRPYf0+Q79sD3ZvvIrUk5B+0FM8/eozbyjxG5oV+7dZ5RZjsZAnfYCgl
QsOsNN1M+71OA3rPjhUK6Mq0db7NFZ60zQoK6zfJ8iaK58gD+MbwNmyaMqFWFQCa
OzDbeBpnrB3ZlcW5/aIpg8NE5ZaNLZOxFIo1axv/Gd6PIIMxpVUlt6GpYzbLz0N+
pW64QckpkSjqRVE+WB4cTrCGmo5fHwcW/VjngSkQDcf4SlwGnt0GVSFxJ95HLZZc
1dn4aGMgkNKiJHSfDibw+3ebdTWbpGpze2ZqALdlG0ttb5oecdPLvwmAWBl4xz90
PBA4Tcwv+/3iQzWxW+dXuTY64ZpZwJzn+eMRd4nGWbSJ7Ao+ebx5Qs/jns3ur+Zd
zM33cncUyLvsEVj5BD2ICyaSTS/r2IEHtsSGy9eNy0j5TwrhsMzkP12zKLV3L+kq
+eCtvbmshe8zKlNUCx1xv2k/KHfzCd+1B0WIj6V6g50drk5M2bZMCyiznKf2jXaE
gXjDLjrr1aglgfs05aojSwqcwsk14rVcMO7/28ngPPzbW+mGEgQ6lt2fG/ZNQkEb
l1RKEXDGH6sGu7jQ7IlUchnFOFtaxi+4F+ScQ0QSwNJ5SHgtkBuemd4t9h0kNYD2
8lCArYSSqZR+cEwjNa3Oj/i4Bn/fseH+3rug2e2+XFvvXf9+yl91samyl3p9+QPO
FxJ4wiKowH0j7cliUPmBCi6/eUGqKc1xklup9LS72mmR+5ZApUGKwLw4CHzTZ+tb
d2+W4WdMUvN7sk3HXsEVAMVyyZ9qm8XgbnIzmOvWDreOGUJxdldu3Gn+/SV3zqd4
Lh71zObQ4gYNjzGOIXfxRN6lM1zJFnvDu9aQZq2YPQo1KVEJl9lSBE8acIMWJQwA
CZP9A3oTPx8gwO147tehC/0IQ4Sts0Nk8X/z1fhIYlywoXhkVOaLCnkVTzdZFLB8
Rr+diAr6BTo6G/ShvFNyLiBkmcS16qWXFbOhYook+Admvj14xSlc/N1w+i/2ANpy
LEPSchREAD0XFKRSWgqASvXy221mjkfuR+SRB/2+1qGIUQY1TeuVinBLqM5gblOg
RD9b+y5R3t1Bs0RP4Fs5FlBK1rIgqbigFb0A8rEtHbRIJKCaZp8F77SY5ng0isBX
+fI7xmkjE7UoTKVMGjnk/dNtDK9sRwO6tbw8+VpsTrU8psmfpW/bnlMvZeWKLktT
JG1D2RGAdOfRpNoehLDesAfUthRnZWAFSyQml9CsRBHjQ7373/F7VwdNFEzwtWHv
MKj9l+9gmJkU9uVih1jG4J4W6gHXIcu8jdYJNLASZWET8RDQlz/6jTtRz0VpvEEX
pi5z+TYD1Ee5x6ZmHkyQ6Tt4KY+a63BN7tsPZlVe4vXUAfKY7hRWyCd5CImEu/N4
lFrIWrN9UR+ceMuBrFLTcuV6pfInmeEtF05Ht1OjHsPSHCO6QOmVPg2rJis4Zr79
lFiStPQeRC9ifbnyheMLYbl589R6OqSllfmpSBK6Ztre89LXVWAX1+WzRLMjzz2W
klz6Wiix1pjkJ7xpu9udn1hGXZydGPsl8laea7u99+GSDd6m9P2iJhr6tWk05kdA
BtVYlN3pIC2JEytc+GX4kUhnPok6ERoVINpKD7USmQisz3wiQ0x6NrMVNRgbgy0k
3GwsdxhYLljKvVn2wysGpEbXGhq/GYlDCwh27WQ3HzvD5rocy1zg0cBy6SJmyFga
ug4bAAmKPJOikR6OcdxxULJxZGu34vfn6Vt9VChOl0ZOvJX2NUbItkO4AyyH68sj
k+5J8NhQebIeUDS8QvYlyRzVKN3G+bVJUvpfhTZmXvey/kR/gHiEj8L4D+lbujeQ
GpxnV9nYe2bsdIE92RFrW4VssQb61wupLp9SLfh5WKcEOSZXpLTM94ME7EuRMm9y
D1NU2WlO3pC+kNfUCrAjHb6g3cvQ3tXvbdj/qn816yHKRHu/237VPXOPiiMGi9r2
yOZ/If1MEE9S+sRmUb4GzozxKw/0HzadVx0vFV412g8U8lBFAdcDaUa58Wmycl00
/o7X5mbDqeoxWDt98j8FvzEANkqGzY3UQYdI4cWaOTjgnsZI2BduN9l/It+GYVSv
QOB53ikgAJkgYOxfGE2e5VBUSi+KcueMknUW9nV5my6aspDrxhCynC4QYoIIfoBK
oL2pkD/FQMLce8Lq8ubNO5Oh2xduG3ilvs7P2tpKM5h3Doge6BHenWOHKUFj3ouM
x1KKpjhOmFUpXLwsWaVZ0PDr7X7c+A5YruqpbQvuEoa7M+gMQIru/s/n9aFRfu+T
T4aR4crBybWaalcyJUiLL2O6f8DgU0VQ5dWgQ0Fq0jjxDlMouAuOfyGaYfOwYgK+
wNHV5J+cnlgGCHMT4sJjrqsQWsPCLAlv+xK09+KTdjz0vUsiO1mG5UN0nvXYCQsa
6Gg3HG7as/W3gJ0mBr89sOz5VhftmjvaeiksVF86GuW3BHORit+lpcJo99O06G1q
dx8lVaeoVn3TvatDNa8/Pe+xXpdBP72UIDvQXaEPakQrtWW9JeK6VMt/Z7XBlZPL
ZBRmktlM7CWyvR9yiO8C/Mw7b8ZUwWRoM2M9oS5NclGaNoXAMAge9qRTX0VVmmS9
J8zHSPZKIuykS8BWlKLXvYCWi6doIOk8mzoGxP3sY4tMoXRz+960cfiOtamVB7Ta
vK/KpzN3sM+nvV973c0NLfXMomwRtnT7xLV6emxZ+nvOGdm7eXeE5rckqn8pX54v
ww0rEAH2ixkzqj3zEpNY85u6NcbJnt6JES0gXGGfewQgeCHOPX07+2oM1zyNyBA7
/uYh/GRD1N+OvH0usaa5LmIXe9vVIgfFjZ5b+eeq4Rs2vsFoZW4ndz5j3x3F3Imj
xFxlE9RspyAyvh3na+1jc2RMxPIipwkV6YQQv9/+6FkErm1AMqal0lFshZCkV3gt
adZjWUC7JP1qi0+kfi1SNBgJ8z+zkOzwJ7sHbIYVAq9JRAtXRNetVa+DPSvo7hf7
kL+8KzhQGyKYQyT8bibZlggPqPWpx1qKgnmVnWvi2GRT4tb2TX13wohWXjkJQKxr
aR7Afk/CkbVvU2VJUO65OMDFS8ZWlW7bjom1vQZa1cm1ekEs7Zc6C7Dc6YddPJwC
jisVzkccm5BTvM5GVKm9/8DThTR/GSTPVJn4H6DGzZUjnj8XrpEEXFJXKf6w85pV
dpQFoMzyOEo4tPNecBjAt8u2mf9xiJZQlDEJ67SsbOTrB+Pz5RmQ2cBNN4VtIKgq
Ebj+Srqm5Eepd9O4exXJPUsiwpgNPHHrVm+/3yObSSp6nmp3TZG61zejOA+FZSBQ
2s1MxcRpE7o974ytDrpFt0n/MKX0xy++I1I7PrItySjZA9fVNgYjix17XBMTqywn
/bsLw35fKvR7T6yEPc3SNyOQpXd152f6zf+l1jQwsTw2EJtucnG0UWI3kIp0KClO
BwNLUTMkBKpgDAlhyGmI/5WiwAsmq895QlhdLkDRGtsKtt7T4vrcFfJnryiOGNW8
46Keajxp7Y6HDesRh+n9sLiW4X+dExvQYd0XxzTZVaQTSMD+/3FLuAD60gtfnefO
kWgSRBWhz/SQnj8qaCte2UHrxlPIbzAbzF5gMQUlGug35tYaeuQvORVEPZZiwQn2
F/MlX4SaCGzNK/tl+41Qd9i4udB2mjwt+U1PVKPI8x43c1WLL6jefoeOTDMJYrWQ
PABdlPDFxwFnQ9X4FX083TLaoaUkOSKQACXT0xSeWgpEflLuGQO7Ttvfs4QrIEbE
dEtj87qT8NdLqBvB+XjGePOSYwjJvj9YcloaJPTF4iYWEX38fgD17oUPNK0BTiSk
ftkbwYi/jl1pe3KkVWYoQDmGKJXCTP1J7uPPrEJbi98uBUKuokJDEZ7NdE0B9bL2
GKeyMfn8J5jqdBaG+EfSk7cRlNUEgTt0vtiKWvPfWDkQ50LEYlLHEkWcz7bq6OBa
Tyzt0U8OKz0l9kj6e/Tk4i33q1On+gkqUqRlR2VWqW8XzFEDYuEhORqtZNzOXpdZ
HjqFOEW68KvpJkaBdY7gmZdo6WZx9IJqNw/XA28YhFgWl3S3x2Wt6b3ONPIIOryu
c0atEeGHnTmVd5K5mhhwVJXlitnG3PxW1/KCHqRkaTnwS4wgWg6wqfh22l0z0oAj
HQfY6Yw1xyv1riYJdtVrTRY1M5IFBV1DoF5fkbVlUVI+NzLc/2tZKCrmzroL3XF7
DCIIw7vV8tD4DntrvOb0ingWtuvCYntV+dYeNdcFiA8ywPzTMdyAImXLLrRx5WIh
x3hWCSlA2phyDf8V1uDkUf648SVDTugEB/Kipjx4NXMP30n3v0zt6cXJliUAUKSu
Tka3VlPqqTIG2ZE++EuhaVf8LZmnzk7vro7MXtosgP3KJrB/UDOFbSibvexm41XZ
u+X7i+97ofWUMhuoh74g1Ush4O3QwYKLgRyRyMPYdnHQCh04sWAwiifPp9XU48P6
kdyl/7BgYA3LECSJbYeJsAYQX4OZxZc1slwnoZoB9rIQDMgQLKq7hhVURe+eACe/
DdpoDsdKqUIJjn9BEBmLJAUFrpozRoTUyrn9Rm8zGgYqjtd6vwficRGylRJ73xaE
HXa8wex8M26930e3+5x2Y9liBV4V4+X5eDaHG5xDeNJIogyHBefehBnwsy4YoAs6
p2bNwagU71P60rPyVxkxu5fSz12Iaup7dCbqIDLJ1z1Smgc7gpOCpe8VqPV+/0mf
yaKsuM+uRlNnNGHTjrXyMiz03mfU7PzMTHt/SvgZDgf/FXMW6e0QpcuKcjb+4q9j
QJU+h4tZHHX9S5CtsvbBF3IdHMrA7XMPqCwda1kYZiy2NsJsrB8nCA4LfvTZLcjQ
vhsZMNv4/fVh8V19YezowesmE0O16tFRfkYsg10aiABL02tfYU1hG7OfHKylPvnX
ly66x3PGcHIolajuAEN2Lnrz0Kb5FNByowuqrFm602it3mqurgjoEsfZvmpUhJL1
FEsaueGWMxdLR4JcxqgHHylc8qW4f0TSLlp2+WfZqa9PborPmYloKh/2Y/+PKek1
AHjzN2kKSLX9Dy02EqPnIfMFOs1pOy4ZSQLO/PIurX2kD50xQsUbuAXAEReY820i
sBe+Y/1Uz/igzl6iQhEpTDoOBHiAykJ8Bi9HPLkDVLW2ozf9zX03AzuTkltCZFyu
Ol69FJY2aZa0dQg4tfZjlM9hbvnDndAS+n9SYTGTEHkvLLRidHzG8kK8YZeNVqOM
1DnB7VT58/ezi0I3pOjGpH182XQBoOPitj8bfIVnCTxdZ27V0j2jGEybPMxSUHk2
eNn08MoWo1Qvy3lvXyYy2vtAxUMHb3ojbIhkDd/1N+iRh/rM55ByMqi3+2UlfSY/
tPiP6BPqB842wdUo3gtZcrNeNaGvGq7LGmWP4rtdApf/0iMogjBOwDmVqXpLKTGD
L6urT5u1lIgFf8PEHqGYr5HmL/bxuDF00Mr30mNHBWyXEpsmqfYewYso3bs9/1A4
4XMZkhHlfntA5gVZiLhJ2sMCHz/7Ji0+tlx2zpnSQQgJ/6QO3bZgOiFUiazOFn35
T/EJ4aDZlPiW916OOqUJbqEItSYU4ZrH/AqX1QMXPHFU9g+ji7VbM6/NIQY5c6pD
jBwKnFv/b+HyhFrlL+hyEavNRKFlpJCMy1cnDcWejlZkhhspeHx2B+5nAG5/7yej
v0MoAv8sBkHpt38atxjaEvAnI9Lkgv5uFQIVn6NEPRViWc6v+3wHG93aWdgTxSK6
00pTX2fvBvWOV0Lkf7RkI5+NZ+MCgRrVDz4BBs0dhKULAQN6RI9qaADjNP6Q1cjG
tzi4I0l6glx1ezsbf/FIPwQfyq0jVaN5v8YDXmaGbOcrxZVRCSkMXV1cCBnpQpQ9
6ftdm+jyGUEYoXrKRMh2N96MpErhNOjOIid/p97MtUnxdTGtHv5LLgG4bPtsdya3
YWZuKOG8ECUJC2a4T4AqvQD9TCTZ2QQqfPhlF3kRxD2szpf4KoX8Kdyv4/azqh1/
Z1OHVuqTI/TsW4PJalhwnBvZ3N2vYqfJDlRXB6qxT8Rcu3hrQ1goBDOfLmEQtMXV
qWP+EUJi8yAYRFOr6Gl0WP0VRez3GB7Vzb7gvaP2AkBwPNTH0/DI4O66EL43uBeg
EZwLj+sPy6lcbCJYeFRPU6wGH00pDso5f0SKGeMIhnMQOpykqpGWSH6AeLjqH9uO
+WWwEVLCrJTGoYvJwoFIxWnhsnMO4UdfjGmH5t+xYJxYvBYUI3RcG4k7e//RbDFd
n0VbaIzCLCKce9C509g+uqm1GtPeDQYiyp5jfpSj01cceWDbAOhN+W+ZwYw/tZAh
j7irfwkgXhW/Y87gh77pwvfSr7fj6ihhAzD8tRnQETfSmmOCD5SuLrHGuCSFHgOj
Gpr+ApSeepKThLMOOneaKpy+Qq/7HLHqj5zrOr0siezya0R91EhDY64v3fjYKbTd
1ondUDE+am5RU5IM2C16COtULdokUwZbLj+uzGgOsNMoNUw2e3MtIIyHJh7ia1LK
0vMjMicRLbn7Bnx0RdbPuAddLEacbWa/i9rkM27JrtPUZq4aR7aTimY/kvLGMx1E
OmOWVBhOyVfzBo3JyDRbcQq4a5eiiWrD8w/6SwjCdo/xwkHhqkckEsE3RWil8IsA
j2Z4BnLXuoknAcpkn7u9nRKxjw+S/B9kxBjjhtt9w2KgGF+PxDPp/U9s4L0/Gu7W
B5wyxbL0yZF2IIKRoa9Mqn7/o7FUx8NBIIBJfleJVyyG77VJ1eDPhvFGvogU/qG/
p4+nlfL5tLjUJweNHsZqBkmpJAi+khD0widpxjoy54H3lmXpFgwHiVq0l87BusDw
tRJlfK/q6FTDoElxkcBcqOmd1A5TStJAcA3UQOkFjLjVHvGfFpmELto+4mo2TpGF
h8m4aJDRgmNrw7aKpD3ZUB+87tneoPii+3q5upQXpasanPChaHULBIw/Nj0DkzMO
OQbMMb0ERVkwhYBL9416iNeBQcWJNxHxx9ZGPrQa7Qxs23UHKqsSGadXtAa1xnyl
x04EsD/01eEjzfMgW5fFQXg06N2XoLUJxkMFX9AakpMORU69GxUwmdkFCHhC5T9/
VTUPKns1DB35n7CGHhfY1YlP5fPrd4vRXKVO5Op6lLhJb1dXHOM02eLIdrzwBsJa
SObagRK9bQECCzcHglLZmwslM6s8SdQ8+HEqeOAB5kvjBVdcSKFAHXnY7awNH3hj
cLDkR0Ra/GTST4JU5u6BTx4soSJaWqMst0nyVzXiYZaQnFcx/BBGKXAqg6XpVyVC
C4pq9ut20gMjNmE1wLp3lQg0U10I8Rd33u5kjBLrtHhZa/IzFoRkDl+zaO+6hP7A
nzabJSJSivFKEyWqHkiMyrp40NA9Xi1fT3jfhNZoR2sOwTubmm9LRRxsBESIlHej
PdnsZf4Si/slqNvYwW6qKlqBNV2uY6PM3UUzektzMz/MpFJUvF0MbKEgau/NL4+N
9JCw/pWCgt42CXRsRQK9O4s7w/GuERXLUxlEr9Fna67ZYxTOqbltZ77+zx0Lc0aq
VlRB1dV8hLTwiRfZGhLH9y44XoWpTIwIl8RMlgNSNb7M290MkzTT1XjTw3spham8
Ys2Xgb3wa6nPfgVnrvEZMJSCsAEWwtcB8dC/qSw+L/S5Txm+Yn/ZYC1bVuz1ebmi
cXth83/lhR3ieYJu2HWGk6PJbRZ+4SiOtfWS99TvSq94fOwbb5valE233K6aYala
cAiqEqC7PaP5ySSVHHECqQzRDeqhIPMGhfXrcmMOszH1wmCthu81OpQNQ4p2Go4j
k6o+CuYoIR7harbJRZzBq7YJIvZ2KJT+a3qkG/wh1nGV4LClmNqqq+BjGfR2Izz5
AzjTa1XpoCQ/pSSQZyC1rF406J4svuENj0eebL6T0LrRT7Y33+7hK4+C0yU0ITQC
BnTaKRrp7LItFVdS855GhMOiWpVGWbNE8GZmF4F7AfROF10HGNREHf+JkNeodk5e
esaQXuMgwssuILuJ+pEQb5lpHTtK7ybMpNHCdrNj3kw2TWH9NAeZI1TuFK3n/t9r
ph0Hvv1R5oInwdpS7ewMyRzhDt4Wwpt8+vNd/hS3YYcTuQt3zLpX+491xHU8t9st
ejnlnRBMKn1SLU/u3PXsnZVQlrS+to0L08yqojklhebtcJhu6lloNiJtVuaDwffs
TDOGN8b4klaKymfw4pm8ptCRJQgO5EOczhy2RIcXhim6ynBnDbz8b1TaicVsjtPq
qjyBFwrE3qYyHh5clYV2s3Ztrrlkxxv2HOn2G7YFOiwZmWGkA6hJF53QE5yph+nl
QzqJrhydjP5NlfTv73LnSH4/pYIc0+yLDrwRlTUoHmyQlv7IA/X4vmMmxcgf25hB
5E4Lpvw9ZpD+xRxEZiriHpx8mamvxmFYbap5tYDikoYyCOHnnzPWtEuTxEcqhVfa
OHVUxD8LOu0VZ6KBFPO4rtadEzB92x21kVKbh2NjuLwSf3f1KHz2VcsakyiFhAns
Vu11mvgvY9ap5Ov5gMwqXv89dy1st4KHw4nimI+Cq0B0fvzdG+VAEeCf/vGnm50+
8+PtGXZbwM6aHdudyXxHsFsGXQpT+nCZp+FPoqaUixcFw1/ZwYhFBI75fc2CQJl7
2X8xAiwy6J5z+QRXCIV6fwHnMYFajg7Fikffoc7n1bbgruO7MxpS08irrlzQ4hkM
D9/OJcRlw3AWxRZT8jbG/4fTLYlI2bMaT+uR6MwpOF+DE2Q33f5IORF1LBHO4Xr8
zx4lMaf5i4HbMXFOf9o1GrZxQT0q8mVKGOMfTqcS8vIqkAkGXUTa9JLq7QLfe8+q
AacOpBoToheeeICrA4FyL3VYgHk8QFLTzYze+QbXrEjUPVfmEV+wCIor88lkKsE8
JPF9OCPy0PBe1qAImEpkItxcJSYWQxFOCdopagdmBFI5kXbJWP5Ciz/B0bM741yT
rBEYFiZaevyJ1pARtpuI1QENPs8asoCNP4o3HNNzjXmZxcx1rXyMeJM1Q7f8uk92
RAshKhAa0vCCid1c+8hct5ku90xKOXwSVHNtU/e3qZjckpB9rH8uHkqElgaUantd
aietwsAgisrw4x+xaLuP+9Yqv0/zTkp5pAusdr34Bx4ndlXijJ25OgBYZIlYl4aV
deCBxuuvws2O1vPhWjzlLOxD5RtW5YFTOdFLXO64bLIPKh2XwYeTQhzSrnrDPMFS
g4np8d1wo+UZAN79upC0X4cxzY62W4JHFPzgKsX9dGDO/1O/FMYJdh6sReAqtSlX
MxpeeDY+hu+3lWlv9UQdu2uY1NraMEEy7CUEpBPDtLS0b//dGooiyV7jbdNDGBJN
mSiiHxLNBqfWbfjSAT8t4ELEv+o4+QkF1/YHFlS8j5siMn6pqgtkbZv8KX3U2qCI
NEY6hpblzCE/a8iO41CVb4rJJIegtr+UTrXWqISWfJlzOXioVJx/EVI3MGQlQRtw
A9a4A2W9M2IykbLGy9ZaeIG8qN4NJmypjzE6WVLzC/xIHODC/KN3Zm3FG1ULPzH5
mNkTbiLuTPobTNeImF3+es5itX6oUGrJJN9bSbIFitEaKSH0p1IES1L7I0FsvFi3
QUeOALS4RVUfghb3dA79poeUvAHPSOhoyfRm9LURQwp0BPS8hZUJHTHEX+cvDQEH
MoaNaGEAEMJtOF9vYa3oxZzQ9GKzLrFpAonVASubcYcEIyr3Z3FjjnJkLYRnbywi
N4qmjDNGFyFtlh4MoRAl+6/osKp8P62VU3puvqLcl+MzQj6Np6hAmBmqA3TYQtJ/
0zK/emyfUJOLhmk+FHqHynqWPtmM3E0NupY3rimLpSP2NCavdU9ei/YfM0yffLZG
oH4MM+nps4JjWFqZa2P6Ei+cIVPPHMZP8DGJ33obcshzzeMyASMM7GUO1nj2/piz
M9Xr1/ED5HguY2Wwtfxi4IbGRNpdqHs+43J4peWmzaMHeP6RpEvlLbFiz7cPT4Lr
jyVGh5a2KllzQ/61kaX96ShHtQS3ygyvYc9s/F0Al0DkT2MWRNHb2xdRewnXv4XR
HPlrreVVHdB21q9fRLIFlXeZst1sHyNU5aqa6pdrEOIB9fIUpIpXKOT6ef/rM513
4XKWj1K5Cy4HD032FptbPFqx+eqmP2Lxp625DcxQr6SyOJ/JA0bIzmGTBQkcy26i
3SPJLtGfSryIdghuc2xtP6gspkEDNu4D1rGzbApHjfsuQ1+kbPgjTsg24aj/YsyD
O5dkEGMh2SisoFD6LqqVuCKqFwfCUDECyqref174KbStFmXFbi6WZ7qdsvs+SUbP
7xntg1FH6xR4klOFj3O8oQ3VICMRDgbtY0byxWXQRpYp+DTKmWtpBXxuNsItXAam
hZXY0K/KKpv1Wvs5IYlc3w8Devj5ql5K8TTmYrcuokUwYxcDtK30IZnOMZ5LHU8L
RBQsIay/L3weSSutQbN6A+m2ahoff2FE2yxrclh9soIHJ+NwDkoPp7vAXwA0E99z
T+SkE0vCvI9K2tGVXaiGKGGwiKW1OOITP32bsk7uGMI2yrRgwtjxrrBul3ROliYJ
wBTIDPxVPXJXdlT5QkyWF3j/2ut7NKp1BHi8og4Ze5txwstPLIb1bBxD2fAP4km9
NC7D+1171sfBszarkujnBcj4FszV7ylu8+4T1ix0NpsWh2HnYwajKiqxMAcoiFU8
xtLWs02akvvTVLqxRmNXkHZaxyqNRLMoGUl7vvQoyzdw/tISE1gWDKIu6T1Ggf6D
i+9rbYBYWo9A0oTLswGWM6volMnwOVDUKBe1JsSkAzuuBwZeYd0NALIjbHt7MlaA
FB5mjga4iTo4VonwZrjZoUQ3Xd1juLuXJAQvJBYYKigyFa4uryjplrDzN2mOug83
AC+TW/ROS/AOifHgY4KZ7zQ0UBUA0kj1ZuGl9VWySXAvT1yV8znpKLaSdSLXvATq
egy/UAi0v+mYIc+g5ujTL0a3uqkAp/yFnsnEk5+SmpcVXihFfLW++5jqmeaR//x5
pBZRDvxMKOxLXYk6vWODJUMwWlrMlssFt5Xrji20gfdM5iZbudZFhTRaBrUE5h1M
DG8tyLsziMrc+kBD1DerIpnJuTaMAHUxsP7aDNtdgWdyP1R0Grumb3PFeZn50gen
IJraqHTX1ZS/xVXEmQBJOpCB3Aoy39zz28L5Bglb438sf6s91AnQPqyiFHe3AFqo
8E3fXT+kCJqLU/1yLnMVJzE/58R81jJKiZ5unhcmCwzQqeHlIEf4FKJpr1x0y84C
8av0V5CSv7MqweGWwZ75ISdhJ54OsdxLiDpJBQizhRWwHnJ5Oio5bbryFr1oFZ+m
pi+9qhv3oEXbfLtwF0TtQB8Wwc448Zh76jsfSmID7aA9aLHKW8FeY1bqnYVEqfWw
sEK8QAyMeSLoT6ylAzPBT5J3/TdAIqsaDssnXLCpOaYZbaZkVC8WQlZN+ZYLnWYQ
vzhZvpOgjI8vWle9oejTXTGXpz5gxOsSB5wHSukR00sb+UOjI+2XypYrAIq75Ry8
SRCFQOkhSy88VmUnBMYu9Tw1UkgjQ+EJQk/M8Nj6+GdhIrNF0mE8+Wslp2HgJjAm
iOWpRaQvq+SwHootD0L7tQ8CoqXwLAGvvT6w17rIemY/5LaKA0Yw3kKHgPRZy8NJ
GjMPLAr7Grr82SmY6pQHqrHJdycQ9kr9+qIeFOVexRuzSA5Ec0cg64T9pjWg0oLr
ahIqOz36l0Fwe4sTaQhYyz0f4vksxAty3lnS/g7uyt/gGc5Gkp1+S6DFKdIul+Oc
vWHyhDvf0sdiRHCcaG0EkCbsSPD4EVVaSVr5+unmqXV8IsDwo65/+kPGShNTS+KL
MvZzfhEnWK2M1QuMO/yMEAKMRKcAZoJlrTktn3PoAhF4Me7zqcnuc3Qmoe83KM4i
Txkfmh9VjYvuq0GbqVsOz5B2QoYCTckDFP7ris3IjOXRjekZmNlfiRfBwohXntKc
BzimwDYpZhcBTtGOhTjyNiRk0JjGdQStB/3VDDmk6IOP3uNG2RwrR/5NubE9Gg2+
YeJ6MSmOo+XOeE3GPoVnXeXSn42m9JH5ue3KLHUFq67BDdLmxX4vs2l/WWwZbndQ
2XlARlBwDiUXTpq20U55AI6IRVMRf3RJxX8W7W2txofhUPX+yER5OAfrOmd4bqRb
ifomNWxdhWFpAxbQsyp7R1LTQcAFxERUku7cbCxngugQjFeLOSS0xHHT8sQB9Sve
Ss/JMpe0f/MTVSkmzpPDLiR4XxBUAyHEVzMlvMoQ2cTOrLHaSJpiCxHJVlGo2UPz
+I/zRsDL8P1VV+MICOeabMStDbn+3n7GKtBIKV0IJ1584CI2tr7qmZFgA7Y5281f
8r3ZACQ78jBcl22VgHiF+Jo1tB5tw/EzRnT33SiROBxqVKaAauNWloe4nlkIBfZX
4guUtIUHkmCTwcPD5bKnmhcT3rfvZPxGrCcR3b4mpwx1RncLxh77wpGBeeVrQGHX
Dq+uyhIHGV0KuNfwTX9CtQM2BIQcjEnFosxAUQWhK5IOlvLmwMmX9iHGzeh+188F
h0Vq9J4shBc7QQy9Kt8j4VRsb9oPQ4eZaf+zvIfYlXTtSGGz7GGNBERGGqgpsWsy
39tAKdh8iPKAN9it8rejwr3qY/zZ9YJ5o2ZydZph6ipO5nEdFKmgEWY2ilFi1E8q
JcfF2kTmGp8+UJU6bwKwJ6pSoJ7UYaUoK4MUxAjxL33w/0ll47istvgeL2343X7m
Ihxz414F+YvtQioiu5lXdON1Kl+wFVPO6xtIRe2VafuePFoOk9HtX2TOmvdAG3KA
bdyhzkR79qRcWIfY1FJozOKVBrwEmxjWANdy6nVI5wq0cY2AjQcNVF9mYNicnGhz
KaBw4CX6YLzTbLdD9KGd8KHIybFfbbqTsZp9ol+mMEXmjL35ksJL89e44z6PZ9fo
jaCpeOz8/Ju+T7tkeztvJzYq+K+xbk7deeqSfUQp8xlDpipRB9fShViu1gKkCMg/
1tvtCCeFCVny2Y9Y7ugnLKRWeY4jX+cyoGZYGXO5Niy2HXyoo0Z2yEZKJqtIm2P+
BtopWwRP80XMak5DRvvxGLTGffyIH2GFpmAzT0iUB6MyeI4LLE5hif+YbjGHc1eu
bzkkhIis63xrHVR5GCvZH7mQg/W1Ht2+7hEBWJDc1mIF8E80A7Re0V6QsqLYO950
WRh5QgAVWi6gaPC9m/9cKxZjThR8Yjevv+Ra4IiZx49OMAZYrtg1vws76ly2nd5a
UmVULQy74zvWbOjvE80+n9yFLpLvyIIGcrGrKM1TB6c584I+k3ssTgypTKtuQsdK
8lWk5//k4jCX50YoaPO84H6lOEMjfT6dxoLWfwebR6GQTES0C/Khfw+O36MC5moz
tOl2c9oiD1S9sxPDqqD3xgsB5LbGjtUwb4M03SX4XAP9y/ApdvB7Soi6vSfL+Isz
Ui16JIU5IGsdvcds1HGCwXpIzzb+LgXbyxjSMfqcQ30MaN44DPPswnuhGLSaMCxT
p2P63KPM6rICxmgxvOB/bPbBUlxDC15grlOseyrbAhFm7udFm0ogZJLN4+6slxjY
i8y1IuGP+Rx5E3XrU47BhA+v+QboZ4pWM0Yuk9zJr73xuXkKvAqNv7IOYkJ/RIA2
PgRa/P8oOnAt003SQMl202RgzFRnuTbvtT/OBPofuAn2hzC+TrvJSGSFK4NiFAWa
mOM1MTtLpY1kbdfC3zicIYbZYO5xAiKRgmpqwVQ3bQ5bfunIX3F4ep1ES0TuCna6
DM24PxQfPiXo2s895euLuDFzLMRpXF5R/CfTgiCfd08trZWZl9VbujMIzM+4v4bw
s+ICcRPuHmRGvY6OVV8RTz1jseKui9NOb/ls+WdaK2/30rA2ajkhObTqwk94Wtqe
lhmf49gQrrUHg7r3yo5apmi5Nwno6bz5ELDCC9Yfc1srqLPo84y07e6oH7ZVyFov
X+HYWml+dzZwm0pBGm3G6AiBdCvvJwZmtAOMkg9ECIDtPA49oRSkHziuVBE6gP4A
0bxVCahP/1rI0VGacJNAqydAUcJviPQgvO6V0rfxbGOwKOhjMCbHTr0sSessNwtF
l1So+sBOBble7mhnnQFF4/fcEZntSxHOdpCS62bRNzdsTtLAYIoXbnh7wrNjfxuA
6t88w71uRLRlYT+HXobTIOu3PpOZFh+b1WUyaqwiJTlBhTO8DeTDWCPsl+pTovhF
sNfHSyVNAcCsIrsl6QijG/9kZ3Feg3K45SsS44A/TuyHtQU0+MXmuxRmt+Wl/rTp
LXTpfeP9JUnfs9jdd4yb6zZWwtJp9I2DZF+mFrHvLzSjLvw6LYYNrLDVe9yTgOJG
bReHWupq9UFQKZF+g8J5+BQiQtKJVQuZUOrzzgRLJN4DjCgilnAztrnoSY7drTEv
EiJA7Efva7dgixfIwutnMvRMUFuCGpJbAesdC55h1VueT/GVVUIGd0/YLXFJvfgQ
2B3vxHoHzl6rShAP3H3eQVIzhi1R9FMu6AUDs/D5m/zYh1seGRmdrlg3vgble1fE
FIIaqwUbWIO1IpsmYEKi8FvkX4aonQGily3qOnWDGdMRmimfRmw4/arpnuwAnxUI
ydSG80sl3Kdi2zVSo4IysQ5TE+wZe4TK39qZUSm+kL3HucjcUjV6g+pgQ2acCLUA
f0Z9LMJ0RR8OsrPpK6Nqr6XJTfQrI2LwNRf+gXeq4EWoy7uNarEMUrDQs+C7a7qA
KHoAHGaGpZlzp2kWYini6k8zI9UVccxRBfviokdZfE7SIs+92ZcHyg9tlyXq0Aqq
ePZH3SO1Zcypkg0DtT6WDKqCNRCA2a82h8Kt1ByoAlUaYBWR6X2XC3YOGhSfpdgl
74GaNcDSlf7eImPuKGdojACEvpITG1xWaGWzBPMq9q3yndQiVrrkitkOg1GBtU7/
YEPIiq8ZgHMnllu2d7uAvpktUG1QUXJUfd4sgH8rDfUxLujrwZOoFyBZ2fS8YoQD
0F0mWdhDt+8eW7TycRT+saITGx/4erMut5lW5HGq7KG6+rtN1xTWw/IqtL7P8UYr
wTVmJTuyMrGvHmz1LFt3jNXqAS6RMer+p5/1/L4+JZr2FAK8RQb6jP/Pw1O1GZvU
u9+HGEf1YuJ5RrruqPu6R3xVHoPxj0FoHLpaPlxjjgWichKcBXD4Oncm8MlLbgAe
5zoY5R2+7L6Gpx0R4HGwZcO5ZVVdsQ1CJEg52vD6neuLcXMiOdxXDVpfUljJO17z
PddbGNaIvF9yHzbheVP/NeTT1Hw69tTzetku7jp2XExdc/lkx3r4PAaoiXRMc5rs
4VEJddXdZgBcJRMARBjRtAofMp1EtvQj8INboIG1GAtdMXHwfPkMDUn89SY4+Vuv
xhatY+eUWBP16xLpUQnhtI2GmgJdhOIng0MOetPJW6N8y0IrCu/s85diVXDPcFb4
lNsaRkQuwLGEJ1pILs9lm6I3KJ7K8zXEoXd18l+mg7MoQ7/4nycujS84vfXT7I07
lhZ+QXYgrJKrPMEYh037tZuR1HvRl8kDDM7o2rcuBApn+whYBNI7NwLKJ2D4crJu
NxPIspfFT8lAURBnD+bWdDemgjkg8bd07wPGHg+7a0zX8hM/GQ3syNC+G1khSxPI
W9CU/5570p6mFG4a/2Js3pKyIjSayCG1lxtC4GOan+XAjoC9RIehHXmj1wuBRZRp
NwLwA7t0g8/MwI9xMfhvTsvthQ1B4obo3EEalzEf899+QKcL14FoEDc1EyZYvKEn
SXvBU+KjKt3+zaS9WF36f0AXIyZDd8/NmpsiLqA5VfDX+v7cWVpf+Z+fcU9vD61G
jILDgyoFmoEJAfjokUHMqdR46FVGyJz60npKj4laYS78NBHxuwaRhvit41y6+VX5
1XVQp0soD3xekOVchM0DVc9NtxU903wAI737U3OKiJVhQ99B5T3wQxtlb0aCwPZs
OJrV9TP8q4XuefnUMJaH7GrYOWyERsoegqSVAmhivl2lj4BkQdFLlcT8muEIXmTE
0xB93GHW+xlVhFBTuN0I3rQ/TlFjM4wS7p3WGiw0aS8HH/lXVOmA45Lyb1CnuWy8
X15FCT65G+bqaHu4/oVqhQrERhAipHcLPba0N5jwirZ1Z67cGrj9nYJopQTXLBP1
WPpNlcwB3dsqAs65oWcvRpLfVAGPEDaDYqFFdjHbz4suSnsXxomdJaOXEAgOVH1m
drXHQoB4ApgTjHSiFj9ttInR7Y4/xlaWrkPfWNv8VW7z2vh/MddtU5NpObnIlo/U
6v7PC9r2NhH+n9Uu0zP2lYixlYUXsm5Ib1jF02TDHkSue8uPouF2Fr5HDU46SlhY
GtxHjhSoyTTqIdVa2Zqf6JdMw8G1BChRPY/qDbhRiS5/J2Tf1XXoUuUXTw1nFynn
+uVcxF1h0FXNwqtoyHP8bdWJfdPyV1/hKvV7QDRvLjCQ7a8OjpH0xmR203MBVmmo
N07+gPbpl0GvTzJG+NUolHkzNI3OgSQNcak38xRWbwq6Vn4rOMfxr1JVGQds8Bia
D2rT++A38dh6wUyZwx21mHIKzDTv/fzI5/G4yt1Plcu4+feIs2cGdUQoM1sHJqIT
JhH4WtxjldoiksqdZXGntI2Te8dcVIpCsxuiOd66wuv9BTzjQULMPL2jb0eM6RXI
RPYv3XEIWZYyjtmCoE3wK4bc8fU3AE+ONJL7yICvji7zSTz7D6UjR3lk9hqGFghf
+Nqfz/NXAXowiTj0wVCqz6UuymYESmwTY7p+5Q4JjB3Trcz42HKstw7fmIFpVA3D
C47VZLcX0zRZgVbjPftxDFLIRtY4sjqyEcx6lJH+eHnBktYaom4XGsByqK6zg01j
UJiD+LBZRvI36fHeiAQIzvmvkG5HqgyRNUS945TLr1LThpdxtFBhS7iOYxOS3ubV
3Bq/BJDo8o3w1i0E+tvDjXjhI8rum9oYJDX7cyZtjRHF6PfaVFazqHNGMV8ul1ja
GRbjAg6O0zeQbQDLA7PepjKKovb6zjBFdOCawJFD0prKqu1KVQn5jLb601ZZMHRT
T/g3sNYvy93rpUtZNbrjIOrm9DlNfqQbNTJxcFLvqEkiaPDelGD32BK7xC9kspDl
QFVn846OMOMWIPEf9ZOcJt4hRqucSh6yRY+pb9RoTuO5mjJQA1naVwdrZxEIVe9N
W83p9vdkyqOtk7kUTfglyhJs16QQB17bgZaxpLH5MriXsW6OiR61vO02d/Ot1JLY
3O6yx4z075AnVQIYu5/vxDyyQ0L2RaUNpuKP0J4cYTmKIQbtG+ldR838v0ATi33r
HEI1EB7iUb5ciaOpQNpR0winj7ZKckbqFtLno2JhSt+FuOMrn4U42OxsnUWfIPia
MwISXjD4E69ya6YezKpvJjNdBxyoARjLZttZ4tg32aPwf6jQtofKZ1mo10E0rjp6
nzwqkfER5UwlH47aiNOaahSPNQUe4TF26XIkyHASKgdd7veA85VLnnWedW0hC4ZZ
axV7bTBGVfM+OBS+AiN8BYEVNaRorOz9cALVgUNPla62Q/SvfNms1Ff9EyNzSR9X
i2q4Yi5UXoAaP9/rzI9elBvCsNYwduH7mzWCogO9Gb6g/YiDJ3S57ysJaJY4SLP0
bG+ag9RBqdZZWEHmcflMxzu4lpdbDd6zI8H0MMsmw+uj4lCe8KwW0BPtlzv4AoFD
gJu9SvHggQivR/MtGqMu2DS16m2n7WJocfLCKHkboumHwxThY6D7YA8zYgVV3WSw
YYepauKovPNClFa3HPMpVn8Wxml4En2Dg1OTH2NocF0j8XcJWtvizviFOqzRPvhO
4/gvq9wpGKdOZnt2Cux27dTWSuPOzq5u3RNm3SvjE+lqNNVhTSSGC5nHbgiAchIF
TMp6jO46posOPrNUkHnpJYSlxPBw0hDGe25au40Ki7800GlOqO7UaSDXu+U9kHCW
mcr5AD70LkHfwD9e7L7rsQXnafGYv1S3V4Y0BCDZMXh1XidBqWRFkGMkNLo/PJoS
Qz8PZVWH2TE++hboo8cJ99PsDHEW7T9u2tPhWgrRKcuW25A0Nk+D45gDNQ1MLrQZ
oxDmFAWaJN0+V1rPP9M8AXNWnN3IU5pMUuMdTdmkb4HvFCk+6G+8MtnN475Vdfqm
TqWNqi24LtssHfZbRanS//jHcUVe5BfbcmRnIDbbXfGMujxIF829iIvVv7WI3ViL
2bTL6EsupPa+MrdQOqve0rXToi3KhjyC8LL5K5u6OE6iW3a6i2bAHsWRH6dNSCnP
7hXcOzvQpcUCe9k1ph3Sm5FN5i+oAVVVx3boVc889CZvqcAopc0E61h0KWEvy5Z1
SVYrdcQOsfI8JN7gepO/9aYvDMjBp+v3ydBf3JjRF5ukZto0j4xsoG3WHo8IP79L
SdYkFNtYUCyfGArCqK1B2taC45uZQ2e82WWonwyHsFor9lcVn4FB1fyl/hO7JBBO
0FAaTDzBmfc6ti41GNzwYVgM7ETxn5Ar+UCTaqhvKxAWtMcbEOnvMDee2e8wnp/1
EBlDTljkBM3V07Dqk+NNq7kBmibkfGCWLnu+GrqxjhGEn6Ai8oDuypQuEvgjameA
OR0wFzDah+iM0XJoZH2aNEICECUd+TOjXKI0t57G153HX8+hHnqeC2xkVuQ2mnuH
EyDLhV+szuwzgxnfPzIx8zJKkVJDwb6437h+eQMuSuADGMmYqChXQanoagqNmnec
J5500tOHJC/gvArkMvL9nr4B+I11yEoVhA7f91XM+7+TytgAQ0JFPASrwOJIYJHa
AnDMNaWRA/Y/+NZsAfIa4JTX4G9xSBBIPvTn3UMjTdC1jFsFKldxw26qXH5ud6gy
PntWqGvXra3J9oYXfe2z7965ffrq8d7bgOJRm2G5ScC+XDXXFrnZaGEmGI6hOGd2
BF6aVCX0WHzGFs169ZAUBTBBqT75ViZFhFuc5W+ZfvtifWjAex295KqICjxOLwDe
NzzoGo0yFvs3QjNLPiDDX/z9ZzNwJlzKWXR4AfAi2OViqBjcOHPZGdKrDVMA67mJ
lVtgGkTfje4CMqxRKEnlJttk4hbYbrzR/AEwENc9n/diJUb1q40zTGU2C9xCLDHs
dx2TkpZVaUsvOYMv6eY3OH9Pkv1N++efxF/Hl+OxZAVZOzvuTeFjsRpyYewpF5VM
Mu8DQbBoRL2HRDqo+i5x01KRfYsesOiTY4xDpF601CboQI9lbxO1OJt1fkBAyjTW
Ge2c2FekV8vsACC4cvj7TJnn0fZfC7cjYxMfFpQbj+k5iOVryyX74IfU4uhtWwNE
jiz7dqYUhXx/wFsZrcwmn98GWb6EL0xiLI431toFarrynfmsaWsjr08mpkDzBtKN
jegk3LEjcrbs2y4FAEK3bUDwmvF3WykMSILH2R6cBPwJexLX4bDwr68J7C2fQd0Z
48A94u/USNPy+mR5H0lAU/CE0mR9FVtyWMg4hspe9i4MRDp3iTAFFcltxIHbHn6q
xYul0gvnYGb6C6kmGWW/z//aeN+tSZlX8QZSokit4ASMYBvPojtOfkI38KR8WYr5
WOF4jDg2B+GrCPjzPQ0lwmnJqHs1FlPCETSqhXLHXFNCy8oA9MRJ0zs42jJ8W+49
LYSIdvdCrlSKjJc2MeDxkA2/SWkDDlZ/3vCk8wTO4Dr/cIRkgC0vJR9WapWHRR3L
HImTScmaYO9ja5J3s7YvVjYo7dY4JXeKPuE3LCt6pgqmYFDGp3/SEaNbX7VGjTWj
vmDkKVWnij6dE3GWYiUWEHfAv9IABrYPfmHpwdi0iV5zEC5UPdabA98APYGBWGhj
UsYsyiWlhS97jIcUayxufNObHvCJt1p9eXdETGn75USislGrE5Wja8KUPXsC/Z1F
g25+O/EtWlb7+7F4DcOwHSr7d++LYEZvPkUqeKr9se10CIquviaN/X35SsAjZwFb
xgufyWQWqNqAb3wUCFGD7BVvaqmVxiwaMt+2u4NqgghYBX9rMYQ/RQuPNMU6avsn
pHHXX77TypprUfRiAVSTzl0dnOi0bgmu9J88xx/+t4jqR5YwZeG5/owjjGnM4NKM
MxVGXk0mvBXjrriXPy/TezO9Yk8vCEw6+uJfM+aW62qSipRpOfConuQ0wdoQCPr3
oxh+wXkrZamLuAuUyl/dTOXTQnMeJ55Fh+dls8GwqXuVEU4RT0yumHqXu1pZjCzA
5EDcAIYA8dmStwDFxeIKD94x7lrs7s5QW68OdxMs37FhaqXyHhHBvBptkoI3u9/o
vPP18orglEJMun5qkFgGrMZF2sdoQruFXSxe9TMR0/t9FldJU2eerqtP+LiVdopf
f4FEEN4z/eDa6iFEbl/e8mxf7q8ytcnc3NDIDC5GixWHe+1hP7ueWiYRI7BZAyj6
V73kmNMcBJ7cVDdYaNjHA83WbTeiMZTqt/HXDk/gMNIN/LR29Wo9wRTIgCH/+BP5
Ia8z00henqRTQ6hL4HqcZ3I1G8jt2PcvUQwONYAPFttPIfuOCje9YrI20GdqrSg/
0PnALzBKcRdZeY33gU9Ne3RqHoZLs/qBejvZ6/PyMVll9oagRs5bVgnKW5EFn7Nw
nxHQYVB9QX4qEbTaeY0N2zIrHg9qjAZnfok5lPWmyhEBSvQEsM2ueRblqRmF8+tp
Q953HwV9SFtnUo3H9ufZ0bEJzU2OwBhI8Fo6+a6Uo1UwtN9K13NVwPsi4O4mhBpE
h+vSdPoDL+pDck85pLE4Y04tcmC3IgTLKQ3G54aqMbzePxbqbnOanMpaXwFI1Ix6
gBNGZdjvmnDFFgI9wB0CmvZxZWu/GlgMPSa6vWSoe8kxsgPVkRRgpV3DeUu6e8fj
cVMDzTEcOtWvMuNKOxlv+uo0eHH4TTUHsmP3HQJrclzn+dN8rjlgj+D3R2624It3
wcUpg9lvMDNEb257z5gCpo52zZzjkA9tP4Ph6+O5HW7E1fxs0ibjcMrWu3fEXz8c
lWazi5bcvXp2Pj7rhG7r01O0s1l/PsxX/bic+Ev1ydSdv+kgBrhcTDss2pXy7boc
ACRgku65Ii14zqhKxHQj/NeIXpoyxXhtQ5SkcwntUMX6ctD00fEoiBvHQI0FjQcC
ylyIdZtiRtZq6vealojrNKfAN7R4roaSpDaLDK2L9y441GUXW8JsLGgoKPH3zbSp
EOsnDA9oJNwOsF5pvLAuHFOubEnzR+w5PTsljph7TF+h7mjfv4OF4OnPJ5juzewM
LhGQet2nCbrGnmg51cHjTd62m7ruQlrwQ4dY0bGLndHyeMgJIXwSbYPTNsvsWP1t
OMA/n76g1sdCcrZ40dbg35tOdr76UlnUXA5c7JlLZLud+MQChAmMn1WrMbv5Ppxb
ekA/Nfwp7Fh4+Z08dShOZvQO2u8ezedhkBcrtimSIOgUa5558MJYYf7uUtksp2Pc
9bh1Ulh6x4Rxgr8Xg+m2dLwVCA61y44M/Vf/GEP/BmZr7CsUl/qFETAcNgweAEvu
FRYDR66q9G1CTVJexyxfnEB/Bwsgzoy/Hka/tlwRyTLbIz/mlpzxHiR7OIB81qdK
5aVBu4N6PW1lgsXL1+x7mICJl9u1IeloRO9uFSlj4UVlT8+mrZx6RgLtuTa46xnv
XxjbRJ1VOz/Pc9BXRrF8uhJBT9qiCqcf9SZ42jHXHobxpA17S8jXqOKnEX/fMi7Q
XzcM3QbmKKV66N0x/LpcGV0FGFmcSGWMApizf+cfVe/Btj2LbGzcnLceaVrb2rnM
dnHW1sr4jh9wBuZIG3Arj8dMFskBSMJsh+YvTYL7AYERi6/H9vHKRMH7UsFsBl0L
j/yMCfLcJDsNOS++o+7ua3ZYqk89jyeCUYxALPMRU59UBP/Is3r6Xn2TXLwVIC47
wsmOfFypsbDcMJSYnw5YDV1RnNiK5wpUxU+XDakZ/tM3DzP+RoUayBll0vr1eTHi
kuDYYbOyxuCxUKiHxIyXMRVE2EceCa8CeJ4Jj0Usyc08DBooNNsBk8cEWRNTULKx
IRiDP3o8bRY7Mo0d5NcrU7fwgnuvdLNZBXyG1f3ylOlEUvgN010LK6SVi9n33kdn
WhpyG8rvK5aGlSMleQUf7e1aQpJMKiV0OzeffE5dI5y0+CDeIgG+ensQqG1sLWTe
dQq4VAjjaGclXTeKc0wTs9ZaQ2FJEp09IsSp7AmvDcx7Z4EPSGjuy2NIPBhNdDx/
BVjyxgKg5spaKbA85SN7cjaL9vQW3uwyuVrmnIVfM9Po+ZvCoRPP6QeNtug5v9Jr
Wa9RzvFPCEvTQ7Sri6e0FquPw8gw24F5Danno4RXYCJhA2IPEjzWI6H1m2cQt7mQ
gfkqqT0tostPjTD0fA9YWQnAU6XzFC2qHQ7zrKTr24c0RJHnE6Xf51DGVq4l4FVA
rz45uiQM3dmxOnetuQAAxxaBJiABc9CAkxw68L9Cbi8Ur/kQ/ei3C8ov7X170Clk
8s+6htY4rlKAhkKhhZfRJOAiUieMIDU6unTqRsiIff3CT8vc7K/AxGHnVRH/A4Ty
pJG8abcJXpESnYLtdfwzMY/gTfidtSHxvwa0Co7ff+UUBVPGE2YmJKQEW/gocmTb
4B72e8kzTyNaFTiZqPoZFuGH6Rq4KsLxbt3EGoWmIzbUP3bX9iCgHKeYW0C9zGSr
pTIIYWzJ6OIG1f66xPBoH9a+H6m8ng8/2tl6Bhf+wA47Cs/YFWXLS3gstG+/czNG
kXv+duTpJkERfNi9rCoZ3HCOtcKrIPmrX39Kcp+VArBqAxEG9VLqaRpvyJpvXY1S
CTjPyr4s6wjME2J0U5top17+G6IJHhIzJUNHOsoDfkMGnaJ52YoZMdW79QdQYzY4
9uecV0L8UoYxVRG1izGjsPVGffAMLiINGeI1cIK3K7Wybuff4/tAg/9pThhKu3UG
T+kPB6t36bVT7u6GDOu4+PIR/cmBfOT4kWMrslA0+UY8Bb/laeJMoJNCmhYi58fd
Tb5qJPqa2rtcbM65qUkraAiOolDt47o/FzV1Blge2Sn4PPjsc1CyDJb1HvcXodnh
0WqX2tZLHLfh72FdATRccHoafP2kdc+91JKeo/R7u6cELvtX0iRKIZzTRwI5plZ1
MoxhFBrU40BVWg7DfXNPA1taoWxlJgMNKbF5RmznIjaxUqqtspWjmZc1/i0wENae
PHFlEhwUtRobTfc087/fh2QTNBx/2Z4mU3UVBu1ZlWQKAdZtdfWNJ+9S0SW8IADg
5TFSa+gFEWXjEvPTyCymKCUaeUWb5O2CqvpGdkMLb9zj3yEgBfLVsO2iDJBXTHFu
o7P4QIydC59Gkb56dixiZqagHlbu7BU1SH1vyfsW272dHyqmQ8/kA4UlJBL/UTiy
PrUMX3NeGv9zH0ZXZcX+jGFgyELKmhQFOCKM77lU9D08aooflw1qjXMrgpuWyJsR
P/XnuT66li4slNQ6i8sDy1qDP2mUWa/b6+9VGBifTT4=
`pragma protect end_protected
