// single_region.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module single_region (
		input  wire  inclk,  //  altclkctrl_input.inclk
		output wire  outclk  // altclkctrl_output.outclk
	);

	single_region_altclkctrl_181_bjorw2i altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
