// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rNNulOy4j37AY+Y60lu2OoWv5FS1RMXfs313w9XhxyJgaa4FY6SKiDaTmhLs9uR9
jJ6sv+wOU4M7Kp6EcGoHyw3PCi6mLc+Y3FUCdCdVZBbpTjARvy+OPicGh+R6FxNg
EIYJDEDTfOiXSD/5XnLR0M0leC2msZMYg635T3rdUrY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3008)
5mKwrZzR2FMZm/XT53QDcmTtH9hOhc6SxLzC+XVWS7bEbHyAKHHrz2uV0DvbbYS1
aiGxSJL4j/U07fZ8qA2VQ+e8TEw2BkqXC12UhZ0TfI/MSMcfOE46yGhs7QR8OYGE
9mquwLjukIuz23ynyxoDzq24HRw5Bb/uBZoCNKK3Pyq83WIualfHwtlrOu16Ee7+
RveiWNN9jjH3nZfndKIsnkz0Pno5f+5+4ek1djIi14ZOCUk0TfPH49fAHKZIACpE
jNbCGel5r+l+/j03a5TnsFdIwugKyJgdZCwcXmUUr57fsgQSH8XhEf6nacUEj+S1
odz4l+FK7ydAdju167AdouZ0E3BhoqsIJaTJpKRJTl/CeOt1RZ8UVMAdCKAx77Gk
IJVxSm1PQ2XgGIgnTXxo+0/kDDYnxqwB+7sxBA6ae+P6i/E6QIKHCTuILw9yfNH2
rDBfNFx6i8oK5upDjv5aKIA0/5VhEQhk3izCF5q/HjAHqcMnU3jQZLMbYKKTK3PP
+iPgX3SAJGZw8ALON9NiZMy/V5xVbnTZNsFKhH2zmZ/KDXSKk2xQlNbhRGKGFM2i
Y9N8QdTF3Px5W4PZ3qto582jtFlCnMr10UIu+dCt96MdccpbzwB17hHHc46Ct8ZC
5UkqzsJtu94nlfYIhDmNNvpnFmCf5Ggep1tp26zL7KpvuyEqgPST5WlhK1IApdQB
PvgxDP7Ap8bNwOrQx0BEzt29UIPlyrBo7AcDogNGD6qNfoAdNi6zR79YkRAXAx5/
yOPF2ZibiRMX0ePMyHR0UqugZ7bOFlE0c+8Q/WE9LNG2bHlpxTth7bG4v7F2dG5g
Lg95w1VLDDbQeCtPuI7sEObvmjaWKdwRrvYl4s4CzJkM9vhaS4lXC8j8bZsouo5Y
xzOlrhlC1DWAj2yik+tT/EzuEWmqfaOUCyadmRwq7YHCWkpgCPixpFXNvEfTtgDM
FgTiDzaM/cjF4xw/+zJnQ0BNHwJYU0jFx/PndRfpYh/MtDrk5/RLvpdKwDiJfPMB
4LkrFMfqP2/2oaYzXBHFSpQomkK+BfgV1ztonSx72zGexQLRowSYlyJEA6VM+TyP
1ngSUemXvrNdOxi0RfH6qnEcXjXGOWO/4kHeRgblieDXn8P8bsquDYvPH9MqAonk
UbG9StiI8iJRbIG/isgBwJU4OSpzP/cPpgWbWeeng1G8bQ5AxqpOqjWAK6552aOn
s3oih2TU/jrqS2ZJI1dVVknvI8rRkip0EK6sCRyRh56FFLAE+TCyZKibjsNkciOO
6H405R8xwdLRXf0/oRDAbUjho/UmFWYb/8PjZkcjDussRhDECLRyU2zZ2a72G4t4
8/6kuF8xi1Tc4VAb9BgOoK8WNmfo4xuWI1LX9GWxyehxR/K7rxnNZXNZO8FLj4M8
libhM1As5sXDcYUdglgyqOZtmS15K8GPfexU013Njm/2/TmPcTwIDMgQWjb/+rRO
vuM+o6evjFWL/j/58UjzJhJBc81gl3PuXTcxxbBo5cdcxzjTKb8cWnHwv/47dre+
nwszXzXw7GiUVHjolW9M++x9TpPacV6cCvMwHuxEt8R49nNHVrRQAdsT0p2fFFVJ
dVaOI+V1/c1B4/HNIIRqV9QKX1sX7/UBxIJiMETEqcDScFlfDC3hKi/V+Gi1Il/n
6GR/3E1vZgN20cO9lElu/b38Lm+AwPM1DsJkmmCf3Lsc3IQfUpSABkTOjuJj60Bc
uMVQtnY9rWkO5PYP1+MclaZrtCzSrfirvRtvjdcNkZof8ElvfPiPwvTpnyoYnZNC
gmnZNDmWF1VgXZMYhw6N45iQypms9UOpJk1xJZu6ct/qX9Lp5D5h0Kue0TwH/LK+
yj3wdhJ4CUlsmjV3PtrHkIhyfiXPkrXRUVHcHyLRkCHb+bX+bFuEOEi28hcwmsI4
4JUnUnjY42wD0n15OdQET+B7i+UXCl4w9Vr/Viteg1QToVdEEb1avjAeyTxnvZKu
pCDy9TMgLCWJ1wujsDVKVAhgSTZfgNygydHpmMIdd1xTEhKhwqSARfW4ShfwDDxa
vJ2LFp3W1djN21JlTO4Z32ox9aaGnS8CO+Xj/1IZVh9OitomxYn0gOXrt1MTmqOy
zk+yXqCCOpLYrt31b9GprUEAAxaDUr3SFj3x9y4SgFWSyZjA5UZjayFPrML+STDh
EMU6fx5p6VPuWdOFHYIIwMV77IVjfMP3FIXEOv8tHSVeOcV5fR3WPTknDGtuWSnK
Zwvi1Mdref5C5WMWetM8KZfjGda6C2Rwd6pvMGAGOWI/oWujVjSIB785RzO7zRFm
Zgyq9JbeN7FURBoj4JBNpmTCsYK47yBkD8bxL01NIwYRYHvde8Bhs75acM2tNZKO
X9CRLDwIBo8trVtxQLAHGhgMRoLTX2uxD2lQAUJoTm+9tLXZ/htZv4YR1JmCMr9w
xvKhvqzRJ1V8agjIc3esCBhHd6YCp4vlSpA6uer3wrGrvmBHcRW+886wdSamRIQT
7BgxFWk29oSbuFzGlOh1sMN4N5bBUDqf6pXzQsAroBOY43ipTF3QV38WxlMVONYM
pzx5499mi4TPjM5vSFctq7kf3h26X6/IqhZ5Wmkc9Pg7ZKtv4tmJkAbVdYzYDFbC
rP5TtAfa3u0yymVrqDQixw4DNBgDCisPbDs5x4gLQoaYIVkKtWl40KAIyib7CJ5l
kpBkRzT0SfaEemce6KM0nf5IDmpVzr8wq2Z7EcYb6DC4EtWDe+cyJXvS0CJUHjjh
T1UhLV27jhmm2CWjb0IbBHCyN5cr0qk589tafE+sOqgIglzHf1wsJb3EiTctQtdz
3CCVEfVzVXtrsbRW6cSMv0icgzmAuBmHA6jTM/6LAzUbgLXZSOw5PzEP3jHOeJRV
NPZbck4a7PqM2Ggg8vNiVZcKxx0aQaazTqAT/YF5cXRAQZfNQoFc2mA4Y0qZex/v
CZjYlkFyMDG0r1WaQqb+Jz2R5b2aqjdt3m0shDxxvEQuN3ezzgl6W/xlAY7iAivH
Fgm/QHs+oW2WKYTNZ8E5ylIATteC3d8LiJV/g+5IMmj8kMUAfZRsrNOnZZUyX1Jv
UHh5wWrZGmsXjXHuVapHq2jSFlwKMJaOzLff65oGcU0BNeaD5p0NSgQCy3un4bDH
E0YAl8XUfKGloKMyBQ3wwYNtA567MumtmIp1yzXxG9ztclsWWKcwMUwVrjzv1MTh
A2XLKJhuF0xvo7NuWwxvsuGjPKLdLwkvxAr9Vju7ClfK/H8ceLglDJDMthcc4mm/
zgGiHtD791hsFPlHYHP3Dm7sABpn1IUqMt9vQk+esjg0HPFHlV1rtYQulJKWzS9N
i9QaxCzON8LC+CtTSeyoH5MCilU/zLdTP06Rkpoxbr1ZncXciyeWhkGOWRU9UNYQ
F2yJ9ZNUw58IpwShhuNRr1LXw3zHUKTGIH49pw3GPNJXpRPm2QPbxd/Ccm/gQZiF
MEldE6IKXd9CGRdNWzs5Rv6GWejuiBpKQyt1dfIFEotrIF0+h3uaobbWqWBscooU
mXz9Ycq4LoqonSOPyrAdKIw66R1Hz6X1OTm44UiZ8i9WXvYblZ23IsPyviGLOT+Y
mWctnMlB2mgMROtm71M1dzo5V3GabxvJzlSsBHYLMwrLKJLVNOeo7T1wHKU5TBHv
2q5T6B3ySlMtAxwxchdIvgZPnU6M+PPYLnkHAr/wUUEOr4VmLB909SpTzT7/02ZW
AMfkPJQ9iuP0JfJ6ExMMx3LLbVVyiDEiAfjYqQeXLWwGMuasA73hF1P5eXgXNPnx
7VhznWMNYiz5p+taXNpM+eiN6sVWwKokiS4zYOW8h3LlDZjrFU6EHShy16HIu0/H
AuQT8UsMja81w5ofYH4HJraV/M3N3viKmR1fiRemh6sdqAwYHJ0ERct0vNz+HjPn
SrHtcsO+v2MIIDxuC0aZ5tfH5j3VhXZUxnb4GgW9C+uOybZktlRP2gx2T8KPYAc+
cVq9C1/jSvYr85Q+an714qZQJdkwbAQiVp6LC7UQCL8=
`pragma protect end_protected
