// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:54 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ry2Xk32zPHCDrHC3OecMG5Y2KHWcyx2fg0t6xD/PjuvP5V9FJoFOQ6LPoH/Cmm/f
dvxuuXel70kXlNUKl1OHvqVJQpCreSpLIY14AwqpOPiPE4Iwod4DP17Ld+76PZrQ
DAFPKoqHVQaIeXJhITRFLr3J5DRsxXwAhMVHMECT2Pg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10544)
4ym2BqxMIOjdL99g/9a9I2IveAYoK4MjRjjFViTgwuilaLhv0zSxAgkdpMRIZdpe
MkClpE0nkX7uVEOdRjUHPWw+Vsgv8F0jl9Vt2v1FJqpAid2Qb08AoUq30gZ1sEDJ
ESSPTifW1L0Tlz0Kg6G9mWSYD0JxuNj32Wrx/CWf6dxSMBDbSwKhd8JDZ31Yvu3f
h/7i6seqXRnY67r6sMliKB5Pi22wTod0OG84rqYy/Gah0ZIampS+Q6gcZMArYc7C
pd8HcNJgzxuKPzd1ngtKiYoNNTKPNUtK9WJfVvkgKSycD2o9UX/pl3pfIF52qsq0
7o0eKzxSXYMAV1ji5d1Q3ywCZfLCTe6BkyFE/jzYA7jXud04eADGPG3Cz5+IwvW0
COyBeRL3YOMm98sSNPsuufoFV1DVh6Ca1Bq37hlMSGfsQNhm/obIzpIFJdaQCcB7
QR2nXsqnwLm2XFoFX8v1i+EMj11OwrDlmBUv4VcR31wCNMBNzbCjz5cTM4yij+7A
e3AXXR3hcOScMCuQI6e2pu+Q+hwKmZn8fTtbBrp2BgB8VjszPApE5wPRg3XrmUEG
+eAsChI03bVYjzIZdYNgRUevsh/hmnhoyEz2j4zmrWwI+1/0b+wGAP+6O0r9Ru1V
7OTeWKozw61XDuUvRnF0vF1X/ZK7+xx4Dm1NCSksfneP/ia2UByTtEXqwoC1xOFX
aww5VxdtOYzSsrJqWIXYDj1lDgVSzEpmFT7w9c9ozc2xs4pan8rgZL0pVKXJIkNd
KsvanFRwuv8UdCMnF6XL/9ReiZO3tNdNpI7KOZsJGbZ8kO2C9uK94SsqR6GpvNHJ
2Pdxil6hdny6Nu3gAvslDesOoJB+ocWvXPJdkasHy0/wm70dr1jiuCmBU2yjfgeQ
G1mJinb7IlTSfP1FdXWn8U09oYbwFY/Y2Bc1/GS82gWQijL3VLGB2/hoD42n4Y3e
tjpPMaaCXLvyoCMT6X0BZaAcIk6IL842hndHvEH25MZLkWQ6os3QSOc9Km5DxEji
ujgKDqxmFg/r4o4Q3/O55mLNQ4xRka38EKgU9SwAo8D/uTs1zcT4tjgXDfBjmy83
cu7j2bQxGswbJKx6Qiv3+B3LIBvA0qZB5rgt1nBqcto/hlChTopG7PLgdT+HG5Kb
nts/w3lRg35MqkJYUlZc2pkcuKpXraqKGvtjlU9o/F5gWOa1L3bZLnxPBdYe6SMo
ztAIQxcyE29qU9M6Dm5Lhg2EMbwFf1mWSNacpZHLXfG+T6Tk2eTkwYlnUI967rRh
W01PGEbF60jMuBozRsR59HbMCN9ZiukzxRqhTjp+yqmBZ5E+Ov+p55LdrpYWhLp3
+fpn1X+6kBB/7XRQObQl0+7vv1it80Mng4fgUgOPStywxvJeacd06dEVkwCOblz8
6eg+m+syyxwEpkGo58K2W8EQL7aZ5E8g+xPGfM8q3eywYttiobg0hlMy5E5Dj/go
9VB/Byz432kkKYjpdZPsm8V1oF0UT7vuTqD6bPrqx36kLRi7ddl5v3WK6P3nJlzu
+9sM9DSR622zPK7mNwMGbNyex3thX8FObu+cGb3OmSp1pNG7d0jpRzuzUwst6IPW
K2RQK33DsF2CXUXLluerYPUOxgpb3XeDxETg618nbh8Tq42L/JYs0yC9jmnbYZiW
+aoKbIVw4SsOryHPexykBhh/pW4iXWgK931m+B7Cxv+vXBe2C59MeTdZWBymu5VJ
ESjXT51LEwgsdyNd9g/USBLnIggKEoRta1sNjf+Vc5zHft51URv2va/2BanPrTgB
HD69JW/6TfW9G+IZPjCfc/ODtzsz4YfaFAajdKrxVxJFECFrMyZwFbmPSCMYtjpw
s826zgidNRBDbsp4o+5uXKyFETOaaP7wuykjTL17rIqEvcM0UjTui5koQHzU4F3F
4sVRJpWbC9DpQpKNKqe0wPhs4Oq3+XPJ07fFw0KkfORapBHGd/udcfGSyUU4s+pw
8O61NJOT2EFPxqWD0u7PNtSK9c5OF4hXG8fUwiCa+0MfCyT9c+UCdbcKMcI5nbfD
QwtmGqpgvByFxMlw8VpFJUwaSQU2FXo8CaLcRR3ic+J9FacTJtB2QU1DopQUqXic
+IEcLRy8c2KUJxVoCCN+ZhEIK0Tz0Nn5EpXQ+GG/OV22QCMCFobgN5yKyn3hPcb/
tdqlKozyLoiTAkwfhCdRRI6cOnXloEPWJBMiGdS0CevJEGFgncX3JQ+NKEH+JOsg
mz7v18sIOgshFYCZanMw7FcRcUi3cKV3hVGa3rUspAkP+Bi+zVfvIqx1nw3xa/mD
hwvupSGva5iLfwe6W5MVlZIzCCzqTTZx0YysRC+Nd7rMUk03E1r3lutJUudrVG+s
fJn/1YVmQL/TbEeD3ij6A5jjXVNDNLFuoUJS/ThgkjYYPjkWcYhM8SUHqOaaWfiP
/PNfFOhTGpxjd2CyYbM9/UUXcmxF4FAL5VZNXGVSOpyog8I2kDBitt45pBrHbIAh
2oWSpXeSiyviUYBko0WON21CLT+gw88xYb63Wt1+tCkbUHgYkmQnwM+0jRXWG3JV
OZabWYry320pWd1G+9/BO6vW/ys4YC0IkdXqcXTfVi0h7JNf+NgbTSj0zDSlv7nG
GHMi9m2Xku1d8Mso0ZDNB875x7Bdg7PHGN2OJ2/8bp/4dzKzTM2AwSVPgacFhKZK
2ztC4igSyUEjaiwZSpsYhN/67CylDoOoxkak4sGeohHaZ2727z8aKwuL0th3I7A1
hizsWAHg7zIOyaD4HkQ/UNJ2WZRd0m2BCI6EJYin1ekoCP4e5wAJTjKY8SdMqraR
nCgMyB0b+zOqEpBXLiSO7PiTA+144NNmsTeAvOQJ9ZaM46G9OiJf2SDDJdZEdiCb
cXdZ5F82OqlfO3bvNrTFbxXm9lezi/TNP3gekYAnJ+bT8tdDMvVk4Fs0nKH6Bkas
ljyUxCHpeun/mNAVZKNhNh/iEcgBzjmXubcDurJa9f7J3qemH8VUYDnyduR6OnAp
w50tmjzq9cPbbOewghuaVeRgJ7qbpVDeffg6LiPLArhVC/AHb4Krn4Mc6ChjAn/3
zfZJrntrtsWFn6JIbgTt8Wkin4hZkPqhNJ6OUtxuhsxnhSkVOvcF1g2isRZJzi+B
BM3mqjTF729pjYbmadK2SvJ4MgEkDqZxMe11Cc3V14qGIUW2MDwIk3B7YkXO+ql2
PyDtEeBHcLef606pEbSIwwYbUr+dhEr08itaTdPQAWbkb3z4Lgsg8DwCQXSKQWLZ
dlHhR2LrHhrul6jPM2RwA4DG7cuxVS1v4R3ljnO6+u7xLzMVVeVjLC/aZx/tzQMD
JxUIqThUznSqEYkONRFJHoC8gXG3KY48FdK5ZPVkVE+IQgf2HCJZPJzQloHnbHq1
eB9lSWjBy/tVcqU8u6QrbVUa4ob0cSkZCOCkR+HH6+7ZiQ7nKvozpS5aLuNjPz3s
J2dkbEtokoWeE4rsUNOZrujDEci1TCOQvHH0bZfZ2IgoG4xF4JawDnBQVHKMCjdF
mSXeEpbXva3ykMse39wzhG5nqGXDzMIP8Z7BTPsUcT5QgWWNJ8iDzP9MiRSp2l/y
zrH28uRr5k3ob7sbtc/g9COTD7psP6AFDQaRjJ410fiLW1R3iDWD+5ruBnCzlAT6
fM3HX1xWE9mXRSRFRV3s2bJYW/iyT/uXxGozSumaY7s7lrXgOWQSbN3n3K4GygSh
nM10amdUnYP2KKwh31dXNbieurOpdn4IVwCRns2gps2wpWIOHdzgmIb+4EWhh+Wj
9Nk3dvEY48D4RxnjpKjxoAsj1wUR2SrDox2jwDg2bGwUtzYaRNvPt+Q7EKmtkW8w
aciSA19gIbwrIJUpg80bYMppw8dUv/sIA+gaK+hdOYRHHHNOhjPE5Oaia6YOXyQ2
eG52GbZucBRY1OHCzc/We9ngvZwFtKBHrgE0kpvE9+QrAo979gydyYtO6RwH9MXj
kKJjIq569G6ZBkk10oGPgr/dFXT+asaA5AhpfSg4w9xJ7MZDDjrpD/A81yTQU7Um
dJLGDTjLiIUd0cco0Df9vDc2cN4V69tu+d9Z8tYuaUg9nfL3IamTwDb6NkpUIMio
7VvUgVZJWkyWc2u2lcCJhX/YI9cLzjD50hsoHspMcWWKGGvWv7d8sjLFsEh45kgT
dY+Sm6wmt2MY6M4VBkJoHFTIvjfUEaQ/k5oAv/eQiJaedsUKdBLkqvIH7M/OL0N5
M/S2xU4xY0oej1VwuepCgduKc5o6zcIoqeTMwiF8A8lh0FgKc8ZDT2IZBCHtN5uv
ULa8MfPYdCTObMky/sN8iJqPCIT5oWEBsvk7dgSr4psjUPGj3LRJhy5kY7v7QZEU
Yx7mrVIY63sWgWRAjnFrmIQZFPkgdN9ZFfnFYF9LO2yfIYUlMXU6LkOtKq7vZLK3
Dph/qkbkzZZ+hIfW3d5L6oqGkMu+DWkWWgpfjUuUx716XOyhvoWoUn2L3ut8Dblq
RVcSFwynIRWip9VH289LxdMA+RZ3/R65RWMnC8ZlqO8+mY4oVflluw5xmg+LZqk1
pvN0odYwz6tOn6kxxAipqAmKXzBIrusK4euhEWKl8z4qq+WYRYx6LULonJFx9F5G
yju4kmHX6xWTuW+aGxzyHIIb3VaFFTAs810x+qBeqRANfOrjKxXd+vJaRo6bJbVJ
54APvKrNZtzKnpZFPfcxyFlYsdGdSp/gew1U27f9SWTjhwGFH6eFd2ZKqmDy9HXb
4AwY1tivCew/DpVYdwNTrmGauQuTfGzYf8CrlTFaBcqUS7E9RMehGjYaJRbYJR5W
/4TEo9XF+UeEwxjvXDMyMRvQExqAAu5T7rN7V3peBQi2WGjDdNlqEMPwJz6fcGzB
0fmKhcHwMKifTkkhrrJ5FpMVVCl8Uj5fx3WiAYrWZTFDKdNo3dKvaTSIXElUpRx4
lu/unyYvNrEvAZZtrZ472n4/mYh+kk9FbLZzHexAVlhamW3lrBD34epC6n0YI5Sa
lOtGndWDGelyiOjXtvqI2P+5gNdbfsBZy673N8Sj2UZjlo14Nwaw3kMlZb1L0L5R
Z4+K16NIQMoMFhBysFdLEVE2R1LRbe7c5aHmEYrHV2OC0qkNQ1x+PIqh9EGpzxZG
C4mYLhnyUa/sKeeWJCN+pMXlU99JhgATffHxjqTckhyja3/G/yIA7bgkC7i3pVuV
F6XD7L+pTb/iZ22/bDaVpMCxgJhzizPI6aVLUlZaaMsdA1IpdSanTW4dk7jdU8v1
lwG0WUyhYzO0f3tUHe2/k62BRheCteifUnRUaujWjufWKTW6c/7kJqwFq2CI3R0H
+rJazLEUe1HWA1dRwmQGkpQFvM0xmnOijuL2QD7C2geQP+RCOrTexWHjWzHsaBrs
AJw4QoMp6MBV9mO43/iyy8QGabQx2PWjnX3OIjNCcOw9DGDkSJwMFUgYG07lrB6Z
hfMs2YWLdXiNMAbWAkluoAB5oq99F646gtKAD9FsRf1ijwZUcTLTW375NUrgaH5L
my8uTO0B7+sEYRK2tFOrKrrD6Ajsq7fY1BZ4gV9mrnliAmBl87K9ucLxD87/Vy8O
0YyzBc363gX7c3V8/GwUcKcQX0EtXdlQrFTQxpT9h3b1FbSYV/XOkUlzAY8dS4GU
1iUB9+WHBMxHapGm4nauUrbp6HKHEYwPNNAH1y3HQ4a6h5fP8s7vw9ptBWem2qXq
7HIGpiKB1HLeAazw0q4LImqbPNTSQehuACZvyN01K4FCd9iL2RIpP0KMaedW05oX
51NjFE1uBhwdge/ULo3stjd6FCwxC48DslBuFcXTdtADWf7qU5TdqDpMrc+Bra71
HAQJD7uiy1ovjRYjsR1NXShg/J0aV6McMOUKQXYeKFwgCWPjVOQdTwhyeu3/n19x
wfG1m7R/9grsU7mbzIJdmn2wzLVNueCOB2cY+g9Ahv3ptkDEkTkRZ2hNcMJgctyz
+C2L3y4ii6jiTU0Jr8M3dGodlRfI90Z8b6G+dmokhdOOw1MpG8fbFIIHYd+23Kii
hUGWJfuSSu7Hypbo2OBL8zGQw+EX4tYkYfNkPncE44JbYd+vhaeQbPbwc9HYTNWP
7ux4rkLBtjo/xNHZ2PQ7jN0xocRfZ5R0j7oNMhJF0famTtrU/nxnlodOE7TduBfH
3oANw2xwwhG3Uh4s56QR+MnYebylRLsNYO3OeqQHhUTJJVfuicQ9u4BtwHJWUFWM
1n0sstpA/DqZiMHWw7+zbTs+l3yaoLBKRyA13z7jX0twvRGe014y6TK6oE1+FfDO
anBBYIqz+36/iHFz14qHmEA11gmR9Kp0aLUDrLlaCtwx3vg/LbVo9tkGlMhLZMJQ
8rf1PCxcEerXeTMblXq/cFw+77ilWAKq6xKQRa4md7Z5d3bRSenB24P0Hyc0ew8/
0Ri7aL2Aj6jSRFenZ2OlzKIMVwuTDBm+VzQABCWE964TeOxUgVeRFcxtR2ahSIYi
wB+p7an5GEhd8N6rUyEFcHYkzo4AR1Zl6qggOvSPrTtdRk5PCPdspb8FW87L/1pC
q0JK+bwc/X9GUpydbh15R3jiM0EeM8LH/qhWCgQr8H3x951VpT5hnDJnGYiQ5FH6
mDxkoJJpx4XD2xvl1BtPSYfPtwArZPaYJd455wKnn0bMIXtsuR24PlH1KXDZ7TC1
kEusDbuyvABjM1L0uUr3LU8OsLTeWRbZODtO76PGmKmx7UjXN+Wg6SK5wVRSZ94y
dPvhbAu7I2UuY3F5KLbJL/863jO18QhfUxOy14itbIMDTuncToGpjkMfgjksVusX
e5wYRPZxRlLaf3vZcJZUQrTL/0aCYjCG1Z60bizdCwdxW+irXWSN9UUG4hjWO2cr
Qm0jbpigsZk/yXiQX03a6tZe5kK6pSr+vhcosBXe+ESJFZo9bhk8K0fFtTEjI0lP
g4C5Kt3WKmYyXvaWsbG7co6nj/DnQ2cWPb668/OssJp0OmZ5yJWqPzQurGt1sqhV
qZlA/tn6OfGshRkPfL6TxN6a32pcikO6kIaS61QtLx27ka1yClDxb6mVTYIbbUFJ
rTZj/krV68nfW+E2w/NWdnGPKgkWV6SLIzGPnFuhsm55fIsGxRjv4LWl/iWjNSas
nFy1hxjfw8Rm13sobNEhSCQHj/DU3TA9dHyS7De+cJBQ18i2iFbIZFkgC24VvxMb
xJ0gnhudSQJ2VXH0eqEbdQmpTcD3KpMtbptSjWNNKRYslwH8cOnRNCK+e2ePWneW
lStBvL4frfCrHGBF5VRbUrkTCfpyNwroB70NWfF9UQtUreRZz4ZR+3wA+BcAFhKi
n29nwPfaF8fTH/8iYbPyt09pNSKXJKmN/Zgz4ku1xCURjM21ZOtv2Y0FVz9Aj3hZ
VQtX169zBZbaKAMoYauaDfPMOxXCNRzPRoA3xLCP0O1RhfJW2I2sH64egNZtWDT3
vQcg0liaKf9xkn9mJX6MJQ36cZbpMOFN9xz1VStB0S+qmyl4+o+z6oSsATLpZs+P
bCBZtSGq4V2NOsEvcvJKVnYBB0zHn1+z2XSYDEsmGCxcJ+PQ8/iGvLd8OsBp9OOa
g/EO6J+4rMz7kP5sWp7z2XNugeywN4ojAcbDMbtedn/f1K2Htl5TszR3HVnrhBx7
IywDM5ygfLXz7DUFocEf8hlO2sPVi0VduWMb9vUHueuovtggCE6/EvLRRsLBl5tj
ZmijHu8nykOgUf4bas+2+t6MCsP2Pe02L4YpxQHbOssKLOszs+Oo1ZU9fvFKc0Pe
DCoX3b3fEeavPtlk3n9ARiYh1Pap2csq3THwdfWLr2xSyLTeLDxkwK9e1wPBPBaY
tabCOShuqXQwfxj2dQF6uYciTr32xzbA2kwSaUZco6YmaYrhqH2thCJqT6QZuIrY
32jbDb2tvX8PrltLcI0aElMp/Vno21kir6b04E7sLFH+EaqovL6UaMPC1+Plq7ga
Cew0Xs12d64koEDML1EEjqRDauHW+hF3wApELljtPY9lIt/8PNvcPUpJId94+XQv
i/oApKNlVHSG19GGhInPl/34mN0Ci4H60fal8LUQmH9Fn3l9GcHT1ILpELZblB/D
oimHyHwD7wr+eoLmC++LDs3k0LhcBANQGgfuqivh0hs/JTEefGnTcGLy+o7qa88y
ZES7izEWL9KXlfak/lO0mLCleIX/zW9fm03PkFz/H1eIw0oxAbbwioBqtNYBaXUx
WGDbW9zORDgfDtcQctSI8oa09lnLUVMjITnowXmclXl9r9UnbwGVr9hTbpKGB/Iv
tOTBzXr3hrlL9PkGqBjrFn8GdVgDEbUatrJOV7QSujuZy9YKrfo4pKr11f3oELK6
5SEyHweTOMYhWZSOZVyLYZmL6tgtvyut82E1QkSSKU8t1tTTpEirxbprazBogArQ
cQc8QMebSaTk3hZESmrtPMS4QKjY4tXLECL5MXaOOQ4QLXYF5xIJ+98qBT8ZukGB
cTxNDkn1+q2x62LcmxtPruSZt5tvGOT1HoC82tvg/ZJwUtV+On/PHSUKH6cfMuCL
AoKiL7q49X6SoDRCV1fxSlOUB38JaHA+1Z+Y41nmPK3SUv+C/rgxzWBVNZ/+dFsr
SYPipsxj47OIosS6793wAFtdJ2A7JqGDYh0DB5L/mkvUDDSahDnl81IJY9NGLTZE
eUznPcwI08PJ+OoYuDyZ2T7O3fLbk1mwDvduY0/glh52vjR+mOyCYtjgptGPy8Nn
EffgSoJCgyi63gtUdhLHf6RL9qd6CmqmfwZTZCDVPnqGkY6fiPK/qzrd5i7VP6cg
KU1kf0SGZfZppA/ARjnJ4Qjt2XNsvktQvxekNSzmq+EuSBTqlAB4EdvEBEJAkDll
nf+zUTmp/JZn/LWfWSMV6yH+6s9NyCAzopC8sNEd8RSP9pvIr5avvMhVQusiNV78
KEYMSlbPFlxxlQpJQaTaRkiRfQHzecaSOiKXYpcl13XKlKaKXUghL7rJ0IU984KY
z/Pjs3xiV2U6s+dFsYyA+OmzKOV8S2x1onv1XETXBJ5HCFemQhAEvqdWfgCKPaAg
8gqzXw4igtPrtcrYRPzpxTE/h3yYUdy4+QTMxYG6mpm41KIP46NADe1dFsIxvycm
zq5j1RN5kL6OGxx7eQpfNpV4/LB3pbRX7SGPcKVIUocRno12EEApAWbpPBJr4JBK
j1lJPEPrxUb/B+AYAIkArb4tpQSBdxitiIz8iNMsI5F15QRV+HDv/QdwlOjIZiQM
BctfdYGQX3BjqZCntTDUn4f+06a3IH9OQC+uGm/2pgp6O0l+jBsxpfRi359RUlww
0fMZ15WXZ8ySBlv5O/c3/sLzJi88X6ZZwR26AECdov8V5oqcUqem65yq4WE/+hWU
zSWmLSh053d631SyzNDsn3Wjn4ALQbNWuOgAGYD1orFbAgtSrVPEg08fFUUZhCUL
hUZE0ravzvDHsyn5zSFuiVDssJFoSAqhO992hrBSUD1/eXpZryLgcO5VKt0j29F+
nbzN2zsYzbDKegHQu9Y/pIRQvTlSER14xgmybCRIaqZzKMDgTurXfRW+x73VqLku
XZDT0EPmJFDyFP7lUubRE00UD+xNNGblrqW/TurcdYVpXA/Ln0O86ZlXdGmA2z7N
0eO+QTAFJrIvYBWPcUKxzRgXjJcpejzbfgI9MVA5woPyr2GtgFBgMOo4VfYDbMEV
Widyw2Buu7Uevjr9Fqd+dVPLYnhd67Gxd/cXEanNyvkKjUkkCu2gn2dS3aydbV1a
PG0M/B6hq5K7f86pJ6Lnz6ODOCjqvYXQwy996/xigW9GSCT8Qp+uCU+tQ+Xe0lIs
hsXPBWVbs4utWY8JF/HeOPYIJ/HYCL103q+xbT0yDpPBMkyBWLLhOuPPDZ2EiZ/Y
on2/aQ/Lp3W9lA0NJCJ60zMqLkOHEa9eXKvx9Uz1PEgPRSO2zn76AMJ/TMNBMTZK
pwh55MQ6Ya12dojszCXq3WchKM4HcgYT5avd6TCwxeIArbGRXtJ2Z6qPqRUbMX1g
HSv9wBRersWGVXfHLVkagXMx9dLSHrs57vLkY8slbu0SiuXNEf0z4dxO3zvWNllp
WynEMPpXPFbohiJgnEjLwQBAZlkK83BVXFTsf2NMjBMcXdRABAOpjSkr487jQYuY
Dajkh0E3ELuptstMMuHZxHuXKrapQpkUi6YX5kTiz0qUVLv7qPhKU20osOYCN9Rj
zXvNt5eZYb69mXoybJsEu9+HcmRtMJmg23w3tqXLRrKTDhHP+0G7+Ckp4hpijBeF
xeTX05i1KYBUjKKxacX+bs8GJ4rsW+ywSW7CX185x1QVPwbwISBkQcVdyStkEdIQ
BW8/gGBr/SUmARPMSFUiY1xFvu2YASR/NGXasVaDG0yC0QAYlmib+Wi0EnwKdHoG
BI6FXe8Pjxwzj1AVIv/Dx51h306HCHvybhVKJegk92Nyk1K4xUhDynD+BVS+bP+/
LJzkYOZYXLT0qMXF8nXs72FfMXX6pgueK5FgDpdady+TpRvixmo/i2mbaFvdP4Gh
FwzVkgvrsqOGW5yHKqyLIS2ZknkgzIN5PhtrNgPTOICOJXnGXszZAEtje54ZKqOm
xHP5L36CgbWozfK6occKF+fvR1bn8AeRcCuPuAskj4I4sSiUVx0zyzmF37D9vNZD
e2QQL2MmzyG2dZEZsBtGdZpgavHhw5DtcqxYByuJMQ4mNYwUCOqxxRe+vGUByH5T
D0ZVC9pyOUbD1BbenDJoctHFbwTZ2SZg4k/zx2lmLSiGbMjwRWVC3ZB/kw8obN9r
0lx6no9sVj7ULFb76fNeN1KYUZCFvG/lanriRZNijmKpNE931pmKMZeQPSwT7iLy
r9KxR4wjHeWAPdrBTDKZnAWyEBcOiOTa4PyiCYmz7FJniCwXCtrlXxUaf5yUPz55
zejGJkgdnCFjzU+Q1Fu62cFRv2FCTYmMwSsaH6S+WR+5R7H+ncEJJEyVgnE6BNGG
V7DFUqBn9NO2rwn2oNGMu2gH25G9TyjUx72McDPqfh93CMkDkCTfSWkK5VURNBhL
yMBuVqEisBGRmK/eBxW9oyNbZGXQFqmgZWpVjNmNtpX3cOgOEXWIT7GMxtNN2ZIg
VyoVQtUX7Dd+WMY2F7nwq0/2A0HqJF7lx25QdpmEZ6c3pMYQtgyb2JVffxSbutnA
Iq0P31DCvGQ+QbwwgYTNVyWsySIMqK71gRYE83TCH8Og1brn2UKZC6tduLjOabrq
yNwwUUR4rCIdR5LNARBBqyqP2u993NRzRNcuD4sVVJUmrG+5yeaPYHbH8lP+ZEfy
XQZk3uaNgiZTLNUIWh9TvaiHi0ygEBS0F0M83++tl1cNvNo7ytWU0xyptqsQjEYR
sTHtmFtMrPU9sWzcWVFcwDoFuIz4Kx32prvJnAtBLBNxqBiRf0Iid7Wd/nDLtX3K
CHTkfBYU8Q0oTkI+jilD/7L0erWyDBG/NiJuqLHTeZ6NqEx7qZFmczC2HUsYM1o4
3hvkW7I+5XP3zTSFizuA/578tsQYH48jV8MpL5N3VQn9kBRMA94DexoMvKUCe46+
3GdxKL3IUXz8b3ljSsNuXSr/nLR7Jsn1VBuIoRNy2K4z59A5mCRK4cTh6FYbA5+o
3SeHZ7nU6v/Db8oYlkO82OG8yxcDBrg7SInPp+yRFmUVMxYim9BenH/0Jl/jIr7R
7R8l9po86rfFPLiVYW3XtnPzr/0MvOvRay87tj2Ybqsg26LCL56UHsD2nGg876j+
3PpeHYHoi2ugxYeuqXK39rPfT1rBQ2pV6irzukGp9t1AmOfRtWK3FjgjBZgKOrZR
NSFxFM5sNHRPFaEap7VnQSPjHPlYKJsgmH6udGF8PNzq95YOZVDr0ESJVpCedTlw
x4LdpolcIukKDtPonHrwzQ06fkTg927UCgt3Qio97v0OmnxXzJpy8xGa9lfh5xVo
c8ETJJJlRlxpc6WDLVIJR112Fp8NBUSxgVhq7KOLVEsGdXCRVfHVMbNEsEhF86m6
Oxz9mL4V5hIkHcSd/VspSvP1nGsGjVFll15SCIZqloFZWKTBWNdy9Bd8ireRKJcj
87riUjNHZPXw2aatNUw1r2meCwqEjLyvycfnViL2LxkjaJStQPE8TrZFDRoMtVsK
QMfwHKcPLQYJHiBbrekEycjXOYHU7ABzAA76gVw2WD92Lyc2j7NIZYyNkHvJIB9j
QEDrAnXDx3D0M3zJ2FykkRhBoMZwHSeraT+H1qjZHIJQHXRlA3N0WHAKk7+nm5OA
W8I7bX4yECsR7UJWrWdfFjFHVbzQPFCAHV9J5VrrXZ2AOnrCOUSk2y1pwl/EchYv
RSP5q4b1w9HacX3C6AjbR+WYLjo+rg/884RjrGaRvN3gU4pEnl502caWZMvUezUx
XBn8soj3x65iLZ7LtaXq8lKWmIBs17MzlqI+hEViPeO+u0Hp20gSpAAQq2+OWuFX
htz27z6Zrdy+GFV92h6sNGCrgMPQ9CzYYJs1vUV1SFcQEgZlcUnnCaSR/Qa7T5Gu
DDIqRyJhK+cc1HZV7XaDeLd5NQo7Ldq4Jf0hAaD7nfk3M6LnBA4QotLq08jtcuLk
Mb7wNteZQKVa/bGOFE5dv1B6FpKpvibevoGGETn/caR0vQjehreclAJEo6MW5FKa
Mda9tFq+f28rEPk0yJSClIcsAW+69r7eOYdhNVHKCSY+Xu3Tm/TYtUwAZW4nymqP
v6d6QGgxEzvjtjgl6raqKDNPqhNXg+Ufrc+WtB7MvkJg4pP5t0bIqrWENljAzcSW
37JvyrK8WC6+TDdNGOgV6hvkIT5kN2KDMu6inEFgbF5AR7oaUrm9jGNxrnFhc3AK
FKG+IzA4bZ34AS7aaW1V+TuJdyFHLzKXb7g1nzB/PunspKXmq0KUSG/AZiwRX6g4
qFrvX9E1VDs8Ij3DndPcM/W65QbWQIJ6ru6bUIyYg+obA6zu/91THCY2mbx8/rYj
JJVJrHqPGiAS20hHd3hIbD/hhxMUhqy3f4i5nqc3OdTlNLI94pwMAlRRnVcAd+PC
uYjhq1LOh94El1Iew2Btmf71lz/4SWCGrgkNQUAXw3JfkJqcY+p6tVxJWierw/8D
X/dbFifndCPqjtJjm/gLb9vXeEbLquV8c0BR5V5dhmDR10JssFMZ3038LiNmknu4
3EFJF5TZQ+6Fa15dQEZMt43mJbFZg7Rgbu4LpxcP3jaQJLo2Rc+syqvtOq801hga
P6ccZvZhqL2p+5iOy/qQ+ElFMF5AqmLIQVwgEd5CSZttGmJFPbP7Zv1wJJTMBWLW
bI/7w1KWVWrmYBBfyijtb9vrYxXX+W1SbvXj1TQFk6x8vSSN7gBQi0bsjA71UfIA
F9cNobXG1IMG3hqmWQepe4r2TvAWJrS6HUxQidj9A7v0a5OEDrrGUZ4Pbb6wP4BF
STMw9OJFKpIjIuulb0HQhwh3eho3DfFhdsjKZHELwLIQnjz6ZezKkeyDsOw8sU6+
i5WgnygjkGZq6bRZVQgVIreJvEXmiVCRaSTVKS5++ds+K2pvBMsKxJl0lxLglo1h
dYhEpv/f+wHoWZujTN0+2yeiUK6aKl2lSitwSkfUcOFXnzoc5w8F/jdMLKY4p7hz
jh461VXsSa/wsSdrE5sxMlozeajD21SbjwtbnHhJe9ptDiW14K/JSEbHRoUBKna5
LWqw+7TTb2hlyariBay1q4Htto/K4K1T+09EHOEbrjZoipWTi0TlsSSABX+O+B/9
7TW8A/5aX+DkbpseyBK1Ya2Rw/yg0m01XhIQ273YzzmIw9Poy+J70qyxQagZ3gp9
hm6TIIFDpy5JA7DY2IGfny4MBujTkqTak0tloGv45pJgZhqTMIFNHaSkuPjjL7Ui
xf50O4MY5gkBhwa1L7R3xdz7XFpQa2j7AD69aUHCnfOzUVeAJ02NRVusr+Dn8bSx
VkbiuBiabifN3G3QQ9U83B0I2zHyOyA9msfan42/foFu/tv3gaFdYqDtLJpsEa21
s+zcTgvEfKRUUDRar5d3FSrNCx+3RWNm3PmHjT05UL4ych9w1p2L2H+OKitrxNqZ
T5TxDZvzo4yb+lqf2ynK0eaH3cGvqxbzs8J0ZJkrDvo=
`pragma protect end_protected
